# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfstp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.935000 2.255000 2.155000 ;
        RECT 0.720000 1.870000 2.255000 1.935000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.070000 1.765000 15.685000 1.935000 ;
        RECT 14.070000 1.935000 14.300000 3.075000 ;
        RECT 14.080000 0.255000 14.270000 1.075000 ;
        RECT 14.080000 1.075000 15.685000 1.255000 ;
        RECT 14.940000 0.255000 15.130000 1.075000 ;
        RECT 14.970000 1.935000 15.160000 3.075000 ;
        RECT 15.035000 1.255000 15.685000 1.765000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.140000 0.550000 1.765000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435000 0.390000 3.695000 1.760000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.305000 0.255000 10.855000 0.665000 ;
        RECT 10.685000 0.665000 10.855000 1.585000 ;
        RECT 10.685000 1.585000 11.895000 1.765000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.205000 0.830000 4.780000 1.775000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.840000 0.085000 ;
        RECT  0.275000  0.085000  0.605000 0.970000 ;
        RECT  1.855000  0.085000  2.185000 0.970000 ;
        RECT  4.410000  0.085000  4.660000 0.660000 ;
        RECT  6.910000  0.085000  7.240000 0.780000 ;
        RECT  7.965000  0.085000  8.135000 0.835000 ;
        RECT  7.965000  0.835000  9.315000 1.185000 ;
        RECT 11.745000  0.085000 12.075000 1.005000 ;
        RECT 13.580000  0.085000 13.910000 1.130000 ;
        RECT 14.440000  0.085000 14.770000 0.905000 ;
        RECT 15.300000  0.085000 15.630000 0.905000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 15.840000 3.415000 ;
        RECT  0.525000 2.665000  0.855000 3.245000 ;
        RECT  2.645000 2.725000  2.855000 3.245000 ;
        RECT  4.350000 2.795000  4.610000 3.245000 ;
        RECT  6.890000 2.435000  7.080000 3.245000 ;
        RECT  8.300000 2.135000  8.630000 3.245000 ;
        RECT 11.340000 2.630000 11.550000 3.245000 ;
        RECT 12.230000 2.460000 12.525000 3.245000 ;
        RECT 13.650000 1.815000 13.900000 3.245000 ;
        RECT 14.470000 2.105000 14.800000 3.245000 ;
        RECT 15.330000 2.105000 15.660000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.095000 2.325000  2.135000 2.495000 ;
      RECT  0.095000 2.495000  0.355000 3.045000 ;
      RECT  1.065000 0.640000  1.395000 1.215000 ;
      RECT  1.065000 1.215000  2.595000 1.540000 ;
      RECT  1.370000 2.665000  1.700000 2.905000 ;
      RECT  1.370000 2.905000  2.475000 3.075000 ;
      RECT  1.870000 2.495000  2.135000 2.735000 ;
      RECT  2.305000 2.385000  3.195000 2.555000 ;
      RECT  2.305000 2.555000  2.475000 2.905000 ;
      RECT  2.355000 0.640000  3.025000 0.970000 ;
      RECT  2.425000 1.540000  2.595000 2.385000 ;
      RECT  2.765000 0.970000  3.025000 1.930000 ;
      RECT  2.765000 1.930000  3.625000 2.100000 ;
      RECT  3.025000 2.555000  3.195000 2.905000 ;
      RECT  3.025000 2.905000  4.180000 3.075000 ;
      RECT  3.365000 2.100000  3.625000 2.735000 ;
      RECT  3.825000 2.025000  4.985000 2.285000 ;
      RECT  3.865000 0.330000  4.240000 0.660000 ;
      RECT  3.865000 0.660000  4.035000 1.945000 ;
      RECT  3.865000 1.945000  4.985000 2.025000 ;
      RECT  3.955000 2.455000  5.590000 2.625000 ;
      RECT  3.955000 2.625000  4.180000 2.905000 ;
      RECT  4.780000 2.795000  5.930000 2.805000 ;
      RECT  4.780000 2.805000  6.720000 3.075000 ;
      RECT  4.830000 0.255000  6.020000 0.425000 ;
      RECT  4.830000 0.425000  5.070000 0.660000 ;
      RECT  5.340000 0.595000  5.680000 0.805000 ;
      RECT  5.340000 0.805000  5.590000 2.455000 ;
      RECT  5.760000 1.295000  6.020000 1.965000 ;
      RECT  5.760000 1.965000  5.930000 2.795000 ;
      RECT  5.850000 0.425000  6.020000 1.295000 ;
      RECT  6.100000 2.305000  6.370000 2.635000 ;
      RECT  6.190000 0.535000  6.450000 0.865000 ;
      RECT  6.190000 0.865000  6.370000 1.355000 ;
      RECT  6.190000 1.355000  8.935000 1.545000 ;
      RECT  6.190000 1.545000  6.370000 2.305000 ;
      RECT  6.540000 2.095000  7.420000 2.265000 ;
      RECT  6.540000 2.265000  6.720000 2.805000 ;
      RECT  6.695000 1.715000  7.780000 1.925000 ;
      RECT  6.785000 0.950000  7.785000 1.185000 ;
      RECT  7.250000 2.265000  7.420000 2.785000 ;
      RECT  7.250000 2.785000  8.120000 2.955000 ;
      RECT  7.590000 1.925000  7.780000 2.615000 ;
      RECT  7.595000 0.735000  7.785000 0.950000 ;
      RECT  7.950000 1.795000  9.690000 1.965000 ;
      RECT  7.950000 1.965000  8.120000 2.785000 ;
      RECT  8.605000 1.545000  8.935000 1.625000 ;
      RECT  8.800000 2.295000 10.630000 2.475000 ;
      RECT  8.800000 2.475000  9.000000 2.635000 ;
      RECT  9.250000 2.645000  9.580000 2.695000 ;
      RECT  9.250000 2.695000 11.120000 3.025000 ;
      RECT  9.360000 1.965000  9.690000 2.015000 ;
      RECT  9.870000 0.835000 10.515000 1.935000 ;
      RECT  9.870000 1.935000 12.465000 2.125000 ;
      RECT 10.300000 2.475000 10.630000 2.525000 ;
      RECT 11.025000 1.175000 12.560000 1.235000 ;
      RECT 11.025000 1.235000 12.990000 1.415000 ;
      RECT 11.770000 2.125000 12.465000 2.255000 ;
      RECT 11.770000 2.255000 12.060000 2.960000 ;
      RECT 12.110000 1.585000 12.465000 1.935000 ;
      RECT 12.265000 0.675000 12.560000 1.175000 ;
      RECT 12.695000 1.415000 12.990000 2.790000 ;
      RECT 13.160000 0.255000 13.410000 1.425000 ;
      RECT 13.160000 1.425000 14.855000 1.595000 ;
      RECT 13.160000 1.595000 13.480000 3.075000 ;
  END
END sky130_fd_sc_lp__sdfstp_4
