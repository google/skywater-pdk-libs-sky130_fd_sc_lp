* NGSPICE file created from sky130_fd_sc_lp__nand3b_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand3b_m A_N B C VGND VNB VPB VPWR Y
M1000 VPWR A_N a_37_47# VPB phighvt w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=1.113e+11p ps=1.37e+06u
M1001 VGND A_N a_37_47# VNB nshort w=420000u l=150000u
+  ad=2.121e+11p pd=1.85e+06u as=1.113e+11p ps=1.37e+06u
M1002 Y C VPWR VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1003 Y a_37_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_323_47# B a_251_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1005 Y a_37_47# a_323_47# VNB nshort w=420000u l=150000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1006 VPWR B Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_251_47# C VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

