* File: sky130_fd_sc_lp__nand4_1.spice
* Created: Wed Sep  2 10:05:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4_1.pex.spice"
.subckt sky130_fd_sc_lp__nand4_1  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1007 A_133_47# N_D_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2226 PD=1.08 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1003 A_211_47# N_C_M1003_g A_133_47# VNB NSHORT L=0.15 W=0.84 AD=0.1764
+ AS=0.1008 PD=1.26 PS=1.08 NRD=22.14 NRS=9.276 M=1 R=5.6 SA=75000.6 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1000 A_325_47# N_B_M1000_g A_211_47# VNB NSHORT L=0.15 W=0.84 AD=0.1764
+ AS=0.1764 PD=1.26 PS=1.26 NRD=22.14 NRS=22.14 M=1 R=5.6 SA=75001.1 SB=75001
+ A=0.126 P=1.98 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g A_325_47# VNB NSHORT L=0.15 W=0.84 AD=0.4284
+ AS=0.1764 PD=2.7 PS=1.26 NRD=34.992 NRS=22.14 M=1 R=5.6 SA=75001.7 SB=75000.4
+ A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3654 PD=1.54 PS=3.1 NRD=0 NRS=3.9006 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3276 AS=0.1764 PD=1.78 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3276 PD=1.54 PS=1.78 NRD=0 NRS=37.5088 M=1 R=8.4 SA=75001.3
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.5796 AS=0.1764 PD=3.44 PS=1.54 NRD=30.4759 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75000.4 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__nand4_1.pxi.spice"
*
.ends
*
*
