* File: sky130_fd_sc_lp__o21a_4.pex.spice
* Created: Fri Aug 28 11:04:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21A_4%A_90_23# 1 2 3 12 16 20 24 28 32 36 40 42 51
+ 53 54 55 56 57 58 60 64 66 69 70 72 74 77 88
c153 72 0 1.8044e-19 $X=4.53 $Y=2.035
c154 66 0 8.01629e-20 $X=4.085 $Y=1.16
r155 85 86 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.705 $Y=1.49
+ $X2=1.815 $Y2=1.49
r156 84 85 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.385 $Y=1.49
+ $X2=1.705 $Y2=1.49
r157 83 84 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.275 $Y=1.49
+ $X2=1.385 $Y2=1.49
r158 82 83 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=0.955 $Y=1.49
+ $X2=1.275 $Y2=1.49
r159 81 82 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.845 $Y=1.49
+ $X2=0.955 $Y2=1.49
r160 70 72 13.9957 $w=2.08e-07 $l=2.65e-07 $layer=LI1_cond $X=4.265 $Y=2.035
+ $X2=4.53 $Y2=2.035
r161 69 70 6.86909 $w=2.1e-07 $l=1.43091e-07 $layer=LI1_cond $X=4.175 $Y=1.93
+ $X2=4.265 $Y2=2.035
r162 68 69 42.2071 $w=1.78e-07 $l=6.85e-07 $layer=LI1_cond $X=4.175 $Y=1.245
+ $X2=4.175 $Y2=1.93
r163 67 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=1.16
+ $X2=3.08 $Y2=1.16
r164 66 68 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.085 $Y=1.16
+ $X2=4.175 $Y2=1.245
r165 66 67 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.085 $Y=1.16
+ $X2=3.245 $Y2=1.16
r166 62 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.075
+ $X2=3.08 $Y2=1.16
r167 62 64 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.08 $Y=1.075
+ $X2=3.08 $Y2=0.68
r168 58 76 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.1 $X2=2.78
+ $Y2=2.015
r169 58 60 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=2.78 $Y=2.1
+ $X2=2.78 $Y2=2.91
r170 56 76 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.685 $Y=2.015
+ $X2=2.78 $Y2=2.015
r171 56 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.685 $Y=2.015
+ $X2=2.345 $Y2=2.015
r172 54 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=1.16
+ $X2=3.08 $Y2=1.16
r173 54 55 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.915 $Y=1.16
+ $X2=2.345 $Y2=1.16
r174 53 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.26 $Y=1.93
+ $X2=2.345 $Y2=2.015
r175 52 74 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.26 $Y=1.585
+ $X2=2.26 $Y2=1.49
r176 52 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.26 $Y=1.585
+ $X2=2.26 $Y2=1.93
r177 51 74 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.26 $Y=1.395
+ $X2=2.26 $Y2=1.49
r178 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.26 $Y=1.245
+ $X2=2.345 $Y2=1.16
r179 50 51 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.26 $Y=1.245
+ $X2=2.26 $Y2=1.395
r180 49 88 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.045 $Y=1.49
+ $X2=2.135 $Y2=1.49
r181 49 86 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.045 $Y=1.49
+ $X2=1.815 $Y2=1.49
r182 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.045
+ $Y=1.49 $X2=2.045 $Y2=1.49
r183 45 81 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.685 $Y=1.49
+ $X2=0.845 $Y2=1.49
r184 45 78 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.685 $Y=1.49
+ $X2=0.525 $Y2=1.49
r185 44 48 79.3876 $w=1.88e-07 $l=1.36e-06 $layer=LI1_cond $X=0.685 $Y=1.49
+ $X2=2.045 $Y2=1.49
r186 44 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.685
+ $Y=1.49 $X2=0.685 $Y2=1.49
r187 42 74 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=1.49
+ $X2=2.26 $Y2=1.49
r188 42 48 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.175 $Y=1.49
+ $X2=2.045 $Y2=1.49
r189 38 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.655
+ $X2=2.135 $Y2=1.49
r190 38 40 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.135 $Y=1.655
+ $X2=2.135 $Y2=2.465
r191 34 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.49
r192 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=0.665
r193 30 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.655
+ $X2=1.705 $Y2=1.49
r194 30 32 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.705 $Y=1.655
+ $X2=1.705 $Y2=2.465
r195 26 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.49
r196 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=0.665
r197 22 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.275 $Y=1.655
+ $X2=1.275 $Y2=1.49
r198 22 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.275 $Y=1.655
+ $X2=1.275 $Y2=2.465
r199 18 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.49
r200 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=0.665
r201 14 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.845 $Y=1.655
+ $X2=0.845 $Y2=1.49
r202 14 16 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.845 $Y=1.655
+ $X2=0.845 $Y2=2.465
r203 10 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.49
r204 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=0.665
r205 3 72 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.835 $X2=4.53 $Y2=2.035
r206 2 76 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=1.835 $X2=2.78 $Y2=2.095
r207 2 60 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=1.835 $X2=2.78 $Y2=2.91
r208 1 64 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.325 $X2=3.08 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%B1 3 7 11 15 17 28 29
r56 27 29 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=3.02 $Y=1.51
+ $X2=3.295 $Y2=1.51
r57 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.51 $X2=3.02 $Y2=1.51
r58 25 27 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.995 $Y=1.51
+ $X2=3.02 $Y2=1.51
r59 24 25 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.865 $Y=1.51
+ $X2=2.995 $Y2=1.51
r60 23 28 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.68 $Y=1.592
+ $X2=3.02 $Y2=1.592
r61 22 24 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.68 $Y=1.51
+ $X2=2.865 $Y2=1.51
r62 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.51 $X2=2.68 $Y2=1.51
r63 19 22 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.565 $Y=1.51
+ $X2=2.68 $Y2=1.51
r64 17 23 1.37605 $w=3.33e-07 $l=4e-08 $layer=LI1_cond $X=2.64 $Y=1.592 $X2=2.68
+ $Y2=1.592
r65 13 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.345
+ $X2=3.295 $Y2=1.51
r66 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.295 $Y=1.345
+ $X2=3.295 $Y2=0.745
r67 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.995 $Y=1.675
+ $X2=2.995 $Y2=1.51
r68 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.995 $Y=1.675
+ $X2=2.995 $Y2=2.465
r69 5 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.345
+ $X2=2.865 $Y2=1.51
r70 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.865 $Y=1.345 $X2=2.865
+ $Y2=0.745
r71 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.565 $Y=1.675
+ $X2=2.565 $Y2=1.51
r72 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.565 $Y=1.675
+ $X2=2.565 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%A1 3 7 11 15 18 20 21 23 24 27 28 31 32 33 34
c88 20 0 5.42069e-20 $X=5.04 $Y=2.31
c89 15 0 1.8044e-19 $X=5.175 $Y=2.465
r90 33 34 15.2014 $w=3.58e-07 $l=3.95e-07 $layer=LI1_cond $X=4.56 $Y=2.405
+ $X2=4.955 $Y2=2.405
r91 32 33 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=2.405
+ $X2=4.56 $Y2=2.405
r92 31 32 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=2.405
+ $X2=4.08 $Y2=2.405
r93 28 41 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.772 $Y=1.51
+ $X2=3.772 $Y2=1.675
r94 28 40 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.772 $Y=1.51
+ $X2=3.772 $Y2=1.345
r95 27 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.75 $Y=1.51
+ $X2=3.75 $Y2=1.675
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.75
+ $Y=1.51 $X2=3.75 $Y2=1.51
r97 24 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.51
+ $X2=5.265 $Y2=1.675
r98 24 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.51
+ $X2=5.265 $Y2=1.345
r99 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.265
+ $Y=1.51 $X2=5.265 $Y2=1.51
r100 21 23 7.33373 $w=2.18e-07 $l=1.4e-07 $layer=LI1_cond $X=5.125 $Y=1.535
+ $X2=5.265 $Y2=1.535
r101 20 34 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.04 $Y=2.31
+ $X2=5.04 $Y2=2.405
r102 19 21 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.04 $Y=1.645
+ $X2=5.125 $Y2=1.535
r103 19 20 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.04 $Y=1.645
+ $X2=5.04 $Y2=2.31
r104 18 31 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.83 $Y=2.31
+ $X2=3.915 $Y2=2.405
r105 18 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.83 $Y=2.31
+ $X2=3.83 $Y2=1.675
r106 15 44 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.175 $Y=2.465
+ $X2=5.175 $Y2=1.675
r107 11 43 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.175 $Y=0.745
+ $X2=5.175 $Y2=1.345
r108 7 41 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.885 $Y=2.465
+ $X2=3.885 $Y2=1.675
r109 3 40 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.805 $Y=0.745
+ $X2=3.805 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%A2 3 7 11 15 17 23 24
c59 11 0 8.01629e-20 $X=4.745 $Y=0.745
c60 3 0 7.08164e-20 $X=4.315 $Y=0.745
r61 22 24 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.61 $Y=1.51
+ $X2=4.745 $Y2=1.51
r62 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.61
+ $Y=1.51 $X2=4.61 $Y2=1.51
r63 19 22 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=4.315 $Y=1.51
+ $X2=4.61 $Y2=1.51
r64 17 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.61 $Y=1.665
+ $X2=4.61 $Y2=1.51
r65 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.675
+ $X2=4.745 $Y2=1.51
r66 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.745 $Y=1.675
+ $X2=4.745 $Y2=2.465
r67 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.345
+ $X2=4.745 $Y2=1.51
r68 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.745 $Y=1.345 $X2=4.745
+ $Y2=0.745
r69 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.675
+ $X2=4.315 $Y2=1.51
r70 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.315 $Y=1.675
+ $X2=4.315 $Y2=2.465
r71 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.345
+ $X2=4.315 $Y2=1.51
r72 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.315 $Y=1.345 $X2=4.315
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%VPWR 1 2 3 4 5 18 24 30 36 38 40 45 46 48 49
+ 50 51 52 64 75 82 85
r89 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 81 82 9.82912 $w=6.08e-07 $l=1.45e-07 $layer=LI1_cond $X=3.67 $Y=3.11
+ $X2=3.815 $Y2=3.11
r91 78 81 1.37255 $w=6.08e-07 $l=7e-08 $layer=LI1_cond $X=3.6 $Y=3.11 $X2=3.67
+ $Y2=3.11
r92 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r93 76 78 3.72549 $w=6.08e-07 $l=1.9e-07 $layer=LI1_cond $X=3.41 $Y=3.11 $X2=3.6
+ $Y2=3.11
r94 74 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r95 73 76 5.68627 $w=6.08e-07 $l=2.9e-07 $layer=LI1_cond $X=3.12 $Y=3.11
+ $X2=3.41 $Y2=3.11
r96 73 75 8.45657 $w=6.08e-07 $l=7.5e-08 $layer=LI1_cond $X=3.12 $Y=3.11
+ $X2=3.045 $Y2=3.11
r97 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 71 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r99 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 68 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r102 67 70 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 67 82 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.815 $Y2=3.33
r104 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r105 64 84 3.9934 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=5.295 $Y=3.33
+ $X2=5.527 $Y2=3.33
r106 64 70 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.295 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 56 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r112 52 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 52 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r114 50 62 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.35 $Y2=3.33
r116 48 59 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.49 $Y2=3.33
r118 47 62 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.655 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=3.33
+ $X2=1.49 $Y2=3.33
r120 45 55 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.24 $Y2=3.33
r121 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.63 $Y2=3.33
r122 44 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.63 $Y2=3.33
r124 40 43 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=5.425 $Y=1.98
+ $X2=5.425 $Y2=2.95
r125 38 84 3.21882 $w=2.6e-07 $l=1.38109e-07 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.527 $Y2=3.33
r126 38 43 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.425 $Y2=2.95
r127 34 76 4.33422 $w=3.3e-07 $l=3.05e-07 $layer=LI1_cond $X=3.41 $Y=2.805
+ $X2=3.41 $Y2=3.11
r128 34 36 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=3.41 $Y=2.805
+ $X2=3.41 $Y2=2.01
r129 33 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.35 $Y2=3.33
r130 33 75 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=3.045 $Y2=3.33
r131 28 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=3.245
+ $X2=2.35 $Y2=3.33
r132 28 30 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=2.35 $Y=3.245
+ $X2=2.35 $Y2=2.38
r133 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.49 $Y=2.18
+ $X2=1.49 $Y2=2.95
r134 22 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=3.245
+ $X2=1.49 $Y2=3.33
r135 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.49 $Y=3.245
+ $X2=1.49 $Y2=2.95
r136 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.63 $Y=2.18
+ $X2=0.63 $Y2=2.95
r137 16 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=3.245
+ $X2=0.63 $Y2=3.33
r138 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.63 $Y=3.245
+ $X2=0.63 $Y2=2.95
r139 5 43 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.835 $X2=5.39 $Y2=2.95
r140 5 40 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.835 $X2=5.39 $Y2=1.98
r141 4 81 300 $w=1.7e-07 $l=1.40329e-06 $layer=licon1_PDIFF $count=2 $X=3.07
+ $Y=1.835 $X2=3.67 $Y2=2.97
r142 4 36 300 $w=1.7e-07 $l=4.1845e-07 $layer=licon1_PDIFF $count=2 $X=3.07
+ $Y=1.835 $X2=3.41 $Y2=2.01
r143 3 30 300 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=2 $X=2.21
+ $Y=1.835 $X2=2.35 $Y2=2.38
r144 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.35
+ $Y=1.835 $X2=1.49 $Y2=2.95
r145 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.35
+ $Y=1.835 $X2=1.49 $Y2=2.18
r146 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.505
+ $Y=1.835 $X2=0.63 $Y2=2.95
r147 1 18 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.505
+ $Y=1.835 $X2=0.63 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%X 1 2 3 4 13 15 16 19 21 25 29 33 37 42 43 44
+ 45 49 51
r56 49 51 3.04419 $w=2.63e-07 $l=7e-08 $layer=LI1_cond $X=0.217 $Y=1.225
+ $X2=0.217 $Y2=1.295
r57 44 49 2.82608 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=1.14
+ $X2=0.217 $Y2=1.225
r58 44 45 15.7863 $w=2.63e-07 $l=3.63e-07 $layer=LI1_cond $X=0.217 $Y=1.302
+ $X2=0.217 $Y2=1.665
r59 44 51 0.304419 $w=2.63e-07 $l=7e-09 $layer=LI1_cond $X=0.217 $Y=1.302
+ $X2=0.217 $Y2=1.295
r60 41 45 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=0.217 $Y=1.755
+ $X2=0.217 $Y2=1.665
r61 37 39 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=1.915 $Y=1.98
+ $X2=1.915 $Y2=2.91
r62 35 37 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.915 $Y=1.925
+ $X2=1.915 $Y2=1.98
r63 31 33 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=1.6 $Y=1.055 $X2=1.6
+ $Y2=0.42
r64 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.155 $Y=1.84
+ $X2=1.06 $Y2=1.84
r65 29 35 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.825 $Y=1.84
+ $X2=1.915 $Y2=1.925
r66 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.825 $Y=1.84
+ $X2=1.155 $Y2=1.84
r67 25 27 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.06 $Y=1.98
+ $X2=1.06 $Y2=2.91
r68 23 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=1.925
+ $X2=1.06 $Y2=1.84
r69 23 25 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.06 $Y=1.925
+ $X2=1.06 $Y2=1.98
r70 22 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.835 $Y=1.14
+ $X2=0.74 $Y2=1.14
r71 21 31 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.505 $Y=1.14
+ $X2=1.6 $Y2=1.055
r72 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.505 $Y=1.14
+ $X2=0.835 $Y2=1.14
r73 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=1.055
+ $X2=0.74 $Y2=1.14
r74 17 19 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.74 $Y=1.055
+ $X2=0.74 $Y2=0.42
r75 16 41 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.35 $Y=1.84
+ $X2=0.217 $Y2=1.755
r76 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.965 $Y=1.84
+ $X2=1.06 $Y2=1.84
r77 15 16 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.965 $Y=1.84
+ $X2=0.35 $Y2=1.84
r78 14 44 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.35 $Y=1.14
+ $X2=0.217 $Y2=1.14
r79 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.645 $Y=1.14
+ $X2=0.74 $Y2=1.14
r80 13 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.645 $Y=1.14
+ $X2=0.35 $Y2=1.14
r81 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.78
+ $Y=1.835 $X2=1.92 $Y2=2.91
r82 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.78
+ $Y=1.835 $X2=1.92 $Y2=1.98
r83 3 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.92
+ $Y=1.835 $X2=1.06 $Y2=2.91
r84 3 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.92
+ $Y=1.835 $X2=1.06 $Y2=1.98
r85 2 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.46
+ $Y=0.245 $X2=1.6 $Y2=0.42
r86 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.245 $X2=0.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%A_792_367# 1 2 11
r14 8 11 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.1 $Y=2.835 $X2=4.96
+ $Y2=2.835
r15 2 11 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=2.835
r16 1 8 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.835 $X2=4.1 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 60 61 67 70 73 76
r88 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r89 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r90 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r91 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r93 61 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r94 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r95 58 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=4.96
+ $Y2=0
r96 58 60 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=5.52
+ $Y2=0
r97 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r98 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r99 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r100 54 73 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.095
+ $Y2=0
r101 54 56 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.56
+ $Y2=0
r102 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.96
+ $Y2=0
r103 53 56 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=4.56 $Y2=0
r104 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r105 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r106 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.03
+ $Y2=0
r107 49 51 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.195 $Y=0
+ $X2=3.6 $Y2=0
r108 48 73 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.095
+ $Y2=0
r109 48 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.6
+ $Y2=0
r110 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r111 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r112 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r113 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.17
+ $Y2=0
r114 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.68
+ $Y2=0
r115 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.03
+ $Y2=0
r116 43 46 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.68 $Y2=0
r117 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r118 42 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r119 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r120 39 64 4.66755 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=0
+ $X2=0.237 $Y2=0
r121 39 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.475 $Y=0 $X2=0.72
+ $Y2=0
r122 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.17
+ $Y2=0
r123 38 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0
+ $X2=0.72 $Y2=0
r124 36 52 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r125 36 71 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r126 32 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r127 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.45
r128 28 73 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.095 $Y=0.085
+ $X2=4.095 $Y2=0
r129 28 30 12.3718 $w=3.38e-07 $l=3.65e-07 $layer=LI1_cond $X=4.095 $Y=0.085
+ $X2=4.095 $Y2=0.45
r130 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r131 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.39
r132 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r133 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.37
r134 16 64 3.09863 $w=3.3e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.237 $Y2=0
r135 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.31 $Y2=0.39
r136 5 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.82
+ $Y=0.325 $X2=4.96 $Y2=0.45
r137 4 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.88
+ $Y=0.325 $X2=4.09 $Y2=0.45
r138 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.89
+ $Y=0.245 $X2=2.03 $Y2=0.39
r139 2 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.245 $X2=1.17 $Y2=0.37
r140 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.185
+ $Y=0.245 $X2=0.31 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_4%A_485_65# 1 2 3 4 15 17 18 22 23 24 27 33 34
+ 37
c61 17 0 7.08164e-20 $X=3.425 $Y=0.34
r62 35 37 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=5.425 $Y=1.085
+ $X2=5.425 $Y2=0.47
r63 33 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.295 $Y=1.17
+ $X2=5.425 $Y2=1.085
r64 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=1.17
+ $X2=4.625 $Y2=1.17
r65 30 34 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.53 $Y=1.085
+ $X2=4.625 $Y2=1.17
r66 30 32 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=4.53 $Y=1.085
+ $X2=4.53 $Y2=1.02
r67 29 39 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.905
+ $X2=4.53 $Y2=0.82
r68 29 32 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=4.53 $Y=0.905
+ $X2=4.53 $Y2=1.02
r69 25 39 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.735
+ $X2=4.53 $Y2=0.82
r70 25 27 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=4.53 $Y=0.735
+ $X2=4.53 $Y2=0.47
r71 23 39 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.435 $Y=0.82
+ $X2=4.53 $Y2=0.82
r72 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.435 $Y=0.82
+ $X2=3.755 $Y2=0.82
r73 20 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.59 $Y=0.735
+ $X2=3.755 $Y2=0.82
r74 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.59 $Y=0.735
+ $X2=3.59 $Y2=0.45
r75 19 22 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.59 $Y=0.425
+ $X2=3.59 $Y2=0.45
r76 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.425 $Y=0.34
+ $X2=3.59 $Y2=0.425
r77 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.425 $Y=0.34
+ $X2=2.745 $Y2=0.34
r78 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.58 $Y=0.425
+ $X2=2.745 $Y2=0.34
r79 13 15 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.58 $Y=0.425
+ $X2=2.58 $Y2=0.45
r80 4 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.25
+ $Y=0.325 $X2=5.39 $Y2=0.47
r81 3 32 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.325 $X2=4.53 $Y2=1.02
r82 3 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.325 $X2=4.53 $Y2=0.47
r83 2 22 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=3.37
+ $Y=0.325 $X2=3.59 $Y2=0.45
r84 1 15 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=2.425
+ $Y=0.325 $X2=2.58 $Y2=0.45
.ends

