* File: sky130_fd_sc_lp__a21bo_4.pex.spice
* Created: Wed Sep  2 09:18:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BO_4%B1_N 3 7 9 10 14
r36 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.375
+ $X2=0.535 $Y2=1.54
r37 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.375
+ $X2=0.535 $Y2=1.21
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.375 $X2=0.535 $Y2=1.375
r39 10 15 9.1564 $w=3.63e-07 $l=2.9e-07 $layer=LI1_cond $X=0.622 $Y=1.665
+ $X2=0.622 $Y2=1.375
r40 9 15 2.5259 $w=3.63e-07 $l=8e-08 $layer=LI1_cond $X=0.622 $Y=1.295 $X2=0.622
+ $Y2=1.375
r41 7 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.585 $Y=2.465
+ $X2=0.585 $Y2=1.54
r42 3 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.55 $Y=0.655
+ $X2=0.55 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%A_188_315# 1 2 3 10 12 13 14 17 19 21 24 28
+ 32 36 40 42 49 51 52 53 56 62 64 68 70
c146 51 0 6.74193e-20 $X=2.735 $Y=1.355
r147 71 72 17.1165 $w=3.52e-07 $l=1.25e-07 $layer=POLY_cond $X=1.32 $Y=1.5
+ $X2=1.445 $Y2=1.5
r148 66 68 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.115 $Y=0.995
+ $X2=5.115 $Y2=0.76
r149 65 70 4.43451 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=1.08
+ $X2=3.78 $Y2=1.08
r150 64 66 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.015 $Y=1.08
+ $X2=5.115 $Y2=0.995
r151 64 65 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=5.015 $Y=1.08
+ $X2=3.945 $Y2=1.08
r152 60 70 1.86336 $w=1.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.74 $Y=0.995
+ $X2=3.78 $Y2=1.08
r153 60 62 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=3.74 $Y=0.995
+ $X2=3.74 $Y2=0.42
r154 56 58 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.78 $Y=1.97
+ $X2=3.78 $Y2=2.65
r155 54 70 1.86336 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=1.165
+ $X2=3.78 $Y2=1.08
r156 54 56 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=3.78 $Y=1.165
+ $X2=3.78 $Y2=1.97
r157 52 70 4.43451 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=1.08
+ $X2=3.78 $Y2=1.08
r158 52 53 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=3.615 $Y=1.08
+ $X2=2.82 $Y2=1.08
r159 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.735 $Y=1.165
+ $X2=2.82 $Y2=1.08
r160 50 51 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.735 $Y=1.165
+ $X2=2.735 $Y2=1.355
r161 49 79 12.3239 $w=3.52e-07 $l=9e-08 $layer=POLY_cond $X=2.53 $Y=1.5 $X2=2.62
+ $Y2=1.5
r162 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.53
+ $Y=1.44 $X2=2.53 $Y2=1.44
r163 45 74 32.8636 $w=3.52e-07 $l=2.4e-07 $layer=POLY_cond $X=1.51 $Y=1.5
+ $X2=1.75 $Y2=1.5
r164 45 72 8.90057 $w=3.52e-07 $l=6.5e-08 $layer=POLY_cond $X=1.51 $Y=1.5
+ $X2=1.445 $Y2=1.5
r165 44 48 62.8485 $w=1.78e-07 $l=1.02e-06 $layer=LI1_cond $X=1.51 $Y=1.445
+ $X2=2.53 $Y2=1.445
r166 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.51
+ $Y=1.44 $X2=1.51 $Y2=1.44
r167 42 51 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.65 $Y=1.445
+ $X2=2.735 $Y2=1.355
r168 42 48 7.39394 $w=1.78e-07 $l=1.2e-07 $layer=LI1_cond $X=2.65 $Y=1.445
+ $X2=2.53 $Y2=1.445
r169 38 79 22.7654 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.62 $Y=1.275
+ $X2=2.62 $Y2=1.5
r170 38 40 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.62 $Y=1.275
+ $X2=2.62 $Y2=0.655
r171 34 49 30.8097 $w=3.52e-07 $l=2.25e-07 $layer=POLY_cond $X=2.305 $Y=1.5
+ $X2=2.53 $Y2=1.5
r172 34 76 17.1165 $w=3.52e-07 $l=1.25e-07 $layer=POLY_cond $X=2.305 $Y=1.5
+ $X2=2.18 $Y2=1.5
r173 34 36 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.305 $Y=1.605
+ $X2=2.305 $Y2=2.465
r174 30 76 22.7654 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.18 $Y=1.275
+ $X2=2.18 $Y2=1.5
r175 30 32 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.18 $Y=1.275
+ $X2=2.18 $Y2=0.655
r176 26 76 41.7642 $w=3.52e-07 $l=3.05e-07 $layer=POLY_cond $X=1.875 $Y=1.5
+ $X2=2.18 $Y2=1.5
r177 26 74 17.1165 $w=3.52e-07 $l=1.25e-07 $layer=POLY_cond $X=1.875 $Y=1.5
+ $X2=1.75 $Y2=1.5
r178 26 28 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.875 $Y=1.605
+ $X2=1.875 $Y2=2.465
r179 22 74 22.7654 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.75 $Y=1.275
+ $X2=1.75 $Y2=1.5
r180 22 24 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.75 $Y=1.275
+ $X2=1.75 $Y2=0.655
r181 19 72 22.7654 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.445 $Y=1.725
+ $X2=1.445 $Y2=1.5
r182 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.445 $Y=1.725
+ $X2=1.445 $Y2=2.465
r183 15 71 22.7654 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.32 $Y=1.275
+ $X2=1.32 $Y2=1.5
r184 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.32 $Y=1.275
+ $X2=1.32 $Y2=0.655
r185 13 71 26.4837 $w=3.52e-07 $l=1.83712e-07 $layer=POLY_cond $X=1.245 $Y=1.65
+ $X2=1.32 $Y2=1.5
r186 13 14 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.245 $Y=1.65
+ $X2=1.09 $Y2=1.65
r187 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.015 $Y=1.725
+ $X2=1.09 $Y2=1.65
r188 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.015 $Y=1.725
+ $X2=1.015 $Y2=2.465
r189 3 58 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=3.64
+ $Y=1.835 $X2=3.78 $Y2=2.65
r190 3 56 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=3.64
+ $Y=1.835 $X2=3.78 $Y2=1.97
r191 2 68 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.235 $X2=5.11 $Y2=0.76
r192 1 62 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.6
+ $Y=0.235 $X2=3.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%A_42_47# 1 2 9 13 17 21 23 27 31 36 39 42 45
+ 48 50 51 53 55
c103 23 0 6.74193e-20 $X=3.45 $Y=1.51
c104 17 0 2.82339e-20 $X=3.955 $Y=0.655
r105 54 55 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.112 $Y=1.705
+ $X2=3.112 $Y2=1.875
r106 50 51 8.17249 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.095
+ $X2=0.272 $Y2=1.93
r107 48 51 55.4545 $w=1.78e-07 $l=9e-07 $layer=LI1_cond $X=0.18 $Y=1.03 $X2=0.18
+ $Y2=1.93
r108 45 54 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.155 $Y=1.51
+ $X2=3.155 $Y2=1.705
r109 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.155
+ $Y=1.51 $X2=3.155 $Y2=1.51
r110 42 55 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.99 $Y=2.37
+ $X2=2.99 $Y2=1.875
r111 40 53 4.19346 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.455 $Y=2.455
+ $X2=0.272 $Y2=2.455
r112 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=2.455
+ $X2=2.99 $Y2=2.37
r113 39 40 159.84 $w=1.68e-07 $l=2.45e-06 $layer=LI1_cond $X=2.905 $Y=2.455
+ $X2=0.455 $Y2=2.455
r114 36 53 2.63236 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.272 $Y=2.37
+ $X2=0.272 $Y2=2.455
r115 35 50 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=0.272 $Y=2.112
+ $X2=0.272 $Y2=2.095
r116 35 36 8.14604 $w=3.63e-07 $l=2.58e-07 $layer=LI1_cond $X=0.272 $Y=2.112
+ $X2=0.272 $Y2=2.37
r117 29 48 8.30054 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.26 $Y=0.86
+ $X2=0.26 $Y2=1.03
r118 29 31 14.914 $w=3.38e-07 $l=4.4e-07 $layer=LI1_cond $X=0.26 $Y=0.86
+ $X2=0.26 $Y2=0.42
r119 26 27 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.955 $Y=1.51
+ $X2=3.995 $Y2=1.51
r120 25 26 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=3.565 $Y=1.51
+ $X2=3.955 $Y2=1.51
r121 24 25 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.525 $Y=1.51
+ $X2=3.565 $Y2=1.51
r122 23 46 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=3.45 $Y=1.51
+ $X2=3.155 $Y2=1.51
r123 23 24 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.45 $Y=1.51
+ $X2=3.525 $Y2=1.51
r124 19 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.675
+ $X2=3.995 $Y2=1.51
r125 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.995 $Y=1.675
+ $X2=3.995 $Y2=2.465
r126 15 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=1.345
+ $X2=3.955 $Y2=1.51
r127 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.955 $Y=1.345
+ $X2=3.955 $Y2=0.655
r128 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.675
+ $X2=3.565 $Y2=1.51
r129 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.565 $Y=1.675
+ $X2=3.565 $Y2=2.465
r130 7 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.345
+ $X2=3.525 $Y2=1.51
r131 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.525 $Y=1.345
+ $X2=3.525 $Y2=0.655
r132 2 53 300 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.495
r133 2 50 600 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.095
r134 1 31 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.235 $X2=0.335 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%A2 3 7 11 15 18 20 23 25 30 31 33 34 35
c87 25 0 2.82339e-20 $X=4.56 $Y=1.48
c88 3 0 1.34732e-19 $X=4.425 $Y=2.465
r89 34 35 15.7161 $w=3.48e-07 $l=3.95e-07 $layer=LI1_cond $X=5.04 $Y=2.03
+ $X2=5.435 $Y2=2.03
r90 33 34 15.7161 $w=3.48e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=2.03
+ $X2=5.04 $Y2=2.03
r91 31 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.51
+ $X2=5.845 $Y2=1.675
r92 31 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.51
+ $X2=5.845 $Y2=1.345
r93 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.845
+ $Y=1.51 $X2=5.845 $Y2=1.51
r94 27 30 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=5.55 $Y=1.492
+ $X2=5.845 $Y2=1.492
r95 23 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.46
+ $X2=4.445 $Y2=1.625
r96 23 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.46
+ $X2=4.445 $Y2=1.295
r97 22 25 4.57003 $w=2.88e-07 $l=1.15e-07 $layer=LI1_cond $X=4.445 $Y=1.48
+ $X2=4.56 $Y2=1.48
r98 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.445
+ $Y=1.46 $X2=4.445 $Y2=1.46
r99 20 35 3.05086 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=5.55 $Y=1.94 $X2=5.55
+ $Y2=2.03
r100 19 27 2.39218 $w=2.3e-07 $l=1.53e-07 $layer=LI1_cond $X=5.55 $Y=1.645
+ $X2=5.55 $Y2=1.492
r101 19 20 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.55 $Y=1.645
+ $X2=5.55 $Y2=1.94
r102 18 33 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.56 $Y=1.94 $X2=4.56
+ $Y2=2.03
r103 17 25 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.56 $Y=1.625
+ $X2=4.56 $Y2=1.48
r104 17 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.56 $Y=1.625
+ $X2=4.56 $Y2=1.94
r105 15 46 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.755 $Y=2.465
+ $X2=5.755 $Y2=1.675
r106 11 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.755 $Y=0.655
+ $X2=5.755 $Y2=1.345
r107 7 42 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.465 $Y=0.655
+ $X2=4.465 $Y2=1.295
r108 3 43 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.425 $Y=2.465
+ $X2=4.425 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%A1 3 7 11 15 17 23 24
c50 23 0 1.34732e-19 $X=5.1 $Y=1.51
r51 22 24 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=5.1 $Y=1.51
+ $X2=5.325 $Y2=1.51
r52 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.1
+ $Y=1.51 $X2=5.1 $Y2=1.51
r53 19 22 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.895 $Y=1.51
+ $X2=5.1 $Y2=1.51
r54 17 23 4.89394 $w=3.63e-07 $l=1.55e-07 $layer=LI1_cond $X=5.082 $Y=1.665
+ $X2=5.082 $Y2=1.51
r55 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.675
+ $X2=5.325 $Y2=1.51
r56 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.325 $Y=1.675
+ $X2=5.325 $Y2=2.465
r57 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.345
+ $X2=5.325 $Y2=1.51
r58 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.325 $Y=1.345
+ $X2=5.325 $Y2=0.655
r59 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=1.675
+ $X2=4.895 $Y2=1.51
r60 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.895 $Y=1.675
+ $X2=4.895 $Y2=2.465
r61 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=1.345
+ $X2=4.895 $Y2=1.51
r62 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.895 $Y=1.345
+ $X2=4.895 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%VPWR 1 2 3 4 5 18 22 26 30 34 36 38 43 48 53
+ 58 65 66 69 72 75 78 81
r92 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r96 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 66 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r98 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r99 63 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.705 $Y=3.33
+ $X2=5.54 $Y2=3.33
r100 63 65 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.705 $Y=3.33 $X2=6
+ $Y2=3.33
r101 62 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r102 62 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 59 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=3.33
+ $X2=4.64 $Y2=3.33
r105 59 61 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.805 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=3.33
+ $X2=5.54 $Y2=3.33
r107 58 61 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.375 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 57 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.52 $Y2=3.33
r111 54 56 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.64 $Y2=3.33
r113 53 56 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 52 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 52 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.66 $Y2=3.33
r118 49 51 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 48 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.52 $Y2=3.33
r120 48 51 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 47 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 47 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r124 44 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r125 44 46 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 43 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.66 $Y2=3.33
r127 43 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 41 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 38 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r131 38 40 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 36 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 36 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 32 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.54 $Y=3.245
+ $X2=5.54 $Y2=3.33
r135 32 34 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.54 $Y=3.245
+ $X2=5.54 $Y2=2.75
r136 28 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=3.245
+ $X2=4.64 $Y2=3.33
r137 28 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.64 $Y=3.245
+ $X2=4.64 $Y2=2.75
r138 24 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=3.33
r139 24 26 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=2.875
r140 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=3.245
+ $X2=1.66 $Y2=3.33
r141 20 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=3.245
+ $X2=1.66 $Y2=2.875
r142 16 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r143 16 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=2.875
r144 5 34 600 $w=1.7e-07 $l=9.8251e-07 $layer=licon1_PDIFF $count=1 $X=5.4
+ $Y=1.835 $X2=5.54 $Y2=2.75
r145 4 30 600 $w=1.7e-07 $l=9.8251e-07 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=1.835 $X2=4.64 $Y2=2.75
r146 3 26 600 $w=1.7e-07 $l=1.10779e-06 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.835 $X2=2.52 $Y2=2.875
r147 2 22 600 $w=1.7e-07 $l=1.10779e-06 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.835 $X2=1.66 $Y2=2.875
r148 1 18 600 $w=1.7e-07 $l=1.10779e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%X 1 2 3 4 14 15 16 19 21 25 27 28 29 30 31
+ 32 39 45
r67 43 45 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.165 $Y=2 $X2=1.2
+ $Y2=2
r68 31 32 15.8461 $w=3.98e-07 $l=5.5e-07 $layer=LI1_cond $X=2.09 $Y=2 $X2=2.64
+ $Y2=2
r69 30 31 11.8125 $w=3.98e-07 $l=4.1e-07 $layer=LI1_cond $X=1.68 $Y=2 $X2=2.09
+ $Y2=2
r70 29 39 2.84813 $w=3.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.08 $Y=2
+ $X2=0.995 $Y2=2.065
r71 29 43 2.84813 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=2 $X2=1.165
+ $Y2=2
r72 29 30 13.109 $w=3.98e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=2 $X2=1.68
+ $Y2=2
r73 29 45 0.720277 $w=3.98e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=2 $X2=1.2
+ $Y2=2
r74 28 39 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=2.065
+ $X2=0.995 $Y2=2.065
r75 23 25 36.0455 $w=1.78e-07 $l=5.85e-07 $layer=LI1_cond $X=2.39 $Y=1.005
+ $X2=2.39 $Y2=0.42
r76 22 27 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.63 $Y=1.09
+ $X2=1.535 $Y2=1.09
r77 21 23 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.3 $Y=1.09
+ $X2=2.39 $Y2=1.005
r78 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.3 $Y=1.09 $X2=1.63
+ $Y2=1.09
r79 17 27 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=1.005
+ $X2=1.535 $Y2=1.09
r80 17 19 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=1.535 $Y=1.005
+ $X2=1.535 $Y2=0.42
r81 15 27 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.44 $Y=1.09
+ $X2=1.535 $Y2=1.09
r82 15 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.44 $Y=1.09
+ $X2=1.165 $Y2=1.09
r83 14 29 3.86674 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.08 $Y=1.8 $X2=1.08
+ $Y2=2
r84 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.08 $Y=1.175
+ $X2=1.165 $Y2=1.09
r85 13 14 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.08 $Y=1.175
+ $X2=1.08 $Y2=1.8
r86 4 31 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.09 $Y2=2.035
r87 3 29 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.835 $X2=1.23 $Y2=2.035
r88 2 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.255
+ $Y=0.235 $X2=2.395 $Y2=0.42
r89 1 19 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.395
+ $Y=0.235 $X2=1.535 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%A_645_367# 1 2 3 4 13 15 17 21 25 29 33 42
+ 44
r54 31 44 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=2.29 $X2=5.985
+ $Y2=2.375
r55 31 33 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=5.985 $Y=2.29
+ $X2=5.985 $Y2=1.98
r56 30 42 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.205 $Y=2.375
+ $X2=5.09 $Y2=2.375
r57 29 44 3.18746 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.835 $Y=2.375
+ $X2=5.985 $Y2=2.375
r58 29 30 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.835 $Y=2.375
+ $X2=5.205 $Y2=2.375
r59 26 40 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.305 $Y=2.375
+ $X2=4.21 $Y2=2.375
r60 25 42 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.975 $Y=2.375
+ $X2=5.09 $Y2=2.375
r61 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=2.375
+ $X2=4.305 $Y2=2.375
r62 23 40 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.21 $Y=2.46 $X2=4.21
+ $Y2=2.375
r63 23 24 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=4.21 $Y=2.46
+ $X2=4.21 $Y2=2.905
r64 19 40 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.21 $Y=2.29 $X2=4.21
+ $Y2=2.375
r65 19 21 19.2632 $w=1.88e-07 $l=3.3e-07 $layer=LI1_cond $X=4.21 $Y=2.29
+ $X2=4.21 $Y2=1.96
r66 18 38 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.445 $Y=2.99 $X2=3.345
+ $Y2=2.99
r67 17 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.115 $Y=2.99
+ $X2=4.21 $Y2=2.905
r68 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.115 $Y=2.99
+ $X2=3.445 $Y2=2.99
r69 13 38 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=2.905
+ $X2=3.345 $Y2=2.99
r70 13 15 38.5409 $w=1.98e-07 $l=6.95e-07 $layer=LI1_cond $X=3.345 $Y=2.905
+ $X2=3.345 $Y2=2.21
r71 4 44 300 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_PDIFF $count=2 $X=5.83
+ $Y=1.835 $X2=5.97 $Y2=2.405
r72 4 33 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.835 $X2=5.97 $Y2=1.98
r73 3 42 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=4.97
+ $Y=1.835 $X2=5.11 $Y2=2.455
r74 2 40 300 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_PDIFF $count=2 $X=4.07
+ $Y=1.835 $X2=4.21 $Y2=2.405
r75 2 21 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.07
+ $Y=1.835 $X2=4.21 $Y2=1.96
r76 1 38 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.835 $X2=3.35 $Y2=2.91
r77 1 15 400 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.835 $X2=3.35 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%VGND 1 2 3 4 5 18 22 24 28 30 32 35 36 37 39
+ 48 52 61 71 75
r87 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r88 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r89 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r90 59 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r91 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r93 56 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r94 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r95 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 53 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.17
+ $Y2=0
r97 53 55 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.56
+ $Y2=0
r98 52 74 4.29523 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=5.855 $Y=0 $X2=6.047
+ $Y2=0
r99 52 58 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.855 $Y=0 $X2=5.52
+ $Y2=0
r100 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r101 48 68 5.34892 $w=8.03e-07 $l=3.6e-07 $layer=LI1_cond $X=3.072 $Y=0
+ $X2=3.072 $Y2=0.36
r102 48 50 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.64
+ $Y2=0
r103 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r104 47 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r105 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r106 44 61 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=0.935
+ $Y2=0
r107 44 46 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.68
+ $Y2=0
r108 42 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r109 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r110 39 61 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.935
+ $Y2=0
r111 39 41 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.24
+ $Y2=0
r112 37 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r113 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r114 37 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r115 35 46 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.68
+ $Y2=0
r116 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.965
+ $Y2=0
r117 34 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.64
+ $Y2=0
r118 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=1.965
+ $Y2=0
r119 30 74 3.06482 $w=2.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.995 $Y=0.085
+ $X2=6.047 $Y2=0
r120 30 32 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.995 $Y=0.085
+ $X2=5.995 $Y2=0.38
r121 26 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0
r122 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0.36
r123 25 48 10.2506 $w=1.7e-07 $l=4.03e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.072 $Y2=0
r124 24 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.17
+ $Y2=0
r125 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.005 $Y=0
+ $X2=3.475 $Y2=0
r126 20 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=0.085
+ $X2=1.965 $Y2=0
r127 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.965 $Y=0.085
+ $X2=1.965 $Y2=0.38
r128 16 61 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0
r129 16 18 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0.38
r130 5 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.83
+ $Y=0.235 $X2=5.97 $Y2=0.38
r131 4 28 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.03
+ $Y=0.235 $X2=4.17 $Y2=0.36
r132 3 68 45.5 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_NDIFF $count=4 $X=2.695
+ $Y=0.235 $X2=3.31 $Y2=0.36
r133 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.825
+ $Y=0.235 $X2=1.965 $Y2=0.38
r134 1 18 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=0.625
+ $Y=0.235 $X2=1.105 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_4%A_908_47# 1 2 9 14 16
r24 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=0.34
+ $X2=4.68 $Y2=0.34
r25 9 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.435 $Y=0.34
+ $X2=5.56 $Y2=0.34
r26 9 10 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.435 $Y=0.34
+ $X2=4.845 $Y2=0.34
r27 2 16 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.4
+ $Y=0.235 $X2=5.54 $Y2=0.42
r28 1 14 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.54
+ $Y=0.235 $X2=4.68 $Y2=0.37
.ends

