* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_1178_399# a_831_47# a_1517_63# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_610_487# a_831_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1149_125# a_1178_399# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1178_399# a_610_487# a_1517_63# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 VPWR a_1517_63# a_1665_381# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_1517_63# a_610_487# a_1670_63# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1047_125# a_610_487# a_1136_451# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_55_119# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_328_119# a_831_47# a_1047_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1517_63# a_831_47# a_1623_493# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1623_493# a_1665_381# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 Q a_1665_381# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_414_487# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VGND a_55_119# a_256_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1047_125# a_831_47# a_1149_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Q a_1665_381# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_256_487# D a_328_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 VPWR a_610_487# a_831_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VGND a_1517_63# a_1665_381# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_328_119# a_610_487# a_1047_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_1665_381# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_55_119# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_464_119# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND CLK a_610_487# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_328_119# a_55_119# a_414_487# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_256_119# D a_328_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1136_451# a_1178_399# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 VGND a_1047_125# a_1178_399# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 a_328_119# SCE a_464_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1670_63# a_1665_381# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VPWR a_1047_125# a_1178_399# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X31 VPWR SCE a_256_487# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 VPWR CLK a_610_487# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 VPWR a_1665_381# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
