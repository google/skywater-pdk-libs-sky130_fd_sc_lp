* File: sky130_fd_sc_lp__or3_2.pxi.spice
* Created: Fri Aug 28 11:23:15 2020
* 
x_PM_SKY130_FD_SC_LP__OR3_2%C N_C_M1006_g N_C_M1009_g C C C N_C_c_64_n
+ PM_SKY130_FD_SC_LP__OR3_2%C
x_PM_SKY130_FD_SC_LP__OR3_2%B N_B_M1001_g N_B_c_93_n N_B_M1008_g B B B
+ N_B_c_95_n PM_SKY130_FD_SC_LP__OR3_2%B
x_PM_SKY130_FD_SC_LP__OR3_2%A N_A_c_130_n N_A_M1002_g N_A_c_125_n N_A_c_126_n
+ N_A_M1003_g A A N_A_c_129_n PM_SKY130_FD_SC_LP__OR3_2%A
x_PM_SKY130_FD_SC_LP__OR3_2%A_35_60# N_A_35_60#_M1006_s N_A_35_60#_M1008_d
+ N_A_35_60#_M1009_s N_A_35_60#_c_170_n N_A_35_60#_M1005_g N_A_35_60#_M1000_g
+ N_A_35_60#_c_172_n N_A_35_60#_M1007_g N_A_35_60#_M1004_g N_A_35_60#_c_174_n
+ N_A_35_60#_c_175_n N_A_35_60#_c_176_n N_A_35_60#_c_177_n N_A_35_60#_c_178_n
+ N_A_35_60#_c_179_n N_A_35_60#_c_180_n N_A_35_60#_c_188_n N_A_35_60#_c_181_n
+ N_A_35_60#_c_241_p N_A_35_60#_c_182_n N_A_35_60#_c_183_n N_A_35_60#_c_184_n
+ PM_SKY130_FD_SC_LP__OR3_2%A_35_60#
x_PM_SKY130_FD_SC_LP__OR3_2%VPWR N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_c_269_n
+ N_VPWR_c_270_n N_VPWR_c_271_n VPWR N_VPWR_c_272_n N_VPWR_c_273_n
+ N_VPWR_c_274_n N_VPWR_c_268_n PM_SKY130_FD_SC_LP__OR3_2%VPWR
x_PM_SKY130_FD_SC_LP__OR3_2%X N_X_M1005_d N_X_M1000_s N_X_c_292_n X X X
+ N_X_c_293_n X PM_SKY130_FD_SC_LP__OR3_2%X
x_PM_SKY130_FD_SC_LP__OR3_2%VGND N_VGND_M1006_d N_VGND_M1003_d N_VGND_M1007_s
+ N_VGND_c_317_n N_VGND_c_318_n VGND N_VGND_c_319_n N_VGND_c_320_n
+ N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n PM_SKY130_FD_SC_LP__OR3_2%VGND
cc_1 VNB N_C_M1006_g 0.0485722f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.51
cc_2 VNB N_C_M1009_g 0.00410587f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.045
cc_3 VNB C 0.00842391f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C_c_64_n 0.0327668f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.415
cc_5 VNB N_B_M1001_g 0.0161185f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.51
cc_6 VNB N_B_c_93_n 0.0471919f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.58
cc_7 VNB N_B_M1008_g 0.0290967f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.045
cc_8 VNB N_B_c_95_n 0.00308781f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.58
cc_9 VNB N_A_c_125_n 0.0109242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_c_126_n 0.00516844f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.58
cc_11 VNB N_A_M1003_g 0.0402682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A 0.00612827f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_A_c_129_n 0.0333316f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.415
cc_14 VNB N_A_35_60#_c_170_n 0.0180467f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_15 VNB N_A_35_60#_M1000_g 0.00360915f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.415
cc_16 VNB N_A_35_60#_c_172_n 0.0186777f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.415
cc_17 VNB N_A_35_60#_M1004_g 0.00593158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_35_60#_c_174_n 0.0150147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_35_60#_c_175_n 0.037265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_35_60#_c_176_n 0.00900833f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.775
cc_21 VNB N_A_35_60#_c_177_n 0.00191899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_35_60#_c_178_n 5.86146e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_35_60#_c_179_n 0.00767351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_35_60#_c_180_n 0.0121587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_35_60#_c_181_n 0.00574803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_35_60#_c_182_n 0.0189305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_35_60#_c_183_n 0.0731534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_35_60#_c_184_n 0.023651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_268_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_292_n 9.01419e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_31 VNB N_X_c_293_n 0.00197987f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.775
cc_32 VNB N_VGND_c_317_n 0.0121431f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_33 VNB N_VGND_c_318_n 0.0148507f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_34 VNB N_VGND_c_319_n 0.0193791f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.665
cc_35 VNB N_VGND_c_320_n 0.0163982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_321_n 0.0153331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_322_n 0.0247102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_323_n 0.197281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_C_M1009_g 0.0278562f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.045
cc_40 VPB C 0.00441444f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_41 VPB C 4.09303e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_42 VPB N_B_M1001_g 0.0234802f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.51
cc_43 VPB N_B_c_95_n 0.00116715f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=1.58
cc_44 VPB N_A_c_130_n 0.0224245f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.25
cc_45 VPB N_A_c_125_n 0.0109242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_c_126_n 0.00195529f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.58
cc_47 VPB A 0.0044923f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_48 VPB N_A_c_129_n 0.0135629f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=1.415
cc_49 VPB N_A_35_60#_M1000_g 0.0245057f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=1.415
cc_50 VPB N_A_35_60#_M1004_g 0.0272217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_35_60#_c_175_n 0.0133967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_35_60#_c_188_n 0.028873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_269_n 0.050046f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_54 VPB N_VPWR_c_270_n 0.0138386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_271_n 0.0548501f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=1.415
cc_56 VPB N_VPWR_c_272_n 0.0503536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_273_n 0.0181698f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.775
cc_58 VPB N_VPWR_c_274_n 0.0134351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_268_n 0.10754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_X_c_293_n 0.00165165f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.775
cc_61 N_C_M1009_g N_B_M1001_g 0.0444618f $X=0.585 $Y=2.045 $X2=0 $Y2=0
cc_62 C N_B_M1001_g 0.00339111f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_63 N_C_M1006_g N_B_c_93_n 0.0100007f $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_64 C N_B_c_93_n 0.00339111f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_C_c_64_n N_B_c_93_n 0.0198232f $X=0.51 $Y=1.415 $X2=0 $Y2=0
cc_66 N_C_M1006_g N_B_M1008_g 0.00881494f $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_67 N_C_M1006_g N_B_c_95_n 4.89415e-19 $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_68 C N_B_c_95_n 0.058339f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_C_M1006_g N_A_35_60#_c_175_n 0.00955913f $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_70 N_C_M1009_g N_A_35_60#_c_175_n 0.00390838f $X=0.585 $Y=2.045 $X2=0 $Y2=0
cc_71 C N_A_35_60#_c_175_n 0.0510017f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 C N_A_35_60#_c_175_n 0.00682423f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_73 N_C_c_64_n N_A_35_60#_c_175_n 0.00813358f $X=0.51 $Y=1.415 $X2=0 $Y2=0
cc_74 N_C_M1006_g N_A_35_60#_c_176_n 0.0150119f $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_75 C N_A_35_60#_c_176_n 0.0267725f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_C_c_64_n N_A_35_60#_c_176_n 0.00141194f $X=0.51 $Y=1.415 $X2=0 $Y2=0
cc_77 N_C_c_64_n N_A_35_60#_c_180_n 0.00171235f $X=0.51 $Y=1.415 $X2=0 $Y2=0
cc_78 N_C_M1009_g N_A_35_60#_c_188_n 7.88459e-19 $X=0.585 $Y=2.045 $X2=0 $Y2=0
cc_79 C N_A_35_60#_c_188_n 0.00242983f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_C_c_64_n N_A_35_60#_c_188_n 0.00279372f $X=0.51 $Y=1.415 $X2=0 $Y2=0
cc_81 C A_132_367# 0.00500727f $X=0.635 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_82 N_C_M1006_g N_VGND_c_320_n 0.00317679f $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_83 N_C_M1006_g N_VGND_c_321_n 0.0116578f $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_84 N_C_M1006_g N_VGND_c_323_n 0.00453221f $X=0.515 $Y=0.51 $X2=0 $Y2=0
cc_85 N_B_c_95_n N_A_c_130_n 0.0190163f $X=1.195 $Y=1.205 $X2=-0.19 $Y2=-0.245
cc_86 N_B_M1001_g N_A_c_126_n 0.0480278f $X=0.96 $Y=2.045 $X2=0 $Y2=0
cc_87 N_B_c_93_n N_A_c_126_n 0.00781326f $X=1.285 $Y=1.015 $X2=0 $Y2=0
cc_88 N_B_c_95_n N_A_c_126_n 0.00542634f $X=1.195 $Y=1.205 $X2=0 $Y2=0
cc_89 N_B_M1008_g N_A_M1003_g 0.0344924f $X=1.285 $Y=0.51 $X2=0 $Y2=0
cc_90 N_B_c_95_n N_A_M1003_g 6.67978e-19 $X=1.195 $Y=1.205 $X2=0 $Y2=0
cc_91 N_B_c_93_n A 0.00174379f $X=1.285 $Y=1.015 $X2=0 $Y2=0
cc_92 N_B_c_95_n A 0.0501448f $X=1.195 $Y=1.205 $X2=0 $Y2=0
cc_93 N_B_M1001_g N_A_c_129_n 0.00253273f $X=0.96 $Y=2.045 $X2=0 $Y2=0
cc_94 N_B_c_93_n N_A_c_129_n 0.00541831f $X=1.285 $Y=1.015 $X2=0 $Y2=0
cc_95 N_B_c_95_n N_A_c_129_n 7.8856e-19 $X=1.195 $Y=1.205 $X2=0 $Y2=0
cc_96 N_B_c_93_n N_A_35_60#_c_176_n 0.0106669f $X=1.285 $Y=1.015 $X2=0 $Y2=0
cc_97 N_B_M1008_g N_A_35_60#_c_176_n 0.0134899f $X=1.285 $Y=0.51 $X2=0 $Y2=0
cc_98 N_B_c_95_n N_A_35_60#_c_176_n 0.0233133f $X=1.195 $Y=1.205 $X2=0 $Y2=0
cc_99 N_B_c_95_n A_207_367# 0.00433061f $X=1.195 $Y=1.205 $X2=-0.19 $Y2=-0.245
cc_100 N_B_c_95_n N_VPWR_c_269_n 0.0163669f $X=1.195 $Y=1.205 $X2=0 $Y2=0
cc_101 N_B_M1008_g N_VGND_c_318_n 0.00317679f $X=1.285 $Y=0.51 $X2=0 $Y2=0
cc_102 N_B_M1008_g N_VGND_c_321_n 0.00762612f $X=1.285 $Y=0.51 $X2=0 $Y2=0
cc_103 N_B_M1008_g N_VGND_c_323_n 0.00398819f $X=1.285 $Y=0.51 $X2=0 $Y2=0
cc_104 N_A_M1003_g N_A_35_60#_c_170_n 0.026908f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_105 A N_A_35_60#_c_170_n 0.00109911f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 A N_A_35_60#_M1000_g 9.35115e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A_c_129_n N_A_35_60#_M1000_g 0.00627085f $X=1.8 $Y=1.415 $X2=0 $Y2=0
cc_108 N_A_M1003_g N_A_35_60#_c_177_n 0.00504915f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_109 N_A_M1003_g N_A_35_60#_c_178_n 0.0126445f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_110 A N_A_35_60#_c_178_n 0.017868f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A_c_129_n N_A_35_60#_c_178_n 9.20375e-19 $X=1.8 $Y=1.415 $X2=0 $Y2=0
cc_112 N_A_M1003_g N_A_35_60#_c_181_n 0.00367301f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_113 A N_A_35_60#_c_181_n 0.00994412f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_114 A N_A_35_60#_c_183_n 0.00156739f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A_c_129_n N_A_35_60#_c_183_n 0.0166368f $X=1.8 $Y=1.415 $X2=0 $Y2=0
cc_116 N_A_c_130_n N_VPWR_c_269_n 0.0156803f $X=1.32 $Y=1.73 $X2=0 $Y2=0
cc_117 N_A_c_125_n N_VPWR_c_269_n 0.0033383f $X=1.635 $Y=1.655 $X2=0 $Y2=0
cc_118 A N_VPWR_c_269_n 0.0408943f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_119 N_A_M1003_g N_X_c_292_n 0.00101933f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_120 A N_X_c_292_n 0.00129542f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_121 A N_X_c_293_n 0.0222237f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A_c_129_n N_X_c_293_n 0.00156165f $X=1.8 $Y=1.415 $X2=0 $Y2=0
cc_123 A N_VGND_M1003_d 0.00145475f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_124 N_A_M1003_g N_VGND_c_317_n 0.0023262f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_125 N_A_M1003_g N_VGND_c_318_n 0.00359419f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_126 N_A_M1003_g N_VGND_c_321_n 4.56217e-19 $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_127 N_A_M1003_g N_VGND_c_323_n 0.00517167f $X=1.715 $Y=0.51 $X2=0 $Y2=0
cc_128 N_A_35_60#_M1000_g N_VPWR_c_269_n 0.00655144f $X=2.335 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_35_60#_M1004_g N_VPWR_c_271_n 0.00860548f $X=2.765 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_35_60#_c_182_n N_VPWR_c_271_n 0.0173406f $X=2.975 $Y=1.415 $X2=0
+ $Y2=0
cc_131 N_A_35_60#_c_183_n N_VPWR_c_271_n 0.0018562f $X=2.975 $Y=1.415 $X2=0
+ $Y2=0
cc_132 N_A_35_60#_M1000_g N_VPWR_c_273_n 0.0054895f $X=2.335 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_35_60#_M1004_g N_VPWR_c_273_n 0.00533769f $X=2.765 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_35_60#_M1000_g N_VPWR_c_268_n 0.0110654f $X=2.335 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_35_60#_M1004_g N_VPWR_c_268_n 0.0104504f $X=2.765 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_35_60#_c_179_n N_X_M1005_d 0.00431761f $X=2.855 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_35_60#_c_170_n N_X_c_292_n 0.00666696f $X=2.305 $Y=1.25 $X2=0 $Y2=0
cc_138 N_A_35_60#_c_172_n N_X_c_292_n 0.00432227f $X=2.735 $Y=1.25 $X2=0 $Y2=0
cc_139 N_A_35_60#_c_179_n N_X_c_292_n 0.016804f $X=2.855 $Y=0.655 $X2=0 $Y2=0
cc_140 N_A_35_60#_c_184_n N_X_c_292_n 0.0101944f $X=3.032 $Y=1.33 $X2=0 $Y2=0
cc_141 N_A_35_60#_M1000_g X 0.0162895f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_35_60#_M1004_g X 0.0172692f $X=2.765 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_35_60#_c_170_n N_X_c_293_n 0.00107932f $X=2.305 $Y=1.25 $X2=0 $Y2=0
cc_144 N_A_35_60#_M1000_g N_X_c_293_n 0.0100639f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_35_60#_c_172_n N_X_c_293_n 7.6484e-19 $X=2.735 $Y=1.25 $X2=0 $Y2=0
cc_146 N_A_35_60#_M1004_g N_X_c_293_n 0.00628532f $X=2.765 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_35_60#_c_182_n N_X_c_293_n 0.0188368f $X=2.975 $Y=1.415 $X2=0 $Y2=0
cc_148 N_A_35_60#_c_183_n N_X_c_293_n 0.0217865f $X=2.975 $Y=1.415 $X2=0 $Y2=0
cc_149 N_A_35_60#_c_184_n N_X_c_293_n 0.01121f $X=3.032 $Y=1.33 $X2=0 $Y2=0
cc_150 N_A_35_60#_c_176_n N_VGND_M1006_d 0.00551246f $X=1.405 $Y=0.785 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_35_60#_c_178_n N_VGND_M1003_d 0.00154372f $X=1.93 $Y=0.72 $X2=0 $Y2=0
cc_152 N_A_35_60#_c_179_n N_VGND_M1003_d 0.00443723f $X=2.855 $Y=0.655 $X2=0
+ $Y2=0
cc_153 N_A_35_60#_c_241_p N_VGND_M1003_d 0.00971702f $X=2.08 $Y=0.72 $X2=0 $Y2=0
cc_154 N_A_35_60#_c_179_n N_VGND_M1007_s 0.00587656f $X=2.855 $Y=0.655 $X2=0
+ $Y2=0
cc_155 N_A_35_60#_c_184_n N_VGND_M1007_s 0.00503428f $X=3.032 $Y=1.33 $X2=0
+ $Y2=0
cc_156 N_A_35_60#_c_170_n N_VGND_c_317_n 0.00395466f $X=2.305 $Y=1.25 $X2=0
+ $Y2=0
cc_157 N_A_35_60#_c_177_n N_VGND_c_317_n 0.0049059f $X=1.5 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_35_60#_c_178_n N_VGND_c_317_n 0.0249029f $X=1.93 $Y=0.72 $X2=0 $Y2=0
cc_159 N_A_35_60#_c_176_n N_VGND_c_318_n 0.00212688f $X=1.405 $Y=0.785 $X2=0
+ $Y2=0
cc_160 N_A_35_60#_c_177_n N_VGND_c_318_n 0.0157184f $X=1.5 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_35_60#_c_178_n N_VGND_c_318_n 0.00310486f $X=1.93 $Y=0.72 $X2=0 $Y2=0
cc_162 N_A_35_60#_c_170_n N_VGND_c_319_n 0.00365477f $X=2.305 $Y=1.25 $X2=0
+ $Y2=0
cc_163 N_A_35_60#_c_172_n N_VGND_c_319_n 0.00365477f $X=2.735 $Y=1.25 $X2=0
+ $Y2=0
cc_164 N_A_35_60#_c_179_n N_VGND_c_319_n 0.0124536f $X=2.855 $Y=0.655 $X2=0
+ $Y2=0
cc_165 N_A_35_60#_c_174_n N_VGND_c_320_n 0.013428f $X=0.3 $Y=0.51 $X2=0 $Y2=0
cc_166 N_A_35_60#_c_176_n N_VGND_c_320_n 0.00212104f $X=1.405 $Y=0.785 $X2=0
+ $Y2=0
cc_167 N_A_35_60#_c_176_n N_VGND_c_321_n 0.0426493f $X=1.405 $Y=0.785 $X2=0
+ $Y2=0
cc_168 N_A_35_60#_c_177_n N_VGND_c_321_n 0.011231f $X=1.5 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_35_60#_c_172_n N_VGND_c_322_n 0.00873062f $X=2.735 $Y=1.25 $X2=0
+ $Y2=0
cc_170 N_A_35_60#_c_179_n N_VGND_c_322_n 0.0278189f $X=2.855 $Y=0.655 $X2=0
+ $Y2=0
cc_171 N_A_35_60#_c_170_n N_VGND_c_323_n 0.00524019f $X=2.305 $Y=1.25 $X2=0
+ $Y2=0
cc_172 N_A_35_60#_c_172_n N_VGND_c_323_n 0.00572792f $X=2.735 $Y=1.25 $X2=0
+ $Y2=0
cc_173 N_A_35_60#_c_174_n N_VGND_c_323_n 0.0113655f $X=0.3 $Y=0.51 $X2=0 $Y2=0
cc_174 N_A_35_60#_c_176_n N_VGND_c_323_n 0.0106309f $X=1.405 $Y=0.785 $X2=0
+ $Y2=0
cc_175 N_A_35_60#_c_177_n N_VGND_c_323_n 0.00975716f $X=1.5 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A_35_60#_c_178_n N_VGND_c_323_n 0.00665853f $X=1.93 $Y=0.72 $X2=0 $Y2=0
cc_177 N_A_35_60#_c_179_n N_VGND_c_323_n 0.0230988f $X=2.855 $Y=0.655 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_268_n N_X_M1000_s 0.00223559f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_273_n X 0.0196054f $X=2.895 $Y=3.33 $X2=0 $Y2=0
cc_180 N_VPWR_c_268_n X 0.0127183f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_271_n N_X_c_293_n 0.00114352f $X=2.98 $Y=1.98 $X2=0 $Y2=0
