* File: sky130_fd_sc_lp__buf_16.pxi.spice
* Created: Fri Aug 28 10:09:57 2020
* 
x_PM_SKY130_FD_SC_LP__BUF_16%A N_A_M1005_g N_A_M1000_g N_A_M1009_g N_A_M1008_g
+ N_A_M1023_g N_A_M1015_g N_A_M1028_g N_A_M1021_g N_A_M1036_g N_A_M1033_g
+ N_A_M1039_g N_A_M1040_g N_A_c_186_n N_A_c_215_p A N_A_c_188_n
+ PM_SKY130_FD_SC_LP__BUF_16%A
x_PM_SKY130_FD_SC_LP__BUF_16%A_130_47# N_A_130_47#_M1005_s N_A_130_47#_M1023_s
+ N_A_130_47#_M1036_s N_A_130_47#_M1000_d N_A_130_47#_M1015_d
+ N_A_130_47#_M1033_d N_A_130_47#_M1001_g N_A_130_47#_c_319_n
+ N_A_130_47#_M1002_g N_A_130_47#_M1003_g N_A_130_47#_c_320_n
+ N_A_130_47#_M1004_g N_A_130_47#_M1007_g N_A_130_47#_M1006_g
+ N_A_130_47#_M1014_g N_A_130_47#_M1010_g N_A_130_47#_M1016_g
+ N_A_130_47#_M1011_g N_A_130_47#_M1017_g N_A_130_47#_M1012_g
+ N_A_130_47#_M1018_g N_A_130_47#_M1013_g N_A_130_47#_M1019_g
+ N_A_130_47#_M1022_g N_A_130_47#_M1020_g N_A_130_47#_M1025_g
+ N_A_130_47#_M1024_g N_A_130_47#_M1027_g N_A_130_47#_M1026_g
+ N_A_130_47#_M1029_g N_A_130_47#_M1032_g N_A_130_47#_M1030_g
+ N_A_130_47#_M1034_g N_A_130_47#_M1031_g N_A_130_47#_M1035_g
+ N_A_130_47#_M1037_g N_A_130_47#_M1042_g N_A_130_47#_M1038_g
+ N_A_130_47#_M1043_g N_A_130_47#_c_304_n N_A_130_47#_M1041_g
+ N_A_130_47#_c_635_p N_A_130_47#_c_461_p N_A_130_47#_c_305_n
+ N_A_130_47#_c_306_n N_A_130_47#_c_336_n N_A_130_47#_c_337_n
+ N_A_130_47#_c_451_p N_A_130_47#_c_636_p N_A_130_47#_c_368_n
+ N_A_130_47#_c_338_n N_A_130_47#_c_452_p N_A_130_47#_c_626_p
+ N_A_130_47#_c_307_n N_A_130_47#_c_339_n N_A_130_47#_c_340_n
+ N_A_130_47#_c_308_n N_A_130_47#_c_341_n N_A_130_47#_c_309_n
+ N_A_130_47#_c_310_n N_A_130_47#_c_311_n N_A_130_47#_c_312_n
+ N_A_130_47#_c_313_n N_A_130_47#_c_314_n N_A_130_47#_c_315_n
+ N_A_130_47#_c_316_n N_A_130_47#_c_317_n N_A_130_47#_c_318_n
+ PM_SKY130_FD_SC_LP__BUF_16%A_130_47#
x_PM_SKY130_FD_SC_LP__BUF_16%VPWR N_VPWR_M1000_s N_VPWR_M1008_s N_VPWR_M1021_s
+ N_VPWR_M1040_s N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1012_d N_VPWR_M1022_d
+ N_VPWR_M1027_d N_VPWR_M1030_d N_VPWR_M1037_d N_VPWR_M1041_d N_VPWR_c_664_n
+ N_VPWR_c_665_n N_VPWR_c_666_n N_VPWR_c_667_n N_VPWR_c_668_n N_VPWR_c_669_n
+ N_VPWR_c_670_n N_VPWR_c_671_n N_VPWR_c_672_n N_VPWR_c_673_n N_VPWR_c_674_n
+ N_VPWR_c_675_n N_VPWR_c_676_n N_VPWR_c_677_n N_VPWR_c_678_n N_VPWR_c_679_n
+ N_VPWR_c_680_n N_VPWR_c_681_n N_VPWR_c_682_n N_VPWR_c_683_n N_VPWR_c_684_n
+ N_VPWR_c_685_n N_VPWR_c_686_n N_VPWR_c_687_n N_VPWR_c_688_n N_VPWR_c_689_n
+ N_VPWR_c_690_n N_VPWR_c_691_n VPWR N_VPWR_c_692_n N_VPWR_c_693_n
+ N_VPWR_c_694_n N_VPWR_c_695_n N_VPWR_c_696_n N_VPWR_c_697_n N_VPWR_c_698_n
+ N_VPWR_c_663_n PM_SKY130_FD_SC_LP__BUF_16%VPWR
x_PM_SKY130_FD_SC_LP__BUF_16%X N_X_M1001_d N_X_M1007_d N_X_M1016_d N_X_M1018_d
+ N_X_M1020_d N_X_M1026_d N_X_M1034_d N_X_M1042_d N_X_M1002_s N_X_M1006_s
+ N_X_M1011_s N_X_M1013_s N_X_M1025_s N_X_M1029_s N_X_M1031_s N_X_M1038_s X
+ N_X_c_862_n N_X_c_863_n N_X_c_864_n N_X_c_865_n N_X_c_866_n N_X_c_867_n
+ N_X_c_868_n N_X_c_869_n N_X_c_878_n PM_SKY130_FD_SC_LP__BUF_16%X
x_PM_SKY130_FD_SC_LP__BUF_16%VGND N_VGND_M1005_d N_VGND_M1009_d N_VGND_M1028_d
+ N_VGND_M1039_d N_VGND_M1003_s N_VGND_M1014_s N_VGND_M1017_s N_VGND_M1019_s
+ N_VGND_M1024_s N_VGND_M1032_s N_VGND_M1035_s N_VGND_M1043_s N_VGND_c_1048_n
+ N_VGND_c_1049_n N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n
+ N_VGND_c_1053_n N_VGND_c_1054_n N_VGND_c_1055_n N_VGND_c_1056_n
+ N_VGND_c_1057_n N_VGND_c_1058_n N_VGND_c_1059_n N_VGND_c_1060_n
+ N_VGND_c_1061_n N_VGND_c_1062_n N_VGND_c_1063_n N_VGND_c_1064_n
+ N_VGND_c_1065_n N_VGND_c_1066_n N_VGND_c_1067_n N_VGND_c_1068_n
+ N_VGND_c_1069_n N_VGND_c_1070_n N_VGND_c_1071_n N_VGND_c_1072_n
+ N_VGND_c_1073_n VGND N_VGND_c_1074_n N_VGND_c_1075_n N_VGND_c_1076_n
+ N_VGND_c_1077_n N_VGND_c_1078_n N_VGND_c_1079_n N_VGND_c_1080_n
+ N_VGND_c_1081_n N_VGND_c_1082_n N_VGND_c_1083_n
+ PM_SKY130_FD_SC_LP__BUF_16%VGND
cc_1 VNB N_A_M1005_g 0.0324974f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.655
cc_2 VNB N_A_M1000_g 7.24268e-19 $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_3 VNB N_A_M1009_g 0.021612f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.655
cc_4 VNB N_A_M1008_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.465
cc_5 VNB N_A_M1023_g 0.0215906f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.655
cc_6 VNB N_A_M1015_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=2.465
cc_7 VNB N_A_M1028_g 0.022112f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=0.655
cc_8 VNB N_A_M1021_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=2.465
cc_9 VNB N_A_M1036_g 0.022109f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=0.655
cc_10 VNB N_A_M1033_g 4.57435e-19 $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=2.465
cc_11 VNB N_A_M1039_g 0.0217866f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.655
cc_12 VNB N_A_M1040_g 4.70146e-19 $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=2.465
cc_13 VNB N_A_c_186_n 0.00806404f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.485
cc_14 VNB A 0.0026033f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_15 VNB N_A_c_188_n 0.135916f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.48
cc_16 VNB N_A_130_47#_M1001_g 0.0225241f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.645
cc_17 VNB N_A_130_47#_M1003_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_130_47#_M1007_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=0.655
cc_19 VNB N_A_130_47#_M1014_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.655
cc_20 VNB N_A_130_47#_M1016_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.48
cc_21 VNB N_A_130_47#_M1017_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.48
cc_22 VNB N_A_130_47#_M1018_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.48
cc_23 VNB N_A_130_47#_M1019_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.48
cc_24 VNB N_A_130_47#_M1020_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_130_47#_M1024_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_130_47#_M1026_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_130_47#_M1032_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_130_47#_M1034_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_130_47#_M1035_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_130_47#_M1042_g 0.0232295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_130_47#_M1043_g 0.0332666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_130_47#_c_304_n 0.296242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_130_47#_c_305_n 0.00249586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_130_47#_c_306_n 0.00402102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_130_47#_c_307_n 0.00134483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_130_47#_c_308_n 0.00303174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_130_47#_c_309_n 0.00312313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_130_47#_c_310_n 0.00359692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_130_47#_c_311_n 0.00179809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_130_47#_c_312_n 0.00107293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_130_47#_c_313_n 0.00107293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_130_47#_c_314_n 0.00107293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_130_47#_c_315_n 0.00107293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_130_47#_c_316_n 0.00107293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_130_47#_c_317_n 0.00107293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_130_47#_c_318_n 0.00107293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VPWR_c_663_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_X_c_862_n 0.0042266f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.48
cc_49 VNB N_X_c_863_n 0.00469444f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_50 VNB N_X_c_864_n 0.00469444f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=1.48
cc_51 VNB N_X_c_865_n 0.00469444f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=1.485
cc_52 VNB N_X_c_866_n 0.00469444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_X_c_867_n 0.00469444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_X_c_868_n 0.00469444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_X_c_869_n 0.0050457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1048_n 0.0140954f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.645
cc_57 VNB N_VGND_c_1049_n 0.0441686f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=2.465
cc_58 VNB N_VGND_c_1050_n 0.00400713f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.655
cc_59 VNB N_VGND_c_1051_n 3.19614e-19 $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=2.465
cc_60 VNB N_VGND_c_1052_n 0.00190253f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.48
cc_61 VNB N_VGND_c_1053_n 0.00529363f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=1.48
cc_62 VNB N_VGND_c_1054_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.485
cc_63 VNB N_VGND_c_1055_n 0.00532497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1056_n 0.00532497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1057_n 0.00532497f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.48
cc_66 VNB N_VGND_c_1058_n 0.00532497f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=1.48
cc_67 VNB N_VGND_c_1059_n 0.00532497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1060_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1061_n 0.00532497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1062_n 0.0109056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1063_n 0.0467359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1064_n 0.0153654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1065_n 0.00432792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1066_n 0.0149952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1067_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1068_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1069_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1070_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1071_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1072_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1073_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1074_n 0.01729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1075_n 0.0151146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1076_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1077_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1078_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1079_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1080_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1081_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1082_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1083_n 0.470958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VPB N_A_M1000_g 0.0272502f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_93 VPB N_A_M1008_g 0.0191131f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.465
cc_94 VPB N_A_M1015_g 0.0191131f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=2.465
cc_95 VPB N_A_M1021_g 0.0191131f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=2.465
cc_96 VPB N_A_M1033_g 0.0190927f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.465
cc_97 VPB N_A_M1040_g 0.0192926f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.465
cc_98 VPB N_A_130_47#_c_319_n 0.0153591f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=2.465
cc_99 VPB N_A_130_47#_c_320_n 0.0157473f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=2.465
cc_100 VPB N_A_130_47#_M1006_g 0.0187408f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.465
cc_101 VPB N_A_130_47#_M1010_g 0.0187408f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.465
cc_102 VPB N_A_130_47#_M1011_g 0.0187408f $X=-0.19 $Y=1.655 $X2=1.89 $Y2=1.48
cc_103 VPB N_A_130_47#_M1012_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_130_47#_M1013_g 0.0187408f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=1.48
cc_105 VPB N_A_130_47#_M1022_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_130_47#_M1025_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_130_47#_M1027_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_130_47#_M1029_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_130_47#_M1030_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_130_47#_M1031_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_130_47#_M1037_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_130_47#_M1038_g 0.019202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_130_47#_c_304_n 0.0490622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_130_47#_M1041_g 0.0276562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_130_47#_c_336_n 0.00240582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_130_47#_c_337_n 0.00309037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_130_47#_c_338_n 0.00240157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_130_47#_c_339_n 0.0012141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_130_47#_c_340_n 0.00210233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_130_47#_c_341_n 0.00210233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_130_47#_c_310_n 0.00126874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_130_47#_c_311_n 0.0102159f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_130_47#_c_312_n 0.00152497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_130_47#_c_313_n 0.00152497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_130_47#_c_314_n 0.00152497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_130_47#_c_315_n 0.00152497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_130_47#_c_316_n 0.00152497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_130_47#_c_317_n 0.00152497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_130_47#_c_318_n 0.00152497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_664_n 0.0140695f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.645
cc_131 VPB N_VPWR_c_665_n 0.0615039f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.465
cc_132 VPB N_VPWR_c_666_n 0.00400996f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=1.645
cc_133 VPB N_VPWR_c_667_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.48
cc_134 VPB N_VPWR_c_668_n 0.00194686f $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.485
cc_135 VPB N_VPWR_c_669_n 0.00397862f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_670_n 0.0166024f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.48
cc_137 VPB N_VPWR_c_671_n 0.00400996f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=1.48
cc_138 VPB N_VPWR_c_672_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_673_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_674_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_675_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_676_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_677_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_678_n 0.0108797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_679_n 0.0510625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_680_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_681_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_682_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_683_n 0.00430203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_684_n 0.0149952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_685_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_686_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_687_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_688_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_689_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_690_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_691_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_692_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_693_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_694_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_695_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_696_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_697_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_698_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_663_n 0.048547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_X_c_862_n 0.0012822f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.48
cc_167 VPB N_X_c_863_n 0.00204925f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_168 VPB N_X_c_864_n 0.00204925f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=1.48
cc_169 VPB N_X_c_865_n 0.00204925f $X=-0.19 $Y=1.655 $X2=2.08 $Y2=1.485
cc_170 VPB N_X_c_866_n 0.00204925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_X_c_867_n 0.00204925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_X_c_868_n 0.00204925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_X_c_869_n 0.00276017f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 N_A_M1039_g N_A_130_47#_M1001_g 0.0208615f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_175 N_A_M1040_g N_A_130_47#_c_319_n 0.0208615f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_c_188_n N_A_130_47#_c_304_n 0.0208615f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_177 N_A_M1009_g N_A_130_47#_c_305_n 0.0143403f $X=1.005 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A_M1023_g N_A_130_47#_c_305_n 0.0142259f $X=1.435 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A_c_186_n N_A_130_47#_c_305_n 0.0429575f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_180 N_A_c_188_n N_A_130_47#_c_305_n 0.00243542f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_181 N_A_M1005_g N_A_130_47#_c_306_n 0.00465535f $X=0.575 $Y=0.655 $X2=0 $Y2=0
cc_182 N_A_c_186_n N_A_130_47#_c_306_n 0.0212043f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_183 N_A_c_188_n N_A_130_47#_c_306_n 0.00253619f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_184 N_A_M1008_g N_A_130_47#_c_336_n 0.013787f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_M1015_g N_A_130_47#_c_336_n 0.0138996f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_c_186_n N_A_130_47#_c_336_n 0.0422336f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_187 N_A_c_188_n N_A_130_47#_c_336_n 0.00240656f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_188 N_A_M1000_g N_A_130_47#_c_337_n 0.00218098f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_c_186_n N_A_130_47#_c_337_n 0.0212044f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_190 N_A_c_188_n N_A_130_47#_c_337_n 0.00250529f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_191 N_A_M1028_g N_A_130_47#_c_368_n 0.0129521f $X=1.865 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_M1036_g N_A_130_47#_c_368_n 0.0129521f $X=2.295 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A_c_186_n N_A_130_47#_c_368_n 0.00528015f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_194 N_A_c_215_p N_A_130_47#_c_368_n 0.00528015f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_195 A N_A_130_47#_c_368_n 0.0229606f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A_c_188_n N_A_130_47#_c_368_n 5.3208e-19 $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_197 N_A_M1021_g N_A_130_47#_c_338_n 0.0139311f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A_M1033_g N_A_130_47#_c_338_n 0.0139311f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A_c_186_n N_A_130_47#_c_338_n 0.00857975f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_200 N_A_c_215_p N_A_130_47#_c_338_n 0.00857975f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_201 A N_A_130_47#_c_338_n 0.0263164f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_202 N_A_c_188_n N_A_130_47#_c_338_n 0.00240522f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_203 N_A_M1039_g N_A_130_47#_c_307_n 0.0149674f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A_c_215_p N_A_130_47#_c_307_n 0.0065206f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_205 N_A_M1040_g N_A_130_47#_c_339_n 0.0145946f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_c_215_p N_A_130_47#_c_339_n 0.0065206f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_207 N_A_c_186_n N_A_130_47#_c_340_n 0.0212044f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_208 N_A_c_188_n N_A_130_47#_c_340_n 0.00250529f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_209 N_A_M1028_g N_A_130_47#_c_308_n 0.00416701f $X=1.865 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A_c_186_n N_A_130_47#_c_308_n 0.0167182f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_211 A N_A_130_47#_c_308_n 8.4662e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_212 N_A_c_188_n N_A_130_47#_c_308_n 0.00253619f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_213 N_A_c_215_p N_A_130_47#_c_341_n 0.0212044f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_214 N_A_c_188_n N_A_130_47#_c_341_n 0.00250529f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_215 N_A_M1036_g N_A_130_47#_c_309_n 0.00410876f $X=2.295 $Y=0.655 $X2=0 $Y2=0
cc_216 N_A_c_215_p N_A_130_47#_c_309_n 0.0175338f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_217 A N_A_130_47#_c_309_n 8.45582e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A_c_188_n N_A_130_47#_c_309_n 0.00253619f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_219 N_A_M1039_g N_A_130_47#_c_310_n 0.00706996f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_220 N_A_c_215_p N_A_130_47#_c_310_n 0.0151451f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_221 A N_A_130_47#_c_310_n 0.00462514f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_222 N_A_c_215_p N_A_130_47#_c_311_n 0.00120198f $X=2.57 $Y=1.48 $X2=0 $Y2=0
cc_223 N_A_c_188_n N_A_130_47#_c_311_n 0.00449786f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_224 N_A_M1000_g N_VPWR_c_665_n 0.00579553f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_c_186_n N_VPWR_c_665_n 0.00807001f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_226 N_A_c_188_n N_VPWR_c_665_n 0.00300963f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_227 N_A_M1008_g N_VPWR_c_666_n 0.0016342f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A_M1015_g N_VPWR_c_666_n 0.0016342f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A_M1021_g N_VPWR_c_667_n 0.0016342f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_M1033_g N_VPWR_c_667_n 0.0016342f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_M1040_g N_VPWR_c_668_n 0.00164679f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_M1015_g N_VPWR_c_680_n 0.00585385f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A_M1021_g N_VPWR_c_680_n 0.00585385f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A_M1033_g N_VPWR_c_682_n 0.00585385f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A_M1040_g N_VPWR_c_682_n 0.00585385f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_M1000_g N_VPWR_c_692_n 0.00585385f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_M1008_g N_VPWR_c_692_n 0.00585385f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_M1000_g N_VPWR_c_663_n 0.01183f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A_M1008_g N_VPWR_c_663_n 0.0106302f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_M1015_g N_VPWR_c_663_n 0.0106302f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A_M1021_g N_VPWR_c_663_n 0.0106302f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_242 N_A_M1033_g N_VPWR_c_663_n 0.0106302f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A_M1040_g N_VPWR_c_663_n 0.0106555f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A_M1040_g N_X_c_878_n 7.3936e-19 $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A_M1005_g N_VGND_c_1049_n 0.0046456f $X=0.575 $Y=0.655 $X2=0 $Y2=0
cc_246 N_A_c_186_n N_VGND_c_1049_n 0.00491721f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_247 N_A_c_188_n N_VGND_c_1049_n 0.00268738f $X=2.725 $Y=1.48 $X2=0 $Y2=0
cc_248 N_A_M1009_g N_VGND_c_1050_n 0.00163936f $X=1.005 $Y=0.655 $X2=0 $Y2=0
cc_249 N_A_M1023_g N_VGND_c_1050_n 0.00158356f $X=1.435 $Y=0.655 $X2=0 $Y2=0
cc_250 N_A_M1023_g N_VGND_c_1051_n 0.00101353f $X=1.435 $Y=0.655 $X2=0 $Y2=0
cc_251 N_A_M1028_g N_VGND_c_1051_n 0.0117144f $X=1.865 $Y=0.655 $X2=0 $Y2=0
cc_252 N_A_M1036_g N_VGND_c_1051_n 0.011764f $X=2.295 $Y=0.655 $X2=0 $Y2=0
cc_253 N_A_M1039_g N_VGND_c_1051_n 0.00101962f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_254 N_A_M1039_g N_VGND_c_1052_n 0.00159771f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_255 N_A_M1036_g N_VGND_c_1064_n 0.00486043f $X=2.295 $Y=0.655 $X2=0 $Y2=0
cc_256 N_A_M1039_g N_VGND_c_1064_n 0.00585385f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_257 N_A_M1005_g N_VGND_c_1074_n 0.00585385f $X=0.575 $Y=0.655 $X2=0 $Y2=0
cc_258 N_A_M1009_g N_VGND_c_1074_n 0.00585385f $X=1.005 $Y=0.655 $X2=0 $Y2=0
cc_259 N_A_M1023_g N_VGND_c_1075_n 0.00583607f $X=1.435 $Y=0.655 $X2=0 $Y2=0
cc_260 N_A_M1028_g N_VGND_c_1075_n 0.00486043f $X=1.865 $Y=0.655 $X2=0 $Y2=0
cc_261 N_A_M1005_g N_VGND_c_1083_n 0.0116446f $X=0.575 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A_M1009_g N_VGND_c_1083_n 0.0106302f $X=1.005 $Y=0.655 $X2=0 $Y2=0
cc_263 N_A_M1023_g N_VGND_c_1083_n 0.0105967f $X=1.435 $Y=0.655 $X2=0 $Y2=0
cc_264 N_A_M1028_g N_VGND_c_1083_n 0.00835506f $X=1.865 $Y=0.655 $X2=0 $Y2=0
cc_265 N_A_M1036_g N_VGND_c_1083_n 0.00835506f $X=2.295 $Y=0.655 $X2=0 $Y2=0
cc_266 N_A_M1039_g N_VGND_c_1083_n 0.0106555f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_267 N_A_130_47#_c_336_n N_VPWR_M1008_s 0.00176461f $X=1.52 $Y=1.84 $X2=0
+ $Y2=0
cc_268 N_A_130_47#_c_338_n N_VPWR_M1021_s 0.00176461f $X=2.38 $Y=1.84 $X2=0
+ $Y2=0
cc_269 N_A_130_47#_c_339_n N_VPWR_M1040_s 0.00180544f $X=2.905 $Y=1.84 $X2=0
+ $Y2=0
cc_270 N_A_130_47#_c_337_n N_VPWR_c_665_n 0.00166618f $X=0.92 $Y=1.84 $X2=0
+ $Y2=0
cc_271 N_A_130_47#_c_336_n N_VPWR_c_666_n 0.0135055f $X=1.52 $Y=1.84 $X2=0 $Y2=0
cc_272 N_A_130_47#_c_338_n N_VPWR_c_667_n 0.0135055f $X=2.38 $Y=1.84 $X2=0 $Y2=0
cc_273 N_A_130_47#_c_319_n N_VPWR_c_668_n 0.0129247f $X=3.155 $Y=1.725 $X2=0
+ $Y2=0
cc_274 N_A_130_47#_c_320_n N_VPWR_c_668_n 7.59601e-19 $X=3.585 $Y=1.725 $X2=0
+ $Y2=0
cc_275 N_A_130_47#_c_339_n N_VPWR_c_668_n 0.0146153f $X=2.905 $Y=1.84 $X2=0
+ $Y2=0
cc_276 N_A_130_47#_c_311_n N_VPWR_c_668_n 0.00142796f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_277 N_A_130_47#_c_320_n N_VPWR_c_669_n 0.00208116f $X=3.585 $Y=1.725 $X2=0
+ $Y2=0
cc_278 N_A_130_47#_M1006_g N_VPWR_c_669_n 0.00211566f $X=4.015 $Y=2.465 $X2=0
+ $Y2=0
cc_279 N_A_130_47#_c_304_n N_VPWR_c_669_n 5.29564e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_280 N_A_130_47#_c_311_n N_VPWR_c_669_n 8.68506e-19 $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_281 N_A_130_47#_c_312_n N_VPWR_c_669_n 0.0171314f $X=3.8 $Y=1.49 $X2=0 $Y2=0
cc_282 N_A_130_47#_M1006_g N_VPWR_c_670_n 0.00585385f $X=4.015 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_130_47#_M1010_g N_VPWR_c_670_n 0.00585385f $X=4.445 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A_130_47#_M1010_g N_VPWR_c_671_n 0.00211566f $X=4.445 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_A_130_47#_M1011_g N_VPWR_c_671_n 0.00211566f $X=4.875 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_130_47#_c_304_n N_VPWR_c_671_n 5.29564e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_287 N_A_130_47#_c_311_n N_VPWR_c_671_n 8.68506e-19 $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_288 N_A_130_47#_c_313_n N_VPWR_c_671_n 0.0171314f $X=4.66 $Y=1.49 $X2=0 $Y2=0
cc_289 N_A_130_47#_M1012_g N_VPWR_c_672_n 0.00211566f $X=5.305 $Y=2.465 $X2=0
+ $Y2=0
cc_290 N_A_130_47#_M1013_g N_VPWR_c_672_n 0.00211566f $X=5.735 $Y=2.465 $X2=0
+ $Y2=0
cc_291 N_A_130_47#_c_304_n N_VPWR_c_672_n 5.29564e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_292 N_A_130_47#_c_311_n N_VPWR_c_672_n 8.68506e-19 $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_293 N_A_130_47#_c_314_n N_VPWR_c_672_n 0.0171314f $X=5.52 $Y=1.49 $X2=0 $Y2=0
cc_294 N_A_130_47#_M1022_g N_VPWR_c_673_n 0.00211566f $X=6.165 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_130_47#_M1025_g N_VPWR_c_673_n 0.00211566f $X=6.595 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_130_47#_c_304_n N_VPWR_c_673_n 5.29564e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_297 N_A_130_47#_c_311_n N_VPWR_c_673_n 8.68506e-19 $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_298 N_A_130_47#_c_315_n N_VPWR_c_673_n 0.0171314f $X=6.38 $Y=1.49 $X2=0 $Y2=0
cc_299 N_A_130_47#_M1027_g N_VPWR_c_674_n 0.00211566f $X=7.025 $Y=2.465 $X2=0
+ $Y2=0
cc_300 N_A_130_47#_M1029_g N_VPWR_c_674_n 0.00211566f $X=7.455 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_A_130_47#_c_304_n N_VPWR_c_674_n 5.29564e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_302 N_A_130_47#_c_311_n N_VPWR_c_674_n 8.68506e-19 $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_303 N_A_130_47#_c_316_n N_VPWR_c_674_n 0.0171314f $X=7.24 $Y=1.49 $X2=0 $Y2=0
cc_304 N_A_130_47#_M1030_g N_VPWR_c_675_n 0.00211566f $X=7.885 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_130_47#_M1031_g N_VPWR_c_675_n 0.00211566f $X=8.315 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A_130_47#_c_304_n N_VPWR_c_675_n 5.29564e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_307 N_A_130_47#_c_311_n N_VPWR_c_675_n 8.68506e-19 $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_308 N_A_130_47#_c_317_n N_VPWR_c_675_n 0.0171314f $X=8.1 $Y=1.49 $X2=0 $Y2=0
cc_309 N_A_130_47#_M1031_g N_VPWR_c_676_n 0.00585385f $X=8.315 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A_130_47#_M1037_g N_VPWR_c_676_n 0.00585385f $X=8.745 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_130_47#_M1037_g N_VPWR_c_677_n 0.00211566f $X=8.745 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A_130_47#_M1038_g N_VPWR_c_677_n 0.00211566f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_313 N_A_130_47#_c_304_n N_VPWR_c_677_n 5.29564e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_314 N_A_130_47#_c_311_n N_VPWR_c_677_n 8.68506e-19 $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_315 N_A_130_47#_c_318_n N_VPWR_c_677_n 0.0171314f $X=8.96 $Y=1.49 $X2=0 $Y2=0
cc_316 N_A_130_47#_M1041_g N_VPWR_c_679_n 0.00411939f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_317 N_A_130_47#_c_451_p N_VPWR_c_680_n 0.0149362f $X=1.65 $Y=2.025 $X2=0
+ $Y2=0
cc_318 N_A_130_47#_c_452_p N_VPWR_c_682_n 0.0149362f $X=2.51 $Y=2.025 $X2=0
+ $Y2=0
cc_319 N_A_130_47#_c_319_n N_VPWR_c_684_n 0.00525069f $X=3.155 $Y=1.725 $X2=0
+ $Y2=0
cc_320 N_A_130_47#_c_320_n N_VPWR_c_684_n 0.00585385f $X=3.585 $Y=1.725 $X2=0
+ $Y2=0
cc_321 N_A_130_47#_M1013_g N_VPWR_c_686_n 0.00585385f $X=5.735 $Y=2.465 $X2=0
+ $Y2=0
cc_322 N_A_130_47#_M1022_g N_VPWR_c_686_n 0.00585385f $X=6.165 $Y=2.465 $X2=0
+ $Y2=0
cc_323 N_A_130_47#_M1025_g N_VPWR_c_688_n 0.00585385f $X=6.595 $Y=2.465 $X2=0
+ $Y2=0
cc_324 N_A_130_47#_M1027_g N_VPWR_c_688_n 0.00585385f $X=7.025 $Y=2.465 $X2=0
+ $Y2=0
cc_325 N_A_130_47#_M1029_g N_VPWR_c_690_n 0.00585385f $X=7.455 $Y=2.465 $X2=0
+ $Y2=0
cc_326 N_A_130_47#_M1030_g N_VPWR_c_690_n 0.00585385f $X=7.885 $Y=2.465 $X2=0
+ $Y2=0
cc_327 N_A_130_47#_c_461_p N_VPWR_c_692_n 0.0149362f $X=0.79 $Y=2.025 $X2=0
+ $Y2=0
cc_328 N_A_130_47#_M1011_g N_VPWR_c_693_n 0.00585385f $X=4.875 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_A_130_47#_M1012_g N_VPWR_c_693_n 0.00585385f $X=5.305 $Y=2.465 $X2=0
+ $Y2=0
cc_330 N_A_130_47#_M1038_g N_VPWR_c_694_n 0.00585385f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_331 N_A_130_47#_M1041_g N_VPWR_c_694_n 0.00585385f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_332 N_A_130_47#_M1000_d N_VPWR_c_663_n 0.003017f $X=0.65 $Y=1.835 $X2=0 $Y2=0
cc_333 N_A_130_47#_M1015_d N_VPWR_c_663_n 0.003017f $X=1.51 $Y=1.835 $X2=0 $Y2=0
cc_334 N_A_130_47#_M1033_d N_VPWR_c_663_n 0.003017f $X=2.37 $Y=1.835 $X2=0 $Y2=0
cc_335 N_A_130_47#_c_319_n N_VPWR_c_663_n 0.00897288f $X=3.155 $Y=1.725 $X2=0
+ $Y2=0
cc_336 N_A_130_47#_c_320_n N_VPWR_c_663_n 0.0106914f $X=3.585 $Y=1.725 $X2=0
+ $Y2=0
cc_337 N_A_130_47#_M1006_g N_VPWR_c_663_n 0.0106914f $X=4.015 $Y=2.465 $X2=0
+ $Y2=0
cc_338 N_A_130_47#_M1010_g N_VPWR_c_663_n 0.0106914f $X=4.445 $Y=2.465 $X2=0
+ $Y2=0
cc_339 N_A_130_47#_M1011_g N_VPWR_c_663_n 0.0106914f $X=4.875 $Y=2.465 $X2=0
+ $Y2=0
cc_340 N_A_130_47#_M1012_g N_VPWR_c_663_n 0.0106914f $X=5.305 $Y=2.465 $X2=0
+ $Y2=0
cc_341 N_A_130_47#_M1013_g N_VPWR_c_663_n 0.0106914f $X=5.735 $Y=2.465 $X2=0
+ $Y2=0
cc_342 N_A_130_47#_M1022_g N_VPWR_c_663_n 0.0106914f $X=6.165 $Y=2.465 $X2=0
+ $Y2=0
cc_343 N_A_130_47#_M1025_g N_VPWR_c_663_n 0.0106914f $X=6.595 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A_130_47#_M1027_g N_VPWR_c_663_n 0.0106914f $X=7.025 $Y=2.465 $X2=0
+ $Y2=0
cc_345 N_A_130_47#_M1029_g N_VPWR_c_663_n 0.0106914f $X=7.455 $Y=2.465 $X2=0
+ $Y2=0
cc_346 N_A_130_47#_M1030_g N_VPWR_c_663_n 0.0106914f $X=7.885 $Y=2.465 $X2=0
+ $Y2=0
cc_347 N_A_130_47#_M1031_g N_VPWR_c_663_n 0.0106914f $X=8.315 $Y=2.465 $X2=0
+ $Y2=0
cc_348 N_A_130_47#_M1037_g N_VPWR_c_663_n 0.0106914f $X=8.745 $Y=2.465 $X2=0
+ $Y2=0
cc_349 N_A_130_47#_M1038_g N_VPWR_c_663_n 0.0105068f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_350 N_A_130_47#_M1041_g N_VPWR_c_663_n 0.0116957f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_351 N_A_130_47#_c_461_p N_VPWR_c_663_n 0.0100304f $X=0.79 $Y=2.025 $X2=0
+ $Y2=0
cc_352 N_A_130_47#_c_451_p N_VPWR_c_663_n 0.0100304f $X=1.65 $Y=2.025 $X2=0
+ $Y2=0
cc_353 N_A_130_47#_c_452_p N_VPWR_c_663_n 0.0100304f $X=2.51 $Y=2.025 $X2=0
+ $Y2=0
cc_354 N_A_130_47#_M1001_g N_X_c_862_n 0.00220648f $X=3.155 $Y=0.655 $X2=0 $Y2=0
cc_355 N_A_130_47#_c_319_n N_X_c_862_n 0.00182909f $X=3.155 $Y=1.725 $X2=0 $Y2=0
cc_356 N_A_130_47#_M1003_g N_X_c_862_n 0.00390855f $X=3.585 $Y=0.655 $X2=0 $Y2=0
cc_357 N_A_130_47#_c_320_n N_X_c_862_n 0.00197192f $X=3.585 $Y=1.725 $X2=0 $Y2=0
cc_358 N_A_130_47#_c_304_n N_X_c_862_n 0.0218339f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_359 N_A_130_47#_c_307_n N_X_c_862_n 0.0126612f $X=2.905 $Y=1.13 $X2=0 $Y2=0
cc_360 N_A_130_47#_c_339_n N_X_c_862_n 0.0100203f $X=2.905 $Y=1.84 $X2=0 $Y2=0
cc_361 N_A_130_47#_c_310_n N_X_c_862_n 0.0372715f $X=3 $Y=1.665 $X2=0 $Y2=0
cc_362 N_A_130_47#_c_311_n N_X_c_862_n 0.0268113f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_363 N_A_130_47#_c_312_n N_X_c_862_n 0.0295923f $X=3.8 $Y=1.49 $X2=0 $Y2=0
cc_364 N_A_130_47#_M1007_g N_X_c_863_n 0.00386542f $X=4.015 $Y=0.655 $X2=0 $Y2=0
cc_365 N_A_130_47#_M1006_g N_X_c_863_n 0.00247666f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_366 N_A_130_47#_M1014_g N_X_c_863_n 0.00386542f $X=4.445 $Y=0.655 $X2=0 $Y2=0
cc_367 N_A_130_47#_M1010_g N_X_c_863_n 0.00247666f $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A_130_47#_c_304_n N_X_c_863_n 0.0207982f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_369 N_A_130_47#_c_311_n N_X_c_863_n 0.0297586f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_370 N_A_130_47#_c_312_n N_X_c_863_n 0.0299092f $X=3.8 $Y=1.49 $X2=0 $Y2=0
cc_371 N_A_130_47#_c_313_n N_X_c_863_n 0.0299092f $X=4.66 $Y=1.49 $X2=0 $Y2=0
cc_372 N_A_130_47#_M1016_g N_X_c_864_n 0.00386542f $X=4.875 $Y=0.655 $X2=0 $Y2=0
cc_373 N_A_130_47#_M1011_g N_X_c_864_n 0.00247666f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A_130_47#_M1017_g N_X_c_864_n 0.00386542f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_375 N_A_130_47#_M1012_g N_X_c_864_n 0.00247666f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A_130_47#_c_304_n N_X_c_864_n 0.0207982f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_377 N_A_130_47#_c_311_n N_X_c_864_n 0.0297586f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_378 N_A_130_47#_c_313_n N_X_c_864_n 0.0299092f $X=4.66 $Y=1.49 $X2=0 $Y2=0
cc_379 N_A_130_47#_c_314_n N_X_c_864_n 0.0299092f $X=5.52 $Y=1.49 $X2=0 $Y2=0
cc_380 N_A_130_47#_M1018_g N_X_c_865_n 0.00386542f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_381 N_A_130_47#_M1013_g N_X_c_865_n 0.00247666f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_382 N_A_130_47#_M1019_g N_X_c_865_n 0.00386542f $X=6.165 $Y=0.655 $X2=0 $Y2=0
cc_383 N_A_130_47#_M1022_g N_X_c_865_n 0.00247666f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_384 N_A_130_47#_c_304_n N_X_c_865_n 0.0207982f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_385 N_A_130_47#_c_311_n N_X_c_865_n 0.0297586f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_386 N_A_130_47#_c_314_n N_X_c_865_n 0.0299092f $X=5.52 $Y=1.49 $X2=0 $Y2=0
cc_387 N_A_130_47#_c_315_n N_X_c_865_n 0.0299092f $X=6.38 $Y=1.49 $X2=0 $Y2=0
cc_388 N_A_130_47#_M1020_g N_X_c_866_n 0.00386542f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_389 N_A_130_47#_M1025_g N_X_c_866_n 0.00247666f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_390 N_A_130_47#_M1024_g N_X_c_866_n 0.00386542f $X=7.025 $Y=0.655 $X2=0 $Y2=0
cc_391 N_A_130_47#_M1027_g N_X_c_866_n 0.00247666f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_392 N_A_130_47#_c_304_n N_X_c_866_n 0.0207982f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_393 N_A_130_47#_c_311_n N_X_c_866_n 0.0297586f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_394 N_A_130_47#_c_315_n N_X_c_866_n 0.0299092f $X=6.38 $Y=1.49 $X2=0 $Y2=0
cc_395 N_A_130_47#_c_316_n N_X_c_866_n 0.0299092f $X=7.24 $Y=1.49 $X2=0 $Y2=0
cc_396 N_A_130_47#_M1026_g N_X_c_867_n 0.00386542f $X=7.455 $Y=0.655 $X2=0 $Y2=0
cc_397 N_A_130_47#_M1029_g N_X_c_867_n 0.00247666f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_398 N_A_130_47#_M1032_g N_X_c_867_n 0.00386542f $X=7.885 $Y=0.655 $X2=0 $Y2=0
cc_399 N_A_130_47#_M1030_g N_X_c_867_n 0.00247666f $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A_130_47#_c_304_n N_X_c_867_n 0.0207982f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_401 N_A_130_47#_c_311_n N_X_c_867_n 0.0297586f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_402 N_A_130_47#_c_316_n N_X_c_867_n 0.0299092f $X=7.24 $Y=1.49 $X2=0 $Y2=0
cc_403 N_A_130_47#_c_317_n N_X_c_867_n 0.0299092f $X=8.1 $Y=1.49 $X2=0 $Y2=0
cc_404 N_A_130_47#_M1034_g N_X_c_868_n 0.00386542f $X=8.315 $Y=0.655 $X2=0 $Y2=0
cc_405 N_A_130_47#_M1031_g N_X_c_868_n 0.00247666f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_406 N_A_130_47#_M1035_g N_X_c_868_n 0.00386542f $X=8.745 $Y=0.655 $X2=0 $Y2=0
cc_407 N_A_130_47#_M1037_g N_X_c_868_n 0.00247666f $X=8.745 $Y=2.465 $X2=0 $Y2=0
cc_408 N_A_130_47#_c_304_n N_X_c_868_n 0.0207982f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_409 N_A_130_47#_c_311_n N_X_c_868_n 0.0297039f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_410 N_A_130_47#_c_317_n N_X_c_868_n 0.0299092f $X=8.1 $Y=1.49 $X2=0 $Y2=0
cc_411 N_A_130_47#_c_318_n N_X_c_868_n 0.0299092f $X=8.96 $Y=1.49 $X2=0 $Y2=0
cc_412 N_A_130_47#_M1042_g N_X_c_869_n 0.00386542f $X=9.175 $Y=0.655 $X2=0 $Y2=0
cc_413 N_A_130_47#_M1038_g N_X_c_869_n 0.00264212f $X=9.175 $Y=2.465 $X2=0 $Y2=0
cc_414 N_A_130_47#_M1043_g N_X_c_869_n 0.00710182f $X=9.605 $Y=0.655 $X2=0 $Y2=0
cc_415 N_A_130_47#_c_304_n N_X_c_869_n 0.0308397f $X=9.605 $Y=1.655 $X2=0 $Y2=0
cc_416 N_A_130_47#_M1041_g N_X_c_869_n 0.00557757f $X=9.605 $Y=2.465 $X2=0 $Y2=0
cc_417 N_A_130_47#_c_311_n N_X_c_869_n 0.00701277f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_418 N_A_130_47#_c_318_n N_X_c_869_n 0.029223f $X=8.96 $Y=1.49 $X2=0 $Y2=0
cc_419 N_A_130_47#_c_319_n N_X_c_878_n 0.00291209f $X=3.155 $Y=1.725 $X2=0 $Y2=0
cc_420 N_A_130_47#_c_320_n N_X_c_878_n 0.00766908f $X=3.585 $Y=1.725 $X2=0 $Y2=0
cc_421 N_A_130_47#_M1006_g N_X_c_878_n 0.00766908f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_422 N_A_130_47#_M1010_g N_X_c_878_n 0.00766908f $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_423 N_A_130_47#_M1011_g N_X_c_878_n 0.00766908f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_424 N_A_130_47#_M1012_g N_X_c_878_n 0.00766908f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_425 N_A_130_47#_M1013_g N_X_c_878_n 0.00766908f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_426 N_A_130_47#_M1022_g N_X_c_878_n 0.00766908f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_427 N_A_130_47#_M1025_g N_X_c_878_n 0.00766908f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_428 N_A_130_47#_M1027_g N_X_c_878_n 0.00766908f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_429 N_A_130_47#_M1029_g N_X_c_878_n 0.00766908f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_430 N_A_130_47#_M1030_g N_X_c_878_n 0.00766908f $X=7.885 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A_130_47#_M1031_g N_X_c_878_n 0.00766908f $X=8.315 $Y=2.465 $X2=0 $Y2=0
cc_432 N_A_130_47#_M1037_g N_X_c_878_n 0.00766908f $X=8.745 $Y=2.465 $X2=0 $Y2=0
cc_433 N_A_130_47#_M1038_g N_X_c_878_n 0.0123908f $X=9.175 $Y=2.465 $X2=0 $Y2=0
cc_434 N_A_130_47#_M1041_g N_X_c_878_n 0.00197372f $X=9.605 $Y=2.465 $X2=0 $Y2=0
cc_435 N_A_130_47#_c_452_p N_X_c_878_n 0.00375391f $X=2.51 $Y=2.025 $X2=0 $Y2=0
cc_436 N_A_130_47#_c_311_n N_X_c_878_n 0.569124f $X=8.96 $Y=1.665 $X2=0 $Y2=0
cc_437 N_A_130_47#_c_312_n N_X_c_878_n 2.75984e-19 $X=3.8 $Y=1.49 $X2=0 $Y2=0
cc_438 N_A_130_47#_c_313_n N_X_c_878_n 2.75984e-19 $X=4.66 $Y=1.49 $X2=0 $Y2=0
cc_439 N_A_130_47#_c_314_n N_X_c_878_n 2.75984e-19 $X=5.52 $Y=1.49 $X2=0 $Y2=0
cc_440 N_A_130_47#_c_315_n N_X_c_878_n 2.75984e-19 $X=6.38 $Y=1.49 $X2=0 $Y2=0
cc_441 N_A_130_47#_c_316_n N_X_c_878_n 2.75984e-19 $X=7.24 $Y=1.49 $X2=0 $Y2=0
cc_442 N_A_130_47#_c_317_n N_X_c_878_n 2.75984e-19 $X=8.1 $Y=1.49 $X2=0 $Y2=0
cc_443 N_A_130_47#_c_318_n N_X_c_878_n 2.75984e-19 $X=8.96 $Y=1.49 $X2=0 $Y2=0
cc_444 N_A_130_47#_c_305_n N_VGND_M1009_d 0.00176461f $X=1.53 $Y=1.13 $X2=0
+ $Y2=0
cc_445 N_A_130_47#_c_368_n N_VGND_M1028_d 0.00333682f $X=2.415 $Y=0.95 $X2=0
+ $Y2=0
cc_446 N_A_130_47#_c_307_n N_VGND_M1039_d 0.00180544f $X=2.905 $Y=1.13 $X2=0
+ $Y2=0
cc_447 N_A_130_47#_c_305_n N_VGND_c_1050_n 0.0135055f $X=1.53 $Y=1.13 $X2=0
+ $Y2=0
cc_448 N_A_130_47#_c_368_n N_VGND_c_1051_n 0.0170777f $X=2.415 $Y=0.95 $X2=0
+ $Y2=0
cc_449 N_A_130_47#_M1001_g N_VGND_c_1052_n 0.00955801f $X=3.155 $Y=0.655 $X2=0
+ $Y2=0
cc_450 N_A_130_47#_M1003_g N_VGND_c_1052_n 6.60089e-19 $X=3.585 $Y=0.655 $X2=0
+ $Y2=0
cc_451 N_A_130_47#_c_307_n N_VGND_c_1052_n 0.0156506f $X=2.905 $Y=1.13 $X2=0
+ $Y2=0
cc_452 N_A_130_47#_M1003_g N_VGND_c_1053_n 0.00196442f $X=3.585 $Y=0.655 $X2=0
+ $Y2=0
cc_453 N_A_130_47#_M1007_g N_VGND_c_1053_n 0.00199892f $X=4.015 $Y=0.655 $X2=0
+ $Y2=0
cc_454 N_A_130_47#_c_304_n N_VGND_c_1053_n 7.55194e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_455 N_A_130_47#_c_311_n N_VGND_c_1053_n 0.00141255f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_456 N_A_130_47#_c_312_n N_VGND_c_1053_n 0.0120942f $X=3.8 $Y=1.49 $X2=0 $Y2=0
cc_457 N_A_130_47#_M1007_g N_VGND_c_1054_n 0.00585385f $X=4.015 $Y=0.655 $X2=0
+ $Y2=0
cc_458 N_A_130_47#_M1014_g N_VGND_c_1054_n 0.00585385f $X=4.445 $Y=0.655 $X2=0
+ $Y2=0
cc_459 N_A_130_47#_M1014_g N_VGND_c_1055_n 0.00199892f $X=4.445 $Y=0.655 $X2=0
+ $Y2=0
cc_460 N_A_130_47#_M1016_g N_VGND_c_1055_n 0.00199892f $X=4.875 $Y=0.655 $X2=0
+ $Y2=0
cc_461 N_A_130_47#_c_304_n N_VGND_c_1055_n 7.55194e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_462 N_A_130_47#_c_311_n N_VGND_c_1055_n 0.00141255f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_463 N_A_130_47#_c_313_n N_VGND_c_1055_n 0.0120942f $X=4.66 $Y=1.49 $X2=0
+ $Y2=0
cc_464 N_A_130_47#_M1017_g N_VGND_c_1056_n 0.00199892f $X=5.305 $Y=0.655 $X2=0
+ $Y2=0
cc_465 N_A_130_47#_M1018_g N_VGND_c_1056_n 0.00199892f $X=5.735 $Y=0.655 $X2=0
+ $Y2=0
cc_466 N_A_130_47#_c_304_n N_VGND_c_1056_n 7.55194e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_467 N_A_130_47#_c_311_n N_VGND_c_1056_n 0.00141255f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_468 N_A_130_47#_c_314_n N_VGND_c_1056_n 0.0120942f $X=5.52 $Y=1.49 $X2=0
+ $Y2=0
cc_469 N_A_130_47#_M1019_g N_VGND_c_1057_n 0.00199892f $X=6.165 $Y=0.655 $X2=0
+ $Y2=0
cc_470 N_A_130_47#_M1020_g N_VGND_c_1057_n 0.00199892f $X=6.595 $Y=0.655 $X2=0
+ $Y2=0
cc_471 N_A_130_47#_c_304_n N_VGND_c_1057_n 7.55194e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_472 N_A_130_47#_c_311_n N_VGND_c_1057_n 0.00141255f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_473 N_A_130_47#_c_315_n N_VGND_c_1057_n 0.0120942f $X=6.38 $Y=1.49 $X2=0
+ $Y2=0
cc_474 N_A_130_47#_M1024_g N_VGND_c_1058_n 0.00199892f $X=7.025 $Y=0.655 $X2=0
+ $Y2=0
cc_475 N_A_130_47#_M1026_g N_VGND_c_1058_n 0.00199892f $X=7.455 $Y=0.655 $X2=0
+ $Y2=0
cc_476 N_A_130_47#_c_304_n N_VGND_c_1058_n 7.55194e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_477 N_A_130_47#_c_311_n N_VGND_c_1058_n 0.00141255f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_478 N_A_130_47#_c_316_n N_VGND_c_1058_n 0.0120942f $X=7.24 $Y=1.49 $X2=0
+ $Y2=0
cc_479 N_A_130_47#_M1032_g N_VGND_c_1059_n 0.00199892f $X=7.885 $Y=0.655 $X2=0
+ $Y2=0
cc_480 N_A_130_47#_M1034_g N_VGND_c_1059_n 0.00199892f $X=8.315 $Y=0.655 $X2=0
+ $Y2=0
cc_481 N_A_130_47#_c_304_n N_VGND_c_1059_n 7.55194e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_482 N_A_130_47#_c_311_n N_VGND_c_1059_n 0.00141255f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_483 N_A_130_47#_c_317_n N_VGND_c_1059_n 0.0120942f $X=8.1 $Y=1.49 $X2=0 $Y2=0
cc_484 N_A_130_47#_M1034_g N_VGND_c_1060_n 0.00585385f $X=8.315 $Y=0.655 $X2=0
+ $Y2=0
cc_485 N_A_130_47#_M1035_g N_VGND_c_1060_n 0.00585385f $X=8.745 $Y=0.655 $X2=0
+ $Y2=0
cc_486 N_A_130_47#_M1035_g N_VGND_c_1061_n 0.00199892f $X=8.745 $Y=0.655 $X2=0
+ $Y2=0
cc_487 N_A_130_47#_M1042_g N_VGND_c_1061_n 0.00199892f $X=9.175 $Y=0.655 $X2=0
+ $Y2=0
cc_488 N_A_130_47#_c_304_n N_VGND_c_1061_n 7.55194e-19 $X=9.605 $Y=1.655 $X2=0
+ $Y2=0
cc_489 N_A_130_47#_c_311_n N_VGND_c_1061_n 0.00141255f $X=8.96 $Y=1.665 $X2=0
+ $Y2=0
cc_490 N_A_130_47#_c_318_n N_VGND_c_1061_n 0.0120942f $X=8.96 $Y=1.49 $X2=0
+ $Y2=0
cc_491 N_A_130_47#_M1043_g N_VGND_c_1063_n 0.00502529f $X=9.605 $Y=0.655 $X2=0
+ $Y2=0
cc_492 N_A_130_47#_c_626_p N_VGND_c_1064_n 0.00651381f $X=2.51 $Y=0.59 $X2=0
+ $Y2=0
cc_493 N_A_130_47#_M1001_g N_VGND_c_1066_n 0.00525069f $X=3.155 $Y=0.655 $X2=0
+ $Y2=0
cc_494 N_A_130_47#_M1003_g N_VGND_c_1066_n 0.00585385f $X=3.585 $Y=0.655 $X2=0
+ $Y2=0
cc_495 N_A_130_47#_M1018_g N_VGND_c_1068_n 0.00585385f $X=5.735 $Y=0.655 $X2=0
+ $Y2=0
cc_496 N_A_130_47#_M1019_g N_VGND_c_1068_n 0.00585385f $X=6.165 $Y=0.655 $X2=0
+ $Y2=0
cc_497 N_A_130_47#_M1020_g N_VGND_c_1070_n 0.00585385f $X=6.595 $Y=0.655 $X2=0
+ $Y2=0
cc_498 N_A_130_47#_M1024_g N_VGND_c_1070_n 0.00585385f $X=7.025 $Y=0.655 $X2=0
+ $Y2=0
cc_499 N_A_130_47#_M1026_g N_VGND_c_1072_n 0.00585385f $X=7.455 $Y=0.655 $X2=0
+ $Y2=0
cc_500 N_A_130_47#_M1032_g N_VGND_c_1072_n 0.00585385f $X=7.885 $Y=0.655 $X2=0
+ $Y2=0
cc_501 N_A_130_47#_c_635_p N_VGND_c_1074_n 0.00713515f $X=0.79 $Y=0.59 $X2=0
+ $Y2=0
cc_502 N_A_130_47#_c_636_p N_VGND_c_1075_n 0.00633629f $X=1.65 $Y=0.59 $X2=0
+ $Y2=0
cc_503 N_A_130_47#_M1016_g N_VGND_c_1076_n 0.00585385f $X=4.875 $Y=0.655 $X2=0
+ $Y2=0
cc_504 N_A_130_47#_M1017_g N_VGND_c_1076_n 0.00585385f $X=5.305 $Y=0.655 $X2=0
+ $Y2=0
cc_505 N_A_130_47#_M1042_g N_VGND_c_1077_n 0.00585385f $X=9.175 $Y=0.655 $X2=0
+ $Y2=0
cc_506 N_A_130_47#_M1043_g N_VGND_c_1077_n 0.00585385f $X=9.605 $Y=0.655 $X2=0
+ $Y2=0
cc_507 N_A_130_47#_M1005_s N_VGND_c_1083_n 0.00325821f $X=0.65 $Y=0.235 $X2=0
+ $Y2=0
cc_508 N_A_130_47#_M1023_s N_VGND_c_1083_n 0.00478158f $X=1.51 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_130_47#_M1036_s N_VGND_c_1083_n 0.00444305f $X=2.37 $Y=0.235 $X2=0
+ $Y2=0
cc_510 N_A_130_47#_M1001_g N_VGND_c_1083_n 0.00897288f $X=3.155 $Y=0.655 $X2=0
+ $Y2=0
cc_511 N_A_130_47#_M1003_g N_VGND_c_1083_n 0.0107375f $X=3.585 $Y=0.655 $X2=0
+ $Y2=0
cc_512 N_A_130_47#_M1007_g N_VGND_c_1083_n 0.0107375f $X=4.015 $Y=0.655 $X2=0
+ $Y2=0
cc_513 N_A_130_47#_M1014_g N_VGND_c_1083_n 0.0107375f $X=4.445 $Y=0.655 $X2=0
+ $Y2=0
cc_514 N_A_130_47#_M1016_g N_VGND_c_1083_n 0.0107375f $X=4.875 $Y=0.655 $X2=0
+ $Y2=0
cc_515 N_A_130_47#_M1017_g N_VGND_c_1083_n 0.0107375f $X=5.305 $Y=0.655 $X2=0
+ $Y2=0
cc_516 N_A_130_47#_M1018_g N_VGND_c_1083_n 0.0107375f $X=5.735 $Y=0.655 $X2=0
+ $Y2=0
cc_517 N_A_130_47#_M1019_g N_VGND_c_1083_n 0.0107375f $X=6.165 $Y=0.655 $X2=0
+ $Y2=0
cc_518 N_A_130_47#_M1020_g N_VGND_c_1083_n 0.0107375f $X=6.595 $Y=0.655 $X2=0
+ $Y2=0
cc_519 N_A_130_47#_M1024_g N_VGND_c_1083_n 0.0107375f $X=7.025 $Y=0.655 $X2=0
+ $Y2=0
cc_520 N_A_130_47#_M1026_g N_VGND_c_1083_n 0.0107375f $X=7.455 $Y=0.655 $X2=0
+ $Y2=0
cc_521 N_A_130_47#_M1032_g N_VGND_c_1083_n 0.0107375f $X=7.885 $Y=0.655 $X2=0
+ $Y2=0
cc_522 N_A_130_47#_M1034_g N_VGND_c_1083_n 0.0107375f $X=8.315 $Y=0.655 $X2=0
+ $Y2=0
cc_523 N_A_130_47#_M1035_g N_VGND_c_1083_n 0.0107375f $X=8.745 $Y=0.655 $X2=0
+ $Y2=0
cc_524 N_A_130_47#_M1042_g N_VGND_c_1083_n 0.0107375f $X=9.175 $Y=0.655 $X2=0
+ $Y2=0
cc_525 N_A_130_47#_M1043_g N_VGND_c_1083_n 0.0117419f $X=9.605 $Y=0.655 $X2=0
+ $Y2=0
cc_526 N_A_130_47#_c_635_p N_VGND_c_1083_n 0.00908616f $X=0.79 $Y=0.59 $X2=0
+ $Y2=0
cc_527 N_A_130_47#_c_636_p N_VGND_c_1083_n 0.00750004f $X=1.65 $Y=0.59 $X2=0
+ $Y2=0
cc_528 N_A_130_47#_c_626_p N_VGND_c_1083_n 0.00785222f $X=2.51 $Y=0.59 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_663_n N_X_M1002_s 0.00388669f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_530 N_VPWR_c_663_n N_X_M1006_s 0.003017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_531 N_VPWR_c_663_n N_X_M1011_s 0.003017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_532 N_VPWR_c_663_n N_X_M1013_s 0.003017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_533 N_VPWR_c_663_n N_X_M1025_s 0.003017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_534 N_VPWR_c_663_n N_X_M1029_s 0.003017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_535 N_VPWR_c_663_n N_X_M1031_s 0.003017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_536 N_VPWR_c_663_n N_X_M1038_s 0.003017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_c_668_n N_X_c_862_n 0.0365253f $X=2.94 $Y=2.26 $X2=0 $Y2=0
cc_538 N_VPWR_c_669_n N_X_c_862_n 0.00820875f $X=3.8 $Y=2.085 $X2=0 $Y2=0
cc_539 N_VPWR_c_684_n N_X_c_862_n 0.0140491f $X=3.67 $Y=3.33 $X2=0 $Y2=0
cc_540 N_VPWR_c_663_n N_X_c_862_n 0.0090585f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_541 N_VPWR_c_669_n N_X_c_863_n 0.00822181f $X=3.8 $Y=2.085 $X2=0 $Y2=0
cc_542 N_VPWR_c_670_n N_X_c_863_n 0.0149362f $X=4.53 $Y=3.33 $X2=0 $Y2=0
cc_543 N_VPWR_c_671_n N_X_c_863_n 0.00822181f $X=4.66 $Y=2.085 $X2=0 $Y2=0
cc_544 N_VPWR_c_663_n N_X_c_863_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_545 N_VPWR_c_671_n N_X_c_864_n 0.00822181f $X=4.66 $Y=2.085 $X2=0 $Y2=0
cc_546 N_VPWR_c_672_n N_X_c_864_n 0.00822181f $X=5.52 $Y=2.085 $X2=0 $Y2=0
cc_547 N_VPWR_c_693_n N_X_c_864_n 0.0149362f $X=5.39 $Y=3.33 $X2=0 $Y2=0
cc_548 N_VPWR_c_663_n N_X_c_864_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_549 N_VPWR_c_672_n N_X_c_865_n 0.00822181f $X=5.52 $Y=2.085 $X2=0 $Y2=0
cc_550 N_VPWR_c_673_n N_X_c_865_n 0.00822181f $X=6.38 $Y=2.085 $X2=0 $Y2=0
cc_551 N_VPWR_c_686_n N_X_c_865_n 0.0149362f $X=6.25 $Y=3.33 $X2=0 $Y2=0
cc_552 N_VPWR_c_663_n N_X_c_865_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_673_n N_X_c_866_n 0.00822181f $X=6.38 $Y=2.085 $X2=0 $Y2=0
cc_554 N_VPWR_c_674_n N_X_c_866_n 0.00822181f $X=7.24 $Y=2.085 $X2=0 $Y2=0
cc_555 N_VPWR_c_688_n N_X_c_866_n 0.0149362f $X=7.11 $Y=3.33 $X2=0 $Y2=0
cc_556 N_VPWR_c_663_n N_X_c_866_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_557 N_VPWR_c_674_n N_X_c_867_n 0.00822181f $X=7.24 $Y=2.085 $X2=0 $Y2=0
cc_558 N_VPWR_c_675_n N_X_c_867_n 0.00822181f $X=8.1 $Y=2.085 $X2=0 $Y2=0
cc_559 N_VPWR_c_690_n N_X_c_867_n 0.0149362f $X=7.97 $Y=3.33 $X2=0 $Y2=0
cc_560 N_VPWR_c_663_n N_X_c_867_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_561 N_VPWR_c_675_n N_X_c_868_n 0.00822181f $X=8.1 $Y=2.085 $X2=0 $Y2=0
cc_562 N_VPWR_c_676_n N_X_c_868_n 0.0149362f $X=8.83 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_c_677_n N_X_c_868_n 0.00822181f $X=8.96 $Y=2.085 $X2=0 $Y2=0
cc_564 N_VPWR_c_663_n N_X_c_868_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_565 N_VPWR_c_677_n N_X_c_869_n 0.00822181f $X=8.96 $Y=2.085 $X2=0 $Y2=0
cc_566 N_VPWR_c_694_n N_X_c_869_n 0.0149362f $X=9.69 $Y=3.33 $X2=0 $Y2=0
cc_567 N_VPWR_c_663_n N_X_c_869_n 0.0100304f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_568 N_VPWR_M1004_d N_X_c_878_n 0.00149321f $X=3.66 $Y=1.835 $X2=0 $Y2=0
cc_569 N_VPWR_M1010_d N_X_c_878_n 0.00149321f $X=4.52 $Y=1.835 $X2=0 $Y2=0
cc_570 N_VPWR_M1012_d N_X_c_878_n 0.00149321f $X=5.38 $Y=1.835 $X2=0 $Y2=0
cc_571 N_VPWR_M1022_d N_X_c_878_n 0.00149321f $X=6.24 $Y=1.835 $X2=0 $Y2=0
cc_572 N_VPWR_M1027_d N_X_c_878_n 0.00149321f $X=7.1 $Y=1.835 $X2=0 $Y2=0
cc_573 N_VPWR_M1030_d N_X_c_878_n 0.00149321f $X=7.96 $Y=1.835 $X2=0 $Y2=0
cc_574 N_VPWR_M1037_d N_X_c_878_n 0.00149321f $X=8.82 $Y=1.835 $X2=0 $Y2=0
cc_575 N_VPWR_c_668_n N_X_c_878_n 0.00167762f $X=2.94 $Y=2.26 $X2=0 $Y2=0
cc_576 N_VPWR_c_669_n N_X_c_878_n 0.025736f $X=3.8 $Y=2.085 $X2=0 $Y2=0
cc_577 N_VPWR_c_671_n N_X_c_878_n 0.025736f $X=4.66 $Y=2.085 $X2=0 $Y2=0
cc_578 N_VPWR_c_672_n N_X_c_878_n 0.025736f $X=5.52 $Y=2.085 $X2=0 $Y2=0
cc_579 N_VPWR_c_673_n N_X_c_878_n 0.025736f $X=6.38 $Y=2.085 $X2=0 $Y2=0
cc_580 N_VPWR_c_674_n N_X_c_878_n 0.025736f $X=7.24 $Y=2.085 $X2=0 $Y2=0
cc_581 N_VPWR_c_675_n N_X_c_878_n 0.025736f $X=8.1 $Y=2.085 $X2=0 $Y2=0
cc_582 N_VPWR_c_677_n N_X_c_878_n 0.025736f $X=8.96 $Y=2.085 $X2=0 $Y2=0
cc_583 N_VPWR_c_679_n N_X_c_878_n 0.00691659f $X=9.82 $Y=2.085 $X2=0 $Y2=0
cc_584 N_X_c_863_n N_VGND_c_1054_n 0.0149362f $X=4.23 $Y=0.47 $X2=0 $Y2=0
cc_585 N_X_c_868_n N_VGND_c_1060_n 0.0149362f $X=8.53 $Y=0.47 $X2=0 $Y2=0
cc_586 N_X_c_862_n N_VGND_c_1066_n 0.0140491f $X=3.37 $Y=0.47 $X2=0 $Y2=0
cc_587 N_X_c_865_n N_VGND_c_1068_n 0.0149362f $X=5.95 $Y=0.47 $X2=0 $Y2=0
cc_588 N_X_c_866_n N_VGND_c_1070_n 0.0149362f $X=6.81 $Y=0.47 $X2=0 $Y2=0
cc_589 N_X_c_867_n N_VGND_c_1072_n 0.0149362f $X=7.67 $Y=0.47 $X2=0 $Y2=0
cc_590 N_X_c_864_n N_VGND_c_1076_n 0.0149362f $X=5.09 $Y=0.47 $X2=0 $Y2=0
cc_591 N_X_c_869_n N_VGND_c_1077_n 0.0149362f $X=9.39 $Y=0.47 $X2=0 $Y2=0
cc_592 N_X_M1001_d N_VGND_c_1083_n 0.00388669f $X=3.23 $Y=0.235 $X2=0 $Y2=0
cc_593 N_X_M1007_d N_VGND_c_1083_n 0.003017f $X=4.09 $Y=0.235 $X2=0 $Y2=0
cc_594 N_X_M1016_d N_VGND_c_1083_n 0.003017f $X=4.95 $Y=0.235 $X2=0 $Y2=0
cc_595 N_X_M1018_d N_VGND_c_1083_n 0.003017f $X=5.81 $Y=0.235 $X2=0 $Y2=0
cc_596 N_X_M1020_d N_VGND_c_1083_n 0.003017f $X=6.67 $Y=0.235 $X2=0 $Y2=0
cc_597 N_X_M1026_d N_VGND_c_1083_n 0.003017f $X=7.53 $Y=0.235 $X2=0 $Y2=0
cc_598 N_X_M1034_d N_VGND_c_1083_n 0.003017f $X=8.39 $Y=0.235 $X2=0 $Y2=0
cc_599 N_X_M1042_d N_VGND_c_1083_n 0.003017f $X=9.25 $Y=0.235 $X2=0 $Y2=0
cc_600 N_X_c_862_n N_VGND_c_1083_n 0.0090585f $X=3.37 $Y=0.47 $X2=0 $Y2=0
cc_601 N_X_c_863_n N_VGND_c_1083_n 0.0100304f $X=4.23 $Y=0.47 $X2=0 $Y2=0
cc_602 N_X_c_864_n N_VGND_c_1083_n 0.0100304f $X=5.09 $Y=0.47 $X2=0 $Y2=0
cc_603 N_X_c_865_n N_VGND_c_1083_n 0.0100304f $X=5.95 $Y=0.47 $X2=0 $Y2=0
cc_604 N_X_c_866_n N_VGND_c_1083_n 0.0100304f $X=6.81 $Y=0.47 $X2=0 $Y2=0
cc_605 N_X_c_867_n N_VGND_c_1083_n 0.0100304f $X=7.67 $Y=0.47 $X2=0 $Y2=0
cc_606 N_X_c_868_n N_VGND_c_1083_n 0.0100304f $X=8.53 $Y=0.47 $X2=0 $Y2=0
cc_607 N_X_c_869_n N_VGND_c_1083_n 0.0100304f $X=9.39 $Y=0.47 $X2=0 $Y2=0
