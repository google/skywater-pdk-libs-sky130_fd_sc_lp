* File: sky130_fd_sc_lp__or3_m.pex.spice
* Created: Wed Sep  2 10:30:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3_M%C 3 5 7 8 9 12 14 15 16 17 22 24
c43 14 0 5.77736e-20 $X=0.667 $Y=1.435
r44 22 24 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.667 $Y=0.93
+ $X2=0.667 $Y2=0.765
r45 16 17 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=0.925
+ $X2=0.705 $Y2=1.295
r46 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=0.93 $X2=0.69 $Y2=0.93
r47 15 16 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=0.555
+ $X2=0.705 $Y2=0.925
r48 10 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.005 $Y=1.825
+ $X2=1.005 $Y2=2.195
r49 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=1.75
+ $X2=1.005 $Y2=1.825
r50 8 9 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=0.93 $Y=1.75 $X2=0.63
+ $Y2=1.75
r51 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.555 $Y=1.675
+ $X2=0.63 $Y2=1.75
r52 7 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.555 $Y=1.675
+ $X2=0.555 $Y2=1.435
r53 5 14 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.667 $Y=1.248
+ $X2=0.667 $Y2=1.435
r54 4 22 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.667 $Y=0.952
+ $X2=0.667 $Y2=0.93
r55 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.667 $Y=0.952
+ $X2=0.667 $Y2=1.248
r56 3 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.555 $Y=0.445
+ $X2=0.555 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_M%B 3 6 9 10 13 14 15 19
c44 6 0 1.35794e-19 $X=1.365 $Y=2.195
r45 14 15 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.215 $Y=0.925
+ $X2=1.215 $Y2=1.295
r46 14 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=0.93 $X2=1.23 $Y2=0.93
r47 12 19 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.23 $Y=1.285
+ $X2=1.23 $Y2=0.93
r48 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.252 $Y=1.285
+ $X2=1.252 $Y2=1.435
r49 10 19 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.23 $Y=0.915
+ $X2=1.23 $Y2=0.93
r50 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.252 $Y=0.765
+ $X2=1.252 $Y2=0.915
r51 6 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.365 $Y=2.195
+ $X2=1.365 $Y2=1.435
r52 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.365 $Y=0.445
+ $X2=1.365 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_M%A 3 7 11 12 13 16 17
r43 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.815
+ $Y=1.16 $X2=1.815 $Y2=1.16
r44 13 17 3.16609 $w=5.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.68 $Y=1.33
+ $X2=1.815 $Y2=1.33
r45 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.815 $Y=1.5
+ $X2=1.815 $Y2=1.16
r46 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.5
+ $X2=1.815 $Y2=1.665
r47 10 16 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=1.16
r48 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.795 $Y=0.445
+ $X2=1.795 $Y2=0.995
r49 3 12 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.725 $Y=2.195
+ $X2=1.725 $Y2=1.665
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_M%A_43_47# 1 2 3 10 14 17 20 22 23 26 28 32 37
+ 39 41 42 44 45 46 47
c96 22 0 5.77736e-20 $X=0.685 $Y=1.88
r97 43 44 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.245 $Y=0.895
+ $X2=2.245 $Y2=1.795
r98 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.16 $Y=0.81
+ $X2=2.245 $Y2=0.895
r99 41 42 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.16 $Y=0.81
+ $X2=1.685 $Y2=0.81
r100 40 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=1.88
+ $X2=1.46 $Y2=1.88
r101 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.16 $Y=1.88
+ $X2=2.245 $Y2=1.795
r102 39 40 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.16 $Y=1.88
+ $X2=1.625 $Y2=1.88
r103 35 42 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.59 $Y=0.725
+ $X2=1.685 $Y2=0.81
r104 35 37 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.59 $Y=0.725
+ $X2=1.59 $Y2=0.51
r105 33 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.46 $Y=2.94 $X2=1.46
+ $Y2=2.85
r106 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.46
+ $Y=2.94 $X2=1.46 $Y2=2.94
r107 30 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=1.965
+ $X2=1.46 $Y2=1.88
r108 30 32 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=1.46 $Y=1.965
+ $X2=1.46 $Y2=2.94
r109 29 45 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.895 $Y=1.88
+ $X2=0.79 $Y2=1.88
r110 28 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=1.88
+ $X2=1.46 $Y2=1.88
r111 28 29 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.295 $Y=1.88
+ $X2=0.895 $Y2=1.88
r112 24 45 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=1.965
+ $X2=0.79 $Y2=1.88
r113 24 26 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=1.965
+ $X2=0.79 $Y2=2.13
r114 22 45 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.685 $Y=1.88
+ $X2=0.79 $Y2=1.88
r115 22 23 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.685 $Y=1.88
+ $X2=0.425 $Y2=1.88
r116 18 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.33 $Y=1.795
+ $X2=0.425 $Y2=1.88
r117 18 20 75.0096 $w=1.88e-07 $l=1.285e-06 $layer=LI1_cond $X=0.33 $Y=1.795
+ $X2=0.33 $Y2=0.51
r118 14 17 897.34 $w=1.5e-07 $l=1.75e-06 $layer=POLY_cond $X=2.265 $Y=0.445
+ $X2=2.265 $Y2=2.195
r119 12 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.265 $Y=2.775
+ $X2=2.265 $Y2=2.195
r120 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=2.85
+ $X2=1.46 $Y2=2.85
r121 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.19 $Y=2.85
+ $X2=2.265 $Y2=2.775
r122 10 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.19 $Y=2.85
+ $X2=1.625 $Y2=2.85
r123 3 26 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.985 $X2=0.79 $Y2=2.13
r124 2 37 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.58 $Y2=0.51
r125 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.235 $X2=0.34 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_M%VPWR 1 6 9 10 11 21 22
c23 22 0 1.35794e-19 $X=2.64 $Y=3.33
r24 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r25 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r26 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r28 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r30 11 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 9 18 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r32 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.97 $Y2=3.33
r33 8 21 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=1.97 $Y2=3.33
r35 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=3.245 $X2=1.97
+ $Y2=3.33
r36 4 6 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=1.97 $Y=3.245
+ $X2=1.97 $Y2=2.26
r37 1 6 600 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=1.985 $X2=1.97 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_M%X 1 2 7 8 9 10 11 12 13 26 38 49
r23 49 50 7.00423 $w=4.08e-07 $l=1.05e-07 $layer=LI1_cond $X=2.52 $Y=2.26
+ $X2=2.52 $Y2=2.155
r24 36 38 1.26488 $w=4.08e-07 $l=4.5e-08 $layer=LI1_cond $X=2.52 $Y=2.36
+ $X2=2.52 $Y2=2.405
r25 23 26 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=0.485 $X2=2.64
+ $Y2=0.555
r26 12 36 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=2.52 $Y=2.34 $X2=2.52
+ $Y2=2.36
r27 12 49 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=2.52 $Y=2.34 $X2=2.52
+ $Y2=2.26
r28 12 13 9.83793 $w=4.08e-07 $l=3.5e-07 $layer=LI1_cond $X=2.52 $Y=2.425
+ $X2=2.52 $Y2=2.775
r29 12 38 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=2.52 $Y=2.425
+ $X2=2.52 $Y2=2.405
r30 11 50 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.64 $Y=2.035
+ $X2=2.64 $Y2=2.155
r31 10 11 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=2.035
r32 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.295 $X2=2.64
+ $Y2=1.665
r33 8 9 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=0.925 $X2=2.64
+ $Y2=1.295
r34 7 23 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.64 $Y=0.38 $X2=2.64
+ $Y2=0.485
r35 7 44 8.45022 $w=2.08e-07 $l=1.6e-07 $layer=LI1_cond $X=2.64 $Y=0.38 $X2=2.48
+ $Y2=0.38
r36 7 8 23.6824 $w=1.68e-07 $l=3.63e-07 $layer=LI1_cond $X=2.64 $Y=0.562
+ $X2=2.64 $Y2=0.925
r37 7 26 0.456684 $w=1.68e-07 $l=7e-09 $layer=LI1_cond $X=2.64 $Y=0.562 $X2=2.64
+ $Y2=0.555
r38 2 49 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.985 $X2=2.48 $Y2=2.26
r39 1 44 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.235 $X2=2.48 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_M%VGND 1 2 9 13 16 17 18 20 30 31 34
r45 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r47 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r48 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.15
+ $Y2=0
r50 25 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.68
+ $Y2=0
r51 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r52 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.15
+ $Y2=0
r54 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r55 18 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r56 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r57 16 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.68
+ $Y2=0
r58 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.01
+ $Y2=0
r59 15 30 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.64
+ $Y2=0
r60 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.01
+ $Y2=0
r61 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=0.085
+ $X2=2.01 $Y2=0
r62 11 13 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.01 $Y=0.085
+ $X2=2.01 $Y2=0.38
r63 7 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085 $X2=1.15
+ $Y2=0
r64 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.38
r65 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.87
+ $Y=0.235 $X2=2.01 $Y2=0.38
r66 1 9 182 $w=1.7e-07 $l=5.88048e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.235 $X2=1.15 $Y2=0.38
.ends

