* File: sky130_fd_sc_lp__a21bo_m.pex.spice
* Created: Wed Sep  2 09:19:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BO_M%A_80_72# 1 2 9 12 15 17 20 21 23 24 26 27 28
+ 29 34
c94 28 0 9.86124e-20 $X=1.91 $Y=1.71
c95 26 0 1.44532e-19 $X=1.805 $Y=2.335
c96 23 0 1.07508e-19 $X=1.7 $Y=2.42
c97 12 0 7.53516e-20 $X=0.577 $Y=1.968
r98 33 34 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.71 $Y=0.495
+ $X2=2.71 $Y2=1.625
r99 29 33 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.625 $Y=0.39
+ $X2=2.71 $Y2=0.495
r100 29 31 22.1818 $w=2.08e-07 $l=4.2e-07 $layer=LI1_cond $X=2.625 $Y=0.39
+ $X2=2.205 $Y2=0.39
r101 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.625 $Y=1.71
+ $X2=2.71 $Y2=1.625
r102 27 28 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.625 $Y=1.71
+ $X2=1.91 $Y2=1.71
r103 26 36 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=2.335
+ $X2=1.805 $Y2=2.42
r104 25 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.805 $Y=1.795
+ $X2=1.91 $Y2=1.71
r105 25 26 28.5195 $w=2.08e-07 $l=5.4e-07 $layer=LI1_cond $X=1.805 $Y=1.795
+ $X2=1.805 $Y2=2.335
r106 23 36 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.7 $Y=2.42
+ $X2=1.805 $Y2=2.42
r107 23 24 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=1.7 $Y=2.42
+ $X2=0.675 $Y2=2.42
r108 21 38 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.64
+ $X2=0.577 $Y2=1.475
r109 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.64 $X2=0.59 $Y2=1.64
r110 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=2.335
+ $X2=0.675 $Y2=2.42
r111 18 20 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.59 $Y=2.335
+ $X2=0.59 $Y2=1.64
r112 15 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.475 $Y=2.855
+ $X2=0.475 $Y2=2.145
r113 12 17 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.577 $Y=1.968
+ $X2=0.577 $Y2=2.145
r114 11 21 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=1.652
+ $X2=0.577 $Y2=1.64
r115 11 12 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.577 $Y=1.652
+ $X2=0.577 $Y2=1.968
r116 9 38 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=0.475 $Y=0.7
+ $X2=0.475 $Y2=1.475
r117 2 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=2.195 $X2=1.805 $Y2=2.34
r118 1 31 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.235 $X2=2.205 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%B1_N 1 3 4 6 8 12 16 19 20 21 22 27 28
c57 8 0 9.86124e-20 $X=1.11 $Y=2.385
r58 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=1.19
+ $X2=1.2 $Y2=1.19
r59 21 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.2
+ $Y2=2.035
r60 20 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r61 20 28 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.295
+ $X2=1.2 $Y2=1.19
r62 18 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.2 $Y=1.53 $X2=1.2
+ $Y2=1.19
r63 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.53 $X2=1.2
+ $Y2=1.695
r64 14 16 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.905 $Y=2.46
+ $X2=1.11 $Y2=2.46
r65 12 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.2 $Y=1.175 $X2=1.2
+ $Y2=1.19
r66 9 12 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.905 $Y=1.1 $X2=1.2
+ $Y2=1.1
r67 8 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.11 $Y=2.385
+ $X2=1.11 $Y2=2.46
r68 8 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.11 $Y=2.385
+ $X2=1.11 $Y2=1.695
r69 4 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.535
+ $X2=0.905 $Y2=2.46
r70 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=2.535
+ $X2=0.905 $Y2=2.855
r71 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.025
+ $X2=0.905 $Y2=1.1
r72 1 3 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.905 $Y=1.025
+ $X2=0.905 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%A_196_98# 1 2 10 12 13 14 17 18 20 24 29 30
+ 32 36 37 40 45 48
c76 32 0 6.783e-20 $X=1.705 $Y=0.76
c77 30 0 1.44532e-19 $X=1.57 $Y=2.94
c78 14 0 1.07508e-19 $X=1.775 $Y=2.01
r79 40 42 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=0.68 $X2=1.12
+ $Y2=0.76
r80 37 48 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=0.93
+ $X2=1.805 $Y2=0.765
r81 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.79
+ $Y=0.93 $X2=1.79 $Y2=0.93
r82 34 36 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=0.845
+ $X2=1.79 $Y2=0.93
r83 33 42 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.225 $Y=0.76
+ $X2=1.12 $Y2=0.76
r84 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=0.76
+ $X2=1.79 $Y2=0.845
r85 32 33 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.705 $Y=0.76
+ $X2=1.225 $Y2=0.76
r86 30 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=2.94
+ $X2=1.57 $Y2=2.775
r87 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=2.94 $X2=1.57 $Y2=2.94
r88 26 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=2.86
+ $X2=1.57 $Y2=2.86
r89 21 23 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.53 $Y=2.01 $X2=1.7
+ $Y2=2.01
r90 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.02 $Y=2.085
+ $X2=2.02 $Y2=2.405
r91 17 48 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.91 $Y=0.445
+ $X2=1.91 $Y2=0.765
r92 14 23 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.775 $Y=2.01
+ $X2=1.7 $Y2=2.01
r93 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.945 $Y=2.01
+ $X2=2.02 $Y2=2.085
r94 13 14 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.945 $Y=2.01
+ $X2=1.775 $Y2=2.01
r95 12 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.7 $Y=1.935 $X2=1.7
+ $Y2=2.01
r96 12 24 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.7 $Y=1.935 $X2=1.7
+ $Y2=1.435
r97 10 24 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.805 $Y=1.255
+ $X2=1.805 $Y2=1.435
r98 9 37 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.805 $Y=0.945
+ $X2=1.805 $Y2=0.93
r99 9 10 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.805 $Y=0.945
+ $X2=1.805 $Y2=1.255
r100 7 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.53 $Y=2.085
+ $X2=1.53 $Y2=2.01
r101 7 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.53 $Y=2.085
+ $X2=1.53 $Y2=2.775
r102 2 26 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.645 $X2=1.12 $Y2=2.86
r103 1 40 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.49 $X2=1.12 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%A1 3 6 9 10 11 12 13 17
c43 17 0 6.783e-20 $X=2.36 $Y=0.93
r44 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.36
+ $Y=0.93 $X2=2.36 $Y2=0.93
r45 13 18 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.26 $Y=1.295
+ $X2=2.26 $Y2=0.93
r46 12 18 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=2.26 $Y=0.925
+ $X2=2.26 $Y2=0.93
r47 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.36 $Y=1.27
+ $X2=2.36 $Y2=0.93
r48 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.27
+ $X2=2.36 $Y2=1.435
r49 9 17 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=0.765
+ $X2=2.36 $Y2=0.93
r50 6 11 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.45 $Y=2.405
+ $X2=2.45 $Y2=1.435
r51 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.42 $Y=0.445 $X2=2.42
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%A2 3 7 11 13 14 15 16 21
r36 15 16 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.665
r37 14 15 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=0.925
+ $X2=3.09 $Y2=1.295
r38 14 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.06
+ $Y=1.005 $X2=3.06 $Y2=1.005
r39 12 21 39.0632 $w=4.2e-07 $l=2.95e-07 $layer=POLY_cond $X=3.015 $Y=1.3
+ $X2=3.015 $Y2=1.005
r40 12 13 52.1105 $w=4.2e-07 $l=2.1e-07 $layer=POLY_cond $X=3.015 $Y=1.3
+ $X2=3.015 $Y2=1.51
r41 11 21 1.98626 $w=4.2e-07 $l=1.5e-08 $layer=POLY_cond $X=3.015 $Y=0.99
+ $X2=3.015 $Y2=1.005
r42 10 11 44.1654 $w=4.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.98 $Y=0.84
+ $X2=2.98 $Y2=0.99
r43 7 13 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=2.88 $Y=2.405
+ $X2=2.88 $Y2=1.51
r44 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.81 $Y=0.445
+ $X2=2.81 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%X 1 2 7 8 9 10 11 12 13
r12 13 39 5.18812 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=0.26 $Y=2.775 $X2=0.26
+ $Y2=2.685
r13 12 39 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.685
r14 11 12 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r15 10 11 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r16 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295 $X2=0.24
+ $Y2=1.665
r17 8 9 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925 $X2=0.24
+ $Y2=1.295
r18 8 37 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.8
r19 7 37 13.3743 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=0.26 $Y=0.555
+ $X2=0.26 $Y2=0.8
r20 2 13 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.645 $X2=0.26 $Y2=2.85
r21 1 7 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.49 $X2=0.26 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%VPWR 1 2 9 11 15 17 19 26 27 30 33
r39 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 27 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 24 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.665 $Y2=3.33
r44 24 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 19 30 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.69 $Y2=3.33
r48 19 21 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 17 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 13 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=3.245
+ $X2=2.665 $Y2=3.33
r52 13 15 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=2.665 $Y=3.245
+ $X2=2.665 $Y2=2.49
r53 12 30 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.69 $Y2=3.33
r54 11 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.665 $Y2=3.33
r55 11 12 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=0.795 $Y2=3.33
r56 7 30 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r57 7 9 17.1645 $w=2.08e-07 $l=3.25e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.92
r58 2 15 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=2.195 $X2=2.665 $Y2=2.49
r59 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.645 $X2=0.69 $Y2=2.92
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%A_419_439# 1 2 9 11 12 15
r19 13 15 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=3.095 $Y=2.145
+ $X2=3.095 $Y2=2.34
r20 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.99 $Y=2.06
+ $X2=3.095 $Y2=2.145
r21 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.99 $Y=2.06
+ $X2=2.34 $Y2=2.06
r22 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.235 $Y=2.145
+ $X2=2.34 $Y2=2.06
r23 7 9 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=2.235 $Y=2.145
+ $X2=2.235 $Y2=2.34
r24 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=2.195 $X2=3.095 $Y2=2.34
r25 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=2.195 $X2=2.235 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_M%VGND 1 2 3 12 16 18 20 23 24 25 31 35 41 45
r48 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r50 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.695
+ $Y2=0
r52 36 38 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.64
+ $Y2=0
r53 35 44 3.51344 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.167
+ $Y2=0
r54 35 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=2.64
+ $Y2=0
r55 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 31 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.695
+ $Y2=0
r57 31 33 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.2
+ $Y2=0
r58 29 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r59 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 25 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r61 25 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r62 25 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r63 23 28 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r64 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.69
+ $Y2=0
r65 22 33 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r66 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.69
+ $Y2=0
r67 18 44 3.33045 $w=1.9e-07 $l=1.32868e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.167 $Y2=0
r68 18 20 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.38
r69 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0
r70 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0.38
r71 10 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r72 10 12 29.0476 $w=2.08e-07 $l=5.5e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.635
r73 3 20 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.235 $X2=3.06 $Y2=0.38
r74 2 16 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.235 $X2=1.695 $Y2=0.38
r75 1 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.49 $X2=0.69 $Y2=0.635
.ends

