* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_lp2 A0 A1 S VGND VNB VPB VPWR X
X0 a_84_259# A1 a_590_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_349_57# A0 a_84_259# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_306_401# A1 a_84_259# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VPWR S a_182_303# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_84_259# A0 a_518_401# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_518_401# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_115_57# a_84_259# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_84_259# a_115_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_776_57# S a_182_303# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_590_57# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 X a_84_259# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VPWR a_182_303# a_306_401# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 VGND a_182_303# a_349_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND S a_776_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
