* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfstp_lp CLK D SET_B VGND VNB VPB VPWR Q
X0 a_904_125# a_943_321# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_2287_74# a_1526_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_1256_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1731_99# a_1526_125# a_2104_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_2374_74# a_1526_125# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_2287_74# a_2532_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_135_409# a_479_409# a_709_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_531_109# a_266_409# a_479_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_709_419# a_479_409# a_904_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_709_419# a_1448_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1731_99# a_1526_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_2532_74# a_2287_74# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_266_409# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_1526_125# a_266_409# a_1683_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_709_419# a_943_321# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 VPWR D a_135_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_2287_74# a_1526_125# a_2374_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1726_419# a_1731_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X18 a_135_409# a_266_409# a_709_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1683_125# a_1731_99# a_1761_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_709_419# a_1448_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_1761_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1526_125# a_479_409# a_1726_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X23 a_373_109# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_2287_74# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_1448_419# a_266_409# a_1526_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 VPWR SET_B a_1526_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 a_709_419# a_266_409# a_881_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 a_2104_47# a_1526_125# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR a_266_409# a_479_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X30 a_266_409# CLK a_373_109# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_881_419# a_943_321# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 VGND a_266_409# a_531_109# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_943_321# a_709_419# a_1256_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_943_321# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X35 a_110_57# D a_135_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VGND D a_110_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_1448_125# a_479_409# a_1526_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
