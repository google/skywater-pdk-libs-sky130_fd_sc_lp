* File: sky130_fd_sc_lp__maj3_0.pex.spice
* Created: Fri Aug 28 10:42:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MAJ3_0%A 1 3 6 9 12 16 20 22 23 27 28
r49 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.07 $X2=1.35 $Y2=1.07
r50 23 28 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.2 $Y=1.24 $X2=1.35
+ $Y2=1.24
r51 22 23 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.24 $X2=1.2
+ $Y2=1.24
r52 18 20 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=0.86 $Y=1.97 $X2=1.06
+ $Y2=1.97
r53 14 27 85.6701 $w=2.93e-07 $l=6.09241e-07 $layer=POLY_cond $X=1.52 $Y=1.575
+ $X2=1.29 $Y2=1.07
r54 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.52 $Y=1.575
+ $X2=1.52 $Y2=2.365
r55 10 27 29.7384 $w=2.93e-07 $l=2.70185e-07 $layer=POLY_cond $X=1.49 $Y=0.905
+ $X2=1.29 $Y2=1.07
r56 10 12 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.49 $Y=0.905
+ $X2=1.49 $Y2=0.495
r57 9 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.06 $Y=1.895
+ $X2=1.06 $Y2=1.97
r58 8 27 85.6701 $w=2.93e-07 $l=6.09241e-07 $layer=POLY_cond $X=1.06 $Y=1.575
+ $X2=1.29 $Y2=1.07
r59 8 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.06 $Y=1.575 $X2=1.06
+ $Y2=1.895
r60 4 27 29.7384 $w=2.93e-07 $l=3.01413e-07 $layer=POLY_cond $X=1.06 $Y=0.905
+ $X2=1.29 $Y2=1.07
r61 4 6 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.06 $Y=0.905 $X2=1.06
+ $Y2=0.495
r62 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.86 $Y=2.045
+ $X2=0.86 $Y2=1.97
r63 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.86 $Y=2.045 $X2=0.86
+ $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_0%B 3 7 11 15 17 18 22
r46 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.21
+ $Y=1.07 $X2=2.21 $Y2=1.07
r47 18 23 7.67632 $w=6.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.64 $Y=1.24
+ $X2=2.21 $Y2=1.24
r48 17 23 0.892596 $w=6.68e-07 $l=5e-08 $layer=LI1_cond $X=2.16 $Y=1.24 $X2=2.21
+ $Y2=1.24
r49 13 22 86.458 $w=2.9e-07 $l=6.02993e-07 $layer=POLY_cond $X=2.31 $Y=1.575
+ $X2=2.095 $Y2=1.07
r50 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.31 $Y=1.575
+ $X2=2.31 $Y2=2.365
r51 9 22 29.9477 $w=2.9e-07 $l=2.85832e-07 $layer=POLY_cond $X=2.31 $Y=0.905
+ $X2=2.095 $Y2=1.07
r52 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.31 $Y=0.905
+ $X2=2.31 $Y2=0.495
r53 5 22 86.458 $w=2.9e-07 $l=6.02993e-07 $layer=POLY_cond $X=1.88 $Y=1.575
+ $X2=2.095 $Y2=1.07
r54 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.88 $Y=1.575 $X2=1.88
+ $Y2=2.365
r55 1 22 29.9477 $w=2.9e-07 $l=2.15e-07 $layer=POLY_cond $X=1.88 $Y=1.07
+ $X2=2.095 $Y2=1.07
r56 1 3 210.234 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.88 $Y=1.07 $X2=1.88
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_0%C 4 5 6 9 13 16 19 21 24
c59 21 0 1.64375e-19 $X=2.64 $Y=2.775
c60 13 0 1.65452e-19 $X=2.67 $Y=0.495
r61 24 27 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.76 $Y=2.9 $X2=2.76
+ $Y2=3.02
r62 24 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=2.9
+ $X2=2.76 $Y2=2.735
r63 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=2.9 $X2=2.76 $Y2=2.9
r64 21 25 3.60138 $w=3.98e-07 $l=1.25e-07 $layer=LI1_cond $X=2.725 $Y=2.775
+ $X2=2.725 $Y2=2.9
r65 17 19 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.5 $Y=1.58 $X2=0.67
+ $Y2=1.58
r66 16 26 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.67 $Y=2.365
+ $X2=2.67 $Y2=2.735
r67 13 16 958.872 $w=1.5e-07 $l=1.87e-06 $layer=POLY_cond $X=2.67 $Y=0.495
+ $X2=2.67 $Y2=2.365
r68 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.67 $Y=1.505
+ $X2=0.67 $Y2=1.58
r69 7 9 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.67 $Y=1.505
+ $X2=0.67 $Y2=0.495
r70 5 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.595 $Y=3.02
+ $X2=2.76 $Y2=3.02
r71 5 6 1035.79 $w=1.5e-07 $l=2.02e-06 $layer=POLY_cond $X=2.595 $Y=3.02
+ $X2=0.575 $Y2=3.02
r72 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.5 $Y=2.945
+ $X2=0.575 $Y2=3.02
r73 2 4 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.5 $Y=2.945 $X2=0.5
+ $Y2=2.365
r74 1 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.5 $Y=1.655 $X2=0.5
+ $Y2=1.58
r75 1 4 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.5 $Y=1.655 $X2=0.5
+ $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_0%A_28_431# 1 2 3 4 14 17 21 23 25 28 30 33 36
+ 38 39 42 43 48 50 54
c101 43 0 9.18356e-20 $X=3.12 $Y=1.27
c102 21 0 1.64375e-19 $X=3.22 $Y=2.255
r103 51 54 8.19054 $w=4.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.78 $Y=0.495
+ $X2=2.095 $Y2=0.495
r104 45 48 6.50043 $w=4.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.205 $Y=0.495
+ $X2=0.455 $Y2=0.495
r105 43 59 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.27
+ $X2=3.125 $Y2=1.105
r106 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.12
+ $Y=1.27 $X2=3.12 $Y2=1.27
r107 40 42 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.12 $Y=1.755
+ $X2=3.12 $Y2=1.27
r108 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.955 $Y=1.84
+ $X2=3.12 $Y2=1.755
r109 38 39 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.955 $Y=1.84
+ $X2=2.26 $Y2=1.84
r110 34 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=1.84
+ $X2=2.26 $Y2=1.84
r111 34 56 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.095 $Y=1.84
+ $X2=1.78 $Y2=1.84
r112 34 36 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.095 $Y=1.925
+ $X2=2.095 $Y2=2.365
r113 33 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=1.755
+ $X2=1.78 $Y2=1.84
r114 32 51 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.78 $Y=0.725
+ $X2=1.78 $Y2=0.495
r115 32 33 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=1.78 $Y=0.725
+ $X2=1.78 $Y2=1.755
r116 31 50 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=1.84
+ $X2=0.285 $Y2=1.84
r117 30 56 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=1.84
+ $X2=1.78 $Y2=1.84
r118 30 31 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=1.695 $Y=1.84
+ $X2=0.45 $Y2=1.84
r119 26 50 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=1.925
+ $X2=0.285 $Y2=1.84
r120 26 28 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.285 $Y=1.925
+ $X2=0.285 $Y2=2.365
r121 25 50 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.205 $Y=1.755
+ $X2=0.285 $Y2=1.84
r122 24 45 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.205 $Y=0.725
+ $X2=0.205 $Y2=0.495
r123 24 25 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.205 $Y=0.725
+ $X2=0.205 $Y2=1.755
r124 21 23 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.22 $Y=2.255
+ $X2=3.22 $Y2=1.775
r125 17 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.1 $Y=0.495
+ $X2=3.1 $Y2=1.105
r126 14 23 47.1551 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=3.125 $Y=1.605
+ $X2=3.125 $Y2=1.775
r127 13 43 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=3.125 $Y=1.275
+ $X2=3.125 $Y2=1.27
r128 13 14 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=3.125 $Y=1.275
+ $X2=3.125 $Y2=1.605
r129 4 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=2.155 $X2=2.095 $Y2=2.365
r130 3 28 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=2.155 $X2=0.285 $Y2=2.365
r131 2 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.285 $X2=2.095 $Y2=0.495
r132 1 48 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.285 $X2=0.455 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_0%VPWR 1 2 9 12 16 18 20 25 32 33 36 39
r50 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r54 30 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.19 $Y2=3.33
r55 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.19 $Y2=3.33
r59 26 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 25 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=3.19 $Y2=3.33
r61 25 28 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 23 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 20 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.19 $Y2=3.33
r65 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 18 40 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 18 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 14 16 5.68539 $w=3.73e-07 $l=1.85e-07 $layer=LI1_cond $X=3.005 $Y=2.292
+ $X2=3.19 $Y2=2.292
r69 12 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=3.245
+ $X2=3.19 $Y2=3.33
r70 11 16 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.19 $Y=2.48
+ $X2=3.19 $Y2=2.292
r71 11 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.19 $Y=2.48
+ $X2=3.19 $Y2=3.245
r72 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245 $X2=1.19
+ $Y2=3.33
r73 7 9 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=1.19 $Y=3.245 $X2=1.19
+ $Y2=2.365
r74 2 14 600 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.155 $X2=3.005 $Y2=2.29
r75 1 9 600 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.155 $X2=1.19 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_0%X 1 2 10 13 14 15
c17 10 0 1.65452e-19 $X=3.59 $Y=0.495
r18 14 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=2.035
r19 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.59 $Y=1.295
+ $X2=3.59 $Y2=1.665
r20 11 13 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=3.59 $Y=0.725
+ $X2=3.59 $Y2=1.295
r21 10 11 4.30706 $w=2.5e-07 $l=2.3e-07 $layer=LI1_cond $X=3.59 $Y=0.495
+ $X2=3.59 $Y2=0.725
r22 8 10 7.15047 $w=4.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.315 $Y=0.495
+ $X2=3.59 $Y2=0.495
r23 2 15 300 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=2 $X=3.295
+ $Y=1.935 $X2=3.55 $Y2=2.08
r24 1 8 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.285 $X2=3.315 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_0%VGND 1 2 9 13 16 17 18 20 33 34 37
c43 13 0 9.18356e-20 $X=2.885 $Y=0.495
r44 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r46 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r47 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.275
+ $Y2=0
r52 25 27 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r53 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r54 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=0 $X2=1.275
+ $Y2=0
r56 20 22 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.11 $Y=0 $X2=0.72
+ $Y2=0
r57 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r58 18 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r59 16 30 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.64
+ $Y2=0
r60 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.845
+ $Y2=0
r61 15 33 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=3.6
+ $Y2=0
r62 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.845
+ $Y2=0
r63 11 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0
r64 11 13 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0.495
r65 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=0.085
+ $X2=1.275 $Y2=0
r66 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.275 $Y=0.085
+ $X2=1.275 $Y2=0.495
r67 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.285 $X2=2.885 $Y2=0.495
r68 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.135
+ $Y=0.285 $X2=1.275 $Y2=0.495
.ends

