* File: sky130_fd_sc_lp__o221ai_4.pxi.spice
* Created: Fri Aug 28 11:08:46 2020
* 
x_PM_SKY130_FD_SC_LP__O221AI_4%C1 N_C1_M1005_g N_C1_M1018_g N_C1_M1001_g
+ N_C1_M1021_g N_C1_M1004_g N_C1_M1032_g N_C1_M1010_g N_C1_M1024_g C1 C1 C1 C1
+ C1 N_C1_c_139_n PM_SKY130_FD_SC_LP__O221AI_4%C1
x_PM_SKY130_FD_SC_LP__O221AI_4%B1 N_B1_M1002_g N_B1_M1011_g N_B1_M1003_g
+ N_B1_M1023_g N_B1_M1015_g N_B1_M1026_g N_B1_M1019_g N_B1_M1036_g N_B1_c_223_n
+ N_B1_c_224_n N_B1_c_225_n B1 N_B1_c_226_n N_B1_c_227_n N_B1_c_228_n
+ PM_SKY130_FD_SC_LP__O221AI_4%B1
x_PM_SKY130_FD_SC_LP__O221AI_4%B2 N_B2_c_344_n N_B2_M1012_g N_B2_M1006_g
+ N_B2_c_346_n N_B2_M1013_g N_B2_M1014_g N_B2_c_348_n N_B2_M1030_g N_B2_M1020_g
+ N_B2_c_350_n N_B2_M1031_g N_B2_M1037_g B2 B2 B2 N_B2_c_353_n
+ PM_SKY130_FD_SC_LP__O221AI_4%B2
x_PM_SKY130_FD_SC_LP__O221AI_4%A1 N_A1_M1007_g N_A1_M1016_g N_A1_c_429_n
+ N_A1_M1022_g N_A1_M1017_g N_A1_c_431_n N_A1_M1027_g N_A1_M1029_g N_A1_c_433_n
+ N_A1_M1035_g N_A1_M1033_g N_A1_c_435_n N_A1_c_436_n N_A1_c_437_n N_A1_c_438_n
+ A1 A1 A1 N_A1_c_440_n N_A1_c_441_n PM_SKY130_FD_SC_LP__O221AI_4%A1
x_PM_SKY130_FD_SC_LP__O221AI_4%A2 N_A2_M1009_g N_A2_M1000_g N_A2_M1025_g
+ N_A2_M1008_g N_A2_M1038_g N_A2_M1028_g N_A2_M1039_g N_A2_M1034_g A2 A2 A2
+ N_A2_c_543_n N_A2_c_544_n PM_SKY130_FD_SC_LP__O221AI_4%A2
x_PM_SKY130_FD_SC_LP__O221AI_4%VPWR N_VPWR_M1001_d N_VPWR_M1004_d N_VPWR_M1024_d
+ N_VPWR_M1023_d N_VPWR_M1036_d N_VPWR_M1017_s N_VPWR_M1033_s N_VPWR_c_622_n
+ N_VPWR_c_623_n N_VPWR_c_624_n N_VPWR_c_625_n N_VPWR_c_626_n N_VPWR_c_627_n
+ N_VPWR_c_628_n N_VPWR_c_629_n N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_632_n
+ N_VPWR_c_633_n N_VPWR_c_634_n VPWR N_VPWR_c_635_n N_VPWR_c_636_n
+ N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n N_VPWR_c_641_n
+ N_VPWR_c_642_n N_VPWR_c_621_n PM_SKY130_FD_SC_LP__O221AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O221AI_4%Y N_Y_M1005_d N_Y_M1021_d N_Y_M1001_s N_Y_M1010_s
+ N_Y_M1006_s N_Y_M1020_s N_Y_M1000_d N_Y_M1028_d N_Y_c_771_n N_Y_c_765_n
+ N_Y_c_766_n N_Y_c_782_n N_Y_c_858_n N_Y_c_784_n N_Y_c_767_n N_Y_c_860_n
+ N_Y_c_768_n N_Y_c_807_n N_Y_c_812_n N_Y_c_837_n N_Y_c_769_n N_Y_c_796_n
+ N_Y_c_800_n N_Y_c_814_n N_Y_c_816_n N_Y_c_840_n Y Y N_Y_c_833_n N_Y_c_834_n
+ PM_SKY130_FD_SC_LP__O221AI_4%Y
x_PM_SKY130_FD_SC_LP__O221AI_4%A_592_367# N_A_592_367#_M1011_s
+ N_A_592_367#_M1026_s N_A_592_367#_M1014_d N_A_592_367#_M1037_d
+ N_A_592_367#_c_906_n N_A_592_367#_c_937_n N_A_592_367#_c_910_n
+ N_A_592_367#_c_922_n N_A_592_367#_c_940_n N_A_592_367#_c_908_n
+ N_A_592_367#_c_909_n N_A_592_367#_c_928_n N_A_592_367#_c_930_n
+ PM_SKY130_FD_SC_LP__O221AI_4%A_592_367#
x_PM_SKY130_FD_SC_LP__O221AI_4%A_1317_367# N_A_1317_367#_M1016_d
+ N_A_1317_367#_M1008_s N_A_1317_367#_M1034_s N_A_1317_367#_M1029_d
+ N_A_1317_367#_c_947_n N_A_1317_367#_c_956_n N_A_1317_367#_c_948_n
+ N_A_1317_367#_c_987_n N_A_1317_367#_c_958_n N_A_1317_367#_c_973_n
+ N_A_1317_367#_c_960_n N_A_1317_367#_c_945_n N_A_1317_367#_c_946_n
+ N_A_1317_367#_c_978_n N_A_1317_367#_c_980_n
+ PM_SKY130_FD_SC_LP__O221AI_4%A_1317_367#
x_PM_SKY130_FD_SC_LP__O221AI_4%A_29_65# N_A_29_65#_M1005_s N_A_29_65#_M1018_s
+ N_A_29_65#_M1032_s N_A_29_65#_M1002_s N_A_29_65#_M1015_s N_A_29_65#_M1013_d
+ N_A_29_65#_M1031_d N_A_29_65#_c_991_n N_A_29_65#_c_992_n N_A_29_65#_c_993_n
+ N_A_29_65#_c_1005_n N_A_29_65#_c_994_n N_A_29_65#_c_995_n N_A_29_65#_c_996_n
+ N_A_29_65#_c_997_n N_A_29_65#_c_998_n N_A_29_65#_c_999_n N_A_29_65#_c_1022_n
+ N_A_29_65#_c_1024_n PM_SKY130_FD_SC_LP__O221AI_4%A_29_65#
x_PM_SKY130_FD_SC_LP__O221AI_4%A_509_47# N_A_509_47#_M1002_d N_A_509_47#_M1003_d
+ N_A_509_47#_M1012_s N_A_509_47#_M1030_s N_A_509_47#_M1019_d
+ N_A_509_47#_M1009_s N_A_509_47#_M1038_s N_A_509_47#_M1022_s
+ N_A_509_47#_M1035_s N_A_509_47#_c_1084_n N_A_509_47#_c_1098_n
+ N_A_509_47#_c_1100_n N_A_509_47#_c_1090_n N_A_509_47#_c_1159_p
+ N_A_509_47#_c_1091_n N_A_509_47#_c_1107_n N_A_509_47#_c_1153_p
+ N_A_509_47#_c_1111_n N_A_509_47#_c_1164_p N_A_509_47#_c_1112_n
+ N_A_509_47#_c_1167_p N_A_509_47#_c_1085_n N_A_509_47#_c_1086_n
+ N_A_509_47#_c_1094_n N_A_509_47#_c_1097_n N_A_509_47#_c_1119_n
+ N_A_509_47#_c_1120_n N_A_509_47#_c_1121_n
+ PM_SKY130_FD_SC_LP__O221AI_4%A_509_47#
x_PM_SKY130_FD_SC_LP__O221AI_4%VGND N_VGND_M1007_d N_VGND_M1025_d N_VGND_M1039_d
+ N_VGND_M1027_d N_VGND_c_1190_n N_VGND_c_1191_n N_VGND_c_1192_n N_VGND_c_1193_n
+ N_VGND_c_1194_n N_VGND_c_1195_n N_VGND_c_1196_n VGND N_VGND_c_1197_n
+ N_VGND_c_1198_n N_VGND_c_1199_n N_VGND_c_1200_n N_VGND_c_1201_n
+ N_VGND_c_1202_n N_VGND_c_1203_n PM_SKY130_FD_SC_LP__O221AI_4%VGND
cc_1 VNB N_C1_M1005_g 0.0265735f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.745
cc_2 VNB N_C1_M1018_g 0.0199436f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.745
cc_3 VNB N_C1_M1021_g 0.0208847f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.745
cc_4 VNB N_C1_M1032_g 0.0245347f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.745
cc_5 VNB C1 0.0116226f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_6 VNB N_C1_c_139_n 0.119725f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=1.51
cc_7 VNB N_B1_M1002_g 0.0277968f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.745
cc_8 VNB N_B1_M1003_g 0.0230101f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=2.465
cc_9 VNB N_B1_M1015_g 0.0232626f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.465
cc_10 VNB N_B1_M1019_g 0.0242112f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.465
cc_11 VNB N_B1_M1036_g 0.00141113f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.465
cc_12 VNB N_B1_c_223_n 0.00165028f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_B1_c_224_n 0.0135487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_225_n 0.00250301f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.51
cc_15 VNB N_B1_c_226_n 0.046913f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.51
cc_16 VNB N_B1_c_227_n 0.0309826f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.51
cc_17 VNB N_B1_c_228_n 0.007778f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.51
cc_18 VNB N_B2_c_344_n 0.016406f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.345
cc_19 VNB N_B2_M1006_g 0.00688016f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.745
cc_20 VNB N_B2_c_346_n 0.0162007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B2_M1014_g 0.00674291f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.345
cc_22 VNB N_B2_c_348_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.745
cc_23 VNB N_B2_M1020_g 0.00674291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B2_c_350_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.745
cc_25 VNB N_B2_M1037_g 0.00675245f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.465
cc_26 VNB B2 0.00332766f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.465
cc_27 VNB N_B2_c_353_n 0.0782106f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.51
cc_28 VNB N_A1_M1016_g 0.00782695f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.745
cc_29 VNB N_A1_c_429_n 0.0155545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_M1017_g 0.00735878f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.345
cc_31 VNB N_A1_c_431_n 0.0159819f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.745
cc_32 VNB N_A1_M1029_g 0.00696422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A1_c_433_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.745
cc_34 VNB N_A1_M1033_g 0.0109923f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.465
cc_35 VNB N_A1_c_435_n 0.0029613f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.465
cc_36 VNB N_A1_c_436_n 0.0328708f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_37 VNB N_A1_c_437_n 0.0263405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_c_438_n 0.00632981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB A1 0.0261514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A1_c_440_n 0.0166215f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.51
cc_41 VNB N_A1_c_441_n 0.0911887f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.51
cc_42 VNB N_A2_M1009_g 0.0224154f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.745
cc_43 VNB N_A2_M1025_g 0.0227022f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=2.465
cc_44 VNB N_A2_M1038_g 0.0226825f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.465
cc_45 VNB N_A2_M1039_g 0.0228429f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.465
cc_46 VNB N_A2_c_543_n 0.0026038f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.51
cc_47 VNB N_A2_c_544_n 0.0647912f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.51
cc_48 VNB N_VPWR_c_621_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_Y_c_765_n 0.00301601f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=1.675
cc_50 VNB N_Y_c_766_n 0.00228543f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.465
cc_51 VNB N_Y_c_767_n 0.00895886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_Y_c_768_n 0.00402485f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.51
cc_53 VNB N_Y_c_769_n 0.00242434f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.51
cc_54 VNB N_A_29_65#_c_991_n 0.0311474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_29_65#_c_992_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.465
cc_56 VNB N_A_29_65#_c_993_n 0.00928796f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.465
cc_57 VNB N_A_29_65#_c_994_n 0.00651951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_29_65#_c_995_n 0.00373666f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_59 VNB N_A_29_65#_c_996_n 0.00879375f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_60 VNB N_A_29_65#_c_997_n 0.00353876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_29_65#_c_998_n 0.00228345f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.51
cc_62 VNB N_A_29_65#_c_999_n 0.00389499f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.51
cc_63 VNB N_A_509_47#_c_1084_n 0.00270842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_509_47#_c_1085_n 0.00740486f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.51
cc_65 VNB N_A_509_47#_c_1086_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.51
cc_66 VNB N_VGND_c_1190_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.745
cc_67 VNB N_VGND_c_1191_n 0.011684f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.675
cc_68 VNB N_VGND_c_1192_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.345
cc_69 VNB N_VGND_c_1193_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.675
cc_70 VNB N_VGND_c_1194_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=1.675
cc_71 VNB N_VGND_c_1195_n 0.149489f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.465
cc_72 VNB N_VGND_c_1196_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1197_n 0.011684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1198_n 0.0123026f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.51
cc_75 VNB N_VGND_c_1199_n 0.0180807f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.51
cc_76 VNB N_VGND_c_1200_n 0.48609f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.51
cc_77 VNB N_VGND_c_1201_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.51
cc_78 VNB N_VGND_c_1202_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.51
cc_79 VNB N_VGND_c_1203_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.51
cc_80 VPB N_C1_M1001_g 0.0235869f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=2.465
cc_81 VPB N_C1_M1004_g 0.0179387f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=2.465
cc_82 VPB N_C1_M1010_g 0.0179304f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=2.465
cc_83 VPB N_C1_M1024_g 0.0178625f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=2.465
cc_84 VPB C1 0.0413848f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_85 VPB N_C1_c_139_n 0.0382296f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=1.51
cc_86 VPB N_B1_M1011_g 0.0177365f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.745
cc_87 VPB N_B1_M1023_g 0.0176451f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.745
cc_88 VPB N_B1_M1026_g 0.0177937f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=0.745
cc_89 VPB N_B1_M1036_g 0.0209135f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=2.465
cc_90 VPB N_B1_c_223_n 0.00564855f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_91 VPB N_B1_c_224_n 0.0130361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_B1_c_225_n 3.91316e-19 $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.51
cc_93 VPB N_B1_c_226_n 0.00839363f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.51
cc_94 VPB N_B1_c_228_n 0.0033785f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=1.51
cc_95 VPB N_B2_M1006_g 0.0188867f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.745
cc_96 VPB N_B2_M1014_g 0.0187375f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.345
cc_97 VPB N_B2_M1020_g 0.0187375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_B2_M1037_g 0.0188867f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=2.465
cc_99 VPB N_A1_M1016_g 0.0223632f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.745
cc_100 VPB N_A1_M1017_g 0.0189105f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.345
cc_101 VPB N_A1_M1029_g 0.0183705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A1_M1033_g 0.027229f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=2.465
cc_103 VPB N_A2_M1000_g 0.0183424f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.745
cc_104 VPB N_A2_M1008_g 0.0181378f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.745
cc_105 VPB N_A2_M1028_g 0.0181347f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=0.745
cc_106 VPB N_A2_M1034_g 0.019089f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=2.465
cc_107 VPB N_A2_c_543_n 0.00977364f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.51
cc_108 VPB N_A2_c_544_n 0.0123278f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.51
cc_109 VPB N_VPWR_c_622_n 0.048246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_623_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_624_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_625_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_113 VPB N_VPWR_c_626_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_627_n 0.00563065f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.51
cc_115 VPB N_VPWR_c_628_n 4.05231e-19 $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.51
cc_116 VPB N_VPWR_c_629_n 0.0124746f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.51
cc_117 VPB N_VPWR_c_630_n 0.0560622f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=1.51
cc_118 VPB N_VPWR_c_631_n 0.0271236f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.51
cc_119 VPB N_VPWR_c_632_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.51
cc_120 VPB N_VPWR_c_633_n 0.0545613f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.51
cc_121 VPB N_VPWR_c_634_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=1.51
cc_122 VPB N_VPWR_c_635_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_636_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.587
cc_124 VPB N_VPWR_c_637_n 0.054581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_638_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_639_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_640_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_641_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_642_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_621_n 0.0752287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_Y_c_768_n 0.00126737f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.51
cc_132 VPB N_A_1317_367#_c_945_n 0.00663276f $X=-0.19 $Y=1.655 $X2=2.455
+ $Y2=1.675
cc_133 VPB N_A_1317_367#_c_946_n 0.00330214f $X=-0.19 $Y=1.655 $X2=2.455
+ $Y2=2.465
cc_134 N_C1_M1024_g N_B1_M1011_g 0.0256771f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_135 N_C1_c_139_n N_B1_c_223_n 3.96787e-19 $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_136 N_C1_c_139_n N_B1_c_226_n 0.0256771f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_137 N_C1_M1001_g N_VPWR_c_622_n 0.0203776f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_138 N_C1_M1004_g N_VPWR_c_622_n 7.28867e-19 $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_139 C1 N_VPWR_c_622_n 0.0257064f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_140 N_C1_c_139_n N_VPWR_c_622_n 0.00181296f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_141 N_C1_M1001_g N_VPWR_c_623_n 0.00486043f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_142 N_C1_M1004_g N_VPWR_c_623_n 0.00486043f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_143 N_C1_M1001_g N_VPWR_c_624_n 6.93132e-19 $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_144 N_C1_M1004_g N_VPWR_c_624_n 0.0149058f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_145 N_C1_M1010_g N_VPWR_c_624_n 0.0147185f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_146 N_C1_M1024_g N_VPWR_c_624_n 6.80491e-19 $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_147 N_C1_M1010_g N_VPWR_c_625_n 6.7059e-19 $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_148 N_C1_M1024_g N_VPWR_c_625_n 0.0138087f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_149 N_C1_M1010_g N_VPWR_c_635_n 0.00486043f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_150 N_C1_M1024_g N_VPWR_c_635_n 0.00486043f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_151 N_C1_M1001_g N_VPWR_c_621_n 0.00824727f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_152 N_C1_M1004_g N_VPWR_c_621_n 0.00824727f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_153 N_C1_M1010_g N_VPWR_c_621_n 0.00824727f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_154 N_C1_M1024_g N_VPWR_c_621_n 0.00824727f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_155 N_C1_M1005_g N_Y_c_771_n 0.00553704f $X=0.485 $Y=0.745 $X2=0 $Y2=0
cc_156 N_C1_M1018_g N_Y_c_771_n 0.00718404f $X=0.915 $Y=0.745 $X2=0 $Y2=0
cc_157 N_C1_M1021_g N_Y_c_771_n 3.83324e-19 $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_158 N_C1_M1018_g N_Y_c_765_n 0.00966312f $X=0.915 $Y=0.745 $X2=0 $Y2=0
cc_159 N_C1_M1021_g N_Y_c_765_n 0.0133983f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_160 C1 N_Y_c_765_n 0.0491972f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_161 N_C1_c_139_n N_Y_c_765_n 0.00516717f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_162 N_C1_M1005_g N_Y_c_766_n 0.00578377f $X=0.485 $Y=0.745 $X2=0 $Y2=0
cc_163 N_C1_M1018_g N_Y_c_766_n 0.00180314f $X=0.915 $Y=0.745 $X2=0 $Y2=0
cc_164 C1 N_Y_c_766_n 0.0275105f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_165 N_C1_c_139_n N_Y_c_766_n 0.00256054f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_166 C1 N_Y_c_782_n 0.0149585f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_167 N_C1_c_139_n N_Y_c_782_n 6.4545e-19 $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_168 N_C1_M1032_g N_Y_c_784_n 0.0100087f $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_169 N_C1_M1032_g N_Y_c_767_n 0.0123156f $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_170 C1 N_Y_c_767_n 0.0313254f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_171 N_C1_c_139_n N_Y_c_767_n 0.0135439f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_172 N_C1_M1032_g N_Y_c_768_n 0.00228383f $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_173 N_C1_M1010_g N_Y_c_768_n 7.78799e-19 $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_174 N_C1_M1024_g N_Y_c_768_n 0.00626971f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_175 C1 N_Y_c_768_n 0.0250004f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_176 N_C1_c_139_n N_Y_c_768_n 0.0125975f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_177 N_C1_M1032_g N_Y_c_769_n 0.00137054f $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_178 C1 N_Y_c_769_n 0.0277112f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_179 N_C1_c_139_n N_Y_c_769_n 0.00534045f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_180 N_C1_M1004_g N_Y_c_796_n 0.0122595f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_181 N_C1_M1010_g N_Y_c_796_n 0.0122129f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_182 C1 N_Y_c_796_n 0.0541337f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_183 N_C1_c_139_n N_Y_c_796_n 5.71535e-19 $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_184 N_C1_M1024_g N_Y_c_800_n 0.0133222f $X=2.455 $Y=2.465 $X2=0 $Y2=0
cc_185 N_C1_c_139_n N_Y_c_800_n 5.86662e-19 $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_186 N_C1_M1005_g N_A_29_65#_c_991_n 0.00354524f $X=0.485 $Y=0.745 $X2=0 $Y2=0
cc_187 C1 N_A_29_65#_c_991_n 0.0174135f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_188 N_C1_c_139_n N_A_29_65#_c_991_n 0.00281956f $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_189 N_C1_M1005_g N_A_29_65#_c_992_n 0.0125492f $X=0.485 $Y=0.745 $X2=0 $Y2=0
cc_190 N_C1_M1018_g N_A_29_65#_c_992_n 0.0116888f $X=0.915 $Y=0.745 $X2=0 $Y2=0
cc_191 N_C1_M1021_g N_A_29_65#_c_1005_n 0.00633387f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_192 N_C1_M1032_g N_A_29_65#_c_1005_n 3.1427e-19 $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_193 N_C1_M1021_g N_A_29_65#_c_994_n 0.00925833f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_194 N_C1_M1032_g N_A_29_65#_c_994_n 0.0133221f $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_195 N_C1_c_139_n N_A_29_65#_c_996_n 5.10906e-19 $X=2.455 $Y=1.51 $X2=0 $Y2=0
cc_196 N_C1_M1021_g N_A_29_65#_c_998_n 0.00132489f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_197 N_C1_M1032_g N_A_509_47#_c_1084_n 8.28001e-19 $X=1.935 $Y=0.745 $X2=0
+ $Y2=0
cc_198 N_C1_M1005_g N_VGND_c_1195_n 0.00302501f $X=0.485 $Y=0.745 $X2=0 $Y2=0
cc_199 N_C1_M1018_g N_VGND_c_1195_n 0.00302501f $X=0.915 $Y=0.745 $X2=0 $Y2=0
cc_200 N_C1_M1021_g N_VGND_c_1195_n 0.00302484f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_201 N_C1_M1032_g N_VGND_c_1195_n 0.00302501f $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_202 N_C1_M1005_g N_VGND_c_1200_n 0.004709f $X=0.485 $Y=0.745 $X2=0 $Y2=0
cc_203 N_C1_M1018_g N_VGND_c_1200_n 0.00442123f $X=0.915 $Y=0.745 $X2=0 $Y2=0
cc_204 N_C1_M1021_g N_VGND_c_1200_n 0.00449574f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_205 N_C1_M1032_g N_VGND_c_1200_n 0.00488475f $X=1.935 $Y=0.745 $X2=0 $Y2=0
cc_206 N_B1_M1015_g N_B2_c_344_n 0.0300315f $X=3.745 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_207 N_B1_M1026_g N_B2_M1006_g 0.0300315f $X=3.745 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B1_c_224_n N_B2_M1006_g 0.0121154f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_209 N_B1_c_224_n N_B2_M1014_g 0.0104915f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_210 N_B1_c_224_n N_B2_M1020_g 0.0104475f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_211 N_B1_M1019_g N_B2_c_350_n 0.0322997f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_212 N_B1_M1036_g N_B2_M1037_g 0.0388603f $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B1_c_224_n N_B2_M1037_g 0.0101665f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_214 N_B1_c_227_n N_B2_M1037_g 0.00601155f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_215 N_B1_c_228_n N_B2_M1037_g 7.19093e-19 $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_216 N_B1_M1015_g B2 9.03374e-19 $X=3.745 $Y=0.655 $X2=0 $Y2=0
cc_217 N_B1_M1019_g B2 0.00267012f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_218 N_B1_c_224_n B2 0.10301f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_219 N_B1_c_225_n B2 0.00179798f $X=3.82 $Y=1.592 $X2=0 $Y2=0
cc_220 N_B1_c_227_n B2 9.70329e-19 $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_221 N_B1_c_228_n B2 0.0125651f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_222 N_B1_M1019_g N_B2_c_353_n 0.00552417f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_223 N_B1_c_224_n N_B2_c_353_n 0.00815866f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_224 N_B1_c_225_n N_B2_c_353_n 0.00134682f $X=3.82 $Y=1.592 $X2=0 $Y2=0
cc_225 N_B1_c_226_n N_B2_c_353_n 0.0300315f $X=3.745 $Y=1.51 $X2=0 $Y2=0
cc_226 N_B1_c_227_n N_B2_c_353_n 0.014411f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_227 N_B1_c_228_n N_B2_c_353_n 6.59738e-19 $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_228 N_B1_M1036_g N_A1_M1016_g 0.0345097f $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_229 N_B1_c_227_n N_A1_M1016_g 0.00382983f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_230 N_B1_c_228_n N_A1_M1016_g 0.00578738f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_231 N_B1_M1019_g N_A1_c_435_n 0.00249135f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_232 N_B1_c_227_n N_A1_c_435_n 2.34651e-19 $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_233 N_B1_c_228_n N_A1_c_435_n 0.0124411f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_234 N_B1_M1019_g N_A1_c_436_n 0.00374816f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_235 N_B1_c_227_n N_A1_c_436_n 0.013774f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_236 N_B1_c_228_n N_A1_c_436_n 0.00147566f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_237 N_B1_M1019_g N_A1_c_440_n 0.0224178f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_238 N_B1_M1011_g N_VPWR_c_625_n 0.013789f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1023_g N_VPWR_c_625_n 6.22777e-19 $X=3.315 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_M1011_g N_VPWR_c_626_n 5.74401e-19 $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B1_M1023_g N_VPWR_c_626_n 0.01058f $X=3.315 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B1_M1026_g N_VPWR_c_626_n 0.0117529f $X=3.745 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1036_g N_VPWR_c_627_n 0.0109857f $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B1_M1026_g N_VPWR_c_633_n 0.00486043f $X=3.745 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_M1036_g N_VPWR_c_633_n 0.00547432f $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B1_M1011_g N_VPWR_c_636_n 0.00486043f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B1_M1023_g N_VPWR_c_636_n 0.00486043f $X=3.315 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B1_M1011_g N_VPWR_c_621_n 0.00824727f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_249 N_B1_M1023_g N_VPWR_c_621_n 0.00824727f $X=3.315 $Y=2.465 $X2=0 $Y2=0
cc_250 N_B1_M1026_g N_VPWR_c_621_n 0.0082726f $X=3.745 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B1_M1036_g N_VPWR_c_621_n 0.0103952f $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_252 N_B1_M1002_g N_Y_c_767_n 0.00392226f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_253 N_B1_M1002_g N_Y_c_768_n 0.00431895f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_254 N_B1_M1011_g N_Y_c_768_n 0.0028437f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B1_c_223_n N_Y_c_768_n 0.030692f $X=3.628 $Y=1.592 $X2=0 $Y2=0
cc_256 N_B1_c_226_n N_Y_c_768_n 0.00121127f $X=3.745 $Y=1.51 $X2=0 $Y2=0
cc_257 N_B1_M1011_g N_Y_c_807_n 0.0142932f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_258 N_B1_M1023_g N_Y_c_807_n 0.0104926f $X=3.315 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B1_M1026_g N_Y_c_807_n 0.010446f $X=3.745 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B1_c_223_n N_Y_c_807_n 0.0933902f $X=3.628 $Y=1.592 $X2=0 $Y2=0
cc_261 N_B1_c_226_n N_Y_c_807_n 0.0010661f $X=3.745 $Y=1.51 $X2=0 $Y2=0
cc_262 N_B1_c_224_n N_Y_c_812_n 0.0335742f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_263 N_B1_M1011_g N_Y_c_800_n 9.36327e-19 $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_264 N_B1_M1026_g N_Y_c_814_n 7.12951e-19 $X=3.745 $Y=2.465 $X2=0 $Y2=0
cc_265 N_B1_c_224_n N_Y_c_814_n 0.0217611f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_266 N_B1_M1036_g N_Y_c_816_n 9.05787e-19 $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_267 N_B1_c_224_n N_Y_c_816_n 0.0217611f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_268 N_B1_M1036_g Y 0.0155792f $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_269 N_B1_c_224_n Y 0.0249102f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_270 N_B1_c_227_n Y 6.02872e-19 $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_271 N_B1_c_228_n Y 0.0233735f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_272 N_B1_M1023_g N_A_592_367#_c_906_n 0.0122129f $X=3.315 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_B1_M1026_g N_A_592_367#_c_906_n 0.0122129f $X=3.745 $Y=2.465 $X2=0
+ $Y2=0
cc_274 N_B1_M1036_g N_A_592_367#_c_908_n 0.00211957f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_275 N_B1_M1036_g N_A_592_367#_c_909_n 0.00751822f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_B1_M1002_g N_A_29_65#_c_995_n 0.00331258f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_277 N_B1_M1002_g N_A_29_65#_c_996_n 0.0286363f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_278 N_B1_M1003_g N_A_29_65#_c_996_n 4.69757e-19 $X=3.315 $Y=0.655 $X2=0 $Y2=0
cc_279 N_B1_c_223_n N_A_29_65#_c_996_n 0.0315446f $X=3.628 $Y=1.592 $X2=0 $Y2=0
cc_280 N_B1_c_226_n N_A_29_65#_c_996_n 0.00247298f $X=3.745 $Y=1.51 $X2=0 $Y2=0
cc_281 N_B1_M1003_g N_A_29_65#_c_997_n 0.0122864f $X=3.315 $Y=0.655 $X2=0 $Y2=0
cc_282 N_B1_M1015_g N_A_29_65#_c_997_n 0.0135672f $X=3.745 $Y=0.655 $X2=0 $Y2=0
cc_283 N_B1_c_223_n N_A_29_65#_c_997_n 0.0473541f $X=3.628 $Y=1.592 $X2=0 $Y2=0
cc_284 N_B1_c_224_n N_A_29_65#_c_997_n 0.00192453f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_285 N_B1_c_226_n N_A_29_65#_c_997_n 0.00240865f $X=3.745 $Y=1.51 $X2=0 $Y2=0
cc_286 N_B1_c_224_n N_A_29_65#_c_999_n 0.00981509f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_287 N_B1_M1019_g N_A_29_65#_c_1022_n 0.00581329f $X=5.895 $Y=0.655 $X2=0
+ $Y2=0
cc_288 N_B1_c_228_n N_A_29_65#_c_1022_n 0.00143411f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_289 N_B1_c_224_n N_A_29_65#_c_1024_n 0.00731876f $X=5.815 $Y=1.7 $X2=0 $Y2=0
cc_290 N_B1_M1002_g N_A_509_47#_c_1084_n 0.0092657f $X=2.885 $Y=0.655 $X2=0
+ $Y2=0
cc_291 N_B1_M1003_g N_A_509_47#_c_1084_n 0.00963386f $X=3.315 $Y=0.655 $X2=0
+ $Y2=0
cc_292 N_B1_M1019_g N_A_509_47#_c_1090_n 0.0150738f $X=5.895 $Y=0.655 $X2=0
+ $Y2=0
cc_293 N_B1_M1019_g N_A_509_47#_c_1091_n 0.00900978f $X=5.895 $Y=0.655 $X2=0
+ $Y2=0
cc_294 N_B1_c_227_n N_A_509_47#_c_1091_n 3.94631e-19 $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_295 N_B1_c_228_n N_A_509_47#_c_1091_n 0.00423796f $X=5.95 $Y=1.46 $X2=0 $Y2=0
cc_296 N_B1_M1002_g N_A_509_47#_c_1094_n 7.61432e-19 $X=2.885 $Y=0.655 $X2=0
+ $Y2=0
cc_297 N_B1_M1003_g N_A_509_47#_c_1094_n 0.00594636f $X=3.315 $Y=0.655 $X2=0
+ $Y2=0
cc_298 N_B1_M1015_g N_A_509_47#_c_1094_n 0.00628307f $X=3.745 $Y=0.655 $X2=0
+ $Y2=0
cc_299 N_B1_M1015_g N_A_509_47#_c_1097_n 0.00873689f $X=3.745 $Y=0.655 $X2=0
+ $Y2=0
cc_300 N_B1_M1019_g N_VGND_c_1190_n 0.00102789f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_301 N_B1_M1002_g N_VGND_c_1195_n 0.00357877f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_302 N_B1_M1003_g N_VGND_c_1195_n 0.00357842f $X=3.315 $Y=0.655 $X2=0 $Y2=0
cc_303 N_B1_M1015_g N_VGND_c_1195_n 0.00357842f $X=3.745 $Y=0.655 $X2=0 $Y2=0
cc_304 N_B1_M1019_g N_VGND_c_1195_n 0.00357877f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_305 N_B1_M1002_g N_VGND_c_1200_n 0.00665089f $X=2.885 $Y=0.655 $X2=0 $Y2=0
cc_306 N_B1_M1003_g N_VGND_c_1200_n 0.00535118f $X=3.315 $Y=0.655 $X2=0 $Y2=0
cc_307 N_B1_M1015_g N_VGND_c_1200_n 0.00537847f $X=3.745 $Y=0.655 $X2=0 $Y2=0
cc_308 N_B1_M1019_g N_VGND_c_1200_n 0.00588745f $X=5.895 $Y=0.655 $X2=0 $Y2=0
cc_309 N_B2_M1006_g N_VPWR_c_626_n 0.00109252f $X=4.175 $Y=2.465 $X2=0 $Y2=0
cc_310 N_B2_M1006_g N_VPWR_c_633_n 0.00357877f $X=4.175 $Y=2.465 $X2=0 $Y2=0
cc_311 N_B2_M1014_g N_VPWR_c_633_n 0.00357877f $X=4.605 $Y=2.465 $X2=0 $Y2=0
cc_312 N_B2_M1020_g N_VPWR_c_633_n 0.00357877f $X=5.035 $Y=2.465 $X2=0 $Y2=0
cc_313 N_B2_M1037_g N_VPWR_c_633_n 0.00357877f $X=5.465 $Y=2.465 $X2=0 $Y2=0
cc_314 N_B2_M1006_g N_VPWR_c_621_n 0.00537654f $X=4.175 $Y=2.465 $X2=0 $Y2=0
cc_315 N_B2_M1014_g N_VPWR_c_621_n 0.0053512f $X=4.605 $Y=2.465 $X2=0 $Y2=0
cc_316 N_B2_M1020_g N_VPWR_c_621_n 0.0053512f $X=5.035 $Y=2.465 $X2=0 $Y2=0
cc_317 N_B2_M1037_g N_VPWR_c_621_n 0.00537654f $X=5.465 $Y=2.465 $X2=0 $Y2=0
cc_318 N_B2_M1006_g N_Y_c_807_n 0.0111034f $X=4.175 $Y=2.465 $X2=0 $Y2=0
cc_319 N_B2_M1014_g N_Y_c_812_n 0.0114269f $X=4.605 $Y=2.465 $X2=0 $Y2=0
cc_320 N_B2_M1020_g N_Y_c_812_n 0.0114269f $X=5.035 $Y=2.465 $X2=0 $Y2=0
cc_321 N_B2_M1006_g N_Y_c_814_n 0.0107562f $X=4.175 $Y=2.465 $X2=0 $Y2=0
cc_322 N_B2_M1014_g N_Y_c_814_n 0.0106171f $X=4.605 $Y=2.465 $X2=0 $Y2=0
cc_323 N_B2_M1020_g N_Y_c_814_n 5.8311e-19 $X=5.035 $Y=2.465 $X2=0 $Y2=0
cc_324 N_B2_M1014_g N_Y_c_816_n 5.8311e-19 $X=4.605 $Y=2.465 $X2=0 $Y2=0
cc_325 N_B2_M1020_g N_Y_c_816_n 0.0106171f $X=5.035 $Y=2.465 $X2=0 $Y2=0
cc_326 N_B2_M1037_g N_Y_c_816_n 0.0106824f $X=5.465 $Y=2.465 $X2=0 $Y2=0
cc_327 N_B2_M1037_g Y 0.0113776f $X=5.465 $Y=2.465 $X2=0 $Y2=0
cc_328 N_B2_M1006_g N_A_592_367#_c_910_n 0.0115031f $X=4.175 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_B2_M1014_g N_A_592_367#_c_910_n 0.0114565f $X=4.605 $Y=2.465 $X2=0
+ $Y2=0
cc_330 N_B2_M1020_g N_A_592_367#_c_908_n 0.0115031f $X=5.035 $Y=2.465 $X2=0
+ $Y2=0
cc_331 N_B2_M1037_g N_A_592_367#_c_908_n 0.0115031f $X=5.465 $Y=2.465 $X2=0
+ $Y2=0
cc_332 N_B2_c_344_n N_A_29_65#_c_999_n 0.00856963f $X=4.175 $Y=1.185 $X2=0 $Y2=0
cc_333 N_B2_c_346_n N_A_29_65#_c_999_n 7.27631e-19 $X=4.605 $Y=1.185 $X2=0 $Y2=0
cc_334 B2 N_A_29_65#_c_999_n 0.00290184f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_335 N_B2_c_348_n N_A_29_65#_c_1022_n 5.32462e-19 $X=5.035 $Y=1.185 $X2=0
+ $Y2=0
cc_336 N_B2_c_350_n N_A_29_65#_c_1022_n 0.00328699f $X=5.465 $Y=1.185 $X2=0
+ $Y2=0
cc_337 N_B2_c_344_n N_A_29_65#_c_1024_n 0.0111868f $X=4.175 $Y=1.185 $X2=0 $Y2=0
cc_338 N_B2_c_346_n N_A_29_65#_c_1024_n 0.0105171f $X=4.605 $Y=1.185 $X2=0 $Y2=0
cc_339 N_B2_c_348_n N_A_29_65#_c_1024_n 0.0105805f $X=5.035 $Y=1.185 $X2=0 $Y2=0
cc_340 N_B2_c_350_n N_A_29_65#_c_1024_n 0.00909778f $X=5.465 $Y=1.185 $X2=0
+ $Y2=0
cc_341 B2 N_A_29_65#_c_1024_n 0.0897293f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_342 N_B2_c_353_n N_A_29_65#_c_1024_n 0.00686781f $X=5.465 $Y=1.35 $X2=0 $Y2=0
cc_343 N_B2_c_346_n N_A_509_47#_c_1098_n 0.00655472f $X=4.605 $Y=1.185 $X2=0
+ $Y2=0
cc_344 N_B2_c_348_n N_A_509_47#_c_1098_n 0.0123829f $X=5.035 $Y=1.185 $X2=0
+ $Y2=0
cc_345 N_B2_c_346_n N_A_509_47#_c_1100_n 0.00577264f $X=4.605 $Y=1.185 $X2=0
+ $Y2=0
cc_346 N_B2_c_350_n N_A_509_47#_c_1090_n 0.0102091f $X=5.465 $Y=1.185 $X2=0
+ $Y2=0
cc_347 N_B2_c_344_n N_A_509_47#_c_1094_n 3.46799e-19 $X=4.175 $Y=1.185 $X2=0
+ $Y2=0
cc_348 N_B2_c_344_n N_A_509_47#_c_1097_n 0.0102183f $X=4.175 $Y=1.185 $X2=0
+ $Y2=0
cc_349 N_B2_c_344_n N_VGND_c_1195_n 0.00357877f $X=4.175 $Y=1.185 $X2=0 $Y2=0
cc_350 N_B2_c_346_n N_VGND_c_1195_n 0.00357877f $X=4.605 $Y=1.185 $X2=0 $Y2=0
cc_351 N_B2_c_348_n N_VGND_c_1195_n 0.00357877f $X=5.035 $Y=1.185 $X2=0 $Y2=0
cc_352 N_B2_c_350_n N_VGND_c_1195_n 0.00357877f $X=5.465 $Y=1.185 $X2=0 $Y2=0
cc_353 N_B2_c_344_n N_VGND_c_1200_n 0.00544013f $X=4.175 $Y=1.185 $X2=0 $Y2=0
cc_354 N_B2_c_346_n N_VGND_c_1200_n 0.00541285f $X=4.605 $Y=1.185 $X2=0 $Y2=0
cc_355 N_B2_c_348_n N_VGND_c_1200_n 0.00541285f $X=5.035 $Y=1.185 $X2=0 $Y2=0
cc_356 N_B2_c_350_n N_VGND_c_1200_n 0.00544013f $X=5.465 $Y=1.185 $X2=0 $Y2=0
cc_357 N_A1_c_435_n N_A2_M1009_g 0.00142999f $X=6.53 $Y=1.16 $X2=0 $Y2=0
cc_358 N_A1_c_436_n N_A2_M1009_g 0.0216425f $X=6.49 $Y=1.35 $X2=0 $Y2=0
cc_359 N_A1_c_437_n N_A2_M1009_g 0.0100319f $X=8.385 $Y=1.297 $X2=0 $Y2=0
cc_360 N_A1_c_440_n N_A2_M1009_g 0.0315617f $X=6.49 $Y=1.185 $X2=0 $Y2=0
cc_361 N_A1_c_437_n N_A2_M1025_g 0.0105073f $X=8.385 $Y=1.297 $X2=0 $Y2=0
cc_362 N_A1_c_437_n N_A2_M1038_g 0.0105539f $X=8.385 $Y=1.297 $X2=0 $Y2=0
cc_363 N_A1_c_429_n N_A2_M1039_g 0.0227472f $X=8.66 $Y=1.185 $X2=0 $Y2=0
cc_364 N_A1_c_437_n N_A2_M1039_g 0.0132193f $X=8.385 $Y=1.297 $X2=0 $Y2=0
cc_365 N_A1_c_438_n N_A2_M1039_g 0.00656433f $X=8.59 $Y=1.297 $X2=0 $Y2=0
cc_366 N_A1_M1016_g N_A2_c_543_n 0.00593249f $X=6.51 $Y=2.465 $X2=0 $Y2=0
cc_367 N_A1_M1017_g N_A2_c_543_n 9.13462e-19 $X=8.695 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A1_c_435_n N_A2_c_543_n 0.00736589f $X=6.53 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A1_c_436_n N_A2_c_543_n 5.45798e-19 $X=6.49 $Y=1.35 $X2=0 $Y2=0
cc_370 N_A1_c_437_n N_A2_c_543_n 0.098195f $X=8.385 $Y=1.297 $X2=0 $Y2=0
cc_371 N_A1_c_438_n N_A2_c_543_n 0.00829041f $X=8.59 $Y=1.297 $X2=0 $Y2=0
cc_372 N_A1_M1016_g N_A2_c_544_n 0.0431221f $X=6.51 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A1_M1017_g N_A2_c_544_n 0.0230361f $X=8.695 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A1_c_437_n N_A2_c_544_n 0.00734707f $X=8.385 $Y=1.297 $X2=0 $Y2=0
cc_375 N_A1_c_441_n N_A2_c_544_n 0.0227472f $X=9.77 $Y=1.35 $X2=0 $Y2=0
cc_376 N_A1_M1016_g N_VPWR_c_627_n 0.00826441f $X=6.51 $Y=2.465 $X2=0 $Y2=0
cc_377 N_A1_M1017_g N_VPWR_c_628_n 0.0168375f $X=8.695 $Y=2.465 $X2=0 $Y2=0
cc_378 N_A1_M1029_g N_VPWR_c_628_n 0.0156786f $X=9.125 $Y=2.465 $X2=0 $Y2=0
cc_379 N_A1_M1033_g N_VPWR_c_628_n 7.59779e-19 $X=9.555 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A1_M1033_g N_VPWR_c_630_n 0.00768161f $X=9.555 $Y=2.465 $X2=0 $Y2=0
cc_381 A1 N_VPWR_c_630_n 0.0175666f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_382 N_A1_c_441_n N_VPWR_c_630_n 0.00214862f $X=9.77 $Y=1.35 $X2=0 $Y2=0
cc_383 N_A1_M1016_g N_VPWR_c_637_n 0.00547432f $X=6.51 $Y=2.465 $X2=0 $Y2=0
cc_384 N_A1_M1017_g N_VPWR_c_637_n 0.00486043f $X=8.695 $Y=2.465 $X2=0 $Y2=0
cc_385 N_A1_M1029_g N_VPWR_c_638_n 0.00486043f $X=9.125 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A1_M1033_g N_VPWR_c_638_n 0.00585385f $X=9.555 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A1_M1016_g N_VPWR_c_621_n 0.0103269f $X=6.51 $Y=2.465 $X2=0 $Y2=0
cc_388 N_A1_M1017_g N_VPWR_c_621_n 0.00835496f $X=8.695 $Y=2.465 $X2=0 $Y2=0
cc_389 N_A1_M1029_g N_VPWR_c_621_n 0.00824727f $X=9.125 $Y=2.465 $X2=0 $Y2=0
cc_390 N_A1_M1033_g N_VPWR_c_621_n 0.011499f $X=9.555 $Y=2.465 $X2=0 $Y2=0
cc_391 N_A1_c_436_n Y 0.00176545f $X=6.49 $Y=1.35 $X2=0 $Y2=0
cc_392 N_A1_M1016_g N_Y_c_833_n 9.08502e-19 $X=6.51 $Y=2.465 $X2=0 $Y2=0
cc_393 N_A1_M1016_g N_Y_c_834_n 0.0172078f $X=6.51 $Y=2.465 $X2=0 $Y2=0
cc_394 N_A1_c_435_n N_Y_c_834_n 0.0071949f $X=6.53 $Y=1.16 $X2=0 $Y2=0
cc_395 N_A1_c_436_n N_Y_c_834_n 2.1514e-19 $X=6.49 $Y=1.35 $X2=0 $Y2=0
cc_396 N_A1_M1016_g N_A_1317_367#_c_947_n 0.00715449f $X=6.51 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_A1_M1016_g N_A_1317_367#_c_948_n 0.0020078f $X=6.51 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_A1_M1017_g N_A_1317_367#_c_945_n 0.0136791f $X=8.695 $Y=2.465 $X2=0
+ $Y2=0
cc_399 N_A1_M1029_g N_A_1317_367#_c_945_n 0.0136563f $X=9.125 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A1_M1033_g N_A_1317_367#_c_945_n 0.00435578f $X=9.555 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A1_c_438_n N_A_1317_367#_c_945_n 0.0504232f $X=8.59 $Y=1.297 $X2=0
+ $Y2=0
cc_402 A1 N_A_1317_367#_c_945_n 0.0198134f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_403 N_A1_c_441_n N_A_1317_367#_c_945_n 0.00173078f $X=9.77 $Y=1.35 $X2=0
+ $Y2=0
cc_404 N_A1_c_438_n N_A_1317_367#_c_946_n 0.0171749f $X=8.59 $Y=1.297 $X2=0
+ $Y2=0
cc_405 N_A1_c_440_n N_A_29_65#_c_1022_n 4.92483e-19 $X=6.49 $Y=1.185 $X2=0 $Y2=0
cc_406 N_A1_c_435_n N_A_509_47#_M1019_d 3.17466e-19 $X=6.53 $Y=1.16 $X2=0 $Y2=0
cc_407 N_A1_c_436_n N_A_509_47#_c_1091_n 0.00228344f $X=6.49 $Y=1.35 $X2=0 $Y2=0
cc_408 N_A1_c_440_n N_A_509_47#_c_1091_n 9.83892e-19 $X=6.49 $Y=1.185 $X2=0
+ $Y2=0
cc_409 N_A1_c_435_n N_A_509_47#_c_1107_n 0.0155824f $X=6.53 $Y=1.16 $X2=0 $Y2=0
cc_410 N_A1_c_436_n N_A_509_47#_c_1107_n 2.66669e-19 $X=6.49 $Y=1.35 $X2=0 $Y2=0
cc_411 N_A1_c_437_n N_A_509_47#_c_1107_n 0.0252905f $X=8.385 $Y=1.297 $X2=0
+ $Y2=0
cc_412 N_A1_c_440_n N_A_509_47#_c_1107_n 0.0124367f $X=6.49 $Y=1.185 $X2=0 $Y2=0
cc_413 N_A1_c_437_n N_A_509_47#_c_1111_n 0.0402256f $X=8.385 $Y=1.297 $X2=0
+ $Y2=0
cc_414 N_A1_c_429_n N_A_509_47#_c_1112_n 0.0105886f $X=8.66 $Y=1.185 $X2=0 $Y2=0
cc_415 N_A1_c_437_n N_A_509_47#_c_1112_n 0.0299082f $X=8.385 $Y=1.297 $X2=0
+ $Y2=0
cc_416 A1 N_A_509_47#_c_1112_n 0.00699294f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_417 N_A1_c_431_n N_A_509_47#_c_1085_n 0.0122595f $X=9.09 $Y=1.185 $X2=0 $Y2=0
cc_418 N_A1_c_433_n N_A_509_47#_c_1085_n 0.0121992f $X=9.52 $Y=1.185 $X2=0 $Y2=0
cc_419 A1 N_A_509_47#_c_1085_n 0.061937f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_420 N_A1_c_441_n N_A_509_47#_c_1085_n 0.00865419f $X=9.77 $Y=1.35 $X2=0 $Y2=0
cc_421 N_A1_c_437_n N_A_509_47#_c_1119_n 0.0145842f $X=8.385 $Y=1.297 $X2=0
+ $Y2=0
cc_422 N_A1_c_437_n N_A_509_47#_c_1120_n 0.0145842f $X=8.385 $Y=1.297 $X2=0
+ $Y2=0
cc_423 A1 N_A_509_47#_c_1121_n 0.0152172f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_424 N_A1_c_441_n N_A_509_47#_c_1121_n 0.00254265f $X=9.77 $Y=1.35 $X2=0 $Y2=0
cc_425 N_A1_c_435_n N_VGND_M1007_d 7.5535e-19 $X=6.53 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_426 N_A1_c_440_n N_VGND_c_1190_n 0.00882183f $X=6.49 $Y=1.185 $X2=0 $Y2=0
cc_427 N_A1_c_429_n N_VGND_c_1193_n 0.00748371f $X=8.66 $Y=1.185 $X2=0 $Y2=0
cc_428 N_A1_c_431_n N_VGND_c_1193_n 5.37623e-19 $X=9.09 $Y=1.185 $X2=0 $Y2=0
cc_429 N_A1_c_429_n N_VGND_c_1194_n 5.75816e-19 $X=8.66 $Y=1.185 $X2=0 $Y2=0
cc_430 N_A1_c_431_n N_VGND_c_1194_n 0.0103296f $X=9.09 $Y=1.185 $X2=0 $Y2=0
cc_431 N_A1_c_433_n N_VGND_c_1194_n 0.0120167f $X=9.52 $Y=1.185 $X2=0 $Y2=0
cc_432 N_A1_c_440_n N_VGND_c_1195_n 0.00365202f $X=6.49 $Y=1.185 $X2=0 $Y2=0
cc_433 N_A1_c_429_n N_VGND_c_1198_n 0.00365202f $X=8.66 $Y=1.185 $X2=0 $Y2=0
cc_434 N_A1_c_431_n N_VGND_c_1198_n 0.00486043f $X=9.09 $Y=1.185 $X2=0 $Y2=0
cc_435 N_A1_c_433_n N_VGND_c_1199_n 0.00486043f $X=9.52 $Y=1.185 $X2=0 $Y2=0
cc_436 N_A1_c_429_n N_VGND_c_1200_n 0.00432244f $X=8.66 $Y=1.185 $X2=0 $Y2=0
cc_437 N_A1_c_431_n N_VGND_c_1200_n 0.00824727f $X=9.09 $Y=1.185 $X2=0 $Y2=0
cc_438 N_A1_c_433_n N_VGND_c_1200_n 0.00925092f $X=9.52 $Y=1.185 $X2=0 $Y2=0
cc_439 N_A1_c_440_n N_VGND_c_1200_n 0.00483706f $X=6.49 $Y=1.185 $X2=0 $Y2=0
cc_440 N_A2_M1034_g N_VPWR_c_628_n 0.00104138f $X=8.23 $Y=2.465 $X2=0 $Y2=0
cc_441 N_A2_M1000_g N_VPWR_c_637_n 0.00357877f $X=6.94 $Y=2.465 $X2=0 $Y2=0
cc_442 N_A2_M1008_g N_VPWR_c_637_n 0.00357877f $X=7.37 $Y=2.465 $X2=0 $Y2=0
cc_443 N_A2_M1028_g N_VPWR_c_637_n 0.00357877f $X=7.8 $Y=2.465 $X2=0 $Y2=0
cc_444 N_A2_M1034_g N_VPWR_c_637_n 0.00357877f $X=8.23 $Y=2.465 $X2=0 $Y2=0
cc_445 N_A2_M1000_g N_VPWR_c_621_n 0.00537654f $X=6.94 $Y=2.465 $X2=0 $Y2=0
cc_446 N_A2_M1008_g N_VPWR_c_621_n 0.0053512f $X=7.37 $Y=2.465 $X2=0 $Y2=0
cc_447 N_A2_M1028_g N_VPWR_c_621_n 0.0053512f $X=7.8 $Y=2.465 $X2=0 $Y2=0
cc_448 N_A2_M1034_g N_VPWR_c_621_n 0.0054589f $X=8.23 $Y=2.465 $X2=0 $Y2=0
cc_449 N_A2_M1008_g N_Y_c_837_n 0.0113002f $X=7.37 $Y=2.465 $X2=0 $Y2=0
cc_450 N_A2_M1028_g N_Y_c_837_n 0.0113002f $X=7.8 $Y=2.465 $X2=0 $Y2=0
cc_451 N_A2_c_544_n N_Y_c_837_n 5.68128e-19 $X=8.23 $Y=1.51 $X2=0 $Y2=0
cc_452 N_A2_M1008_g N_Y_c_840_n 5.6266e-19 $X=7.37 $Y=2.465 $X2=0 $Y2=0
cc_453 N_A2_M1028_g N_Y_c_840_n 0.0108085f $X=7.8 $Y=2.465 $X2=0 $Y2=0
cc_454 N_A2_M1034_g N_Y_c_840_n 0.0116093f $X=8.23 $Y=2.465 $X2=0 $Y2=0
cc_455 N_A2_c_543_n N_Y_c_840_n 0.0204377f $X=8.05 $Y=1.51 $X2=0 $Y2=0
cc_456 N_A2_c_544_n N_Y_c_840_n 6.50093e-19 $X=8.23 $Y=1.51 $X2=0 $Y2=0
cc_457 N_A2_M1000_g N_Y_c_833_n 0.0101371f $X=6.94 $Y=2.465 $X2=0 $Y2=0
cc_458 N_A2_M1008_g N_Y_c_833_n 0.00988739f $X=7.37 $Y=2.465 $X2=0 $Y2=0
cc_459 N_A2_M1028_g N_Y_c_833_n 5.1737e-19 $X=7.8 $Y=2.465 $X2=0 $Y2=0
cc_460 N_A2_M1000_g N_Y_c_834_n 0.0126312f $X=6.94 $Y=2.465 $X2=0 $Y2=0
cc_461 N_A2_M1008_g N_Y_c_834_n 0.00105834f $X=7.37 $Y=2.465 $X2=0 $Y2=0
cc_462 N_A2_c_543_n N_Y_c_834_n 0.0595573f $X=8.05 $Y=1.51 $X2=0 $Y2=0
cc_463 N_A2_c_544_n N_Y_c_834_n 5.72225e-19 $X=8.23 $Y=1.51 $X2=0 $Y2=0
cc_464 N_A2_M1000_g N_A_1317_367#_c_956_n 0.0115031f $X=6.94 $Y=2.465 $X2=0
+ $Y2=0
cc_465 N_A2_M1008_g N_A_1317_367#_c_956_n 0.0115031f $X=7.37 $Y=2.465 $X2=0
+ $Y2=0
cc_466 N_A2_M1028_g N_A_1317_367#_c_958_n 0.0114565f $X=7.8 $Y=2.465 $X2=0 $Y2=0
cc_467 N_A2_M1034_g N_A_1317_367#_c_958_n 0.0115031f $X=8.23 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_A2_M1034_g N_A_1317_367#_c_960_n 0.0082428f $X=8.23 $Y=2.465 $X2=0
+ $Y2=0
cc_469 N_A2_M1034_g N_A_1317_367#_c_946_n 0.00382078f $X=8.23 $Y=2.465 $X2=0
+ $Y2=0
cc_470 N_A2_c_543_n N_A_1317_367#_c_946_n 0.00525951f $X=8.05 $Y=1.51 $X2=0
+ $Y2=0
cc_471 N_A2_M1009_g N_A_509_47#_c_1107_n 0.0098539f $X=6.94 $Y=0.655 $X2=0 $Y2=0
cc_472 N_A2_M1025_g N_A_509_47#_c_1111_n 0.00990046f $X=7.37 $Y=0.655 $X2=0
+ $Y2=0
cc_473 N_A2_M1038_g N_A_509_47#_c_1111_n 0.00990046f $X=7.8 $Y=0.655 $X2=0 $Y2=0
cc_474 N_A2_M1039_g N_A_509_47#_c_1112_n 0.0098539f $X=8.23 $Y=0.655 $X2=0 $Y2=0
cc_475 N_A2_M1009_g N_VGND_c_1190_n 0.00754158f $X=6.94 $Y=0.655 $X2=0 $Y2=0
cc_476 N_A2_M1025_g N_VGND_c_1190_n 5.37623e-19 $X=7.37 $Y=0.655 $X2=0 $Y2=0
cc_477 N_A2_M1009_g N_VGND_c_1191_n 0.00365202f $X=6.94 $Y=0.655 $X2=0 $Y2=0
cc_478 N_A2_M1025_g N_VGND_c_1191_n 0.00365202f $X=7.37 $Y=0.655 $X2=0 $Y2=0
cc_479 N_A2_M1009_g N_VGND_c_1192_n 5.37623e-19 $X=6.94 $Y=0.655 $X2=0 $Y2=0
cc_480 N_A2_M1025_g N_VGND_c_1192_n 0.00758038f $X=7.37 $Y=0.655 $X2=0 $Y2=0
cc_481 N_A2_M1038_g N_VGND_c_1192_n 0.00758038f $X=7.8 $Y=0.655 $X2=0 $Y2=0
cc_482 N_A2_M1039_g N_VGND_c_1192_n 5.37623e-19 $X=8.23 $Y=0.655 $X2=0 $Y2=0
cc_483 N_A2_M1038_g N_VGND_c_1193_n 5.37623e-19 $X=7.8 $Y=0.655 $X2=0 $Y2=0
cc_484 N_A2_M1039_g N_VGND_c_1193_n 0.00754158f $X=8.23 $Y=0.655 $X2=0 $Y2=0
cc_485 N_A2_M1038_g N_VGND_c_1197_n 0.00365202f $X=7.8 $Y=0.655 $X2=0 $Y2=0
cc_486 N_A2_M1039_g N_VGND_c_1197_n 0.00365202f $X=8.23 $Y=0.655 $X2=0 $Y2=0
cc_487 N_A2_M1009_g N_VGND_c_1200_n 0.00432244f $X=6.94 $Y=0.655 $X2=0 $Y2=0
cc_488 N_A2_M1025_g N_VGND_c_1200_n 0.00432244f $X=7.37 $Y=0.655 $X2=0 $Y2=0
cc_489 N_A2_M1038_g N_VGND_c_1200_n 0.00432244f $X=7.8 $Y=0.655 $X2=0 $Y2=0
cc_490 N_A2_M1039_g N_VGND_c_1200_n 0.00432244f $X=8.23 $Y=0.655 $X2=0 $Y2=0
cc_491 N_VPWR_c_621_n N_Y_M1001_s 0.00571434f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_492 N_VPWR_c_621_n N_Y_M1010_s 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_493 N_VPWR_c_621_n N_Y_M1006_s 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_494 N_VPWR_c_621_n N_Y_M1020_s 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_495 N_VPWR_c_621_n N_Y_M1000_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_496 N_VPWR_c_621_n N_Y_M1028_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_497 N_VPWR_c_623_n N_Y_c_858_n 0.0120977f $X=1.645 $Y=3.33 $X2=0 $Y2=0
cc_498 N_VPWR_c_621_n N_Y_c_858_n 0.00691495f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_499 N_VPWR_c_635_n N_Y_c_860_n 0.0124525f $X=2.505 $Y=3.33 $X2=0 $Y2=0
cc_500 N_VPWR_c_621_n N_Y_c_860_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_501 N_VPWR_M1024_d N_Y_c_768_n 0.00114647f $X=2.53 $Y=1.835 $X2=0 $Y2=0
cc_502 N_VPWR_M1024_d N_Y_c_807_n 0.005464f $X=2.53 $Y=1.835 $X2=0 $Y2=0
cc_503 N_VPWR_M1023_d N_Y_c_807_n 0.00334477f $X=3.39 $Y=1.835 $X2=0 $Y2=0
cc_504 N_VPWR_M1004_d N_Y_c_796_n 0.00332836f $X=1.67 $Y=1.835 $X2=0 $Y2=0
cc_505 N_VPWR_c_624_n N_Y_c_796_n 0.0170777f $X=1.81 $Y=2.38 $X2=0 $Y2=0
cc_506 N_VPWR_M1024_d N_Y_c_800_n 0.00117565f $X=2.53 $Y=1.835 $X2=0 $Y2=0
cc_507 N_VPWR_c_625_n N_Y_c_800_n 0.0170826f $X=2.67 $Y=2.42 $X2=0 $Y2=0
cc_508 N_VPWR_M1036_d Y 0.0142641f $X=5.97 $Y=1.835 $X2=0 $Y2=0
cc_509 N_VPWR_c_627_n Y 0.026707f $X=6.215 $Y=2.435 $X2=0 $Y2=0
cc_510 N_VPWR_c_621_n N_A_592_367#_M1011_s 0.00536646f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_511 N_VPWR_c_621_n N_A_592_367#_M1026_s 0.00376627f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_621_n N_A_592_367#_M1014_d 0.00223565f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_621_n N_A_592_367#_M1037_d 0.00223562f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_514 N_VPWR_M1023_d N_A_592_367#_c_906_n 0.00344712f $X=3.39 $Y=1.835 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_626_n N_A_592_367#_c_906_n 0.0170777f $X=3.53 $Y=2.75 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_633_n N_A_592_367#_c_910_n 0.0361172f $X=6.05 $Y=3.33 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_621_n N_A_592_367#_c_910_n 0.023676f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_518 N_VPWR_c_633_n N_A_592_367#_c_922_n 0.0125234f $X=6.05 $Y=3.33 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_621_n N_A_592_367#_c_922_n 0.00738676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_627_n N_A_592_367#_c_908_n 0.0121156f $X=6.215 $Y=2.435 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_633_n N_A_592_367#_c_908_n 0.0519089f $X=6.05 $Y=3.33 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_621_n N_A_592_367#_c_908_n 0.0335966f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_627_n N_A_592_367#_c_909_n 0.0396f $X=6.215 $Y=2.435 $X2=0 $Y2=0
cc_524 N_VPWR_c_636_n N_A_592_367#_c_928_n 0.0124525f $X=3.365 $Y=3.33 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_621_n N_A_592_367#_c_928_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_633_n N_A_592_367#_c_930_n 0.0125234f $X=6.05 $Y=3.33 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_621_n N_A_592_367#_c_930_n 0.00738676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_621_n N_A_1317_367#_M1016_d 0.00223562f $X=9.84 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_529 N_VPWR_c_621_n N_A_1317_367#_M1008_s 0.00223565f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_621_n N_A_1317_367#_M1034_s 0.00404775f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_621_n N_A_1317_367#_M1029_d 0.0041489f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_637_n N_A_1317_367#_c_956_n 0.0361172f $X=8.745 $Y=3.33 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_621_n N_A_1317_367#_c_956_n 0.023676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_637_n N_A_1317_367#_c_948_n 0.015759f $X=8.745 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_621_n N_A_1317_367#_c_948_n 0.00991594f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_637_n N_A_1317_367#_c_958_n 0.0379702f $X=8.745 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_621_n N_A_1317_367#_c_958_n 0.0249919f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_637_n N_A_1317_367#_c_973_n 0.0129414f $X=8.745 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_621_n N_A_1317_367#_c_973_n 0.00738676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_M1017_s N_A_1317_367#_c_945_n 0.00176461f $X=8.77 $Y=1.835 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_628_n N_A_1317_367#_c_945_n 0.0170777f $X=8.91 $Y=2.115 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_630_n N_A_1317_367#_c_945_n 0.00166618f $X=9.77 $Y=1.98 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_638_n N_A_1317_367#_c_978_n 0.0136943f $X=9.64 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_621_n N_A_1317_367#_c_978_n 0.00866972f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_637_n N_A_1317_367#_c_980_n 0.0125234f $X=8.745 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_621_n N_A_1317_367#_c_980_n 0.00738676f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_Y_c_807_n N_A_592_367#_M1011_s 0.00334047f $X=4.225 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_548 N_Y_c_807_n N_A_592_367#_M1026_s 0.00353353f $X=4.225 $Y=2.04 $X2=0 $Y2=0
cc_549 N_Y_c_812_n N_A_592_367#_M1014_d 0.00344507f $X=5.085 $Y=2.045 $X2=0
+ $Y2=0
cc_550 Y N_A_592_367#_M1037_d 0.00353977f $X=6.395 $Y=1.95 $X2=0 $Y2=0
cc_551 N_Y_c_807_n N_A_592_367#_c_906_n 0.0323235f $X=4.225 $Y=2.04 $X2=0 $Y2=0
cc_552 N_Y_c_807_n N_A_592_367#_c_937_n 0.0135055f $X=4.225 $Y=2.04 $X2=0 $Y2=0
cc_553 N_Y_M1006_s N_A_592_367#_c_910_n 0.00332344f $X=4.25 $Y=1.835 $X2=0 $Y2=0
cc_554 N_Y_c_814_n N_A_592_367#_c_910_n 0.0159805f $X=4.39 $Y=2.04 $X2=0 $Y2=0
cc_555 N_Y_c_812_n N_A_592_367#_c_940_n 0.0129902f $X=5.085 $Y=2.045 $X2=0 $Y2=0
cc_556 N_Y_M1020_s N_A_592_367#_c_908_n 0.00332344f $X=5.11 $Y=1.835 $X2=0 $Y2=0
cc_557 N_Y_c_816_n N_A_592_367#_c_908_n 0.0159805f $X=5.25 $Y=2.04 $X2=0 $Y2=0
cc_558 Y N_A_592_367#_c_909_n 0.015351f $X=6.395 $Y=1.95 $X2=0 $Y2=0
cc_559 N_Y_c_807_n N_A_592_367#_c_928_n 0.0135055f $X=4.225 $Y=2.04 $X2=0 $Y2=0
cc_560 N_Y_c_834_n N_A_1317_367#_M1016_d 0.0078731f $X=7.32 $Y=2.042 $X2=-0.19
+ $Y2=-0.245
cc_561 N_Y_c_837_n N_A_1317_367#_M1008_s 0.00344607f $X=7.85 $Y=2.035 $X2=0
+ $Y2=0
cc_562 N_Y_c_834_n N_A_1317_367#_c_947_n 0.0153796f $X=7.32 $Y=2.042 $X2=0 $Y2=0
cc_563 N_Y_M1000_d N_A_1317_367#_c_956_n 0.00332344f $X=7.015 $Y=1.835 $X2=0
+ $Y2=0
cc_564 N_Y_c_833_n N_A_1317_367#_c_956_n 0.0158272f $X=7.155 $Y=2.035 $X2=0
+ $Y2=0
cc_565 N_Y_c_837_n N_A_1317_367#_c_987_n 0.0135055f $X=7.85 $Y=2.035 $X2=0 $Y2=0
cc_566 N_Y_M1028_d N_A_1317_367#_c_958_n 0.00332344f $X=7.875 $Y=1.835 $X2=0
+ $Y2=0
cc_567 N_Y_c_840_n N_A_1317_367#_c_958_n 0.0159805f $X=8.015 $Y=2.035 $X2=0
+ $Y2=0
cc_568 N_Y_c_840_n N_A_1317_367#_c_960_n 0.0512449f $X=8.015 $Y=2.035 $X2=0
+ $Y2=0
cc_569 N_Y_c_765_n N_A_29_65#_M1018_s 0.00274146f $X=1.535 $Y=1.17 $X2=0 $Y2=0
cc_570 N_Y_c_767_n N_A_29_65#_M1032_s 0.00258276f $X=2.46 $Y=1.17 $X2=0 $Y2=0
cc_571 N_Y_c_766_n N_A_29_65#_c_991_n 0.00497809f $X=0.865 $Y=1.17 $X2=0 $Y2=0
cc_572 N_Y_M1005_d N_A_29_65#_c_992_n 0.00176461f $X=0.56 $Y=0.325 $X2=0 $Y2=0
cc_573 N_Y_c_771_n N_A_29_65#_c_992_n 0.0159436f $X=0.7 $Y=0.7 $X2=0 $Y2=0
cc_574 N_Y_c_765_n N_A_29_65#_c_992_n 0.00272017f $X=1.535 $Y=1.17 $X2=0 $Y2=0
cc_575 N_Y_c_765_n N_A_29_65#_c_1005_n 0.0192603f $X=1.535 $Y=1.17 $X2=0 $Y2=0
cc_576 N_Y_M1021_d N_A_29_65#_c_994_n 0.00261503f $X=1.5 $Y=0.325 $X2=0 $Y2=0
cc_577 N_Y_c_765_n N_A_29_65#_c_994_n 0.00293866f $X=1.535 $Y=1.17 $X2=0 $Y2=0
cc_578 N_Y_c_784_n N_A_29_65#_c_994_n 0.018928f $X=1.7 $Y=0.7 $X2=0 $Y2=0
cc_579 N_Y_c_767_n N_A_29_65#_c_994_n 0.00315715f $X=2.46 $Y=1.17 $X2=0 $Y2=0
cc_580 N_Y_c_767_n N_A_29_65#_c_995_n 0.0202513f $X=2.46 $Y=1.17 $X2=0 $Y2=0
cc_581 N_Y_c_767_n N_A_29_65#_c_996_n 0.0390813f $X=2.46 $Y=1.17 $X2=0 $Y2=0
cc_582 N_A_29_65#_c_996_n N_A_509_47#_M1002_d 0.00895634f $X=2.81 $Y=0.785
+ $X2=-0.19 $Y2=-0.245
cc_583 N_A_29_65#_c_997_n N_A_509_47#_M1003_d 0.00177993f $X=3.865 $Y=1.117
+ $X2=0 $Y2=0
cc_584 N_A_29_65#_c_1024_n N_A_509_47#_M1012_s 0.00331141f $X=5.515 $Y=0.845
+ $X2=0 $Y2=0
cc_585 N_A_29_65#_c_1024_n N_A_509_47#_M1030_s 0.00331141f $X=5.515 $Y=0.845
+ $X2=0 $Y2=0
cc_586 N_A_29_65#_M1002_s N_A_509_47#_c_1084_n 0.00335455f $X=2.96 $Y=0.235
+ $X2=0 $Y2=0
cc_587 N_A_29_65#_c_994_n N_A_509_47#_c_1084_n 0.0146291f $X=2.035 $Y=0.34 $X2=0
+ $Y2=0
cc_588 N_A_29_65#_c_995_n N_A_509_47#_c_1084_n 0.00473042f $X=2.175 $Y=0.655
+ $X2=0 $Y2=0
cc_589 N_A_29_65#_c_996_n N_A_509_47#_c_1084_n 0.0419143f $X=2.81 $Y=0.785 $X2=0
+ $Y2=0
cc_590 N_A_29_65#_c_997_n N_A_509_47#_c_1084_n 0.00352369f $X=3.865 $Y=1.117
+ $X2=0 $Y2=0
cc_591 N_A_29_65#_M1013_d N_A_509_47#_c_1098_n 0.00330409f $X=4.68 $Y=0.235
+ $X2=0 $Y2=0
cc_592 N_A_29_65#_c_1024_n N_A_509_47#_c_1100_n 0.0593348f $X=5.515 $Y=0.845
+ $X2=0 $Y2=0
cc_593 N_A_29_65#_M1031_d N_A_509_47#_c_1090_n 0.00355031f $X=5.54 $Y=0.235
+ $X2=0 $Y2=0
cc_594 N_A_29_65#_c_1022_n N_A_509_47#_c_1090_n 0.0124003f $X=5.68 $Y=0.83 $X2=0
+ $Y2=0
cc_595 N_A_29_65#_c_1024_n N_A_509_47#_c_1090_n 0.00270524f $X=5.515 $Y=0.845
+ $X2=0 $Y2=0
cc_596 N_A_29_65#_c_1022_n N_A_509_47#_c_1091_n 0.0193773f $X=5.68 $Y=0.83 $X2=0
+ $Y2=0
cc_597 N_A_29_65#_c_997_n N_A_509_47#_c_1094_n 0.0171894f $X=3.865 $Y=1.117
+ $X2=0 $Y2=0
cc_598 N_A_29_65#_M1015_s N_A_509_47#_c_1097_n 0.00333487f $X=3.82 $Y=0.235
+ $X2=0 $Y2=0
cc_599 N_A_29_65#_c_997_n N_A_509_47#_c_1097_n 0.00326378f $X=3.865 $Y=1.117
+ $X2=0 $Y2=0
cc_600 N_A_29_65#_c_999_n N_A_509_47#_c_1097_n 0.0136982f $X=3.99 $Y=0.9 $X2=0
+ $Y2=0
cc_601 N_A_29_65#_c_1024_n N_A_509_47#_c_1097_n 0.00306864f $X=5.515 $Y=0.845
+ $X2=0 $Y2=0
cc_602 N_A_29_65#_c_992_n N_VGND_c_1195_n 0.0422287f $X=1.035 $Y=0.34 $X2=0
+ $Y2=0
cc_603 N_A_29_65#_c_993_n N_VGND_c_1195_n 0.0186386f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_604 N_A_29_65#_c_994_n N_VGND_c_1195_n 0.0623021f $X=2.035 $Y=0.34 $X2=0
+ $Y2=0
cc_605 N_A_29_65#_c_996_n N_VGND_c_1195_n 0.00341695f $X=2.81 $Y=0.785 $X2=0
+ $Y2=0
cc_606 N_A_29_65#_c_998_n N_VGND_c_1195_n 0.0234966f $X=1.2 $Y=0.34 $X2=0 $Y2=0
cc_607 N_A_29_65#_M1002_s N_VGND_c_1200_n 0.00225186f $X=2.96 $Y=0.235 $X2=0
+ $Y2=0
cc_608 N_A_29_65#_M1015_s N_VGND_c_1200_n 0.00225186f $X=3.82 $Y=0.235 $X2=0
+ $Y2=0
cc_609 N_A_29_65#_M1013_d N_VGND_c_1200_n 0.00225186f $X=4.68 $Y=0.235 $X2=0
+ $Y2=0
cc_610 N_A_29_65#_M1031_d N_VGND_c_1200_n 0.00225186f $X=5.54 $Y=0.235 $X2=0
+ $Y2=0
cc_611 N_A_29_65#_c_992_n N_VGND_c_1200_n 0.0238173f $X=1.035 $Y=0.34 $X2=0
+ $Y2=0
cc_612 N_A_29_65#_c_993_n N_VGND_c_1200_n 0.0101082f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_613 N_A_29_65#_c_994_n N_VGND_c_1200_n 0.0347633f $X=2.035 $Y=0.34 $X2=0
+ $Y2=0
cc_614 N_A_29_65#_c_996_n N_VGND_c_1200_n 0.0060615f $X=2.81 $Y=0.785 $X2=0
+ $Y2=0
cc_615 N_A_29_65#_c_998_n N_VGND_c_1200_n 0.0127407f $X=1.2 $Y=0.34 $X2=0 $Y2=0
cc_616 N_A_509_47#_c_1107_n N_VGND_M1007_d 0.0034577f $X=7.06 $Y=0.82 $X2=-0.19
+ $Y2=-0.245
cc_617 N_A_509_47#_c_1111_n N_VGND_M1025_d 0.00335437f $X=7.92 $Y=0.82 $X2=0
+ $Y2=0
cc_618 N_A_509_47#_c_1112_n N_VGND_M1039_d 0.00349176f $X=8.76 $Y=0.82 $X2=0
+ $Y2=0
cc_619 N_A_509_47#_c_1085_n N_VGND_M1027_d 0.00329816f $X=9.64 $Y=0.955 $X2=0
+ $Y2=0
cc_620 N_A_509_47#_c_1107_n N_VGND_c_1190_n 0.016459f $X=7.06 $Y=0.82 $X2=0
+ $Y2=0
cc_621 N_A_509_47#_c_1107_n N_VGND_c_1191_n 0.00196209f $X=7.06 $Y=0.82 $X2=0
+ $Y2=0
cc_622 N_A_509_47#_c_1153_p N_VGND_c_1191_n 0.0124139f $X=7.155 $Y=0.42 $X2=0
+ $Y2=0
cc_623 N_A_509_47#_c_1111_n N_VGND_c_1191_n 0.00196209f $X=7.92 $Y=0.82 $X2=0
+ $Y2=0
cc_624 N_A_509_47#_c_1111_n N_VGND_c_1192_n 0.016459f $X=7.92 $Y=0.82 $X2=0
+ $Y2=0
cc_625 N_A_509_47#_c_1112_n N_VGND_c_1193_n 0.016459f $X=8.76 $Y=0.82 $X2=0
+ $Y2=0
cc_626 N_A_509_47#_c_1085_n N_VGND_c_1194_n 0.0170777f $X=9.64 $Y=0.955 $X2=0
+ $Y2=0
cc_627 N_A_509_47#_c_1084_n N_VGND_c_1195_n 0.0500591f $X=3.365 $Y=0.37 $X2=0
+ $Y2=0
cc_628 N_A_509_47#_c_1159_p N_VGND_c_1195_n 0.0227821f $X=6.225 $Y=0.445 $X2=0
+ $Y2=0
cc_629 N_A_509_47#_c_1107_n N_VGND_c_1195_n 0.00196761f $X=7.06 $Y=0.82 $X2=0
+ $Y2=0
cc_630 N_A_509_47#_c_1094_n N_VGND_c_1195_n 0.0188892f $X=3.53 $Y=0.38 $X2=0
+ $Y2=0
cc_631 N_A_509_47#_c_1097_n N_VGND_c_1195_n 0.133361f $X=4.285 $Y=0.43 $X2=0
+ $Y2=0
cc_632 N_A_509_47#_c_1111_n N_VGND_c_1197_n 0.00196209f $X=7.92 $Y=0.82 $X2=0
+ $Y2=0
cc_633 N_A_509_47#_c_1164_p N_VGND_c_1197_n 0.0124139f $X=8.015 $Y=0.42 $X2=0
+ $Y2=0
cc_634 N_A_509_47#_c_1112_n N_VGND_c_1197_n 0.00196209f $X=8.76 $Y=0.82 $X2=0
+ $Y2=0
cc_635 N_A_509_47#_c_1112_n N_VGND_c_1198_n 0.00181088f $X=8.76 $Y=0.82 $X2=0
+ $Y2=0
cc_636 N_A_509_47#_c_1167_p N_VGND_c_1198_n 0.0124525f $X=8.875 $Y=0.42 $X2=0
+ $Y2=0
cc_637 N_A_509_47#_c_1086_n N_VGND_c_1199_n 0.0178111f $X=9.735 $Y=0.42 $X2=0
+ $Y2=0
cc_638 N_A_509_47#_M1002_d N_VGND_c_1200_n 0.00215176f $X=2.545 $Y=0.235 $X2=0
+ $Y2=0
cc_639 N_A_509_47#_M1003_d N_VGND_c_1200_n 0.00223559f $X=3.39 $Y=0.235 $X2=0
+ $Y2=0
cc_640 N_A_509_47#_M1012_s N_VGND_c_1200_n 0.00223577f $X=4.25 $Y=0.235 $X2=0
+ $Y2=0
cc_641 N_A_509_47#_M1030_s N_VGND_c_1200_n 0.00223577f $X=5.11 $Y=0.235 $X2=0
+ $Y2=0
cc_642 N_A_509_47#_M1019_d N_VGND_c_1200_n 0.00400243f $X=5.97 $Y=0.235 $X2=0
+ $Y2=0
cc_643 N_A_509_47#_M1009_s N_VGND_c_1200_n 0.00266476f $X=7.015 $Y=0.235 $X2=0
+ $Y2=0
cc_644 N_A_509_47#_M1038_s N_VGND_c_1200_n 0.00266476f $X=7.875 $Y=0.235 $X2=0
+ $Y2=0
cc_645 N_A_509_47#_M1022_s N_VGND_c_1200_n 0.00400223f $X=8.735 $Y=0.235 $X2=0
+ $Y2=0
cc_646 N_A_509_47#_M1035_s N_VGND_c_1200_n 0.00371702f $X=9.595 $Y=0.235 $X2=0
+ $Y2=0
cc_647 N_A_509_47#_c_1084_n N_VGND_c_1200_n 0.031218f $X=3.365 $Y=0.37 $X2=0
+ $Y2=0
cc_648 N_A_509_47#_c_1159_p N_VGND_c_1200_n 0.0128285f $X=6.225 $Y=0.445 $X2=0
+ $Y2=0
cc_649 N_A_509_47#_c_1107_n N_VGND_c_1200_n 0.00896404f $X=7.06 $Y=0.82 $X2=0
+ $Y2=0
cc_650 N_A_509_47#_c_1153_p N_VGND_c_1200_n 0.00730033f $X=7.155 $Y=0.42 $X2=0
+ $Y2=0
cc_651 N_A_509_47#_c_1111_n N_VGND_c_1200_n 0.00891615f $X=7.92 $Y=0.82 $X2=0
+ $Y2=0
cc_652 N_A_509_47#_c_1164_p N_VGND_c_1200_n 0.00730033f $X=8.015 $Y=0.42 $X2=0
+ $Y2=0
cc_653 N_A_509_47#_c_1112_n N_VGND_c_1200_n 0.00839284f $X=8.76 $Y=0.82 $X2=0
+ $Y2=0
cc_654 N_A_509_47#_c_1167_p N_VGND_c_1200_n 0.00730901f $X=8.875 $Y=0.42 $X2=0
+ $Y2=0
cc_655 N_A_509_47#_c_1086_n N_VGND_c_1200_n 0.0100304f $X=9.735 $Y=0.42 $X2=0
+ $Y2=0
cc_656 N_A_509_47#_c_1094_n N_VGND_c_1200_n 0.0124024f $X=3.53 $Y=0.38 $X2=0
+ $Y2=0
cc_657 N_A_509_47#_c_1097_n N_VGND_c_1200_n 0.0853926f $X=4.285 $Y=0.43 $X2=0
+ $Y2=0
cc_658 N_A_509_47#_c_1121_n N_VGND_c_1200_n 5.15613e-19 $X=8.865 $Y=0.82 $X2=0
+ $Y2=0
