# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor4bb_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nor4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.795000 1.375000 9.495000 1.760000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.785000 1.355000 7.475000 1.525000 ;
        RECT 5.785000 1.525000 6.205000 1.830000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.345000 1.285000 1.760000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.375000 0.475000 1.760000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.587200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 0.255000 2.365000 0.655000 ;
        RECT 2.025000 0.655000 4.245000 0.825000 ;
        RECT 2.195000 1.685000 5.615000 1.855000 ;
        RECT 2.195000 1.855000 2.385000 2.735000 ;
        RECT 3.055000 0.255000 3.385000 0.655000 ;
        RECT 3.055000 1.855000 5.615000 1.865000 ;
        RECT 3.055000 1.865000 3.285000 2.735000 ;
        RECT 4.055000 0.255000 4.245000 0.655000 ;
        RECT 4.060000 0.825000 4.245000 0.995000 ;
        RECT 4.060000 0.995000 6.350000 1.005000 ;
        RECT 4.060000 1.005000 8.965000 1.165000 ;
        RECT 4.915000 0.255000 5.105000 0.985000 ;
        RECT 4.915000 0.985000 6.350000 0.995000 ;
        RECT 5.250000 1.165000 8.965000 1.175000 ;
        RECT 5.250000 1.175000 5.615000 1.685000 ;
        RECT 6.160000 0.255000 6.350000 0.985000 ;
        RECT 7.020000 0.255000 7.210000 1.005000 ;
        RECT 7.880000 0.255000 8.070000 1.005000 ;
        RECT 8.740000 0.255000 8.965000 1.005000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
        RECT 0.575000  0.085000 0.905000 0.855000 ;
        RECT 1.525000  0.085000 1.855000 0.815000 ;
        RECT 2.535000  0.085000 2.865000 0.485000 ;
        RECT 3.555000  0.085000 3.885000 0.485000 ;
        RECT 4.415000  0.085000 4.745000 0.825000 ;
        RECT 5.275000  0.085000 5.990000 0.815000 ;
        RECT 6.520000  0.085000 6.850000 0.835000 ;
        RECT 7.380000  0.085000 7.710000 0.835000 ;
        RECT 8.240000  0.085000 8.570000 0.835000 ;
        RECT 9.135000  0.085000 9.430000 1.095000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.600000 3.415000 ;
        RECT 0.575000 2.650000 0.905000 3.245000 ;
        RECT 7.810000 2.270000 8.140000 3.245000 ;
        RECT 8.670000 2.270000 9.000000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.145000 0.255000 0.395000 1.025000 ;
      RECT 0.145000 1.025000 0.825000 1.195000 ;
      RECT 0.145000 1.930000 0.825000 2.310000 ;
      RECT 0.145000 2.310000 2.025000 2.480000 ;
      RECT 0.145000 2.480000 0.405000 3.075000 ;
      RECT 0.645000 1.195000 0.825000 1.930000 ;
      RECT 1.005000 1.930000 1.635000 2.140000 ;
      RECT 1.075000 0.255000 1.335000 0.995000 ;
      RECT 1.075000 0.995000 3.890000 1.165000 ;
      RECT 1.075000 1.165000 1.635000 1.175000 ;
      RECT 1.455000 1.175000 1.635000 1.930000 ;
      RECT 1.695000 2.650000 2.025000 2.905000 ;
      RECT 1.695000 2.905000 3.675000 3.075000 ;
      RECT 1.820000 1.335000 3.510000 1.515000 ;
      RECT 1.820000 1.515000 2.025000 2.310000 ;
      RECT 2.555000 2.025000 2.885000 2.905000 ;
      RECT 3.455000 2.035000 5.465000 2.205000 ;
      RECT 3.455000 2.205000 3.675000 2.905000 ;
      RECT 3.720000 1.165000 3.890000 1.335000 ;
      RECT 3.720000 1.335000 5.070000 1.515000 ;
      RECT 3.845000 2.375000 4.175000 2.905000 ;
      RECT 3.845000 2.905000 7.275000 3.075000 ;
      RECT 4.345000 2.205000 4.535000 2.735000 ;
      RECT 4.705000 2.375000 5.035000 2.885000 ;
      RECT 4.705000 2.885000 7.275000 2.905000 ;
      RECT 5.205000 2.205000 5.465000 2.715000 ;
      RECT 5.655000 2.035000 6.775000 2.205000 ;
      RECT 5.655000 2.205000 5.915000 2.715000 ;
      RECT 6.085000 2.375000 6.415000 2.885000 ;
      RECT 6.515000 1.705000 7.625000 1.875000 ;
      RECT 6.515000 1.875000 6.775000 2.035000 ;
      RECT 6.585000 2.205000 6.775000 2.715000 ;
      RECT 6.945000 2.055000 7.275000 2.885000 ;
      RECT 7.445000 1.875000 7.625000 1.930000 ;
      RECT 7.445000 1.930000 9.430000 2.100000 ;
      RECT 7.445000 2.100000 7.640000 3.075000 ;
      RECT 8.310000 2.100000 8.500000 3.075000 ;
      RECT 9.170000 2.100000 9.430000 3.075000 ;
  END
END sky130_fd_sc_lp__nor4bb_4
