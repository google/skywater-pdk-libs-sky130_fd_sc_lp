* File: sky130_fd_sc_lp__a21o_2.pex.spice
* Created: Wed Sep  2 09:20:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21O_2%A_86_269# 1 2 9 13 17 21 24 27 28 29 30 31 33
+ 37 40 42 48
r80 41 48 2.02521 $w=2.38e-07 $l=1e-08 $layer=POLY_cond $X=1.115 $Y=1.585
+ $X2=1.105 $Y2=1.585
r81 40 42 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=1.51
+ $X2=1.155 $Y2=1.345
r82 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.51 $X2=1.115 $Y2=1.51
r83 35 37 32.9809 $w=1.88e-07 $l=5.65e-07 $layer=LI1_cond $X=1.8 $Y=0.985
+ $X2=1.8 $Y2=0.42
r84 31 44 2.68365 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.662 $Y=2.1
+ $X2=1.662 $Y2=2.015
r85 31 33 29.6342 $w=3.13e-07 $l=8.1e-07 $layer=LI1_cond $X=1.662 $Y=2.1
+ $X2=1.662 $Y2=2.91
r86 29 44 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.505 $Y=2.015
+ $X2=1.662 $Y2=2.015
r87 29 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.505 $Y=2.015
+ $X2=1.325 $Y2=2.015
r88 27 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.705 $Y=1.07
+ $X2=1.8 $Y2=0.985
r89 27 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.705 $Y=1.07
+ $X2=1.325 $Y2=1.07
r90 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.24 $Y=1.155
+ $X2=1.325 $Y2=1.07
r91 25 42 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.24 $Y=1.155
+ $X2=1.24 $Y2=1.345
r92 24 30 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.155 $Y=1.93
+ $X2=1.325 $Y2=2.015
r93 23 40 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=1.155 $Y=1.515
+ $X2=1.155 $Y2=1.51
r94 23 24 14.0666 $w=3.38e-07 $l=4.15e-07 $layer=LI1_cond $X=1.155 $Y=1.515
+ $X2=1.155 $Y2=1.93
r95 19 48 13.5836 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.105 $Y=1.345
+ $X2=1.105 $Y2=1.585
r96 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.105 $Y=1.345
+ $X2=1.105 $Y2=0.655
r97 15 48 34.4286 $w=2.38e-07 $l=1.7e-07 $layer=POLY_cond $X=0.935 $Y=1.585
+ $X2=1.105 $Y2=1.585
r98 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.935 $Y=1.675
+ $X2=0.935 $Y2=2.465
r99 11 15 52.6555 $w=2.38e-07 $l=3.60555e-07 $layer=POLY_cond $X=0.675 $Y=1.345
+ $X2=0.935 $Y2=1.585
r100 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.675 $Y=1.345
+ $X2=0.675 $Y2=0.655
r101 7 11 34.4286 $w=2.38e-07 $l=2.33238e-07 $layer=POLY_cond $X=0.505 $Y=1.495
+ $X2=0.675 $Y2=1.345
r102 7 9 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.505 $Y=1.495
+ $X2=0.505 $Y2=2.465
r103 2 44 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.835 $X2=1.67 $Y2=2.095
r104 2 33 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.835 $X2=1.67 $Y2=2.91
r105 1 37 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.67
+ $Y=0.235 $X2=1.81 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_2%B1 3 7 9 13 14
c38 14 0 1.7811e-19 $X=1.685 $Y=1.51
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.685
+ $Y=1.51 $X2=1.685 $Y2=1.51
r40 11 13 15.2211 $w=2.85e-07 $l=9e-08 $layer=POLY_cond $X=1.595 $Y=1.51
+ $X2=1.685 $Y2=1.51
r41 9 14 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=1.657 $Y=1.665
+ $X2=1.657 $Y2=1.51
r42 5 13 33.8246 $w=2.85e-07 $l=2.70185e-07 $layer=POLY_cond $X=1.885 $Y=1.675
+ $X2=1.685 $Y2=1.51
r43 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.885 $Y=1.675
+ $X2=1.885 $Y2=2.465
r44 1 11 17.7656 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.345
+ $X2=1.595 $Y2=1.51
r45 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.595 $Y=1.345
+ $X2=1.595 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_2%A1 3 6 8 9 10 21 23
c37 21 0 1.7811e-19 $X=2.335 $Y=1.35
r38 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.35
+ $X2=2.335 $Y2=1.515
r39 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.35
+ $X2=2.335 $Y2=1.185
r40 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.335
+ $Y=1.35 $X2=2.335 $Y2=1.35
r41 10 22 0.981855 $w=6.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.4 $Y=1.295
+ $X2=2.4 $Y2=1.35
r42 9 10 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.4 $Y=0.925 $X2=2.4
+ $Y2=1.295
r43 8 9 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.4 $Y=0.555 $X2=2.4
+ $Y2=0.925
r44 6 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.315 $Y=2.465
+ $X2=2.315 $Y2=1.515
r45 3 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.245 $Y=0.655
+ $X2=2.245 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_2%A2 1 3 6 8 13
r23 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.35 $X2=2.99 $Y2=1.35
r24 10 13 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.785 $Y=1.35
+ $X2=2.99 $Y2=1.35
r25 8 14 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.35 $X2=2.99
+ $Y2=1.35
r26 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.515
+ $X2=2.785 $Y2=1.35
r27 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.785 $Y=1.515
+ $X2=2.785 $Y2=2.465
r28 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.185
+ $X2=2.785 $Y2=1.35
r29 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.785 $Y=1.185
+ $X2=2.785 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_2%VPWR 1 2 3 10 12 18 22 27 28 29 31 41 42 48
r48 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.15 $Y2=3.33
r54 36 38 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 32 45 4.34571 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.207 $Y2=3.33
r59 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.15 $Y2=3.33
r61 31 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 29 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 29 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 27 38 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.55 $Y2=3.33
r66 26 41 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.715 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=3.33
+ $X2=2.55 $Y2=3.33
r68 22 25 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.55 $Y=2.11
+ $X2=2.55 $Y2=2.95
r69 20 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=3.245
+ $X2=2.55 $Y2=3.33
r70 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.55 $Y=3.245
+ $X2=2.55 $Y2=2.95
r71 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=3.33
r72 16 18 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=2.385
r73 12 15 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=0.27 $Y=1.98
+ $X2=0.27 $Y2=2.95
r74 10 45 3.09214 $w=2.9e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.207 $Y2=3.33
r75 10 15 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.95
r76 3 25 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.835 $X2=2.55 $Y2=2.95
r77 3 22 400 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.835 $X2=2.55 $Y2=2.11
r78 2 18 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=2.385
r79 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.95
r80 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_2%X 1 2 9 14 16 17 18 19 20
r21 20 38 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.7 $Y=2.775
+ $X2=0.7 $Y2=2.91
r22 19 20 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=2.405 $X2=0.7
+ $Y2=2.775
r23 18 19 21.2951 $w=2.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.7 $Y=1.98 $X2=0.7
+ $Y2=2.405
r24 17 18 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.7 $Y=1.665
+ $X2=0.7 $Y2=1.98
r25 16 17 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=1.295 $X2=0.7
+ $Y2=1.665
r26 12 16 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.7 $Y=1.155 $X2=0.7
+ $Y2=1.295
r27 12 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.7 $Y=1.07 $X2=0.89
+ $Y2=1.07
r28 7 14 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=0.985
+ $X2=0.89 $Y2=1.07
r29 7 9 32.9809 $w=1.88e-07 $l=5.65e-07 $layer=LI1_cond $X=0.89 $Y=0.985
+ $X2=0.89 $Y2=0.42
r30 2 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.91
r31 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=1.98
r32 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.75
+ $Y=0.235 $X2=0.89 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_2%A_392_367# 1 2 9 13 14 17
r21 17 19 48.7169 $w=2.18e-07 $l=9.3e-07 $layer=LI1_cond $X=2.995 $Y=1.98
+ $X2=2.995 $Y2=2.91
r22 15 17 6.54797 $w=2.18e-07 $l=1.25e-07 $layer=LI1_cond $X=2.995 $Y=1.855
+ $X2=2.995 $Y2=1.98
r23 13 15 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.885 $Y=1.77
+ $X2=2.995 $Y2=1.855
r24 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.885 $Y=1.77
+ $X2=2.215 $Y2=1.77
r25 9 11 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=2.102 $Y=1.98
+ $X2=2.102 $Y2=2.91
r26 7 14 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=2.102 $Y=1.855
+ $X2=2.215 $Y2=1.77
r27 7 9 6.40246 $w=2.23e-07 $l=1.25e-07 $layer=LI1_cond $X=2.102 $Y=1.855
+ $X2=2.102 $Y2=1.98
r28 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.835 $X2=3 $Y2=2.91
r29 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.835 $X2=3 $Y2=1.98
r30 1 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=2.91
r31 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_2%VGND 1 2 3 12 14 18 20 22 24 25 26 31 40 44
r44 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r47 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r49 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.32
+ $Y2=0
r50 32 34 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.68
+ $Y2=0
r51 31 43 4.09313 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.132
+ $Y2=0
r52 31 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r53 30 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r54 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 26 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r56 26 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r57 26 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 24 29 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.24
+ $Y2=0
r59 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.46
+ $Y2=0
r60 20 43 3.19156 $w=2.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.132 $Y2=0
r61 20 22 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0.38
r62 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=0.085
+ $X2=1.32 $Y2=0
r63 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.32 $Y=0.085
+ $X2=1.32 $Y2=0.36
r64 15 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.46
+ $Y2=0
r65 14 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.32
+ $Y2=0
r66 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=0.625
+ $Y2=0
r67 10 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.46 $Y=0.085
+ $X2=0.46 $Y2=0
r68 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.46 $Y=0.085
+ $X2=0.46 $Y2=0.38
r69 3 22 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=2.86
+ $Y=0.235 $X2=3.01 $Y2=0.38
r70 2 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.18
+ $Y=0.235 $X2=1.32 $Y2=0.36
r71 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.335
+ $Y=0.235 $X2=0.46 $Y2=0.38
.ends

