* File: sky130_fd_sc_lp__xor2_m.pxi.spice
* Created: Fri Aug 28 11:36:46 2020
* 
x_PM_SKY130_FD_SC_LP__XOR2_M%A N_A_c_70_n N_A_M1002_g N_A_M1009_g N_A_M1008_g
+ N_A_c_74_n N_A_M1007_g N_A_c_76_n A A N_A_c_78_n PM_SKY130_FD_SC_LP__XOR2_M%A
x_PM_SKY130_FD_SC_LP__XOR2_M%B N_B_M1000_g N_B_M1004_g N_B_c_119_n N_B_c_120_n
+ N_B_M1005_g N_B_c_126_n N_B_c_127_n N_B_M1006_g B B B N_B_c_122_n N_B_c_123_n
+ PM_SKY130_FD_SC_LP__XOR2_M%B
x_PM_SKY130_FD_SC_LP__XOR2_M%A_41_535# N_A_41_535#_M1000_d N_A_41_535#_M1004_s
+ N_A_41_535#_M1001_g N_A_41_535#_M1003_g N_A_41_535#_c_191_n
+ N_A_41_535#_c_192_n N_A_41_535#_c_193_n N_A_41_535#_c_184_n
+ N_A_41_535#_c_185_n N_A_41_535#_c_186_n N_A_41_535#_c_187_n
+ N_A_41_535#_c_197_n N_A_41_535#_c_188_n N_A_41_535#_c_189_n
+ PM_SKY130_FD_SC_LP__XOR2_M%A_41_535#
x_PM_SKY130_FD_SC_LP__XOR2_M%VPWR N_VPWR_M1002_d N_VPWR_M1005_d N_VPWR_c_250_n
+ N_VPWR_c_251_n N_VPWR_c_252_n N_VPWR_c_253_n VPWR N_VPWR_c_254_n
+ N_VPWR_c_255_n N_VPWR_c_249_n N_VPWR_c_257_n PM_SKY130_FD_SC_LP__XOR2_M%VPWR
x_PM_SKY130_FD_SC_LP__XOR2_M%A_282_535# N_A_282_535#_M1008_d
+ N_A_282_535#_M1001_s N_A_282_535#_c_292_n N_A_282_535#_c_293_n
+ N_A_282_535#_c_294_n N_A_282_535#_c_295_n
+ PM_SKY130_FD_SC_LP__XOR2_M%A_282_535#
x_PM_SKY130_FD_SC_LP__XOR2_M%X N_X_M1006_d N_X_M1001_d N_X_c_322_n N_X_c_316_n X
+ X X X X PM_SKY130_FD_SC_LP__XOR2_M%X
x_PM_SKY130_FD_SC_LP__XOR2_M%VGND N_VGND_M1000_s N_VGND_M1009_d N_VGND_M1003_d
+ N_VGND_c_344_n N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n
+ VGND N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n
+ PM_SKY130_FD_SC_LP__XOR2_M%VGND
cc_1 VNB N_A_M1009_g 0.0373998f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.99
cc_2 VNB N_A_M1007_g 0.0319542f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=0.99
cc_3 VNB N_B_M1000_g 0.0575617f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.885
cc_4 VNB N_B_c_119_n 0.0898429f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.99
cc_5 VNB N_B_c_120_n 0.0100709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B_M1006_g 0.0331629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_122_n 0.0409285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_123_n 0.0133478f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.2
cc_9 VNB N_A_41_535#_M1003_g 0.0371246f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.78
cc_10 VNB N_A_41_535#_c_184_n 0.00233604f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.78
cc_11 VNB N_A_41_535#_c_185_n 0.00766907f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_12 VNB N_A_41_535#_c_186_n 0.00803677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_41_535#_c_187_n 0.0251251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_41_535#_c_188_n 5.16948e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.2
cc_15 VNB N_A_41_535#_c_189_n 0.012192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_249_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.995
cc_17 VNB N_X_c_316_n 0.0031675f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.885
cc_18 VNB X 0.0199906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB X 0.0134841f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.78
cc_20 VNB N_VGND_c_344_n 0.0130327f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.885
cc_21 VNB N_VGND_c_345_n 0.0314738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_346_n 0.0107611f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=0.99
cc_23 VNB N_VGND_c_347_n 0.0136522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_348_n 0.0492997f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.35
cc_25 VNB N_VGND_c_349_n 0.0199579f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_26 VNB N_VGND_c_350_n 0.0415057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_351_n 0.00628644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_352_n 0.236872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_A_c_70_n 0.0187485f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.5
cc_30 VPB N_A_M1002_g 0.0187687f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.885
cc_31 VPB N_A_M1009_g 0.0025117f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.99
cc_32 VPB N_A_M1008_g 0.0196005f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.885
cc_33 VPB N_A_c_74_n 0.0238812f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.78
cc_34 VPB N_A_M1007_g 0.00235679f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=0.99
cc_35 VPB N_A_c_76_n 0.018643f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.78
cc_36 VPB A 0.0110071f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_37 VPB N_A_c_78_n 0.047907f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.995
cc_38 VPB N_B_M1000_g 0.0693878f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.885
cc_39 VPB N_B_M1005_g 0.0431359f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.885
cc_40 VPB N_B_c_126_n 0.0200822f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.78
cc_41 VPB N_B_c_127_n 0.00873493f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=1.78
cc_42 VPB N_B_M1006_g 0.0248215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_41_535#_M1001_g 0.0346322f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.5
cc_44 VPB N_A_41_535#_c_191_n 0.0284186f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=0.99
cc_45 VPB N_A_41_535#_c_192_n 0.0201261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_41_535#_c_193_n 0.0464988f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.5
cc_47 VPB N_A_41_535#_c_184_n 0.00186127f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.78
cc_48 VPB N_A_41_535#_c_185_n 0.00323487f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_49 VPB N_A_41_535#_c_187_n 0.0187157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_41_535#_c_197_n 0.00195113f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.995
cc_51 VPB N_A_41_535#_c_188_n 8.49936e-19 $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.2
cc_52 VPB N_A_41_535#_c_189_n 0.00543279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_250_n 4.09336e-19 $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.5
cc_54 VPB N_VPWR_c_251_n 0.00433998f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.78
cc_55 VPB N_VPWR_c_252_n 0.0153555f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=0.99
cc_56 VPB N_VPWR_c_253_n 0.00401177f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=0.99
cc_57 VPB N_VPWR_c_254_n 0.0297839f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.35
cc_58 VPB N_VPWR_c_255_n 0.037794f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.995
cc_59 VPB N_VPWR_c_249_n 0.0652074f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.995
cc_60 VPB N_VPWR_c_257_n 0.00436274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_282_535#_c_292_n 0.00136178f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.5
cc_62 VPB N_A_282_535#_c_293_n 0.0186171f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.885
cc_63 VPB N_A_282_535#_c_294_n 0.00484272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_282_535#_c_295_n 0.0130392f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.78
cc_65 VPB X 0.0453112f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.78
cc_66 VPB X 0.0122453f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=0.99
cc_67 N_A_c_70_n N_B_M1000_g 0.0539835f $X=0.905 $Y=2.5 $X2=0 $Y2=0
cc_68 N_A_M1009_g N_B_M1000_g 0.0557829f $X=0.975 $Y=0.99 $X2=0 $Y2=0
cc_69 A N_B_M1000_g 0.00526056f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_70 N_A_M1009_g N_B_c_119_n 0.00930902f $X=0.975 $Y=0.99 $X2=0 $Y2=0
cc_71 N_A_M1007_g N_B_c_119_n 0.00825049f $X=1.71 $Y=0.99 $X2=0 $Y2=0
cc_72 N_A_c_70_n N_B_M1005_g 0.0186056f $X=0.905 $Y=2.5 $X2=0 $Y2=0
cc_73 N_A_c_74_n N_B_c_127_n 0.0060701f $X=1.635 $Y=1.78 $X2=0 $Y2=0
cc_74 A N_B_c_127_n 0.00173646f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_75 N_A_c_78_n N_B_c_127_n 0.0186056f $X=1.065 $Y=1.995 $X2=0 $Y2=0
cc_76 N_A_M1007_g N_B_M1006_g 0.0791381f $X=1.71 $Y=0.99 $X2=0 $Y2=0
cc_77 N_A_c_78_n N_B_M1006_g 0.0042528f $X=1.065 $Y=1.995 $X2=0 $Y2=0
cc_78 N_A_M1009_g N_B_c_123_n 0.00403102f $X=0.975 $Y=0.99 $X2=0 $Y2=0
cc_79 N_A_M1007_g N_B_c_123_n 0.0276463f $X=1.71 $Y=0.99 $X2=0 $Y2=0
cc_80 A N_A_41_535#_c_193_n 0.0439528f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_81 A N_A_41_535#_c_184_n 0.00155805f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_82 N_A_M1009_g N_A_41_535#_c_186_n 0.00913264f $X=0.975 $Y=0.99 $X2=0 $Y2=0
cc_83 N_A_M1009_g N_A_41_535#_c_187_n 0.0129459f $X=0.975 $Y=0.99 $X2=0 $Y2=0
cc_84 N_A_c_74_n N_A_41_535#_c_187_n 0.0153309f $X=1.635 $Y=1.78 $X2=0 $Y2=0
cc_85 N_A_M1007_g N_A_41_535#_c_187_n 0.00820936f $X=1.71 $Y=0.99 $X2=0 $Y2=0
cc_86 N_A_c_76_n N_A_41_535#_c_187_n 0.0170487f $X=1.155 $Y=1.78 $X2=0 $Y2=0
cc_87 A N_A_41_535#_c_187_n 0.0302583f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_88 A N_A_41_535#_c_197_n 0.0185886f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_89 N_A_c_70_n N_VPWR_c_250_n 0.00241335f $X=0.905 $Y=2.5 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_VPWR_c_250_n 0.00958161f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_91 N_A_M1008_g N_VPWR_c_250_n 0.00771798f $X=1.335 $Y=2.885 $X2=0 $Y2=0
cc_92 A N_VPWR_c_250_n 0.0109568f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_93 N_A_M1008_g N_VPWR_c_252_n 0.00486043f $X=1.335 $Y=2.885 $X2=0 $Y2=0
cc_94 N_A_M1002_g N_VPWR_c_254_n 0.00486043f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_95 N_A_M1002_g N_VPWR_c_249_n 0.00445138f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_96 N_A_M1008_g N_VPWR_c_249_n 0.00838234f $X=1.335 $Y=2.885 $X2=0 $Y2=0
cc_97 A N_VPWR_c_249_n 0.013004f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_98 N_A_M1008_g N_A_282_535#_c_292_n 0.001666f $X=1.335 $Y=2.885 $X2=0 $Y2=0
cc_99 N_A_c_74_n N_A_282_535#_c_293_n 0.00131838f $X=1.635 $Y=1.78 $X2=0 $Y2=0
cc_100 N_A_c_70_n N_A_282_535#_c_294_n 0.00421179f $X=0.905 $Y=2.5 $X2=0 $Y2=0
cc_101 N_A_c_74_n N_A_282_535#_c_294_n 0.0054282f $X=1.635 $Y=1.78 $X2=0 $Y2=0
cc_102 A N_A_282_535#_c_294_n 0.00459387f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_103 N_A_M1009_g N_VGND_c_346_n 0.00756372f $X=0.975 $Y=0.99 $X2=0 $Y2=0
cc_104 N_A_M1007_g N_VGND_c_346_n 0.0015332f $X=1.71 $Y=0.99 $X2=0 $Y2=0
cc_105 N_A_c_76_n N_VGND_c_346_n 0.00121536f $X=1.155 $Y=1.78 $X2=0 $Y2=0
cc_106 N_B_c_126_n N_A_41_535#_M1001_g 4.79799e-19 $X=1.995 $Y=2.17 $X2=0 $Y2=0
cc_107 N_B_M1006_g N_A_41_535#_M1003_g 0.0157219f $X=2.07 $Y=0.99 $X2=0 $Y2=0
cc_108 N_B_c_123_n N_A_41_535#_M1003_g 0.00334149f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_109 N_B_c_126_n N_A_41_535#_c_191_n 0.00944528f $X=1.995 $Y=2.17 $X2=0 $Y2=0
cc_110 N_B_M1000_g N_A_41_535#_c_193_n 0.0282361f $X=0.545 $Y=0.99 $X2=0 $Y2=0
cc_111 N_B_M1000_g N_A_41_535#_c_184_n 0.0208302f $X=0.545 $Y=0.99 $X2=0 $Y2=0
cc_112 N_B_M1000_g N_A_41_535#_c_186_n 0.00913264f $X=0.545 $Y=0.99 $X2=0 $Y2=0
cc_113 N_B_c_119_n N_A_41_535#_c_186_n 0.00420384f $X=1.995 $Y=0.335 $X2=0 $Y2=0
cc_114 N_B_c_127_n N_A_41_535#_c_187_n 0.00670019f $X=1.84 $Y=2.17 $X2=0 $Y2=0
cc_115 N_B_M1006_g N_A_41_535#_c_187_n 0.0150797f $X=2.07 $Y=0.99 $X2=0 $Y2=0
cc_116 N_B_c_123_n N_A_41_535#_c_187_n 0.0500474f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_117 N_B_M1006_g N_A_41_535#_c_188_n 0.00262123f $X=2.07 $Y=0.99 $X2=0 $Y2=0
cc_118 N_B_M1006_g N_A_41_535#_c_189_n 0.00944528f $X=2.07 $Y=0.99 $X2=0 $Y2=0
cc_119 N_B_M1000_g N_VPWR_c_250_n 0.00204405f $X=0.545 $Y=0.99 $X2=0 $Y2=0
cc_120 N_B_M1005_g N_VPWR_c_250_n 7.58747e-19 $X=1.765 $Y=2.885 $X2=0 $Y2=0
cc_121 N_B_M1005_g N_VPWR_c_251_n 0.00321113f $X=1.765 $Y=2.885 $X2=0 $Y2=0
cc_122 N_B_M1005_g N_VPWR_c_252_n 0.00437852f $X=1.765 $Y=2.885 $X2=0 $Y2=0
cc_123 N_B_M1000_g N_VPWR_c_254_n 0.00585385f $X=0.545 $Y=0.99 $X2=0 $Y2=0
cc_124 N_B_M1000_g N_VPWR_c_249_n 0.0118816f $X=0.545 $Y=0.99 $X2=0 $Y2=0
cc_125 N_B_M1005_g N_VPWR_c_249_n 0.00732232f $X=1.765 $Y=2.885 $X2=0 $Y2=0
cc_126 N_B_M1005_g N_A_282_535#_c_292_n 0.00170909f $X=1.765 $Y=2.885 $X2=0
+ $Y2=0
cc_127 N_B_M1005_g N_A_282_535#_c_293_n 0.0154423f $X=1.765 $Y=2.885 $X2=0 $Y2=0
cc_128 N_B_c_126_n N_A_282_535#_c_293_n 0.0112534f $X=1.995 $Y=2.17 $X2=0 $Y2=0
cc_129 N_B_M1005_g N_A_282_535#_c_295_n 0.00437921f $X=1.765 $Y=2.885 $X2=0
+ $Y2=0
cc_130 N_B_c_123_n N_X_M1006_d 0.00488566f $X=2.16 $Y=0.43 $X2=-0.19 $Y2=-0.245
cc_131 N_B_M1006_g N_X_c_322_n 9.61618e-19 $X=2.07 $Y=0.99 $X2=0 $Y2=0
cc_132 N_B_c_123_n N_X_c_322_n 0.0249265f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_133 N_B_M1006_g N_X_c_316_n 6.27847e-19 $X=2.07 $Y=0.99 $X2=0 $Y2=0
cc_134 N_B_c_123_n N_X_c_316_n 0.0151747f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_135 N_B_c_120_n N_VGND_c_345_n 0.0156657f $X=0.62 $Y=0.335 $X2=0 $Y2=0
cc_136 N_B_M1000_g N_VGND_c_346_n 0.00498409f $X=0.545 $Y=0.99 $X2=0 $Y2=0
cc_137 N_B_c_119_n N_VGND_c_346_n 0.0254786f $X=1.995 $Y=0.335 $X2=0 $Y2=0
cc_138 N_B_c_122_n N_VGND_c_346_n 5.75798e-19 $X=2.16 $Y=0.335 $X2=0 $Y2=0
cc_139 N_B_c_123_n N_VGND_c_346_n 0.0446952f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_140 N_B_c_122_n N_VGND_c_348_n 0.00665377f $X=2.16 $Y=0.335 $X2=0 $Y2=0
cc_141 N_B_c_123_n N_VGND_c_348_n 0.020191f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_142 N_B_c_120_n N_VGND_c_349_n 0.0191381f $X=0.62 $Y=0.335 $X2=0 $Y2=0
cc_143 N_B_c_119_n N_VGND_c_350_n 0.0235142f $X=1.995 $Y=0.335 $X2=0 $Y2=0
cc_144 N_B_c_123_n N_VGND_c_350_n 0.0414165f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_145 N_B_c_120_n N_VGND_c_352_n 0.0478156f $X=0.62 $Y=0.335 $X2=0 $Y2=0
cc_146 N_B_c_123_n N_VGND_c_352_n 0.0246682f $X=2.16 $Y=0.43 $X2=0 $Y2=0
cc_147 N_A_41_535#_M1001_g N_VPWR_c_251_n 0.0050558f $X=2.715 $Y=2.665 $X2=0
+ $Y2=0
cc_148 N_A_41_535#_c_193_n N_VPWR_c_254_n 0.00935935f $X=0.33 $Y=2.835 $X2=0
+ $Y2=0
cc_149 N_A_41_535#_M1001_g N_VPWR_c_255_n 0.00494486f $X=2.715 $Y=2.665 $X2=0
+ $Y2=0
cc_150 N_A_41_535#_M1004_s N_VPWR_c_249_n 0.00418801f $X=0.205 $Y=2.675 $X2=0
+ $Y2=0
cc_151 N_A_41_535#_M1001_g N_VPWR_c_249_n 0.00519032f $X=2.715 $Y=2.665 $X2=0
+ $Y2=0
cc_152 N_A_41_535#_c_193_n N_VPWR_c_249_n 0.00777327f $X=0.33 $Y=2.835 $X2=0
+ $Y2=0
cc_153 N_A_41_535#_M1001_g N_A_282_535#_c_295_n 5.17804e-19 $X=2.715 $Y=2.665
+ $X2=0 $Y2=0
cc_154 N_A_41_535#_M1003_g N_X_c_322_n 2.36833e-19 $X=2.725 $Y=0.99 $X2=0 $Y2=0
cc_155 N_A_41_535#_c_187_n N_X_c_316_n 0.014967f $X=2.685 $Y=1.645 $X2=0 $Y2=0
cc_156 N_A_41_535#_c_189_n N_X_c_316_n 2.64547e-19 $X=2.77 $Y=1.725 $X2=0 $Y2=0
cc_157 N_A_41_535#_M1003_g X 0.016663f $X=2.725 $Y=0.99 $X2=0 $Y2=0
cc_158 N_A_41_535#_c_187_n X 0.00459567f $X=2.685 $Y=1.645 $X2=0 $Y2=0
cc_159 N_A_41_535#_c_188_n X 0.0125585f $X=2.77 $Y=1.725 $X2=0 $Y2=0
cc_160 N_A_41_535#_c_189_n X 0.00453617f $X=2.77 $Y=1.725 $X2=0 $Y2=0
cc_161 N_A_41_535#_M1001_g X 0.00887595f $X=2.715 $Y=2.665 $X2=0 $Y2=0
cc_162 N_A_41_535#_M1003_g X 0.00571493f $X=2.725 $Y=0.99 $X2=0 $Y2=0
cc_163 N_A_41_535#_c_188_n X 0.0471564f $X=2.77 $Y=1.725 $X2=0 $Y2=0
cc_164 N_A_41_535#_c_189_n X 0.0163625f $X=2.77 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A_41_535#_M1001_g X 0.00659395f $X=2.715 $Y=2.665 $X2=0 $Y2=0
cc_166 N_A_41_535#_c_192_n X 0.002907f $X=2.77 $Y=2.23 $X2=0 $Y2=0
cc_167 N_A_41_535#_c_188_n X 0.00247029f $X=2.77 $Y=1.725 $X2=0 $Y2=0
cc_168 N_A_41_535#_c_185_n N_VGND_c_345_n 0.00829174f $X=0.435 $Y=1.645 $X2=0
+ $Y2=0
cc_169 N_A_41_535#_c_187_n N_VGND_c_346_n 0.0107963f $X=2.685 $Y=1.645 $X2=0
+ $Y2=0
cc_170 N_A_41_535#_M1003_g N_VGND_c_348_n 0.0100687f $X=2.725 $Y=0.99 $X2=0
+ $Y2=0
cc_171 N_A_41_535#_M1003_g N_VGND_c_350_n 0.00342259f $X=2.725 $Y=0.99 $X2=0
+ $Y2=0
cc_172 N_A_41_535#_M1003_g N_VGND_c_352_n 0.00428633f $X=2.725 $Y=0.99 $X2=0
+ $Y2=0
cc_173 A_124_535# N_VPWR_c_249_n 0.00350399f $X=0.62 $Y=2.675 $X2=3.12 $Y2=3.33
cc_174 N_VPWR_c_249_n N_A_282_535#_M1008_d 0.00442034f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_175 N_VPWR_c_252_n N_A_282_535#_c_292_n 0.00776392f $X=1.875 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_249_n N_A_282_535#_c_292_n 0.00690901f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_251_n N_A_282_535#_c_293_n 0.0148498f $X=1.98 $Y=2.95 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_252_n N_A_282_535#_c_293_n 0.00305343f $X=1.875 $Y=3.33 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_255_n N_A_282_535#_c_293_n 0.00379351f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_249_n N_A_282_535#_c_293_n 0.0125811f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_255_n N_A_282_535#_c_295_n 0.0053567f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_249_n N_A_282_535#_c_295_n 0.00767485f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_255_n X 0.0112481f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_249_n X 0.0143844f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_185 N_A_282_535#_c_295_n X 0.00377258f $X=2.46 $Y=2.52 $X2=0 $Y2=0
cc_186 X N_VGND_c_348_n 0.0274985f $X=3.035 $Y=1.21 $X2=0 $Y2=0
