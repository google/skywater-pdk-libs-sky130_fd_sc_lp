* File: sky130_fd_sc_lp__a21oi_1.pex.spice
* Created: Wed Sep  2 09:20:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21OI_1%A2 3 6 8 9 13 15
c25 8 0 2.16691e-19 $X=0.24 $Y=1.295
r26 13 16 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.377 $Y=1.46
+ $X2=0.377 $Y2=1.625
r27 13 15 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.377 $Y=1.46
+ $X2=0.377 $Y2=1.295
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.46 $X2=0.37 $Y2=1.46
r29 9 14 7.87503 $w=2.98e-07 $l=2.05e-07 $layer=LI1_cond $X=0.305 $Y=1.665
+ $X2=0.305 $Y2=1.46
r30 8 14 6.33844 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.305 $Y=1.295
+ $X2=0.305 $Y2=1.46
r31 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.625
r32 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.765
+ $X2=0.475 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_1%A1 3 7 9 10 11 12 19 31
c42 7 0 1.06063e-19 $X=0.975 $Y=2.465
c43 3 0 1.10627e-19 $X=0.865 $Y=0.765
r44 31 33 2.91866 $w=1.88e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.295 $X2=0.72
+ $Y2=1.345
r45 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.675
r46 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.345
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.51 $X2=0.925 $Y2=1.51
r48 12 20 4.52224 $w=3.93e-07 $l=1.55e-07 $layer=LI1_cond $X=0.822 $Y=1.665
+ $X2=0.822 $Y2=1.51
r49 11 20 4.31801 $w=3.93e-07 $l=1.48e-07 $layer=LI1_cond $X=0.822 $Y=1.362
+ $X2=0.822 $Y2=1.51
r50 11 33 3.61119 $w=3.93e-07 $l=1.7e-08 $layer=LI1_cond $X=0.822 $Y=1.362
+ $X2=0.822 $Y2=1.345
r51 11 31 1.05072 $w=1.88e-07 $l=1.8e-08 $layer=LI1_cond $X=0.72 $Y=1.277
+ $X2=0.72 $Y2=1.295
r52 10 11 20.5474 $w=1.88e-07 $l=3.52e-07 $layer=LI1_cond $X=0.72 $Y=0.925
+ $X2=0.72 $Y2=1.277
r53 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=0.555
+ $X2=0.72 $Y2=0.925
r54 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.975 $Y=2.465
+ $X2=0.975 $Y2=1.675
r55 3 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.865 $Y=0.765
+ $X2=0.865 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_1%B1 1 3 6 8 9 15
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.46 $X2=1.65 $Y2=1.46
r30 12 15 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.405 $Y=1.46
+ $X2=1.65 $Y2=1.46
r31 9 16 7.74593 $w=3.03e-07 $l=2.05e-07 $layer=LI1_cond $X=1.682 $Y=1.665
+ $X2=1.682 $Y2=1.46
r32 8 16 6.23453 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.682 $Y=1.295
+ $X2=1.682 $Y2=1.46
r33 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.625
+ $X2=1.405 $Y2=1.46
r34 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.405 $Y=1.625
+ $X2=1.405 $Y2=2.465
r35 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.295
+ $X2=1.405 $Y2=1.46
r36 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.405 $Y=1.295
+ $X2=1.405 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_1%A_27_367# 1 2 7 9 11 15 20
r28 13 20 1.49886 $w=2.95e-07 $l=9.31128e-08 $layer=LI1_cond $X=1.207 $Y=2.47
+ $X2=1.19 $Y2=2.385
r29 13 15 17.189 $w=2.93e-07 $l=4.4e-07 $layer=LI1_cond $X=1.207 $Y=2.47
+ $X2=1.207 $Y2=2.91
r30 12 18 2.69408 $w=5.4e-07 $l=1.48e-07 $layer=LI1_cond $X=0.39 $Y=2.2
+ $X2=0.242 $Y2=2.2
r31 11 20 11.6884 $w=5.4e-07 $l=5.24404e-07 $layer=LI1_cond $X=0.75 $Y=2.2
+ $X2=1.19 $Y2=2.385
r32 11 12 7.97386 $w=5.38e-07 $l=3.6e-07 $layer=LI1_cond $X=0.75 $Y=2.2 $X2=0.39
+ $Y2=2.2
r33 7 18 4.91488 $w=2.95e-07 $l=2.7e-07 $layer=LI1_cond $X=0.242 $Y=2.47
+ $X2=0.242 $Y2=2.2
r34 7 9 0.390659 $w=2.93e-07 $l=1e-08 $layer=LI1_cond $X=0.242 $Y=2.47 $X2=0.242
+ $Y2=2.48
r35 2 20 600 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.385
r36 2 15 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.91
r37 1 18 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.015
r38 1 9 300 $w=1.7e-07 $l=7.04734e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_1%VPWR 1 6 8 10 17 18 21
r29 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r31 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r32 15 17 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=1.68 $Y2=3.33
r33 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r36 10 12 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r37 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r40 4 6 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.765
r41 1 6 600 $w=1.7e-07 $l=1.01373e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.725 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_1%Y 1 2 8 9 10 11 12 13 27
r34 20 27 1.62879 $w=3.73e-07 $l=5.3e-08 $layer=LI1_cond $X=1.172 $Y=0.978
+ $X2=1.172 $Y2=0.925
r35 13 34 5.0187 $w=3.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.68 $Y=2.775
+ $X2=1.68 $Y2=2.91
r36 12 13 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.405
+ $X2=1.68 $Y2=2.775
r37 11 38 21.2576 $w=1.78e-07 $l=3.45e-07 $layer=LI1_cond $X=1.62 $Y=2.04
+ $X2=1.275 $Y2=2.04
r38 11 12 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.68 $Y=2.13
+ $X2=1.68 $Y2=2.405
r39 10 37 8.73886 $w=3.73e-07 $l=1.71e-07 $layer=LI1_cond $X=1.172 $Y=0.994
+ $X2=1.172 $Y2=1.165
r40 10 20 0.491709 $w=3.73e-07 $l=1.6e-08 $layer=LI1_cond $X=1.172 $Y=0.994
+ $X2=1.172 $Y2=0.978
r41 10 27 0.491709 $w=3.73e-07 $l=1.6e-08 $layer=LI1_cond $X=1.172 $Y=0.909
+ $X2=1.172 $Y2=0.925
r42 9 10 12.8766 $w=3.73e-07 $l=4.19e-07 $layer=LI1_cond $X=1.172 $Y=0.49
+ $X2=1.172 $Y2=0.909
r43 8 38 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.275 $Y=1.95 $X2=1.275
+ $Y2=2.04
r44 8 37 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.275 $Y=1.95
+ $X2=1.275 $Y2=1.165
r45 2 11 400 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2.115
r46 2 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2.91
r47 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.94
+ $Y=0.345 $X2=1.15 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_1%VGND 1 2 7 9 11 13 15 17 27
r26 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r27 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r29 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r30 18 23 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r31 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=1.2
+ $Y2=0
r32 17 26 4.28421 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.725
+ $Y2=0
r33 17 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.2
+ $Y2=0
r34 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r35 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r36 11 26 3.07584 $w=2.8e-07 $l=1.09087e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.725 $Y2=0
r37 11 13 16.6693 $w=2.78e-07 $l=4.05e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.49
r38 7 23 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r39 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.49
r40 2 13 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=1.48
+ $Y=0.345 $X2=1.645 $Y2=0.49
r41 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.49
.ends

