* NGSPICE file created from sky130_fd_sc_lp__a21o_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_792_49# A1 a_134_269# VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=4.704e+11p ps=4.48e+06u
M1001 VPWR a_134_269# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.7766e+12p pd=1.542e+07u as=7.056e+11p ps=6.16e+06u
M1002 X a_134_269# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=1.5204e+12p ps=1.202e+07u
M1003 a_792_49# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_134_269# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_529_367# B1 a_134_269# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3734e+12p pd=1.226e+07u as=3.528e+11p ps=3.08e+06u
M1006 VGND A2 a_792_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_529_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_134_269# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 a_134_269# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_134_269# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_134_269# B1 a_529_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_134_269# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_529_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_529_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_134_269# A1 a_792_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A2 a_529_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_134_269# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_134_269# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_134_269# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

