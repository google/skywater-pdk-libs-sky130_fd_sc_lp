* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_355_463# D a_380_50# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VPWR RESET_B a_380_50# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_937_333# a_865_255# a_1445_69# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_225_50# a_35_74# a_308_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_2408_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_1818_119# a_1445_69# a_1641_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR CLK a_865_255# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND CLK a_865_255# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_2408_367# a_1445_69# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_380_50# a_865_255# a_809_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_35_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_380_50# a_35_74# a_513_463# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1599_113# a_1641_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_2408_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR RESET_B a_809_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_512_81# SCD a_225_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_757_317# a_865_255# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_1641_21# a_1445_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 VGND a_809_463# a_937_333# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_380_50# a_757_317# a_809_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_1578_533# a_1641_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR RESET_B a_1641_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_809_463# a_757_317# a_991_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR SCE a_355_463# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_308_50# D a_380_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_757_317# a_865_255# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_35_74# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_809_463# a_865_255# a_895_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_895_463# a_937_333# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VPWR a_809_463# a_937_333# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X30 a_380_50# SCE a_512_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_225_50# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_2408_367# a_1445_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 a_1085_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND RESET_B a_1818_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1445_69# a_757_317# a_1578_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X36 a_991_119# a_937_333# a_1085_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_937_333# a_757_317# a_1445_69# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 a_1445_69# a_865_255# a_1599_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_513_463# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
