* File: sky130_fd_sc_lp__nor3b_2.pxi.spice
* Created: Wed Sep  2 10:09:41 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3B_2%C_N N_C_N_M1012_g N_C_N_M1001_g N_C_N_c_79_n
+ N_C_N_c_84_n C_N C_N N_C_N_c_80_n N_C_N_c_81_n PM_SKY130_FD_SC_LP__NOR3B_2%C_N
x_PM_SKY130_FD_SC_LP__NOR3B_2%A_27_131# N_A_27_131#_M1012_s N_A_27_131#_M1001_s
+ N_A_27_131#_M1006_g N_A_27_131#_c_112_n N_A_27_131#_M1000_g
+ N_A_27_131#_M1009_g N_A_27_131#_c_114_n N_A_27_131#_M1004_g
+ N_A_27_131#_c_115_n N_A_27_131#_c_116_n N_A_27_131#_c_117_n
+ N_A_27_131#_c_124_n N_A_27_131#_c_118_n N_A_27_131#_c_119_n
+ N_A_27_131#_c_125_n N_A_27_131#_c_126_n N_A_27_131#_c_120_n
+ N_A_27_131#_c_163_p N_A_27_131#_c_121_n PM_SKY130_FD_SC_LP__NOR3B_2%A_27_131#
x_PM_SKY130_FD_SC_LP__NOR3B_2%B N_B_M1002_g N_B_M1003_g N_B_M1010_g N_B_M1007_g
+ B N_B_c_201_n N_B_c_202_n PM_SKY130_FD_SC_LP__NOR3B_2%B
x_PM_SKY130_FD_SC_LP__NOR3B_2%A N_A_M1005_g N_A_M1011_g N_A_M1008_g N_A_M1013_g
+ A A A N_A_c_257_n PM_SKY130_FD_SC_LP__NOR3B_2%A
x_PM_SKY130_FD_SC_LP__NOR3B_2%VPWR N_VPWR_M1001_d N_VPWR_M1008_d N_VPWR_M1013_d
+ N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_299_n VPWR
+ N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n
+ N_VPWR_c_295_n PM_SKY130_FD_SC_LP__NOR3B_2%VPWR
x_PM_SKY130_FD_SC_LP__NOR3B_2%A_217_365# N_A_217_365#_M1006_d
+ N_A_217_365#_M1009_d N_A_217_365#_M1010_s N_A_217_365#_c_357_n
+ N_A_217_365#_c_353_n N_A_217_365#_c_364_n N_A_217_365#_c_354_n
+ N_A_217_365#_c_355_n N_A_217_365#_c_356_n N_A_217_365#_c_384_n
+ PM_SKY130_FD_SC_LP__NOR3B_2%A_217_365#
x_PM_SKY130_FD_SC_LP__NOR3B_2%Y N_Y_M1000_s N_Y_M1003_s N_Y_M1005_d N_Y_M1006_s
+ N_Y_c_395_n N_Y_c_446_p N_Y_c_396_n N_Y_c_447_p N_Y_c_397_n Y Y Y Y Y Y
+ N_Y_c_442_p Y Y PM_SKY130_FD_SC_LP__NOR3B_2%Y
x_PM_SKY130_FD_SC_LP__NOR3B_2%A_472_365# N_A_472_365#_M1002_d
+ N_A_472_365#_M1008_s N_A_472_365#_c_455_n N_A_472_365#_c_459_n
+ N_A_472_365#_c_454_n N_A_472_365#_c_468_n N_A_472_365#_c_474_n
+ PM_SKY130_FD_SC_LP__NOR3B_2%A_472_365#
x_PM_SKY130_FD_SC_LP__NOR3B_2%VGND N_VGND_M1012_d N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_M1011_s N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n
+ VGND N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n
+ N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n N_VGND_c_491_n N_VGND_c_492_n
+ PM_SKY130_FD_SC_LP__NOR3B_2%VGND
cc_1 VNB N_C_N_M1012_g 0.0439005f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.865
cc_2 VNB N_C_N_c_79_n 0.00344356f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_3 VNB N_C_N_c_80_n 0.0192606f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_4 VNB N_C_N_c_81_n 0.0110114f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_5 VNB N_A_27_131#_M1006_g 0.00771862f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_6 VNB N_A_27_131#_c_112_n 0.0207384f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_7 VNB N_A_27_131#_M1009_g 0.00623531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_131#_c_114_n 0.0171939f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_9 VNB N_A_27_131#_c_115_n 0.0583266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_131#_c_116_n 0.0479651f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.035
cc_11 VNB N_A_27_131#_c_117_n 0.0163722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_131#_c_118_n 0.010654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_131#_c_119_n 0.00964142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_131#_c_120_n 0.00249854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_131#_c_121_n 0.00497423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1003_g 0.0246385f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.75
cc_17 VNB N_B_M1007_g 0.0231529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB B 0.00282983f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_19 VNB N_B_c_201_n 0.046252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_c_202_n 0.00219549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_M1005_g 0.0236035f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.865
cc_22 VNB N_A_M1011_g 0.0342108f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.75
cc_23 VNB A 0.0404476f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_24 VNB N_A_c_257_n 0.066206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_295_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_395_n 0.00614791f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_27 VNB N_Y_c_396_n 0.00892285f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_28 VNB N_Y_c_397_n 0.00183474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB Y 0.00428826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 0.00161876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_480_n 0.0179461f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_VGND_c_481_n 0.00496801f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_33 VNB N_VGND_c_482_n 3.22989e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_483_n 0.0396624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_484_n 0.0178681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_485_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_486_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_487_n 0.0209183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_488_n 0.275151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_489_n 0.0410673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_490_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_491_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_492_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_C_N_M1001_g 0.0489863f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.75
cc_45 VPB N_C_N_c_79_n 0.0264006f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_46 VPB N_C_N_c_84_n 0.0197068f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_47 VPB N_C_N_c_81_n 0.0212656f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_48 VPB N_A_27_131#_M1006_g 0.0239697f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_49 VPB N_A_27_131#_M1009_g 0.0193798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_27_131#_c_124_n 0.0179496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_27_131#_c_125_n 0.014576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_27_131#_c_126_n 0.00969337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_131#_c_120_n 0.0141157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B_M1002_g 0.0190502f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.865
cc_55 VPB N_B_M1010_g 0.0240116f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_56 VPB B 0.00488962f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_57 VPB N_B_c_201_n 0.0141602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_M1008_g 0.0235869f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_59 VPB N_A_M1013_g 0.0235869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB A 0.0165391f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_61 VPB N_A_c_257_n 0.0200722f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_296_n 0.00980564f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_63 VPB N_VPWR_c_297_n 0.0156931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_298_n 0.0104993f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_65 VPB N_VPWR_c_299_n 0.0483636f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.615
cc_66 VPB N_VPWR_c_300_n 0.0169178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_301_n 0.065101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_302_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_303_n 0.00613202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_304_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_295_n 0.0721267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_217_365#_c_353_n 0.00205645f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_73 VPB N_A_217_365#_c_354_n 0.00301082f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_74 VPB N_A_217_365#_c_355_n 0.00285541f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.615
cc_75 VPB N_A_217_365#_c_356_n 0.00982738f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.035
cc_76 VPB Y 0.00168374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_472_365#_c_454_n 0.0248437f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_78 N_C_N_M1012_g N_A_27_131#_c_115_n 0.0172269f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_79 N_C_N_M1012_g N_A_27_131#_c_117_n 0.00169164f $X=0.475 $Y=0.865 $X2=0
+ $Y2=0
cc_80 N_C_N_M1001_g N_A_27_131#_c_124_n 0.00313661f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_81 N_C_N_M1012_g N_A_27_131#_c_118_n 0.0184816f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_82 N_C_N_c_80_n N_A_27_131#_c_118_n 3.11195e-19 $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_83 N_C_N_c_81_n N_A_27_131#_c_118_n 0.00881452f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_84 N_C_N_c_80_n N_A_27_131#_c_119_n 0.00103736f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_85 N_C_N_c_81_n N_A_27_131#_c_119_n 0.0234625f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_86 N_C_N_M1001_g N_A_27_131#_c_125_n 0.0171445f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_87 N_C_N_c_84_n N_A_27_131#_c_125_n 3.02199e-19 $X=0.385 $Y=2.12 $X2=0 $Y2=0
cc_88 N_C_N_c_81_n N_A_27_131#_c_125_n 0.00901834f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_89 N_C_N_c_84_n N_A_27_131#_c_126_n 0.0010133f $X=0.385 $Y=2.12 $X2=0 $Y2=0
cc_90 N_C_N_c_81_n N_A_27_131#_c_126_n 0.0241777f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_91 N_C_N_c_80_n N_A_27_131#_c_120_n 0.0194903f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_92 N_C_N_c_81_n N_A_27_131#_c_120_n 0.0316862f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_93 N_C_N_M1012_g N_A_27_131#_c_121_n 0.00485883f $X=0.475 $Y=0.865 $X2=0
+ $Y2=0
cc_94 N_C_N_c_81_n N_A_27_131#_c_121_n 0.00376433f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_95 N_C_N_M1001_g N_VPWR_c_296_n 0.0138465f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_96 N_C_N_M1001_g N_VPWR_c_300_n 0.00383152f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_97 N_C_N_M1001_g N_VPWR_c_295_n 0.00391732f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_98 N_C_N_M1001_g N_A_217_365#_c_357_n 6.08235e-19 $X=0.475 $Y=2.75 $X2=0
+ $Y2=0
cc_99 N_C_N_M1001_g N_A_217_365#_c_353_n 0.00438951f $X=0.475 $Y=2.75 $X2=0
+ $Y2=0
cc_100 N_C_N_M1012_g N_VGND_c_484_n 0.00333215f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_101 N_C_N_M1012_g N_VGND_c_488_n 0.00387424f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_102 N_C_N_M1012_g N_VGND_c_489_n 0.014794f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_103 N_A_27_131#_c_114_n N_B_M1003_g 0.0189504f $X=2.02 $Y=1.185 $X2=0 $Y2=0
cc_104 N_A_27_131#_M1009_g N_B_c_201_n 0.0261923f $X=1.855 $Y=2.455 $X2=0 $Y2=0
cc_105 N_A_27_131#_c_116_n N_B_c_201_n 0.00381172f $X=1.855 $Y=1.35 $X2=0 $Y2=0
cc_106 N_A_27_131#_M1009_g N_B_c_202_n 3.69966e-19 $X=1.855 $Y=2.455 $X2=0 $Y2=0
cc_107 N_A_27_131#_c_116_n N_B_c_202_n 9.12271e-19 $X=1.855 $Y=1.35 $X2=0 $Y2=0
cc_108 N_A_27_131#_M1006_g N_VPWR_c_296_n 0.00221845f $X=1.425 $Y=2.455 $X2=0
+ $Y2=0
cc_109 N_A_27_131#_c_125_n N_VPWR_c_296_n 0.0246736f $X=0.755 $Y=2.385 $X2=0
+ $Y2=0
cc_110 N_A_27_131#_c_124_n N_VPWR_c_300_n 0.00864257f $X=0.26 $Y=2.75 $X2=0
+ $Y2=0
cc_111 N_A_27_131#_M1006_g N_VPWR_c_301_n 0.00351226f $X=1.425 $Y=2.455 $X2=0
+ $Y2=0
cc_112 N_A_27_131#_M1009_g N_VPWR_c_301_n 0.00351226f $X=1.855 $Y=2.455 $X2=0
+ $Y2=0
cc_113 N_A_27_131#_M1006_g N_VPWR_c_295_n 0.00660267f $X=1.425 $Y=2.455 $X2=0
+ $Y2=0
cc_114 N_A_27_131#_M1009_g N_VPWR_c_295_n 0.00532831f $X=1.855 $Y=2.455 $X2=0
+ $Y2=0
cc_115 N_A_27_131#_c_124_n N_VPWR_c_295_n 0.00911154f $X=0.26 $Y=2.75 $X2=0
+ $Y2=0
cc_116 N_A_27_131#_c_125_n N_VPWR_c_295_n 0.00867721f $X=0.755 $Y=2.385 $X2=0
+ $Y2=0
cc_117 N_A_27_131#_M1006_g N_A_217_365#_c_353_n 0.00357735f $X=1.425 $Y=2.455
+ $X2=0 $Y2=0
cc_118 N_A_27_131#_c_115_n N_A_217_365#_c_353_n 0.00452483f $X=1.35 $Y=1.35
+ $X2=0 $Y2=0
cc_119 N_A_27_131#_c_125_n N_A_217_365#_c_353_n 0.0143312f $X=0.755 $Y=2.385
+ $X2=0 $Y2=0
cc_120 N_A_27_131#_c_120_n N_A_217_365#_c_353_n 0.0371818f $X=0.84 $Y=2.3 $X2=0
+ $Y2=0
cc_121 N_A_27_131#_c_163_p N_A_217_365#_c_353_n 0.0117884f $X=1.34 $Y=1.35 $X2=0
+ $Y2=0
cc_122 N_A_27_131#_M1006_g N_A_217_365#_c_364_n 0.0114688f $X=1.425 $Y=2.455
+ $X2=0 $Y2=0
cc_123 N_A_27_131#_M1009_g N_A_217_365#_c_364_n 0.0114222f $X=1.855 $Y=2.455
+ $X2=0 $Y2=0
cc_124 N_A_27_131#_M1009_g N_A_217_365#_c_354_n 8.28776e-19 $X=1.855 $Y=2.455
+ $X2=0 $Y2=0
cc_125 N_A_27_131#_c_116_n N_A_217_365#_c_354_n 0.0027782f $X=1.855 $Y=1.35
+ $X2=0 $Y2=0
cc_126 N_A_27_131#_c_114_n N_Y_c_395_n 0.0165519f $X=2.02 $Y=1.185 $X2=0 $Y2=0
cc_127 N_A_27_131#_c_112_n Y 0.00269561f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_128 N_A_27_131#_c_116_n Y 0.00285063f $X=1.855 $Y=1.35 $X2=0 $Y2=0
cc_129 N_A_27_131#_c_121_n Y 0.00194046f $X=0.84 $Y=1.312 $X2=0 $Y2=0
cc_130 N_A_27_131#_M1006_g Y 0.00385692f $X=1.425 $Y=2.455 $X2=0 $Y2=0
cc_131 N_A_27_131#_c_112_n Y 2.92164e-19 $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_132 N_A_27_131#_M1009_g Y 0.00823136f $X=1.855 $Y=2.455 $X2=0 $Y2=0
cc_133 N_A_27_131#_c_114_n Y 4.46199e-19 $X=2.02 $Y=1.185 $X2=0 $Y2=0
cc_134 N_A_27_131#_c_116_n Y 0.0233752f $X=1.855 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A_27_131#_c_120_n Y 0.00839295f $X=0.84 $Y=2.3 $X2=0 $Y2=0
cc_136 N_A_27_131#_c_163_p Y 0.0253322f $X=1.34 $Y=1.35 $X2=0 $Y2=0
cc_137 N_A_27_131#_c_121_n Y 6.33252e-19 $X=0.84 $Y=1.312 $X2=0 $Y2=0
cc_138 N_A_27_131#_M1006_g Y 0.00295174f $X=1.425 $Y=2.455 $X2=0 $Y2=0
cc_139 N_A_27_131#_M1009_g Y 0.00166729f $X=1.855 $Y=2.455 $X2=0 $Y2=0
cc_140 N_A_27_131#_c_116_n Y 2.04e-19 $X=1.855 $Y=1.35 $X2=0 $Y2=0
cc_141 N_A_27_131#_M1006_g Y 0.00804084f $X=1.425 $Y=2.455 $X2=0 $Y2=0
cc_142 N_A_27_131#_M1009_g Y 0.00764419f $X=1.855 $Y=2.455 $X2=0 $Y2=0
cc_143 N_A_27_131#_c_112_n N_VGND_c_480_n 0.00526846f $X=1.485 $Y=1.185 $X2=0
+ $Y2=0
cc_144 N_A_27_131#_c_114_n N_VGND_c_480_n 0.00585385f $X=2.02 $Y=1.185 $X2=0
+ $Y2=0
cc_145 N_A_27_131#_c_114_n N_VGND_c_481_n 0.0032219f $X=2.02 $Y=1.185 $X2=0
+ $Y2=0
cc_146 N_A_27_131#_c_117_n N_VGND_c_484_n 0.00423683f $X=0.26 $Y=0.865 $X2=0
+ $Y2=0
cc_147 N_A_27_131#_c_112_n N_VGND_c_488_n 0.00924047f $X=1.485 $Y=1.185 $X2=0
+ $Y2=0
cc_148 N_A_27_131#_c_114_n N_VGND_c_488_n 0.0110388f $X=2.02 $Y=1.185 $X2=0
+ $Y2=0
cc_149 N_A_27_131#_c_117_n N_VGND_c_488_n 0.00740463f $X=0.26 $Y=0.865 $X2=0
+ $Y2=0
cc_150 N_A_27_131#_c_112_n N_VGND_c_489_n 0.0133926f $X=1.485 $Y=1.185 $X2=0
+ $Y2=0
cc_151 N_A_27_131#_c_114_n N_VGND_c_489_n 0.00112166f $X=2.02 $Y=1.185 $X2=0
+ $Y2=0
cc_152 N_A_27_131#_c_115_n N_VGND_c_489_n 0.011717f $X=1.35 $Y=1.35 $X2=0 $Y2=0
cc_153 N_A_27_131#_c_118_n N_VGND_c_489_n 0.0161414f $X=0.755 $Y=1.195 $X2=0
+ $Y2=0
cc_154 N_A_27_131#_c_163_p N_VGND_c_489_n 0.0290303f $X=1.34 $Y=1.35 $X2=0 $Y2=0
cc_155 N_A_27_131#_c_121_n N_VGND_c_489_n 0.0156279f $X=0.84 $Y=1.312 $X2=0
+ $Y2=0
cc_156 N_B_M1007_g N_A_M1005_g 0.0246319f $X=2.97 $Y=0.655 $X2=0 $Y2=0
cc_157 B N_A_M1005_g 0.0026318f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_158 N_B_c_201_n N_A_M1005_g 0.0210437f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_159 B N_A_M1008_g 2.31424e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_160 B A 0.0367458f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_161 N_B_c_201_n A 2.98678e-19 $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_162 N_B_M1002_g N_VPWR_c_301_n 0.00351226f $X=2.285 $Y=2.455 $X2=0 $Y2=0
cc_163 N_B_M1010_g N_VPWR_c_301_n 0.00351226f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_164 N_B_M1002_g N_VPWR_c_295_n 0.00532831f $X=2.285 $Y=2.455 $X2=0 $Y2=0
cc_165 N_B_M1010_g N_VPWR_c_295_n 0.00660267f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_166 N_B_M1002_g N_A_217_365#_c_354_n 0.00116087f $X=2.285 $Y=2.455 $X2=0
+ $Y2=0
cc_167 N_B_M1002_g N_A_217_365#_c_355_n 0.0114688f $X=2.285 $Y=2.455 $X2=0 $Y2=0
cc_168 N_B_M1010_g N_A_217_365#_c_355_n 0.0114688f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_169 N_B_M1003_g N_Y_c_395_n 0.0148296f $X=2.54 $Y=0.655 $X2=0 $Y2=0
cc_170 N_B_c_201_n N_Y_c_395_n 0.00852745f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_171 N_B_c_202_n N_Y_c_395_n 0.0129835f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_172 N_B_M1007_g N_Y_c_396_n 0.013286f $X=2.97 $Y=0.655 $X2=0 $Y2=0
cc_173 N_B_c_201_n N_Y_c_396_n 0.00145734f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_174 N_B_c_202_n N_Y_c_396_n 0.0277185f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_175 N_B_c_201_n N_Y_c_397_n 0.00266482f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_176 N_B_c_202_n N_Y_c_397_n 0.0193992f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_177 N_B_M1003_g Y 5.37516e-19 $X=2.54 $Y=0.655 $X2=0 $Y2=0
cc_178 N_B_c_201_n Y 9.48256e-19 $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_179 N_B_c_202_n Y 0.00843263f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_180 N_B_M1002_g Y 7.74836e-19 $X=2.285 $Y=2.455 $X2=0 $Y2=0
cc_181 N_B_M1002_g N_A_472_365#_c_455_n 0.00362131f $X=2.285 $Y=2.455 $X2=0
+ $Y2=0
cc_182 N_B_M1010_g N_A_472_365#_c_455_n 0.00400136f $X=2.715 $Y=2.455 $X2=0
+ $Y2=0
cc_183 N_B_c_201_n N_A_472_365#_c_455_n 0.00264974f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_184 N_B_c_202_n N_A_472_365#_c_455_n 0.0152151f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_185 N_B_M1002_g N_A_472_365#_c_459_n 0.0068358f $X=2.285 $Y=2.455 $X2=0 $Y2=0
cc_186 N_B_M1010_g N_A_472_365#_c_459_n 0.0127128f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_187 N_B_M1010_g N_A_472_365#_c_454_n 0.0136016f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_188 B N_A_472_365#_c_454_n 0.0284067f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_189 N_B_c_201_n N_A_472_365#_c_454_n 0.00292343f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_190 N_B_c_202_n N_A_472_365#_c_454_n 0.00865492f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_191 N_B_M1003_g N_VGND_c_481_n 0.00174472f $X=2.54 $Y=0.655 $X2=0 $Y2=0
cc_192 N_B_M1003_g N_VGND_c_482_n 6.27404e-19 $X=2.54 $Y=0.655 $X2=0 $Y2=0
cc_193 N_B_M1007_g N_VGND_c_482_n 0.010132f $X=2.97 $Y=0.655 $X2=0 $Y2=0
cc_194 N_B_M1003_g N_VGND_c_485_n 0.00585385f $X=2.54 $Y=0.655 $X2=0 $Y2=0
cc_195 N_B_M1007_g N_VGND_c_485_n 0.00486043f $X=2.97 $Y=0.655 $X2=0 $Y2=0
cc_196 N_B_M1003_g N_VGND_c_488_n 0.0107631f $X=2.54 $Y=0.655 $X2=0 $Y2=0
cc_197 N_B_M1007_g N_VGND_c_488_n 0.00824727f $X=2.97 $Y=0.655 $X2=0 $Y2=0
cc_198 N_A_M1008_g N_VPWR_c_297_n 0.0175702f $X=3.89 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A_M1013_g N_VPWR_c_297_n 6.80491e-19 $X=4.32 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A_M1008_g N_VPWR_c_299_n 7.4416e-19 $X=3.89 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A_M1013_g N_VPWR_c_299_n 0.0206425f $X=4.32 $Y=2.465 $X2=0 $Y2=0
cc_202 A N_VPWR_c_299_n 0.0262188f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_M1008_g N_VPWR_c_302_n 0.00486043f $X=3.89 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A_M1013_g N_VPWR_c_302_n 0.00486043f $X=4.32 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A_M1008_g N_VPWR_c_295_n 0.00824727f $X=3.89 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_M1013_g N_VPWR_c_295_n 0.00824727f $X=4.32 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_M1005_g N_Y_c_396_n 0.0148035f $X=3.4 $Y=0.655 $X2=0 $Y2=0
cc_208 N_A_M1011_g N_Y_c_396_n 0.00253213f $X=3.83 $Y=0.655 $X2=0 $Y2=0
cc_209 A N_Y_c_396_n 0.0308272f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A_c_257_n N_Y_c_396_n 7.70942e-19 $X=4.32 $Y=1.51 $X2=0 $Y2=0
cc_211 N_A_M1008_g N_A_472_365#_c_454_n 0.0143f $X=3.89 $Y=2.465 $X2=0 $Y2=0
cc_212 A N_A_472_365#_c_454_n 0.0451172f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A_c_257_n N_A_472_365#_c_454_n 0.00465161f $X=4.32 $Y=1.51 $X2=0 $Y2=0
cc_214 A N_A_472_365#_c_468_n 0.0152412f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_215 N_A_c_257_n N_A_472_365#_c_468_n 6.52992e-19 $X=4.32 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A_M1005_g N_VGND_c_482_n 0.010132f $X=3.4 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A_M1011_g N_VGND_c_482_n 6.27404e-19 $X=3.83 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A_M1011_g N_VGND_c_483_n 0.00702716f $X=3.83 $Y=0.655 $X2=0 $Y2=0
cc_219 A N_VGND_c_483_n 0.0203314f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_220 N_A_c_257_n N_VGND_c_483_n 0.00212584f $X=4.32 $Y=1.51 $X2=0 $Y2=0
cc_221 N_A_M1005_g N_VGND_c_486_n 0.00486043f $X=3.4 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A_M1011_g N_VGND_c_486_n 0.00585385f $X=3.83 $Y=0.655 $X2=0 $Y2=0
cc_223 N_A_M1005_g N_VGND_c_488_n 0.00824727f $X=3.4 $Y=0.655 $X2=0 $Y2=0
cc_224 N_A_M1011_g N_VGND_c_488_n 0.0118358f $X=3.83 $Y=0.655 $X2=0 $Y2=0
cc_225 N_VPWR_c_295_n N_A_217_365#_M1006_d 0.00247091f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_226 N_VPWR_c_295_n N_A_217_365#_M1009_d 0.00223565f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_295_n N_A_217_365#_M1010_s 0.00212303f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_296_n N_A_217_365#_c_357_n 0.0114889f $X=0.69 $Y=2.765 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_301_n N_A_217_365#_c_357_n 0.0143128f $X=3.51 $Y=3.33 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_295_n N_A_217_365#_c_357_n 0.00815375f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_296_n N_A_217_365#_c_353_n 0.0163475f $X=0.69 $Y=2.765 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_301_n N_A_217_365#_c_364_n 0.0361172f $X=3.51 $Y=3.33 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_295_n N_A_217_365#_c_364_n 0.023676f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_234 N_VPWR_c_297_n N_A_217_365#_c_355_n 0.0080981f $X=3.675 $Y=2.365 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_301_n N_A_217_365#_c_355_n 0.0540354f $X=3.51 $Y=3.33 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_295_n N_A_217_365#_c_355_n 0.0337842f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_297_n N_A_217_365#_c_356_n 0.0284588f $X=3.675 $Y=2.365 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_301_n N_A_217_365#_c_384_n 0.0125234f $X=3.51 $Y=3.33 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_295_n N_A_217_365#_c_384_n 0.0073762f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_295_n N_Y_M1006_s 0.00225186f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_c_295_n N_A_472_365#_M1002_d 0.00225186f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_242 N_VPWR_c_295_n N_A_472_365#_M1008_s 0.00571434f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_VPWR_M1008_d N_A_472_365#_c_454_n 0.00479121f $X=3.55 $Y=1.835 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_297_n N_A_472_365#_c_454_n 0.0220026f $X=3.675 $Y=2.365 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_302_n N_A_472_365#_c_474_n 0.0120977f $X=4.37 $Y=3.33 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_295_n N_A_472_365#_c_474_n 0.00691495f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_247 N_A_217_365#_c_364_n N_Y_M1006_s 0.00332344f $X=1.975 $Y=2.99 $X2=0 $Y2=0
cc_248 N_A_217_365#_c_354_n N_Y_c_395_n 0.00585765f $X=2.07 $Y=1.97 $X2=0 $Y2=0
cc_249 N_A_217_365#_c_353_n Y 0.00152483f $X=1.21 $Y=1.97 $X2=0 $Y2=0
cc_250 N_A_217_365#_c_354_n Y 0.0354498f $X=2.07 $Y=1.97 $X2=0 $Y2=0
cc_251 N_A_217_365#_c_364_n Y 0.0159805f $X=1.975 $Y=2.99 $X2=0 $Y2=0
cc_252 N_A_217_365#_c_355_n N_A_472_365#_M1002_d 0.00332344f $X=2.835 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_253 N_A_217_365#_c_355_n N_A_472_365#_c_459_n 0.0159805f $X=2.835 $Y=2.99
+ $X2=0 $Y2=0
cc_254 N_A_217_365#_M1010_s N_A_472_365#_c_454_n 0.0048182f $X=2.79 $Y=1.825
+ $X2=0 $Y2=0
cc_255 N_A_217_365#_c_356_n N_A_472_365#_c_454_n 0.0202165f $X=2.93 $Y=2.425
+ $X2=0 $Y2=0
cc_256 N_Y_c_395_n N_VGND_M1004_d 0.0027754f $X=2.62 $Y=1.075 $X2=0 $Y2=0
cc_257 N_Y_c_396_n N_VGND_M1007_d 0.00176461f $X=3.52 $Y=1.08 $X2=0 $Y2=0
cc_258 N_Y_c_442_p N_VGND_c_480_n 0.0210771f $X=1.76 $Y=0.42 $X2=0 $Y2=0
cc_259 N_Y_c_395_n N_VGND_c_481_n 0.0209082f $X=2.62 $Y=1.075 $X2=0 $Y2=0
cc_260 N_Y_c_396_n N_VGND_c_482_n 0.0170777f $X=3.52 $Y=1.08 $X2=0 $Y2=0
cc_261 N_Y_c_396_n N_VGND_c_483_n 0.00166417f $X=3.52 $Y=1.08 $X2=0 $Y2=0
cc_262 N_Y_c_446_p N_VGND_c_485_n 0.0138717f $X=2.755 $Y=0.42 $X2=0 $Y2=0
cc_263 N_Y_c_447_p N_VGND_c_486_n 0.0138717f $X=3.615 $Y=0.42 $X2=0 $Y2=0
cc_264 N_Y_M1000_s N_VGND_c_488_n 0.00504451f $X=1.56 $Y=0.235 $X2=0 $Y2=0
cc_265 N_Y_M1003_s N_VGND_c_488_n 0.00397496f $X=2.615 $Y=0.235 $X2=0 $Y2=0
cc_266 N_Y_M1005_d N_VGND_c_488_n 0.00397496f $X=3.475 $Y=0.235 $X2=0 $Y2=0
cc_267 N_Y_c_446_p N_VGND_c_488_n 0.00886411f $X=2.755 $Y=0.42 $X2=0 $Y2=0
cc_268 N_Y_c_447_p N_VGND_c_488_n 0.00886411f $X=3.615 $Y=0.42 $X2=0 $Y2=0
cc_269 N_Y_c_442_p N_VGND_c_488_n 0.0127519f $X=1.76 $Y=0.42 $X2=0 $Y2=0
