# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sdfstp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.950000 2.255000 2.225000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.390000 0.255000 14.590000 0.965000 ;
        RECT 14.390000 0.965000 15.275000 1.135000 ;
        RECT 14.390000 1.825000 15.275000 1.995000 ;
        RECT 14.390000 1.995000 14.590000 3.075000 ;
        RECT 14.555000 1.135000 15.275000 1.825000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.150000 0.550000 1.780000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435000 0.265000 3.765000 1.380000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.315000 0.265000 11.040000 0.500000 ;
        RECT  8.315000 0.500000  9.925000 0.640000 ;
        RECT 10.870000 0.500000 11.040000 1.585000 ;
        RECT 10.870000 1.585000 12.090000 1.765000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.305000 0.780000 4.685000 1.825000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.245000 15.360000 3.415000 ;
      RECT  0.155000  2.395000  2.245000 2.645000 ;
      RECT  0.155000  2.645000  0.415000 3.065000 ;
      RECT  0.405000  0.085000  0.735000 0.980000 ;
      RECT  0.585000  2.815000  0.915000 3.245000 ;
      RECT  1.195000  0.650000  1.525000 1.150000 ;
      RECT  1.195000  1.150000  2.595000 1.405000 ;
      RECT  1.430000  2.815000  2.595000 3.075000 ;
      RECT  1.985000  0.085000  2.620000 0.980000 ;
      RECT  2.425000  1.405000  2.595000 1.950000 ;
      RECT  2.425000  1.950000  3.365000 2.120000 ;
      RECT  2.425000  2.120000  2.595000 2.815000 ;
      RECT  2.765000  2.300000  3.025000 3.245000 ;
      RECT  2.790000  0.650000  3.085000 1.550000 ;
      RECT  2.790000  1.550000  3.785000 1.780000 ;
      RECT  3.195000  2.120000  3.365000 2.800000 ;
      RECT  3.195000  2.800000  4.320000 2.970000 ;
      RECT  3.535000  1.780000  3.785000 2.630000 ;
      RECT  3.965000  0.280000  4.230000 0.610000 ;
      RECT  3.965000  0.610000  4.135000 1.995000 ;
      RECT  3.965000  1.995000  5.135000 2.185000 ;
      RECT  3.965000  2.185000  4.305000 2.325000 ;
      RECT  4.150000  2.495000  5.740000 2.525000 ;
      RECT  4.150000  2.525000  4.830000 2.665000 ;
      RECT  4.150000  2.665000  4.320000 2.800000 ;
      RECT  4.400000  0.085000  4.655000 0.610000 ;
      RECT  4.500000  2.835000  4.830000 3.245000 ;
      RECT  4.660000  2.355000  5.740000 2.495000 ;
      RECT  4.825000  0.255000  6.070000 0.425000 ;
      RECT  4.825000  0.425000  5.120000 0.610000 ;
      RECT  4.855000  1.245000  5.135000 1.995000 ;
      RECT  5.000000  2.705000  6.790000 3.035000 ;
      RECT  5.380000  0.595000  5.710000 2.185000 ;
      RECT  5.380000  2.185000  5.740000 2.355000 ;
      RECT  5.880000  0.425000  6.070000 1.375000 ;
      RECT  5.880000  1.375000  6.090000 1.705000 ;
      RECT  5.910000  1.705000  6.090000 2.705000 ;
      RECT  6.240000  0.325000  6.430000 0.715000 ;
      RECT  6.260000  0.715000  6.430000 1.225000 ;
      RECT  6.260000  1.225000  9.085000 1.415000 ;
      RECT  6.260000  1.415000  6.450000 2.385000 ;
      RECT  6.620000  1.935000  7.650000 2.105000 ;
      RECT  6.620000  2.105000  6.790000 2.705000 ;
      RECT  6.825000  0.725000  7.795000 1.055000 ;
      RECT  6.845000  1.585000  8.010000 1.765000 ;
      RECT  6.950000  0.085000  7.280000 0.555000 ;
      RECT  6.980000  2.275000  7.310000 3.245000 ;
      RECT  7.480000  2.105000  7.650000 2.565000 ;
      RECT  7.480000  2.565000  8.350000 2.735000 ;
      RECT  7.820000  1.765000  8.010000 2.385000 ;
      RECT  7.965000  0.085000  8.135000 0.810000 ;
      RECT  7.965000  0.810000  9.540000 1.010000 ;
      RECT  8.180000  1.735000  9.910000 1.905000 ;
      RECT  8.180000  1.905000  8.350000 2.565000 ;
      RECT  8.520000  2.075000  8.745000 3.245000 ;
      RECT  8.915000  2.075000  9.210000 2.275000 ;
      RECT  8.915000  2.275000 10.840000 2.445000 ;
      RECT  8.915000  2.445000  9.210000 2.755000 ;
      RECT  9.420000  2.615000  9.750000 2.795000 ;
      RECT  9.420000  2.795000 11.360000 2.965000 ;
      RECT  9.610000  1.905000  9.910000 2.095000 ;
      RECT 10.080000  1.915000 10.700000 1.935000 ;
      RECT 10.080000  1.935000 12.760000 2.105000 ;
      RECT 10.095000  0.670000 10.700000 1.915000 ;
      RECT 10.510000  2.445000 10.840000 2.615000 ;
      RECT 11.060000  2.275000 11.360000 2.795000 ;
      RECT 11.220000  1.235000 13.200000 1.415000 ;
      RECT 11.530000  2.275000 11.785000 3.245000 ;
      RECT 11.885000  0.085000 12.215000 0.995000 ;
      RECT 11.955000  2.105000 12.760000 2.255000 ;
      RECT 11.955000  2.255000 12.250000 2.550000 ;
      RECT 12.425000  0.665000 12.755000 1.235000 ;
      RECT 12.440000  2.460000 12.760000 3.245000 ;
      RECT 12.500000  1.585000 12.760000 1.935000 ;
      RECT 12.930000  1.415000 13.200000 2.790000 ;
      RECT 13.390000  0.700000 13.670000 1.315000 ;
      RECT 13.390000  1.315000 14.335000 1.645000 ;
      RECT 13.390000  1.645000 13.685000 2.485000 ;
      RECT 13.840000  0.085000 14.170000 1.095000 ;
      RECT 13.855000  1.825000 14.220000 3.245000 ;
      RECT 14.760000  0.085000 15.090000 0.795000 ;
      RECT 14.760000  2.165000 15.090000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfstp_2
