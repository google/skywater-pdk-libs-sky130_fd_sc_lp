* File: sky130_fd_sc_lp__invlp_1.pxi.spice
* Created: Fri Aug 28 10:39:45 2020
* 
x_PM_SKY130_FD_SC_LP__INVLP_1%A N_A_c_23_n N_A_M1003_g N_A_M1000_g N_A_c_25_n
+ N_A_c_26_n N_A_M1001_g N_A_M1002_g N_A_c_28_n N_A_c_29_n N_A_c_30_n A
+ PM_SKY130_FD_SC_LP__INVLP_1%A
x_PM_SKY130_FD_SC_LP__INVLP_1%VPWR N_VPWR_M1000_s N_VPWR_c_57_n N_VPWR_c_58_n
+ VPWR N_VPWR_c_59_n N_VPWR_c_56_n PM_SKY130_FD_SC_LP__INVLP_1%VPWR
x_PM_SKY130_FD_SC_LP__INVLP_1%Y N_Y_M1001_d N_Y_M1002_d Y Y Y Y Y Y Y N_Y_c_75_n
+ PM_SKY130_FD_SC_LP__INVLP_1%Y
x_PM_SKY130_FD_SC_LP__INVLP_1%VGND N_VGND_M1003_s N_VGND_c_91_n N_VGND_c_92_n
+ VGND N_VGND_c_93_n N_VGND_c_94_n PM_SKY130_FD_SC_LP__INVLP_1%VGND
cc_1 VNB N_A_c_23_n 0.0206088f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.185
cc_2 VNB N_A_M1000_g 0.010756f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_3 VNB N_A_c_25_n 0.00779456f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.26
cc_4 VNB N_A_c_26_n 0.0195654f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.185
cc_5 VNB N_A_M1002_g 0.018812f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_6 VNB N_A_c_28_n 0.0494845f $X=-0.19 $Y=-0.245 $X2=0.47 $Y2=1.35
cc_7 VNB N_A_c_29_n 0.00974826f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.35
cc_8 VNB N_A_c_30_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.26
cc_9 VNB A 0.00998322f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_VPWR_c_56_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_11 VNB N_Y_c_75_n 0.0555506f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.35
cc_12 VNB N_VGND_c_91_n 0.0125985f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.515
cc_13 VNB N_VGND_c_92_n 0.0321429f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_14 VNB N_VGND_c_93_n 0.0279551f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_15 VNB N_VGND_c_94_n 0.111965f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.335
cc_16 VPB N_A_M1000_g 0.0255645f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_17 VPB N_A_M1002_g 0.0234886f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_18 VPB N_VPWR_c_57_n 0.0135296f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.515
cc_19 VPB N_VPWR_c_58_n 0.0539213f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_20 VPB N_VPWR_c_59_n 0.0270004f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_21 VPB N_VPWR_c_56_n 0.049042f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_22 VPB N_Y_c_75_n 0.0547566f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.35
cc_23 N_A_M1000_g N_VPWR_c_58_n 0.0317724f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_24 N_A_M1002_g N_VPWR_c_58_n 0.00466134f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_25 N_A_c_28_n N_VPWR_c_58_n 0.00376879f $X=0.47 $Y=1.35 $X2=0 $Y2=0
cc_26 A N_VPWR_c_58_n 0.0143153f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_27 N_A_M1000_g N_VPWR_c_59_n 0.00486043f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_28 N_A_M1002_g N_VPWR_c_59_n 0.0054895f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_29 N_A_M1000_g N_VPWR_c_56_n 0.00814425f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_30 N_A_M1002_g N_VPWR_c_56_n 0.0107696f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_31 N_A_c_23_n N_Y_c_75_n 0.00299127f $X=0.545 $Y=1.185 $X2=0 $Y2=0
cc_32 N_A_c_26_n N_Y_c_75_n 0.0203563f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_33 N_A_M1002_g N_Y_c_75_n 0.0416428f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_34 N_A_c_29_n N_Y_c_75_n 0.0055523f $X=0.56 $Y=1.35 $X2=0 $Y2=0
cc_35 N_A_c_30_n N_Y_c_75_n 0.00731937f $X=0.935 $Y=1.26 $X2=0 $Y2=0
cc_36 A N_Y_c_75_n 0.00989672f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_37 N_A_c_23_n N_VGND_c_92_n 0.021395f $X=0.545 $Y=1.185 $X2=0 $Y2=0
cc_38 N_A_c_26_n N_VGND_c_92_n 0.00332397f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_39 N_A_c_28_n N_VGND_c_92_n 0.00212401f $X=0.47 $Y=1.35 $X2=0 $Y2=0
cc_40 A N_VGND_c_92_n 0.0232978f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_41 N_A_c_23_n N_VGND_c_93_n 0.00486043f $X=0.545 $Y=1.185 $X2=0 $Y2=0
cc_42 N_A_c_26_n N_VGND_c_93_n 0.0054895f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_43 N_A_c_23_n N_VGND_c_94_n 0.00823808f $X=0.545 $Y=1.185 $X2=0 $Y2=0
cc_44 N_A_c_26_n N_VGND_c_94_n 0.0108635f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_45 N_VPWR_c_56_n A_130_367# 0.00899413f $X=1.2 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_46 N_VPWR_c_56_n N_Y_M1002_d 0.00231914f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_47 N_VPWR_c_58_n N_Y_c_75_n 0.0421563f $X=0.36 $Y=1.98 $X2=0 $Y2=0
cc_48 N_VPWR_c_59_n N_Y_c_75_n 0.0210192f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_49 N_VPWR_c_56_n N_Y_c_75_n 0.0125689f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_50 N_Y_c_75_n N_VGND_c_92_n 0.0239189f $X=1.15 $Y=0.42 $X2=0 $Y2=0
cc_51 N_Y_c_75_n N_VGND_c_93_n 0.0210192f $X=1.15 $Y=0.42 $X2=0 $Y2=0
cc_52 N_Y_M1001_d N_VGND_c_94_n 0.00231914f $X=1.01 $Y=0.235 $X2=0 $Y2=0
cc_53 N_Y_c_75_n N_VGND_c_94_n 0.0125689f $X=1.15 $Y=0.42 $X2=0 $Y2=0
cc_54 N_VGND_c_94_n A_124_47# 0.010279f $X=1.2 $Y=0 $X2=-0.19 $Y2=-0.245
