# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__o22ai_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o22ai_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.035000 2.845000 1.705000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.035000 2.275000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.450000 0.845000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.450000 1.415000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.437600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.165000 1.100000 1.170000 1.270000 ;
        RECT 0.165000 1.270000 0.335000 1.960000 ;
        RECT 0.165000 1.960000 1.315000 2.130000 ;
        RECT 0.840000 0.615000 1.170000 1.100000 ;
        RECT 1.085000 2.130000 1.315000 2.235000 ;
        RECT 1.085000 2.235000 1.640000 3.065000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 3.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.290000  2.310000 0.620000 3.245000 ;
      RECT 0.330000  0.265000 1.765000 0.435000 ;
      RECT 0.330000  0.435000 0.660000 0.920000 ;
      RECT 1.350000  0.435000 1.765000 0.945000 ;
      RECT 1.595000  0.945000 1.765000 1.885000 ;
      RECT 1.595000  1.885000 3.195000 2.055000 ;
      RECT 1.945000  0.085000 2.275000 0.855000 ;
      RECT 2.640000  0.485000 3.195000 0.855000 ;
      RECT 2.740000  2.235000 3.070000 3.245000 ;
      RECT 3.025000  0.855000 3.195000 1.885000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__o22ai_lp
END LIBRARY
