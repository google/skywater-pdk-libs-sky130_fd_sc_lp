* File: sky130_fd_sc_lp__and3_0.pxi.spice
* Created: Fri Aug 28 10:05:43 2020
* 
x_PM_SKY130_FD_SC_LP__AND3_0%A N_A_c_66_n N_A_M1005_g N_A_M1007_g N_A_c_67_n
+ N_A_c_68_n N_A_c_73_n A A A N_A_c_70_n N_A_c_71_n PM_SKY130_FD_SC_LP__AND3_0%A
x_PM_SKY130_FD_SC_LP__AND3_0%B N_B_M1003_g N_B_M1002_g N_B_c_109_n N_B_c_114_n B
+ B N_B_c_111_n PM_SKY130_FD_SC_LP__AND3_0%B
x_PM_SKY130_FD_SC_LP__AND3_0%C N_C_c_157_n N_C_M1001_g N_C_M1000_g N_C_c_158_n
+ N_C_c_159_n N_C_c_165_n N_C_c_166_n N_C_c_167_n C C C N_C_c_161_n N_C_c_162_n
+ C PM_SKY130_FD_SC_LP__AND3_0%C
x_PM_SKY130_FD_SC_LP__AND3_0%A_68_65# N_A_68_65#_M1005_s N_A_68_65#_M1007_s
+ N_A_68_65#_M1002_d N_A_68_65#_c_219_n N_A_68_65#_M1004_g N_A_68_65#_M1006_g
+ N_A_68_65#_c_222_n N_A_68_65#_c_223_n N_A_68_65#_c_233_n N_A_68_65#_c_224_n
+ N_A_68_65#_c_225_n N_A_68_65#_c_234_n N_A_68_65#_c_226_n N_A_68_65#_c_227_n
+ N_A_68_65#_c_228_n N_A_68_65#_c_229_n N_A_68_65#_c_230_n N_A_68_65#_c_235_n
+ N_A_68_65#_c_292_p N_A_68_65#_c_236_n PM_SKY130_FD_SC_LP__AND3_0%A_68_65#
x_PM_SKY130_FD_SC_LP__AND3_0%VPWR N_VPWR_M1007_d N_VPWR_M1000_d N_VPWR_c_320_n
+ N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n VPWR
+ N_VPWR_c_325_n N_VPWR_c_319_n N_VPWR_c_327_n PM_SKY130_FD_SC_LP__AND3_0%VPWR
x_PM_SKY130_FD_SC_LP__AND3_0%X N_X_M1006_d N_X_M1004_d X X X X X X X X
+ PM_SKY130_FD_SC_LP__AND3_0%X
x_PM_SKY130_FD_SC_LP__AND3_0%VGND N_VGND_M1001_d VGND N_VGND_c_371_n
+ N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n PM_SKY130_FD_SC_LP__AND3_0%VGND
cc_1 VNB N_A_c_66_n 0.0221631f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.345
cc_2 VNB N_A_c_67_n 0.0185117f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.525
cc_3 VNB N_A_c_68_n 0.0074722f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=2.155
cc_4 VNB A 0.00896295f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_5 VNB N_A_c_70_n 0.0187808f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.02
cc_6 VNB N_A_c_71_n 0.0206354f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.855
cc_7 VNB N_B_M1003_g 0.0346546f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.525
cc_8 VNB N_B_c_109_n 0.0150682f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.525
cc_9 VNB B 0.00496147f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=2.305
cc_10 VNB N_B_c_111_n 0.015327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_c_157_n 0.0206309f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.035
cc_12 VNB N_C_c_158_n 0.026119f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.305
cc_13 VNB N_C_c_159_n 0.0173601f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.525
cc_14 VNB C 0.00499652f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.02
cc_15 VNB N_C_c_161_n 0.0170606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C_c_162_n 0.0128015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_68_65#_c_219_n 0.0239081f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.525
cc_18 VNB N_A_68_65#_M1004_g 0.00173748f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_19 VNB N_A_68_65#_M1006_g 0.0308944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_68_65#_c_222_n 0.0229154f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.02
cc_21 VNB N_A_68_65#_c_223_n 0.0462903f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.02
cc_22 VNB N_A_68_65#_c_224_n 7.92559e-19 $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.02
cc_23 VNB N_A_68_65#_c_225_n 0.0156131f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.295
cc_24 VNB N_A_68_65#_c_226_n 7.73304e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_68_65#_c_227_n 0.0179995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_68_65#_c_228_n 7.30704e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_68_65#_c_229_n 0.0066793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_68_65#_c_230_n 0.0223693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_319_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB X 0.0632329f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.535
cc_31 VNB N_VGND_c_371_n 0.0162788f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB N_VGND_c_372_n 0.181292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_373_n 0.0404941f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.02
cc_34 VNB N_VGND_c_374_n 0.0227126f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.295
cc_35 VPB N_A_c_68_n 0.030179f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=2.155
cc_36 VPB N_A_c_73_n 0.0319865f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=2.305
cc_37 VPB A 0.00475245f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_38 VPB N_B_M1002_g 0.0365396f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.535
cc_39 VPB N_B_c_109_n 0.00580495f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.525
cc_40 VPB N_B_c_114_n 0.0152609f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=2.155
cc_41 VPB B 0.00328376f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=2.305
cc_42 VPB N_C_M1000_g 0.0213262f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.535
cc_43 VPB N_C_c_159_n 0.00314667f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.525
cc_44 VPB N_C_c_165_n 0.0137663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_C_c_166_n 0.0126119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_C_c_167_n 0.0179855f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.02
cc_47 VPB C 5.38506e-19 $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.02
cc_48 VPB C 0.00830162f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.855
cc_49 VPB N_A_68_65#_M1004_g 0.0645753f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_50 VPB N_A_68_65#_c_223_n 0.0216517f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.02
cc_51 VPB N_A_68_65#_c_233_n 0.0283302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_68_65#_c_234_n 0.0139824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_68_65#_c_235_n 0.0148087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_68_65#_c_236_n 0.00257275f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_320_n 0.0156478f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.625
cc_56 VPB N_VPWR_c_321_n 0.0175917f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.525
cc_57 VPB N_VPWR_c_322_n 0.0295271f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_58 VPB N_VPWR_c_323_n 0.0248753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_324_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_325_n 0.018524f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.295
cc_61 VPB N_VPWR_c_319_n 0.0672018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_327_n 0.0116111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB X 0.04124f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.535
cc_64 VPB X 0.0229888f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=2.305
cc_65 VPB X 0.0116595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 A N_B_M1003_g 0.00916133f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A_c_71_n N_B_M1003_g 0.0265428f $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_68 N_A_c_68_n N_B_M1002_g 0.0117282f $X=0.697 $Y=2.155 $X2=0 $Y2=0
cc_69 N_A_c_73_n N_B_M1002_g 0.0167964f $X=0.697 $Y=2.305 $X2=0 $Y2=0
cc_70 N_A_c_66_n N_B_c_109_n 0.0265428f $X=0.605 $Y=1.345 $X2=0 $Y2=0
cc_71 N_A_c_67_n N_B_c_114_n 0.0265428f $X=0.605 $Y=1.525 $X2=0 $Y2=0
cc_72 N_A_c_66_n B 6.74786e-19 $X=0.605 $Y=1.345 $X2=0 $Y2=0
cc_73 N_A_c_68_n B 4.96571e-19 $X=0.697 $Y=2.155 $X2=0 $Y2=0
cc_74 A B 0.0529376f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_75 N_A_c_70_n N_B_c_111_n 0.0265428f $X=0.59 $Y=1.02 $X2=0 $Y2=0
cc_76 N_A_c_68_n N_A_68_65#_c_223_n 0.00972899f $X=0.697 $Y=2.155 $X2=0 $Y2=0
cc_77 A N_A_68_65#_c_223_n 0.0766385f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A_c_70_n N_A_68_65#_c_223_n 0.0165659f $X=0.59 $Y=1.02 $X2=0 $Y2=0
cc_79 N_A_c_71_n N_A_68_65#_c_223_n 0.00419675f $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_80 N_A_c_73_n N_A_68_65#_c_233_n 0.00572564f $X=0.697 $Y=2.305 $X2=0 $Y2=0
cc_81 A N_A_68_65#_c_224_n 0.0249256f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_82 N_A_c_70_n N_A_68_65#_c_224_n 0.00387137f $X=0.59 $Y=1.02 $X2=0 $Y2=0
cc_83 N_A_c_71_n N_A_68_65#_c_224_n 0.0107029f $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_84 N_A_c_68_n N_A_68_65#_c_234_n 0.00428405f $X=0.697 $Y=2.155 $X2=0 $Y2=0
cc_85 N_A_c_73_n N_A_68_65#_c_234_n 0.0101878f $X=0.697 $Y=2.305 $X2=0 $Y2=0
cc_86 A N_A_68_65#_c_234_n 0.0132846f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A_c_71_n N_A_68_65#_c_226_n 8.56711e-19 $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_88 A N_A_68_65#_c_228_n 0.0107738f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A_c_71_n N_A_68_65#_c_228_n 2.03747e-19 $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_90 N_A_c_67_n N_A_68_65#_c_235_n 0.00269047f $X=0.605 $Y=1.525 $X2=0 $Y2=0
cc_91 N_A_c_68_n N_A_68_65#_c_235_n 0.00175777f $X=0.697 $Y=2.155 $X2=0 $Y2=0
cc_92 N_A_c_73_n N_A_68_65#_c_235_n 0.00263212f $X=0.697 $Y=2.305 $X2=0 $Y2=0
cc_93 A N_A_68_65#_c_235_n 0.00879175f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_94 N_A_c_73_n N_VPWR_c_320_n 0.00363299f $X=0.697 $Y=2.305 $X2=0 $Y2=0
cc_95 N_A_c_73_n N_VPWR_c_323_n 0.00490845f $X=0.697 $Y=2.305 $X2=0 $Y2=0
cc_96 N_A_c_73_n N_VPWR_c_319_n 0.00506877f $X=0.697 $Y=2.305 $X2=0 $Y2=0
cc_97 N_A_c_71_n N_VGND_c_372_n 0.00478647f $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_98 N_A_c_71_n N_VGND_c_373_n 0.00320551f $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_99 N_B_M1003_g N_C_c_157_n 0.0492513f $X=1.07 $Y=0.535 $X2=-0.19 $Y2=-0.245
cc_100 N_B_c_109_n N_C_c_159_n 0.0144397f $X=1.16 $Y=1.75 $X2=0 $Y2=0
cc_101 N_B_M1002_g N_C_c_165_n 0.00810762f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_102 N_B_M1002_g N_C_c_166_n 0.0174118f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_103 N_B_c_114_n N_C_c_167_n 0.0144397f $X=1.16 $Y=1.915 $X2=0 $Y2=0
cc_104 B C 0.0480206f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_111_n C 0.00153225f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B_M1002_g C 0.00121896f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_107 N_B_c_109_n C 5.29116e-19 $X=1.16 $Y=1.75 $X2=0 $Y2=0
cc_108 B C 0.0144933f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B_c_111_n N_C_c_161_n 0.0144397f $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B_M1003_g N_C_c_162_n 0.00773232f $X=1.07 $Y=0.535 $X2=0 $Y2=0
cc_111 B N_C_c_162_n 0.00246218f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B_M1003_g N_A_68_65#_c_224_n 0.0132272f $X=1.07 $Y=0.535 $X2=0 $Y2=0
cc_113 B N_A_68_65#_c_224_n 0.00191969f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B_M1002_g N_A_68_65#_c_234_n 0.0145298f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_115 N_B_c_114_n N_A_68_65#_c_234_n 0.0025531f $X=1.16 $Y=1.915 $X2=0 $Y2=0
cc_116 B N_A_68_65#_c_234_n 0.0258561f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B_M1003_g N_A_68_65#_c_226_n 0.00368329f $X=1.07 $Y=0.535 $X2=0 $Y2=0
cc_118 B N_A_68_65#_c_227_n 0.00830815f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B_c_111_n N_A_68_65#_c_227_n 3.689e-19 $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B_M1003_g N_A_68_65#_c_228_n 0.00468409f $X=1.07 $Y=0.535 $X2=0 $Y2=0
cc_121 B N_A_68_65#_c_228_n 0.0153413f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B_c_111_n N_A_68_65#_c_228_n 7.31855e-19 $X=1.16 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B_M1002_g N_A_68_65#_c_236_n 0.00213184f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_124 N_B_M1002_g N_VPWR_c_320_n 0.00191337f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_125 N_B_M1002_g N_VPWR_c_321_n 0.00490845f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_126 N_B_M1002_g N_VPWR_c_319_n 0.00506877f $X=1.145 $Y=2.625 $X2=0 $Y2=0
cc_127 N_B_M1003_g N_VGND_c_372_n 0.00430609f $X=1.07 $Y=0.535 $X2=0 $Y2=0
cc_128 N_B_M1003_g N_VGND_c_373_n 0.00320497f $X=1.07 $Y=0.535 $X2=0 $Y2=0
cc_129 N_B_M1003_g N_VGND_c_374_n 0.00131637f $X=1.07 $Y=0.535 $X2=0 $Y2=0
cc_130 C N_A_68_65#_c_219_n 0.00179749f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_C_c_161_n N_A_68_65#_c_219_n 0.0128213f $X=1.73 $Y=1.375 $X2=0 $Y2=0
cc_132 N_C_c_162_n N_A_68_65#_c_219_n 0.00412894f $X=1.715 $Y=1.21 $X2=0 $Y2=0
cc_133 N_C_M1000_g N_A_68_65#_M1004_g 0.00520316f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_134 N_C_c_159_n N_A_68_65#_M1004_g 0.0075214f $X=1.715 $Y=1.7 $X2=0 $Y2=0
cc_135 N_C_c_165_n N_A_68_65#_M1004_g 0.00663505f $X=1.592 $Y=2.125 $X2=0 $Y2=0
cc_136 C N_A_68_65#_M1004_g 4.5959e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 C N_A_68_65#_M1004_g 0.00348259f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_138 N_C_c_158_n N_A_68_65#_M1006_g 0.00128655f $X=1.625 $Y=1.005 $X2=0 $Y2=0
cc_139 N_C_c_159_n N_A_68_65#_c_222_n 0.0128213f $X=1.715 $Y=1.7 $X2=0 $Y2=0
cc_140 N_C_c_157_n N_A_68_65#_c_224_n 0.0024816f $X=1.43 $Y=0.855 $X2=0 $Y2=0
cc_141 N_C_c_165_n N_A_68_65#_c_234_n 2.19445e-19 $X=1.592 $Y=2.125 $X2=0 $Y2=0
cc_142 N_C_c_166_n N_A_68_65#_c_234_n 0.00303623f $X=1.592 $Y=2.275 $X2=0 $Y2=0
cc_143 C N_A_68_65#_c_234_n 0.00713451f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_144 N_C_c_157_n N_A_68_65#_c_226_n 0.00345123f $X=1.43 $Y=0.855 $X2=0 $Y2=0
cc_145 N_C_c_157_n N_A_68_65#_c_227_n 0.00430415f $X=1.43 $Y=0.855 $X2=0 $Y2=0
cc_146 N_C_c_158_n N_A_68_65#_c_227_n 0.020593f $X=1.625 $Y=1.005 $X2=0 $Y2=0
cc_147 C N_A_68_65#_c_227_n 0.0291506f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_C_c_161_n N_A_68_65#_c_227_n 0.00111493f $X=1.73 $Y=1.375 $X2=0 $Y2=0
cc_149 N_C_c_158_n N_A_68_65#_c_229_n 0.00100196f $X=1.625 $Y=1.005 $X2=0 $Y2=0
cc_150 C N_A_68_65#_c_229_n 0.0285663f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_151 N_C_c_161_n N_A_68_65#_c_229_n 0.0014674f $X=1.73 $Y=1.375 $X2=0 $Y2=0
cc_152 N_C_c_158_n N_A_68_65#_c_230_n 0.00412894f $X=1.625 $Y=1.005 $X2=0 $Y2=0
cc_153 N_C_c_166_n N_A_68_65#_c_236_n 0.00340232f $X=1.592 $Y=2.275 $X2=0 $Y2=0
cc_154 N_C_M1000_g N_VPWR_c_321_n 0.00490845f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_155 N_C_M1000_g N_VPWR_c_322_n 0.00370693f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_156 N_C_c_166_n N_VPWR_c_322_n 8.61462e-19 $X=1.592 $Y=2.275 $X2=0 $Y2=0
cc_157 N_C_c_167_n N_VPWR_c_322_n 8.79542e-19 $X=1.715 $Y=1.88 $X2=0 $Y2=0
cc_158 C N_VPWR_c_322_n 0.0188265f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_159 N_C_M1000_g N_VPWR_c_319_n 0.00506877f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_160 C X 0.00336792f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_161 C X 0.0137067f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_162 N_C_c_157_n N_VGND_c_372_n 0.00403983f $X=1.43 $Y=0.855 $X2=0 $Y2=0
cc_163 N_C_c_157_n N_VGND_c_373_n 0.00414769f $X=1.43 $Y=0.855 $X2=0 $Y2=0
cc_164 N_C_c_157_n N_VGND_c_374_n 0.010971f $X=1.43 $Y=0.855 $X2=0 $Y2=0
cc_165 N_C_c_158_n N_VGND_c_374_n 0.00137447f $X=1.625 $Y=1.005 $X2=0 $Y2=0
cc_166 N_A_68_65#_c_234_n N_VPWR_c_320_n 0.0155785f $X=1.225 $Y=2.18 $X2=0 $Y2=0
cc_167 N_A_68_65#_c_292_p N_VPWR_c_321_n 0.00512477f $X=1.36 $Y=2.625 $X2=0
+ $Y2=0
cc_168 N_A_68_65#_M1004_g N_VPWR_c_322_n 0.0090162f $X=2.345 $Y=2.735 $X2=0
+ $Y2=0
cc_169 N_A_68_65#_c_236_n N_VPWR_c_322_n 0.00254124f $X=1.355 $Y=2.46 $X2=0
+ $Y2=0
cc_170 N_A_68_65#_c_233_n N_VPWR_c_323_n 0.0110039f $X=0.5 $Y=2.625 $X2=0 $Y2=0
cc_171 N_A_68_65#_M1004_g N_VPWR_c_325_n 0.00545548f $X=2.345 $Y=2.735 $X2=0
+ $Y2=0
cc_172 N_A_68_65#_M1004_g N_VPWR_c_319_n 0.0120531f $X=2.345 $Y=2.735 $X2=0
+ $Y2=0
cc_173 N_A_68_65#_c_233_n N_VPWR_c_319_n 0.0152283f $X=0.5 $Y=2.625 $X2=0 $Y2=0
cc_174 N_A_68_65#_c_292_p N_VPWR_c_319_n 0.00832937f $X=1.36 $Y=2.625 $X2=0
+ $Y2=0
cc_175 N_A_68_65#_M1004_g X 0.0231014f $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_176 N_A_68_65#_M1006_g X 0.0246475f $X=2.405 $Y=0.535 $X2=0 $Y2=0
cc_177 N_A_68_65#_c_227_n X 0.014009f $X=2.105 $Y=0.915 $X2=0 $Y2=0
cc_178 N_A_68_65#_c_229_n X 0.0475921f $X=2.27 $Y=1.12 $X2=0 $Y2=0
cc_179 N_A_68_65#_M1004_g X 7.06088e-19 $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_180 N_A_68_65#_c_224_n A_157_65# 0.00456566f $X=1.09 $Y=0.52 $X2=-0.19
+ $Y2=-0.245
cc_181 N_A_68_65#_c_224_n A_229_65# 0.00357971f $X=1.09 $Y=0.52 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_68_65#_c_226_n A_229_65# 8.23851e-19 $X=1.175 $Y=0.83 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_68_65#_M1006_g N_VGND_c_371_n 0.00414769f $X=2.405 $Y=0.535 $X2=0
+ $Y2=0
cc_184 N_A_68_65#_M1006_g N_VGND_c_372_n 0.00818536f $X=2.405 $Y=0.535 $X2=0
+ $Y2=0
cc_185 N_A_68_65#_c_224_n N_VGND_c_372_n 0.0318499f $X=1.09 $Y=0.52 $X2=0 $Y2=0
cc_186 N_A_68_65#_c_225_n N_VGND_c_372_n 0.00620247f $X=0.325 $Y=0.52 $X2=0
+ $Y2=0
cc_187 N_A_68_65#_c_227_n N_VGND_c_372_n 0.00970208f $X=2.105 $Y=0.915 $X2=0
+ $Y2=0
cc_188 N_A_68_65#_c_224_n N_VGND_c_373_n 0.0313118f $X=1.09 $Y=0.52 $X2=0 $Y2=0
cc_189 N_A_68_65#_c_225_n N_VGND_c_373_n 0.00702119f $X=0.325 $Y=0.52 $X2=0
+ $Y2=0
cc_190 N_A_68_65#_M1006_g N_VGND_c_374_n 0.0134927f $X=2.405 $Y=0.535 $X2=0
+ $Y2=0
cc_191 N_A_68_65#_c_224_n N_VGND_c_374_n 0.0206746f $X=1.09 $Y=0.52 $X2=0 $Y2=0
cc_192 N_A_68_65#_c_227_n N_VGND_c_374_n 0.0669735f $X=2.105 $Y=0.915 $X2=0
+ $Y2=0
cc_193 N_A_68_65#_c_230_n N_VGND_c_374_n 0.00115966f $X=2.27 $Y=1.12 $X2=0 $Y2=0
cc_194 N_VPWR_c_325_n X 0.024468f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_319_n X 0.0140441f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_322_n X 0.00245941f $X=1.79 $Y=2.56 $X2=0 $Y2=0
cc_197 X N_VGND_c_371_n 0.0117077f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_198 X N_VGND_c_372_n 0.00992777f $X=2.555 $Y=0.47 $X2=0 $Y2=0
