* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a32oi_0 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR A3 a_37_397# VPB phighvt w=640000u l=150000u
+  ad=5.664e+11p pd=4.33e+06u as=5.28e+11p ps=5.49e+06u
M1001 Y B2 a_37_397# VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1002 Y B1 a_141_47# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=1.008e+11p ps=1.32e+06u
M1003 VPWR A1 a_37_397# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_447_47# A2 a_333_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.764e+11p ps=1.68e+06u
M1005 a_141_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.499e+11p ps=2.87e+06u
M1006 a_37_397# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A3 a_447_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_37_397# B1 Y VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_333_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
