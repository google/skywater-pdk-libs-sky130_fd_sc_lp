# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__xnor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.425000 1.655000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.185000 0.440000 1.920000 ;
        RECT 0.085000 1.920000 1.995000 2.090000 ;
        RECT 1.825000 1.425000 2.465000 1.845000 ;
        RECT 1.825000 1.845000 1.995000 1.920000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.657300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 2.355000 3.275000 2.555000 ;
        RECT 2.505000 2.555000 2.765000 3.075000 ;
        RECT 3.015000 0.255000 3.275000 1.175000 ;
        RECT 3.015000 1.845000 3.275000 2.355000 ;
        RECT 3.095000 1.175000 3.275000 1.845000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 3.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.125000  0.265000 0.455000 0.845000 ;
      RECT 0.125000  0.845000 0.780000 1.015000 ;
      RECT 0.125000  2.260000 0.385000 3.245000 ;
      RECT 0.555000  2.260000 2.335000 2.430000 ;
      RECT 0.555000  2.430000 0.815000 3.075000 ;
      RECT 0.610000  1.015000 0.780000 1.085000 ;
      RECT 0.610000  1.085000 2.845000 1.255000 ;
      RECT 0.950000  0.085000 1.280000 0.915000 ;
      RECT 0.985000  2.600000 1.825000 3.245000 ;
      RECT 1.470000  0.255000 1.800000 0.745000 ;
      RECT 1.470000  0.745000 2.835000 0.915000 ;
      RECT 1.970000  0.085000 2.300000 0.575000 ;
      RECT 2.165000  2.015000 2.845000 2.185000 ;
      RECT 2.165000  2.185000 2.335000 2.260000 ;
      RECT 2.505000  0.255000 2.835000 0.745000 ;
      RECT 2.675000  1.255000 2.845000 1.345000 ;
      RECT 2.675000  1.345000 2.925000 1.675000 ;
      RECT 2.675000  1.675000 2.845000 2.015000 ;
      RECT 2.935000  2.725000 3.265000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__xnor2_1
END LIBRARY
