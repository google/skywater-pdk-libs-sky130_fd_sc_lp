# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.580000 1.210000 2.075000 1.790000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.775000 0.255000 8.065000 3.075000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.425000 2.155000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 0.670000 ;
      RECT 0.095000  2.325000 0.425000 3.245000 ;
      RECT 0.595000  0.400000 0.855000 0.955000 ;
      RECT 0.595000  0.955000 1.010000 1.625000 ;
      RECT 0.595000  1.625000 0.795000 2.990000 ;
      RECT 1.045000  2.045000 2.075000 2.130000 ;
      RECT 1.045000  2.130000 1.340000 2.715000 ;
      RECT 1.180000  0.855000 1.410000 1.960000 ;
      RECT 1.180000  1.960000 2.075000 2.045000 ;
      RECT 1.510000  2.300000 1.735000 3.245000 ;
      RECT 1.710000  0.085000 2.040000 1.040000 ;
      RECT 1.905000  2.130000 2.075000 2.605000 ;
      RECT 1.905000  2.605000 3.495000 2.880000 ;
      RECT 2.245000  0.860000 2.575000 1.190000 ;
      RECT 2.245000  1.190000 2.425000 2.435000 ;
      RECT 2.595000  1.575000 2.775000 2.605000 ;
      RECT 2.755000  0.860000 3.125000 1.105000 ;
      RECT 2.755000  1.105000 4.240000 1.190000 ;
      RECT 2.945000  1.190000 4.240000 1.275000 ;
      RECT 2.945000  1.275000 3.155000 2.435000 ;
      RECT 3.325000  2.285000 4.930000 2.455000 ;
      RECT 3.325000  2.455000 3.495000 2.605000 ;
      RECT 3.370000  1.445000 3.700000 1.855000 ;
      RECT 3.370000  1.855000 4.580000 2.115000 ;
      RECT 3.570000  0.085000 4.240000 0.935000 ;
      RECT 3.760000  2.635000 4.090000 3.245000 ;
      RECT 3.980000  1.275000 4.240000 1.675000 ;
      RECT 4.410000  0.575000 4.685000 1.245000 ;
      RECT 4.410000  1.245000 4.580000 1.855000 ;
      RECT 4.760000  1.425000 5.035000 1.595000 ;
      RECT 4.760000  1.595000 4.930000 2.285000 ;
      RECT 4.855000  1.195000 5.035000 1.425000 ;
      RECT 4.990000  0.640000 5.395000 0.970000 ;
      RECT 5.110000  1.875000 5.375000 2.755000 ;
      RECT 5.205000  0.970000 5.395000 1.125000 ;
      RECT 5.205000  1.125000 6.595000 1.295000 ;
      RECT 5.205000  1.295000 5.375000 1.875000 ;
      RECT 5.790000  1.465000 6.120000 1.625000 ;
      RECT 5.790000  1.625000 7.605000 1.655000 ;
      RECT 5.790000  1.655000 6.935000 1.795000 ;
      RECT 5.975000  0.085000 6.305000 0.945000 ;
      RECT 5.980000  1.965000 6.360000 3.245000 ;
      RECT 6.335000  1.295000 6.595000 1.455000 ;
      RECT 6.475000  0.415000 6.935000 0.945000 ;
      RECT 6.540000  1.795000 6.935000 2.750000 ;
      RECT 6.765000  0.945000 7.170000 1.270000 ;
      RECT 6.765000  1.270000 7.605000 1.625000 ;
      RECT 7.305000  1.825000 7.605000 3.245000 ;
      RECT 7.340000  0.085000 7.605000 1.095000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__dfxtp_1
END LIBRARY
