* NGSPICE file created from sky130_fd_sc_lp__sdfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_225_50# SCD a_512_81# VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_894_463# a_864_255# a_808_463# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.289e+11p ps=2.77e+06u
M1002 VPWR a_864_255# a_756_265# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.72075e+12p pd=2.2e+07u as=3.339e+11p ps=3.05e+06u
M1003 a_308_50# a_35_74# a_225_50# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VPWR a_936_333# a_894_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1085_119# a_936_333# a_991_119# VNB nshort w=420000u l=150000u
+  ad=1.554e+11p pd=1.62e+06u as=1.344e+11p ps=1.48e+06u
M1006 VGND a_864_255# a_756_265# VNB nshort w=840000u l=150000u
+  ad=1.6517e+12p pd=1.461e+07u as=2.394e+11p ps=2.25e+06u
M1007 a_332_468# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1008 a_864_255# CLK VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1009 a_1406_69# a_864_255# a_936_333# VPB phighvt w=840000u l=150000u
+  ad=4.3735e+11p pd=3.33e+06u as=2.352e+11p ps=2.24e+06u
M1010 VPWR a_2431_47# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1011 VGND a_1406_69# a_2431_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 VPWR SCD a_490_468# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1013 a_808_463# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1635_21# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1015 a_1406_69# a_756_265# a_936_333# VNB nshort w=640000u l=150000u
+  ad=3.88e+11p pd=2.85e+06u as=1.792e+11p ps=1.84e+06u
M1016 a_808_463# a_756_265# a_380_50# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.95e+11p ps=3.87e+06u
M1017 VGND a_1635_21# a_1593_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1018 a_490_468# a_35_74# a_380_50# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND RESET_B a_225_50# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_864_255# CLK VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1021 a_1569_534# a_756_265# a_1406_69# VPB phighvt w=420000u l=150000u
+  ad=1.848e+11p pd=1.72e+06u as=0p ps=0u
M1022 VPWR SCE a_35_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1023 VGND SCE a_35_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1024 Q a_2431_47# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1025 a_936_333# a_808_463# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_380_50# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1593_113# a_864_255# a_1406_69# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_1406_69# a_2431_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1029 Q a_2431_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_936_333# a_808_463# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_808_463# a_864_255# a_380_50# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=4.1875e+11p ps=3.77e+06u
M1032 a_380_50# D a_332_468# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_380_50# D a_308_50# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1809_119# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1035 VPWR a_1635_21# a_1569_534# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_991_119# a_756_265# a_808_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND RESET_B a_1085_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_1406_69# a_1635_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_512_81# SCE a_380_50# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1635_21# a_1406_69# a_1809_119# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1041 VGND a_2431_47# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

