* NGSPICE file created from sky130_fd_sc_lp__dlrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 VPWR a_267_464# a_414_47# VPB phighvt w=640000u l=150000u
+  ad=2.4044e+12p pd=1.823e+07u as=1.696e+11p ps=1.81e+06u
M1001 VGND D a_49_70# VNB nshort w=420000u l=150000u
+  ad=1.1865e+12p pd=1.156e+07u as=1.113e+11p ps=1.37e+06u
M1002 VGND a_267_464# a_414_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 Q a_857_21# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1004 a_651_469# a_49_70# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1005 Q a_857_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR D a_49_70# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1007 VPWR RESET_B a_857_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1008 Q a_857_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1009 a_671_47# a_414_47# a_599_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=8.82e+10p ps=1.26e+06u
M1010 VPWR a_857_21# a_828_469# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=9.45e+10p ps=1.29e+06u
M1011 VGND a_857_21# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_599_47# a_49_70# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1083_73# a_671_47# a_857_21# VNB nshort w=840000u l=150000u
+  ad=3.024e+11p pd=2.4e+06u as=2.226e+11p ps=2.21e+06u
M1014 a_857_21# a_671_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_857_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_828_469# a_414_47# a_671_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.158e+11p ps=2.03e+06u
M1017 a_779_47# a_267_464# a_671_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1018 VPWR a_857_21# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_857_21# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_671_47# a_267_464# a_651_469# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND RESET_B a_1083_73# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_267_464# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1023 VPWR a_857_21# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_857_21# a_779_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_267_464# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

