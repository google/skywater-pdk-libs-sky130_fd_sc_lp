* File: sky130_fd_sc_lp__a211oi_m.pex.spice
* Created: Wed Sep  2 09:18:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211OI_M%A2 3 6 9 10 13 14 15 19
r28 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.925
+ $X2=0.29 $Y2=1.295
r29 14 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=0.93 $X2=0.29 $Y2=0.93
r30 12 19 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.29 $Y=1.285
+ $X2=0.29 $Y2=0.93
r31 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.337 $Y=1.285
+ $X2=0.337 $Y2=1.435
r32 10 19 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.29 $Y=0.915
+ $X2=0.29 $Y2=0.93
r33 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.337 $Y=0.765
+ $X2=0.337 $Y2=0.915
r34 6 13 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.475 $Y=2.055
+ $X2=0.475 $Y2=1.435
r35 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_M%A1 3 7 11 12 13 16 17
r37 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.08 $X2=0.925 $Y2=1.08
r38 13 17 4.80777 $w=5.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.25
+ $X2=0.925 $Y2=1.25
r39 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.925 $Y=1.42
+ $X2=0.925 $Y2=1.08
r40 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.42
+ $X2=0.925 $Y2=1.585
r41 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=0.915
+ $X2=0.925 $Y2=1.08
r42 7 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.015 $Y=2.055 $X2=1.015
+ $Y2=1.585
r43 3 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.835 $Y=0.445 $X2=0.835
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_M%B1 3 7 11 12 13 16
r36 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.465
+ $Y=1.08 $X2=1.465 $Y2=1.08
r37 13 17 5.04229 $w=5.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.25
+ $X2=1.465 $Y2=1.25
r38 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.465 $Y=1.42
+ $X2=1.465 $Y2=1.08
r39 11 12 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.42
+ $X2=1.465 $Y2=1.585
r40 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=0.915
+ $X2=1.465 $Y2=1.08
r41 7 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.495 $Y=2.055 $X2=1.495
+ $Y2=1.585
r42 3 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.375 $Y=0.445 $X2=1.375
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_M%C1 3 6 7 8 9 10
r29 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.825
+ $Y=2.78 $X2=1.825 $Y2=2.78
r30 10 16 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=1.85 $Y=2.775
+ $X2=1.825 $Y2=2.775
r31 9 10 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.047 $Y=2.405
+ $X2=2.047 $Y2=2.775
r32 8 16 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=2.775
+ $X2=1.825 $Y2=2.775
r33 7 15 2.54577 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=1.84 $Y=2.775
+ $X2=1.825 $Y2=2.775
r34 3 6 825.553 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=1.915 $Y=0.445
+ $X2=1.915 $Y2=2.055
r35 1 7 32.5671 $w=3.4e-07 $l=2.04083e-07 $layer=POLY_cond $X=1.915 $Y=2.605
+ $X2=1.84 $Y2=2.775
r36 1 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.915 $Y=2.605
+ $X2=1.915 $Y2=2.055
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_M%A_27_369# 1 2 11 12 15
r19 13 15 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.23 $Y=1.855
+ $X2=1.23 $Y2=1.97
r20 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.125 $Y=1.77
+ $X2=1.23 $Y2=1.855
r21 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.125 $Y=1.77
+ $X2=0.365 $Y2=1.77
r22 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.26 $Y=1.855
+ $X2=0.365 $Y2=1.77
r23 7 9 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.26 $Y=1.855
+ $X2=0.26 $Y2=1.99
r24 2 15 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.845 $X2=1.23 $Y2=1.97
r25 1 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_M%VPWR 1 6 8 10 20 21 24
r18 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r19 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r20 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r21 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.71 $Y2=3.33
r22 15 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=1.2 $Y2=3.33
r23 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r24 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r25 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.71 $Y2=3.33
r26 10 12 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 8 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r28 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.72
+ $Y2=3.33
r29 8 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=3.245 $X2=0.71
+ $Y2=3.33
r31 4 6 38.5894 $w=3.28e-07 $l=1.105e-06 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=2.14
r32 1 6 600 $w=1.7e-07 $l=3.66367e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.845 $X2=0.71 $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_M%Y 1 2 3 12 14 15 18 21 22 23 24 25
r38 24 25 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.99
r39 23 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=1.295
+ $X2=2.13 $Y2=1.665
r40 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=0.925
+ $X2=2.13 $Y2=1.295
r41 20 22 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.13 $Y=0.815
+ $X2=2.13 $Y2=0.925
r42 20 21 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.815 $X2=2.13
+ $Y2=0.73
r43 16 21 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=2.16 $Y=0.645
+ $X2=2.13 $Y2=0.73
r44 16 18 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.16 $Y=0.645
+ $X2=2.16 $Y2=0.51
r45 14 21 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=0.73
+ $X2=2.13 $Y2=0.73
r46 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.965 $Y=0.73
+ $X2=1.265 $Y2=0.73
r47 10 15 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.16 $Y=0.645
+ $X2=1.265 $Y2=0.73
r48 10 12 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.16 $Y=0.645
+ $X2=1.16 $Y2=0.51
r49 3 25 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.845 $X2=2.13 $Y2=1.99
r50 2 18 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.235 $X2=2.13 $Y2=0.51
r51 1 12 182 $w=1.7e-07 $l=3.79967e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.16 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_M%VGND 1 2 7 9 13 15 17 24 25 31
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r39 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 25 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r41 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.61
+ $Y2=0
r43 22 24 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=2.16
+ $Y2=0
r44 18 28 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r45 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=1.2
+ $Y2=0
r46 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.61
+ $Y2=0
r47 17 20 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.2
+ $Y2=0
r48 15 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r49 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r50 15 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0
r52 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0.36
r53 7 28 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r54 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r55 2 13 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.61 $Y2=0.36
r56 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

