* File: sky130_fd_sc_lp__busdrivernovlp_20.pex.spice
* Created: Fri Aug 28 10:13:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%TE_B 3 5 7 9 10 11 12 14 15 17 19
+ 22 26 29 30 31 34 35 36 37 38 39 40 42 43 44 46 47 48 50 53 57 58 60 66 72
c203 39 0 1.45114e-19 $X=3.335 $Y=0.935
c204 5 0 3.30551e-20 $X=0.93 $Y=0.955
r205 67 72 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.67 $Y=1.16 $X2=0.67
+ $Y2=1.08
r206 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.16 $X2=0.67 $Y2=1.16
r207 64 66 29.8306 $w=3.07e-07 $l=1.9e-07 $layer=POLY_cond $X=0.48 $Y=1.14
+ $X2=0.67 $Y2=1.14
r208 60 67 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.67 $Y=1.295
+ $X2=0.67 $Y2=1.16
r209 58 71 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.125 $Y=1.16
+ $X2=6.125 $Y2=1.325
r210 58 70 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.125 $Y=1.16
+ $X2=6.125 $Y2=0.995
r211 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.115
+ $Y=1.16 $X2=6.115 $Y2=1.16
r212 54 57 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.9 $Y=1.16
+ $X2=6.115 $Y2=1.16
r213 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.64
+ $Y=0.43 $X2=2.64 $Y2=0.43
r214 50 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.9 $Y=0.995
+ $X2=5.9 $Y2=1.16
r215 49 50 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.9 $Y=0.815
+ $X2=5.9 $Y2=0.995
r216 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.815 $Y=0.73
+ $X2=5.9 $Y2=0.815
r217 47 48 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=5.815 $Y=0.73
+ $X2=4.205 $Y2=0.73
r218 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.12 $Y=0.645
+ $X2=4.205 $Y2=0.73
r219 45 46 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.12 $Y=0.435
+ $X2=4.12 $Y2=0.645
r220 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.035 $Y=0.35
+ $X2=4.12 $Y2=0.435
r221 43 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.035 $Y=0.35
+ $X2=3.505 $Y2=0.35
r222 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=0.435
+ $X2=3.505 $Y2=0.35
r223 41 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.42 $Y=0.435
+ $X2=3.42 $Y2=0.85
r224 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.935
+ $X2=3.42 $Y2=0.85
r225 39 40 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.335 $Y=0.935
+ $X2=2.805 $Y2=0.935
r226 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.64 $Y=0.85
+ $X2=2.805 $Y2=0.935
r227 37 52 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.435
+ $X2=2.64 $Y2=0.35
r228 37 38 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.64 $Y=0.435
+ $X2=2.64 $Y2=0.85
r229 35 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0.35
+ $X2=2.64 $Y2=0.35
r230 35 36 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.475 $Y=0.35
+ $X2=1.74 $Y2=0.35
r231 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.655 $Y=0.435
+ $X2=1.74 $Y2=0.35
r232 33 34 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.655 $Y=0.435
+ $X2=1.655 $Y2=0.995
r233 32 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=1.08
+ $X2=0.67 $Y2=1.08
r234 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=1.08
+ $X2=1.655 $Y2=0.995
r235 31 32 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.57 $Y=1.08
+ $X2=0.835 $Y2=1.08
r236 28 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.64 $Y=0.77
+ $X2=2.64 $Y2=0.43
r237 28 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=0.77
+ $X2=2.64 $Y2=0.935
r238 26 71 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.225 $Y=2.285
+ $X2=6.225 $Y2=1.325
r239 22 70 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.115 $Y=0.445
+ $X2=6.115 $Y2=0.995
r240 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.985 $Y=1.185
+ $X2=3.985 $Y2=0.655
r241 16 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.63 $Y=1.26
+ $X2=3.555 $Y2=1.26
r242 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.91 $Y=1.26
+ $X2=3.985 $Y2=1.185
r243 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.91 $Y=1.26
+ $X2=3.63 $Y2=1.26
r244 12 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.555 $Y=1.185
+ $X2=3.555 $Y2=1.26
r245 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.555 $Y=1.185
+ $X2=3.555 $Y2=0.655
r246 10 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.48 $Y=1.26
+ $X2=3.555 $Y2=1.26
r247 10 11 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.48 $Y=1.26
+ $X2=2.805 $Y2=1.26
r248 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.73 $Y=1.185
+ $X2=2.805 $Y2=1.26
r249 9 29 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.73 $Y=1.185
+ $X2=2.73 $Y2=0.935
r250 5 66 40.8208 $w=3.07e-07 $l=3.40147e-07 $layer=POLY_cond $X=0.93 $Y=0.955
+ $X2=0.67 $Y2=1.14
r251 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.93 $Y=0.955
+ $X2=0.93 $Y2=0.635
r252 1 64 19.5117 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.14
r253 1 3 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=2.255
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A_27_367# 1 2 7 9 12 14 16 17 18
+ 21 24 27 29 30 31 33 35 40
c105 29 0 3.30551e-20 $X=0.55 $Y=0.73
c106 17 0 1.14036e-19 $X=1.875 $Y=1.64
c107 14 0 3.92328e-20 $X=1.44 $Y=1.715
c108 12 0 9.82022e-20 $X=1.44 $Y=0.635
r109 41 47 29.2588 $w=3.13e-07 $l=1.9e-07 $layer=POLY_cond $X=1.25 $Y=1.53
+ $X2=1.44 $Y2=1.53
r110 40 43 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=1.51
+ $X2=1.25 $Y2=1.675
r111 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.51 $X2=1.25 $Y2=1.51
r112 35 37 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.715 $Y=0.61
+ $X2=0.715 $Y2=0.73
r113 32 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.43 $Y=1.675
+ $X2=0.265 $Y2=1.675
r114 31 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=1.675
+ $X2=1.25 $Y2=1.675
r115 31 32 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.085 $Y=1.675
+ $X2=0.43 $Y2=1.675
r116 29 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0.73
+ $X2=0.715 $Y2=0.73
r117 29 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.55 $Y=0.73
+ $X2=0.27 $Y2=0.73
r118 25 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=1.76
+ $X2=0.265 $Y2=1.675
r119 25 27 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.265 $Y=1.76
+ $X2=0.265 $Y2=1.98
r120 24 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.185 $Y=1.59
+ $X2=0.265 $Y2=1.675
r121 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.185 $Y=0.815
+ $X2=0.27 $Y2=0.73
r122 23 24 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.185 $Y=0.815
+ $X2=0.185 $Y2=1.59
r123 19 21 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.95 $Y=1.715
+ $X2=1.95 $Y2=2.675
r124 18 47 24.674 $w=3.13e-07 $l=1.42653e-07 $layer=POLY_cond $X=1.515 $Y=1.64
+ $X2=1.44 $Y2=1.53
r125 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.875 $Y=1.64
+ $X2=1.95 $Y2=1.715
r126 17 18 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.875 $Y=1.64
+ $X2=1.515 $Y2=1.64
r127 14 47 19.9686 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.44 $Y=1.715
+ $X2=1.44 $Y2=1.53
r128 14 16 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.44 $Y=1.715 $X2=1.44
+ $Y2=2.465
r129 10 47 19.9686 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.44 $Y=1.345
+ $X2=1.44 $Y2=1.53
r130 10 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.44 $Y=1.345
+ $X2=1.44 $Y2=0.635
r131 7 41 36.9585 $w=3.13e-07 $l=3.19374e-07 $layer=POLY_cond $X=1.01 $Y=1.715
+ $X2=1.25 $Y2=1.53
r132 7 9 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.01 $Y=1.715 $X2=1.01
+ $Y2=2.465
r133 2 27 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.835 $X2=0.265 $Y2=1.98
r134 1 35 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.425 $X2=0.715 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A_217_367# 1 2 3 12 14 15 20 22 24
+ 25 26 27 29 30 32 34 35 37 39 40 42 44 45 47 49 50 52 54 55 57 59 60 62 64 65
+ 67 69 70 72 74 75 77 79 80 82 83 85 86 88 89 91 92 94 95 97 98 100 101 103 104
+ 105 106 107 108 109 110 111 112 113 114 116 118 121 123 126 130 131 133 137
+ 141 144 145 146 149 160 168 169 170 175 180 185 190 191 208
c502 168 0 3.75487e-20 $X=2.4 $Y=1.74
c503 145 0 5.44897e-19 $X=2.305 $Y=1.665
c504 144 0 3.02269e-19 $X=9.215 $Y=1.665
c505 123 0 6.94902e-20 $X=1.765 $Y=1.635
c506 26 0 3.81595e-20 $X=9.165 $Y=1.65
r507 190 192 40.8145 $w=3.72e-07 $l=3.15e-07 $layer=POLY_cond $X=16.945 $Y=1.535
+ $X2=17.26 $Y2=1.535
r508 190 191 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=16.945
+ $Y=1.51 $X2=16.945 $Y2=1.51
r509 188 190 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=16.83 $Y=1.535
+ $X2=16.945 $Y2=1.535
r510 187 188 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=16.4 $Y=1.535
+ $X2=16.83 $Y2=1.535
r511 186 187 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=15.97 $Y=1.535
+ $X2=16.4 $Y2=1.535
r512 184 186 29.1532 $w=3.72e-07 $l=2.25e-07 $layer=POLY_cond $X=15.745 $Y=1.535
+ $X2=15.97 $Y2=1.535
r513 184 185 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.745
+ $Y=1.51 $X2=15.745 $Y2=1.51
r514 182 184 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=15.54 $Y=1.535
+ $X2=15.745 $Y2=1.535
r515 181 182 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=15.11 $Y=1.535
+ $X2=15.54 $Y2=1.535
r516 179 181 29.1532 $w=3.72e-07 $l=2.25e-07 $layer=POLY_cond $X=14.885 $Y=1.535
+ $X2=15.11 $Y2=1.535
r517 179 180 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.885
+ $Y=1.51 $X2=14.885 $Y2=1.51
r518 177 179 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=14.68 $Y=1.535
+ $X2=14.885 $Y2=1.535
r519 176 177 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=14.25 $Y=1.535
+ $X2=14.68 $Y2=1.535
r520 174 176 29.1532 $w=3.72e-07 $l=2.25e-07 $layer=POLY_cond $X=14.025 $Y=1.535
+ $X2=14.25 $Y2=1.535
r521 174 175 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.025
+ $Y=1.51 $X2=14.025 $Y2=1.51
r522 168 171 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=1.74
+ $X2=2.4 $Y2=1.905
r523 168 170 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=1.74
+ $X2=2.4 $Y2=1.575
r524 168 169 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=1.74 $X2=2.4 $Y2=1.74
r525 165 169 7.79116 $w=3.53e-07 $l=2.4e-07 $layer=LI1_cond $X=2.16 $Y=1.727
+ $X2=2.4 $Y2=1.727
r526 165 208 6.8759 $w=3.53e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.727
+ $X2=2.045 $Y2=1.727
r527 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.665
r528 160 191 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.965 $Y=1.665
+ $X2=16.965 $Y2=1.665
r529 157 160 0.782757 $w=2.3e-07 $l=1.22e-06 $layer=MET1_cond $X=15.745 $Y=1.665
+ $X2=16.965 $Y2=1.665
r530 157 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.745 $Y=1.665
+ $X2=15.745 $Y2=1.665
r531 154 157 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=14.885 $Y=1.665
+ $X2=15.745 $Y2=1.665
r532 154 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.885 $Y=1.665
+ $X2=14.885 $Y2=1.665
r533 151 154 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=14.025 $Y=1.665
+ $X2=14.885 $Y2=1.665
r534 151 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.025 $Y=1.665
+ $X2=14.025 $Y2=1.665
r535 148 151 2.99308 $w=2.3e-07 $l=4.665e-06 $layer=MET1_cond $X=9.36 $Y=1.665
+ $X2=14.025 $Y2=1.665
r536 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.665
r537 146 148 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=9.33 $Y=1.665
+ $X2=9.36 $Y2=1.665
r538 145 164 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=1.665
+ $X2=2.16 $Y2=1.665
r539 144 146 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=9.33 $Y2=1.665
r540 144 145 8.55196 $w=1.4e-07 $l=6.91e-06 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=2.305 $Y2=1.665
r541 141 149 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=9.04 $Y=1.665
+ $X2=9.36 $Y2=1.665
r542 141 142 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.955 $Y=1.665
+ $X2=8.955 $Y2=1.87
r543 137 139 12.2323 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=8.862 $Y=0.815
+ $X2=8.862 $Y2=1.095
r544 133 141 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.955 $Y=1.55
+ $X2=8.955 $Y2=1.665
r545 133 139 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=8.955 $Y=1.55
+ $X2=8.955 $Y2=1.095
r546 130 142 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=1.87
+ $X2=8.955 $Y2=1.87
r547 130 131 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.87 $Y=1.87
+ $X2=8.025 $Y2=1.87
r548 126 128 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=7.86 $Y=1.98
+ $X2=7.86 $Y2=2.9
r549 124 131 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.86 $Y=1.955
+ $X2=8.025 $Y2=1.87
r550 124 126 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=7.86 $Y=1.955
+ $X2=7.86 $Y2=1.98
r551 123 208 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.765 $Y=1.635
+ $X2=2.045 $Y2=1.635
r552 120 123 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=1.72
+ $X2=1.765 $Y2=1.635
r553 120 121 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.68 $Y=1.72
+ $X2=1.68 $Y2=1.94
r554 119 135 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=2.025
+ $X2=1.225 $Y2=2.025
r555 118 121 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.595 $Y=2.025
+ $X2=1.68 $Y2=1.94
r556 118 119 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.595 $Y=2.025
+ $X2=1.39 $Y2=2.025
r557 114 135 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=2.11
+ $X2=1.225 $Y2=2.025
r558 114 116 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.225 $Y=2.11
+ $X2=1.225 $Y2=2.9
r559 101 192 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=17.26 $Y=1.725
+ $X2=17.26 $Y2=1.535
r560 101 103 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=17.26 $Y=1.725
+ $X2=17.26 $Y2=2.465
r561 98 188 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=16.83 $Y=1.725
+ $X2=16.83 $Y2=1.535
r562 98 100 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=16.83 $Y=1.725
+ $X2=16.83 $Y2=2.465
r563 95 187 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=16.4 $Y=1.725
+ $X2=16.4 $Y2=1.535
r564 95 97 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=16.4 $Y=1.725
+ $X2=16.4 $Y2=2.465
r565 92 186 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=15.97 $Y=1.725
+ $X2=15.97 $Y2=1.535
r566 92 94 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=15.97 $Y=1.725
+ $X2=15.97 $Y2=2.465
r567 89 182 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=15.54 $Y=1.725
+ $X2=15.54 $Y2=1.535
r568 89 91 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=15.54 $Y=1.725
+ $X2=15.54 $Y2=2.465
r569 86 181 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=15.11 $Y=1.725
+ $X2=15.11 $Y2=1.535
r570 86 88 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=15.11 $Y=1.725
+ $X2=15.11 $Y2=2.465
r571 83 177 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=14.68 $Y=1.725
+ $X2=14.68 $Y2=1.535
r572 83 85 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=14.68 $Y=1.725
+ $X2=14.68 $Y2=2.465
r573 80 176 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=14.25 $Y=1.725
+ $X2=14.25 $Y2=1.535
r574 80 82 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=14.25 $Y=1.725
+ $X2=14.25 $Y2=2.465
r575 77 174 26.5618 $w=3.72e-07 $l=2.84561e-07 $layer=POLY_cond $X=13.82
+ $Y=1.725 $X2=14.025 $Y2=1.535
r576 77 79 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=13.82 $Y=1.725
+ $X2=13.82 $Y2=2.465
r577 76 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.465 $Y=1.65
+ $X2=13.39 $Y2=1.65
r578 75 77 27.4257 $w=3.72e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.745 $Y=1.65
+ $X2=13.82 $Y2=1.725
r579 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=13.745 $Y=1.65
+ $X2=13.465 $Y2=1.65
r580 72 113 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.39 $Y=1.725
+ $X2=13.39 $Y2=1.65
r581 72 74 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=13.39 $Y=1.725
+ $X2=13.39 $Y2=2.465
r582 71 112 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.035 $Y=1.65
+ $X2=12.96 $Y2=1.65
r583 70 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.315 $Y=1.65
+ $X2=13.39 $Y2=1.65
r584 70 71 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=13.315 $Y=1.65
+ $X2=13.035 $Y2=1.65
r585 67 112 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.96 $Y=1.725
+ $X2=12.96 $Y2=1.65
r586 67 69 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.96 $Y=1.725
+ $X2=12.96 $Y2=2.465
r587 66 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.605 $Y=1.65
+ $X2=12.53 $Y2=1.65
r588 65 112 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.885 $Y=1.65
+ $X2=12.96 $Y2=1.65
r589 65 66 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.885 $Y=1.65
+ $X2=12.605 $Y2=1.65
r590 62 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.53 $Y=1.725
+ $X2=12.53 $Y2=1.65
r591 62 64 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.53 $Y=1.725
+ $X2=12.53 $Y2=2.465
r592 61 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.175 $Y=1.65
+ $X2=12.1 $Y2=1.65
r593 60 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.455 $Y=1.65
+ $X2=12.53 $Y2=1.65
r594 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.455 $Y=1.65
+ $X2=12.175 $Y2=1.65
r595 57 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.1 $Y=1.725
+ $X2=12.1 $Y2=1.65
r596 57 59 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.1 $Y=1.725
+ $X2=12.1 $Y2=2.465
r597 56 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.745 $Y=1.65
+ $X2=11.67 $Y2=1.65
r598 55 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.025 $Y=1.65
+ $X2=12.1 $Y2=1.65
r599 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.025 $Y=1.65
+ $X2=11.745 $Y2=1.65
r600 52 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.67 $Y=1.725
+ $X2=11.67 $Y2=1.65
r601 52 54 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=11.67 $Y=1.725
+ $X2=11.67 $Y2=2.465
r602 51 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.315 $Y=1.65
+ $X2=11.24 $Y2=1.65
r603 50 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.595 $Y=1.65
+ $X2=11.67 $Y2=1.65
r604 50 51 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=11.595 $Y=1.65
+ $X2=11.315 $Y2=1.65
r605 47 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.24 $Y=1.725
+ $X2=11.24 $Y2=1.65
r606 47 49 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=11.24 $Y=1.725
+ $X2=11.24 $Y2=2.465
r607 46 107 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.885 $Y=1.65
+ $X2=10.81 $Y2=1.65
r608 45 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.165 $Y=1.65
+ $X2=11.24 $Y2=1.65
r609 45 46 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=11.165 $Y=1.65
+ $X2=10.885 $Y2=1.65
r610 42 107 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.81 $Y=1.725
+ $X2=10.81 $Y2=1.65
r611 42 44 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=10.81 $Y=1.725
+ $X2=10.81 $Y2=2.465
r612 41 106 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.455 $Y=1.65
+ $X2=10.38 $Y2=1.65
r613 40 107 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.735 $Y=1.65
+ $X2=10.81 $Y2=1.65
r614 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.735 $Y=1.65
+ $X2=10.455 $Y2=1.65
r615 37 106 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.38 $Y=1.725
+ $X2=10.38 $Y2=1.65
r616 37 39 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=10.38 $Y=1.725
+ $X2=10.38 $Y2=2.465
r617 36 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.025 $Y=1.65
+ $X2=9.95 $Y2=1.65
r618 35 106 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.305 $Y=1.65
+ $X2=10.38 $Y2=1.65
r619 35 36 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.305 $Y=1.65
+ $X2=10.025 $Y2=1.65
r620 32 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.95 $Y=1.725
+ $X2=9.95 $Y2=1.65
r621 32 34 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.95 $Y=1.725
+ $X2=9.95 $Y2=2.465
r622 31 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.595 $Y=1.65
+ $X2=9.52 $Y2=1.65
r623 30 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.875 $Y=1.65
+ $X2=9.95 $Y2=1.65
r624 30 31 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.875 $Y=1.65
+ $X2=9.595 $Y2=1.65
r625 27 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.52 $Y=1.725
+ $X2=9.52 $Y2=1.65
r626 27 29 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.52 $Y=1.725
+ $X2=9.52 $Y2=2.465
r627 25 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.445 $Y=1.65
+ $X2=9.52 $Y2=1.65
r628 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.445 $Y=1.65
+ $X2=9.165 $Y2=1.65
r629 22 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.09 $Y=1.725
+ $X2=9.165 $Y2=1.65
r630 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.09 $Y=1.725
+ $X2=9.09 $Y2=2.465
r631 20 171 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.38 $Y=2.675
+ $X2=2.38 $Y2=1.905
r632 16 170 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.34 $Y=1.325
+ $X2=2.34 $Y2=1.575
r633 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.265 $Y=1.25
+ $X2=2.34 $Y2=1.325
r634 14 15 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.265 $Y=1.25
+ $X2=1.905 $Y2=1.25
r635 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.83 $Y=1.175
+ $X2=1.905 $Y2=1.25
r636 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.83 $Y=1.175
+ $X2=1.83 $Y2=0.635
r637 3 128 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=7.72
+ $Y=1.835 $X2=7.86 $Y2=2.9
r638 3 126 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.72
+ $Y=1.835 $X2=7.86 $Y2=1.98
r639 2 135 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.225 $Y2=2.105
r640 2 116 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.225 $Y2=2.9
r641 1 137 182 $w=1.7e-07 $l=6.81175e-07 $layer=licon1_NDIFF $count=1 $X=8.63
+ $Y=0.235 $X2=8.85 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A_381_85# 1 2 7 9 11 12 14 16 17
+ 20 24 26 27 28 29 33 35 37 38
c115 38 0 1.45114e-19 $X=2.965 $Y=1.65
c116 37 0 1.87795e-19 $X=2.965 $Y=1.575
c117 35 0 1.87887e-19 $X=2.965 $Y=1.74
c118 29 0 1.32904e-19 $X=2.33 $Y=2.17
c119 27 0 1.51585e-19 $X=2.245 $Y=1.285
c120 20 0 9.82022e-20 $X=2.16 $Y=0.78
c121 9 0 6.10011e-20 $X=3.675 $Y=1.725
r122 36 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.965 $Y=1.74
+ $X2=2.965 $Y2=1.65
r123 35 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=1.74
+ $X2=2.965 $Y2=1.575
r124 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.74 $X2=2.965 $Y2=1.74
r125 33 35 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.965 $Y=2.085
+ $X2=2.965 $Y2=1.74
r126 30 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.885 $Y=1.37
+ $X2=2.885 $Y2=1.575
r127 28 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.8 $Y=2.17
+ $X2=2.965 $Y2=2.085
r128 28 29 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.8 $Y=2.17
+ $X2=2.33 $Y2=2.17
r129 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.8 $Y=1.285
+ $X2=2.885 $Y2=1.37
r130 26 27 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.8 $Y=1.285
+ $X2=2.245 $Y2=1.285
r131 22 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.165 $Y=2.255
+ $X2=2.33 $Y2=2.17
r132 22 24 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.165 $Y=2.255
+ $X2=2.165 $Y2=2.4
r133 18 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.12 $Y=1.2
+ $X2=2.245 $Y2=1.285
r134 18 20 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=2.12 $Y=1.2 $X2=2.12
+ $Y2=0.78
r135 14 16 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.105 $Y=1.725
+ $X2=4.105 $Y2=2.465
r136 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.75 $Y=1.65
+ $X2=3.675 $Y2=1.65
r137 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.03 $Y=1.65
+ $X2=4.105 $Y2=1.725
r138 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.03 $Y=1.65
+ $X2=3.75 $Y2=1.65
r139 9 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.675 $Y=1.725
+ $X2=3.675 $Y2=1.65
r140 9 11 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.675 $Y=1.725
+ $X2=3.675 $Y2=2.465
r141 8 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.13 $Y=1.65
+ $X2=2.965 $Y2=1.65
r142 7 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.6 $Y=1.65
+ $X2=3.675 $Y2=1.65
r143 7 8 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.6 $Y=1.65 $X2=3.13
+ $Y2=1.65
r144 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=2.255 $X2=2.165 $Y2=2.4
r145 1 20 182 $w=1.7e-07 $l=4.65349e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.425 $X2=2.16 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A_726_47# 1 2 3 12 16 20 24 28 32
+ 34 36 37 39 40 42 43 45 46 47 48 50 51 53 55 56 58 60 61 63 65 66 68 70 71 73
+ 75 78 79 80 81 82 83 84 87 91 93 95 99 100 101 102 103 104 105 119 130 131 132
+ 135 140 145 150 155 176
c333 131 0 1.51162e-19 $X=6.675 $Y=1.16
c334 103 0 4.45833e-21 $X=9.6 $Y=1.295
c335 79 0 1.44143e-19 $X=6.675 $Y=1.665
r336 154 155 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.185
+ $Y=1.2 $X2=13.185 $Y2=1.2
r337 152 154 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=12.96 $Y=1.175
+ $X2=13.185 $Y2=1.175
r338 151 152 60.25 $w=3.44e-07 $l=4.3e-07 $layer=POLY_cond $X=12.53 $Y=1.175
+ $X2=12.96 $Y2=1.175
r339 149 151 28.7238 $w=3.44e-07 $l=2.05e-07 $layer=POLY_cond $X=12.325 $Y=1.175
+ $X2=12.53 $Y2=1.175
r340 149 150 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.325
+ $Y=1.2 $X2=12.325 $Y2=1.2
r341 147 149 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=12.1 $Y=1.175
+ $X2=12.325 $Y2=1.175
r342 144 145 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.445
+ $Y=1.2 $X2=11.445 $Y2=1.2
r343 139 140 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.605
+ $Y=1.2 $X2=10.605 $Y2=1.2
r344 134 135 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.745
+ $Y=1.2 $X2=9.745 $Y2=1.2
r345 132 134 97.9223 $w=3.3e-07 $l=5.6e-07 $layer=POLY_cond $X=10.305 $Y=1.2
+ $X2=9.745 $Y2=1.2
r346 130 131 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.675
+ $Y=1.16 $X2=6.675 $Y2=1.16
r347 128 131 3.48112 $w=6.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.48 $Y=1.33
+ $X2=6.675 $Y2=1.33
r348 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.295
+ $X2=6.48 $Y2=1.295
r349 124 176 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=5.535 $Y=1.295
+ $X2=5.535 $Y2=1.08
r350 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r351 119 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.185 $Y=1.295
+ $X2=13.185 $Y2=1.295
r352 116 119 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=12.325 $Y=1.295
+ $X2=13.185 $Y2=1.295
r353 116 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.325 $Y=1.295
+ $X2=12.325 $Y2=1.295
r354 113 116 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=11.465 $Y=1.295
+ $X2=12.325 $Y2=1.295
r355 113 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.465 $Y=1.295
+ $X2=11.465 $Y2=1.295
r356 110 113 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=10.605 $Y=1.295
+ $X2=11.465 $Y2=1.295
r357 110 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.605 $Y=1.295
+ $X2=10.605 $Y2=1.295
r358 107 110 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.745 $Y=1.295
+ $X2=10.605 $Y2=1.295
r359 107 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.745 $Y=1.295
+ $X2=9.745 $Y2=1.295
r360 105 107 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=9.715 $Y=1.295
+ $X2=9.745 $Y2=1.295
r361 104 127 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.295
+ $X2=6.48 $Y2=1.295
r362 103 105 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=9.6 $Y=1.295
+ $X2=9.715 $Y2=1.295
r363 103 104 3.68192 $w=1.4e-07 $l=2.975e-06 $layer=MET1_cond $X=9.6 $Y=1.295
+ $X2=6.625 $Y2=1.295
r364 102 123 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.295
+ $X2=5.52 $Y2=1.295
r365 101 127 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.295
+ $X2=6.48 $Y2=1.295
r366 101 102 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=6.335 $Y=1.295
+ $X2=5.665 $Y2=1.295
r367 96 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=1.08
+ $X2=3.77 $Y2=1.08
r368 96 98 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=3.855 $Y=1.08
+ $X2=5.08 $Y2=1.08
r369 95 176 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.435 $Y=1.08
+ $X2=5.535 $Y2=1.08
r370 95 98 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.435 $Y=1.08
+ $X2=5.08 $Y2=1.08
r371 91 100 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=3.83 $Y=1.96
+ $X2=3.83 $Y2=1.815
r372 91 93 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=3.83 $Y=1.96
+ $X2=3.83 $Y2=1.98
r373 89 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=1.165
+ $X2=3.77 $Y2=1.08
r374 89 100 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.77 $Y=1.165
+ $X2=3.77 $Y2=1.815
r375 85 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=0.995
+ $X2=3.77 $Y2=1.08
r376 85 87 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.77 $Y=0.995
+ $X2=3.77 $Y2=0.855
r377 78 130 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.675 $Y=1.5
+ $X2=6.675 $Y2=1.16
r378 78 79 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.675 $Y=1.5
+ $X2=6.675 $Y2=1.665
r379 77 130 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.675 $Y=0.995
+ $X2=6.675 $Y2=1.16
r380 73 75 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=15.97 $Y=0.985
+ $X2=15.97 $Y2=0.555
r381 72 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.615 $Y=1.06
+ $X2=15.54 $Y2=1.06
r382 71 73 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.895 $Y=1.06
+ $X2=15.97 $Y2=0.985
r383 71 72 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=15.895 $Y=1.06
+ $X2=15.615 $Y2=1.06
r384 68 84 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.54 $Y=0.985
+ $X2=15.54 $Y2=1.06
r385 68 70 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=15.54 $Y=0.985
+ $X2=15.54 $Y2=0.555
r386 67 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.185 $Y=1.06
+ $X2=15.11 $Y2=1.06
r387 66 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.465 $Y=1.06
+ $X2=15.54 $Y2=1.06
r388 66 67 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=15.465 $Y=1.06
+ $X2=15.185 $Y2=1.06
r389 63 83 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.11 $Y=0.985
+ $X2=15.11 $Y2=1.06
r390 63 65 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=15.11 $Y=0.985
+ $X2=15.11 $Y2=0.555
r391 62 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.755 $Y=1.06
+ $X2=14.68 $Y2=1.06
r392 61 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.035 $Y=1.06
+ $X2=15.11 $Y2=1.06
r393 61 62 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=15.035 $Y=1.06
+ $X2=14.755 $Y2=1.06
r394 58 82 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.68 $Y=0.985
+ $X2=14.68 $Y2=1.06
r395 58 60 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=14.68 $Y=0.985
+ $X2=14.68 $Y2=0.555
r396 57 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.325 $Y=1.06
+ $X2=14.25 $Y2=1.06
r397 56 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.605 $Y=1.06
+ $X2=14.68 $Y2=1.06
r398 56 57 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=14.605 $Y=1.06
+ $X2=14.325 $Y2=1.06
r399 53 81 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.25 $Y=0.985
+ $X2=14.25 $Y2=1.06
r400 53 55 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=14.25 $Y=0.985
+ $X2=14.25 $Y2=0.555
r401 52 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.895 $Y=1.06
+ $X2=13.82 $Y2=1.06
r402 51 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.175 $Y=1.06
+ $X2=14.25 $Y2=1.06
r403 51 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=14.175 $Y=1.06
+ $X2=13.895 $Y2=1.06
r404 48 80 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.82 $Y=0.985
+ $X2=13.82 $Y2=1.06
r405 48 50 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.82 $Y=0.985
+ $X2=13.82 $Y2=0.555
r406 46 80 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.745 $Y=1.06
+ $X2=13.82 $Y2=1.06
r407 46 47 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=13.745 $Y=1.06
+ $X2=13.465 $Y2=1.06
r408 43 47 26.108 $w=3.44e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.39 $Y=0.985
+ $X2=13.465 $Y2=1.06
r409 43 154 28.7238 $w=3.44e-07 $l=2.84561e-07 $layer=POLY_cond $X=13.39
+ $Y=0.985 $X2=13.185 $Y2=1.175
r410 43 45 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.39 $Y=0.985
+ $X2=13.39 $Y2=0.555
r411 40 152 22.2144 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=12.96 $Y=0.985
+ $X2=12.96 $Y2=1.175
r412 40 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.96 $Y=0.985
+ $X2=12.96 $Y2=0.555
r413 37 151 22.2144 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=12.53 $Y=0.985
+ $X2=12.53 $Y2=1.175
r414 37 39 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.53 $Y=0.985
+ $X2=12.53 $Y2=0.555
r415 34 147 22.2144 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=12.1 $Y=0.985
+ $X2=12.1 $Y2=1.175
r416 34 36 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.1 $Y=0.985
+ $X2=12.1 $Y2=0.555
r417 30 147 60.25 $w=3.44e-07 $l=4.3e-07 $layer=POLY_cond $X=11.67 $Y=1.175
+ $X2=12.1 $Y2=1.175
r418 30 144 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=11.67 $Y=1.175
+ $X2=11.445 $Y2=1.175
r419 30 32 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.67 $Y=1.035
+ $X2=11.67 $Y2=0.555
r420 26 144 28.7238 $w=3.44e-07 $l=2.05e-07 $layer=POLY_cond $X=11.24 $Y=1.175
+ $X2=11.445 $Y2=1.175
r421 26 28 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.24 $Y=1.035
+ $X2=11.24 $Y2=0.555
r422 22 26 60.25 $w=3.44e-07 $l=4.3e-07 $layer=POLY_cond $X=10.81 $Y=1.175
+ $X2=11.24 $Y2=1.175
r423 22 139 28.7238 $w=3.44e-07 $l=2.05e-07 $layer=POLY_cond $X=10.81 $Y=1.175
+ $X2=10.605 $Y2=1.175
r424 22 24 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.81 $Y=1.035
+ $X2=10.81 $Y2=0.555
r425 18 139 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=10.38 $Y=1.175
+ $X2=10.605 $Y2=1.175
r426 18 132 10.5087 $w=3.44e-07 $l=8.66025e-08 $layer=POLY_cond $X=10.38
+ $Y=1.175 $X2=10.305 $Y2=1.2
r427 18 20 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.38 $Y=1.035
+ $X2=10.38 $Y2=0.555
r428 16 79 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.615 $Y=2.285
+ $X2=6.615 $Y2=1.665
r429 12 77 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.615 $Y=0.445
+ $X2=6.615 $Y2=0.995
r430 3 93 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.75
+ $Y=1.835 $X2=3.89 $Y2=1.98
r431 2 98 182 $w=1.7e-07 $l=9.5751e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.235 $X2=5.08 $Y2=1.08
r432 1 87 182 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.235 $X2=3.77 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A 3 7 9 11 14 16 17 19 20 21 23 24
+ 25 28 30 32 33 37 39 41 42 43 44 45 54 65
c162 43 0 1.08533e-19 $X=8.06 $Y=1.65
c163 42 0 1.69365e-19 $X=7.63 $Y=1.65
c164 25 0 1.51162e-19 $X=7.2 $Y=1.65
c165 14 0 9.77732e-20 $X=5.395 $Y=0.655
r166 65 66 1.41962 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=5.09 $Y=1.665
+ $X2=5.09 $Y2=1.675
r167 53 55 46.7612 $w=2.68e-07 $l=2.6e-07 $layer=POLY_cond $X=5.135 $Y=1.53
+ $X2=5.395 $Y2=1.53
r168 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.135
+ $Y=1.51 $X2=5.135 $Y2=1.51
r169 51 53 16.1866 $w=2.68e-07 $l=9e-08 $layer=POLY_cond $X=5.045 $Y=1.53
+ $X2=5.135 $Y2=1.53
r170 44 65 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=5.09 $Y=1.627
+ $X2=5.09 $Y2=1.665
r171 44 54 4.08593 $w=3.28e-07 $l=1.17e-07 $layer=LI1_cond $X=5.09 $Y=1.627
+ $X2=5.09 $Y2=1.51
r172 44 45 16.1843 $w=2.28e-07 $l=3.23e-07 $layer=LI1_cond $X=5.04 $Y=1.712
+ $X2=5.04 $Y2=2.035
r173 44 66 1.85393 $w=2.28e-07 $l=3.7e-08 $layer=LI1_cond $X=5.04 $Y=1.712
+ $X2=5.04 $Y2=1.675
r174 39 43 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.075 $Y=1.725
+ $X2=8.06 $Y2=1.65
r175 39 41 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.075 $Y=1.725
+ $X2=8.075 $Y2=2.465
r176 35 43 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.045 $Y=1.575
+ $X2=8.06 $Y2=1.65
r177 35 37 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=8.045 $Y=1.575
+ $X2=8.045 $Y2=0.655
r178 34 42 12.05 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.72 $Y=1.65 $X2=7.63
+ $Y2=1.65
r179 33 43 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.97 $Y=1.65 $X2=8.06
+ $Y2=1.65
r180 33 34 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.97 $Y=1.65
+ $X2=7.72 $Y2=1.65
r181 30 42 12.05 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.645 $Y=1.725
+ $X2=7.63 $Y2=1.65
r182 30 32 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.645 $Y=1.725
+ $X2=7.645 $Y2=2.465
r183 26 42 12.05 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.615 $Y=1.575
+ $X2=7.63 $Y2=1.65
r184 26 28 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=7.615 $Y=1.575
+ $X2=7.615 $Y2=0.655
r185 24 42 12.05 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.54 $Y=1.65 $X2=7.63
+ $Y2=1.65
r186 24 25 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.54 $Y=1.65 $X2=7.2
+ $Y2=1.65
r187 22 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.125 $Y=1.725
+ $X2=7.2 $Y2=1.65
r188 22 23 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=7.125 $Y=1.725
+ $X2=7.125 $Y2=3.075
r189 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.05 $Y=3.15
+ $X2=7.125 $Y2=3.075
r190 20 21 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=7.05 $Y=3.15
+ $X2=5.79 $Y2=3.15
r191 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.715 $Y=3.075
+ $X2=5.79 $Y2=3.15
r192 18 19 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=5.715 $Y=1.715
+ $X2=5.715 $Y2=3.075
r193 17 55 22.7584 $w=2.68e-07 $l=1.42653e-07 $layer=POLY_cond $X=5.47 $Y=1.64
+ $X2=5.395 $Y2=1.53
r194 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.64 $Y=1.64
+ $X2=5.715 $Y2=1.715
r195 16 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.64 $Y=1.64
+ $X2=5.47 $Y2=1.64
r196 12 55 16.3317 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.395 $Y=1.345
+ $X2=5.395 $Y2=1.53
r197 12 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.395 $Y=1.345
+ $X2=5.395 $Y2=0.655
r198 9 51 16.3317 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.045 $Y=1.715
+ $X2=5.045 $Y2=1.53
r199 9 11 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.045 $Y=1.715 $X2=5.045
+ $Y2=2.465
r200 5 51 50.3582 $w=2.68e-07 $l=3.60832e-07 $layer=POLY_cond $X=4.765 $Y=1.345
+ $X2=5.045 $Y2=1.53
r201 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.765 $Y=1.345
+ $X2=4.765 $Y2=0.655
r202 1 5 26.9776 $w=2.68e-07 $l=2.12132e-07 $layer=POLY_cond $X=4.615 $Y=1.495
+ $X2=4.765 $Y2=1.345
r203 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=4.615 $Y=1.495
+ $X2=4.615 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A_1238_47# 1 2 9 10 12 14 17 19 20
+ 24 26 29 33 35 37 38 39
c126 29 0 3.37012e-20 $X=8.525 $Y=1.44
c127 26 0 3.19487e-19 $X=7.105 $Y=1.845
c128 20 0 9.77732e-20 $X=6.495 $Y=0.73
c129 12 0 7.99176e-20 $X=9.065 $Y=1.185
r130 38 39 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.525 $Y=1.26
+ $X2=8.525 $Y2=1.185
r131 33 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.83 $Y=1.93
+ $X2=7.105 $Y2=1.93
r132 30 38 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.525 $Y=1.44
+ $X2=8.525 $Y2=1.26
r133 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.525
+ $Y=1.44 $X2=8.525 $Y2=1.44
r134 27 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.19 $Y=1.44
+ $X2=7.105 $Y2=1.44
r135 27 29 46.6216 $w=3.28e-07 $l=1.335e-06 $layer=LI1_cond $X=7.19 $Y=1.44
+ $X2=8.525 $Y2=1.44
r136 26 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.105 $Y=1.845
+ $X2=7.105 $Y2=1.93
r137 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.105 $Y=1.605
+ $X2=7.105 $Y2=1.44
r138 25 26 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.105 $Y=1.605
+ $X2=7.105 $Y2=1.845
r139 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.105 $Y=1.275
+ $X2=7.105 $Y2=1.44
r140 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.105 $Y=0.815
+ $X2=7.105 $Y2=1.275
r141 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.02 $Y=0.73
+ $X2=7.105 $Y2=0.815
r142 19 20 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.02 $Y=0.73
+ $X2=6.495 $Y2=0.73
r143 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.33 $Y=0.645
+ $X2=6.495 $Y2=0.73
r144 15 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=6.33 $Y=0.645
+ $X2=6.33 $Y2=0.47
r145 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.065 $Y=1.185
+ $X2=9.065 $Y2=0.655
r146 11 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.69 $Y=1.26
+ $X2=8.525 $Y2=1.26
r147 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.99 $Y=1.26
+ $X2=9.065 $Y2=1.185
r148 10 11 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=8.99 $Y=1.26 $X2=8.69
+ $Y2=1.26
r149 9 39 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.555 $Y=0.655
+ $X2=8.555 $Y2=1.185
r150 2 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.69
+ $Y=1.865 $X2=6.83 $Y2=2.01
r151 1 17 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=6.19
+ $Y=0.235 $X2=6.33 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13
+ 14 15 16 17 54 60 64 68 72 76 80 86 90 94 96 100 104 108 112 116 118 122 124
+ 126 129 130 132 133 135 136 138 139 140 141 143 144 146 147 149 150 151 152
+ 153 155 160 165 177 185 212 218 221 224 227 230 233 236 240
r274 239 240 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r275 236 237 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r276 233 234 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r277 230 231 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r278 227 228 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r279 224 225 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r280 221 222 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r281 218 219 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r282 216 240 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=3.33
+ $X2=17.52 $Y2=3.33
r283 216 237 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=3.33
+ $X2=16.56 $Y2=3.33
r284 215 216 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r285 213 236 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.7 $Y=3.33
+ $X2=16.615 $Y2=3.33
r286 213 215 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=16.7 $Y=3.33
+ $X2=17.04 $Y2=3.33
r287 212 239 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=17.39 $Y=3.33
+ $X2=17.575 $Y2=3.33
r288 212 215 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=17.39 $Y=3.33
+ $X2=17.04 $Y2=3.33
r289 211 237 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.56 $Y2=3.33
r290 210 211 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r291 208 211 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.6 $Y2=3.33
r292 207 208 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r293 205 208 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.64 $Y2=3.33
r294 204 205 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r295 202 205 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r296 202 234 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r297 201 202 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r298 199 233 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.4 $Y=3.33
+ $X2=12.315 $Y2=3.33
r299 199 201 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.4 $Y=3.33
+ $X2=12.72 $Y2=3.33
r300 198 234 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r301 197 198 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r302 195 198 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r303 194 195 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r304 192 195 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r305 191 192 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r306 189 230 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.875 $Y=3.33
+ $X2=8.54 $Y2=3.33
r307 189 191 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.875 $Y=3.33
+ $X2=9.36 $Y2=3.33
r308 188 231 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r309 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r310 185 230 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.205 $Y=3.33
+ $X2=8.54 $Y2=3.33
r311 185 187 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.205 $Y=3.33
+ $X2=7.92 $Y2=3.33
r312 184 188 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r313 184 228 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6 $Y2=3.33
r314 183 184 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r315 181 227 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.01 $Y2=3.33
r316 181 183 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.96 $Y2=3.33
r317 180 228 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r318 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r319 177 227 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6.01 $Y2=3.33
r320 177 179 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.52 $Y2=3.33
r321 176 180 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r322 175 176 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r323 173 176 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r324 173 225 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r325 172 175 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r326 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r327 170 224 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.76 $Y=3.33
+ $X2=2.635 $Y2=3.33
r328 170 172 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.76 $Y=3.33
+ $X2=3.12 $Y2=3.33
r329 169 225 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r330 169 222 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r331 168 169 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r332 166 221 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=1.695 $Y2=3.33
r333 166 168 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=2.16 $Y2=3.33
r334 165 224 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.51 $Y=3.33
+ $X2=2.635 $Y2=3.33
r335 165 168 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.51 $Y=3.33
+ $X2=2.16 $Y2=3.33
r336 164 222 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r337 164 219 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r338 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r339 161 218 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.88 $Y=3.33
+ $X2=0.755 $Y2=3.33
r340 161 163 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r341 160 221 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.695 $Y2=3.33
r342 160 163 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.2 $Y2=3.33
r343 158 219 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r344 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r345 155 218 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.63 $Y=3.33
+ $X2=0.755 $Y2=3.33
r346 155 157 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=3.33
+ $X2=0.24 $Y2=3.33
r347 153 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r348 153 231 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r349 151 210 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=15.67 $Y=3.33
+ $X2=15.6 $Y2=3.33
r350 151 152 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.67 $Y=3.33
+ $X2=15.755 $Y2=3.33
r351 149 207 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=14.81 $Y=3.33
+ $X2=14.64 $Y2=3.33
r352 149 150 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.81 $Y=3.33
+ $X2=14.895 $Y2=3.33
r353 148 210 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=14.98 $Y=3.33
+ $X2=15.6 $Y2=3.33
r354 148 150 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.98 $Y=3.33
+ $X2=14.895 $Y2=3.33
r355 146 204 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=13.95 $Y=3.33
+ $X2=13.68 $Y2=3.33
r356 146 147 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.95 $Y=3.33
+ $X2=14.035 $Y2=3.33
r357 145 207 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=14.12 $Y=3.33
+ $X2=14.64 $Y2=3.33
r358 145 147 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.12 $Y=3.33
+ $X2=14.035 $Y2=3.33
r359 143 201 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.09 $Y=3.33
+ $X2=12.72 $Y2=3.33
r360 143 144 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.09 $Y=3.33
+ $X2=13.175 $Y2=3.33
r361 142 204 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=13.26 $Y=3.33
+ $X2=13.68 $Y2=3.33
r362 142 144 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.26 $Y=3.33
+ $X2=13.175 $Y2=3.33
r363 140 197 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.28 $Y2=3.33
r364 140 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.455 $Y2=3.33
r365 138 194 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.51 $Y=3.33
+ $X2=10.32 $Y2=3.33
r366 138 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.51 $Y=3.33
+ $X2=10.595 $Y2=3.33
r367 137 197 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=10.68 $Y=3.33
+ $X2=11.28 $Y2=3.33
r368 137 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.68 $Y=3.33
+ $X2=10.595 $Y2=3.33
r369 135 191 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.57 $Y=3.33
+ $X2=9.36 $Y2=3.33
r370 135 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.57 $Y=3.33
+ $X2=9.695 $Y2=3.33
r371 134 194 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=9.82 $Y=3.33
+ $X2=10.32 $Y2=3.33
r372 134 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.82 $Y=3.33
+ $X2=9.695 $Y2=3.33
r373 132 183 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=6.96 $Y2=3.33
r374 132 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.39 $Y2=3.33
r375 131 187 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.92 $Y2=3.33
r376 131 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.39 $Y2=3.33
r377 129 175 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=4.56 $Y2=3.33
r378 129 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=4.83 $Y2=3.33
r379 128 179 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.995 $Y=3.33
+ $X2=5.52 $Y2=3.33
r380 128 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=3.33
+ $X2=4.83 $Y2=3.33
r381 124 239 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=17.515
+ $Y=3.245 $X2=17.575 $Y2=3.33
r382 124 126 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=17.515 $Y=3.245
+ $X2=17.515 $Y2=2.455
r383 120 236 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.615 $Y=3.245
+ $X2=16.615 $Y2=3.33
r384 120 122 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=16.615 $Y=3.245
+ $X2=16.615 $Y2=2.455
r385 119 152 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.84 $Y=3.33
+ $X2=15.755 $Y2=3.33
r386 118 236 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.53 $Y=3.33
+ $X2=16.615 $Y2=3.33
r387 118 119 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.53 $Y=3.33
+ $X2=15.84 $Y2=3.33
r388 114 152 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.755 $Y=3.245
+ $X2=15.755 $Y2=3.33
r389 114 116 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=15.755 $Y=3.245
+ $X2=15.755 $Y2=2.455
r390 110 150 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.895 $Y=3.245
+ $X2=14.895 $Y2=3.33
r391 110 112 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=14.895 $Y=3.245
+ $X2=14.895 $Y2=2.455
r392 106 147 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.035 $Y=3.245
+ $X2=14.035 $Y2=3.33
r393 106 108 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=14.035 $Y=3.245
+ $X2=14.035 $Y2=2.455
r394 102 144 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.175 $Y=3.245
+ $X2=13.175 $Y2=3.33
r395 102 104 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=13.175 $Y=3.245
+ $X2=13.175 $Y2=2.455
r396 98 233 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.315 $Y=3.245
+ $X2=12.315 $Y2=3.33
r397 98 100 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=12.315 $Y=3.245
+ $X2=12.315 $Y2=2.455
r398 97 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.54 $Y=3.33
+ $X2=11.455 $Y2=3.33
r399 96 233 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.23 $Y=3.33
+ $X2=12.315 $Y2=3.33
r400 96 97 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.23 $Y=3.33
+ $X2=11.54 $Y2=3.33
r401 92 141 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.455 $Y=3.245
+ $X2=11.455 $Y2=3.33
r402 92 94 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=11.455 $Y=3.245
+ $X2=11.455 $Y2=2.455
r403 88 139 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.595 $Y=3.245
+ $X2=10.595 $Y2=3.33
r404 88 90 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=10.595 $Y=3.245
+ $X2=10.595 $Y2=2.455
r405 84 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.695 $Y=3.245
+ $X2=9.695 $Y2=3.33
r406 84 86 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=9.695 $Y=3.245
+ $X2=9.695 $Y2=2.475
r407 80 83 12.1393 $w=6.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.54 $Y=2.27
+ $X2=8.54 $Y2=2.95
r408 78 230 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.54 $Y=3.245
+ $X2=8.54 $Y2=3.33
r409 78 83 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.54 $Y=3.245
+ $X2=8.54 $Y2=2.95
r410 74 133 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=3.33
r411 74 76 41.2575 $w=2.48e-07 $l=8.95e-07 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=2.35
r412 70 227 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r413 70 72 43.1293 $w=3.28e-07 $l=1.235e-06 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.01
r414 66 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=3.33
r415 66 68 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=2.895
r416 62 224 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=3.33
r417 62 64 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=2.6
r418 58 221 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=3.245
+ $X2=1.695 $Y2=3.33
r419 58 60 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.695 $Y=3.245
+ $X2=1.695 $Y2=2.455
r420 54 57 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=0.755 $Y=2.105
+ $X2=0.755 $Y2=2.95
r421 52 218 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=3.245
+ $X2=0.755 $Y2=3.33
r422 52 57 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.755 $Y=3.245
+ $X2=0.755 $Y2=2.95
r423 17 126 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=17.335
+ $Y=1.835 $X2=17.475 $Y2=2.455
r424 16 122 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=16.475
+ $Y=1.835 $X2=16.615 $Y2=2.455
r425 15 116 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=15.615
+ $Y=1.835 $X2=15.755 $Y2=2.455
r426 14 112 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=14.755
+ $Y=1.835 $X2=14.895 $Y2=2.455
r427 13 108 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=13.895
+ $Y=1.835 $X2=14.035 $Y2=2.455
r428 12 104 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=13.035
+ $Y=1.835 $X2=13.175 $Y2=2.455
r429 11 100 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=12.175
+ $Y=1.835 $X2=12.315 $Y2=2.455
r430 10 94 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=11.315
+ $Y=1.835 $X2=11.455 $Y2=2.455
r431 9 90 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=10.455
+ $Y=1.835 $X2=10.595 $Y2=2.455
r432 8 86 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=9.595
+ $Y=1.835 $X2=9.735 $Y2=2.475
r433 7 83 200 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=3 $X=8.15
+ $Y=1.835 $X2=8.37 $Y2=2.95
r434 7 80 200 $w=1.7e-07 $l=5.33784e-07 $layer=licon1_PDIFF $count=3 $X=8.15
+ $Y=1.835 $X2=8.37 $Y2=2.27
r435 6 76 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.285
+ $Y=1.835 $X2=7.43 $Y2=2.35
r436 5 72 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.865
+ $Y=1.865 $X2=6.01 $Y2=2.01
r437 4 68 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=4.69
+ $Y=1.835 $X2=4.83 $Y2=2.895
r438 3 64 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=2.455
+ $Y=2.255 $X2=2.595 $Y2=2.6
r439 2 60 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=1.835 $X2=1.655 $Y2=2.455
r440 1 57 600 $w=1.7e-07 $l=1.22916e-06 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.835 $X2=0.795 $Y2=2.95
r441 1 54 300 $w=1.7e-07 $l=3.71079e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.835 $X2=0.795 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A_658_367# 1 2 3 10 12 14 18 21 22
+ 26 33 35
c55 33 0 6.10011e-20 $X=4.32 $Y=2.44
r56 24 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.46 $Y=2.33 $X2=5.46
+ $Y2=2.415
r57 24 26 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=5.46 $Y=2.33
+ $X2=5.46 $Y2=2.02
r58 23 33 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=2.415
+ $X2=4.32 $Y2=2.415
r59 22 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.335 $Y=2.415
+ $X2=5.46 $Y2=2.415
r60 22 23 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=5.335 $Y=2.415
+ $X2=4.485 $Y2=2.415
r61 20 33 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.32 $Y=2.5 $X2=4.32
+ $Y2=2.415
r62 20 21 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.32 $Y=2.5
+ $X2=4.32 $Y2=2.895
r63 16 33 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.32 $Y=2.33 $X2=4.32
+ $Y2=2.415
r64 16 18 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.32 $Y=2.33
+ $X2=4.32 $Y2=1.98
r65 15 31 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=2.98
+ $X2=3.42 $Y2=2.98
r66 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.155 $Y=2.98
+ $X2=4.32 $Y2=2.895
r67 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.155 $Y=2.98
+ $X2=3.505 $Y2=2.98
r68 10 31 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.895
+ $X2=3.42 $Y2=2.98
r69 10 12 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.42 $Y=2.895
+ $X2=3.42 $Y2=1.98
r70 3 35 300 $w=1.7e-07 $l=7.60345e-07 $layer=licon1_PDIFF $count=2 $X=5.12
+ $Y=1.835 $X2=5.42 $Y2=2.46
r71 3 26 600 $w=1.7e-07 $l=3.81445e-07 $layer=licon1_PDIFF $count=1 $X=5.12
+ $Y=1.835 $X2=5.42 $Y2=2.02
r72 2 33 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=2.44
r73 2 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=1.98
r74 1 31 400 $w=1.7e-07 $l=1.12813e-06 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.835 $X2=3.42 $Y2=2.9
r75 1 12 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.835 $X2=3.42 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 55 57 59 63 67 69 72 82 92 102 112 122 132 142 143 154
r265 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.165 $Y=2.035
+ $X2=10.165 $Y2=2.035
r266 151 155 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.305 $Y=2.035
+ $X2=10.165 $Y2=2.035
r267 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.305 $Y=2.035
+ $X2=9.305 $Y2=2.035
r268 142 147 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=17.045 $Y=2.035
+ $X2=17.045 $Y2=2.9
r269 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.045 $Y=2.035
+ $X2=17.045 $Y2=2.035
r270 136 143 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=16.185 $Y=2.035
+ $X2=17.045 $Y2=2.035
r271 135 139 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=16.185 $Y=2.035
+ $X2=16.185 $Y2=2.9
r272 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.185 $Y=2.035
+ $X2=16.185 $Y2=2.035
r273 132 135 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=16.185 $Y=0.36
+ $X2=16.185 $Y2=2.035
r274 126 136 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=15.325 $Y=2.035
+ $X2=16.185 $Y2=2.035
r275 125 129 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=15.325 $Y=2.035
+ $X2=15.325 $Y2=2.9
r276 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.325 $Y=2.035
+ $X2=15.325 $Y2=2.035
r277 122 125 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=15.325 $Y=0.36
+ $X2=15.325 $Y2=2.035
r278 116 126 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=14.465 $Y=2.035
+ $X2=15.325 $Y2=2.035
r279 115 119 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=14.465 $Y=2.035
+ $X2=14.465 $Y2=2.9
r280 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.465 $Y=2.035
+ $X2=14.465 $Y2=2.035
r281 112 115 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=14.465 $Y=0.36
+ $X2=14.465 $Y2=2.035
r282 106 116 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=13.605 $Y=2.035
+ $X2=14.465 $Y2=2.035
r283 105 109 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=13.605 $Y=2.035
+ $X2=13.605 $Y2=2.9
r284 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.605 $Y=2.035
+ $X2=13.605 $Y2=2.035
r285 102 105 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=13.605 $Y=0.36
+ $X2=13.605 $Y2=2.035
r286 95 99 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=12.745 $Y=2.035
+ $X2=12.745 $Y2=2.9
r287 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.745 $Y=2.035
+ $X2=12.745 $Y2=2.035
r288 92 95 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=12.745 $Y=0.36
+ $X2=12.745 $Y2=2.035
r289 86 96 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=11.885 $Y=2.035
+ $X2=12.745 $Y2=2.035
r290 85 89 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=11.885 $Y=2.035
+ $X2=11.885 $Y2=2.9
r291 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.885 $Y=2.035
+ $X2=11.885 $Y2=2.035
r292 82 85 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=11.885 $Y=0.36
+ $X2=11.885 $Y2=2.035
r293 76 86 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=11.025 $Y=2.035
+ $X2=11.885 $Y2=2.035
r294 76 155 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=11.025 $Y=2.035
+ $X2=10.165 $Y2=2.035
r295 75 79 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=11.025 $Y=2.035
+ $X2=11.025 $Y2=2.9
r296 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.025 $Y=2.035
+ $X2=11.025 $Y2=2.035
r297 72 75 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=11.025 $Y=0.36
+ $X2=11.025 $Y2=2.035
r298 69 106 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=13.175 $Y=2.035
+ $X2=13.605 $Y2=2.035
r299 69 96 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=13.175 $Y=2.035
+ $X2=12.745 $Y2=2.035
r300 65 154 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=10.165 $Y=2.13
+ $X2=10.165 $Y2=2.04
r301 65 67 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=10.165 $Y=2.13
+ $X2=10.165 $Y2=2.9
r302 61 154 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=10.165 $Y=1.95
+ $X2=10.165 $Y2=2.04
r303 61 63 55.5268 $w=3.28e-07 $l=1.59e-06 $layer=LI1_cond $X=10.165 $Y=1.95
+ $X2=10.165 $Y2=0.36
r304 60 150 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=2.04
+ $X2=9.305 $Y2=2.04
r305 59 154 3.59259 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10 $Y=2.04
+ $X2=10.165 $Y2=2.04
r306 59 60 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=10 $Y=2.04 $X2=9.39
+ $Y2=2.04
r307 55 150 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.305 $Y=2.13
+ $X2=9.305 $Y2=2.04
r308 55 57 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=9.305 $Y=2.13
+ $X2=9.305 $Y2=2.9
r309 18 147 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=16.905
+ $Y=1.835 $X2=17.045 $Y2=2.9
r310 18 142 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=16.905
+ $Y=1.835 $X2=17.045 $Y2=2.105
r311 17 139 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=16.045
+ $Y=1.835 $X2=16.185 $Y2=2.9
r312 17 135 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=16.045
+ $Y=1.835 $X2=16.185 $Y2=2.105
r313 16 129 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=15.185
+ $Y=1.835 $X2=15.325 $Y2=2.9
r314 16 125 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=15.185
+ $Y=1.835 $X2=15.325 $Y2=2.105
r315 15 119 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=14.325
+ $Y=1.835 $X2=14.465 $Y2=2.9
r316 15 115 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=14.325
+ $Y=1.835 $X2=14.465 $Y2=2.105
r317 14 109 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.835 $X2=13.605 $Y2=2.9
r318 14 105 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.835 $X2=13.605 $Y2=2.105
r319 13 99 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=12.605
+ $Y=1.835 $X2=12.745 $Y2=2.9
r320 13 95 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=12.605
+ $Y=1.835 $X2=12.745 $Y2=2.105
r321 12 89 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=11.745
+ $Y=1.835 $X2=11.885 $Y2=2.9
r322 12 85 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=11.745
+ $Y=1.835 $X2=11.885 $Y2=2.105
r323 11 79 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=10.885
+ $Y=1.835 $X2=11.025 $Y2=2.9
r324 11 75 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=10.885
+ $Y=1.835 $X2=11.025 $Y2=2.105
r325 10 154 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=10.025
+ $Y=1.835 $X2=10.165 $Y2=2.105
r326 10 67 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=10.025
+ $Y=1.835 $X2=10.165 $Y2=2.9
r327 9 150 400 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.835 $X2=9.305 $Y2=2.125
r328 9 57 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.835 $X2=9.305 $Y2=2.9
r329 8 132 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=16.045
+ $Y=0.235 $X2=16.185 $Y2=0.36
r330 7 122 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=15.185
+ $Y=0.235 $X2=15.325 $Y2=0.36
r331 6 112 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.325
+ $Y=0.235 $X2=14.465 $Y2=0.36
r332 5 102 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=13.465
+ $Y=0.235 $X2=13.605 $Y2=0.36
r333 4 92 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=12.605
+ $Y=0.235 $X2=12.745 $Y2=0.36
r334 3 82 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=11.745
+ $Y=0.235 $X2=11.885 $Y2=0.36
r335 2 72 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=10.885
+ $Y=0.235 $X2=11.025 $Y2=0.36
r336 1 63 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=10.02
+ $Y=0.235 $X2=10.165 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13
+ 42 46 50 54 58 62 66 70 72 76 80 84 88 92 95 96 98 99 101 102 103 104 106 107
+ 109 110 112 113 115 116 117 119 124 132 144 172 173 176 179 182 185 188
r241 188 189 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r242 185 186 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r243 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r244 179 180 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r245 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r246 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r247 170 173 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=17.52 $Y2=0
r248 169 172 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=16.08 $Y=0
+ $X2=17.52 $Y2=0
r249 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r250 167 170 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.08 $Y2=0
r251 166 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r252 164 167 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.6 $Y2=0
r253 163 164 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r254 161 164 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.64 $Y2=0
r255 160 161 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r256 158 161 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r257 158 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r258 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r259 155 188 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.4 $Y=0
+ $X2=12.315 $Y2=0
r260 155 157 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.4 $Y=0
+ $X2=12.72 $Y2=0
r261 154 189 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r262 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r263 151 154 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r264 150 151 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r265 148 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.995 $Y=0
+ $X2=7.87 $Y2=0
r266 148 150 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=7.995 $Y=0
+ $X2=10.32 $Y2=0
r267 147 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r268 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r269 144 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.87 $Y2=0
r270 144 146 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r271 143 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r272 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r273 140 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.48 $Y2=0
r274 140 183 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=4.56 $Y2=0
r275 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r276 137 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.55 $Y2=0
r277 137 139 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=5.52 $Y2=0
r278 136 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r279 136 180 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=3.12 $Y2=0
r280 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r281 133 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=0
+ $X2=3.07 $Y2=0
r282 133 135 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.155 $Y=0
+ $X2=4.08 $Y2=0
r283 132 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=0
+ $X2=4.55 $Y2=0
r284 132 135 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.385 $Y=0
+ $X2=4.08 $Y2=0
r285 131 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r286 130 131 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r287 128 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.64 $Y2=0
r288 128 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=1.2 $Y2=0
r289 127 130 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r290 127 128 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r291 125 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0
+ $X2=1.225 $Y2=0
r292 125 127 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.39 $Y=0
+ $X2=1.68 $Y2=0
r293 124 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=3.07 $Y2=0
r294 124 130 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=2.64 $Y2=0
r295 122 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.2 $Y2=0
r296 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r297 119 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0
+ $X2=1.225 $Y2=0
r298 119 121 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=0
+ $X2=0.72 $Y2=0
r299 117 151 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r300 117 186 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=7.92 $Y2=0
r301 115 166 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=15.67 $Y=0 $X2=15.6
+ $Y2=0
r302 115 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.67 $Y=0
+ $X2=15.755 $Y2=0
r303 114 169 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=15.84 $Y=0
+ $X2=16.08 $Y2=0
r304 114 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.84 $Y=0
+ $X2=15.755 $Y2=0
r305 112 163 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=14.81 $Y=0
+ $X2=14.64 $Y2=0
r306 112 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.81 $Y=0
+ $X2=14.895 $Y2=0
r307 111 166 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=14.98 $Y=0
+ $X2=15.6 $Y2=0
r308 111 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.98 $Y=0
+ $X2=14.895 $Y2=0
r309 109 160 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=13.95 $Y=0
+ $X2=13.68 $Y2=0
r310 109 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.95 $Y=0
+ $X2=14.035 $Y2=0
r311 108 163 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=14.12 $Y=0
+ $X2=14.64 $Y2=0
r312 108 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.12 $Y=0
+ $X2=14.035 $Y2=0
r313 106 157 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.09 $Y=0
+ $X2=12.72 $Y2=0
r314 106 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.09 $Y=0
+ $X2=13.175 $Y2=0
r315 105 160 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=13.26 $Y=0
+ $X2=13.68 $Y2=0
r316 105 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.26 $Y=0
+ $X2=13.175 $Y2=0
r317 103 153 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=11.37 $Y=0
+ $X2=11.28 $Y2=0
r318 103 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.37 $Y=0
+ $X2=11.455 $Y2=0
r319 101 150 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.51 $Y=0
+ $X2=10.32 $Y2=0
r320 101 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.51 $Y=0
+ $X2=10.595 $Y2=0
r321 100 153 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=10.68 $Y=0
+ $X2=11.28 $Y2=0
r322 100 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.68 $Y=0
+ $X2=10.595 $Y2=0
r323 98 142 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.675 $Y=0
+ $X2=6.48 $Y2=0
r324 98 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.84
+ $Y2=0
r325 97 146 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.44 $Y2=0
r326 97 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=6.84
+ $Y2=0
r327 95 139 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.545 $Y=0
+ $X2=5.52 $Y2=0
r328 95 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.545 $Y=0 $X2=5.71
+ $Y2=0
r329 94 142 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.875 $Y=0
+ $X2=6.48 $Y2=0
r330 94 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=0 $X2=5.71
+ $Y2=0
r331 90 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.755 $Y=0.085
+ $X2=15.755 $Y2=0
r332 90 92 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.755 $Y=0.085
+ $X2=15.755 $Y2=0.36
r333 86 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.895 $Y=0.085
+ $X2=14.895 $Y2=0
r334 86 88 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=14.895 $Y=0.085
+ $X2=14.895 $Y2=0.36
r335 82 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.035 $Y=0.085
+ $X2=14.035 $Y2=0
r336 82 84 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=14.035 $Y=0.085
+ $X2=14.035 $Y2=0.36
r337 78 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.175 $Y=0.085
+ $X2=13.175 $Y2=0
r338 78 80 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.175 $Y=0.085
+ $X2=13.175 $Y2=0.36
r339 74 188 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.315 $Y=0.085
+ $X2=12.315 $Y2=0
r340 74 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.315 $Y=0.085
+ $X2=12.315 $Y2=0.36
r341 73 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.54 $Y=0
+ $X2=11.455 $Y2=0
r342 72 188 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.23 $Y=0
+ $X2=12.315 $Y2=0
r343 72 73 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.23 $Y=0 $X2=11.54
+ $Y2=0
r344 68 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.455 $Y=0.085
+ $X2=11.455 $Y2=0
r345 68 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.455 $Y=0.085
+ $X2=11.455 $Y2=0.36
r346 64 102 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.595 $Y=0.085
+ $X2=10.595 $Y2=0
r347 64 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=0.085
+ $X2=10.595 $Y2=0.36
r348 60 185 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0
r349 60 62 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0.48
r350 56 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0
r351 56 58 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0.38
r352 52 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=0.085
+ $X2=5.71 $Y2=0
r353 52 54 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.71 $Y=0.085
+ $X2=5.71 $Y2=0.3
r354 48 182 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=0.085
+ $X2=4.55 $Y2=0
r355 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.55 $Y=0.085
+ $X2=4.55 $Y2=0.38
r356 44 179 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0
r357 44 46 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.44
r358 40 176 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0
r359 40 42 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0.61
r360 13 92 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=15.615
+ $Y=0.235 $X2=15.755 $Y2=0.36
r361 12 88 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.755
+ $Y=0.235 $X2=14.895 $Y2=0.36
r362 11 84 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=13.895
+ $Y=0.235 $X2=14.035 $Y2=0.36
r363 10 80 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=13.035
+ $Y=0.235 $X2=13.175 $Y2=0.36
r364 9 76 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=12.175
+ $Y=0.235 $X2=12.315 $Y2=0.36
r365 8 70 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=11.315
+ $Y=0.235 $X2=11.455 $Y2=0.36
r366 7 66 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=10.455
+ $Y=0.235 $X2=10.595 $Y2=0.36
r367 6 62 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=7.69
+ $Y=0.235 $X2=7.83 $Y2=0.48
r368 5 58 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=6.69
+ $Y=0.235 $X2=6.84 $Y2=0.38
r369 4 54 182 $w=1.7e-07 $l=2.70555e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.235 $X2=5.71 $Y2=0.3
r370 3 50 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.55 $Y2=0.38
r371 2 46 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=2.925
+ $Y=0.235 $X2=3.07 $Y2=0.44
r372 1 42 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.425 $X2=1.225 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP_20%A_1451_47# 1 2 3 11 12 13 14 15 16
+ 21 27
c52 12 0 1.88451e-19 $X=8.175 $Y=1.01
r53 17 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.505 $Y=0.35
+ $X2=8.34 $Y2=0.35
r54 16 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.22 $Y=0.35
+ $X2=9.345 $Y2=0.35
r55 16 17 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.22 $Y=0.35
+ $X2=8.505 $Y2=0.35
r56 14 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.34 $Y=0.435 $X2=8.34
+ $Y2=0.35
r57 14 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=8.34 $Y=0.435
+ $X2=8.34 $Y2=0.925
r58 12 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.175 $Y=1.01
+ $X2=8.34 $Y2=0.925
r59 12 13 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.175 $Y=1.01
+ $X2=7.565 $Y2=1.01
r60 11 13 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=7.462 $Y=0.925
+ $X2=7.565 $Y2=1.01
r61 11 21 24.8869 $w=2.03e-07 $l=4.6e-07 $layer=LI1_cond $X=7.462 $Y=0.925
+ $X2=7.462 $Y2=0.465
r62 3 27 91 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=2 $X=9.14
+ $Y=0.235 $X2=9.305 $Y2=0.43
r63 2 25 91 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=2 $X=8.12
+ $Y=0.235 $X2=8.34 $Y2=0.43
r64 1 21 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=7.255
+ $Y=0.235 $X2=7.4 $Y2=0.38
.ends

