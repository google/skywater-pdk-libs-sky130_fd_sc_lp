# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand2b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.365000 0.495000 1.760000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.425000 5.180000 1.760000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.016000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.765000 3.080000 1.930000 ;
        RECT 1.435000 1.930000 4.515000 1.935000 ;
        RECT 1.435000 1.935000 1.695000 3.075000 ;
        RECT 1.475000 0.605000 1.805000 1.085000 ;
        RECT 1.475000 1.085000 2.805000 1.255000 ;
        RECT 2.365000 1.935000 4.515000 2.100000 ;
        RECT 2.365000 2.100000 3.690000 2.120000 ;
        RECT 2.365000 2.120000 2.665000 3.075000 ;
        RECT 2.475000 0.605000 2.805000 1.085000 ;
        RECT 2.620000 1.255000 2.805000 1.440000 ;
        RECT 2.620000 1.440000 3.080000 1.765000 ;
        RECT 3.360000 2.120000 3.690000 3.075000 ;
        RECT 4.295000 2.100000 4.515000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.095000  0.255000 0.345000 1.025000 ;
      RECT 0.095000  1.025000 0.835000 1.195000 ;
      RECT 0.095000  1.930000 0.835000 2.100000 ;
      RECT 0.095000  2.100000 0.355000 3.075000 ;
      RECT 0.525000  0.085000 0.855000 0.855000 ;
      RECT 0.525000  2.270000 1.265000 3.245000 ;
      RECT 0.665000  1.195000 0.835000 1.425000 ;
      RECT 0.665000  1.425000 2.450000 1.595000 ;
      RECT 0.665000  1.595000 0.835000 1.930000 ;
      RECT 1.005000  1.800000 1.265000 2.270000 ;
      RECT 1.045000  0.255000 3.165000 0.425000 ;
      RECT 1.045000  0.425000 1.305000 1.185000 ;
      RECT 1.865000  2.105000 2.195000 3.245000 ;
      RECT 1.975000  0.425000 2.305000 0.915000 ;
      RECT 2.835000  2.290000 3.165000 3.245000 ;
      RECT 2.975000  0.425000 3.165000 1.085000 ;
      RECT 2.975000  1.085000 4.955000 1.255000 ;
      RECT 3.335000  0.085000 3.665000 0.915000 ;
      RECT 3.835000  0.285000 4.025000 1.075000 ;
      RECT 3.835000  1.075000 4.955000 1.085000 ;
      RECT 3.860000  2.270000 4.125000 3.245000 ;
      RECT 4.195000  0.085000 4.525000 0.905000 ;
      RECT 4.685000  1.930000 5.015000 3.245000 ;
      RECT 4.695000  0.305000 4.955000 1.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_lp__nand2b_4
END LIBRARY
