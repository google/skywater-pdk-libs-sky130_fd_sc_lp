* File: sky130_fd_sc_lp__o2bb2ai_0.spice
* Created: Fri Aug 28 11:12:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2ai_0  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1003 A_117_56# N_A1_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_195_56#_M1000_d N_A2_N_M1000_g A_117_56# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_400_47#_M1009_d N_A_195_56#_M1009_g N_Y_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=11.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_B2_M1007_g N_A_400_47#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_400_47#_M1002_d N_B1_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_195_56#_M1005_d N_A1_N_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A2_N_M1001_g N_A_195_56#_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1006 N_Y_M1006_d N_A_195_56#_M1006_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1004 A_486_483# N_B2_M1004_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g A_486_483# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_83 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o2bb2ai_0.pxi.spice"
*
.ends
*
*
