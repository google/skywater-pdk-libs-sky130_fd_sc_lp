* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__einvp_4 A TE VGND VNB VPB VPWR Z
X0 a_301_367# a_35_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR a_35_47# a_301_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 Z A a_301_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_301_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR a_35_47# a_301_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_301_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_35_47# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_301_367# a_35_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_35_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Z A a_301_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
