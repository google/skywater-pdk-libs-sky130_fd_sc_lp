* File: sky130_fd_sc_lp__a221o_2.pex.spice
* Created: Fri Aug 28 09:52:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221O_2%A_86_27# 1 2 3 10 12 15 17 19 22 26 27 29 30
+ 33 36 37 38 41 48
c101 37 0 4.51811e-20 $X=3.31 $Y=1.165
r102 50 52 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.505 $Y=1.38
+ $X2=0.935 $Y2=1.38
r103 45 48 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.67 $Y=2.095
+ $X2=2.975 $Y2=2.095
r104 39 41 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=3.44 $Y=1.075
+ $X2=3.44 $Y2=0.42
r105 38 44 5.76111 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=1.165
+ $X2=2.67 $Y2=1.165
r106 37 39 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=3.31 $Y=1.165
+ $X2=3.44 $Y2=1.075
r107 37 38 34.197 $w=1.78e-07 $l=5.55e-07 $layer=LI1_cond $X=3.31 $Y=1.165
+ $X2=2.755 $Y2=1.165
r108 36 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=1.93
+ $X2=2.67 $Y2=2.095
r109 35 44 0.787725 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.67 $Y=1.255
+ $X2=2.67 $Y2=1.165
r110 35 36 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.67 $Y=1.255
+ $X2=2.67 $Y2=1.93
r111 31 44 27.6628 $w=1.72e-07 $l=3.9e-07 $layer=LI1_cond $X=2.28 $Y=1.165
+ $X2=2.67 $Y2=1.165
r112 31 33 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=2.28 $Y=1.075
+ $X2=2.28 $Y2=0.42
r113 29 31 11.7035 $w=1.72e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.115 $Y=1.16
+ $X2=2.28 $Y2=1.165
r114 29 30 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.115 $Y=1.16
+ $X2=1.235 $Y2=1.16
r115 27 52 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.07 $Y=1.38
+ $X2=0.935 $Y2=1.38
r116 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.38 $X2=1.07 $Y2=1.38
r117 24 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.11 $Y=1.245
+ $X2=1.235 $Y2=1.16
r118 24 26 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.11 $Y=1.245
+ $X2=1.11 $Y2=1.38
r119 20 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.545
+ $X2=0.935 $Y2=1.38
r120 20 22 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.935 $Y=1.545
+ $X2=0.935 $Y2=2.465
r121 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.215
+ $X2=0.935 $Y2=1.38
r122 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=1.215
+ $X2=0.935 $Y2=0.685
r123 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.545
+ $X2=0.505 $Y2=1.38
r124 13 15 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.505 $Y=1.545
+ $X2=0.505 $Y2=2.465
r125 10 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.215
+ $X2=0.505 $Y2=1.38
r126 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.505 $Y=1.215
+ $X2=0.505 $Y2=0.685
r127 3 48 600 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.835 $X2=2.975 $Y2=2.095
r128 2 41 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.265
+ $Y=0.245 $X2=3.405 $Y2=0.42
r129 1 33 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=2.14
+ $Y=0.265 $X2=2.28 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%A2 1 3 7 9 13
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.51 $X2=1.61 $Y2=1.51
r40 9 13 4.58022 $w=3.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.64 $Y=1.665
+ $X2=1.64 $Y2=1.51
r41 5 12 55.3704 $w=2.88e-07 $l=3.0801e-07 $layer=POLY_cond $X=1.705 $Y=1.245
+ $X2=1.612 $Y2=1.51
r42 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.705 $Y=1.245
+ $X2=1.705 $Y2=0.685
r43 1 12 38.6342 $w=2.88e-07 $l=1.73292e-07 $layer=POLY_cond $X=1.595 $Y=1.675
+ $X2=1.612 $Y2=1.51
r44 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.595 $Y=1.675
+ $X2=1.595 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%A1 3 7 9 10 17 18
r39 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.51 $X2=2.24 $Y2=1.51
r40 15 17 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.065 $Y=1.51
+ $X2=2.24 $Y2=1.51
r41 13 15 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.06 $Y=1.51
+ $X2=2.065 $Y2=1.51
r42 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.24 $Y=1.665
+ $X2=2.24 $Y2=2.035
r43 9 18 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.24 $Y=1.665
+ $X2=2.24 $Y2=1.51
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.345
+ $X2=2.065 $Y2=1.51
r45 5 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.065 $Y=1.345
+ $X2=2.065 $Y2=0.685
r46 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.675
+ $X2=2.06 $Y2=1.51
r47 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.06 $Y=1.675 $X2=2.06
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%C1 3 7 9 12 13
c32 13 0 1.41378e-19 $X=3.1 $Y=1.51
r33 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.51 $X2=3.1
+ $Y2=1.675
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.51 $X2=3.1
+ $Y2=1.345
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.51 $X2=3.1 $Y2=1.51
r36 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.1 $Y=1.665 $X2=3.1
+ $Y2=1.51
r37 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.19 $Y=2.465
+ $X2=3.19 $Y2=1.675
r38 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.19 $Y=0.665
+ $X2=3.19 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%B1 3 7 9 12 13
c36 7 0 1.41378e-19 $X=3.62 $Y=2.465
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.51
+ $X2=3.64 $Y2=1.675
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.51
+ $X2=3.64 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.64
+ $Y=1.51 $X2=3.64 $Y2=1.51
r40 9 13 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.62 $Y=1.665
+ $X2=3.62 $Y2=1.51
r41 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.62 $Y=2.465
+ $X2=3.62 $Y2=1.675
r42 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.62 $Y=0.665
+ $X2=3.62 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%B2 3 6 8 10 17 19
c28 17 0 4.51811e-20 $X=4.18 $Y=1.36
r29 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.18 $Y=1.36
+ $X2=4.18 $Y2=1.525
r30 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.18 $Y=1.36
+ $X2=4.18 $Y2=1.195
r31 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.18
+ $Y=1.36 $X2=4.18 $Y2=1.36
r32 10 18 8.41685 $w=5.38e-07 $l=3.8e-07 $layer=LI1_cond $X=4.56 $Y=1.48
+ $X2=4.18 $Y2=1.48
r33 8 18 2.21496 $w=5.38e-07 $l=1e-07 $layer=LI1_cond $X=4.08 $Y=1.48 $X2=4.18
+ $Y2=1.48
r34 6 20 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.09 $Y=2.465 $X2=4.09
+ $Y2=1.525
r35 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.09 $Y=0.665
+ $X2=4.09 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%VPWR 1 2 3 10 12 18 22 26 28 30 40 41 47 50
r57 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r62 38 41 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r63 37 40 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=3.33
+ $X2=2.275 $Y2=3.33
r66 35 37 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.44 $Y=3.33 $X2=2.64
+ $Y2=3.33
r67 34 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 34 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 31 44 4.43563 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r71 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 30 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.27 $Y2=3.33
r73 30 33 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 28 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r75 28 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 24 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=3.245
+ $X2=2.275 $Y2=3.33
r77 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.275 $Y=3.245
+ $X2=2.275 $Y2=2.95
r78 23 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.27 $Y2=3.33
r79 22 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=3.33
+ $X2=2.275 $Y2=3.33
r80 22 23 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.11 $Y=3.33
+ $X2=1.435 $Y2=3.33
r81 18 21 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=1.27 $Y=2.005
+ $X2=1.27 $Y2=2.95
r82 16 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=3.245
+ $X2=1.27 $Y2=3.33
r83 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.27 $Y=3.245
+ $X2=1.27 $Y2=2.95
r84 12 15 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=0.275 $Y=1.98
+ $X2=0.275 $Y2=2.95
r85 10 44 3.08204 $w=3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.212 $Y2=3.33
r86 10 15 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.95
r87 3 26 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=1.835 $X2=2.275 $Y2=2.95
r88 2 21 400 $w=1.7e-07 $l=1.23819e-06 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.835 $X2=1.27 $Y2=2.95
r89 2 18 400 $w=1.7e-07 $l=3.34365e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.835 $X2=1.27 $Y2=2.005
r90 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.95
r91 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%X 1 2 7 8 9 10 11 12 13 22
r18 13 40 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=0.705 $Y=2.775
+ $X2=0.705 $Y2=2.91
r19 12 13 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=2.405
+ $X2=0.705 $Y2=2.775
r20 11 12 22.2631 $w=2.18e-07 $l=4.25e-07 $layer=LI1_cond $X=0.705 $Y=1.98
+ $X2=0.705 $Y2=2.405
r21 10 11 16.5009 $w=2.18e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.98
r22 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.665
r23 8 9 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=0.925
+ $X2=0.705 $Y2=1.295
r24 7 8 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=0.555
+ $X2=0.705 $Y2=0.925
r25 7 22 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=0.705 $Y=0.555
+ $X2=0.705 $Y2=0.42
r26 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.91
r27 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=1.98
r28 1 22 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.265 $X2=0.72 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%A_334_367# 1 2 9 13 17 20
r33 15 17 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.835 $Y=2.43
+ $X2=3.835 $Y2=2.085
r34 14 20 3.15366 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.94 $Y=2.515
+ $X2=1.792 $Y2=2.515
r35 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.67 $Y=2.515
+ $X2=3.835 $Y2=2.43
r36 13 14 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=3.67 $Y=2.515
+ $X2=1.94 $Y2=2.515
r37 7 20 3.37808 $w=2.77e-07 $l=9.31128e-08 $layer=LI1_cond $X=1.775 $Y=2.43
+ $X2=1.792 $Y2=2.515
r38 7 9 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=1.775 $Y=2.43
+ $X2=1.775 $Y2=2.085
r39 2 17 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=3.695
+ $Y=1.835 $X2=3.835 $Y2=2.085
r40 1 20 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.67
+ $Y=1.835 $X2=1.81 $Y2=2.525
r41 1 9 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.835 $X2=1.81 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%A_653_367# 1 2 7 11 13
r16 11 16 3.43112 $w=3e-07 $l=1.52e-07 $layer=LI1_cond $X=4.32 $Y=2.77 $X2=4.32
+ $Y2=2.922
r17 11 13 26.3141 $w=2.98e-07 $l=6.85e-07 $layer=LI1_cond $X=4.32 $Y=2.77
+ $X2=4.32 $Y2=2.085
r18 7 16 3.38598 $w=3.05e-07 $l=1.5e-07 $layer=LI1_cond $X=4.17 $Y=2.922
+ $X2=4.32 $Y2=2.922
r19 7 9 28.9055 $w=3.03e-07 $l=7.65e-07 $layer=LI1_cond $X=4.17 $Y=2.922
+ $X2=3.405 $Y2=2.922
r20 2 16 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.165
+ $Y=1.835 $X2=4.305 $Y2=2.91
r21 2 13 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=4.165
+ $Y=1.835 $X2=4.305 $Y2=2.085
r22 1 9 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.835 $X2=3.405 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_2%VGND 1 2 3 4 13 15 19 23 27 30 31 32 34 39
+ 52 53 59 62
r59 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r60 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r62 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r63 50 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r64 50 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r65 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r66 47 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=2.975
+ $Y2=0
r67 47 49 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=4.08
+ $Y2=0
r68 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r69 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r70 43 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r71 42 45 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r72 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r73 40 59 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.32
+ $Y2=0
r74 40 42 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.68
+ $Y2=0
r75 39 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.975
+ $Y2=0
r76 39 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.64
+ $Y2=0
r77 38 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r78 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r79 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r80 35 56 4.43563 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r81 35 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r82 34 59 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.32
+ $Y2=0
r83 34 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r84 32 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r85 32 43 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r86 30 49 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.08
+ $Y2=0
r87 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.305
+ $Y2=0
r88 29 52 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.56
+ $Y2=0
r89 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.305
+ $Y2=0
r90 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=0.085
+ $X2=4.305 $Y2=0
r91 25 27 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.305 $Y=0.085
+ $X2=4.305 $Y2=0.39
r92 21 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=0.085
+ $X2=2.975 $Y2=0
r93 21 23 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.975 $Y=0.085
+ $X2=2.975 $Y2=0.39
r94 17 59 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=0.085
+ $X2=1.32 $Y2=0
r95 17 19 5.44483 $w=6.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.32 $Y=0.085
+ $X2=1.32 $Y2=0.39
r96 13 56 3.08204 $w=3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.212 $Y2=0
r97 13 15 12.4848 $w=2.98e-07 $l=3.25e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.41
r98 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.165
+ $Y=0.245 $X2=4.305 $Y2=0.39
r99 3 23 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.245 $X2=2.975 $Y2=0.39
r100 2 19 45.5 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=4 $X=1.01
+ $Y=0.265 $X2=1.49 $Y2=0.39
r101 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.265 $X2=0.29 $Y2=0.41
.ends

