# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux2_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__mux2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.935000 2.135000 1.185000 ;
        RECT 1.965000 1.185000 2.135000 1.550000 ;
        RECT 1.965000 1.550000 2.650000 2.005000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.360000 0.470000 2.735000 1.380000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.955000 0.785000 3.275000 1.850000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.255000 0.835000 1.095000 ;
        RECT 0.580000 1.095000 0.750000 1.850000 ;
        RECT 0.580000 1.850000 0.805000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.125000  0.085000 0.410000 1.095000 ;
      RECT 0.125000  1.815000 0.410000 3.245000 ;
      RECT 0.930000  1.275000 1.175000 1.605000 ;
      RECT 0.985000  2.855000 1.315000 3.245000 ;
      RECT 1.005000  0.595000 2.190000 0.765000 ;
      RECT 1.005000  0.765000 1.175000 1.275000 ;
      RECT 1.005000  1.605000 1.175000 2.515000 ;
      RECT 1.005000  2.515000 2.415000 2.685000 ;
      RECT 1.045000  0.085000 1.375000 0.425000 ;
      RECT 1.420000  1.395000 1.750000 2.175000 ;
      RECT 1.420000  2.175000 3.745000 2.345000 ;
      RECT 1.930000  0.255000 2.190000 0.595000 ;
      RECT 2.085000  2.685000 2.415000 2.845000 ;
      RECT 2.905000  0.085000 3.235000 0.615000 ;
      RECT 2.985000  2.515000 3.315000 3.245000 ;
      RECT 3.445000  0.275000 3.745000 2.175000 ;
      RECT 3.485000  2.345000 3.745000 2.895000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2_2
