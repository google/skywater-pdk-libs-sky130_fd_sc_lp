* File: sky130_fd_sc_lp__buflp_8.pxi.spice
* Created: Fri Aug 28 10:12:46 2020
* 
x_PM_SKY130_FD_SC_LP__BUFLP_8%A N_A_c_152_n N_A_M1003_g N_A_M1020_g N_A_c_154_n
+ N_A_M1006_g N_A_M1026_g N_A_M1041_g N_A_c_157_n N_A_M1008_g N_A_M1009_g
+ N_A_c_159_n N_A_M1000_g N_A_M1018_g N_A_c_161_n N_A_M1024_g N_A_M1042_g
+ N_A_c_163_n N_A_M1027_g A A A A N_A_c_165_n N_A_c_166_n A
+ PM_SKY130_FD_SC_LP__BUFLP_8%A
x_PM_SKY130_FD_SC_LP__BUFLP_8%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1006_s
+ N_A_27_47#_M1020_s N_A_27_47#_M1026_s N_A_27_47#_M1002_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1005_g N_A_27_47#_M1012_g N_A_27_47#_M1007_g N_A_27_47#_M1013_g
+ N_A_27_47#_M1014_g N_A_27_47#_M1019_g N_A_27_47#_M1021_g N_A_27_47#_M1022_g
+ N_A_27_47#_M1023_g N_A_27_47#_M1029_g N_A_27_47#_M1034_g N_A_27_47#_M1040_g
+ N_A_27_47#_M1004_g N_A_27_47#_M1010_g N_A_27_47#_M1011_g N_A_27_47#_M1017_g
+ N_A_27_47#_M1015_g N_A_27_47#_M1025_g N_A_27_47#_M1028_g N_A_27_47#_M1016_g
+ N_A_27_47#_M1031_g N_A_27_47#_M1030_g N_A_27_47#_M1033_g N_A_27_47#_M1032_g
+ N_A_27_47#_M1036_g N_A_27_47#_M1037_g N_A_27_47#_M1039_g N_A_27_47#_M1038_g
+ N_A_27_47#_M1043_g N_A_27_47#_M1035_g N_A_27_47#_c_304_n N_A_27_47#_c_326_n
+ N_A_27_47#_c_305_n N_A_27_47#_c_337_n N_A_27_47#_c_328_n N_A_27_47#_c_368_p
+ N_A_27_47#_c_329_n N_A_27_47#_c_306_n N_A_27_47#_c_307_n N_A_27_47#_c_308_n
+ N_A_27_47#_c_331_n N_A_27_47#_c_356_n N_A_27_47#_c_332_n N_A_27_47#_c_309_n
+ PM_SKY130_FD_SC_LP__BUFLP_8%A_27_47#
x_PM_SKY130_FD_SC_LP__BUFLP_8%A_114_367# N_A_114_367#_M1020_d
+ N_A_114_367#_M1041_d N_A_114_367#_M1018_s N_A_114_367#_c_665_n
+ N_A_114_367#_c_667_n N_A_114_367#_c_670_n N_A_114_367#_c_672_n
+ N_A_114_367#_c_674_n N_A_114_367#_c_678_n N_A_114_367#_c_680_n
+ N_A_114_367#_c_682_n PM_SKY130_FD_SC_LP__BUFLP_8%A_114_367#
x_PM_SKY130_FD_SC_LP__BUFLP_8%VPWR N_VPWR_M1009_d N_VPWR_M1042_d N_VPWR_M1005_d
+ N_VPWR_M1014_d N_VPWR_M1023_d N_VPWR_M1035_d N_VPWR_c_708_n N_VPWR_c_709_n
+ N_VPWR_c_710_n N_VPWR_c_711_n N_VPWR_c_712_n N_VPWR_c_713_n N_VPWR_c_714_n
+ N_VPWR_c_715_n N_VPWR_c_716_n N_VPWR_c_717_n N_VPWR_c_718_n N_VPWR_c_719_n
+ N_VPWR_c_720_n N_VPWR_c_721_n VPWR N_VPWR_c_722_n N_VPWR_c_723_n
+ N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_707_n PM_SKY130_FD_SC_LP__BUFLP_8%VPWR
x_PM_SKY130_FD_SC_LP__BUFLP_8%A_636_367# N_A_636_367#_M1002_s
+ N_A_636_367#_M1007_s N_A_636_367#_M1021_s N_A_636_367#_M1034_s
+ N_A_636_367#_M1011_d N_A_636_367#_M1016_d N_A_636_367#_M1032_d
+ N_A_636_367#_M1038_d N_A_636_367#_c_854_n N_A_636_367#_c_848_n
+ N_A_636_367#_c_849_n N_A_636_367#_c_868_n N_A_636_367#_c_850_n
+ N_A_636_367#_c_876_n N_A_636_367#_c_851_n N_A_636_367#_c_885_n
+ N_A_636_367#_c_887_n N_A_636_367#_c_891_n N_A_636_367#_c_893_n
+ N_A_636_367#_c_895_n N_A_636_367#_c_897_n N_A_636_367#_c_899_n
+ N_A_636_367#_c_901_n N_A_636_367#_c_903_n N_A_636_367#_c_969_p
+ N_A_636_367#_c_852_n N_A_636_367#_c_853_n N_A_636_367#_c_913_n
+ N_A_636_367#_c_914_n N_A_636_367#_c_915_n
+ PM_SKY130_FD_SC_LP__BUFLP_8%A_636_367#
x_PM_SKY130_FD_SC_LP__BUFLP_8%X N_X_M1010_s N_X_M1025_s N_X_M1031_s N_X_M1036_s
+ N_X_M1004_s N_X_M1015_s N_X_M1030_s N_X_M1037_s N_X_c_988_n N_X_c_1100_p
+ N_X_c_979_n N_X_c_980_n N_X_c_970_n N_X_c_971_n N_X_c_1005_n N_X_c_1007_n
+ N_X_c_972_n N_X_c_981_n N_X_c_1017_n N_X_c_973_n N_X_c_982_n N_X_c_1027_n
+ N_X_c_974_n N_X_c_983_n N_X_c_984_n N_X_c_975_n N_X_c_976_n N_X_c_985_n
+ N_X_c_977_n N_X_c_986_n X X PM_SKY130_FD_SC_LP__BUFLP_8%X
x_PM_SKY130_FD_SC_LP__BUFLP_8%A_114_47# N_A_114_47#_M1003_d N_A_114_47#_M1008_d
+ N_A_114_47#_M1024_d N_A_114_47#_c_1118_n N_A_114_47#_c_1143_p
+ N_A_114_47#_c_1120_n N_A_114_47#_c_1126_n N_A_114_47#_c_1128_n
+ N_A_114_47#_c_1131_n PM_SKY130_FD_SC_LP__BUFLP_8%A_114_47#
x_PM_SKY130_FD_SC_LP__BUFLP_8%VGND N_VGND_M1000_s N_VGND_M1027_s N_VGND_M1012_d
+ N_VGND_M1019_d N_VGND_M1029_d N_VGND_M1043_d N_VGND_c_1154_n N_VGND_c_1155_n
+ N_VGND_c_1156_n N_VGND_c_1157_n N_VGND_c_1158_n N_VGND_c_1159_n
+ N_VGND_c_1160_n N_VGND_c_1161_n N_VGND_c_1162_n N_VGND_c_1163_n
+ N_VGND_c_1164_n N_VGND_c_1165_n N_VGND_c_1166_n N_VGND_c_1167_n
+ N_VGND_c_1168_n VGND N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n
+ N_VGND_c_1172_n PM_SKY130_FD_SC_LP__BUFLP_8%VGND
x_PM_SKY130_FD_SC_LP__BUFLP_8%A_644_47# N_A_644_47#_M1001_s N_A_644_47#_M1013_s
+ N_A_644_47#_M1022_s N_A_644_47#_M1040_s N_A_644_47#_M1017_d
+ N_A_644_47#_M1028_d N_A_644_47#_M1033_d N_A_644_47#_M1039_d
+ N_A_644_47#_c_1304_n N_A_644_47#_c_1298_n N_A_644_47#_c_1299_n
+ N_A_644_47#_c_1312_n N_A_644_47#_c_1300_n N_A_644_47#_c_1318_n
+ N_A_644_47#_c_1301_n N_A_644_47#_c_1325_n N_A_644_47#_c_1327_n
+ N_A_644_47#_c_1331_n N_A_644_47#_c_1333_n N_A_644_47#_c_1335_n
+ N_A_644_47#_c_1337_n N_A_644_47#_c_1373_n N_A_644_47#_c_1302_n
+ N_A_644_47#_c_1303_n N_A_644_47#_c_1345_n N_A_644_47#_c_1349_n
+ N_A_644_47#_c_1351_n PM_SKY130_FD_SC_LP__BUFLP_8%A_644_47#
cc_1 VNB N_A_c_152_n 0.0192154f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_2 VNB N_A_M1020_g 0.00759806f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_A_c_154_n 0.0167424f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.185
cc_4 VNB N_A_M1026_g 0.00706305f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_5 VNB N_A_M1041_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_6 VNB N_A_c_157_n 0.0167469f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.185
cc_7 VNB N_A_M1009_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_8 VNB N_A_c_159_n 0.0159015f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.185
cc_9 VNB N_A_M1018_g 0.00706452f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_10 VNB N_A_c_161_n 0.0161347f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=1.185
cc_11 VNB N_A_M1042_g 0.00740668f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_12 VNB N_A_c_163_n 0.016367f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=1.185
cc_13 VNB A 0.00298504f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_14 VNB N_A_c_165_n 0.128247f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=1.35
cc_15 VNB N_A_c_166_n 0.0114419f $X=-0.19 $Y=-0.245 $X2=2.088 $Y2=1.347
cc_16 VNB N_A_27_47#_M1002_g 0.00314208f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.515
cc_17 VNB N_A_27_47#_M1001_g 0.0205385f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.185
cc_18 VNB N_A_27_47#_M1005_g 0.0029978f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_19 VNB N_A_27_47#_M1012_g 0.0198735f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.655
cc_20 VNB N_A_27_47#_M1007_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_21 VNB N_A_27_47#_M1013_g 0.0200684f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=0.655
cc_22 VNB N_A_27_47#_M1014_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_M1019_g 0.0212847f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_24 VNB N_A_27_47#_M1021_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_M1022_g 0.0215022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_M1023_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.35
cc_27 VNB N_A_27_47#_M1029_g 0.0198735f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.35
cc_28 VNB N_A_27_47#_M1034_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.35
cc_29 VNB N_A_27_47#_M1040_g 0.0200684f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.35
cc_30 VNB N_A_27_47#_M1004_g 0.00316367f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=1.35
cc_31 VNB N_A_27_47#_M1010_g 0.020168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_M1011_g 0.00332682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_M1017_g 0.0200726f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.347
cc_34 VNB N_A_27_47#_M1015_g 0.00332682f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.295
cc_35 VNB N_A_27_47#_M1025_g 0.0200726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_M1028_g 0.0209398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_M1016_g 0.00332682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_M1031_g 0.0218154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_M1030_g 0.00332682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_47#_M1033_g 0.0217951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_47#_M1032_g 0.00332682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_M1036_g 0.0218154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_M1037_g 0.00332682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_47#_M1039_g 0.0215119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_47#_M1038_g 0.00315587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_47#_M1043_g 0.024631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_47#_M1035_g 0.0036596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_47#_c_304_n 0.0215853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_47#_c_305_n 0.0254327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_47#_c_306_n 0.00686822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_27_47#_c_307_n 0.00319044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_47#_c_308_n 0.0115555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_27_47#_c_309_n 0.363003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VPWR_c_707_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_X_c_970_n 0.00324651f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=0.655
cc_56 VNB N_X_c_971_n 0.00137838f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.515
cc_57 VNB N_X_c_972_n 0.00312561f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_58 VNB N_X_c_973_n 0.00312561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_X_c_974_n 0.0104463f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.35
cc_60 VNB N_X_c_975_n 0.00176907f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_61 VNB N_X_c_976_n 0.00232363f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.35
cc_62 VNB N_X_c_977_n 0.00232363f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=1.35
cc_63 VNB X 0.0243502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1154_n 0.00238736f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.655
cc_65 VNB N_VGND_c_1155_n 0.00604227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1156_n 0.00171822f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.515
cc_67 VNB N_VGND_c_1157_n 0.0158404f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_68 VNB N_VGND_c_1158_n 0.00221438f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=0.655
cc_69 VNB N_VGND_c_1159_n 0.0171133f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_70 VNB N_VGND_c_1160_n 0.00231715f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=0.655
cc_71 VNB N_VGND_c_1161_n 0.011122f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_72 VNB N_VGND_c_1162_n 0.0229175f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_73 VNB N_VGND_c_1163_n 0.0478878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1164_n 0.00357001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1165_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1166_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_77 VNB N_VGND_c_1167_n 0.0158404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1168_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.35
cc_79 VNB N_VGND_c_1169_n 0.0995368f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=1.35
cc_80 VNB N_VGND_c_1170_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1171_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.347
cc_82 VNB N_VGND_c_1172_n 0.488968f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.347
cc_83 VNB N_A_644_47#_c_1298_n 0.00275044f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=1.515
cc_84 VNB N_A_644_47#_c_1299_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.465
cc_85 VNB N_A_644_47#_c_1300_n 0.00348765f $X=-0.19 $Y=-0.245 $X2=2.285
+ $Y2=0.655
cc_86 VNB N_A_644_47#_c_1301_n 0.00505471f $X=-0.19 $Y=-0.245 $X2=2.715
+ $Y2=0.655
cc_87 VNB N_A_644_47#_c_1302_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.35
cc_88 VNB N_A_644_47#_c_1303_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.35
cc_89 VPB N_A_M1020_g 0.0235442f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_90 VPB N_A_M1026_g 0.018509f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_91 VPB N_A_M1041_g 0.0185278f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_92 VPB N_A_M1009_g 0.0185278f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_93 VPB N_A_M1018_g 0.0185268f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_94 VPB N_A_M1042_g 0.0189936f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_95 VPB N_A_27_47#_M1002_g 0.0201436f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.515
cc_96 VPB N_A_27_47#_M1005_g 0.0191875f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_97 VPB N_A_27_47#_M1007_g 0.0191926f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_98 VPB N_A_27_47#_M1014_g 0.0191926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_27_47#_M1021_g 0.0191926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_27_47#_M1023_g 0.0191926f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.35
cc_101 VPB N_A_27_47#_M1034_g 0.0191926f $X=-0.19 $Y=1.655 $X2=1.72 $Y2=1.35
cc_102 VPB N_A_27_47#_M1004_g 0.0203231f $X=-0.19 $Y=1.655 $X2=2.4 $Y2=1.35
cc_103 VPB N_A_27_47#_M1011_g 0.0208763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_27_47#_M1015_g 0.0208806f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.295
cc_105 VPB N_A_27_47#_M1016_g 0.0208763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_27_47#_M1030_g 0.0208806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_27_47#_M1032_g 0.0208763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_27_47#_M1037_g 0.0208806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_27_47#_M1038_g 0.0200024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_27_47#_M1035_g 0.0232333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_326_n 0.0449052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_27_47#_c_305_n 0.00130682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_27_47#_c_328_n 0.00356615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_27_47#_c_329_n 0.00911742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_27_47#_c_306_n 0.00213042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_331_n 0.00875086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_332_n 0.00127131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_708_n 0.0047158f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.655
cc_119 VPB N_VPWR_c_709_n 0.00472864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_710_n 0.0047158f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_121 VPB N_VPWR_c_711_n 0.0185788f $X=-0.19 $Y=1.655 $X2=2.285 $Y2=0.655
cc_122 VPB N_VPWR_c_712_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_713_n 0.0047158f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_124 VPB N_VPWR_c_714_n 0.0116157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_715_n 0.0403716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_716_n 0.0490546f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.35
cc_127 VPB N_VPWR_c_717_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.35
cc_128 VPB N_VPWR_c_718_n 0.0185788f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=1.35
cc_129 VPB N_VPWR_c_719_n 0.00324402f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=1.35
cc_130 VPB N_VPWR_c_720_n 0.0195335f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=1.35
cc_131 VPB N_VPWR_c_721_n 0.00324402f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.35
cc_132 VPB N_VPWR_c_722_n 0.0185788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_723_n 0.102743f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.347
cc_134 VPB N_VPWR_c_724_n 0.00324402f $X=-0.19 $Y=1.655 $X2=2.4 $Y2=1.347
cc_135 VPB N_VPWR_c_725_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_707_n 0.0474947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_636_367#_c_848_n 0.00225436f $X=-0.19 $Y=1.655 $X2=2.215
+ $Y2=2.465
cc_138 VPB N_A_636_367#_c_849_n 0.00230427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_636_367#_c_850_n 0.00225436f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_636_367#_c_851_n 0.00455863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_636_367#_c_852_n 0.00230427f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.347
cc_142 VPB N_A_636_367#_c_853_n 0.00230427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_X_c_979_n 0.00307912f $X=-0.19 $Y=1.655 $X2=2.285 $Y2=1.185
cc_144 VPB N_X_c_980_n 0.00297779f $X=-0.19 $Y=1.655 $X2=2.285 $Y2=0.655
cc_145 VPB N_X_c_981_n 0.00307912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_X_c_982_n 0.00307912f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.35
cc_147 VPB N_X_c_983_n 0.0109427f $X=-0.19 $Y=1.655 $X2=1.72 $Y2=1.35
cc_148 VPB N_X_c_984_n 0.00231148f $X=-0.19 $Y=1.655 $X2=1.72 $Y2=1.35
cc_149 VPB N_X_c_985_n 0.00230209f $X=-0.19 $Y=1.655 $X2=2.4 $Y2=1.35
cc_150 VPB N_X_c_986_n 0.00230209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB X 0.00474806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 N_A_c_163_n N_A_27_47#_M1001_g 0.0216249f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_153 A N_A_27_47#_M1001_g 3.21428e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A_c_152_n N_A_27_47#_c_305_n 0.0199154f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_155 N_A_c_166_n N_A_27_47#_c_305_n 0.0265665f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_156 N_A_c_152_n N_A_27_47#_c_337_n 0.0113847f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A_c_154_n N_A_27_47#_c_337_n 0.0105208f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_158 N_A_c_165_n N_A_27_47#_c_337_n 6.95778e-19 $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_159 N_A_c_166_n N_A_27_47#_c_337_n 0.0328179f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_160 N_A_M1020_g N_A_27_47#_c_328_n 0.016986f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A_M1026_g N_A_27_47#_c_328_n 0.0140549f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_c_165_n N_A_27_47#_c_328_n 0.00224206f $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_163 N_A_c_166_n N_A_27_47#_c_328_n 0.0383999f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_164 N_A_M1041_g N_A_27_47#_c_329_n 0.0140243f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_M1009_g N_A_27_47#_c_329_n 0.0104915f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A_M1018_g N_A_27_47#_c_329_n 0.0104388f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_M1042_g N_A_27_47#_c_329_n 0.0165384f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_168 A N_A_27_47#_c_329_n 0.0354834f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_169 N_A_c_165_n N_A_27_47#_c_329_n 0.00863949f $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_170 N_A_c_166_n N_A_27_47#_c_329_n 0.0637422f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_171 N_A_M1042_g N_A_27_47#_c_306_n 0.00420569f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_172 A N_A_27_47#_c_306_n 0.0149286f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A_c_165_n N_A_27_47#_c_306_n 0.00244123f $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_174 N_A_c_152_n N_A_27_47#_c_308_n 7.92899e-19 $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A_c_157_n N_A_27_47#_c_356_n 0.005522f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_176 N_A_c_165_n N_A_27_47#_c_356_n 0.0012621f $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_177 N_A_c_166_n N_A_27_47#_c_356_n 0.0244274f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_178 N_A_c_165_n N_A_27_47#_c_332_n 0.00232957f $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_179 N_A_c_166_n N_A_27_47#_c_332_n 0.0143528f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_180 N_A_M1042_g N_A_27_47#_c_309_n 0.0230227f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_c_165_n N_A_27_47#_c_309_n 0.0137964f $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_182 N_A_M1020_g N_A_114_367#_c_665_n 0.00206773f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_M1026_g N_A_114_367#_c_665_n 5.89773e-19 $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_M1020_g N_A_114_367#_c_667_n 0.0101651f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_M1026_g N_A_114_367#_c_667_n 0.0108604f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_M1041_g N_A_114_367#_c_667_n 6.46727e-19 $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_M1026_g N_A_114_367#_c_670_n 0.0105205f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_M1041_g N_A_114_367#_c_670_n 0.0105205f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_M1041_g N_A_114_367#_c_672_n 0.0021125f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_M1009_g N_A_114_367#_c_672_n 7.32094e-19 $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_M1026_g N_A_114_367#_c_674_n 5.95697e-19 $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_A_M1041_g N_A_114_367#_c_674_n 0.00910881f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A_M1009_g N_A_114_367#_c_674_n 0.0104892f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_M1018_g N_A_114_367#_c_674_n 5.95697e-19 $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_M1009_g N_A_114_367#_c_678_n 0.01115f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_M1018_g N_A_114_367#_c_678_n 0.01115f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_M1018_g N_A_114_367#_c_680_n 7.32094e-19 $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_M1042_g N_A_114_367#_c_680_n 0.00212147f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_M1009_g N_A_114_367#_c_682_n 6.46727e-19 $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_M1018_g N_A_114_367#_c_682_n 0.0104833f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A_M1042_g N_A_114_367#_c_682_n 0.00932771f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_A_M1009_g N_VPWR_c_708_n 0.00284434f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A_M1018_g N_VPWR_c_708_n 0.00284434f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A_M1042_g N_VPWR_c_709_n 0.00276193f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A_M1020_g N_VPWR_c_716_n 0.00547432f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_M1026_g N_VPWR_c_716_n 0.00357842f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_M1041_g N_VPWR_c_716_n 0.00357842f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_M1009_g N_VPWR_c_716_n 0.00547432f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A_M1018_g N_VPWR_c_718_n 0.0054895f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A_M1042_g N_VPWR_c_718_n 0.0054895f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_M1020_g N_VPWR_c_707_n 0.0108268f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_M1026_g N_VPWR_c_707_n 0.00535118f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_M1041_g N_VPWR_c_707_n 0.00535118f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A_M1009_g N_VPWR_c_707_n 0.00975595f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_M1018_g N_VPWR_c_707_n 0.00979301f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_M1042_g N_VPWR_c_707_n 0.00988926f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_M1042_g N_A_636_367#_c_854_n 6.97104e-19 $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_218 N_A_M1042_g N_A_636_367#_c_849_n 3.84262e-19 $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_219 N_A_c_154_n N_A_114_47#_c_1118_n 0.00922208f $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_220 N_A_c_157_n N_A_114_47#_c_1118_n 0.0118963f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_221 N_A_c_159_n N_A_114_47#_c_1120_n 0.0113307f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_222 N_A_c_161_n N_A_114_47#_c_1120_n 0.0109736f $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_223 N_A_c_163_n N_A_114_47#_c_1120_n 0.00323025f $X=2.715 $Y=1.185 $X2=0
+ $Y2=0
cc_224 A N_A_114_47#_c_1120_n 0.0330373f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_225 N_A_c_165_n N_A_114_47#_c_1120_n 0.00150992f $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_226 N_A_c_166_n N_A_114_47#_c_1120_n 0.0236456f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_227 N_A_c_165_n N_A_114_47#_c_1126_n 7.75366e-19 $X=2.715 $Y=1.35 $X2=0 $Y2=0
cc_228 N_A_c_166_n N_A_114_47#_c_1126_n 0.0145739f $X=2.088 $Y=1.347 $X2=0 $Y2=0
cc_229 N_A_c_159_n N_A_114_47#_c_1128_n 4.5114e-19 $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_230 N_A_c_161_n N_A_114_47#_c_1128_n 0.00745542f $X=2.285 $Y=1.185 $X2=0
+ $Y2=0
cc_231 N_A_c_163_n N_A_114_47#_c_1128_n 0.00604218f $X=2.715 $Y=1.185 $X2=0
+ $Y2=0
cc_232 N_A_c_152_n N_A_114_47#_c_1131_n 0.00546947f $X=0.495 $Y=1.185 $X2=0
+ $Y2=0
cc_233 N_A_c_154_n N_A_114_47#_c_1131_n 0.00589857f $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_234 N_A_c_157_n N_A_114_47#_c_1131_n 8.27749e-19 $X=1.425 $Y=1.185 $X2=0
+ $Y2=0
cc_235 N_A_c_157_n N_VGND_c_1154_n 0.00107091f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_236 N_A_c_159_n N_VGND_c_1154_n 0.00882762f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_237 N_A_c_161_n N_VGND_c_1154_n 0.00286449f $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_238 N_A_c_163_n N_VGND_c_1155_n 0.00384911f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_239 N_A_c_152_n N_VGND_c_1163_n 0.0054895f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_240 N_A_c_154_n N_VGND_c_1163_n 0.00359361f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_241 N_A_c_157_n N_VGND_c_1163_n 0.00357877f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_242 N_A_c_159_n N_VGND_c_1163_n 0.00486043f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_243 N_A_c_161_n N_VGND_c_1165_n 0.0054895f $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_244 N_A_c_163_n N_VGND_c_1165_n 0.0054895f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_245 N_A_c_152_n N_VGND_c_1172_n 0.00722852f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_246 N_A_c_154_n N_VGND_c_1172_n 0.00559711f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_247 N_A_c_157_n N_VGND_c_1172_n 0.00553549f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_248 N_A_c_159_n N_VGND_c_1172_n 0.00440581f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_249 N_A_c_161_n N_VGND_c_1172_n 0.00599734f $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_250 N_A_c_163_n N_VGND_c_1172_n 0.00981835f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_328_n N_A_114_367#_M1020_d 0.00176461f $X=1.055 $Y=1.77
+ $X2=-0.19 $Y2=-0.245
cc_252 N_A_27_47#_c_329_n N_A_114_367#_M1041_d 0.00176461f $X=2.815 $Y=1.77
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_329_n N_A_114_367#_M1018_s 0.00176461f $X=2.815 $Y=1.77
+ $X2=0 $Y2=0
cc_254 N_A_27_47#_c_328_n N_A_114_367#_c_667_n 0.0170777f $X=1.055 $Y=1.77 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1026_s N_A_114_367#_c_670_n 0.00332344f $X=1 $Y=1.835 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_368_p N_A_114_367#_c_670_n 0.0126348f $X=1.14 $Y=1.98 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_329_n N_A_114_367#_c_672_n 0.01723f $X=2.815 $Y=1.77 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_329_n N_A_114_367#_c_678_n 0.0289344f $X=2.815 $Y=1.77 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_329_n N_A_114_367#_c_680_n 0.01723f $X=2.815 $Y=1.77 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_329_n N_VPWR_M1009_d 0.00176891f $X=2.815 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_261 N_A_27_47#_c_329_n N_VPWR_M1042_d 4.50532e-19 $X=2.815 $Y=1.77 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_306_n N_VPWR_M1042_d 0.00282238f $X=2.985 $Y=1.43 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1002_g N_VPWR_c_709_n 0.00620388f $X=3.105 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_329_n N_VPWR_c_709_n 0.00309162f $X=2.815 $Y=1.77 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_306_n N_VPWR_c_709_n 0.0114205f $X=2.985 $Y=1.43 $X2=0 $Y2=0
cc_266 N_A_27_47#_M1005_g N_VPWR_c_710_n 0.00271808f $X=3.535 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_M1007_g N_VPWR_c_710_n 0.00271808f $X=3.965 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1007_g N_VPWR_c_711_n 0.0054895f $X=3.965 $Y=2.465 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1014_g N_VPWR_c_711_n 0.0054895f $X=4.395 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1014_g N_VPWR_c_712_n 0.00271808f $X=4.395 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1021_g N_VPWR_c_712_n 0.00271808f $X=4.825 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1023_g N_VPWR_c_713_n 0.00271808f $X=5.255 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1034_g N_VPWR_c_713_n 0.00271808f $X=5.685 $Y=2.465 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1038_g N_VPWR_c_715_n 0.00109254f $X=9.615 $Y=2.465 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1035_g N_VPWR_c_715_n 0.0165757f $X=10.045 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_326_n N_VPWR_c_716_n 0.0174288f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_277 N_A_27_47#_M1002_g N_VPWR_c_720_n 0.0054895f $X=3.105 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1005_g N_VPWR_c_720_n 0.0054895f $X=3.535 $Y=2.465 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1021_g N_VPWR_c_722_n 0.0054895f $X=4.825 $Y=2.465 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1023_g N_VPWR_c_722_n 0.0054895f $X=5.255 $Y=2.465 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_M1034_g N_VPWR_c_723_n 0.00547432f $X=5.685 $Y=2.465 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1004_g N_VPWR_c_723_n 0.00357842f $X=6.115 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1011_g N_VPWR_c_723_n 0.00357877f $X=6.615 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_M1015_g N_VPWR_c_723_n 0.00357842f $X=7.115 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1016_g N_VPWR_c_723_n 0.00357877f $X=7.615 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1030_g N_VPWR_c_723_n 0.00357842f $X=8.115 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1032_g N_VPWR_c_723_n 0.00357877f $X=8.615 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1037_g N_VPWR_c_723_n 0.00357842f $X=9.115 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_M1038_g N_VPWR_c_723_n 0.00357877f $X=9.615 $Y=2.465 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1035_g N_VPWR_c_723_n 0.00486043f $X=10.045 $Y=2.465 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_M1020_s N_VPWR_c_707_n 0.00423245f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_M1026_s N_VPWR_c_707_n 0.00225186f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_293 N_A_27_47#_M1002_g N_VPWR_c_707_n 0.00997125f $X=3.105 $Y=2.465 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1005_g N_VPWR_c_707_n 0.00979301f $X=3.535 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1007_g N_VPWR_c_707_n 0.00979301f $X=3.965 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_M1014_g N_VPWR_c_707_n 0.00979301f $X=4.395 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_M1021_g N_VPWR_c_707_n 0.00979301f $X=4.825 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1023_g N_VPWR_c_707_n 0.00979301f $X=5.255 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1034_g N_VPWR_c_707_n 0.00975595f $X=5.685 $Y=2.465 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_M1004_g N_VPWR_c_707_n 0.00553547f $X=6.115 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1011_g N_VPWR_c_707_n 0.0057905f $X=6.615 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1015_g N_VPWR_c_707_n 0.00570659f $X=7.115 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_M1016_g N_VPWR_c_707_n 0.0057905f $X=7.615 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_M1030_g N_VPWR_c_707_n 0.00570659f $X=8.115 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_M1032_g N_VPWR_c_707_n 0.0057905f $X=8.615 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1037_g N_VPWR_c_707_n 0.00570659f $X=9.115 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_M1038_g N_VPWR_c_707_n 0.00553549f $X=9.615 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_M1035_g N_VPWR_c_707_n 0.00824727f $X=10.045 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_326_n N_VPWR_c_707_n 0.00963639f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_310 N_A_27_47#_M1002_g N_A_636_367#_c_854_n 0.0153072f $X=3.105 $Y=2.465
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_M1005_g N_A_636_367#_c_854_n 0.014976f $X=3.535 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_M1007_g N_A_636_367#_c_854_n 7.24315e-19 $X=3.965 $Y=2.465
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_M1005_g N_A_636_367#_c_848_n 0.01115f $X=3.535 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_M1007_g N_A_636_367#_c_848_n 0.01115f $X=3.965 $Y=2.465 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_307_n N_A_636_367#_c_848_n 0.0388321f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_309_n N_A_636_367#_c_848_n 0.00239965f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_M1002_g N_A_636_367#_c_849_n 0.00372308f $X=3.105 $Y=2.465
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_M1005_g N_A_636_367#_c_849_n 0.00157732f $X=3.535 $Y=2.465
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_306_n N_A_636_367#_c_849_n 0.00639807f $X=2.985 $Y=1.43
+ $X2=0 $Y2=0
cc_320 N_A_27_47#_c_307_n N_A_636_367#_c_849_n 0.0276081f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_309_n N_A_636_367#_c_849_n 0.00248733f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_M1005_g N_A_636_367#_c_868_n 7.24315e-19 $X=3.535 $Y=2.465
+ $X2=0 $Y2=0
cc_323 N_A_27_47#_M1007_g N_A_636_367#_c_868_n 0.014976f $X=3.965 $Y=2.465 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1014_g N_A_636_367#_c_868_n 0.014976f $X=4.395 $Y=2.465 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1021_g N_A_636_367#_c_868_n 7.24315e-19 $X=4.825 $Y=2.465
+ $X2=0 $Y2=0
cc_326 N_A_27_47#_M1014_g N_A_636_367#_c_850_n 0.01115f $X=4.395 $Y=2.465 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_M1021_g N_A_636_367#_c_850_n 0.01115f $X=4.825 $Y=2.465 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_307_n N_A_636_367#_c_850_n 0.0388321f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_309_n N_A_636_367#_c_850_n 0.00239965f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_M1014_g N_A_636_367#_c_876_n 7.24315e-19 $X=4.395 $Y=2.465
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_M1021_g N_A_636_367#_c_876_n 0.014976f $X=4.825 $Y=2.465 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_M1023_g N_A_636_367#_c_876_n 0.014976f $X=5.255 $Y=2.465 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_M1034_g N_A_636_367#_c_876_n 7.24315e-19 $X=5.685 $Y=2.465
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_M1023_g N_A_636_367#_c_851_n 0.01115f $X=5.255 $Y=2.465 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_M1034_g N_A_636_367#_c_851_n 0.0127273f $X=5.685 $Y=2.465
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_M1004_g N_A_636_367#_c_851_n 0.0029339f $X=6.115 $Y=2.465
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_307_n N_A_636_367#_c_851_n 0.0664403f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_309_n N_A_636_367#_c_851_n 0.00536003f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_M1034_g N_A_636_367#_c_885_n 0.00197018f $X=5.685 $Y=2.465
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_M1004_g N_A_636_367#_c_885_n 5.89773e-19 $X=6.115 $Y=2.465
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_M1023_g N_A_636_367#_c_887_n 6.73286e-19 $X=5.255 $Y=2.465
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_M1034_g N_A_636_367#_c_887_n 0.0130117f $X=5.685 $Y=2.465
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_M1004_g N_A_636_367#_c_887_n 0.0133459f $X=6.115 $Y=2.465
+ $X2=0 $Y2=0
cc_344 N_A_27_47#_M1011_g N_A_636_367#_c_887_n 7.43959e-19 $X=6.615 $Y=2.465
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_M1004_g N_A_636_367#_c_891_n 0.0109138f $X=6.115 $Y=2.465
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_M1011_g N_A_636_367#_c_891_n 0.0143648f $X=6.615 $Y=2.465
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_M1015_g N_A_636_367#_c_893_n 0.0131712f $X=7.115 $Y=2.465
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_M1016_g N_A_636_367#_c_893_n 7.04111e-19 $X=7.615 $Y=2.465
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_M1015_g N_A_636_367#_c_895_n 0.0109138f $X=7.115 $Y=2.465
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_M1016_g N_A_636_367#_c_895_n 0.0143648f $X=7.615 $Y=2.465
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_M1030_g N_A_636_367#_c_897_n 0.0131712f $X=8.115 $Y=2.465
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_M1032_g N_A_636_367#_c_897_n 7.04111e-19 $X=8.615 $Y=2.465
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_M1030_g N_A_636_367#_c_899_n 0.0109138f $X=8.115 $Y=2.465
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_M1032_g N_A_636_367#_c_899_n 0.0143648f $X=8.615 $Y=2.465
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_M1037_g N_A_636_367#_c_901_n 0.0130573f $X=9.115 $Y=2.465
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_M1038_g N_A_636_367#_c_901_n 9.72084e-19 $X=9.615 $Y=2.465
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_M1037_g N_A_636_367#_c_903_n 0.0109138f $X=9.115 $Y=2.465
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_M1038_g N_A_636_367#_c_903_n 0.0118963f $X=9.615 $Y=2.465
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_M1007_g N_A_636_367#_c_852_n 0.00157732f $X=3.965 $Y=2.465
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_M1014_g N_A_636_367#_c_852_n 0.00157732f $X=4.395 $Y=2.465
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_307_n N_A_636_367#_c_852_n 0.0276081f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_309_n N_A_636_367#_c_852_n 0.00248733f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_M1021_g N_A_636_367#_c_853_n 0.00157732f $X=4.825 $Y=2.465
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_M1023_g N_A_636_367#_c_853_n 0.00157732f $X=5.255 $Y=2.465
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_307_n N_A_636_367#_c_853_n 0.0276081f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_309_n N_A_636_367#_c_853_n 0.00272398f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_M1015_g N_A_636_367#_c_913_n 5.89773e-19 $X=7.115 $Y=2.465
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_M1030_g N_A_636_367#_c_914_n 5.89773e-19 $X=8.115 $Y=2.465
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_M1037_g N_A_636_367#_c_915_n 5.89773e-19 $X=9.115 $Y=2.465
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_M1011_g N_X_c_988_n 0.0125612f $X=6.615 $Y=2.465 $X2=0 $Y2=0
cc_371 N_A_27_47#_M1015_g N_X_c_988_n 7.27325e-19 $X=7.115 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A_27_47#_M1011_g N_X_c_979_n 0.0115433f $X=6.615 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A_27_47#_M1015_g N_X_c_979_n 0.0151263f $X=7.115 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A_27_47#_c_307_n N_X_c_979_n 0.0492574f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_375 N_A_27_47#_c_309_n N_X_c_979_n 0.00416609f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_376 N_A_27_47#_M1004_g N_X_c_980_n 0.00115862f $X=6.115 $Y=2.465 $X2=0 $Y2=0
cc_377 N_A_27_47#_M1011_g N_X_c_980_n 0.00158254f $X=6.615 $Y=2.465 $X2=0 $Y2=0
cc_378 N_A_27_47#_c_307_n N_X_c_980_n 0.02772f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_379 N_A_27_47#_c_309_n N_X_c_980_n 0.00459133f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_380 N_A_27_47#_M1017_g N_X_c_970_n 0.0103102f $X=6.705 $Y=0.655 $X2=0 $Y2=0
cc_381 N_A_27_47#_M1025_g N_X_c_970_n 0.0104187f $X=7.135 $Y=0.655 $X2=0 $Y2=0
cc_382 N_A_27_47#_c_307_n N_X_c_970_n 0.0506643f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_309_n N_X_c_970_n 0.00232085f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_384 N_A_27_47#_M1010_g N_X_c_971_n 3.08854e-19 $X=6.275 $Y=0.655 $X2=0 $Y2=0
cc_385 N_A_27_47#_c_307_n N_X_c_971_n 0.013984f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_386 N_A_27_47#_c_309_n N_X_c_971_n 0.00266022f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_387 N_A_27_47#_M1016_g N_X_c_1005_n 0.0125612f $X=7.615 $Y=2.465 $X2=0 $Y2=0
cc_388 N_A_27_47#_M1030_g N_X_c_1005_n 7.27325e-19 $X=8.115 $Y=2.465 $X2=0 $Y2=0
cc_389 N_A_27_47#_M1028_g N_X_c_1007_n 0.00585188f $X=7.565 $Y=0.655 $X2=0 $Y2=0
cc_390 N_A_27_47#_M1031_g N_X_c_1007_n 5.88195e-19 $X=8.065 $Y=0.655 $X2=0 $Y2=0
cc_391 N_A_27_47#_M1028_g N_X_c_972_n 0.00906883f $X=7.565 $Y=0.655 $X2=0 $Y2=0
cc_392 N_A_27_47#_M1031_g N_X_c_972_n 0.0112452f $X=8.065 $Y=0.655 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_307_n N_X_c_972_n 0.0492951f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_309_n N_X_c_972_n 0.00400849f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_395 N_A_27_47#_M1016_g N_X_c_981_n 0.0115433f $X=7.615 $Y=2.465 $X2=0 $Y2=0
cc_396 N_A_27_47#_M1030_g N_X_c_981_n 0.0150578f $X=8.115 $Y=2.465 $X2=0 $Y2=0
cc_397 N_A_27_47#_c_307_n N_X_c_981_n 0.0492574f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_398 N_A_27_47#_c_309_n N_X_c_981_n 0.00400849f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_399 N_A_27_47#_M1032_g N_X_c_1017_n 0.0125612f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A_27_47#_M1037_g N_X_c_1017_n 7.27325e-19 $X=9.115 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A_27_47#_M1033_g N_X_c_973_n 0.00962761f $X=8.565 $Y=0.655 $X2=0 $Y2=0
cc_402 N_A_27_47#_M1036_g N_X_c_973_n 0.0112452f $X=9.065 $Y=0.655 $X2=0 $Y2=0
cc_403 N_A_27_47#_c_307_n N_X_c_973_n 0.049329f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_404 N_A_27_47#_c_309_n N_X_c_973_n 0.00400849f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_405 N_A_27_47#_M1032_g N_X_c_982_n 0.0115433f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_406 N_A_27_47#_M1037_g N_X_c_982_n 0.0150578f $X=9.115 $Y=2.465 $X2=0 $Y2=0
cc_407 N_A_27_47#_c_307_n N_X_c_982_n 0.0492574f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_408 N_A_27_47#_c_309_n N_X_c_982_n 0.00400849f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_409 N_A_27_47#_M1038_g N_X_c_1027_n 0.0123462f $X=9.615 $Y=2.465 $X2=0 $Y2=0
cc_410 N_A_27_47#_M1035_g N_X_c_1027_n 9.49435e-19 $X=10.045 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_M1039_g N_X_c_974_n 0.00958336f $X=9.565 $Y=0.655 $X2=0 $Y2=0
cc_412 N_A_27_47#_M1043_g N_X_c_974_n 0.0161614f $X=10.045 $Y=0.655 $X2=0 $Y2=0
cc_413 N_A_27_47#_c_307_n N_X_c_974_n 0.0224562f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_414 N_A_27_47#_c_309_n N_X_c_974_n 0.00385554f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_415 N_A_27_47#_M1038_g N_X_c_983_n 0.01115f $X=9.615 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A_27_47#_M1035_g N_X_c_983_n 0.0151297f $X=10.045 $Y=2.465 $X2=0 $Y2=0
cc_417 N_A_27_47#_c_307_n N_X_c_983_n 0.0186645f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_418 N_A_27_47#_c_309_n N_X_c_983_n 0.00253752f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_419 N_A_27_47#_M1016_g N_X_c_984_n 0.00173883f $X=7.615 $Y=2.465 $X2=0 $Y2=0
cc_420 N_A_27_47#_c_307_n N_X_c_984_n 0.02772f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_421 N_A_27_47#_c_309_n N_X_c_984_n 0.00423635f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_422 N_A_27_47#_M1028_g N_X_c_975_n 0.00138961f $X=7.565 $Y=0.655 $X2=0 $Y2=0
cc_423 N_A_27_47#_c_307_n N_X_c_975_n 0.0204548f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_424 N_A_27_47#_c_309_n N_X_c_975_n 0.00230524f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_425 N_A_27_47#_M1031_g N_X_c_976_n 4.44647e-19 $X=8.065 $Y=0.655 $X2=0 $Y2=0
cc_426 N_A_27_47#_M1033_g N_X_c_976_n 0.00792922f $X=8.565 $Y=0.655 $X2=0 $Y2=0
cc_427 N_A_27_47#_M1036_g N_X_c_976_n 6.69159e-19 $X=9.065 $Y=0.655 $X2=0 $Y2=0
cc_428 N_A_27_47#_c_307_n N_X_c_976_n 0.026869f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_429 N_A_27_47#_c_309_n N_X_c_976_n 0.00411613f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_430 N_A_27_47#_M1032_g N_X_c_985_n 0.00173883f $X=8.615 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A_27_47#_c_307_n N_X_c_985_n 0.02772f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_309_n N_X_c_985_n 0.00415747f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_433 N_A_27_47#_M1036_g N_X_c_977_n 4.44647e-19 $X=9.065 $Y=0.655 $X2=0 $Y2=0
cc_434 N_A_27_47#_M1039_g N_X_c_977_n 0.00777721f $X=9.565 $Y=0.655 $X2=0 $Y2=0
cc_435 N_A_27_47#_M1043_g N_X_c_977_n 9.35553e-19 $X=10.045 $Y=0.655 $X2=0 $Y2=0
cc_436 N_A_27_47#_c_307_n N_X_c_977_n 0.026869f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_437 N_A_27_47#_c_309_n N_X_c_977_n 0.00411613f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_438 N_A_27_47#_M1038_g N_X_c_986_n 0.00173883f $X=9.615 $Y=2.465 $X2=0 $Y2=0
cc_439 N_A_27_47#_c_307_n N_X_c_986_n 0.02772f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_440 N_A_27_47#_c_309_n N_X_c_986_n 0.00415747f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_441 N_A_27_47#_M1039_g X 9.64082e-19 $X=9.565 $Y=0.655 $X2=0 $Y2=0
cc_442 N_A_27_47#_M1038_g X 9.96541e-19 $X=9.615 $Y=2.465 $X2=0 $Y2=0
cc_443 N_A_27_47#_M1043_g X 0.00796462f $X=10.045 $Y=0.655 $X2=0 $Y2=0
cc_444 N_A_27_47#_M1035_g X 0.00785246f $X=10.045 $Y=2.465 $X2=0 $Y2=0
cc_445 N_A_27_47#_c_307_n X 0.0261204f $X=9.655 $Y=1.43 $X2=0 $Y2=0
cc_446 N_A_27_47#_c_309_n X 0.0153009f $X=10.045 $Y=1.43 $X2=0 $Y2=0
cc_447 N_A_27_47#_c_337_n N_A_114_47#_M1003_d 0.00328233f $X=1.045 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_448 N_A_27_47#_M1006_s N_A_114_47#_c_1118_n 0.00472489f $X=1 $Y=0.235 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_337_n N_A_114_47#_c_1118_n 0.00352531f $X=1.045 $Y=0.925
+ $X2=0 $Y2=0
cc_450 N_A_27_47#_c_356_n N_A_114_47#_c_1118_n 0.018913f $X=1.21 $Y=0.765 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_329_n N_A_114_47#_c_1120_n 0.00170365f $X=2.815 $Y=1.77
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_c_337_n N_A_114_47#_c_1131_n 0.0160355f $X=1.045 $Y=0.925
+ $X2=0 $Y2=0
cc_453 N_A_27_47#_M1001_g N_VGND_c_1155_n 0.00222426f $X=3.145 $Y=0.655 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_306_n N_VGND_c_1155_n 0.0127937f $X=2.985 $Y=1.43 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_307_n N_VGND_c_1155_n 0.00256539f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_M1001_g N_VGND_c_1156_n 6.79703e-19 $X=3.145 $Y=0.655 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_M1012_g N_VGND_c_1156_n 0.0105033f $X=3.575 $Y=0.655 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_M1013_g N_VGND_c_1156_n 0.00199874f $X=4.005 $Y=0.655 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_M1013_g N_VGND_c_1157_n 0.0054895f $X=4.005 $Y=0.655 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_M1019_g N_VGND_c_1157_n 0.00486043f $X=4.435 $Y=0.655 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_M1013_g N_VGND_c_1158_n 6.85661e-19 $X=4.005 $Y=0.655 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_M1019_g N_VGND_c_1158_n 0.01152f $X=4.435 $Y=0.655 $X2=0 $Y2=0
cc_463 N_A_27_47#_M1022_g N_VGND_c_1158_n 0.00629085f $X=4.985 $Y=0.655 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_M1022_g N_VGND_c_1159_n 0.0054895f $X=4.985 $Y=0.655 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_M1029_g N_VGND_c_1159_n 0.00486043f $X=5.415 $Y=0.655 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_M1022_g N_VGND_c_1160_n 6.94749e-19 $X=4.985 $Y=0.655 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_M1029_g N_VGND_c_1160_n 0.0105873f $X=5.415 $Y=0.655 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_M1040_g N_VGND_c_1160_n 0.00336952f $X=5.845 $Y=0.655 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_M1039_g N_VGND_c_1162_n 0.00108379f $X=9.565 $Y=0.655 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_M1043_g N_VGND_c_1162_n 0.0126962f $X=10.045 $Y=0.655 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_304_n N_VGND_c_1163_n 0.0174288f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_472 N_A_27_47#_M1001_g N_VGND_c_1167_n 0.0054895f $X=3.145 $Y=0.655 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_M1012_g N_VGND_c_1167_n 0.00486043f $X=3.575 $Y=0.655 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_M1040_g N_VGND_c_1169_n 0.00547432f $X=5.845 $Y=0.655 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_M1010_g N_VGND_c_1169_n 0.00357842f $X=6.275 $Y=0.655 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_M1017_g N_VGND_c_1169_n 0.00359361f $X=6.705 $Y=0.655 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_M1025_g N_VGND_c_1169_n 0.00359361f $X=7.135 $Y=0.655 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_M1028_g N_VGND_c_1169_n 0.00357877f $X=7.565 $Y=0.655 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_M1031_g N_VGND_c_1169_n 0.00359361f $X=8.065 $Y=0.655 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_M1033_g N_VGND_c_1169_n 0.00357877f $X=8.565 $Y=0.655 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_M1036_g N_VGND_c_1169_n 0.00359361f $X=9.065 $Y=0.655 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_M1039_g N_VGND_c_1169_n 0.00357877f $X=9.565 $Y=0.655 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_M1043_g N_VGND_c_1169_n 0.00564095f $X=10.045 $Y=0.655 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_M1003_s N_VGND_c_1172_n 0.00266928f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_M1006_s N_VGND_c_1172_n 0.00280678f $X=1 $Y=0.235 $X2=0 $Y2=0
cc_486 N_A_27_47#_M1001_g N_VGND_c_1172_n 0.00981835f $X=3.145 $Y=0.655 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_M1012_g N_VGND_c_1172_n 0.00824727f $X=3.575 $Y=0.655 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_M1013_g N_VGND_c_1172_n 0.00990036f $X=4.005 $Y=0.655 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_M1019_g N_VGND_c_1172_n 0.00824727f $X=4.435 $Y=0.655 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_M1022_g N_VGND_c_1172_n 0.0103112f $X=4.985 $Y=0.655 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_M1029_g N_VGND_c_1172_n 0.00824727f $X=5.415 $Y=0.655 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_M1040_g N_VGND_c_1172_n 0.0098633f $X=5.845 $Y=0.655 $X2=0
+ $Y2=0
cc_493 N_A_27_47#_M1010_g N_VGND_c_1172_n 0.00535118f $X=6.275 $Y=0.655 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_M1017_g N_VGND_c_1172_n 0.00541283f $X=6.705 $Y=0.655 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_M1025_g N_VGND_c_1172_n 0.00541283f $X=7.135 $Y=0.655 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_M1028_g N_VGND_c_1172_n 0.00560622f $X=7.565 $Y=0.655 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_M1031_g N_VGND_c_1172_n 0.0057814f $X=8.065 $Y=0.655 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_M1033_g N_VGND_c_1172_n 0.0057905f $X=8.565 $Y=0.655 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_M1036_g N_VGND_c_1172_n 0.0057814f $X=9.065 $Y=0.655 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_M1039_g N_VGND_c_1172_n 0.00574036f $X=9.565 $Y=0.655 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_M1043_g N_VGND_c_1172_n 0.00972484f $X=10.045 $Y=0.655 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_c_304_n N_VGND_c_1172_n 0.00963639f $X=0.28 $Y=0.42 $X2=0
+ $Y2=0
cc_503 N_A_27_47#_c_337_n N_VGND_c_1172_n 0.0062047f $X=1.045 $Y=0.925 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_M1001_g N_A_644_47#_c_1304_n 0.00820863f $X=3.145 $Y=0.655
+ $X2=0 $Y2=0
cc_505 N_A_27_47#_M1012_g N_A_644_47#_c_1298_n 0.0124899f $X=3.575 $Y=0.655
+ $X2=0 $Y2=0
cc_506 N_A_27_47#_M1013_g N_A_644_47#_c_1298_n 0.01115f $X=4.005 $Y=0.655 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_307_n N_A_644_47#_c_1298_n 0.0447482f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_309_n N_A_644_47#_c_1298_n 0.00239965f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_509 N_A_27_47#_M1001_g N_A_644_47#_c_1299_n 0.00235582f $X=3.145 $Y=0.655
+ $X2=0 $Y2=0
cc_510 N_A_27_47#_c_307_n N_A_644_47#_c_1299_n 0.0209731f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_c_309_n N_A_644_47#_c_1299_n 0.00248733f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_512 N_A_27_47#_M1012_g N_A_644_47#_c_1312_n 7.17209e-19 $X=3.575 $Y=0.655
+ $X2=0 $Y2=0
cc_513 N_A_27_47#_M1013_g N_A_644_47#_c_1312_n 0.00962188f $X=4.005 $Y=0.655
+ $X2=0 $Y2=0
cc_514 N_A_27_47#_M1019_g N_A_644_47#_c_1300_n 0.0131221f $X=4.435 $Y=0.655
+ $X2=0 $Y2=0
cc_515 N_A_27_47#_M1022_g N_A_644_47#_c_1300_n 0.0117822f $X=4.985 $Y=0.655
+ $X2=0 $Y2=0
cc_516 N_A_27_47#_c_307_n N_A_644_47#_c_1300_n 0.053767f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_309_n N_A_644_47#_c_1300_n 0.00556291f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_518 N_A_27_47#_M1019_g N_A_644_47#_c_1318_n 9.68862e-19 $X=4.435 $Y=0.655
+ $X2=0 $Y2=0
cc_519 N_A_27_47#_M1022_g N_A_644_47#_c_1318_n 0.0103283f $X=4.985 $Y=0.655
+ $X2=0 $Y2=0
cc_520 N_A_27_47#_M1029_g N_A_644_47#_c_1301_n 0.0124899f $X=5.415 $Y=0.655
+ $X2=0 $Y2=0
cc_521 N_A_27_47#_M1040_g N_A_644_47#_c_1301_n 0.0121254f $X=5.845 $Y=0.655
+ $X2=0 $Y2=0
cc_522 N_A_27_47#_M1010_g N_A_644_47#_c_1301_n 0.00233572f $X=6.275 $Y=0.655
+ $X2=0 $Y2=0
cc_523 N_A_27_47#_c_307_n N_A_644_47#_c_1301_n 0.0723563f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_524 N_A_27_47#_c_309_n N_A_644_47#_c_1301_n 0.00536003f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_525 N_A_27_47#_M1040_g N_A_644_47#_c_1325_n 0.00197018f $X=5.845 $Y=0.655
+ $X2=0 $Y2=0
cc_526 N_A_27_47#_M1010_g N_A_644_47#_c_1325_n 5.89773e-19 $X=6.275 $Y=0.655
+ $X2=0 $Y2=0
cc_527 N_A_27_47#_M1029_g N_A_644_47#_c_1327_n 6.48194e-19 $X=5.415 $Y=0.655
+ $X2=0 $Y2=0
cc_528 N_A_27_47#_M1040_g N_A_644_47#_c_1327_n 0.00800443f $X=5.845 $Y=0.655
+ $X2=0 $Y2=0
cc_529 N_A_27_47#_M1010_g N_A_644_47#_c_1327_n 0.00779336f $X=6.275 $Y=0.655
+ $X2=0 $Y2=0
cc_530 N_A_27_47#_M1017_g N_A_644_47#_c_1327_n 5.97847e-19 $X=6.705 $Y=0.655
+ $X2=0 $Y2=0
cc_531 N_A_27_47#_M1010_g N_A_644_47#_c_1331_n 0.0105205f $X=6.275 $Y=0.655
+ $X2=0 $Y2=0
cc_532 N_A_27_47#_M1017_g N_A_644_47#_c_1331_n 0.00865392f $X=6.705 $Y=0.655
+ $X2=0 $Y2=0
cc_533 N_A_27_47#_M1025_g N_A_644_47#_c_1333_n 0.00860735f $X=7.135 $Y=0.655
+ $X2=0 $Y2=0
cc_534 N_A_27_47#_M1028_g N_A_644_47#_c_1333_n 0.0100905f $X=7.565 $Y=0.655
+ $X2=0 $Y2=0
cc_535 N_A_27_47#_M1031_g N_A_644_47#_c_1335_n 0.00899305f $X=8.065 $Y=0.655
+ $X2=0 $Y2=0
cc_536 N_A_27_47#_M1033_g N_A_644_47#_c_1335_n 0.0104838f $X=8.565 $Y=0.655
+ $X2=0 $Y2=0
cc_537 N_A_27_47#_M1036_g N_A_644_47#_c_1337_n 0.00905372f $X=9.065 $Y=0.655
+ $X2=0 $Y2=0
cc_538 N_A_27_47#_M1039_g N_A_644_47#_c_1337_n 0.0100786f $X=9.565 $Y=0.655
+ $X2=0 $Y2=0
cc_539 N_A_27_47#_M1013_g N_A_644_47#_c_1302_n 9.7541e-19 $X=4.005 $Y=0.655
+ $X2=0 $Y2=0
cc_540 N_A_27_47#_c_307_n N_A_644_47#_c_1302_n 0.0209731f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_541 N_A_27_47#_c_309_n N_A_644_47#_c_1302_n 0.00248733f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_542 N_A_27_47#_M1022_g N_A_644_47#_c_1303_n 9.7541e-19 $X=4.985 $Y=0.655
+ $X2=0 $Y2=0
cc_543 N_A_27_47#_c_307_n N_A_644_47#_c_1303_n 0.0209731f $X=9.655 $Y=1.43 $X2=0
+ $Y2=0
cc_544 N_A_27_47#_c_309_n N_A_644_47#_c_1303_n 0.00272398f $X=10.045 $Y=1.43
+ $X2=0 $Y2=0
cc_545 N_A_27_47#_M1010_g N_A_644_47#_c_1345_n 6.29653e-19 $X=6.275 $Y=0.655
+ $X2=0 $Y2=0
cc_546 N_A_27_47#_M1017_g N_A_644_47#_c_1345_n 0.00735618f $X=6.705 $Y=0.655
+ $X2=0 $Y2=0
cc_547 N_A_27_47#_M1025_g N_A_644_47#_c_1345_n 0.00755965f $X=7.135 $Y=0.655
+ $X2=0 $Y2=0
cc_548 N_A_27_47#_M1028_g N_A_644_47#_c_1345_n 6.67164e-19 $X=7.565 $Y=0.655
+ $X2=0 $Y2=0
cc_549 N_A_27_47#_M1031_g N_A_644_47#_c_1349_n 0.00779673f $X=8.065 $Y=0.655
+ $X2=0 $Y2=0
cc_550 N_A_27_47#_M1033_g N_A_644_47#_c_1349_n 6.59874e-19 $X=8.565 $Y=0.655
+ $X2=0 $Y2=0
cc_551 N_A_27_47#_M1036_g N_A_644_47#_c_1351_n 0.00768151f $X=9.065 $Y=0.655
+ $X2=0 $Y2=0
cc_552 N_A_27_47#_M1039_g N_A_644_47#_c_1351_n 9.49589e-19 $X=9.565 $Y=0.655
+ $X2=0 $Y2=0
cc_553 N_A_114_367#_c_678_n N_VPWR_M1009_d 0.00341793f $X=2.265 $Y=2.11
+ $X2=0.495 $Y2=1.185
cc_554 N_A_114_367#_c_678_n N_VPWR_c_708_n 0.0135055f $X=2.265 $Y=2.11 $X2=1.425
+ $Y2=0.655
cc_555 N_A_114_367#_c_665_n N_VPWR_c_716_n 0.01906f $X=0.71 $Y=2.905 $X2=0.7
+ $Y2=1.35
cc_556 N_A_114_367#_c_670_n N_VPWR_c_716_n 0.0298674f $X=1.405 $Y=2.99 $X2=0.7
+ $Y2=1.35
cc_557 N_A_114_367#_c_674_n N_VPWR_c_716_n 0.01906f $X=1.57 $Y=2.905 $X2=0.7
+ $Y2=1.35
cc_558 N_A_114_367#_c_682_n N_VPWR_c_718_n 0.0189236f $X=2.43 $Y=2.91 $X2=1.38
+ $Y2=1.35
cc_559 N_A_114_367#_M1020_d N_VPWR_c_707_n 0.00223559f $X=0.57 $Y=1.835 $X2=0
+ $Y2=0
cc_560 N_A_114_367#_M1041_d N_VPWR_c_707_n 0.00223559f $X=1.43 $Y=1.835 $X2=0
+ $Y2=0
cc_561 N_A_114_367#_M1018_s N_VPWR_c_707_n 0.00223559f $X=2.29 $Y=1.835 $X2=0
+ $Y2=0
cc_562 N_A_114_367#_c_665_n N_VPWR_c_707_n 0.0124545f $X=0.71 $Y=2.905 $X2=0
+ $Y2=0
cc_563 N_A_114_367#_c_670_n N_VPWR_c_707_n 0.0187823f $X=1.405 $Y=2.99 $X2=0
+ $Y2=0
cc_564 N_A_114_367#_c_674_n N_VPWR_c_707_n 0.0124545f $X=1.57 $Y=2.905 $X2=0
+ $Y2=0
cc_565 N_A_114_367#_c_682_n N_VPWR_c_707_n 0.0123859f $X=2.43 $Y=2.91 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_707_n N_A_636_367#_M1002_s 0.00223559f $X=10.32 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_567 N_VPWR_c_707_n N_A_636_367#_M1007_s 0.00223559f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_707_n N_A_636_367#_M1021_s 0.00223559f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_707_n N_A_636_367#_M1034_s 0.00223559f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_707_n N_A_636_367#_M1011_d 0.00280658f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_707_n N_A_636_367#_M1016_d 0.00280658f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_707_n N_A_636_367#_M1032_d 0.00280658f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_707_n N_A_636_367#_M1038_d 0.00411415f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_709_n N_A_636_367#_c_854_n 0.0658787f $X=2.86 $Y=2.19 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_720_n N_A_636_367#_c_854_n 0.0189236f $X=3.665 $Y=3.33 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_707_n N_A_636_367#_c_854_n 0.0123859f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_577 N_VPWR_M1005_d N_A_636_367#_c_848_n 0.00176461f $X=3.61 $Y=1.835 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_710_n N_A_636_367#_c_848_n 0.0135055f $X=3.75 $Y=2.27 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_711_n N_A_636_367#_c_868_n 0.0189236f $X=4.525 $Y=3.33 $X2=0
+ $Y2=0
cc_580 N_VPWR_c_707_n N_A_636_367#_c_868_n 0.0123859f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_581 N_VPWR_M1014_d N_A_636_367#_c_850_n 0.00176461f $X=4.47 $Y=1.835 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_712_n N_A_636_367#_c_850_n 0.0135055f $X=4.61 $Y=2.27 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_722_n N_A_636_367#_c_876_n 0.0189236f $X=5.385 $Y=3.33 $X2=0
+ $Y2=0
cc_584 N_VPWR_c_707_n N_A_636_367#_c_876_n 0.0123859f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_585 N_VPWR_M1023_d N_A_636_367#_c_851_n 0.00176461f $X=5.33 $Y=1.835 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_713_n N_A_636_367#_c_851_n 0.0135055f $X=5.47 $Y=2.27 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_723_n N_A_636_367#_c_885_n 0.01906f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_707_n N_A_636_367#_c_885_n 0.0124545f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_723_n N_A_636_367#_c_891_n 0.0374555f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_707_n N_A_636_367#_c_891_n 0.0239316f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_591 N_VPWR_c_723_n N_A_636_367#_c_895_n 0.0374555f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_707_n N_A_636_367#_c_895_n 0.0239316f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_593 N_VPWR_c_723_n N_A_636_367#_c_899_n 0.0374555f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_707_n N_A_636_367#_c_899_n 0.0239316f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_723_n N_A_636_367#_c_903_n 0.0495958f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_707_n N_A_636_367#_c_903_n 0.030825f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_723_n N_A_636_367#_c_913_n 0.0207136f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_707_n N_A_636_367#_c_913_n 0.0126421f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_VPWR_c_723_n N_A_636_367#_c_914_n 0.0207136f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_707_n N_A_636_367#_c_914_n 0.0126421f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_723_n N_A_636_367#_c_915_n 0.0207136f $X=10.095 $Y=3.33 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_707_n N_A_636_367#_c_915_n 0.0126421f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_707_n N_X_M1004_s 0.00281482f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_604 N_VPWR_c_707_n N_X_M1015_s 0.00281482f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_605 N_VPWR_c_707_n N_X_M1030_s 0.00281482f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_606 N_VPWR_c_707_n N_X_M1037_s 0.00281482f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_607 N_VPWR_M1035_d N_X_c_983_n 0.00310428f $X=10.12 $Y=1.835 $X2=0 $Y2=0
cc_608 N_VPWR_c_715_n N_X_c_983_n 0.0243264f $X=10.26 $Y=2.27 $X2=0 $Y2=0
cc_609 N_A_636_367#_c_891_n N_X_M1004_s 0.00472489f $X=6.735 $Y=2.99 $X2=0 $Y2=0
cc_610 N_A_636_367#_c_895_n N_X_M1015_s 0.00472489f $X=7.735 $Y=2.99 $X2=0 $Y2=0
cc_611 N_A_636_367#_c_899_n N_X_M1030_s 0.00472489f $X=8.735 $Y=2.99 $X2=0 $Y2=0
cc_612 N_A_636_367#_c_903_n N_X_M1037_s 0.00472489f $X=9.745 $Y=2.99 $X2=0 $Y2=0
cc_613 N_A_636_367#_c_891_n N_X_c_988_n 0.0196355f $X=6.735 $Y=2.99 $X2=0 $Y2=0
cc_614 N_A_636_367#_M1011_d N_X_c_979_n 0.00250873f $X=6.69 $Y=1.835 $X2=0 $Y2=0
cc_615 N_A_636_367#_c_893_n N_X_c_979_n 0.0209867f $X=6.9 $Y=2.27 $X2=0 $Y2=0
cc_616 N_A_636_367#_c_851_n N_X_c_980_n 0.0104256f $X=5.735 $Y=1.85 $X2=0 $Y2=0
cc_617 N_A_636_367#_c_895_n N_X_c_1005_n 0.0196355f $X=7.735 $Y=2.99 $X2=0 $Y2=0
cc_618 N_A_636_367#_M1016_d N_X_c_981_n 0.00250873f $X=7.69 $Y=1.835 $X2=0 $Y2=0
cc_619 N_A_636_367#_c_897_n N_X_c_981_n 0.0209867f $X=7.9 $Y=2.27 $X2=0 $Y2=0
cc_620 N_A_636_367#_c_899_n N_X_c_1017_n 0.0196355f $X=8.735 $Y=2.99 $X2=0 $Y2=0
cc_621 N_A_636_367#_M1032_d N_X_c_982_n 0.00250873f $X=8.69 $Y=1.835 $X2=0 $Y2=0
cc_622 N_A_636_367#_c_901_n N_X_c_982_n 0.0209867f $X=8.9 $Y=2.27 $X2=0 $Y2=0
cc_623 N_A_636_367#_c_903_n N_X_c_1027_n 0.0196355f $X=9.745 $Y=2.99 $X2=0 $Y2=0
cc_624 N_A_636_367#_M1038_d N_X_c_983_n 0.00176461f $X=9.69 $Y=1.835 $X2=0 $Y2=0
cc_625 N_A_636_367#_c_969_p N_X_c_983_n 0.0135055f $X=9.83 $Y=2.27 $X2=0 $Y2=0
cc_626 N_X_c_974_n N_VGND_M1043_d 0.00378225f $X=9.995 $Y=1.01 $X2=0 $Y2=0
cc_627 N_X_c_974_n N_VGND_c_1162_n 0.0236357f $X=9.995 $Y=1.01 $X2=0 $Y2=0
cc_628 N_X_M1010_s N_VGND_c_1172_n 0.00225186f $X=6.35 $Y=0.235 $X2=0 $Y2=0
cc_629 N_X_M1025_s N_VGND_c_1172_n 0.00225186f $X=7.21 $Y=0.235 $X2=0 $Y2=0
cc_630 N_X_M1031_s N_VGND_c_1172_n 0.00281482f $X=8.14 $Y=0.235 $X2=0 $Y2=0
cc_631 N_X_M1036_s N_VGND_c_1172_n 0.00281482f $X=9.14 $Y=0.235 $X2=0 $Y2=0
cc_632 N_X_c_970_n N_A_644_47#_M1017_d 0.00176461f $X=7.265 $Y=1.01 $X2=0 $Y2=0
cc_633 N_X_c_972_n N_A_644_47#_M1028_d 0.00250873f $X=8.185 $Y=1.01 $X2=0 $Y2=0
cc_634 N_X_c_973_n N_A_644_47#_M1033_d 0.00250873f $X=9.185 $Y=1.01 $X2=0 $Y2=0
cc_635 N_X_c_974_n N_A_644_47#_M1039_d 0.00229612f $X=9.995 $Y=1.01 $X2=0 $Y2=0
cc_636 N_X_c_971_n N_A_644_47#_c_1301_n 0.00772305f $X=6.575 $Y=1.01 $X2=0 $Y2=0
cc_637 N_X_M1010_s N_A_644_47#_c_1331_n 0.00332344f $X=6.35 $Y=0.235 $X2=0 $Y2=0
cc_638 N_X_c_1100_p N_A_644_47#_c_1331_n 0.0123414f $X=6.49 $Y=0.845 $X2=0 $Y2=0
cc_639 N_X_c_970_n N_A_644_47#_c_1331_n 0.00350153f $X=7.265 $Y=1.01 $X2=0 $Y2=0
cc_640 N_X_M1025_s N_A_644_47#_c_1333_n 0.00332344f $X=7.21 $Y=0.235 $X2=0 $Y2=0
cc_641 N_X_c_970_n N_A_644_47#_c_1333_n 0.00350153f $X=7.265 $Y=1.01 $X2=0 $Y2=0
cc_642 N_X_c_1007_n N_A_644_47#_c_1333_n 0.0140107f $X=7.35 $Y=0.845 $X2=0 $Y2=0
cc_643 N_X_c_972_n N_A_644_47#_c_1333_n 0.00350153f $X=8.185 $Y=1.01 $X2=0 $Y2=0
cc_644 N_X_M1031_s N_A_644_47#_c_1335_n 0.00472489f $X=8.14 $Y=0.235 $X2=0 $Y2=0
cc_645 N_X_c_972_n N_A_644_47#_c_1335_n 0.00351559f $X=8.185 $Y=1.01 $X2=0 $Y2=0
cc_646 N_X_c_973_n N_A_644_47#_c_1335_n 0.00351559f $X=9.185 $Y=1.01 $X2=0 $Y2=0
cc_647 N_X_c_976_n N_A_644_47#_c_1335_n 0.0192149f $X=8.35 $Y=0.805 $X2=0 $Y2=0
cc_648 N_X_M1036_s N_A_644_47#_c_1337_n 0.00472489f $X=9.14 $Y=0.235 $X2=0 $Y2=0
cc_649 N_X_c_973_n N_A_644_47#_c_1337_n 0.00351559f $X=9.185 $Y=1.01 $X2=0 $Y2=0
cc_650 N_X_c_974_n N_A_644_47#_c_1337_n 0.00350153f $X=9.995 $Y=1.01 $X2=0 $Y2=0
cc_651 N_X_c_977_n N_A_644_47#_c_1337_n 0.0192149f $X=9.35 $Y=0.845 $X2=0 $Y2=0
cc_652 N_X_c_974_n N_A_644_47#_c_1373_n 0.0171413f $X=9.995 $Y=1.01 $X2=0 $Y2=0
cc_653 N_X_c_970_n N_A_644_47#_c_1345_n 0.0167374f $X=7.265 $Y=1.01 $X2=0 $Y2=0
cc_654 N_X_c_972_n N_A_644_47#_c_1349_n 0.0205104f $X=8.185 $Y=1.01 $X2=0 $Y2=0
cc_655 N_X_c_973_n N_A_644_47#_c_1351_n 0.0205104f $X=9.185 $Y=1.01 $X2=0 $Y2=0
cc_656 N_A_114_47#_c_1120_n N_VGND_M1000_s 0.00330371f $X=2.335 $Y=0.892
+ $X2=0.495 $Y2=1.185
cc_657 N_A_114_47#_c_1120_n N_VGND_c_1154_n 0.0152022f $X=2.335 $Y=0.892
+ $X2=1.425 $Y2=0.655
cc_658 N_A_114_47#_c_1118_n N_VGND_c_1163_n 0.0378082f $X=1.555 $Y=0.34 $X2=0
+ $Y2=0
cc_659 N_A_114_47#_c_1143_p N_VGND_c_1163_n 0.0118138f $X=1.64 $Y=0.425 $X2=0
+ $Y2=0
cc_660 N_A_114_47#_c_1131_n N_VGND_c_1163_n 0.0184671f $X=0.71 $Y=0.34 $X2=0
+ $Y2=0
cc_661 N_A_114_47#_c_1128_n N_VGND_c_1165_n 0.0189236f $X=2.5 $Y=0.42 $X2=0
+ $Y2=0
cc_662 N_A_114_47#_M1003_d N_VGND_c_1172_n 0.00225167f $X=0.57 $Y=0.235 $X2=2.16
+ $Y2=1.347
cc_663 N_A_114_47#_M1008_d N_VGND_c_1172_n 0.0025412f $X=1.5 $Y=0.235 $X2=2.16
+ $Y2=1.347
cc_664 N_A_114_47#_M1024_d N_VGND_c_1172_n 0.00223559f $X=2.36 $Y=0.235 $X2=2.16
+ $Y2=1.347
cc_665 N_A_114_47#_c_1118_n N_VGND_c_1172_n 0.0242404f $X=1.555 $Y=0.34 $X2=2.16
+ $Y2=1.347
cc_666 N_A_114_47#_c_1143_p N_VGND_c_1172_n 0.00658808f $X=1.64 $Y=0.425
+ $X2=2.16 $Y2=1.347
cc_667 N_A_114_47#_c_1120_n N_VGND_c_1172_n 0.0125005f $X=2.335 $Y=0.892
+ $X2=2.16 $Y2=1.347
cc_668 N_A_114_47#_c_1128_n N_VGND_c_1172_n 0.0123859f $X=2.5 $Y=0.42 $X2=2.16
+ $Y2=1.347
cc_669 N_A_114_47#_c_1131_n N_VGND_c_1172_n 0.0123739f $X=0.71 $Y=0.34 $X2=2.16
+ $Y2=1.347
cc_670 N_VGND_c_1172_n N_A_644_47#_M1001_s 0.0041489f $X=10.32 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_671 N_VGND_c_1172_n N_A_644_47#_M1013_s 0.0041489f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_672 N_VGND_c_1172_n N_A_644_47#_M1022_s 0.0041489f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_673 N_VGND_c_1172_n N_A_644_47#_M1040_s 0.00223559f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_674 N_VGND_c_1172_n N_A_644_47#_M1017_d 0.00225167f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_675 N_VGND_c_1172_n N_A_644_47#_M1028_d 0.00280658f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_676 N_VGND_c_1172_n N_A_644_47#_M1033_d 0.00280658f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_677 N_VGND_c_1172_n N_A_644_47#_M1039_d 0.00352348f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_678 N_VGND_c_1167_n N_A_644_47#_c_1304_n 0.0153332f $X=3.625 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_1172_n N_A_644_47#_c_1304_n 0.00945339f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_680 N_VGND_M1012_d N_A_644_47#_c_1298_n 0.00176461f $X=3.65 $Y=0.235 $X2=0
+ $Y2=0
cc_681 N_VGND_c_1156_n N_A_644_47#_c_1298_n 0.0153337f $X=3.79 $Y=0.485 $X2=0
+ $Y2=0
cc_682 N_VGND_c_1155_n N_A_644_47#_c_1299_n 0.00752767f $X=2.93 $Y=0.38 $X2=0
+ $Y2=0
cc_683 N_VGND_c_1157_n N_A_644_47#_c_1312_n 0.0153332f $X=4.485 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1172_n N_A_644_47#_c_1312_n 0.00945339f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_685 N_VGND_M1019_d N_A_644_47#_c_1300_n 0.00444361f $X=4.51 $Y=0.235 $X2=0
+ $Y2=0
cc_686 N_VGND_c_1158_n N_A_644_47#_c_1300_n 0.0219238f $X=4.65 $Y=0.485 $X2=0
+ $Y2=0
cc_687 N_VGND_c_1158_n N_A_644_47#_c_1318_n 0.0312008f $X=4.65 $Y=0.485 $X2=0
+ $Y2=0
cc_688 N_VGND_c_1159_n N_A_644_47#_c_1318_n 0.0153332f $X=5.465 $Y=0 $X2=0 $Y2=0
cc_689 N_VGND_c_1172_n N_A_644_47#_c_1318_n 0.00945339f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_690 N_VGND_M1029_d N_A_644_47#_c_1301_n 0.00176461f $X=5.49 $Y=0.235 $X2=0
+ $Y2=0
cc_691 N_VGND_c_1160_n N_A_644_47#_c_1301_n 0.0153337f $X=5.63 $Y=0.485 $X2=0
+ $Y2=0
cc_692 N_VGND_c_1169_n N_A_644_47#_c_1325_n 0.01906f $X=10.115 $Y=0 $X2=0 $Y2=0
cc_693 N_VGND_c_1172_n N_A_644_47#_c_1325_n 0.0124545f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_694 N_VGND_c_1169_n N_A_644_47#_c_1331_n 0.0298936f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_695 N_VGND_c_1172_n N_A_644_47#_c_1331_n 0.0187857f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_696 N_VGND_c_1169_n N_A_644_47#_c_1333_n 0.0330447f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_697 N_VGND_c_1172_n N_A_644_47#_c_1333_n 0.0213073f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_698 N_VGND_c_1169_n N_A_644_47#_c_1335_n 0.0374817f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_699 N_VGND_c_1172_n N_A_644_47#_c_1335_n 0.0239391f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_700 N_VGND_c_1169_n N_A_644_47#_c_1337_n 0.0538929f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_701 N_VGND_c_1172_n N_A_644_47#_c_1337_n 0.0339442f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_702 N_VGND_c_1169_n N_A_644_47#_c_1345_n 0.0186595f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_703 N_VGND_c_1172_n N_A_644_47#_c_1345_n 0.0124318f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_704 N_VGND_c_1169_n N_A_644_47#_c_1349_n 0.0202403f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_705 N_VGND_c_1172_n N_A_644_47#_c_1349_n 0.0125416f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_706 N_VGND_c_1169_n N_A_644_47#_c_1351_n 0.0202403f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_707 N_VGND_c_1172_n N_A_644_47#_c_1351_n 0.0125416f $X=10.32 $Y=0 $X2=0 $Y2=0
