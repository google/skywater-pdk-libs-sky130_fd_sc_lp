* File: sky130_fd_sc_lp__a2bb2oi_lp.spice
* Created: Wed Sep  2 09:24:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2oi_lp  VNB VPB B1 B2 A2_N A1_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 A_170_47# N_B1_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_B2_M1001_g A_170_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1006 A_334_47# N_A_296_146#_M1006_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_296_146#_M1004_g A_334_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.0441 PD=0.71 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1011 A_494_47# N_A2_N_M1011_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0609 PD=0.63 PS=0.71 NRD=14.28 NRS=2.856 M=1 R=2.8 SA=75001.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_A_296_146#_M1012_d N_A2_N_M1012_g A_494_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_652_47# N_A1_N_M1005_g N_A_296_146#_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A1_N_M1000_g A_652_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_A_27_409#_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 N_A_27_409#_M1007_d N_B2_M1007_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1002 N_Y_M1002_d N_A_296_146#_M1002_g N_A_27_409#_M1007_d VPB PHIGHVT L=0.25
+ W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1008 N_A_296_146#_M1008_d N_A2_N_M1008_g N_A_456_339#_M1008_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A1_N_M1009_g N_A_456_339#_M1009_s VPB PHIGHVT L=0.25 W=1
+ AD=0.28 AS=0.285 PD=2.56 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=8.9307 P=13.41
*
.include "sky130_fd_sc_lp__a2bb2oi_lp.pxi.spice"
*
.ends
*
*
