* File: sky130_fd_sc_lp__nor3_4.pex.spice
* Created: Wed Sep  2 10:09:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31 32
+ 47
r73 45 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.685 $Y=1.35
+ $X2=1.775 $Y2=1.35
r74 43 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.345 $Y=1.35
+ $X2=1.685 $Y2=1.35
r75 42 43 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.915 $Y=1.35
+ $X2=1.345 $Y2=1.35
r76 41 42 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.485 $Y=1.35
+ $X2=0.915 $Y2=1.35
r77 38 41 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.325 $Y=1.35
+ $X2=0.485 $Y2=1.35
r78 32 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.685
+ $Y=1.35 $X2=1.685 $Y2=1.35
r79 31 32 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.362
+ $X2=1.68 $Y2=1.362
r80 30 31 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.362
+ $X2=1.2 $Y2=1.362
r81 29 30 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.362
+ $X2=0.72 $Y2=1.362
r82 29 38 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.325
+ $Y=1.35 $X2=0.325 $Y2=1.35
r83 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.515
+ $X2=1.775 $Y2=1.35
r84 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.775 $Y=1.515
+ $X2=1.775 $Y2=2.465
r85 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.185
+ $X2=1.775 $Y2=1.35
r86 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.775 $Y=1.185
+ $X2=1.775 $Y2=0.655
r87 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.515
+ $X2=1.345 $Y2=1.35
r88 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.345 $Y=1.515
+ $X2=1.345 $Y2=2.465
r89 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.185
+ $X2=1.345 $Y2=1.35
r90 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.345 $Y=1.185
+ $X2=1.345 $Y2=0.655
r91 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.515
+ $X2=0.915 $Y2=1.35
r92 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.915 $Y=1.515
+ $X2=0.915 $Y2=2.465
r93 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.185
+ $X2=0.915 $Y2=1.35
r94 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.915 $Y=1.185
+ $X2=0.915 $Y2=0.655
r95 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.515
+ $X2=0.485 $Y2=1.35
r96 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.485 $Y=1.515
+ $X2=0.485 $Y2=2.465
r97 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.185
+ $X2=0.485 $Y2=1.35
r98 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.485 $Y=1.185
+ $X2=0.485 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_4%B 1 3 6 8 10 13 15 17 20 24 27 29 31 35 37 38
+ 39 53 56 70
r125 51 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.975 $Y=1.35
+ $X2=3.065 $Y2=1.35
r126 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.35 $X2=2.975 $Y2=1.35
r127 49 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.975 $Y2=1.35
r128 47 49 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.295 $Y=1.35
+ $X2=2.635 $Y2=1.35
r129 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=1.35 $X2=2.295 $Y2=1.35
r130 44 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.295 $Y2=1.35
r131 39 70 7.9186 $w=4.38e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.295
+ $X2=3.25 $Y2=1.295
r132 39 52 3.03847 $w=4.73e-07 $l=6e-08 $layer=LI1_cond $X=3.035 $Y=1.362
+ $X2=2.975 $Y2=1.362
r133 38 52 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=2.64 $Y=1.362
+ $X2=2.975 $Y2=1.362
r134 38 48 13.0358 $w=3.03e-07 $l=3.45e-07 $layer=LI1_cond $X=2.64 $Y=1.362
+ $X2=2.295 $Y2=1.362
r135 37 48 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.16 $Y=1.362
+ $X2=2.295 $Y2=1.362
r136 35 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.235 $Y=1.35
+ $X2=5.235 $Y2=1.515
r137 35 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.235 $Y=1.35
+ $X2=5.235 $Y2=1.185
r138 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.235
+ $Y=1.35 $X2=5.235 $Y2=1.35
r139 31 34 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=5.2 $Y=1.16 $X2=5.2
+ $Y2=1.35
r140 29 31 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.07 $Y=1.16 $X2=5.2
+ $Y2=1.16
r141 29 70 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=5.07 $Y=1.16
+ $X2=3.25 $Y2=1.16
r142 27 57 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.215 $Y=2.465
+ $X2=5.215 $Y2=1.515
r143 24 56 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.215 $Y=0.655
+ $X2=5.215 $Y2=1.185
r144 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.515
+ $X2=3.065 $Y2=1.35
r145 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.065 $Y=1.515
+ $X2=3.065 $Y2=2.465
r146 15 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.185
+ $X2=3.065 $Y2=1.35
r147 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.065 $Y=1.185
+ $X2=3.065 $Y2=0.655
r148 11 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.515
+ $X2=2.635 $Y2=1.35
r149 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.635 $Y=1.515
+ $X2=2.635 $Y2=2.465
r150 8 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.185
+ $X2=2.635 $Y2=1.35
r151 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.635 $Y=1.185
+ $X2=2.635 $Y2=0.655
r152 4 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.515
+ $X2=2.205 $Y2=1.35
r153 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.205 $Y=1.515
+ $X2=2.205 $Y2=2.465
r154 1 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.185
+ $X2=2.205 $Y2=1.35
r155 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.205 $Y=1.185
+ $X2=2.205 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_4%C 3 7 11 15 19 23 27 31 35 38 39 50 52 59 61
c95 31 0 1.28803e-19 $X=4.785 $Y=2.465
c96 23 0 1.19111e-20 $X=4.355 $Y=2.465
r97 52 59 0.658539 $w=3.48e-07 $l=2e-08 $layer=LI1_cond $X=4.06 $Y=1.59 $X2=4.08
+ $Y2=1.59
r98 46 48 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.925 $Y=1.51
+ $X2=4.355 $Y2=1.51
r99 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.925
+ $Y=1.51 $X2=3.925 $Y2=1.51
r100 43 46 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.495 $Y=1.51
+ $X2=3.925 $Y2=1.51
r101 39 61 5.40486 $w=3.48e-07 $l=1.23e-07 $layer=LI1_cond $X=4.112 $Y=1.59
+ $X2=4.235 $Y2=1.59
r102 39 59 1.05366 $w=3.48e-07 $l=3.2e-08 $layer=LI1_cond $X=4.112 $Y=1.59
+ $X2=4.08 $Y2=1.59
r103 39 52 1.08659 $w=3.48e-07 $l=3.3e-08 $layer=LI1_cond $X=4.027 $Y=1.59
+ $X2=4.06 $Y2=1.59
r104 39 47 3.35855 $w=3.48e-07 $l=1.02e-07 $layer=LI1_cond $X=4.027 $Y=1.59
+ $X2=3.925 $Y2=1.59
r105 38 47 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=3.6 $Y=1.59
+ $X2=3.925 $Y2=1.59
r106 36 50 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.605 $Y=1.51
+ $X2=4.785 $Y2=1.51
r107 36 48 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.605 $Y=1.51
+ $X2=4.355 $Y2=1.51
r108 35 61 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.605 $Y=1.53
+ $X2=4.235 $Y2=1.53
r109 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.605
+ $Y=1.51 $X2=4.605 $Y2=1.51
r110 29 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.675
+ $X2=4.785 $Y2=1.51
r111 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.785 $Y=1.675
+ $X2=4.785 $Y2=2.465
r112 25 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.345
+ $X2=4.785 $Y2=1.51
r113 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.785 $Y=1.345
+ $X2=4.785 $Y2=0.655
r114 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.675
+ $X2=4.355 $Y2=1.51
r115 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.355 $Y=1.675
+ $X2=4.355 $Y2=2.465
r116 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.345
+ $X2=4.355 $Y2=1.51
r117 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.355 $Y=1.345
+ $X2=4.355 $Y2=0.655
r118 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=1.675
+ $X2=3.925 $Y2=1.51
r119 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.925 $Y=1.675
+ $X2=3.925 $Y2=2.465
r120 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=1.345
+ $X2=3.925 $Y2=1.51
r121 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.925 $Y=1.345
+ $X2=3.925 $Y2=0.655
r122 5 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.675
+ $X2=3.495 $Y2=1.51
r123 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.495 $Y=1.675
+ $X2=3.495 $Y2=2.465
r124 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.345
+ $X2=3.495 $Y2=1.51
r125 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.495 $Y=1.345
+ $X2=3.495 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_4%A_29_367# 1 2 3 4 5 18 22 23 26 30 34 38 43
+ 44 45 48 50 51 53
c77 48 0 1.28803e-19 $X=5.45 $Y=2.95
r78 53 55 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.45 $Y=2.24
+ $X2=5.45 $Y2=2.41
r79 46 55 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=2.495
+ $X2=5.45 $Y2=2.41
r80 46 48 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.45 $Y=2.495
+ $X2=5.45 $Y2=2.95
r81 44 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=2.41
+ $X2=5.45 $Y2=2.41
r82 44 45 148.096 $w=1.68e-07 $l=2.27e-06 $layer=LI1_cond $X=5.285 $Y=2.41
+ $X2=3.015 $Y2=2.41
r83 41 45 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.885 $Y=2.325
+ $X2=3.015 $Y2=2.41
r84 41 43 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=2.885 $Y=2.325
+ $X2=2.885 $Y2=1.98
r85 40 43 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.885 $Y=1.875
+ $X2=2.885 $Y2=1.98
r86 39 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.085 $Y=1.79
+ $X2=1.99 $Y2=1.79
r87 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.755 $Y=1.79
+ $X2=2.885 $Y2=1.875
r88 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.755 $Y=1.79
+ $X2=2.085 $Y2=1.79
r89 34 36 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.99 $Y=1.98
+ $X2=1.99 $Y2=2.91
r90 32 51 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=1.875
+ $X2=1.99 $Y2=1.79
r91 32 34 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=1.99 $Y=1.875
+ $X2=1.99 $Y2=1.98
r92 31 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.225 $Y=1.79
+ $X2=1.13 $Y2=1.79
r93 30 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.895 $Y=1.79
+ $X2=1.99 $Y2=1.79
r94 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.895 $Y=1.79
+ $X2=1.225 $Y2=1.79
r95 26 28 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.13 $Y=1.98
+ $X2=1.13 $Y2=2.91
r96 24 50 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=1.875
+ $X2=1.13 $Y2=1.79
r97 24 26 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=1.13 $Y=1.875
+ $X2=1.13 $Y2=1.98
r98 22 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.035 $Y=1.79
+ $X2=1.13 $Y2=1.79
r99 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.035 $Y=1.79
+ $X2=0.365 $Y2=1.79
r100 18 20 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.235 $Y=1.98
+ $X2=0.235 $Y2=2.91
r101 16 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.235 $Y=1.875
+ $X2=0.365 $Y2=1.79
r102 16 18 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=0.235 $Y=1.875
+ $X2=0.235 $Y2=1.98
r103 5 53 400 $w=1.7e-07 $l=4.78357e-07 $layer=licon1_PDIFF $count=1 $X=5.29
+ $Y=1.835 $X2=5.45 $Y2=2.24
r104 5 48 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=5.29
+ $Y=1.835 $X2=5.45 $Y2=2.95
r105 4 43 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=1.98
r106 3 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=1.99 $Y2=2.91
r107 3 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=1.99 $Y2=1.98
r108 2 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=2.91
r109 2 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=1.98
r110 1 20 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.91
r111 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_4%VPWR 1 2 9 15 19 21 26 33 34 37 40
r68 40 41 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 33 34 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r71 31 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=1.56 $Y2=3.33
r72 31 33 247.588 $w=1.68e-07 $l=3.795e-06 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r76 27 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=0.7 $Y2=3.33
r77 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.56 $Y2=3.33
r79 26 29 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.2 $Y2=3.33
r80 24 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r82 21 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.7 $Y2=3.33
r83 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 19 34 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 19 41 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.68 $Y2=3.33
r86 15 18 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.56 $Y=2.19
+ $X2=1.56 $Y2=2.95
r87 13 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=3.245
+ $X2=1.56 $Y2=3.33
r88 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.56 $Y=3.245
+ $X2=1.56 $Y2=2.95
r89 9 12 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.7 $Y=2.19 $X2=0.7
+ $Y2=2.95
r90 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=3.33
r91 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=2.95
r92 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.835 $X2=1.56 $Y2=2.95
r93 2 15 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.835 $X2=1.56 $Y2=2.19
r94 1 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.95
r95 1 9 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_4%A_456_367# 1 2 3 4 13 15 23
r31 21 23 24.7775 $w=3.98e-07 $l=8.6e-07 $layer=LI1_cond $X=4.14 $Y=2.875 $X2=5
+ $Y2=2.875
r32 19 21 24.7775 $w=3.98e-07 $l=8.6e-07 $layer=LI1_cond $X=3.28 $Y=2.875
+ $X2=4.14 $Y2=2.875
r33 17 26 3.11842 $w=4e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=2.875
+ $X2=2.42 $Y2=2.875
r34 17 19 20.0237 $w=3.98e-07 $l=6.95e-07 $layer=LI1_cond $X=2.585 $Y=2.875
+ $X2=3.28 $Y2=2.875
r35 13 26 3.77991 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=2.42 $Y=2.675 $X2=2.42
+ $Y2=2.875
r36 13 15 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.42 $Y=2.675
+ $X2=2.42 $Y2=2.14
r37 4 23 600 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=4.86
+ $Y=1.835 $X2=5 $Y2=2.84
r38 3 21 600 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=1.835 $X2=4.14 $Y2=2.84
r39 2 19 600 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.835 $X2=3.28 $Y2=2.84
r40 1 26 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=2.95
r41 1 15 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_4%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 41 45 47
+ 49 55 57 59 63 65 68 69 72 73 74 75 81 82 85 88 90
c144 59 0 1.19111e-20 $X=5.5 $Y=1.9
r145 85 88 2.48781 $w=3.13e-07 $l=6.8e-08 $layer=LI1_cond $X=2.708 $Y=0.882
+ $X2=2.64 $Y2=0.882
r146 82 90 7.8772 $w=3.13e-07 $l=1.49e-07 $layer=LI1_cond $X=2.716 $Y=0.882
+ $X2=2.865 $Y2=0.882
r147 82 85 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=2.716 $Y=0.882
+ $X2=2.708 $Y2=0.882
r148 82 88 0.329269 $w=3.13e-07 $l=9e-09 $layer=LI1_cond $X=2.631 $Y=0.882
+ $X2=2.64 $Y2=0.882
r149 78 79 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=4.57 $Y=1.98
+ $X2=4.57 $Y2=2.045
r150 75 78 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.57 $Y=1.9 $X2=4.57
+ $Y2=1.98
r151 70 82 3.14635 $w=3.13e-07 $l=8.6e-08 $layer=LI1_cond $X=2.545 $Y=0.882
+ $X2=2.631 $Y2=0.882
r152 70 72 4.76034 $w=2.42e-07 $l=1.1e-07 $layer=LI1_cond $X=2.545 $Y=0.882
+ $X2=2.435 $Y2=0.882
r153 67 68 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.585 $Y=0.895
+ $X2=5.585 $Y2=1.815
r154 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0.81 $X2=5
+ $Y2=0.81
r155 65 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.5 $Y=0.81
+ $X2=5.585 $Y2=0.895
r156 65 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.5 $Y=0.81
+ $X2=5.165 $Y2=0.81
r157 61 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.725 $X2=5
+ $Y2=0.81
r158 61 63 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5 $Y=0.725 $X2=5
+ $Y2=0.42
r159 60 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=1.9
+ $X2=4.57 $Y2=1.9
r160 59 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.5 $Y=1.9
+ $X2=5.585 $Y2=1.815
r161 59 60 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.5 $Y=1.9
+ $X2=4.735 $Y2=1.9
r162 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0.81
+ $X2=4.14 $Y2=0.81
r163 57 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.81 $X2=5
+ $Y2=0.81
r164 57 58 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.835 $Y=0.81
+ $X2=4.305 $Y2=0.81
r165 53 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.725
+ $X2=4.14 $Y2=0.81
r166 53 55 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.14 $Y=0.725
+ $X2=4.14 $Y2=0.42
r167 49 79 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=2.045
+ $X2=4.57 $Y2=2.045
r168 49 51 36.4067 $w=2.18e-07 $l=6.95e-07 $layer=LI1_cond $X=4.405 $Y=2.045
+ $X2=3.71 $Y2=2.045
r169 48 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=0.81
+ $X2=3.28 $Y2=0.81
r170 47 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0.81
+ $X2=4.14 $Y2=0.81
r171 47 48 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.975 $Y=0.81
+ $X2=3.445 $Y2=0.81
r172 43 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=0.725
+ $X2=3.28 $Y2=0.81
r173 43 45 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.28 $Y=0.725
+ $X2=3.28 $Y2=0.42
r174 41 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0.81
+ $X2=3.28 $Y2=0.81
r175 41 90 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.115 $Y=0.81
+ $X2=2.865 $Y2=0.81
r176 37 72 1.69544 $w=2.2e-07 $l=1.57e-07 $layer=LI1_cond $X=2.435 $Y=0.725
+ $X2=2.435 $Y2=0.882
r177 37 39 15.9771 $w=2.18e-07 $l=3.05e-07 $layer=LI1_cond $X=2.435 $Y=0.725
+ $X2=2.435 $Y2=0.42
r178 36 69 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.655 $Y=0.955
+ $X2=1.56 $Y2=0.955
r179 35 72 4.76034 $w=2.42e-07 $l=1.4188e-07 $layer=LI1_cond $X=2.325 $Y=0.955
+ $X2=2.435 $Y2=0.882
r180 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.325 $Y=0.955
+ $X2=1.655 $Y2=0.955
r181 31 69 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=0.87
+ $X2=1.56 $Y2=0.955
r182 31 33 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.56 $Y=0.87
+ $X2=1.56 $Y2=0.42
r183 29 69 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.465 $Y=0.955
+ $X2=1.56 $Y2=0.955
r184 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.465 $Y=0.955
+ $X2=0.795 $Y2=0.955
r185 25 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.685 $Y=0.87
+ $X2=0.795 $Y2=0.955
r186 25 27 23.5727 $w=2.18e-07 $l=4.5e-07 $layer=LI1_cond $X=0.685 $Y=0.87
+ $X2=0.685 $Y2=0.42
r187 8 78 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.835 $X2=4.57 $Y2=1.98
r188 7 51 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.835 $X2=3.71 $Y2=2.04
r189 6 63 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=0.235 $X2=5 $Y2=0.42
r190 5 55 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4
+ $Y=0.235 $X2=4.14 $Y2=0.42
r191 4 45 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.235 $X2=3.28 $Y2=0.42
r192 3 72 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.235 $X2=2.42 $Y2=0.875
r193 3 39 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.235 $X2=2.42 $Y2=0.42
r194 2 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.235 $X2=1.56 $Y2=0.42
r195 1 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.235 $X2=0.7 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46 48
+ 51 52 54 55 57 58 59 61 76 80 89 92 96
r110 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r111 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r112 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r113 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r114 84 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r115 84 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r116 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r117 81 92 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.57
+ $Y2=0
r118 81 83 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.665 $Y=0
+ $X2=5.04 $Y2=0
r119 80 95 4.03428 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=5.335 $Y=0
+ $X2=5.547 $Y2=0
r120 80 83 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.04
+ $Y2=0
r121 79 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r122 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r123 76 92 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.57
+ $Y2=0
r124 76 78 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.08 $Y2=0
r125 75 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r126 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r127 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r128 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r129 69 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r130 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r131 66 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=0 $X2=1.13
+ $Y2=0
r132 66 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.295 $Y=0
+ $X2=1.68 $Y2=0
r133 65 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r134 65 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r135 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r136 62 86 4.47533 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.202 $Y2=0
r137 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.72 $Y2=0
r138 61 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.13
+ $Y2=0
r139 61 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.72
+ $Y2=0
r140 59 75 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r141 59 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r142 57 74 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.6
+ $Y2=0
r143 57 58 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.71
+ $Y2=0
r144 56 78 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=4.08 $Y2=0
r145 56 58 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.71
+ $Y2=0
r146 54 71 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.64
+ $Y2=0
r147 54 55 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.83
+ $Y2=0
r148 53 74 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.6
+ $Y2=0
r149 53 55 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.83
+ $Y2=0
r150 51 68 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=1.68 $Y2=0
r151 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.99
+ $Y2=0
r152 50 71 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.155 $Y=0
+ $X2=2.64 $Y2=0
r153 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=1.99
+ $Y2=0
r154 46 95 3.17794 $w=2.6e-07 $l=1.19143e-07 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.547 $Y2=0
r155 46 48 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.465 $Y2=0.38
r156 42 92 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0
r157 42 44 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0.39
r158 38 58 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.71 $Y2=0
r159 38 40 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.71 $Y2=0.39
r160 34 55 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0
r161 34 36 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0.39
r162 30 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0
r163 30 32 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0.57
r164 26 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0
r165 26 28 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0.57
r166 22 86 3.04234 $w=3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.202 $Y2=0
r167 22 24 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.38
r168 7 48 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.235 $X2=5.43 $Y2=0.38
r169 6 44 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.235 $X2=4.57 $Y2=0.39
r170 5 40 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.71 $Y2=0.39
r171 4 36 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.235 $X2=2.85 $Y2=0.39
r172 3 32 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=1.85
+ $Y=0.235 $X2=1.99 $Y2=0.57
r173 2 28 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.235 $X2=1.13 $Y2=0.57
r174 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends

