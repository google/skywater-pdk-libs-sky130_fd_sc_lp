* File: sky130_fd_sc_lp__or4_4.pex.spice
* Created: Wed Sep  2 10:32:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4_4%D 1 3 6 8 9 10 11
r28 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.375 $X2=0.37 $Y2=1.375
r29 11 16 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.375
r30 10 16 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.375
r31 8 15 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.555 $Y=1.375
+ $X2=0.37 $Y2=1.375
r32 8 9 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.555 $Y=1.375
+ $X2=0.63 $Y2=1.375
r33 4 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.54 $X2=0.63
+ $Y2=1.375
r34 4 6 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.63 $Y=1.54 $X2=0.63
+ $Y2=2.465
r35 1 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.21 $X2=0.63
+ $Y2=1.375
r36 1 3 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.63 $Y=1.21 $X2=0.63
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_4%C 3 7 9 10 14
c38 3 0 6.93714e-20 $X=0.99 $Y=2.465
r39 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=1.51
+ $X2=1.08 $Y2=1.675
r40 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=1.51
+ $X2=1.08 $Y2=1.345
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.51 $X2=1.08 $Y2=1.51
r42 10 15 4.12815 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=1.2 $Y=1.592
+ $X2=1.08 $Y2=1.592
r43 9 15 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=0.72 $Y=1.592
+ $X2=1.08 $Y2=1.592
r44 7 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.06 $Y=0.665
+ $X2=1.06 $Y2=1.345
r45 3 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.99 $Y=2.465
+ $X2=0.99 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_4%B 3 7 9 12 13
c34 13 0 6.93714e-20 $X=1.62 $Y=1.51
c35 3 0 7.73246e-20 $X=1.53 $Y=2.465
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.51
+ $X2=1.62 $Y2=1.675
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.51
+ $X2=1.62 $Y2=1.345
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.51 $X2=1.62 $Y2=1.51
r39 9 13 5.3322 $w=3.33e-07 $l=1.55e-07 $layer=LI1_cond $X=1.662 $Y=1.665
+ $X2=1.662 $Y2=1.51
r40 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.64 $Y=0.665
+ $X2=1.64 $Y2=1.345
r41 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.53 $Y=2.465
+ $X2=1.53 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_4%A 3 7 9 12 13
c40 13 0 7.73246e-20 $X=2.16 $Y=1.51
r41 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.51
+ $X2=2.16 $Y2=1.675
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.51
+ $X2=2.16 $Y2=1.345
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.51 $X2=2.16 $Y2=1.51
r44 9 13 7.00505 $w=2.53e-07 $l=1.55e-07 $layer=LI1_cond $X=2.127 $Y=1.665
+ $X2=2.127 $Y2=1.51
r45 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.07 $Y=2.465
+ $X2=2.07 $Y2=1.675
r46 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.07 $Y=0.665
+ $X2=2.07 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_4%A_58_367# 1 2 3 12 16 20 24 28 32 36 40 42 44
+ 46 50 52 53 56 58 61 63 69 70 74 75
r152 80 81 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.505 $Y=1.51
+ $X2=3.935 $Y2=1.51
r153 79 80 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.075 $Y=1.51
+ $X2=3.505 $Y2=1.51
r154 70 81 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4.095 $Y=1.51
+ $X2=3.935 $Y2=1.51
r155 69 70 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.095
+ $Y=1.51 $X2=4.095 $Y2=1.51
r156 67 79 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.735 $Y=1.51
+ $X2=3.075 $Y2=1.51
r157 67 76 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.735 $Y=1.51
+ $X2=2.645 $Y2=1.51
r158 66 69 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.735 $Y=1.51
+ $X2=4.095 $Y2=1.51
r159 66 67 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.735
+ $Y=1.51 $X2=2.735 $Y2=1.51
r160 64 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.51
+ $X2=2.51 $Y2=1.51
r161 64 66 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.595 $Y=1.51
+ $X2=2.735 $Y2=1.51
r162 62 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.595
+ $X2=2.51 $Y2=1.51
r163 62 63 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.51 $Y=1.595
+ $X2=2.51 $Y2=1.93
r164 61 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.425
+ $X2=2.51 $Y2=1.51
r165 60 61 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.51 $Y=1.165
+ $X2=2.51 $Y2=1.425
r166 59 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=1.08
+ $X2=1.855 $Y2=1.08
r167 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.425 $Y=1.08
+ $X2=2.51 $Y2=1.165
r168 58 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.425 $Y=1.08
+ $X2=2.02 $Y2=1.08
r169 54 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=1.08
r170 54 56 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=0.37
r171 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.69 $Y=1.08
+ $X2=1.855 $Y2=1.08
r172 52 53 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.69 $Y=1.08
+ $X2=1.01 $Y2=1.08
r173 48 53 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.88 $Y=0.995
+ $X2=1.01 $Y2=1.08
r174 48 50 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=0.88 $Y=0.995
+ $X2=0.88 $Y2=0.42
r175 47 73 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=2.015
+ $X2=0.415 $Y2=2.015
r176 46 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.425 $Y=2.015
+ $X2=2.51 $Y2=1.93
r177 46 47 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=2.425 $Y=2.015
+ $X2=0.58 $Y2=2.015
r178 42 73 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=2.1
+ $X2=0.415 $Y2=2.015
r179 42 44 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.415 $Y=2.1
+ $X2=0.415 $Y2=2.95
r180 38 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=1.675
+ $X2=3.935 $Y2=1.51
r181 38 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.935 $Y=1.675
+ $X2=3.935 $Y2=2.465
r182 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=1.345
+ $X2=3.935 $Y2=1.51
r183 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.935 $Y=1.345
+ $X2=3.935 $Y2=0.665
r184 30 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.675
+ $X2=3.505 $Y2=1.51
r185 30 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.505 $Y=1.675
+ $X2=3.505 $Y2=2.465
r186 26 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.345
+ $X2=3.505 $Y2=1.51
r187 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.505 $Y=1.345
+ $X2=3.505 $Y2=0.665
r188 22 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.675
+ $X2=3.075 $Y2=1.51
r189 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.075 $Y=1.675
+ $X2=3.075 $Y2=2.465
r190 18 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.345
+ $X2=3.075 $Y2=1.51
r191 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.075 $Y=1.345
+ $X2=3.075 $Y2=0.665
r192 14 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.675
+ $X2=2.645 $Y2=1.51
r193 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.645 $Y=1.675
+ $X2=2.645 $Y2=2.465
r194 10 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.345
+ $X2=2.645 $Y2=1.51
r195 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.645 $Y=1.345
+ $X2=2.645 $Y2=0.665
r196 3 73 400 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.29
+ $Y=1.835 $X2=0.415 $Y2=2.035
r197 3 44 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.29
+ $Y=1.835 $X2=0.415 $Y2=2.95
r198 2 56 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.715
+ $Y=0.245 $X2=1.855 $Y2=0.37
r199 1 50 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.705
+ $Y=0.245 $X2=0.845 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_4%VPWR 1 2 3 12 16 22 27 28 30 31 32 44 50 51 54
r55 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 51 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 48 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.15 $Y2=3.33
r59 48 50 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.56 $Y2=3.33
r60 47 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 44 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.15 $Y2=3.33
r63 44 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 43 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r65 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r67 36 40 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r68 35 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 32 43 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r71 32 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 30 42 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=3.29 $Y2=3.33
r74 29 46 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.455 $Y=3.33
+ $X2=3.6 $Y2=3.33
r75 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=3.33
+ $X2=3.29 $Y2=3.33
r76 27 39 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.35 $Y2=3.33
r78 26 42 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.35 $Y2=3.33
r80 22 25 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.15 $Y=2.19
+ $X2=4.15 $Y2=2.95
r81 20 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=3.33
r82 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=2.95
r83 16 19 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=3.29 $Y=2.19
+ $X2=3.29 $Y2=2.97
r84 14 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=3.245
+ $X2=3.29 $Y2=3.33
r85 14 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.29 $Y=3.245
+ $X2=3.29 $Y2=2.97
r86 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=3.245
+ $X2=2.35 $Y2=3.33
r87 10 12 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=2.35 $Y=3.245
+ $X2=2.35 $Y2=2.395
r88 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.835 $X2=4.15 $Y2=2.95
r89 3 22 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.835 $X2=4.15 $Y2=2.19
r90 2 19 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=2.97
r91 2 16 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=2.19
r92 1 12 300 $w=1.7e-07 $l=6.54523e-07 $layer=licon1_PDIFF $count=2 $X=2.145
+ $Y=1.835 $X2=2.35 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41 42
+ 44 45 46 47 61
r65 59 61 1.61746 $w=2.83e-07 $l=4e-08 $layer=LI1_cond $X=4.572 $Y=1.255
+ $X2=4.572 $Y2=1.295
r66 46 53 3.43356 $w=2.72e-07 $l=9.12688e-08 $layer=LI1_cond $X=4.572 $Y=1.17
+ $X2=4.585 $Y2=1.085
r67 46 59 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=4.572 $Y=1.17
+ $X2=4.572 $Y2=1.255
r68 46 47 14.0719 $w=2.83e-07 $l=3.48e-07 $layer=LI1_cond $X=4.572 $Y=1.317
+ $X2=4.572 $Y2=1.665
r69 46 61 0.889605 $w=2.83e-07 $l=2.2e-08 $layer=LI1_cond $X=4.572 $Y=1.317
+ $X2=4.572 $Y2=1.295
r70 45 53 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=4.585 $Y=0.925
+ $X2=4.585 $Y2=1.085
r71 44 45 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=4.585 $Y=0.555
+ $X2=4.585 $Y2=0.925
r72 43 47 4.04366 $w=2.83e-07 $l=1e-07 $layer=LI1_cond $X=4.572 $Y=1.765
+ $X2=4.572 $Y2=1.665
r73 40 41 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.85 $Y=1.17
+ $X2=3.737 $Y2=1.17
r74 39 46 3.08518 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.43 $Y=1.17
+ $X2=4.572 $Y2=1.17
r75 39 40 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.43 $Y=1.17
+ $X2=3.85 $Y2=1.17
r76 38 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.815 $Y=1.85
+ $X2=3.72 $Y2=1.85
r77 37 43 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=4.43 $Y=1.85
+ $X2=4.572 $Y2=1.765
r78 37 38 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.43 $Y=1.85
+ $X2=3.815 $Y2=1.85
r79 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.72 $Y=1.98
+ $X2=3.72 $Y2=2.91
r80 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.935
+ $X2=3.72 $Y2=1.85
r81 31 33 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=3.72 $Y=1.935
+ $X2=3.72 $Y2=1.98
r82 27 41 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.737 $Y=1.085
+ $X2=3.737 $Y2=1.17
r83 27 29 34.0611 $w=2.23e-07 $l=6.65e-07 $layer=LI1_cond $X=3.737 $Y=1.085
+ $X2=3.737 $Y2=0.42
r84 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.625 $Y=1.85
+ $X2=3.72 $Y2=1.85
r85 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.625 $Y=1.85
+ $X2=2.955 $Y2=1.85
r86 23 41 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.625 $Y=1.17
+ $X2=3.737 $Y2=1.17
r87 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.625 $Y=1.17
+ $X2=2.955 $Y2=1.17
r88 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.86 $Y=1.98
+ $X2=2.86 $Y2=2.91
r89 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.86 $Y=1.935
+ $X2=2.955 $Y2=1.85
r90 17 19 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=2.86 $Y=1.935
+ $X2=2.86 $Y2=1.98
r91 13 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.86 $Y=1.085
+ $X2=2.955 $Y2=1.17
r92 13 15 38.8182 $w=1.88e-07 $l=6.65e-07 $layer=LI1_cond $X=2.86 $Y=1.085
+ $X2=2.86 $Y2=0.42
r93 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=2.91
r94 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=1.98
r95 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.91
r96 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=1.98
r97 2 29 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.58
+ $Y=0.245 $X2=3.72 $Y2=0.42
r98 1 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.72
+ $Y=0.245 $X2=2.86 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_4%VGND 1 2 3 4 5 16 18 20 24 28 32 34 38 41 42
+ 43 44 45 56 57 63 66
r66 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r67 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r69 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r70 57 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r71 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r72 54 66 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.152
+ $Y2=0
r73 54 56 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.56
+ $Y2=0
r74 53 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r75 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r76 50 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r77 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.355
+ $Y2=0
r79 47 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=2.16
+ $Y2=0
r80 45 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r81 45 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r82 43 52 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.12
+ $Y2=0
r83 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.29
+ $Y2=0
r84 41 49 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.16
+ $Y2=0
r85 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.355
+ $Y2=0
r86 40 52 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.52 $Y=0 $X2=3.12
+ $Y2=0
r87 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.52 $Y=0 $X2=2.355
+ $Y2=0
r88 36 66 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.152 $Y=0.085
+ $X2=4.152 $Y2=0
r89 36 38 13.264 $w=2.63e-07 $l=3.05e-07 $layer=LI1_cond $X=4.152 $Y=0.085
+ $X2=4.152 $Y2=0.39
r90 35 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.29
+ $Y2=0
r91 34 66 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.152
+ $Y2=0
r92 34 35 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=3.455
+ $Y2=0
r93 30 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0
r94 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0.39
r95 26 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=0.085
+ $X2=2.355 $Y2=0
r96 26 28 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=0.085
+ $X2=2.355 $Y2=0.37
r97 22 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=0.085
+ $X2=1.355 $Y2=0
r98 22 24 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.355 $Y=0.085
+ $X2=1.355 $Y2=0.37
r99 21 60 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.29
+ $Y2=0
r100 20 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=1.355
+ $Y2=0
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=0.58
+ $Y2=0
r102 16 60 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.29 $Y2=0
r103 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.415 $Y2=0.39
r104 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.01
+ $Y=0.245 $X2=4.15 $Y2=0.39
r105 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.245 $X2=3.29 $Y2=0.39
r106 3 28 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=2.145
+ $Y=0.245 $X2=2.355 $Y2=0.37
r107 2 24 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=1.135
+ $Y=0.245 $X2=1.355 $Y2=0.37
r108 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.29
+ $Y=0.245 $X2=0.415 $Y2=0.39
.ends

