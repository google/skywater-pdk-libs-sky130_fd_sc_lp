* File: sky130_fd_sc_lp__mux4_lp.spice
* Created: Wed Sep  2 10:02:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux4_lp.pex.spice"
.subckt sky130_fd_sc_lp__mux4_lp  VNB VPB S1 A3 S0 A2 A1 A0 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A0	A0
* A1	A1
* A2	A2
* S0	S0
* A3	A3
* S1	S1
* VPB	VPB
* VNB	VNB
MM1006 A_114_47# N_A_84_21#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_84_21#_M1026_g A_114_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_A_84_21#_M1016_d N_S1_M1016_g N_A_245_411#_M1016_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_470_57#_M1025_d N_A_320_366#_M1025_g N_A_84_21#_M1016_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_684_101# N_S1_M1017_g N_A_320_366#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1533 PD=0.63 PS=1.57 NRD=14.28 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_S1_M1007_g A_684_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.13545 AS=0.0441 PD=1.065 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1027 A_915_101# N_A3_M1027_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.13545 PD=0.745 PS=1.065 NRD=30.708 NRS=104.28 M=1 R=2.8
+ SA=75001.4 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_245_411#_M1003_d N_S0_M1003_g A_915_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.099225 AS=0.06825 PD=1.05 PS=0.745 NRD=0 NRS=30.708 M=1 R=2.8 SA=75001.9
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 A_1112_47# N_A_946_317#_M1011_g N_A_245_411#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.099225 PD=0.66 PS=1.05 NRD=18.564 NRS=51.78 M=1 R=2.8
+ SA=75001 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A2_M1012_g A_1112_47# VNB NSHORT L=0.15 W=0.42 AD=0.2037
+ AS=0.0504 PD=1.39 PS=0.66 NRD=174.276 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1018 A_1414_47# N_A1_M1018_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.2037 PD=0.66 PS=1.39 NRD=18.564 NRS=22.848 M=1 R=2.8 SA=75002.5
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1019 N_A_470_57#_M1019_d N_S0_M1019_g A_1414_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=31.428 NRS=18.564 M=1 R=2.8 SA=75002.9
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1024 A_1600_47# N_A_946_317#_M1024_g N_A_470_57#_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1512 AS=0.0819 PD=1.14 PS=0.81 NRD=87.132 NRS=0 M=1 R=2.8
+ SA=75003.4 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A0_M1000_g A_1600_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1512 PD=0.7 PS=1.14 NRD=0 NRS=87.132 M=1 R=2.8 SA=75004.3 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1014 A_1860_47# N_S0_M1014_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1020 N_A_946_317#_M1020_d N_S0_M1020_g A_1860_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75005.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_84_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1013 N_A_84_21#_M1013_d N_A_320_366#_M1013_g N_A_245_411#_M1013_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.2375 AS=0.375 PD=1.475 PS=2.75 NRD=15.7403 NRS=17.73 M=1 R=4
+ SA=125000 SB=125001 A=0.25 P=2.5 MULT=1
MM1001 N_A_470_57#_M1001_d N_S1_M1001_g N_A_84_21#_M1013_d VPB PHIGHVT L=0.25
+ W=1 AD=0.34 AS=0.2375 PD=2.68 PS=1.475 NRD=10.8153 NRS=22.6353 M=1 R=4
+ SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1022 N_VPWR_M1022_d N_S1_M1022_g N_A_320_366#_M1022_s VPB PHIGHVT L=0.25 W=1
+ AD=0.2316 AS=0.4868 PD=1.52 PS=3.57 NRD=16.7253 NRS=85.0449 M=1 R=4 SA=125000
+ SB=125006 A=0.25 P=2.5 MULT=1
MM1002 A_898_419# N_A3_M1002_g N_VPWR_M1022_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.2316 PD=1.24 PS=1.52 NRD=12.7853 NRS=16.7253 M=1 R=4 SA=125001 SB=125005
+ A=0.25 P=2.5 MULT=1
MM1015 N_A_245_411#_M1015_d N_A_946_317#_M1015_g A_898_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.41 AS=0.12 PD=1.82 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125005 A=0.25 P=2.5 MULT=1
MM1008 A_1210_419# N_S0_M1008_g N_A_245_411#_M1015_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1525 AS=0.41 PD=1.305 PS=1.82 NRD=19.1878 NRS=106.36 M=1 R=4 SA=125002
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A2_M1009_g A_1210_419# VPB PHIGHVT L=0.25 W=1 AD=0.155
+ AS=0.1525 PD=1.31 PS=1.305 NRD=0 NRS=19.1878 M=1 R=4 SA=125003 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1010 A_1433_419# N_A1_M1010_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.155 PD=1.24 PS=1.31 NRD=12.7853 NRS=5.8903 M=1 R=4 SA=125004 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1023 N_A_470_57#_M1023_d N_A_946_317#_M1023_g A_1433_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.2833 AS=0.12 PD=1.595 PS=1.24 NRD=15.7403 NRS=12.7853 M=1 R=4
+ SA=125004 SB=125002 A=0.25 P=2.5 MULT=1
MM1004 A_1692_419# N_S0_M1004_g N_A_470_57#_M1023_d VPB PHIGHVT L=0.25 W=1
+ AD=0.145 AS=0.2833 PD=1.29 PS=1.595 NRD=17.7103 NRS=38.3953 M=1 R=4 SA=125005
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1021 N_VPWR_M1021_d N_A0_M1021_g A_1692_419# VPB PHIGHVT L=0.25 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=1.9503 NRS=17.7103 M=1 R=4 SA=125005 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1028 N_A_946_317#_M1028_d N_S0_M1028_g N_VPWR_M1021_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.145 PD=2.57 PS=1.29 NRD=0 NRS=0 M=1 R=4 SA=125006 SB=125000
+ A=0.25 P=2.5 MULT=1
DX29_noxref VNB VPB NWDIODE A=19.6423 P=24.97
c_128 VNB 0 1.01928e-19 $X=0 $Y=0
c_1542 A_1433_419# 0 1.3249e-19 $X=7.165 $Y=2.095
*
.include "sky130_fd_sc_lp__mux4_lp.pxi.spice"
*
.ends
*
*
