* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VGND B1 a_157_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_832_21# A2_N a_1241_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_157_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_73_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR B2 a_73_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR A1_N a_1241_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_1241_367# A2_N a_832_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 Y B2 a_157_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND a_832_21# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_73_367# a_832_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_73_367# a_832_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND A1_N a_832_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR B1 a_73_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND B1 a_157_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VGND a_832_21# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_157_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_832_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR B2 a_73_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_73_367# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_832_21# A2_N a_1241_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR B1 a_73_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_157_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 Y B2 a_157_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Y a_832_21# a_73_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 Y a_832_21# a_73_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 Y a_832_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VGND A2_N a_832_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_73_367# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_1241_367# A2_N a_832_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_1241_367# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 Y a_832_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_832_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_157_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 VGND A2_N a_832_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_73_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 a_1241_367# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 a_832_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 VPWR A1_N a_1241_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 VGND A1_N a_832_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 a_832_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
