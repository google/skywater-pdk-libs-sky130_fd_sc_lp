* File: sky130_fd_sc_lp__xor2_1.pxi.spice
* Created: Fri Aug 28 11:36:13 2020
* 
x_PM_SKY130_FD_SC_LP__XOR2_1%B N_B_c_62_n N_B_M1008_g N_B_M1001_g N_B_M1003_g
+ N_B_M1004_g N_B_c_65_n N_B_c_66_n N_B_c_72_n N_B_c_67_n N_B_c_68_n B B
+ N_B_c_76_n B PM_SKY130_FD_SC_LP__XOR2_1%B
x_PM_SKY130_FD_SC_LP__XOR2_1%A N_A_M1006_g N_A_c_151_n N_A_M1009_g N_A_M1007_g
+ N_A_c_153_n N_A_M1002_g A A A N_A_c_155_n PM_SKY130_FD_SC_LP__XOR2_1%A
x_PM_SKY130_FD_SC_LP__XOR2_1%A_42_367# N_A_42_367#_M1008_d N_A_42_367#_M1001_s
+ N_A_42_367#_c_201_n N_A_42_367#_M1000_g N_A_42_367#_c_202_n
+ N_A_42_367#_M1005_g N_A_42_367#_c_213_n N_A_42_367#_c_214_n
+ N_A_42_367#_c_226_n N_A_42_367#_c_229_n N_A_42_367#_c_204_n
+ N_A_42_367#_c_231_n N_A_42_367#_c_232_n N_A_42_367#_c_205_n
+ N_A_42_367#_c_206_n N_A_42_367#_c_215_n N_A_42_367#_c_207_n
+ N_A_42_367#_c_208_n N_A_42_367#_c_237_n N_A_42_367#_c_209_n
+ N_A_42_367#_c_210_n N_A_42_367#_c_211_n PM_SKY130_FD_SC_LP__XOR2_1%A_42_367#
x_PM_SKY130_FD_SC_LP__XOR2_1%VPWR N_VPWR_M1006_d N_VPWR_M1004_d N_VPWR_c_313_n
+ N_VPWR_c_314_n N_VPWR_c_315_n VPWR N_VPWR_c_316_n N_VPWR_c_317_n
+ N_VPWR_c_312_n N_VPWR_c_319_n PM_SKY130_FD_SC_LP__XOR2_1%VPWR
x_PM_SKY130_FD_SC_LP__XOR2_1%A_293_367# N_A_293_367#_M1007_d
+ N_A_293_367#_M1005_d N_A_293_367#_c_360_n N_A_293_367#_c_364_n
+ N_A_293_367#_c_361_n PM_SKY130_FD_SC_LP__XOR2_1%A_293_367#
x_PM_SKY130_FD_SC_LP__XOR2_1%X N_X_M1003_d N_X_M1005_s N_X_c_390_n N_X_c_396_n X
+ PM_SKY130_FD_SC_LP__XOR2_1%X
x_PM_SKY130_FD_SC_LP__XOR2_1%VGND N_VGND_M1008_s N_VGND_M1009_d N_VGND_M1000_d
+ N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n
+ VGND N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n
+ PM_SKY130_FD_SC_LP__XOR2_1%VGND
cc_1 VNB N_B_c_62_n 0.0188568f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.295
cc_2 VNB N_B_M1001_g 0.00158573f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_3 VNB N_B_M1003_g 0.0206262f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.765
cc_4 VNB N_B_c_65_n 0.0419246f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_5 VNB N_B_c_66_n 0.00908743f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.46
cc_6 VNB N_B_c_67_n 0.00486247f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.51
cc_7 VNB N_B_c_68_n 0.0376929f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.51
cc_8 VNB B 0.0245085f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A_M1006_g 0.0015007f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.765
cc_10 VNB N_A_c_151_n 0.0159414f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_11 VNB N_A_M1007_g 0.00152408f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.765
cc_12 VNB N_A_c_153_n 0.0155429f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.675
cc_13 VNB A 0.0116868f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.46
cc_14 VNB N_A_c_155_n 0.0412846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_42_367#_c_201_n 0.0208696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_42_367#_c_202_n 0.0095374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_42_367#_M1005_g 0.00189699f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=2.465
cc_18 VNB N_A_42_367#_c_204_n 0.00202722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_42_367#_c_205_n 0.00710512f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_20 VNB N_A_42_367#_c_206_n 8.92719e-19 $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_21 VNB N_A_42_367#_c_207_n 0.0017594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_42_367#_c_208_n 0.0012087f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.51
cc_23 VNB N_A_42_367#_c_209_n 0.0263893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_42_367#_c_210_n 0.0496187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_42_367#_c_211_n 0.0140741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_312_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_390_n 0.0079052f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.345
cc_28 VNB X 0.00456676f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=2.465
cc_29 VNB N_VGND_c_422_n 0.0126248f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.765
cc_30 VNB N_VGND_c_423_n 0.0366605f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.675
cc_31 VNB N_VGND_c_424_n 0.00278994f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_32 VNB N_VGND_c_425_n 0.011635f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.81
cc_33 VNB N_VGND_c_426_n 0.0378088f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.725
cc_34 VNB N_VGND_c_427_n 0.0166314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_428_n 0.0400766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_429_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_430_n 0.219287f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_38 VPB N_B_M1001_g 0.0230759f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.465
cc_39 VPB N_B_M1004_g 0.0224119f $X=-0.19 $Y=1.655 $X2=1.82 $Y2=2.465
cc_40 VPB N_B_c_72_n 0.00848067f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.81
cc_41 VPB N_B_c_67_n 8.2756e-19 $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.51
cc_42 VPB N_B_c_68_n 0.0110481f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.51
cc_43 VPB B 0.00329297f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_44 VPB N_B_c_76_n 0.0112332f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.725
cc_45 VPB N_A_M1006_g 0.0185601f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.765
cc_46 VPB N_A_M1007_g 0.019258f $X=-0.19 $Y=1.655 $X2=1.8 $Y2=0.765
cc_47 VPB N_A_42_367#_M1005_g 0.0269486f $X=-0.19 $Y=1.655 $X2=1.82 $Y2=2.465
cc_48 VPB N_A_42_367#_c_213_n 0.00745873f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.46
cc_49 VPB N_A_42_367#_c_214_n 0.0327625f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.81
cc_50 VPB N_A_42_367#_c_215_n 0.0155808f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_51 VPB N_A_42_367#_c_208_n 0.021493f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.51
cc_52 VPB N_VPWR_c_313_n 0.00251047f $X=-0.19 $Y=1.655 $X2=1.8 $Y2=0.765
cc_53 VPB N_VPWR_c_314_n 0.0293871f $X=-0.19 $Y=1.655 $X2=1.82 $Y2=1.675
cc_54 VPB N_VPWR_c_315_n 0.00414335f $X=-0.19 $Y=1.655 $X2=1.82 $Y2=2.465
cc_55 VPB N_VPWR_c_316_n 0.0178035f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=1.725
cc_56 VPB N_VPWR_c_317_n 0.0306123f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_57 VPB N_VPWR_c_312_n 0.050363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_319_n 0.0142123f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_59 VPB N_A_293_367#_c_360_n 0.00724251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_293_367#_c_361_n 0.015084f $X=-0.19 $Y=1.655 $X2=1.82 $Y2=2.465
cc_61 VPB X 0.0115599f $X=-0.19 $Y=1.655 $X2=1.82 $Y2=2.465
cc_62 N_B_M1001_g N_A_M1006_g 0.084263f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_63 N_B_c_72_n N_A_M1006_g 0.0103161f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_64 N_B_c_62_n N_A_c_151_n 0.0150394f $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_65 N_B_M1004_g N_A_M1007_g 0.0387159f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_66 N_B_c_72_n N_A_M1007_g 0.010566f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_67 N_B_c_67_n N_A_M1007_g 2.10386e-19 $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_68 N_B_c_68_n N_A_M1007_g 0.00273475f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_69 N_B_M1003_g N_A_c_153_n 0.0564963f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_70 N_B_c_62_n A 0.00312863f $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_71 N_B_M1003_g A 0.00448239f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_72 N_B_c_72_n A 0.0865599f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_73 N_B_c_67_n A 0.0159835f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_74 N_B_c_68_n A 0.00622761f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_75 B A 0.027914f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B_M1003_g N_A_c_155_n 0.0210318f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_77 N_B_c_66_n N_A_c_155_n 0.0222729f $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_78 N_B_c_72_n N_A_c_155_n 0.00488238f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_79 N_B_c_67_n N_A_c_155_n 4.76257e-19 $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_80 B N_A_c_155_n 5.4586e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_B_c_76_n N_A_42_367#_M1001_s 0.00258458f $X=0.27 $Y=1.725 $X2=0 $Y2=0
cc_82 N_B_M1003_g N_A_42_367#_c_201_n 0.0157614f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_83 N_B_c_68_n N_A_42_367#_c_202_n 0.00477363f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_84 N_B_c_72_n N_A_42_367#_M1005_g 3.26904e-19 $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_85 N_B_M1001_g N_A_42_367#_c_213_n 7.32094e-19 $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_c_65_n N_A_42_367#_c_213_n 0.00117599f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_87 N_B_c_72_n N_A_42_367#_c_213_n 0.00186226f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_88 N_B_c_76_n N_A_42_367#_c_213_n 0.0225137f $X=0.27 $Y=1.725 $X2=0 $Y2=0
cc_89 N_B_M1001_g N_A_42_367#_c_214_n 0.0142963f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_90 N_B_M1001_g N_A_42_367#_c_226_n 0.0108536f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_A_42_367#_c_226_n 0.011714f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_92 N_B_c_72_n N_A_42_367#_c_226_n 0.0736585f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_93 N_B_c_62_n N_A_42_367#_c_229_n 0.00301723f $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_94 N_B_c_62_n N_A_42_367#_c_204_n 0.00661374f $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_95 N_B_M1003_g N_A_42_367#_c_231_n 0.0108833f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_96 N_B_M1003_g N_A_42_367#_c_232_n 0.0113328f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_97 N_B_M1003_g N_A_42_367#_c_205_n 0.00325562f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_98 N_B_M1003_g N_A_42_367#_c_206_n 0.00361471f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_99 N_B_c_72_n N_A_42_367#_c_215_n 2.40539e-19 $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_100 N_B_c_68_n N_A_42_367#_c_215_n 0.00201699f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_101 N_B_c_72_n N_A_42_367#_c_237_n 0.0132447f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_102 N_B_c_68_n N_A_42_367#_c_237_n 7.35175e-19 $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_c_68_n N_A_42_367#_c_210_n 0.00286745f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_104 N_B_c_72_n A_125_367# 0.00134267f $X=1.935 $Y=1.81 $X2=-0.19 $Y2=-0.245
cc_105 N_B_c_72_n N_VPWR_M1006_d 0.00198204f $X=1.935 $Y=1.81 $X2=-0.19
+ $Y2=-0.245
cc_106 N_B_c_72_n N_VPWR_M1004_d 0.00271869f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_107 N_B_M1001_g N_VPWR_c_313_n 0.00307183f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B_M1001_g N_VPWR_c_314_n 0.0054895f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_109 N_B_M1004_g N_VPWR_c_316_n 0.00409076f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_110 N_B_M1001_g N_VPWR_c_312_n 0.0109356f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_111 N_B_M1004_g N_VPWR_c_312_n 0.00709144f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B_M1004_g N_VPWR_c_319_n 0.0087173f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B_c_72_n N_A_293_367#_M1007_d 0.00176891f $X=1.935 $Y=1.81 $X2=-0.19
+ $Y2=-0.245
cc_114 N_B_M1004_g N_A_293_367#_c_360_n 0.0116867f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B_M1004_g N_A_293_367#_c_364_n 0.0188776f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B_M1003_g N_X_c_390_n 0.00183937f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_117 N_B_c_67_n N_X_c_390_n 0.016121f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_118 N_B_c_68_n N_X_c_390_n 0.00227487f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_119 N_B_M1003_g N_X_c_396_n 0.00744433f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_120 N_B_c_67_n N_X_c_396_n 0.00592675f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_121 N_B_c_68_n N_X_c_396_n 0.00402209f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_122 N_B_M1004_g X 0.00486041f $X=1.82 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B_c_72_n X 0.00932626f $X=1.935 $Y=1.81 $X2=0 $Y2=0
cc_124 N_B_c_67_n X 0.0122686f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_125 N_B_c_68_n X 0.00136561f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_126 N_B_c_62_n N_VGND_c_423_n 0.00351453f $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_127 N_B_c_65_n N_VGND_c_423_n 0.00161388f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_128 B N_VGND_c_423_n 0.0233037f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B_c_62_n N_VGND_c_424_n 4.86336e-19 $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_130 N_B_M1003_g N_VGND_c_424_n 7.55247e-19 $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_131 N_B_c_62_n N_VGND_c_427_n 0.00453633f $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_132 N_B_M1003_g N_VGND_c_428_n 0.00291319f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_133 N_B_c_62_n N_VGND_c_430_n 0.00882554f $X=0.55 $Y=1.295 $X2=0 $Y2=0
cc_134 N_B_M1003_g N_VGND_c_430_n 0.00410425f $X=1.8 $Y=0.765 $X2=0 $Y2=0
cc_135 N_A_M1006_g N_A_42_367#_c_214_n 0.00273619f $X=0.94 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_M1006_g N_A_42_367#_c_226_n 0.0141633f $X=0.94 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_M1007_g N_A_42_367#_c_226_n 0.0144132f $X=1.39 $Y=2.465 $X2=0 $Y2=0
cc_138 A N_A_42_367#_c_229_n 0.0173818f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A_c_151_n N_A_42_367#_c_204_n 3.5044e-19 $X=0.98 $Y=1.295 $X2=0 $Y2=0
cc_140 N_A_c_151_n N_A_42_367#_c_231_n 0.012081f $X=0.98 $Y=1.295 $X2=0 $Y2=0
cc_141 N_A_c_153_n N_A_42_367#_c_231_n 0.0138635f $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_142 A N_A_42_367#_c_231_n 0.0589612f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A_c_155_n N_A_42_367#_c_231_n 5.63199e-19 $X=1.41 $Y=1.46 $X2=0 $Y2=0
cc_144 N_A_c_153_n N_A_42_367#_c_206_n 9.18629e-19 $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_145 N_A_M1006_g N_VPWR_c_313_n 0.0163675f $X=0.94 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1007_g N_VPWR_c_313_n 0.00294729f $X=1.39 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1006_g N_VPWR_c_314_n 0.00486043f $X=0.94 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_M1007_g N_VPWR_c_316_n 0.0054895f $X=1.39 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_VPWR_c_312_n 0.00827383f $X=0.94 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_VPWR_c_312_n 0.00984228f $X=1.39 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_M1007_g N_A_293_367#_c_364_n 0.0081466f $X=1.39 $Y=2.465 $X2=0 $Y2=0
cc_152 A N_X_c_390_n 0.00456373f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A_c_151_n N_VGND_c_424_n 0.00858164f $X=0.98 $Y=1.295 $X2=0 $Y2=0
cc_154 N_A_c_153_n N_VGND_c_424_n 0.00974467f $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_155 N_A_c_151_n N_VGND_c_427_n 0.00400407f $X=0.98 $Y=1.295 $X2=0 $Y2=0
cc_156 N_A_c_153_n N_VGND_c_428_n 0.00400407f $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_157 N_A_c_151_n N_VGND_c_430_n 0.00775088f $X=0.98 $Y=1.295 $X2=0 $Y2=0
cc_158 N_A_c_153_n N_VGND_c_430_n 0.00772763f $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_159 N_A_42_367#_c_226_n A_125_367# 0.00615027f $X=1.94 $Y=2.15 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_42_367#_c_226_n N_VPWR_M1006_d 0.00379439f $X=1.94 $Y=2.15 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_42_367#_c_215_n N_VPWR_M1004_d 0.00689232f $X=3.065 $Y=2.32 $X2=0
+ $Y2=0
cc_162 N_A_42_367#_c_237_n N_VPWR_M1004_d 0.0108213f $X=2.025 $Y=2.15 $X2=0
+ $Y2=0
cc_163 N_A_42_367#_c_214_n N_VPWR_c_313_n 0.0209623f $X=0.335 $Y=2.91 $X2=0
+ $Y2=0
cc_164 N_A_42_367#_c_226_n N_VPWR_c_313_n 0.0169188f $X=1.94 $Y=2.15 $X2=0 $Y2=0
cc_165 N_A_42_367#_c_214_n N_VPWR_c_314_n 0.0210467f $X=0.335 $Y=2.91 $X2=0
+ $Y2=0
cc_166 N_A_42_367#_M1005_g N_VPWR_c_317_n 0.0041378f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_42_367#_M1001_s N_VPWR_c_312_n 0.00215158f $X=0.21 $Y=1.835 $X2=0
+ $Y2=0
cc_168 N_A_42_367#_M1005_g N_VPWR_c_312_n 0.00824063f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_42_367#_c_214_n N_VPWR_c_312_n 0.0125689f $X=0.335 $Y=2.91 $X2=0
+ $Y2=0
cc_170 N_A_42_367#_M1005_g N_VPWR_c_319_n 0.00645297f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_42_367#_c_226_n N_A_293_367#_M1007_d 0.00353353f $X=1.94 $Y=2.15
+ $X2=-0.19 $Y2=-0.245
cc_172 N_A_42_367#_c_215_n N_A_293_367#_M1005_d 0.003826f $X=3.065 $Y=2.32 $X2=0
+ $Y2=0
cc_173 N_A_42_367#_c_208_n N_A_293_367#_M1005_d 0.0067942f $X=3.15 $Y=2.235
+ $X2=0 $Y2=0
cc_174 N_A_42_367#_M1005_g N_A_293_367#_c_360_n 0.0109325f $X=2.885 $Y=2.465
+ $X2=0 $Y2=0
cc_175 N_A_42_367#_c_226_n N_A_293_367#_c_360_n 0.00486113f $X=1.94 $Y=2.15
+ $X2=0 $Y2=0
cc_176 N_A_42_367#_c_215_n N_A_293_367#_c_360_n 0.055896f $X=3.065 $Y=2.32 $X2=0
+ $Y2=0
cc_177 N_A_42_367#_c_237_n N_A_293_367#_c_360_n 0.0120849f $X=2.025 $Y=2.15
+ $X2=0 $Y2=0
cc_178 N_A_42_367#_c_226_n N_A_293_367#_c_364_n 0.017057f $X=1.94 $Y=2.15 $X2=0
+ $Y2=0
cc_179 N_A_42_367#_M1005_g N_A_293_367#_c_361_n 0.00919175f $X=2.885 $Y=2.465
+ $X2=0 $Y2=0
cc_180 N_A_42_367#_c_215_n N_A_293_367#_c_361_n 0.0199094f $X=3.065 $Y=2.32
+ $X2=0 $Y2=0
cc_181 N_A_42_367#_c_205_n N_X_M1003_d 0.00891592f $X=2.625 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_42_367#_c_215_n N_X_M1005_s 0.00582966f $X=3.065 $Y=2.32 $X2=0 $Y2=0
cc_183 N_A_42_367#_c_201_n N_X_c_390_n 0.00823363f $X=2.53 $Y=1.295 $X2=0 $Y2=0
cc_184 N_A_42_367#_c_207_n N_X_c_390_n 0.00327316f $X=2.71 $Y=1.23 $X2=0 $Y2=0
cc_185 N_A_42_367#_c_209_n N_X_c_390_n 0.019902f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_186 N_A_42_367#_c_210_n N_X_c_390_n 0.00119782f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_187 N_A_42_367#_c_231_n N_X_c_396_n 0.0142468f $X=1.7 $Y=0.955 $X2=0 $Y2=0
cc_188 N_A_42_367#_c_232_n N_X_c_396_n 0.0206978f $X=1.785 $Y=0.87 $X2=0 $Y2=0
cc_189 N_A_42_367#_c_205_n N_X_c_396_n 0.0269225f $X=2.625 $Y=0.34 $X2=0 $Y2=0
cc_190 N_A_42_367#_c_202_n X 0.0101612f $X=2.605 $Y=1.37 $X2=0 $Y2=0
cc_191 N_A_42_367#_M1005_g X 0.0049892f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A_42_367#_c_215_n X 0.0301594f $X=3.065 $Y=2.32 $X2=0 $Y2=0
cc_193 N_A_42_367#_c_208_n X 0.0244972f $X=3.15 $Y=2.235 $X2=0 $Y2=0
cc_194 N_A_42_367#_c_209_n X 0.0181886f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_195 N_A_42_367#_c_210_n X 0.00433895f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_196 N_A_42_367#_c_211_n X 0.00131192f $X=2.81 $Y=1.46 $X2=0 $Y2=0
cc_197 N_A_42_367#_c_231_n N_VGND_M1009_d 0.00333177f $X=1.7 $Y=0.955 $X2=0
+ $Y2=0
cc_198 N_A_42_367#_c_205_n N_VGND_M1000_d 9.31758e-19 $X=2.625 $Y=0.34 $X2=0
+ $Y2=0
cc_199 N_A_42_367#_c_207_n N_VGND_M1000_d 0.0153476f $X=2.71 $Y=1.23 $X2=0 $Y2=0
cc_200 N_A_42_367#_c_204_n N_VGND_c_423_n 0.0196794f $X=0.765 $Y=0.5 $X2=0 $Y2=0
cc_201 N_A_42_367#_c_204_n N_VGND_c_424_n 0.0140568f $X=0.765 $Y=0.5 $X2=0 $Y2=0
cc_202 N_A_42_367#_c_231_n N_VGND_c_424_n 0.0170777f $X=1.7 $Y=0.955 $X2=0 $Y2=0
cc_203 N_A_42_367#_c_206_n N_VGND_c_424_n 0.00622828f $X=1.87 $Y=0.34 $X2=0
+ $Y2=0
cc_204 N_A_42_367#_c_201_n N_VGND_c_426_n 0.0027687f $X=2.53 $Y=1.295 $X2=0
+ $Y2=0
cc_205 N_A_42_367#_c_205_n N_VGND_c_426_n 0.0144885f $X=2.625 $Y=0.34 $X2=0
+ $Y2=0
cc_206 N_A_42_367#_c_207_n N_VGND_c_426_n 0.047457f $X=2.71 $Y=1.23 $X2=0 $Y2=0
cc_207 N_A_42_367#_c_209_n N_VGND_c_426_n 0.0225031f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_208 N_A_42_367#_c_210_n N_VGND_c_426_n 0.00165489f $X=3.07 $Y=1.46 $X2=0
+ $Y2=0
cc_209 N_A_42_367#_c_204_n N_VGND_c_427_n 0.0122069f $X=0.765 $Y=0.5 $X2=0 $Y2=0
cc_210 N_A_42_367#_c_201_n N_VGND_c_428_n 0.0029147f $X=2.53 $Y=1.295 $X2=0
+ $Y2=0
cc_211 N_A_42_367#_c_205_n N_VGND_c_428_n 0.060316f $X=2.625 $Y=0.34 $X2=0 $Y2=0
cc_212 N_A_42_367#_c_206_n N_VGND_c_428_n 0.0116772f $X=1.87 $Y=0.34 $X2=0 $Y2=0
cc_213 N_A_42_367#_c_201_n N_VGND_c_430_n 0.00442169f $X=2.53 $Y=1.295 $X2=0
+ $Y2=0
cc_214 N_A_42_367#_c_204_n N_VGND_c_430_n 0.00951044f $X=0.765 $Y=0.5 $X2=0
+ $Y2=0
cc_215 N_A_42_367#_c_205_n N_VGND_c_430_n 0.0342827f $X=2.625 $Y=0.34 $X2=0
+ $Y2=0
cc_216 N_A_42_367#_c_206_n N_VGND_c_430_n 0.00594574f $X=1.87 $Y=0.34 $X2=0
+ $Y2=0
cc_217 N_A_42_367#_c_231_n A_297_69# 0.00615027f $X=1.7 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_218 A_125_367# N_VPWR_c_312_n 0.010279f $X=0.625 $Y=1.835 $X2=0 $Y2=0
cc_219 N_VPWR_c_312_n N_A_293_367#_M1007_d 0.00223559f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_220 N_VPWR_c_312_n N_A_293_367#_M1005_d 0.00235821f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_221 N_VPWR_M1004_d N_A_293_367#_c_360_n 0.00802286f $X=1.895 $Y=1.835 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_316_n N_A_293_367#_c_360_n 0.00319198f $X=1.965 $Y=3.33 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_317_n N_A_293_367#_c_360_n 0.0120807f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_312_n N_A_293_367#_c_360_n 0.0252535f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_319_n N_A_293_367#_c_360_n 0.0247015f $X=2.13 $Y=3.02 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_316_n N_A_293_367#_c_364_n 0.0189076f $X=1.965 $Y=3.33 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_312_n N_A_293_367#_c_364_n 0.012381f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_228 N_VPWR_c_319_n N_A_293_367#_c_364_n 0.0111743f $X=2.13 $Y=3.02 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_317_n N_A_293_367#_c_361_n 0.0102426f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_312_n N_A_293_367#_c_361_n 0.0113007f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_319_n N_A_293_367#_c_361_n 2.89412e-19 $X=2.13 $Y=3.02 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_312_n N_X_M1005_s 0.00314825f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_233 N_A_293_367#_c_360_n N_X_M1005_s 0.00714213f $X=2.935 $Y=2.66 $X2=0 $Y2=0
