* NGSPICE file created from sky130_fd_sc_lp__ebufn_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__ebufn_2 A TE_B VGND VNB VPB VPWR Z
M1000 a_39_367# TE_B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.071e+12p pd=9.26e+06u as=7.272e+11p ps=6.13e+06u
M1001 Z a_96_21# a_27_47# VNB nshort w=840000u l=150000u
+  ad=2.436e+11p pd=2.26e+06u as=8.232e+11p ps=7e+06u
M1002 Z a_96_21# a_39_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1003 VPWR TE_B a_39_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_47# a_284_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.06e+06u
M1005 a_96_21# A VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1006 VPWR TE_B a_284_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.56e+11p ps=2.08e+06u
M1007 VGND a_284_21# a_27_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND TE_B a_284_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1009 a_27_47# a_96_21# Z VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_39_367# a_96_21# Z VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_96_21# A VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
.ends

