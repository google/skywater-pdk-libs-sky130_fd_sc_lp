* File: sky130_fd_sc_lp__and2_lp.spice
* Created: Wed Sep  2 09:30:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2_lp.pex.spice"
.subckt sky130_fd_sc_lp__and2_lp  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1002 A_177_174# N_B_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_213_468#_M1007_d N_A_M1007_g A_177_174# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_494_92# N_A_213_468#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_213_468#_M1001_g A_494_92# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_141_468# N_B_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_213_468#_M1005_d N_B_M1005_g A_141_468# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 A_299_468# N_A_M1004_g N_A_213_468#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_299_468# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.4 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1009 A_457_468# N_A_213_468#_M1009_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_213_468#_M1006_g A_457_468# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_311 A_494_92# 0 6.97414e-20 $X=2.47 $Y=0.46
*
.include "sky130_fd_sc_lp__and2_lp.pxi.spice"
*
.ends
*
*
