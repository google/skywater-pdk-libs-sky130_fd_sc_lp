* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and2b_lp A_N B VGND VNB VPB VPWR X
X0 a_108_127# a_378_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VGND B a_313_153# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A_N a_378_159# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_510_47# A_N a_378_159# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_138_153# a_108_127# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A_N a_510_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR B a_108_127# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 X a_108_127# a_138_153# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_108_127# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_313_153# a_378_159# a_108_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
