* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or2b_lp A B_N VGND VNB VPB VPWR X
M1000 X a_290_409# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=8.5e+11p ps=5.7e+06u
M1001 a_439_57# A a_290_409# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1002 VGND B_N a_117_57# VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_597_57# a_290_409# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1004 X a_290_409# a_597_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1005 a_397_409# a_30_57# a_290_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=2.85e+11p ps=2.57e+06u
M1006 a_117_57# B_N a_30_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1007 a_275_57# a_30_57# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1008 a_290_409# a_30_57# a_275_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_439_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_397_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B_N a_30_57# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
.ends
