* File: sky130_fd_sc_lp__a2bb2o_m.pex.spice
* Created: Wed Sep  2 09:24:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%A_85_345# 1 2 9 13 17 18 21 22 24 25 28 32
+ 35 36 37
c80 37 0 1.22636e-19 $X=2.21 $Y=1.38
c81 32 0 1.22636e-19 $X=2.21 $Y=0.9
r82 35 36 4.65272 $w=1.92e-07 $l=9.58123e-08 $layer=LI1_cond $X=2.13 $Y=1.6
+ $X2=2.107 $Y2=1.685
r83 35 37 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.13 $Y=1.6 $X2=2.13
+ $Y2=1.38
r84 30 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.215
+ $X2=2.21 $Y2=1.38
r85 30 32 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.21 $Y=1.215
+ $X2=2.21 $Y2=0.9
r86 26 36 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=2.107 $Y=1.77
+ $X2=2.107 $Y2=1.685
r87 26 28 26.801 $w=2.13e-07 $l=5e-07 $layer=LI1_cond $X=2.107 $Y=1.77 $X2=2.107
+ $Y2=2.27
r88 24 36 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2 $Y=1.685 $X2=2.107
+ $Y2=1.685
r89 24 25 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=2 $Y=1.685
+ $X2=0.675 $Y2=1.685
r90 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.89 $X2=0.59 $Y2=1.89
r91 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=1.77
+ $X2=0.675 $Y2=1.685
r92 19 21 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.59 $Y=1.77
+ $X2=0.59 $Y2=1.89
r93 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=2.23
+ $X2=0.59 $Y2=1.89
r94 17 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=2.23
+ $X2=0.59 $Y2=2.395
r95 16 22 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.725
+ $X2=0.59 $Y2=1.89
r96 13 18 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.61 $Y=2.885
+ $X2=0.61 $Y2=2.395
r97 9 16 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.545 $Y=0.835
+ $X2=0.545 $Y2=1.725
r98 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=2.145 $X2=2.105 $Y2=2.27
r99 1 32 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.625 $X2=2.21 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%A1_N 3 6 8 9 10 15 17
r39 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.32
+ $X2=1.065 $Y2=1.485
r40 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.32
+ $X2=1.065 $Y2=1.155
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.065
+ $Y=1.32 $X2=1.065 $Y2=1.32
r42 9 10 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.307 $X2=1.68
+ $Y2=1.307
r43 9 16 7.67832 $w=1.93e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=1.307
+ $X2=1.065 $Y2=1.307
r44 8 16 19.6224 $w=1.93e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=1.307
+ $X2=1.065 $Y2=1.307
r45 6 18 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=1.04 $Y=2.885
+ $X2=1.04 $Y2=1.485
r46 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.975 $Y=0.835
+ $X2=0.975 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%A2_N 3 7 9 11 18
r39 18 21 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=2.035
+ $X2=1.52 $Y2=2.2
r40 18 20 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=2.035
+ $X2=1.52 $Y2=1.87
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=2.035 $X2=1.55 $Y2=2.035
r42 11 19 2.87945 $w=5.38e-07 $l=1.3e-07 $layer=LI1_cond $X=1.68 $Y=2.22
+ $X2=1.55 $Y2=2.22
r43 9 19 7.75236 $w=5.38e-07 $l=3.5e-07 $layer=LI1_cond $X=1.2 $Y=2.22 $X2=1.55
+ $Y2=2.22
r44 7 20 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=1.565 $Y=0.835
+ $X2=1.565 $Y2=1.87
r45 3 21 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.4 $Y=2.885 $X2=1.4
+ $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%A_210_125# 1 2 10 11 12 16 19 20 26 27 29
r67 29 32 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.27 $Y=0.35
+ $X2=1.27 $Y2=0.595
r68 27 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=2.9
+ $X2=2.23 $Y2=2.735
r69 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=2.9 $X2=2.23 $Y2=2.9
r70 23 26 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.615 $Y=2.9
+ $X2=2.23 $Y2=2.9
r71 20 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=0.35
+ $X2=2.085 $Y2=0.515
r72 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.085
+ $Y=0.35 $X2=2.085 $Y2=0.35
r73 17 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.35
+ $X2=1.27 $Y2=0.35
r74 17 19 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.435 $Y=0.35
+ $X2=2.085 $Y2=0.35
r75 16 38 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.32 $Y=2.355
+ $X2=2.32 $Y2=2.735
r76 13 16 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.32 $Y=1.305
+ $X2=2.32 $Y2=2.355
r77 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.245 $Y=1.23
+ $X2=2.32 $Y2=1.305
r78 11 12 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.245 $Y=1.23
+ $X2=2.07 $Y2=1.23
r79 10 36 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.995 $Y=0.835
+ $X2=1.995 $Y2=0.515
r80 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.995 $Y=1.155
+ $X2=2.07 $Y2=1.23
r81 8 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.995 $Y=1.155
+ $X2=1.995 $Y2=0.835
r82 2 23 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=2.675 $X2=1.615 $Y2=2.96
r83 1 32 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.625 $X2=1.27 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%B2 3 6 9 10 11 12 13 14 15 21
c44 21 0 1.22636e-19 $X=2.77 $Y=1.32
c45 10 0 2.62727e-19 $X=2.77 $Y=1.66
r46 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=1.32 $X2=2.77 $Y2=1.32
r47 15 22 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=2.705 $Y=1.665
+ $X2=2.705 $Y2=1.32
r48 14 22 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=2.705 $Y=1.295
+ $X2=2.705 $Y2=1.32
r49 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.705 $Y=0.925
+ $X2=2.705 $Y2=1.295
r50 12 13 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.705 $Y=0.555
+ $X2=2.705 $Y2=0.925
r51 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.77 $Y=1.66
+ $X2=2.77 $Y2=1.32
r52 10 11 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.66
+ $X2=2.77 $Y2=1.825
r53 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.155
+ $X2=2.77 $Y2=1.32
r54 6 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.75 $Y=2.355
+ $X2=2.75 $Y2=1.825
r55 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.68 $Y=0.835 $X2=2.68
+ $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%B1 3 6 9 10 11 12 14 21
c28 10 0 1.4009e-19 $X=3.31 $Y=1.66
r29 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.31
+ $Y=1.32 $X2=3.31 $Y2=1.32
r30 14 22 6.42338 $w=5.38e-07 $l=2.9e-07 $layer=LI1_cond $X=3.6 $Y=1.48 $X2=3.31
+ $Y2=1.48
r31 12 22 4.20842 $w=5.38e-07 $l=1.9e-07 $layer=LI1_cond $X=3.12 $Y=1.48
+ $X2=3.31 $Y2=1.48
r32 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.31 $Y=1.66
+ $X2=3.31 $Y2=1.32
r33 10 11 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.66
+ $X2=3.31 $Y2=1.825
r34 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.155
+ $X2=3.31 $Y2=1.32
r35 6 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.25 $Y=2.355
+ $X2=3.25 $Y2=1.825
r36 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.22 $Y=0.835 $X2=3.22
+ $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%X 1 2 7 8 9 10 11 12 13 25
r19 25 41 3.08081 $w=1.78e-07 $l=5e-08 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=0.875
r20 13 46 1.54806 $w=3.33e-07 $l=4.5e-08 $layer=LI1_cond $X=0.312 $Y=2.775
+ $X2=0.312 $Y2=2.82
r21 13 43 6.57974 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=0.312 $Y=2.775
+ $X2=0.312 $Y2=2.655
r22 12 43 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.235 $Y=2.405
+ $X2=0.235 $Y2=2.655
r23 11 12 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=2.035
+ $X2=0.235 $Y2=2.405
r24 10 11 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=2.035
r25 9 10 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r26 8 41 2.99287 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=0.31 $Y=0.857
+ $X2=0.31 $Y2=0.875
r27 8 39 3.03826 $w=3.28e-07 $l=8.7e-08 $layer=LI1_cond $X=0.31 $Y=0.857
+ $X2=0.31 $Y2=0.77
r28 8 9 21.7505 $w=1.78e-07 $l=3.53e-07 $layer=LI1_cond $X=0.235 $Y=0.942
+ $X2=0.235 $Y2=1.295
r29 8 25 1.04747 $w=1.78e-07 $l=1.7e-08 $layer=LI1_cond $X=0.235 $Y=0.942
+ $X2=0.235 $Y2=0.925
r30 7 39 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.31 $Y=0.555
+ $X2=0.31 $Y2=0.77
r31 2 46 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.25
+ $Y=2.675 $X2=0.375 $Y2=2.82
r32 1 39 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.625 $X2=0.31 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%VPWR 1 2 11 15 18 19 20 30 31 34
r40 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.825 $Y2=3.33
r48 22 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 18 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.985 $Y2=3.33
r53 17 30 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.15 $Y=3.33 $X2=3.6
+ $Y2=3.33
r54 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=2.985 $Y2=3.33
r55 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=3.245
+ $X2=2.985 $Y2=3.33
r56 13 15 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=2.985 $Y=3.245
+ $X2=2.985 $Y2=2.44
r57 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=3.33
r58 9 11 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=2.95
r59 2 15 600 $w=1.7e-07 $l=3.66367e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=2.145 $X2=2.985 $Y2=2.44
r60 1 11 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.675 $X2=0.825 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%A_479_429# 1 2 11 12
r14 13 15 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=3.465 $Y=2.175
+ $X2=3.465 $Y2=2.29
r15 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.36 $Y=2.09
+ $X2=3.465 $Y2=2.175
r16 11 12 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.36 $Y=2.09
+ $X2=2.64 $Y2=2.09
r17 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.535 $Y=2.175
+ $X2=2.64 $Y2=2.09
r18 7 9 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.535 $Y=2.175
+ $X2=2.535 $Y2=2.29
r19 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=2.145 $X2=3.465 $Y2=2.29
r20 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=2.145 $X2=2.535 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_M%VGND 1 2 3 13 14 16 18 23 27 29 38 42
r44 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 36 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r47 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r49 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r50 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 30 38 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.76
+ $Y2=0
r52 30 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r53 29 41 4.51706 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.555
+ $Y2=0
r54 29 35 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.12
+ $Y2=0
r55 27 36 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r56 27 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r57 23 25 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=1.77 $Y=0.865 $X2=1.77
+ $Y2=0.945
r58 16 41 3.24911 $w=3.3e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.435 $Y=0.085
+ $X2=3.555 $Y2=0
r59 16 18 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.435 $Y=0.085
+ $X2=3.435 $Y2=0.77
r60 15 21 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.865 $Y=0.945
+ $X2=0.76 $Y2=0.945
r61 14 25 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.675 $Y=0.945 $X2=1.77
+ $Y2=0.945
r62 14 15 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.675 $Y=0.945
+ $X2=0.865 $Y2=0.945
r63 13 21 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.86 $X2=0.76
+ $Y2=0.945
r64 12 38 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0
r65 12 13 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.86
r66 3 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.295
+ $Y=0.625 $X2=3.435 $Y2=0.77
r67 2 23 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.625 $X2=1.78 $Y2=0.865
r68 1 21 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.625 $X2=0.76 $Y2=0.865
.ends

