* File: sky130_fd_sc_lp__a21oi_1.pxi.spice
* Created: Fri Aug 28 09:51:37 2020
* 
x_PM_SKY130_FD_SC_LP__A21OI_1%A2 N_A2_M1002_g N_A2_M1005_g A2 A2 N_A2_c_41_n
+ N_A2_c_42_n PM_SKY130_FD_SC_LP__A21OI_1%A2
x_PM_SKY130_FD_SC_LP__A21OI_1%A1 N_A1_M1000_g N_A1_M1004_g A1 A1 A1 A1
+ N_A1_c_67_n A1 PM_SKY130_FD_SC_LP__A21OI_1%A1
x_PM_SKY130_FD_SC_LP__A21OI_1%B1 N_B1_c_106_n N_B1_M1003_g N_B1_M1001_g B1 B1
+ N_B1_c_109_n PM_SKY130_FD_SC_LP__A21OI_1%B1
x_PM_SKY130_FD_SC_LP__A21OI_1%A_27_367# N_A_27_367#_M1005_s N_A_27_367#_M1004_d
+ N_A_27_367#_c_135_n N_A_27_367#_c_136_n N_A_27_367#_c_139_n
+ N_A_27_367#_c_145_n N_A_27_367#_c_142_n PM_SKY130_FD_SC_LP__A21OI_1%A_27_367#
x_PM_SKY130_FD_SC_LP__A21OI_1%VPWR N_VPWR_M1005_d N_VPWR_c_164_n VPWR
+ N_VPWR_c_165_n N_VPWR_c_166_n N_VPWR_c_163_n N_VPWR_c_168_n
+ PM_SKY130_FD_SC_LP__A21OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A21OI_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_192_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__A21OI_1%Y
x_PM_SKY130_FD_SC_LP__A21OI_1%VGND N_VGND_M1002_s N_VGND_M1003_d N_VGND_c_226_n
+ N_VGND_c_227_n N_VGND_c_228_n N_VGND_c_229_n VGND N_VGND_c_230_n
+ N_VGND_c_231_n PM_SKY130_FD_SC_LP__A21OI_1%VGND
cc_1 VNB N_A2_M1005_g 0.00176105f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB A2 0.0186705f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A2_c_41_n 0.038188f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.46
cc_4 VNB N_A2_c_42_n 0.0200313f $X=-0.19 $Y=-0.245 $X2=0.377 $Y2=1.295
cc_5 VNB N_A1_M1000_g 0.0200878f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_6 VNB A1 0.00101183f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB A1 0.00389956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A1_c_67_n 0.0244135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_106_n 0.0195782f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_10 VNB N_B1_M1001_g 0.00141511f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_11 VNB B1 0.0206912f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_B1_c_109_n 0.0507303f $X=-0.19 $Y=-0.245 $X2=0.377 $Y2=1.295
cc_13 VNB N_VPWR_c_163_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_192_n 0.00313247f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB Y 0.00311435f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_VGND_c_226_n 0.0111997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_227_n 0.0371145f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_VGND_c_228_n 0.0110956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_229_n 0.0378643f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.46
cc_20 VNB N_VGND_c_230_n 0.0303048f $X=-0.19 $Y=-0.245 $X2=0.305 $Y2=1.295
cc_21 VNB N_VGND_c_231_n 0.138598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A2_M1005_g 0.0268644f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_23 VPB A2 0.00614643f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_24 VPB N_A1_M1004_g 0.0196694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB A1 0.00317393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_A1_c_67_n 0.00658433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_B1_M1001_g 0.023828f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_28 VPB B1 0.00818083f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_29 VPB N_A_27_367#_c_135_n 0.0244208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_A_27_367#_c_136_n 0.0233583f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_31 VPB N_VPWR_c_164_n 0.00561441f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_32 VPB N_VPWR_c_165_n 0.0172072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_166_n 0.0291384f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=1.295
cc_34 VPB N_VPWR_c_163_n 0.0444715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_168_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=1.665
cc_36 VPB N_Y_c_192_n 0.00136245f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_37 VPB Y 0.00868018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB Y 0.0389236f $X=-0.19 $Y=1.655 $X2=0.377 $Y2=1.46
cc_39 N_A2_c_42_n N_A1_M1000_g 0.056198f $X=0.377 $Y=1.295 $X2=0 $Y2=0
cc_40 N_A2_M1005_g N_A1_M1004_g 0.038793f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_41 A2 A1 0.0423376f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_42 N_A2_c_42_n A1 0.00609778f $X=0.377 $Y=1.295 $X2=0 $Y2=0
cc_43 N_A2_c_41_n A1 0.00609778f $X=0.37 $Y=1.46 $X2=0 $Y2=0
cc_44 A2 N_A1_c_67_n 2.74873e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_45 N_A2_c_41_n N_A1_c_67_n 0.0202647f $X=0.37 $Y=1.46 $X2=0 $Y2=0
cc_46 A2 N_A_27_367#_c_135_n 0.0190485f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A2_c_41_n N_A_27_367#_c_135_n 9.44165e-19 $X=0.37 $Y=1.46 $X2=0 $Y2=0
cc_48 N_A2_M1005_g N_A_27_367#_c_139_n 0.0263244f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_49 A2 N_A_27_367#_c_139_n 0.00480872f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A2_M1005_g N_VPWR_c_164_n 0.0040372f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_51 N_A2_M1005_g N_VPWR_c_165_n 0.00585385f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_52 N_A2_M1005_g N_VPWR_c_163_n 0.00739333f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_53 A2 N_VGND_c_227_n 0.0214592f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A2_c_41_n N_VGND_c_227_n 0.00109483f $X=0.37 $Y=1.46 $X2=0 $Y2=0
cc_55 N_A2_c_42_n N_VGND_c_227_n 0.0149878f $X=0.377 $Y=1.295 $X2=0 $Y2=0
cc_56 N_A2_c_42_n N_VGND_c_230_n 0.00400407f $X=0.377 $Y=1.295 $X2=0 $Y2=0
cc_57 N_A2_c_42_n N_VGND_c_231_n 0.00772763f $X=0.377 $Y=1.295 $X2=0 $Y2=0
cc_58 N_A1_M1000_g N_B1_c_106_n 0.0190034f $X=0.865 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_59 A1 N_B1_c_106_n 3.81247e-19 $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_60 N_A1_M1004_g N_B1_M1001_g 0.0327063f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_61 A1 N_B1_c_109_n 3.60304e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A1_c_67_n N_B1_c_109_n 0.0172057f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_63 A1 N_A_27_367#_c_139_n 0.010664f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A1_M1004_g N_A_27_367#_c_142_n 0.0242457f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_65 A1 N_A_27_367#_c_142_n 0.0194273f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A1_c_67_n N_A_27_367#_c_142_n 7.34134e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_67 N_A1_M1004_g N_VPWR_c_164_n 0.0040372f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A1_M1004_g N_VPWR_c_166_n 0.00585385f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A1_M1004_g N_VPWR_c_163_n 0.00648359f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A1_M1000_g N_Y_c_192_n 0.00137212f $X=0.865 $Y=0.765 $X2=0 $Y2=0
cc_71 N_A1_M1004_g N_Y_c_192_n 0.00441608f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_72 A1 N_Y_c_192_n 0.00713215f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_73 A1 N_Y_c_192_n 0.0308213f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A1_c_67_n N_Y_c_192_n 0.00215547f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_75 N_A1_M1000_g Y 0.00497666f $X=0.865 $Y=0.765 $X2=0 $Y2=0
cc_76 A1 Y 0.00218229f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A1_c_67_n Y 0.00346416f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_78 N_A1_M1004_g Y 0.00119064f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A1_M1000_g N_VGND_c_227_n 0.00131311f $X=0.865 $Y=0.765 $X2=0 $Y2=0
cc_80 A1 N_VGND_c_227_n 0.0440046f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_81 N_A1_M1000_g N_VGND_c_230_n 0.00454441f $X=0.865 $Y=0.765 $X2=0 $Y2=0
cc_82 A1 N_VGND_c_230_n 0.00643088f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_83 N_A1_M1000_g N_VGND_c_231_n 0.00871269f $X=0.865 $Y=0.765 $X2=0 $Y2=0
cc_84 A1 N_VGND_c_231_n 0.00674245f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 A1 A_110_69# 0.00877995f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_86 N_B1_M1001_g N_A_27_367#_c_145_n 0.00797855f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_87 N_B1_M1001_g N_A_27_367#_c_142_n 0.00267973f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_88 N_B1_M1001_g N_VPWR_c_166_n 0.0054895f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_89 N_B1_M1001_g N_VPWR_c_163_n 0.0109065f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_90 N_B1_c_106_n N_Y_c_192_n 0.00374383f $X=1.405 $Y=1.295 $X2=0 $Y2=0
cc_91 N_B1_M1001_g N_Y_c_192_n 0.0109857f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_92 B1 N_Y_c_192_n 0.0413505f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_93 N_B1_c_109_n N_Y_c_192_n 0.00761881f $X=1.65 $Y=1.46 $X2=0 $Y2=0
cc_94 N_B1_c_106_n Y 0.00931015f $X=1.405 $Y=1.295 $X2=0 $Y2=0
cc_95 N_B1_c_106_n Y 0.00622739f $X=1.405 $Y=1.295 $X2=0 $Y2=0
cc_96 N_B1_M1001_g Y 0.0148933f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_97 B1 Y 0.024812f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_98 N_B1_c_109_n Y 0.00136683f $X=1.65 $Y=1.46 $X2=0 $Y2=0
cc_99 N_B1_c_106_n N_VGND_c_229_n 0.0047964f $X=1.405 $Y=1.295 $X2=0 $Y2=0
cc_100 B1 N_VGND_c_229_n 0.0250133f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B1_c_109_n N_VGND_c_229_n 0.00175401f $X=1.65 $Y=1.46 $X2=0 $Y2=0
cc_102 N_B1_c_106_n N_VGND_c_230_n 0.00447387f $X=1.405 $Y=1.295 $X2=0 $Y2=0
cc_103 N_B1_c_106_n N_VGND_c_231_n 0.00869612f $X=1.405 $Y=1.295 $X2=0 $Y2=0
cc_104 N_A_27_367#_c_139_n N_VPWR_M1005_d 0.00376629f $X=0.75 $Y=2.2 $X2=-0.19
+ $Y2=1.655
cc_105 N_A_27_367#_c_142_n N_VPWR_M1005_d 0.00187796f $X=1.19 $Y=2.385 $X2=-0.19
+ $Y2=1.655
cc_106 N_A_27_367#_c_139_n N_VPWR_c_164_n 0.0122951f $X=0.75 $Y=2.2 $X2=0 $Y2=0
cc_107 N_A_27_367#_c_142_n N_VPWR_c_164_n 0.00806336f $X=1.19 $Y=2.385 $X2=0
+ $Y2=0
cc_108 N_A_27_367#_c_136_n N_VPWR_c_165_n 0.0190529f $X=0.26 $Y=2.48 $X2=0 $Y2=0
cc_109 N_A_27_367#_c_145_n N_VPWR_c_166_n 0.0169299f $X=1.19 $Y=2.91 $X2=0 $Y2=0
cc_110 N_A_27_367#_M1005_s N_VPWR_c_163_n 0.00220592f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_111 N_A_27_367#_M1004_d N_VPWR_c_163_n 0.0022898f $X=1.05 $Y=1.835 $X2=0
+ $Y2=0
cc_112 N_A_27_367#_c_136_n N_VPWR_c_163_n 0.0113912f $X=0.26 $Y=2.48 $X2=0 $Y2=0
cc_113 N_A_27_367#_c_139_n N_VPWR_c_163_n 0.00585868f $X=0.75 $Y=2.2 $X2=0 $Y2=0
cc_114 N_A_27_367#_c_145_n N_VPWR_c_163_n 0.0112082f $X=1.19 $Y=2.91 $X2=0 $Y2=0
cc_115 N_A_27_367#_c_142_n N_VPWR_c_163_n 0.00558016f $X=1.19 $Y=2.385 $X2=0
+ $Y2=0
cc_116 N_A_27_367#_M1004_d N_Y_c_192_n 0.00148118f $X=1.05 $Y=1.835 $X2=0 $Y2=0
cc_117 N_A_27_367#_c_142_n N_Y_c_192_n 0.00157198f $X=1.19 $Y=2.385 $X2=0 $Y2=0
cc_118 N_A_27_367#_M1004_d Y 0.00264591f $X=1.05 $Y=1.835 $X2=0 $Y2=0
cc_119 N_A_27_367#_c_142_n Y 0.0241071f $X=1.19 $Y=2.385 $X2=0 $Y2=0
cc_120 N_VPWR_c_163_n N_Y_M1001_d 0.00371702f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_121 N_VPWR_c_166_n Y 0.0213954f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_122 N_VPWR_c_163_n Y 0.0119743f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_123 Y N_VGND_c_227_n 9.80941e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_124 Y N_VGND_c_229_n 0.0280914f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_125 Y N_VGND_c_230_n 0.0184038f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_126 Y N_VGND_c_231_n 0.0138415f $X=1.115 $Y=0.47 $X2=0 $Y2=0
