* File: sky130_fd_sc_lp__nand4b_4.pxi.spice
* Created: Wed Sep  2 10:06:17 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4B_4%A_N N_A_N_M1027_g N_A_N_M1000_g A_N N_A_N_c_138_n
+ N_A_N_c_139_n PM_SKY130_FD_SC_LP__NAND4B_4%A_N
x_PM_SKY130_FD_SC_LP__NAND4B_4%A_27_51# N_A_27_51#_M1027_s N_A_27_51#_M1000_s
+ N_A_27_51#_M1007_g N_A_27_51#_M1001_g N_A_27_51#_M1008_g N_A_27_51#_M1005_g
+ N_A_27_51#_M1021_g N_A_27_51#_M1018_g N_A_27_51#_M1026_g N_A_27_51#_M1020_g
+ N_A_27_51#_c_174_n N_A_27_51#_c_175_n N_A_27_51#_c_176_n N_A_27_51#_c_185_n
+ N_A_27_51#_c_186_n N_A_27_51#_c_177_n N_A_27_51#_c_178_n N_A_27_51#_c_179_n
+ N_A_27_51#_c_206_n N_A_27_51#_c_180_n PM_SKY130_FD_SC_LP__NAND4B_4%A_27_51#
x_PM_SKY130_FD_SC_LP__NAND4B_4%B N_B_M1009_g N_B_M1002_g N_B_M1017_g N_B_M1011_g
+ N_B_M1029_g N_B_M1013_g N_B_M1033_g N_B_M1023_g B B N_B_c_293_n N_B_c_301_n
+ N_B_c_294_n PM_SKY130_FD_SC_LP__NAND4B_4%B
x_PM_SKY130_FD_SC_LP__NAND4B_4%C N_C_M1004_g N_C_M1003_g N_C_M1010_g N_C_M1014_g
+ N_C_M1019_g N_C_M1025_g N_C_M1031_g N_C_M1028_g C C N_C_c_385_p N_C_c_373_n
+ N_C_c_380_n C PM_SKY130_FD_SC_LP__NAND4B_4%C
x_PM_SKY130_FD_SC_LP__NAND4B_4%D N_D_M1006_g N_D_M1012_g N_D_M1016_g N_D_M1015_g
+ N_D_M1022_g N_D_M1024_g N_D_M1030_g N_D_M1032_g D D D N_D_c_462_n N_D_c_470_n
+ N_D_c_463_n PM_SKY130_FD_SC_LP__NAND4B_4%D
x_PM_SKY130_FD_SC_LP__NAND4B_4%VPWR N_VPWR_M1000_d N_VPWR_M1008_d N_VPWR_M1026_d
+ N_VPWR_M1017_d N_VPWR_M1033_d N_VPWR_M1010_d N_VPWR_M1031_d N_VPWR_M1016_d
+ N_VPWR_M1030_d N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n
+ N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n
+ N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n
+ N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n
+ VPWR N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n
+ N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_537_n
+ PM_SKY130_FD_SC_LP__NAND4B_4%VPWR
x_PM_SKY130_FD_SC_LP__NAND4B_4%Y N_Y_M1001_s N_Y_M1018_s N_Y_M1007_s N_Y_M1021_s
+ N_Y_M1009_s N_Y_M1029_s N_Y_M1004_s N_Y_M1019_s N_Y_M1006_s N_Y_M1022_s
+ N_Y_c_789_n N_Y_c_832_p N_Y_c_688_n N_Y_c_689_n N_Y_c_683_n N_Y_c_684_n
+ N_Y_c_794_n N_Y_c_836_p N_Y_c_685_n N_Y_c_796_n N_Y_c_686_n N_Y_c_691_n
+ N_Y_c_757_n N_Y_c_692_n N_Y_c_805_n N_Y_c_770_n N_Y_c_775_n N_Y_c_809_n
+ N_Y_c_693_n N_Y_c_687_n N_Y_c_694_n N_Y_c_695_n N_Y_c_761_n N_Y_c_696_n Y Y Y
+ Y Y N_Y_c_742_n N_Y_c_746_n N_Y_c_767_n Y N_Y_c_823_n N_Y_c_825_n
+ PM_SKY130_FD_SC_LP__NAND4B_4%Y
x_PM_SKY130_FD_SC_LP__NAND4B_4%VGND N_VGND_M1027_d N_VGND_M1012_d N_VGND_M1024_d
+ N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n VGND N_VGND_c_852_n
+ N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n N_VGND_c_857_n
+ N_VGND_c_858_n N_VGND_c_859_n PM_SKY130_FD_SC_LP__NAND4B_4%VGND
x_PM_SKY130_FD_SC_LP__NAND4B_4%A_217_51# N_A_217_51#_M1001_d N_A_217_51#_M1005_d
+ N_A_217_51#_M1020_d N_A_217_51#_M1011_s N_A_217_51#_M1023_s
+ N_A_217_51#_c_946_n N_A_217_51#_c_948_n N_A_217_51#_c_941_n
+ N_A_217_51#_c_942_n N_A_217_51#_c_943_n N_A_217_51#_c_944_n
+ PM_SKY130_FD_SC_LP__NAND4B_4%A_217_51#
x_PM_SKY130_FD_SC_LP__NAND4B_4%A_644_51# N_A_644_51#_M1002_d N_A_644_51#_M1013_d
+ N_A_644_51#_M1003_s N_A_644_51#_M1025_s N_A_644_51#_c_1005_n
+ N_A_644_51#_c_1002_n N_A_644_51#_c_1012_n N_A_644_51#_c_1013_n
+ N_A_644_51#_c_1003_n N_A_644_51#_c_1004_n N_A_644_51#_c_1023_n
+ N_A_644_51#_c_1008_n PM_SKY130_FD_SC_LP__NAND4B_4%A_644_51#
x_PM_SKY130_FD_SC_LP__NAND4B_4%A_1025_65# N_A_1025_65#_M1003_d
+ N_A_1025_65#_M1014_d N_A_1025_65#_M1028_d N_A_1025_65#_M1015_s
+ N_A_1025_65#_M1032_s N_A_1025_65#_c_1048_n N_A_1025_65#_c_1049_n
+ N_A_1025_65#_c_1050_n N_A_1025_65#_c_1051_n N_A_1025_65#_c_1052_n
+ N_A_1025_65#_c_1053_n N_A_1025_65#_c_1054_n N_A_1025_65#_c_1055_n
+ N_A_1025_65#_c_1056_n PM_SKY130_FD_SC_LP__NAND4B_4%A_1025_65#
cc_1 VNB N_A_N_M1027_g 0.0308041f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.675
cc_2 VNB N_A_N_M1000_g 0.0017668f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.465
cc_3 VNB N_A_N_c_138_n 0.00131484f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_4 VNB N_A_N_c_139_n 0.0874108f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.46
cc_5 VNB N_A_27_51#_M1001_g 0.0281965f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_6 VNB N_A_27_51#_M1005_g 0.0219833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_51#_M1018_g 0.0219833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_51#_M1020_g 0.0222121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_51#_c_174_n 0.0306079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_51#_c_175_n 0.00304001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_51#_c_176_n 0.00927731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_51#_c_177_n 0.0021887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_51#_c_178_n 0.0101068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_51#_c_179_n 2.75597e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_51#_c_180_n 0.0782018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1002_g 0.0233683f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.465
cc_17 VNB N_B_M1011_g 0.0231395f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_18 VNB N_B_M1013_g 0.0219833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_M1023_g 0.0276978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B 0.00159314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_293_n 0.0789081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_294_n 0.00123923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_M1003_g 0.0232185f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.465
cc_24 VNB N_C_M1014_g 0.0190024f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_25 VNB N_C_M1025_g 0.0199436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C_M1028_g 0.0206615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_c_373_n 0.0939361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_D_M1012_g 0.0194936f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.465
cc_29 VNB N_D_M1015_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_30 VNB N_D_M1024_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_D_M1032_g 0.0262168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB D 0.0122645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_D_c_462_n 0.0871209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_D_c_463_n 7.70431e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_537_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_683_n 0.0030484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_684_n 0.00371821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_685_n 0.0229175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_686_n 0.00868064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_687_n 0.00142194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_849_n 0.00907985f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_42 VNB N_VGND_c_850_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.46
cc_43 VNB N_VGND_c_851_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_44 VNB N_VGND_c_852_n 0.0156016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_853_n 0.147694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_854_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_855_n 0.0184219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_856_n 0.484889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_857_n 0.00528596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_858_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_859_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_217_51#_c_941_n 0.00310253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_217_51#_c_942_n 0.0133661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_217_51#_c_943_n 0.00120749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_217_51#_c_944_n 0.00120749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_644_51#_c_1002_n 0.00846753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_644_51#_c_1003_n 0.0053764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_644_51#_c_1004_n 0.00185609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1025_65#_c_1048_n 0.00753147f $X=-0.19 $Y=-0.245 $X2=0.825
+ $Y2=1.46
cc_60 VNB N_A_1025_65#_c_1049_n 0.00478913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1025_65#_c_1050_n 0.00311304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1025_65#_c_1051_n 0.00346371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1025_65#_c_1052_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1025_65#_c_1053_n 0.0120506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1025_65#_c_1054_n 0.030705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1025_65#_c_1055_n 0.00203674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1025_65#_c_1056_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VPB N_A_N_M1000_g 0.0248482f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=2.465
cc_69 VPB N_A_N_c_138_n 0.0171058f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_70 VPB N_A_27_51#_M1007_g 0.0191448f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_71 VPB N_A_27_51#_M1008_g 0.0191009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_27_51#_M1021_g 0.0191009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_27_51#_M1026_g 0.0184222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_27_51#_c_185_n 0.00688215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_27_51#_c_186_n 0.038182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_27_51#_c_179_n 0.00354111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_27_51#_c_180_n 0.0184048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_B_M1009_g 0.0184188f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.675
cc_79 VPB N_B_M1017_g 0.0179962f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_80 VPB N_B_M1029_g 0.0176757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_B_M1033_g 0.0204982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB B 0.00410879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_B_c_293_n 0.0194854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_B_c_301_n 0.00313112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_C_M1004_g 0.0213869f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.675
cc_86 VPB N_C_M1010_g 0.0179328f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_87 VPB N_C_M1019_g 0.0179221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_C_M1031_g 0.0213617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB C 0.00102559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_C_c_373_n 0.0234113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_C_c_380_n 0.00547511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_D_M1006_g 0.0210174f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.675
cc_93 VPB N_D_M1016_g 0.0182038f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_94 VPB N_D_M1022_g 0.0179162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_D_M1030_g 0.0235869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB D 0.0148584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_D_c_462_n 0.0213349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_D_c_470_n 0.00302056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_538_n 0.0069107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_539_n 0.0043704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_540_n 3.19588e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_541_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_542_n 3.12649e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_543_n 0.00174197f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_544_n 3.26939e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_545_n 0.00357855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_546_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_547_n 0.0141676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_548_n 0.0482205f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_549_n 0.0290052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_550_n 0.00439477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_551_n 0.0168265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_552_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_553_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_554_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_555_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_556_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_557_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_558_n 0.0163147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_559_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_560_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_561_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_562_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_563_n 0.0101061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_564_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_537_n 0.0644019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_Y_c_688_n 0.002757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_Y_c_689_n 0.00292381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_Y_c_686_n 0.00340976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_Y_c_691_n 0.00173326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_Y_c_692_n 0.00796461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_Y_c_693_n 0.00185325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_Y_c_694_n 0.00388183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_Y_c_695_n 0.00342814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_Y_c_696_n 0.0019754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 N_A_N_M1000_g N_A_27_51#_M1007_g 0.0191958f $X=0.825 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_N_c_139_n N_A_27_51#_M1001_g 0.00158544f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_138 N_A_N_M1027_g N_A_27_51#_c_175_n 0.0188426f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_139 N_A_N_c_138_n N_A_27_51#_c_175_n 0.00664973f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_140 N_A_N_c_139_n N_A_27_51#_c_175_n 0.00354696f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_141 N_A_N_c_138_n N_A_27_51#_c_176_n 0.0205034f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_142 N_A_N_c_139_n N_A_27_51#_c_176_n 0.00610489f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_143 N_A_N_M1000_g N_A_27_51#_c_185_n 0.00167014f $X=0.825 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_N_c_139_n N_A_27_51#_c_185_n 0.0064724f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_145 N_A_N_M1000_g N_A_27_51#_c_186_n 0.0108164f $X=0.825 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_N_M1027_g N_A_27_51#_c_177_n 0.00402317f $X=0.475 $Y=0.675 $X2=0
+ $Y2=0
cc_147 N_A_N_c_138_n N_A_27_51#_c_177_n 0.00437295f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_148 N_A_N_c_139_n N_A_27_51#_c_177_n 0.01363f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_149 N_A_N_c_139_n N_A_27_51#_c_178_n 0.00586342f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_150 N_A_N_M1000_g N_A_27_51#_c_179_n 0.009139f $X=0.825 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_N_c_138_n N_A_27_51#_c_179_n 0.0128113f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_152 N_A_N_c_139_n N_A_27_51#_c_179_n 0.00480559f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_153 N_A_N_c_138_n N_A_27_51#_c_206_n 0.0135702f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_154 N_A_N_c_139_n N_A_27_51#_c_206_n 0.0104855f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_155 N_A_N_c_139_n N_A_27_51#_c_180_n 0.0230238f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_156 N_A_N_M1000_g N_VPWR_c_538_n 0.00386211f $X=0.825 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_N_M1000_g N_VPWR_c_549_n 0.0054895f $X=0.825 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_N_M1000_g N_VPWR_c_537_n 0.0111148f $X=0.825 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_N_M1027_g N_VGND_c_849_n 0.01295f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_160 N_A_N_c_139_n N_VGND_c_849_n 0.00107744f $X=0.825 $Y=1.46 $X2=0 $Y2=0
cc_161 N_A_N_M1027_g N_VGND_c_852_n 0.00469214f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_162 N_A_N_M1027_g N_VGND_c_856_n 0.0091141f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_163 N_A_N_M1027_g N_A_217_51#_c_942_n 0.00345707f $X=0.475 $Y=0.675 $X2=0
+ $Y2=0
cc_164 N_A_27_51#_M1026_g N_B_M1009_g 0.0198158f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_27_51#_M1020_g N_B_M1002_g 0.0232711f $X=2.715 $Y=0.675 $X2=0 $Y2=0
cc_166 N_A_27_51#_c_178_n N_B_c_293_n 2.08417e-19 $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A_27_51#_c_180_n N_B_c_293_n 0.0243672f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_168 N_A_27_51#_c_178_n N_B_c_294_n 0.0119872f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A_27_51#_c_180_n N_B_c_294_n 2.84673e-19 $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A_27_51#_M1007_g N_VPWR_c_538_n 0.00267794f $X=1.265 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_27_51#_c_178_n N_VPWR_c_538_n 0.0158134f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A_27_51#_c_179_n N_VPWR_c_538_n 0.0475375f $X=0.61 $Y=1.93 $X2=0 $Y2=0
cc_173 N_A_27_51#_c_180_n N_VPWR_c_538_n 0.00160119f $X=2.715 $Y=1.51 $X2=0
+ $Y2=0
cc_174 N_A_27_51#_M1008_g N_VPWR_c_539_n 0.00178561f $X=1.695 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_27_51#_M1021_g N_VPWR_c_539_n 0.00172953f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_27_51#_M1021_g N_VPWR_c_540_n 7.37737e-19 $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_27_51#_M1026_g N_VPWR_c_540_n 0.0142861f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_27_51#_c_186_n N_VPWR_c_549_n 0.0210467f $X=0.61 $Y=2.91 $X2=0 $Y2=0
cc_179 N_A_27_51#_M1007_g N_VPWR_c_551_n 0.00585385f $X=1.265 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_27_51#_M1008_g N_VPWR_c_551_n 0.00585385f $X=1.695 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_27_51#_M1021_g N_VPWR_c_553_n 0.00585385f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_27_51#_M1026_g N_VPWR_c_553_n 0.00486043f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_27_51#_M1000_s N_VPWR_c_537_n 0.00215158f $X=0.485 $Y=1.835 $X2=0
+ $Y2=0
cc_184 N_A_27_51#_M1007_g N_VPWR_c_537_n 0.0105855f $X=1.265 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_27_51#_M1008_g N_VPWR_c_537_n 0.0107298f $X=1.695 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_27_51#_M1021_g N_VPWR_c_537_n 0.0107298f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_27_51#_M1026_g N_VPWR_c_537_n 0.00824727f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_27_51#_c_186_n N_VPWR_c_537_n 0.0125689f $X=0.61 $Y=2.91 $X2=0 $Y2=0
cc_189 N_A_27_51#_M1008_g N_Y_c_688_n 0.014097f $X=1.695 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_27_51#_M1021_g N_Y_c_688_n 0.0142104f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_27_51#_c_178_n N_Y_c_688_n 0.0447045f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_192 N_A_27_51#_c_180_n N_Y_c_688_n 0.00508846f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_193 N_A_27_51#_M1007_g N_Y_c_689_n 8.43785e-19 $X=1.265 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_27_51#_c_178_n N_Y_c_689_n 0.0208722f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A_27_51#_c_179_n N_Y_c_689_n 0.00129273f $X=0.61 $Y=1.93 $X2=0 $Y2=0
cc_196 N_A_27_51#_c_180_n N_Y_c_689_n 0.00298081f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A_27_51#_M1005_g N_Y_c_683_n 0.0123543f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_198 N_A_27_51#_M1018_g N_Y_c_683_n 0.0126682f $X=2.285 $Y=0.675 $X2=0 $Y2=0
cc_199 N_A_27_51#_c_178_n N_Y_c_683_n 0.0469373f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A_27_51#_c_180_n N_Y_c_683_n 0.002812f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A_27_51#_M1001_g N_Y_c_684_n 0.00276154f $X=1.425 $Y=0.675 $X2=0 $Y2=0
cc_202 N_A_27_51#_c_175_n N_Y_c_684_n 0.00287254f $X=0.605 $Y=1.11 $X2=0 $Y2=0
cc_203 N_A_27_51#_c_177_n N_Y_c_684_n 0.00198353f $X=0.73 $Y=1.425 $X2=0 $Y2=0
cc_204 N_A_27_51#_c_178_n N_Y_c_684_n 0.0181088f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_205 N_A_27_51#_c_180_n N_Y_c_684_n 0.00299082f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_206 N_A_27_51#_M1020_g N_Y_c_685_n 0.0126682f $X=2.715 $Y=0.675 $X2=0 $Y2=0
cc_207 N_A_27_51#_c_178_n N_Y_c_685_n 0.0141266f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_208 N_A_27_51#_c_180_n N_Y_c_685_n 2.46815e-19 $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_209 N_A_27_51#_c_178_n N_Y_c_693_n 0.0177796f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A_27_51#_c_180_n N_Y_c_693_n 0.00289569f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_211 N_A_27_51#_c_178_n N_Y_c_687_n 0.0152915f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_212 N_A_27_51#_c_180_n N_Y_c_687_n 0.00290477f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_213 N_A_27_51#_M1026_g N_Y_c_694_n 0.0131017f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A_27_51#_c_178_n N_Y_c_694_n 0.0189254f $X=2.635 $Y=1.51 $X2=0 $Y2=0
cc_215 N_A_27_51#_c_180_n N_Y_c_694_n 0.00254423f $X=2.715 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A_27_51#_c_175_n N_VGND_M1027_d 0.00262874f $X=0.605 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_27_51#_M1001_g N_VGND_c_849_n 0.00216676f $X=1.425 $Y=0.675 $X2=0
+ $Y2=0
cc_218 N_A_27_51#_c_175_n N_VGND_c_849_n 0.0240994f $X=0.605 $Y=1.11 $X2=0 $Y2=0
cc_219 N_A_27_51#_c_174_n N_VGND_c_852_n 0.0174563f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_220 N_A_27_51#_M1001_g N_VGND_c_853_n 0.00344705f $X=1.425 $Y=0.675 $X2=0
+ $Y2=0
cc_221 N_A_27_51#_M1005_g N_VGND_c_853_n 0.00344672f $X=1.855 $Y=0.675 $X2=0
+ $Y2=0
cc_222 N_A_27_51#_M1018_g N_VGND_c_853_n 0.00344672f $X=2.285 $Y=0.675 $X2=0
+ $Y2=0
cc_223 N_A_27_51#_M1020_g N_VGND_c_853_n 0.00344672f $X=2.715 $Y=0.675 $X2=0
+ $Y2=0
cc_224 N_A_27_51#_M1001_g N_VGND_c_856_n 0.00640155f $X=1.425 $Y=0.675 $X2=0
+ $Y2=0
cc_225 N_A_27_51#_M1005_g N_VGND_c_856_n 0.00520181f $X=1.855 $Y=0.675 $X2=0
+ $Y2=0
cc_226 N_A_27_51#_M1018_g N_VGND_c_856_n 0.00520181f $X=2.285 $Y=0.675 $X2=0
+ $Y2=0
cc_227 N_A_27_51#_M1020_g N_VGND_c_856_n 0.0052252f $X=2.715 $Y=0.675 $X2=0
+ $Y2=0
cc_228 N_A_27_51#_c_174_n N_VGND_c_856_n 0.00963638f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_229 N_A_27_51#_M1001_g N_A_217_51#_c_946_n 0.0121676f $X=1.425 $Y=0.675 $X2=0
+ $Y2=0
cc_230 N_A_27_51#_M1005_g N_A_217_51#_c_946_n 0.00850487f $X=1.855 $Y=0.675
+ $X2=0 $Y2=0
cc_231 N_A_27_51#_M1018_g N_A_217_51#_c_948_n 0.00850487f $X=2.285 $Y=0.675
+ $X2=0 $Y2=0
cc_232 N_A_27_51#_M1020_g N_A_217_51#_c_948_n 0.00850487f $X=2.715 $Y=0.675
+ $X2=0 $Y2=0
cc_233 N_A_27_51#_M1001_g N_A_217_51#_c_942_n 0.00368923f $X=1.425 $Y=0.675
+ $X2=0 $Y2=0
cc_234 N_A_27_51#_c_175_n N_A_217_51#_c_942_n 0.00730031f $X=0.605 $Y=1.11 $X2=0
+ $Y2=0
cc_235 N_A_27_51#_c_178_n N_A_217_51#_c_942_n 0.0153918f $X=2.635 $Y=1.51 $X2=0
+ $Y2=0
cc_236 N_A_27_51#_c_180_n N_A_217_51#_c_942_n 0.00597059f $X=2.715 $Y=1.51 $X2=0
+ $Y2=0
cc_237 N_A_27_51#_M1001_g N_A_217_51#_c_943_n 5.29781e-19 $X=1.425 $Y=0.675
+ $X2=0 $Y2=0
cc_238 N_A_27_51#_M1005_g N_A_217_51#_c_943_n 0.00732047f $X=1.855 $Y=0.675
+ $X2=0 $Y2=0
cc_239 N_A_27_51#_M1018_g N_A_217_51#_c_943_n 0.00722371f $X=2.285 $Y=0.675
+ $X2=0 $Y2=0
cc_240 N_A_27_51#_M1020_g N_A_217_51#_c_943_n 5.22442e-19 $X=2.715 $Y=0.675
+ $X2=0 $Y2=0
cc_241 N_A_27_51#_M1018_g N_A_217_51#_c_944_n 5.21592e-19 $X=2.285 $Y=0.675
+ $X2=0 $Y2=0
cc_242 N_A_27_51#_M1020_g N_A_217_51#_c_944_n 0.00722425f $X=2.715 $Y=0.675
+ $X2=0 $Y2=0
cc_243 N_B_M1033_g N_C_M1004_g 0.0107702f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B_c_293_n N_C_c_373_n 0.00998174f $X=4.535 $Y=1.51 $X2=0 $Y2=0
cc_245 N_B_M1009_g N_VPWR_c_540_n 0.0118908f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B_M1017_g N_VPWR_c_540_n 6.94733e-19 $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B_M1009_g N_VPWR_c_541_n 0.00564095f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B_M1017_g N_VPWR_c_541_n 0.00486043f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_249 N_B_M1009_g N_VPWR_c_542_n 6.80168e-19 $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_250 N_B_M1017_g N_VPWR_c_542_n 0.014522f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B_M1029_g N_VPWR_c_542_n 0.0144755f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_252 N_B_M1033_g N_VPWR_c_542_n 6.72004e-19 $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_253 N_B_M1029_g N_VPWR_c_543_n 6.85039e-19 $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_254 N_B_M1033_g N_VPWR_c_543_n 0.0168837f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B_M1029_g N_VPWR_c_557_n 0.00486043f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B_M1033_g N_VPWR_c_557_n 0.00486043f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_257 N_B_M1009_g N_VPWR_c_537_n 0.00948291f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_258 N_B_M1017_g N_VPWR_c_537_n 0.00824727f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B_M1029_g N_VPWR_c_537_n 0.00824727f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B_M1033_g N_VPWR_c_537_n 0.00824727f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_261 N_B_M1002_g N_Y_c_685_n 0.0128724f $X=3.145 $Y=0.675 $X2=0 $Y2=0
cc_262 N_B_M1011_g N_Y_c_685_n 0.011353f $X=3.655 $Y=0.675 $X2=0 $Y2=0
cc_263 N_B_M1013_g N_Y_c_685_n 0.010883f $X=4.085 $Y=0.675 $X2=0 $Y2=0
cc_264 N_B_M1023_g N_Y_c_685_n 0.012699f $X=4.515 $Y=0.675 $X2=0 $Y2=0
cc_265 N_B_c_293_n N_Y_c_685_n 0.0152941f $X=4.535 $Y=1.51 $X2=0 $Y2=0
cc_266 N_B_c_294_n N_Y_c_685_n 0.122816f $X=3.845 $Y=1.602 $X2=0 $Y2=0
cc_267 N_B_M1033_g N_Y_c_686_n 0.00266279f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_268 N_B_M1023_g N_Y_c_686_n 0.0026801f $X=4.515 $Y=0.675 $X2=0 $Y2=0
cc_269 B N_Y_c_686_n 0.0274866f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_270 N_B_c_293_n N_Y_c_686_n 0.00272364f $X=4.535 $Y=1.51 $X2=0 $Y2=0
cc_271 N_B_M1009_g N_Y_c_694_n 0.0135814f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_272 N_B_c_294_n N_Y_c_694_n 0.0482584f $X=3.845 $Y=1.602 $X2=0 $Y2=0
cc_273 N_B_M1017_g N_Y_c_695_n 0.0169443f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_274 N_B_M1029_g N_Y_c_695_n 0.00453506f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_275 N_B_c_293_n N_Y_c_695_n 0.00273522f $X=4.535 $Y=1.51 $X2=0 $Y2=0
cc_276 N_B_c_293_n Y 6.2064e-19 $X=4.535 $Y=1.51 $X2=0 $Y2=0
cc_277 N_B_c_301_n Y 0.01544f $X=4.2 $Y=1.602 $X2=0 $Y2=0
cc_278 N_B_M1033_g Y 6.75854e-19 $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_279 N_B_M1029_g N_Y_c_742_n 0.0122129f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_280 N_B_c_293_n N_Y_c_742_n 0.00249942f $X=4.535 $Y=1.51 $X2=0 $Y2=0
cc_281 N_B_c_301_n N_Y_c_742_n 0.0136881f $X=4.2 $Y=1.602 $X2=0 $Y2=0
cc_282 N_B_c_294_n N_Y_c_742_n 0.00643745f $X=3.845 $Y=1.602 $X2=0 $Y2=0
cc_283 N_B_M1033_g N_Y_c_746_n 0.0135479f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_284 B N_Y_c_746_n 0.030169f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_285 N_B_c_293_n N_Y_c_746_n 0.00123604f $X=4.535 $Y=1.51 $X2=0 $Y2=0
cc_286 N_B_M1002_g N_VGND_c_853_n 0.00344672f $X=3.145 $Y=0.675 $X2=0 $Y2=0
cc_287 N_B_M1011_g N_VGND_c_853_n 0.00344705f $X=3.655 $Y=0.675 $X2=0 $Y2=0
cc_288 N_B_M1013_g N_VGND_c_853_n 0.00344705f $X=4.085 $Y=0.675 $X2=0 $Y2=0
cc_289 N_B_M1023_g N_VGND_c_853_n 0.00344705f $X=4.515 $Y=0.675 $X2=0 $Y2=0
cc_290 N_B_M1002_g N_VGND_c_856_n 0.00540404f $X=3.145 $Y=0.675 $X2=0 $Y2=0
cc_291 N_B_M1011_g N_VGND_c_856_n 0.00538067f $X=3.655 $Y=0.675 $X2=0 $Y2=0
cc_292 N_B_M1013_g N_VGND_c_856_n 0.00520183f $X=4.085 $Y=0.675 $X2=0 $Y2=0
cc_293 N_B_M1023_g N_VGND_c_856_n 0.00640155f $X=4.515 $Y=0.675 $X2=0 $Y2=0
cc_294 N_B_M1002_g N_A_217_51#_c_941_n 0.0111138f $X=3.145 $Y=0.675 $X2=0 $Y2=0
cc_295 N_B_M1011_g N_A_217_51#_c_941_n 0.0106741f $X=3.655 $Y=0.675 $X2=0 $Y2=0
cc_296 N_B_M1013_g N_A_217_51#_c_941_n 0.0099928f $X=4.085 $Y=0.675 $X2=0 $Y2=0
cc_297 N_B_M1023_g N_A_217_51#_c_941_n 0.0101957f $X=4.515 $Y=0.675 $X2=0 $Y2=0
cc_298 N_B_M1002_g N_A_217_51#_c_944_n 0.00692766f $X=3.145 $Y=0.675 $X2=0 $Y2=0
cc_299 N_B_M1011_g N_A_217_51#_c_944_n 5.86881e-19 $X=3.655 $Y=0.675 $X2=0 $Y2=0
cc_300 N_B_M1011_g N_A_644_51#_c_1005_n 0.00977011f $X=3.655 $Y=0.675 $X2=0
+ $Y2=0
cc_301 N_B_M1013_g N_A_644_51#_c_1005_n 0.00977011f $X=4.085 $Y=0.675 $X2=0
+ $Y2=0
cc_302 N_B_M1023_g N_A_644_51#_c_1002_n 0.00995388f $X=4.515 $Y=0.675 $X2=0
+ $Y2=0
cc_303 N_B_M1023_g N_A_644_51#_c_1008_n 0.00290211f $X=4.515 $Y=0.675 $X2=0
+ $Y2=0
cc_304 N_C_M1031_g N_D_M1006_g 0.00830302f $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_305 N_C_M1028_g N_D_M1012_g 0.0150434f $X=6.855 $Y=0.745 $X2=0 $Y2=0
cc_306 N_C_c_385_p N_D_c_462_n 4.15796e-19 $X=6.755 $Y=1.51 $X2=0 $Y2=0
cc_307 N_C_c_373_n N_D_c_462_n 0.0255616f $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_308 N_C_c_385_p N_D_c_463_n 0.00924264f $X=6.755 $Y=1.51 $X2=0 $Y2=0
cc_309 N_C_c_373_n N_D_c_463_n 7.17453e-19 $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_310 N_C_M1004_g N_VPWR_c_543_n 0.0168837f $X=5.145 $Y=2.465 $X2=0 $Y2=0
cc_311 N_C_M1010_g N_VPWR_c_543_n 6.85039e-19 $X=5.575 $Y=2.465 $X2=0 $Y2=0
cc_312 N_C_M1004_g N_VPWR_c_544_n 6.72004e-19 $X=5.145 $Y=2.465 $X2=0 $Y2=0
cc_313 N_C_M1010_g N_VPWR_c_544_n 0.0144755f $X=5.575 $Y=2.465 $X2=0 $Y2=0
cc_314 N_C_M1019_g N_VPWR_c_544_n 0.0147187f $X=6.005 $Y=2.465 $X2=0 $Y2=0
cc_315 N_C_M1031_g N_VPWR_c_544_n 7.36076e-19 $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_316 N_C_M1031_g N_VPWR_c_545_n 0.00543883f $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_317 N_C_M1004_g N_VPWR_c_555_n 0.00486043f $X=5.145 $Y=2.465 $X2=0 $Y2=0
cc_318 N_C_M1010_g N_VPWR_c_555_n 0.00486043f $X=5.575 $Y=2.465 $X2=0 $Y2=0
cc_319 N_C_M1019_g N_VPWR_c_558_n 0.00486043f $X=6.005 $Y=2.465 $X2=0 $Y2=0
cc_320 N_C_M1031_g N_VPWR_c_558_n 0.00488225f $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_321 N_C_M1004_g N_VPWR_c_537_n 0.00824727f $X=5.145 $Y=2.465 $X2=0 $Y2=0
cc_322 N_C_M1010_g N_VPWR_c_537_n 0.00824727f $X=5.575 $Y=2.465 $X2=0 $Y2=0
cc_323 N_C_M1019_g N_VPWR_c_537_n 0.00824727f $X=6.005 $Y=2.465 $X2=0 $Y2=0
cc_324 N_C_M1031_g N_VPWR_c_537_n 0.00907196f $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_325 N_C_M1003_g N_Y_c_685_n 0.00345902f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_326 N_C_M1003_g N_Y_c_686_n 0.00248999f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_327 N_C_c_373_n N_Y_c_686_n 0.00923467f $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_328 N_C_c_380_n N_Y_c_686_n 0.0250457f $X=5.923 $Y=1.587 $X2=0 $Y2=0
cc_329 N_C_M1019_g N_Y_c_691_n 0.00397821f $X=6.005 $Y=2.465 $X2=0 $Y2=0
cc_330 N_C_M1031_g N_Y_c_691_n 0.0111895f $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_331 N_C_c_385_p N_Y_c_691_n 0.0193352f $X=6.755 $Y=1.51 $X2=0 $Y2=0
cc_332 N_C_c_373_n N_Y_c_691_n 0.00271404f $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_333 N_C_M1031_g N_Y_c_757_n 0.0141598f $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_334 N_C_M1031_g N_Y_c_692_n 0.00955919f $X=6.435 $Y=2.465 $X2=0 $Y2=0
cc_335 N_C_c_385_p N_Y_c_692_n 0.0350493f $X=6.755 $Y=1.51 $X2=0 $Y2=0
cc_336 N_C_c_373_n N_Y_c_692_n 0.0115467f $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_337 N_C_M1010_g N_Y_c_761_n 0.0131606f $X=5.575 $Y=2.465 $X2=0 $Y2=0
cc_338 N_C_M1019_g N_Y_c_761_n 0.0131606f $X=6.005 $Y=2.465 $X2=0 $Y2=0
cc_339 N_C_c_373_n N_Y_c_761_n 5.7877e-19 $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_340 N_C_c_380_n N_Y_c_761_n 0.0414289f $X=5.923 $Y=1.587 $X2=0 $Y2=0
cc_341 N_C_c_373_n Y 6.52992e-19 $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_342 N_C_c_380_n Y 0.0153757f $X=5.923 $Y=1.587 $X2=0 $Y2=0
cc_343 N_C_M1004_g N_Y_c_767_n 0.018881f $X=5.145 $Y=2.465 $X2=0 $Y2=0
cc_344 N_C_M1028_g N_VGND_c_850_n 5.18213e-19 $X=6.855 $Y=0.745 $X2=0 $Y2=0
cc_345 N_C_M1003_g N_VGND_c_853_n 0.00302501f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_346 N_C_M1014_g N_VGND_c_853_n 0.00302473f $X=5.915 $Y=0.745 $X2=0 $Y2=0
cc_347 N_C_M1025_g N_VGND_c_853_n 0.00302473f $X=6.345 $Y=0.745 $X2=0 $Y2=0
cc_348 N_C_M1028_g N_VGND_c_853_n 0.00302501f $X=6.855 $Y=0.745 $X2=0 $Y2=0
cc_349 N_C_M1003_g N_VGND_c_856_n 0.0048466f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_350 N_C_M1014_g N_VGND_c_856_n 0.0043467f $X=5.915 $Y=0.745 $X2=0 $Y2=0
cc_351 N_C_M1025_g N_VGND_c_856_n 0.00442121f $X=6.345 $Y=0.745 $X2=0 $Y2=0
cc_352 N_C_M1028_g N_VGND_c_856_n 0.00443098f $X=6.855 $Y=0.745 $X2=0 $Y2=0
cc_353 N_C_M1003_g N_A_217_51#_c_941_n 6.62212e-19 $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_354 N_C_M1003_g N_A_644_51#_c_1002_n 0.0109232f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_355 N_C_c_373_n N_A_644_51#_c_1002_n 0.00844955f $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_356 N_C_c_380_n N_A_644_51#_c_1002_n 0.00809776f $X=5.923 $Y=1.587 $X2=0
+ $Y2=0
cc_357 N_C_M1003_g N_A_644_51#_c_1012_n 9.04736e-19 $X=5.485 $Y=0.745 $X2=0
+ $Y2=0
cc_358 N_C_M1003_g N_A_644_51#_c_1013_n 0.00717434f $X=5.485 $Y=0.745 $X2=0
+ $Y2=0
cc_359 N_C_M1014_g N_A_644_51#_c_1003_n 0.0121896f $X=5.915 $Y=0.745 $X2=0 $Y2=0
cc_360 N_C_M1025_g N_A_644_51#_c_1003_n 0.0131595f $X=6.345 $Y=0.745 $X2=0 $Y2=0
cc_361 N_C_M1028_g N_A_644_51#_c_1003_n 0.00355738f $X=6.855 $Y=0.745 $X2=0
+ $Y2=0
cc_362 N_C_c_385_p N_A_644_51#_c_1003_n 0.026411f $X=6.755 $Y=1.51 $X2=0 $Y2=0
cc_363 N_C_c_373_n N_A_644_51#_c_1003_n 0.00746175f $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_364 N_C_c_380_n N_A_644_51#_c_1003_n 0.0486126f $X=5.923 $Y=1.587 $X2=0 $Y2=0
cc_365 N_C_M1003_g N_A_644_51#_c_1004_n 0.00585102f $X=5.485 $Y=0.745 $X2=0
+ $Y2=0
cc_366 N_C_c_373_n N_A_644_51#_c_1004_n 0.00293063f $X=6.855 $Y=1.51 $X2=0 $Y2=0
cc_367 N_C_c_380_n N_A_644_51#_c_1004_n 0.0217414f $X=5.923 $Y=1.587 $X2=0 $Y2=0
cc_368 N_C_M1028_g N_A_644_51#_c_1023_n 0.00506713f $X=6.855 $Y=0.745 $X2=0
+ $Y2=0
cc_369 N_C_M1003_g N_A_1025_65#_c_1048_n 0.012159f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_370 N_C_M1014_g N_A_1025_65#_c_1048_n 0.0110429f $X=5.915 $Y=0.745 $X2=0
+ $Y2=0
cc_371 N_C_M1025_g N_A_1025_65#_c_1049_n 0.00896715f $X=6.345 $Y=0.745 $X2=0
+ $Y2=0
cc_372 N_C_M1028_g N_A_1025_65#_c_1049_n 0.012573f $X=6.855 $Y=0.745 $X2=0 $Y2=0
cc_373 N_C_M1028_g N_A_1025_65#_c_1051_n 6.54275e-19 $X=6.855 $Y=0.745 $X2=0
+ $Y2=0
cc_374 N_C_M1003_g N_A_1025_65#_c_1055_n 7.61432e-19 $X=5.485 $Y=0.745 $X2=0
+ $Y2=0
cc_375 N_C_M1014_g N_A_1025_65#_c_1055_n 0.00688639f $X=5.915 $Y=0.745 $X2=0
+ $Y2=0
cc_376 N_C_M1025_g N_A_1025_65#_c_1055_n 0.0083414f $X=6.345 $Y=0.745 $X2=0
+ $Y2=0
cc_377 N_C_M1028_g N_A_1025_65#_c_1055_n 4.17863e-19 $X=6.855 $Y=0.745 $X2=0
+ $Y2=0
cc_378 N_D_M1006_g N_VPWR_c_545_n 0.0153615f $X=7.235 $Y=2.465 $X2=0 $Y2=0
cc_379 N_D_M1016_g N_VPWR_c_545_n 7.34156e-19 $X=7.665 $Y=2.465 $X2=0 $Y2=0
cc_380 N_D_M1006_g N_VPWR_c_546_n 6.90148e-19 $X=7.235 $Y=2.465 $X2=0 $Y2=0
cc_381 N_D_M1016_g N_VPWR_c_546_n 0.0151034f $X=7.665 $Y=2.465 $X2=0 $Y2=0
cc_382 N_D_M1022_g N_VPWR_c_546_n 0.0149184f $X=8.095 $Y=2.465 $X2=0 $Y2=0
cc_383 N_D_M1030_g N_VPWR_c_546_n 6.77662e-19 $X=8.525 $Y=2.465 $X2=0 $Y2=0
cc_384 N_D_M1022_g N_VPWR_c_548_n 7.26038e-19 $X=8.095 $Y=2.465 $X2=0 $Y2=0
cc_385 N_D_M1030_g N_VPWR_c_548_n 0.0204592f $X=8.525 $Y=2.465 $X2=0 $Y2=0
cc_386 D N_VPWR_c_548_n 0.0257064f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_387 N_D_c_462_n N_VPWR_c_548_n 0.00180524f $X=8.575 $Y=1.51 $X2=0 $Y2=0
cc_388 N_D_M1006_g N_VPWR_c_559_n 0.00486043f $X=7.235 $Y=2.465 $X2=0 $Y2=0
cc_389 N_D_M1016_g N_VPWR_c_559_n 0.00486043f $X=7.665 $Y=2.465 $X2=0 $Y2=0
cc_390 N_D_M1022_g N_VPWR_c_560_n 0.00486043f $X=8.095 $Y=2.465 $X2=0 $Y2=0
cc_391 N_D_M1030_g N_VPWR_c_560_n 0.00486043f $X=8.525 $Y=2.465 $X2=0 $Y2=0
cc_392 N_D_M1006_g N_VPWR_c_537_n 0.00824727f $X=7.235 $Y=2.465 $X2=0 $Y2=0
cc_393 N_D_M1016_g N_VPWR_c_537_n 0.00824727f $X=7.665 $Y=2.465 $X2=0 $Y2=0
cc_394 N_D_M1022_g N_VPWR_c_537_n 0.00824727f $X=8.095 $Y=2.465 $X2=0 $Y2=0
cc_395 N_D_M1030_g N_VPWR_c_537_n 0.00824727f $X=8.525 $Y=2.465 $X2=0 $Y2=0
cc_396 N_D_M1006_g N_Y_c_692_n 0.0142305f $X=7.235 $Y=2.465 $X2=0 $Y2=0
cc_397 N_D_c_463_n N_Y_c_692_n 0.00999737f $X=7.785 $Y=1.587 $X2=0 $Y2=0
cc_398 N_D_M1016_g N_Y_c_770_n 0.0121665f $X=7.665 $Y=2.465 $X2=0 $Y2=0
cc_399 N_D_M1022_g N_Y_c_770_n 0.0123204f $X=8.095 $Y=2.465 $X2=0 $Y2=0
cc_400 N_D_c_462_n N_Y_c_770_n 5.71109e-19 $X=8.575 $Y=1.51 $X2=0 $Y2=0
cc_401 N_D_c_470_n N_Y_c_770_n 0.0271006f $X=8.11 $Y=1.587 $X2=0 $Y2=0
cc_402 N_D_c_463_n N_Y_c_770_n 0.00578606f $X=7.785 $Y=1.587 $X2=0 $Y2=0
cc_403 D N_Y_c_775_n 0.014749f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_404 N_D_c_462_n N_Y_c_775_n 6.48348e-19 $X=8.575 $Y=1.51 $X2=0 $Y2=0
cc_405 N_D_M1016_g N_Y_c_696_n 0.00590633f $X=7.665 $Y=2.465 $X2=0 $Y2=0
cc_406 N_D_M1022_g N_Y_c_696_n 8.88758e-19 $X=8.095 $Y=2.465 $X2=0 $Y2=0
cc_407 N_D_c_462_n N_Y_c_696_n 0.00278273f $X=8.575 $Y=1.51 $X2=0 $Y2=0
cc_408 N_D_c_463_n N_Y_c_696_n 0.0203476f $X=7.785 $Y=1.587 $X2=0 $Y2=0
cc_409 N_D_M1012_g N_VGND_c_850_n 0.0101653f $X=7.285 $Y=0.745 $X2=0 $Y2=0
cc_410 N_D_M1015_g N_VGND_c_850_n 0.0101212f $X=7.715 $Y=0.745 $X2=0 $Y2=0
cc_411 N_D_M1024_g N_VGND_c_850_n 5.09471e-19 $X=8.145 $Y=0.745 $X2=0 $Y2=0
cc_412 N_D_M1015_g N_VGND_c_851_n 5.06642e-19 $X=7.715 $Y=0.745 $X2=0 $Y2=0
cc_413 N_D_M1024_g N_VGND_c_851_n 0.0100302f $X=8.145 $Y=0.745 $X2=0 $Y2=0
cc_414 N_D_M1032_g N_VGND_c_851_n 0.0123299f $X=8.575 $Y=0.745 $X2=0 $Y2=0
cc_415 N_D_M1012_g N_VGND_c_853_n 0.00414769f $X=7.285 $Y=0.745 $X2=0 $Y2=0
cc_416 N_D_M1015_g N_VGND_c_854_n 0.00414769f $X=7.715 $Y=0.745 $X2=0 $Y2=0
cc_417 N_D_M1024_g N_VGND_c_854_n 0.00414769f $X=8.145 $Y=0.745 $X2=0 $Y2=0
cc_418 N_D_M1032_g N_VGND_c_855_n 0.00414769f $X=8.575 $Y=0.745 $X2=0 $Y2=0
cc_419 N_D_M1012_g N_VGND_c_856_n 0.0078848f $X=7.285 $Y=0.745 $X2=0 $Y2=0
cc_420 N_D_M1015_g N_VGND_c_856_n 0.00787505f $X=7.715 $Y=0.745 $X2=0 $Y2=0
cc_421 N_D_M1024_g N_VGND_c_856_n 0.00787505f $X=8.145 $Y=0.745 $X2=0 $Y2=0
cc_422 N_D_M1032_g N_VGND_c_856_n 0.00825675f $X=8.575 $Y=0.745 $X2=0 $Y2=0
cc_423 N_D_M1012_g N_A_1025_65#_c_1049_n 5.73473e-19 $X=7.285 $Y=0.745 $X2=0
+ $Y2=0
cc_424 N_D_M1012_g N_A_1025_65#_c_1050_n 0.0129943f $X=7.285 $Y=0.745 $X2=0
+ $Y2=0
cc_425 N_D_M1015_g N_A_1025_65#_c_1050_n 0.013227f $X=7.715 $Y=0.745 $X2=0 $Y2=0
cc_426 N_D_c_462_n N_A_1025_65#_c_1050_n 0.00383837f $X=8.575 $Y=1.51 $X2=0
+ $Y2=0
cc_427 N_D_c_463_n N_A_1025_65#_c_1050_n 0.0417955f $X=7.785 $Y=1.587 $X2=0
+ $Y2=0
cc_428 N_D_M1015_g N_A_1025_65#_c_1052_n 8.28776e-19 $X=7.715 $Y=0.745 $X2=0
+ $Y2=0
cc_429 N_D_M1024_g N_A_1025_65#_c_1052_n 8.28776e-19 $X=8.145 $Y=0.745 $X2=0
+ $Y2=0
cc_430 N_D_M1024_g N_A_1025_65#_c_1053_n 0.0132834f $X=8.145 $Y=0.745 $X2=0
+ $Y2=0
cc_431 N_D_M1032_g N_A_1025_65#_c_1053_n 0.0139276f $X=8.575 $Y=0.745 $X2=0
+ $Y2=0
cc_432 D N_A_1025_65#_c_1053_n 0.0212076f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_433 N_D_c_462_n N_A_1025_65#_c_1053_n 0.00899916f $X=8.575 $Y=1.51 $X2=0
+ $Y2=0
cc_434 N_D_c_470_n N_A_1025_65#_c_1053_n 0.0469381f $X=8.11 $Y=1.587 $X2=0 $Y2=0
cc_435 N_D_M1032_g N_A_1025_65#_c_1054_n 0.00354556f $X=8.575 $Y=0.745 $X2=0
+ $Y2=0
cc_436 N_D_c_462_n N_A_1025_65#_c_1056_n 0.00276801f $X=8.575 $Y=1.51 $X2=0
+ $Y2=0
cc_437 N_D_c_470_n N_A_1025_65#_c_1056_n 0.0153331f $X=8.11 $Y=1.587 $X2=0 $Y2=0
cc_438 N_VPWR_c_537_n N_Y_M1007_s 0.00258346f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_c_537_n N_Y_M1021_s 0.00397496f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_440 N_VPWR_c_537_n N_Y_M1009_s 0.00467071f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_441 N_VPWR_c_537_n N_Y_M1029_s 0.00536646f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_442 N_VPWR_c_537_n N_Y_M1004_s 0.00536646f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_443 N_VPWR_c_537_n N_Y_M1019_s 0.00380103f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_444 N_VPWR_c_537_n N_Y_M1006_s 0.00571434f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_445 N_VPWR_c_537_n N_Y_M1022_s 0.00536646f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_446 N_VPWR_c_551_n N_Y_c_789_n 0.015291f $X=1.785 $Y=3.33 $X2=0 $Y2=0
cc_447 N_VPWR_c_537_n N_Y_c_789_n 0.0104192f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_448 N_VPWR_M1008_d N_Y_c_688_n 0.00267852f $X=1.77 $Y=1.835 $X2=0 $Y2=0
cc_449 N_VPWR_c_539_n N_Y_c_688_n 0.0191765f $X=1.95 $Y=2.21 $X2=0 $Y2=0
cc_450 N_VPWR_c_538_n N_Y_c_689_n 0.0016373f $X=1.05 $Y=1.98 $X2=0 $Y2=0
cc_451 N_VPWR_c_553_n N_Y_c_794_n 0.0138717f $X=2.685 $Y=3.33 $X2=0 $Y2=0
cc_452 N_VPWR_c_537_n N_Y_c_794_n 0.00886411f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_453 N_VPWR_c_541_n N_Y_c_796_n 0.0131621f $X=3.565 $Y=3.33 $X2=0 $Y2=0
cc_454 N_VPWR_c_537_n N_Y_c_796_n 0.00808656f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_455 N_VPWR_M1033_d N_Y_c_686_n 0.00125729f $X=4.45 $Y=1.835 $X2=0 $Y2=0
cc_456 N_VPWR_c_545_n N_Y_c_691_n 0.00129069f $X=6.68 $Y=2.27 $X2=0 $Y2=0
cc_457 N_VPWR_c_545_n N_Y_c_757_n 0.0770387f $X=6.68 $Y=2.27 $X2=0 $Y2=0
cc_458 N_VPWR_c_558_n N_Y_c_757_n 0.0184149f $X=6.595 $Y=3.33 $X2=0 $Y2=0
cc_459 N_VPWR_c_537_n N_Y_c_757_n 0.0112195f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_460 N_VPWR_M1031_d N_Y_c_692_n 0.00808513f $X=6.51 $Y=1.835 $X2=0 $Y2=0
cc_461 N_VPWR_c_545_n N_Y_c_692_n 0.0430348f $X=6.68 $Y=2.27 $X2=0 $Y2=0
cc_462 N_VPWR_c_559_n N_Y_c_805_n 0.0120977f $X=7.715 $Y=3.33 $X2=0 $Y2=0
cc_463 N_VPWR_c_537_n N_Y_c_805_n 0.00691495f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_464 N_VPWR_M1016_d N_Y_c_770_n 0.00336779f $X=7.74 $Y=1.835 $X2=0 $Y2=0
cc_465 N_VPWR_c_546_n N_Y_c_770_n 0.0170777f $X=7.88 $Y=2.355 $X2=0 $Y2=0
cc_466 N_VPWR_c_560_n N_Y_c_809_n 0.0124525f $X=8.575 $Y=3.33 $X2=0 $Y2=0
cc_467 N_VPWR_c_537_n N_Y_c_809_n 0.00730901f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_M1026_d N_Y_c_694_n 0.00197722f $X=2.71 $Y=1.835 $X2=0 $Y2=0
cc_469 N_VPWR_c_540_n N_Y_c_694_n 0.0171813f $X=2.85 $Y=2.2 $X2=0 $Y2=0
cc_470 N_VPWR_M1017_d N_Y_c_695_n 0.00185637f $X=3.59 $Y=1.835 $X2=0 $Y2=0
cc_471 N_VPWR_c_542_n N_Y_c_695_n 0.0172287f $X=3.73 $Y=2.375 $X2=0 $Y2=0
cc_472 N_VPWR_M1010_d N_Y_c_761_n 0.00334509f $X=5.65 $Y=1.835 $X2=0 $Y2=0
cc_473 N_VPWR_c_544_n N_Y_c_761_n 0.0172684f $X=5.79 $Y=2.375 $X2=0 $Y2=0
cc_474 N_VPWR_M1033_d Y 0.00208419f $X=4.45 $Y=1.835 $X2=0 $Y2=0
cc_475 N_VPWR_c_543_n Y 0.0119464f $X=4.93 $Y=2.375 $X2=0 $Y2=0
cc_476 N_VPWR_M1017_d N_Y_c_742_n 0.00330294f $X=3.59 $Y=1.835 $X2=0 $Y2=0
cc_477 N_VPWR_M1033_d N_Y_c_746_n 0.0147803f $X=4.45 $Y=1.835 $X2=0 $Y2=0
cc_478 N_VPWR_c_543_n N_Y_c_746_n 0.0320963f $X=4.93 $Y=2.375 $X2=0 $Y2=0
cc_479 N_VPWR_c_543_n N_Y_c_767_n 0.00180677f $X=4.93 $Y=2.375 $X2=0 $Y2=0
cc_480 N_VPWR_c_557_n N_Y_c_823_n 0.0124525f $X=4.425 $Y=3.33 $X2=0 $Y2=0
cc_481 N_VPWR_c_537_n N_Y_c_823_n 0.00730901f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_482 N_VPWR_c_555_n N_Y_c_825_n 0.0124525f $X=5.625 $Y=3.33 $X2=0 $Y2=0
cc_483 N_VPWR_c_537_n N_Y_c_825_n 0.00730901f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_484 N_Y_c_683_n N_A_217_51#_M1005_d 0.00176773f $X=2.405 $Y=1.165 $X2=0 $Y2=0
cc_485 N_Y_c_685_n N_A_217_51#_M1020_d 0.00176773f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_486 N_Y_c_685_n N_A_217_51#_M1011_s 0.00177204f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_487 N_Y_c_685_n N_A_217_51#_M1023_s 0.00230978f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_488 N_Y_M1001_s N_A_217_51#_c_946_n 0.00332344f $X=1.5 $Y=0.255 $X2=0 $Y2=0
cc_489 N_Y_c_832_p N_A_217_51#_c_946_n 0.0126057f $X=1.64 $Y=0.76 $X2=0 $Y2=0
cc_490 N_Y_c_683_n N_A_217_51#_c_946_n 0.00277205f $X=2.405 $Y=1.165 $X2=0 $Y2=0
cc_491 N_Y_M1018_s N_A_217_51#_c_948_n 0.00332344f $X=2.36 $Y=0.255 $X2=0 $Y2=0
cc_492 N_Y_c_683_n N_A_217_51#_c_948_n 0.00277205f $X=2.405 $Y=1.165 $X2=0 $Y2=0
cc_493 N_Y_c_836_p N_A_217_51#_c_948_n 0.0126057f $X=2.5 $Y=0.76 $X2=0 $Y2=0
cc_494 N_Y_c_685_n N_A_217_51#_c_948_n 0.00277205f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_495 N_Y_c_685_n N_A_217_51#_c_941_n 0.00328698f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_496 N_Y_c_684_n N_A_217_51#_c_942_n 0.00166618f $X=1.735 $Y=1.165 $X2=0 $Y2=0
cc_497 N_Y_c_683_n N_A_217_51#_c_943_n 0.0170813f $X=2.405 $Y=1.165 $X2=0 $Y2=0
cc_498 N_Y_c_685_n N_A_217_51#_c_944_n 0.0170813f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_499 N_Y_c_685_n N_A_644_51#_M1002_d 0.00262603f $X=4.88 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_500 N_Y_c_685_n N_A_644_51#_M1013_d 0.00177204f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_501 N_Y_c_685_n N_A_644_51#_c_1005_n 0.0910297f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_502 N_Y_c_685_n N_A_644_51#_c_1002_n 0.0144144f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_503 N_Y_c_685_n N_A_644_51#_c_1004_n 0.0073386f $X=4.88 $Y=1.165 $X2=0 $Y2=0
cc_504 N_Y_c_692_n N_A_1025_65#_c_1050_n 0.00137146f $X=7.355 $Y=1.85 $X2=0
+ $Y2=0
cc_505 N_Y_c_692_n N_A_1025_65#_c_1051_n 0.00735974f $X=7.355 $Y=1.85 $X2=0
+ $Y2=0
cc_506 N_VGND_c_853_n N_A_217_51#_c_946_n 0.0317578f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_856_n N_A_217_51#_c_946_n 0.0199763f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_853_n N_A_217_51#_c_948_n 0.0298674f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_856_n N_A_217_51#_c_948_n 0.0187823f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_c_853_n N_A_217_51#_c_941_n 0.104273f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_856_n N_A_217_51#_c_941_n 0.0656567f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_849_n N_A_217_51#_c_942_n 0.0466946f $X=0.69 $Y=0.4 $X2=0 $Y2=0
cc_513 N_VGND_c_853_n N_A_217_51#_c_942_n 0.0191601f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_856_n N_A_217_51#_c_942_n 0.0114689f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_c_853_n N_A_217_51#_c_943_n 0.0190111f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_856_n N_A_217_51#_c_943_n 0.012566f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_853_n N_A_217_51#_c_944_n 0.0190111f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_856_n N_A_217_51#_c_944_n 0.012566f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_853_n N_A_644_51#_c_1002_n 0.00320672f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_856_n N_A_644_51#_c_1002_n 0.00713532f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_853_n N_A_1025_65#_c_1048_n 0.0567626f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_856_n N_A_1025_65#_c_1048_n 0.031484f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_850_n N_A_1025_65#_c_1049_n 0.0100029f $X=7.5 $Y=0.45 $X2=0
+ $Y2=0
cc_524 N_VGND_c_853_n N_A_1025_65#_c_1049_n 0.0567354f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_856_n N_A_1025_65#_c_1049_n 0.0317249f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_M1012_d N_A_1025_65#_c_1050_n 0.00176461f $X=7.36 $Y=0.325 $X2=0
+ $Y2=0
cc_527 N_VGND_c_850_n N_A_1025_65#_c_1050_n 0.0170777f $X=7.5 $Y=0.45 $X2=0
+ $Y2=0
cc_528 N_VGND_c_850_n N_A_1025_65#_c_1052_n 0.0232405f $X=7.5 $Y=0.45 $X2=0
+ $Y2=0
cc_529 N_VGND_c_851_n N_A_1025_65#_c_1052_n 0.0228652f $X=8.36 $Y=0.45 $X2=0
+ $Y2=0
cc_530 N_VGND_c_854_n N_A_1025_65#_c_1052_n 0.0102275f $X=8.195 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_856_n N_A_1025_65#_c_1052_n 0.00712543f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_M1024_d N_A_1025_65#_c_1053_n 0.00180746f $X=8.22 $Y=0.325 $X2=0
+ $Y2=0
cc_533 N_VGND_c_851_n N_A_1025_65#_c_1053_n 0.0163515f $X=8.36 $Y=0.45 $X2=0
+ $Y2=0
cc_534 N_VGND_c_851_n N_A_1025_65#_c_1054_n 0.0229007f $X=8.36 $Y=0.45 $X2=0
+ $Y2=0
cc_535 N_VGND_c_855_n N_A_1025_65#_c_1054_n 0.0140356f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_856_n N_A_1025_65#_c_1054_n 0.00977851f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_853_n N_A_1025_65#_c_1055_n 0.0234016f $X=7.335 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_856_n N_A_1025_65#_c_1055_n 0.0125857f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_539 N_A_217_51#_c_941_n N_A_644_51#_M1002_d 0.00499647f $X=4.73 $Y=0.4
+ $X2=-0.19 $Y2=-0.245
cc_540 N_A_217_51#_c_941_n N_A_644_51#_M1013_d 0.0033716f $X=4.73 $Y=0.4 $X2=0
+ $Y2=0
cc_541 N_A_217_51#_M1011_s N_A_644_51#_c_1005_n 0.00337308f $X=3.73 $Y=0.255
+ $X2=0 $Y2=0
cc_542 N_A_217_51#_c_941_n N_A_644_51#_c_1005_n 0.0642882f $X=4.73 $Y=0.4 $X2=0
+ $Y2=0
cc_543 N_A_217_51#_M1023_s N_A_644_51#_c_1002_n 0.00534915f $X=4.59 $Y=0.255
+ $X2=0 $Y2=0
cc_544 N_A_217_51#_c_941_n N_A_644_51#_c_1002_n 0.0220541f $X=4.73 $Y=0.4 $X2=0
+ $Y2=0
cc_545 N_A_217_51#_c_941_n N_A_1025_65#_c_1048_n 0.0208109f $X=4.73 $Y=0.4 $X2=0
+ $Y2=0
cc_546 N_A_644_51#_c_1002_n N_A_1025_65#_M1003_d 0.00681515f $X=5.53 $Y=0.815
+ $X2=-0.19 $Y2=-0.245
cc_547 N_A_644_51#_c_1003_n N_A_1025_65#_M1014_d 0.00176773f $X=6.475 $Y=1.165
+ $X2=0 $Y2=0
cc_548 N_A_644_51#_M1003_s N_A_1025_65#_c_1048_n 0.00179574f $X=5.56 $Y=0.325
+ $X2=0 $Y2=0
cc_549 N_A_644_51#_c_1002_n N_A_1025_65#_c_1048_n 0.0264133f $X=5.53 $Y=0.815
+ $X2=0 $Y2=0
cc_550 N_A_644_51#_c_1012_n N_A_1025_65#_c_1048_n 0.0154348f $X=5.662 $Y=0.905
+ $X2=0 $Y2=0
cc_551 N_A_644_51#_c_1003_n N_A_1025_65#_c_1048_n 0.00353778f $X=6.475 $Y=1.165
+ $X2=0 $Y2=0
cc_552 N_A_644_51#_M1025_s N_A_1025_65#_c_1049_n 0.00261964f $X=6.42 $Y=0.325
+ $X2=0 $Y2=0
cc_553 N_A_644_51#_c_1003_n N_A_1025_65#_c_1049_n 0.00282518f $X=6.475 $Y=1.165
+ $X2=0 $Y2=0
cc_554 N_A_644_51#_c_1023_n N_A_1025_65#_c_1049_n 0.0204539f $X=6.64 $Y=0.69
+ $X2=0 $Y2=0
cc_555 N_A_644_51#_c_1003_n N_A_1025_65#_c_1051_n 0.0108938f $X=6.475 $Y=1.165
+ $X2=0 $Y2=0
cc_556 N_A_644_51#_c_1003_n N_A_1025_65#_c_1055_n 0.0170813f $X=6.475 $Y=1.165
+ $X2=0 $Y2=0
