* File: sky130_fd_sc_lp__o2bb2ai_4.spice
* Created: Fri Aug 28 11:12:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2ai_4.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2ai_4  VNB VPB B1 B2 A1_N A2_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2_N	A2_N
* A1_N	A1_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1017 N_A_35_65#_M1017_d N_B1_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005.2 A=0.126 P=1.98 MULT=1
MM1019 N_A_35_65#_M1019_d N_B1_M1019_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.8 A=0.126 P=1.98 MULT=1
MM1034 N_A_35_65#_M1019_d N_B1_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1010 N_A_35_65#_M1010_d N_B2_M1010_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1015 N_A_35_65#_M1010_d N_B2_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1029 N_A_35_65#_M1029_d N_B2_M1029_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1030 N_A_35_65#_M1029_d N_B2_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8 SB=75002.7
+ A=0.126 P=1.98 MULT=1
MM1039 N_A_35_65#_M1039_d N_B1_M1039_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1428 AS=0.1512 PD=1.18 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75003.3
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1011 N_A_35_65#_M1039_d N_A_804_39#_M1011_g N_Y_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1428 AS=0.126 PD=1.18 PS=1.14 NRD=8.568 NRS=2.856 M=1 R=5.6
+ SA=75003.8 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1023 N_A_35_65#_M1023_d N_A_804_39#_M1023_g N_Y_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1512 AS=0.126 PD=1.2 PS=1.14 NRD=11.424 NRS=0 M=1 R=5.6 SA=75004.2
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1027 N_A_35_65#_M1023_d N_A_804_39#_M1027_g N_Y_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75004.7
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1031 N_A_35_65#_M1031_d N_A_804_39#_M1031_g N_Y_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1512 PD=2.21 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75005.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_1235_65#_M1003_d N_A1_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1004 N_A_1235_65#_M1004_d N_A1_N_M1004_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1024 N_A_1235_65#_M1004_d N_A1_N_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1035 N_A_1235_65#_M1035_d N_A1_N_M1035_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1001 N_A_1235_65#_M1035_d N_A2_N_M1001_g N_A_804_39#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1016 N_A_1235_65#_M1016_d N_A2_N_M1016_g N_A_804_39#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1018 N_A_1235_65#_M1016_d N_A2_N_M1018_g N_A_804_39#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1020 N_A_1235_65#_M1020_d N_A2_N_M1020_g N_A_804_39#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2898 AS=0.1176 PD=2.37 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75003.2 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g N_A_132_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75009.1 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_B1_M1012_g N_A_132_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75008.7 A=0.189 P=2.82 MULT=1
MM1036 N_VPWR_M1012_d N_B1_M1036_g N_A_132_367#_M1036_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1953 PD=1.54 PS=1.57 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.1 SB=75008.3 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g N_A_132_367#_M1036_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1953 PD=1.54 PS=1.57 NRD=0 NRS=1.5563 M=1 R=8.4 SA=75001.5
+ SB=75007.8 A=0.189 P=2.82 MULT=1
MM1021 N_Y_M1005_d N_B2_M1021_g N_A_132_367#_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75007.4 A=0.189 P=2.82 MULT=1
MM1032 N_Y_M1032_d N_B2_M1032_g N_A_132_367#_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75006.9 A=0.189 P=2.82 MULT=1
MM1037 N_Y_M1032_d N_B2_M1037_g N_A_132_367#_M1037_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75006.5 A=0.189 P=2.82 MULT=1
MM1038 N_VPWR_M1038_d N_B1_M1038_g N_A_132_367#_M1037_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75003.2 SB=75006.1 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A_804_39#_M1002_g N_VPWR_M1038_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1002_d N_A_804_39#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1013 N_Y_M1013_d N_A_804_39#_M1013_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1025 N_Y_M1013_d N_A_804_39#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.39375 PD=1.54 PS=1.885 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1025_s N_A1_N_M1000_g N_A_804_39#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.39375 AS=0.1764 PD=1.885 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A1_N_M1006_g N_A_804_39#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.2
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1006_d N_A1_N_M1022_g N_A_804_39#_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.6
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_A1_N_M1026_g N_A_804_39#_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3906 AS=0.1764 PD=1.88 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.1
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1007 N_A_804_39#_M1007_d N_A2_N_M1007_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75007.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1014 N_A_804_39#_M1007_d N_A2_N_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1028 N_A_804_39#_M1028_d N_A2_N_M1028_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.7
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1033 N_A_804_39#_M1028_d N_A2_N_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75009.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.5079 P=24.65
*
.include "sky130_fd_sc_lp__o2bb2ai_4.pxi.spice"
*
.ends
*
*
