* File: sky130_fd_sc_lp__a41o_lp.pxi.spice
* Created: Fri Aug 28 10:03:02 2020
* 
x_PM_SKY130_FD_SC_LP__A41O_LP%A4 N_A4_M1002_g N_A4_M1010_g N_A4_c_82_n
+ N_A4_c_83_n A4 N_A4_c_84_n N_A4_c_85_n PM_SKY130_FD_SC_LP__A41O_LP%A4
x_PM_SKY130_FD_SC_LP__A41O_LP%A3 N_A3_M1005_g N_A3_M1006_g N_A3_c_116_n
+ N_A3_c_117_n N_A3_c_118_n A3 A3 A3 N_A3_c_120_n PM_SKY130_FD_SC_LP__A41O_LP%A3
x_PM_SKY130_FD_SC_LP__A41O_LP%A2 N_A2_M1007_g N_A2_M1001_g N_A2_c_163_n
+ N_A2_c_164_n N_A2_c_165_n A2 A2 A2 N_A2_c_167_n PM_SKY130_FD_SC_LP__A41O_LP%A2
x_PM_SKY130_FD_SC_LP__A41O_LP%A1 N_A1_M1000_g N_A1_c_209_n N_A1_M1012_g
+ N_A1_c_210_n A1 N_A1_c_212_n PM_SKY130_FD_SC_LP__A41O_LP%A1
x_PM_SKY130_FD_SC_LP__A41O_LP%B1 N_B1_M1008_g N_B1_M1003_g N_B1_M1004_g
+ N_B1_c_253_n N_B1_c_254_n B1 N_B1_c_255_n N_B1_c_256_n
+ PM_SKY130_FD_SC_LP__A41O_LP%B1
x_PM_SKY130_FD_SC_LP__A41O_LP%A_428_47# N_A_428_47#_M1000_d N_A_428_47#_M1003_d
+ N_A_428_47#_c_302_n N_A_428_47#_M1009_g N_A_428_47#_M1013_g
+ N_A_428_47#_c_304_n N_A_428_47#_M1011_g N_A_428_47#_c_305_n
+ N_A_428_47#_c_306_n N_A_428_47#_c_307_n N_A_428_47#_c_311_n
+ N_A_428_47#_c_312_n N_A_428_47#_c_313_n N_A_428_47#_c_308_n
+ N_A_428_47#_c_309_n PM_SKY130_FD_SC_LP__A41O_LP%A_428_47#
x_PM_SKY130_FD_SC_LP__A41O_LP%A_27_409# N_A_27_409#_M1002_s N_A_27_409#_M1006_d
+ N_A_27_409#_M1012_d N_A_27_409#_c_376_n N_A_27_409#_c_377_n
+ N_A_27_409#_c_378_n N_A_27_409#_c_379_n N_A_27_409#_c_380_n
+ N_A_27_409#_c_381_n N_A_27_409#_c_382_n PM_SKY130_FD_SC_LP__A41O_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__A41O_LP%VPWR N_VPWR_M1002_d N_VPWR_M1001_d N_VPWR_M1013_s
+ N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n
+ N_VPWR_c_434_n N_VPWR_c_435_n VPWR N_VPWR_c_436_n N_VPWR_c_428_n
+ N_VPWR_c_438_n PM_SKY130_FD_SC_LP__A41O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A41O_LP%X N_X_M1011_d N_X_M1013_d X X X X X X X
+ PM_SKY130_FD_SC_LP__A41O_LP%X
x_PM_SKY130_FD_SC_LP__A41O_LP%VGND N_VGND_M1010_s N_VGND_M1004_d N_VGND_c_500_n
+ N_VGND_c_501_n N_VGND_c_502_n VGND N_VGND_c_503_n N_VGND_c_504_n
+ N_VGND_c_505_n N_VGND_c_506_n PM_SKY130_FD_SC_LP__A41O_LP%VGND
cc_1 VNB N_A4_M1002_g 0.00325018f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_2 VNB N_A4_M1010_g 0.0257452f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_3 VNB N_A4_c_82_n 0.0317193f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=0.975
cc_4 VNB N_A4_c_83_n 0.0521067f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.263
cc_5 VNB N_A4_c_84_n 0.0351025f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_6 VNB N_A4_c_85_n 0.00713249f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_7 VNB N_A3_M1006_g 0.0145405f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_8 VNB N_A3_c_116_n 0.0159077f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.975
cc_9 VNB N_A3_c_117_n 0.0222264f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=0.825
cc_10 VNB N_A3_c_118_n 0.0131674f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=0.975
cc_11 VNB A3 0.00780765f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.263
cc_12 VNB N_A3_c_120_n 0.0155401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_M1001_g 0.0141233f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_14 VNB N_A2_c_163_n 0.0180434f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.975
cc_15 VNB N_A2_c_164_n 0.021369f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=0.825
cc_16 VNB N_A2_c_165_n 0.0126863f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=0.975
cc_17 VNB A2 0.00793839f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.263
cc_18 VNB N_A2_c_167_n 0.0155687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1000_g 0.0365899f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_20 VNB N_A1_c_209_n 0.00565132f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.825
cc_21 VNB N_A1_c_210_n 0.0252751f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=0.975
cc_22 VNB A1 0.00528672f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.263
cc_23 VNB N_A1_c_212_n 0.0168049f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.99
cc_24 VNB N_B1_M1008_g 0.03154f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_25 VNB N_B1_M1004_g 0.0287268f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=0.975
cc_26 VNB N_B1_c_253_n 0.0155013f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.99
cc_27 VNB N_B1_c_254_n 0.0100863f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_28 VNB N_B1_c_255_n 0.025357f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_29 VNB N_B1_c_256_n 0.00414282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_428_47#_c_302_n 0.0150623f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_31 VNB N_A_428_47#_M1013_g 0.0168629f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.263
cc_32 VNB N_A_428_47#_c_304_n 0.0186281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_428_47#_c_305_n 9.01586e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_428_47#_c_306_n 0.0185452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_428_47#_c_307_n 0.0112891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_428_47#_c_308_n 0.0019748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_428_47#_c_309_n 0.083643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_428_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB X 0.0170291f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_40 VNB X 0.041708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_500_n 0.0129109f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_42 VNB N_VGND_c_501_n 0.0201255f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.975
cc_43 VNB N_VGND_c_502_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_44 VNB N_VGND_c_503_n 0.0708653f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_45 VNB N_VGND_c_504_n 0.0267352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_505_n 0.230537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_506_n 0.00436611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_A4_M1002_g 0.0463652f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_49 VPB N_A3_M1006_g 0.0374403f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.445
cc_50 VPB N_A2_M1001_g 0.0381061f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.445
cc_51 VPB N_A1_c_209_n 0.00898349f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.825
cc_52 VPB N_A1_M1012_g 0.0337675f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.445
cc_53 VPB A1 7.45984e-19 $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.263
cc_54 VPB N_B1_M1003_g 0.0303112f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.445
cc_55 VPB N_B1_c_254_n 0.0266987f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_56 VPB N_B1_c_256_n 0.00187008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_428_47#_M1013_g 0.0519989f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.263
cc_58 VPB N_A_428_47#_c_311_n 0.0120153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_428_47#_c_312_n 0.0172972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_428_47#_c_313_n 0.00447011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_428_47#_c_308_n 0.00467045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_27_409#_c_376_n 0.0493899f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.263
cc_63 VPB N_A_27_409#_c_377_n 0.00528639f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_64 VPB N_A_27_409#_c_378_n 0.00962049f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_65 VPB N_A_27_409#_c_379_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_66 VPB N_A_27_409#_c_380_n 0.0168179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_27_409#_c_381_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_27_409#_c_382_n 0.00911724f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_429_n 0.0043312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_430_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_71 VPB N_VPWR_c_431_n 0.0112915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_432_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_433_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_434_n 0.0348535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_435_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_436_n 0.0189248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_428_n 0.0659721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_438_n 0.0239038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.0573842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 N_A4_c_83_n N_A3_M1006_g 0.0348419f $X=0.337 $Y=1.263 $X2=0 $Y2=0
cc_81 N_A4_c_85_n N_A3_M1006_g 2.89575e-19 $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_82 N_A4_M1010_g N_A3_c_116_n 0.0240643f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A4_c_84_n N_A3_c_117_n 0.00865959f $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_84 N_A4_c_83_n N_A3_c_118_n 0.00865959f $X=0.337 $Y=1.263 $X2=0 $Y2=0
cc_85 N_A4_M1010_g A3 0.0148571f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A4_c_82_n A3 0.00453461f $X=0.372 $Y=0.975 $X2=0 $Y2=0
cc_87 N_A4_c_83_n A3 0.0013412f $X=0.337 $Y=1.263 $X2=0 $Y2=0
cc_88 N_A4_c_84_n A3 0.0046185f $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_89 N_A4_c_85_n A3 0.0477673f $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_90 N_A4_c_82_n N_A3_c_120_n 0.0240643f $X=0.372 $Y=0.975 $X2=0 $Y2=0
cc_91 N_A4_c_85_n N_A3_c_120_n 4.16987e-19 $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_92 N_A4_M1002_g N_A_27_409#_c_376_n 0.0256336f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_93 N_A4_M1002_g N_A_27_409#_c_377_n 0.0225965f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_94 N_A4_M1002_g N_A_27_409#_c_378_n 0.00461429f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_95 N_A4_c_83_n N_A_27_409#_c_378_n 0.00237073f $X=0.337 $Y=1.263 $X2=0 $Y2=0
cc_96 N_A4_c_85_n N_A_27_409#_c_378_n 0.027138f $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_97 N_A4_M1002_g N_A_27_409#_c_382_n 0.00111611f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_98 N_A4_M1002_g N_VPWR_c_429_n 0.0237304f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_99 N_A4_M1002_g N_VPWR_c_428_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_100 N_A4_M1002_g N_VPWR_c_438_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_101 N_A4_M1010_g N_VGND_c_501_n 0.00488289f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A4_c_82_n N_VGND_c_501_n 0.00192442f $X=0.372 $Y=0.975 $X2=0 $Y2=0
cc_103 N_A4_c_85_n N_VGND_c_501_n 0.0200956f $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_104 N_A4_M1010_g N_VGND_c_503_n 0.00554661f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A4_M1010_g N_VGND_c_505_n 0.010819f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A4_c_82_n N_VGND_c_505_n 0.0014344f $X=0.372 $Y=0.975 $X2=0 $Y2=0
cc_107 N_A4_c_85_n N_VGND_c_505_n 0.00373188f $X=0.27 $Y=0.99 $X2=0 $Y2=0
cc_108 N_A3_M1006_g N_A2_M1001_g 0.03628f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_109 N_A3_c_116_n N_A2_c_163_n 0.0205025f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_110 A3 N_A2_c_163_n 0.00240735f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_111 N_A3_c_117_n N_A2_c_164_n 0.0135694f $X=1.045 $Y=1.27 $X2=0 $Y2=0
cc_112 N_A3_c_118_n N_A2_c_165_n 0.0135694f $X=1.045 $Y=1.435 $X2=0 $Y2=0
cc_113 N_A3_c_116_n A2 3.22049e-19 $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_114 A3 A2 0.0675829f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A3_c_120_n A2 0.00232522f $X=1.045 $Y=0.93 $X2=0 $Y2=0
cc_116 A3 N_A2_c_167_n 0.00232033f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A3_c_120_n N_A2_c_167_n 0.0135694f $X=1.045 $Y=0.93 $X2=0 $Y2=0
cc_118 N_A3_M1006_g N_A_27_409#_c_376_n 0.00105115f $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_119 N_A3_M1006_g N_A_27_409#_c_377_n 0.018952f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_120 N_A3_c_118_n N_A_27_409#_c_377_n 4.53543e-19 $X=1.045 $Y=1.435 $X2=0
+ $Y2=0
cc_121 A3 N_A_27_409#_c_377_n 0.0346014f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_122 N_A3_M1006_g N_A_27_409#_c_379_n 0.0166398f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_123 N_A3_M1006_g N_A_27_409#_c_382_n 0.010514f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_124 A3 N_A_27_409#_c_382_n 0.00215679f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A3_M1006_g N_VPWR_c_429_n 0.022456f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_126 N_A3_M1006_g N_VPWR_c_430_n 8.7471e-19 $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_127 N_A3_M1006_g N_VPWR_c_432_n 0.00769046f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_128 N_A3_M1006_g N_VPWR_c_428_n 0.0134474f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_129 N_A3_c_116_n N_VGND_c_503_n 0.00393362f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_130 A3 N_VGND_c_503_n 0.0159678f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_131 N_A3_c_120_n N_VGND_c_503_n 4.68218e-19 $X=1.045 $Y=0.93 $X2=0 $Y2=0
cc_132 N_A3_c_116_n N_VGND_c_505_n 0.0058113f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_133 A3 N_VGND_c_505_n 0.0198089f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_134 A3 A_128_47# 0.00175001f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_135 A3 A_206_47# 0.00375483f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_136 N_A2_c_163_n N_A1_M1000_g 0.0179759f $X=1.585 $Y=0.765 $X2=0 $Y2=0
cc_137 A2 N_A1_M1000_g 0.0109344f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_138 N_A2_c_167_n N_A1_M1000_g 0.0114898f $X=1.585 $Y=0.93 $X2=0 $Y2=0
cc_139 N_A2_M1001_g N_A1_M1012_g 0.0300833f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_140 N_A2_M1001_g N_A1_c_210_n 0.0160792f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_141 N_A2_c_165_n N_A1_c_210_n 0.0114898f $X=1.585 $Y=1.435 $X2=0 $Y2=0
cc_142 N_A2_M1001_g A1 0.0018844f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_143 N_A2_c_164_n A1 4.20122e-19 $X=1.585 $Y=1.27 $X2=0 $Y2=0
cc_144 A2 A1 0.0259387f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_145 N_A2_c_164_n N_A1_c_212_n 0.0114898f $X=1.585 $Y=1.27 $X2=0 $Y2=0
cc_146 A2 N_A_428_47#_c_305_n 0.0112455f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_147 A2 N_A_428_47#_c_307_n 0.0075595f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_148 N_A2_M1001_g N_A_27_409#_c_379_n 0.0173671f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_149 N_A2_M1001_g N_A_27_409#_c_380_n 0.0208818f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_150 A2 N_A_27_409#_c_380_n 0.00971598f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 N_A2_M1001_g N_A_27_409#_c_381_n 9.47842e-19 $X=1.605 $Y=2.545 $X2=0
+ $Y2=0
cc_152 N_A2_M1001_g N_A_27_409#_c_382_n 0.0107186f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_153 N_A2_c_165_n N_A_27_409#_c_382_n 4.43215e-19 $X=1.585 $Y=1.435 $X2=0
+ $Y2=0
cc_154 A2 N_A_27_409#_c_382_n 0.00559457f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A2_M1001_g N_VPWR_c_429_n 9.45383e-19 $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_156 N_A2_M1001_g N_VPWR_c_430_n 0.0189972f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_157 N_A2_M1001_g N_VPWR_c_432_n 0.00769046f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_158 N_A2_M1001_g N_VPWR_c_428_n 0.0134474f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_159 N_A2_c_163_n N_VGND_c_503_n 0.00394642f $X=1.585 $Y=0.765 $X2=0 $Y2=0
cc_160 A2 N_VGND_c_503_n 0.0107238f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_161 N_A2_c_167_n N_VGND_c_503_n 4.70867e-19 $X=1.585 $Y=0.93 $X2=0 $Y2=0
cc_162 N_A2_c_163_n N_VGND_c_505_n 0.00623283f $X=1.585 $Y=0.765 $X2=0 $Y2=0
cc_163 A2 N_VGND_c_505_n 0.0122628f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_164 A2 A_314_47# 0.00550164f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_165 N_A1_M1000_g N_B1_M1008_g 0.0207188f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A1_c_212_n N_B1_c_253_n 0.00798507f $X=2.155 $Y=1.24 $X2=0 $Y2=0
cc_167 N_A1_M1012_g N_B1_c_254_n 0.0217693f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_168 N_A1_c_210_n N_B1_c_254_n 0.00862587f $X=2.155 $Y=1.58 $X2=0 $Y2=0
cc_169 A1 N_B1_c_255_n 5.34947e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A1_c_212_n N_B1_c_255_n 0.00862587f $X=2.155 $Y=1.24 $X2=0 $Y2=0
cc_171 A1 N_B1_c_256_n 0.0473754f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A1_c_212_n N_B1_c_256_n 0.00482803f $X=2.155 $Y=1.24 $X2=0 $Y2=0
cc_173 N_A1_M1000_g N_A_428_47#_c_305_n 0.00812509f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_174 N_A1_M1000_g N_A_428_47#_c_307_n 0.00229105f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_175 A1 N_A_428_47#_c_307_n 0.00542506f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A1_c_212_n N_A_428_47#_c_307_n 4.91333e-19 $X=2.155 $Y=1.24 $X2=0 $Y2=0
cc_177 N_A1_M1012_g N_A_428_47#_c_311_n 2.53923e-19 $X=2.155 $Y=2.545 $X2=0
+ $Y2=0
cc_178 N_A1_M1012_g N_A_27_409#_c_379_n 2.23645e-19 $X=2.155 $Y=2.545 $X2=0
+ $Y2=0
cc_179 N_A1_c_209_n N_A_27_409#_c_380_n 5.7112e-19 $X=2.155 $Y=1.745 $X2=0 $Y2=0
cc_180 N_A1_M1012_g N_A_27_409#_c_380_n 0.0206823f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_181 A1 N_A_27_409#_c_380_n 0.0246384f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A1_M1012_g N_A_27_409#_c_381_n 0.0179471f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_183 N_A1_M1012_g N_A_27_409#_c_382_n 0.00154414f $X=2.155 $Y=2.545 $X2=0
+ $Y2=0
cc_184 A1 N_A_27_409#_c_382_n 0.00223727f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A1_M1012_g N_VPWR_c_430_n 0.0171497f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_186 N_A1_M1012_g N_VPWR_c_434_n 0.00840515f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_187 N_A1_M1012_g N_VPWR_c_428_n 0.0146909f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_188 N_A1_M1000_g N_VGND_c_503_n 0.00585385f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A1_M1000_g N_VGND_c_505_n 0.011682f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_190 N_B1_M1004_g N_A_428_47#_c_302_n 0.0152538f $X=2.995 $Y=0.445 $X2=0 $Y2=0
cc_191 N_B1_c_255_n N_A_428_47#_M1013_g 0.0044919f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_192 N_B1_c_256_n N_A_428_47#_M1013_g 2.32594e-19 $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_193 N_B1_M1008_g N_A_428_47#_c_305_n 0.00881509f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_B1_M1004_g N_A_428_47#_c_305_n 0.00166179f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_195 N_B1_M1008_g N_A_428_47#_c_306_n 0.00838196f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_B1_M1004_g N_A_428_47#_c_306_n 0.0137461f $X=2.995 $Y=0.445 $X2=0 $Y2=0
cc_197 N_B1_c_253_n N_A_428_47#_c_306_n 7.77439e-19 $X=2.815 $Y=1.225 $X2=0
+ $Y2=0
cc_198 N_B1_c_256_n N_A_428_47#_c_306_n 0.0300491f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_199 N_B1_M1008_g N_A_428_47#_c_307_n 0.00302441f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_B1_c_256_n N_A_428_47#_c_307_n 0.00511128f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_201 N_B1_M1003_g N_A_428_47#_c_311_n 0.0168f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_202 N_B1_M1003_g N_A_428_47#_c_313_n 0.00622019f $X=2.685 $Y=2.545 $X2=0
+ $Y2=0
cc_203 N_B1_c_254_n N_A_428_47#_c_313_n 0.00869635f $X=2.865 $Y=1.54 $X2=0 $Y2=0
cc_204 N_B1_c_256_n N_A_428_47#_c_313_n 0.0172898f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_205 N_B1_M1004_g N_A_428_47#_c_308_n 0.00264563f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_B1_c_254_n N_A_428_47#_c_308_n 0.00488753f $X=2.865 $Y=1.54 $X2=0 $Y2=0
cc_207 N_B1_c_255_n N_A_428_47#_c_308_n 0.00331259f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_208 N_B1_c_256_n N_A_428_47#_c_308_n 0.0312314f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_209 N_B1_M1004_g N_A_428_47#_c_309_n 0.0353386f $X=2.995 $Y=0.445 $X2=0 $Y2=0
cc_210 N_B1_c_256_n N_A_428_47#_c_309_n 0.00132582f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_211 N_B1_M1003_g N_A_27_409#_c_380_n 0.0047165f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_212 N_B1_c_256_n N_A_27_409#_c_380_n 0.00525347f $X=2.825 $Y=1.24 $X2=0 $Y2=0
cc_213 N_B1_M1003_g N_A_27_409#_c_381_n 0.0173747f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_214 N_B1_M1003_g N_VPWR_c_430_n 8.5838e-19 $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_215 N_B1_M1003_g N_VPWR_c_431_n 0.00332836f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_216 N_B1_M1003_g N_VPWR_c_434_n 0.00826654f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_217 N_B1_M1003_g N_VPWR_c_428_n 0.0158042f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_218 N_B1_M1008_g N_VGND_c_502_n 0.0020441f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_219 N_B1_M1004_g N_VGND_c_502_n 0.0101025f $X=2.995 $Y=0.445 $X2=0 $Y2=0
cc_220 N_B1_M1008_g N_VGND_c_503_n 0.00426341f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_221 N_B1_M1004_g N_VGND_c_503_n 0.00364083f $X=2.995 $Y=0.445 $X2=0 $Y2=0
cc_222 N_B1_M1008_g N_VGND_c_505_n 0.00623968f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_223 N_B1_M1004_g N_VGND_c_505_n 0.00416707f $X=2.995 $Y=0.445 $X2=0 $Y2=0
cc_224 N_A_428_47#_c_313_n N_A_27_409#_c_380_n 0.0126166f $X=3.115 $Y=2.01 $X2=0
+ $Y2=0
cc_225 N_A_428_47#_c_311_n N_A_27_409#_c_381_n 0.0638481f $X=2.95 $Y=2.19 $X2=0
+ $Y2=0
cc_226 N_A_428_47#_c_312_n N_VPWR_M1013_s 0.00287554f $X=3.325 $Y=2.01 $X2=0
+ $Y2=0
cc_227 N_A_428_47#_M1013_g N_VPWR_c_431_n 0.022264f $X=3.775 $Y=2.545 $X2=0
+ $Y2=0
cc_228 N_A_428_47#_c_311_n N_VPWR_c_431_n 0.0532606f $X=2.95 $Y=2.19 $X2=0 $Y2=0
cc_229 N_A_428_47#_c_312_n N_VPWR_c_431_n 0.0216833f $X=3.325 $Y=2.01 $X2=0
+ $Y2=0
cc_230 N_A_428_47#_c_311_n N_VPWR_c_434_n 0.0220321f $X=2.95 $Y=2.19 $X2=0 $Y2=0
cc_231 N_A_428_47#_M1013_g N_VPWR_c_436_n 0.00769046f $X=3.775 $Y=2.545 $X2=0
+ $Y2=0
cc_232 N_A_428_47#_M1013_g N_VPWR_c_428_n 0.014085f $X=3.775 $Y=2.545 $X2=0
+ $Y2=0
cc_233 N_A_428_47#_c_311_n N_VPWR_c_428_n 0.0125808f $X=2.95 $Y=2.19 $X2=0 $Y2=0
cc_234 N_A_428_47#_c_302_n X 0.00141229f $X=3.425 $Y=0.765 $X2=0 $Y2=0
cc_235 N_A_428_47#_c_304_n X 0.008729f $X=3.785 $Y=0.765 $X2=0 $Y2=0
cc_236 N_A_428_47#_c_309_n X 7.4405e-19 $X=3.49 $Y=0.93 $X2=0 $Y2=0
cc_237 N_A_428_47#_M1013_g X 0.0468136f $X=3.775 $Y=2.545 $X2=0 $Y2=0
cc_238 N_A_428_47#_c_304_n X 0.00313171f $X=3.785 $Y=0.765 $X2=0 $Y2=0
cc_239 N_A_428_47#_c_306_n X 0.0113826f $X=3.325 $Y=0.81 $X2=0 $Y2=0
cc_240 N_A_428_47#_c_312_n X 0.0110302f $X=3.325 $Y=2.01 $X2=0 $Y2=0
cc_241 N_A_428_47#_c_308_n X 0.0627755f $X=3.49 $Y=0.93 $X2=0 $Y2=0
cc_242 N_A_428_47#_c_309_n X 0.0263924f $X=3.49 $Y=0.93 $X2=0 $Y2=0
cc_243 N_A_428_47#_c_302_n N_VGND_c_502_n 0.0101015f $X=3.425 $Y=0.765 $X2=0
+ $Y2=0
cc_244 N_A_428_47#_c_304_n N_VGND_c_502_n 0.0020441f $X=3.785 $Y=0.765 $X2=0
+ $Y2=0
cc_245 N_A_428_47#_c_305_n N_VGND_c_502_n 0.00936806f $X=2.42 $Y=0.47 $X2=0
+ $Y2=0
cc_246 N_A_428_47#_c_306_n N_VGND_c_502_n 0.0199436f $X=3.325 $Y=0.81 $X2=0
+ $Y2=0
cc_247 N_A_428_47#_c_305_n N_VGND_c_503_n 0.0196636f $X=2.42 $Y=0.47 $X2=0 $Y2=0
cc_248 N_A_428_47#_c_306_n N_VGND_c_503_n 0.00652017f $X=3.325 $Y=0.81 $X2=0
+ $Y2=0
cc_249 N_A_428_47#_c_302_n N_VGND_c_504_n 0.00363971f $X=3.425 $Y=0.765 $X2=0
+ $Y2=0
cc_250 N_A_428_47#_c_304_n N_VGND_c_504_n 0.00549284f $X=3.785 $Y=0.765 $X2=0
+ $Y2=0
cc_251 N_A_428_47#_c_306_n N_VGND_c_504_n 0.00446428f $X=3.325 $Y=0.81 $X2=0
+ $Y2=0
cc_252 N_A_428_47#_M1000_d N_VGND_c_505_n 0.00743588f $X=2.14 $Y=0.235 $X2=0
+ $Y2=0
cc_253 N_A_428_47#_c_302_n N_VGND_c_505_n 0.00416497f $X=3.425 $Y=0.765 $X2=0
+ $Y2=0
cc_254 N_A_428_47#_c_304_n N_VGND_c_505_n 0.0109412f $X=3.785 $Y=0.765 $X2=0
+ $Y2=0
cc_255 N_A_428_47#_c_305_n N_VGND_c_505_n 0.0125545f $X=2.42 $Y=0.47 $X2=0 $Y2=0
cc_256 N_A_428_47#_c_306_n N_VGND_c_505_n 0.0196691f $X=3.325 $Y=0.81 $X2=0
+ $Y2=0
cc_257 N_A_27_409#_c_380_n N_VPWR_M1001_d 0.00202522f $X=2.255 $Y=2.01 $X2=0
+ $Y2=0
cc_258 N_A_27_409#_c_376_n N_VPWR_c_429_n 0.0685263f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_259 N_A_27_409#_c_377_n N_VPWR_c_429_n 0.0262011f $X=1.175 $Y=1.76 $X2=0
+ $Y2=0
cc_260 N_A_27_409#_c_382_n N_VPWR_c_429_n 0.0684934f $X=1.34 $Y=1.76 $X2=0 $Y2=0
cc_261 N_A_27_409#_c_379_n N_VPWR_c_430_n 0.0520536f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_262 N_A_27_409#_c_380_n N_VPWR_c_430_n 0.0164557f $X=2.255 $Y=2.01 $X2=0
+ $Y2=0
cc_263 N_A_27_409#_c_381_n N_VPWR_c_430_n 0.0482418f $X=2.42 $Y=2.19 $X2=0 $Y2=0
cc_264 N_A_27_409#_c_379_n N_VPWR_c_432_n 0.021949f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_265 N_A_27_409#_c_381_n N_VPWR_c_434_n 0.021949f $X=2.42 $Y=2.19 $X2=0 $Y2=0
cc_266 N_A_27_409#_c_376_n N_VPWR_c_428_n 0.0125808f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_267 N_A_27_409#_c_379_n N_VPWR_c_428_n 0.0124703f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_268 N_A_27_409#_c_381_n N_VPWR_c_428_n 0.0124703f $X=2.42 $Y=2.19 $X2=0 $Y2=0
cc_269 N_A_27_409#_c_376_n N_VPWR_c_438_n 0.0220321f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_270 N_VPWR_c_431_n X 0.0520536f $X=3.51 $Y=2.44 $X2=0 $Y2=0
cc_271 N_VPWR_c_436_n X 0.0220321f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_428_n X 0.0125808f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_273 X N_VGND_c_502_n 0.0094508f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_274 X N_VGND_c_504_n 0.0224313f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_275 N_X_M1011_d N_VGND_c_505_n 0.00232985f $X=3.86 $Y=0.235 $X2=0 $Y2=0
cc_276 X N_VGND_c_505_n 0.0141088f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_277 N_VGND_c_505_n A_128_47# 0.00219029f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_278 N_VGND_c_505_n A_206_47# 0.0106378f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_279 N_VGND_c_505_n A_314_47# 0.010459f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_280 N_VGND_c_505_n A_542_47# 0.00271994f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_281 N_VGND_c_505_n A_700_47# 0.00436087f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
