* File: sky130_fd_sc_lp__o22a_lp.spice
* Created: Wed Sep  2 10:20:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o22a_lp  VNB VPB A1 A2 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A1_M1007_g N_A_30_173#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.08085 AS=0.1197 PD=0.805 PS=1.41 NRD=4.284 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_30_173#_M1004_d N_A2_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.08085 PD=0.7 PS=0.805 NRD=0 NRS=25.704 M=1 R=2.8 SA=75000.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_232_419#_M1005_d N_B2_M1005_g N_A_30_173#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.125025 AS=0.0588 PD=1.085 PS=0.7 NRD=69.336 NRS=0 M=1 R=2.8
+ SA=75001.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_30_173#_M1003_d N_B1_M1003_g N_A_232_419#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.125025 PD=1.41 PS=1.085 NRD=0 NRS=69.336 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 A_612_47# N_A_232_419#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_232_419#_M1000_g A_612_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_134_419# N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1001 N_A_232_419#_M1001_d N_A2_M1001_g A_134_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1006 A_338_419# N_B2_M1006_g N_A_232_419#_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=18.6953 NRS=0 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g A_338_419# VPB PHIGHVT L=0.25 W=1 AD=0.41
+ AS=0.15 PD=1.82 PS=1.3 NRD=0.9653 NRS=18.6953 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1002 N_X_M1002_d N_A_232_419#_M1002_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.41 PD=2.57 PS=1.82 NRD=0 NRS=105.375 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=7.5401 P=12.69
*
.include "sky130_fd_sc_lp__o22a_lp.pxi.spice"
*
.ends
*
*
