* NGSPICE file created from sky130_fd_sc_lp__a31o_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 a_269_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.749e+11p pd=6.27e+06u as=1.2726e+12p ps=7.06e+06u
M1001 VPWR a_80_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1002 a_269_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=7.644e+11p ps=5.18e+06u
M1003 a_347_47# A2 a_269_47# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1004 VGND a_80_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1005 a_269_367# A3 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_80_21# B1 a_269_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1007 a_80_21# A1 a_347_47# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1008 VGND B1 a_80_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_269_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

