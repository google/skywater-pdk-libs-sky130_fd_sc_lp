* File: sky130_fd_sc_lp__sdfbbn_1.pex.spice
* Created: Wed Sep  2 10:33:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%SCD 2 5 9 11 12 15 16
c32 5 0 1.17915e-19 $X=0.495 $Y=2.69
r33 15 17 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.415 $Y=1.38
+ $X2=0.415 $Y2=1.215
r34 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.38 $X2=0.385 $Y2=1.38
r35 12 16 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.55
+ $X2=0.385 $Y2=1.55
r36 9 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.535 $Y=0.805
+ $X2=0.535 $Y2=1.215
r37 5 11 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.495 $Y=2.69
+ $X2=0.495 $Y2=1.885
r38 2 11 44.2525 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=0.415 $Y=1.69
+ $X2=0.415 $Y2=1.885
r39 1 15 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.415 $Y=1.41 $X2=0.415
+ $Y2=1.38
r40 1 2 39.929 $w=3.9e-07 $l=2.8e-07 $layer=POLY_cond $X=0.415 $Y=1.41 $X2=0.415
+ $Y2=1.69
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%D 3 7 10 15 16 17 22
c49 15 0 1.41106e-19 $X=1.68 $Y=0.925
r50 22 24 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.315
+ $X2=1.62 $Y2=1.15
r51 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.655 $Y=1.295
+ $X2=1.655 $Y2=1.665
r52 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.655
+ $Y=1.315 $X2=1.655 $Y2=1.315
r53 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.655 $Y=0.925
+ $X2=1.655 $Y2=1.295
r54 10 11 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.62 $Y=1.86
+ $X2=1.285 $Y2=1.86
r55 9 22 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=1.62 $Y=1.35 $X2=1.62
+ $Y2=1.315
r56 9 10 60.4817 $w=4e-07 $l=4.35e-07 $layer=POLY_cond $X=1.62 $Y=1.35 $X2=1.62
+ $Y2=1.785
r57 7 24 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.495 $Y=0.805
+ $X2=1.495 $Y2=1.15
r58 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.285 $Y=1.935
+ $X2=1.285 $Y2=1.86
r59 1 3 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.285 $Y=1.935
+ $X2=1.285 $Y2=2.69
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_328_429# 1 2 7 9 10 11 14 17 19 20 23 26
+ 29 32 35
c73 11 0 1.41106e-19 $X=1.79 $Y=2.22
r74 32 34 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.26 $Y=0.805
+ $X2=3.26 $Y2=1.035
r75 27 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.505
+ $X2=3.18 $Y2=1.34
r76 27 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.18 $Y=1.505
+ $X2=3.18 $Y2=2.2
r77 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.175
+ $X2=3.18 $Y2=1.34
r78 26 34 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.18 $Y=1.175
+ $X2=3.18 $Y2=1.035
r79 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.34 $X2=2.515 $Y2=1.34
r80 20 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=1.34
+ $X2=3.18 $Y2=1.34
r81 20 22 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=3.095 $Y=1.34
+ $X2=2.515 $Y2=1.34
r82 18 23 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.21 $Y=1.34
+ $X2=2.515 $Y2=1.34
r83 18 19 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=1.34
+ $X2=2.135 $Y2=1.34
r84 16 19 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.505
+ $X2=2.135 $Y2=1.34
r85 16 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.135 $Y=1.505
+ $X2=2.135 $Y2=2.145
r86 12 19 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.175
+ $X2=2.135 $Y2=1.34
r87 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.135 $Y=1.175
+ $X2=2.135 $Y2=0.805
r88 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.06 $Y=2.22
+ $X2=2.135 $Y2=2.145
r89 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.06 $Y=2.22
+ $X2=1.79 $Y2=2.22
r90 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.715 $Y=2.295
+ $X2=1.79 $Y2=2.22
r91 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.715 $Y=2.295
+ $X2=1.715 $Y2=2.69
r92 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.04
+ $Y=2.055 $X2=3.18 $Y2=2.2
r93 1 32 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=3.04
+ $Y=0.595 $X2=3.26 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%SCE 4 7 9 10 13 15 17 20 21
r65 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.38
+ $X2=1.015 $Y2=1.545
r66 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.38
+ $X2=1.015 $Y2=1.215
r67 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.015
+ $Y=1.38 $X2=1.015 $Y2=1.38
r68 17 21 7.41049 $w=4.58e-07 $l=2.85e-07 $layer=LI1_cond $X=1.08 $Y=1.665
+ $X2=1.08 $Y2=1.38
r69 13 15 805.043 $w=1.5e-07 $l=1.57e-06 $layer=POLY_cond $X=2.965 $Y=0.805
+ $X2=2.965 $Y2=2.375
r70 11 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.965 $Y=0.255
+ $X2=2.965 $Y2=0.805
r71 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.89 $Y=0.18
+ $X2=2.965 $Y2=0.255
r72 9 10 969.128 $w=1.5e-07 $l=1.89e-06 $layer=POLY_cond $X=2.89 $Y=0.18 $X2=1
+ $Y2=0.18
r73 7 23 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=0.925 $Y=2.69
+ $X2=0.925 $Y2=1.545
r74 4 22 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.925 $Y=0.805
+ $X2=0.925 $Y2=1.215
r75 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=1 $Y2=0.18
r76 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=0.925 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%CLK_N 3 6 7 9 12 13 16 18 21 22
r49 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.025
+ $Y=1.035 $X2=4.025 $Y2=1.035
r50 18 22 8.94433 $w=3.33e-07 $l=2.6e-07 $layer=LI1_cond $X=4.027 $Y=1.295
+ $X2=4.027 $Y2=1.035
r51 14 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.115 $Y=1.855
+ $X2=4.365 $Y2=1.855
r52 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.025 $Y=1.375
+ $X2=4.025 $Y2=1.035
r53 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.375
+ $X2=4.025 $Y2=1.54
r54 11 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=0.87
+ $X2=4.025 $Y2=1.035
r55 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.365 $Y=1.93
+ $X2=4.365 $Y2=1.855
r56 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.365 $Y=1.93
+ $X2=4.365 $Y2=2.375
r57 6 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.115 $Y=1.78
+ $X2=4.115 $Y2=1.855
r58 6 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.115 $Y=1.78
+ $X2=4.115 $Y2=1.54
r59 3 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.115 $Y=0.46
+ $X2=4.115 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_838_50# 1 2 10 14 15 16 17 18 21 26 29 30
+ 32 33 34 38 43 46 50 51 53 54 56 57 58 60 61 62 63 64 65 66 69 70 73 77 79 80
+ 84 93
c249 84 0 2.25888e-20 $X=11.365 $Y=1.51
c250 70 0 3.07529e-20 $X=12.265 $Y=1.865
c251 50 0 4.10494e-20 $X=7.21 $Y=1.215
r252 84 93 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.365 $Y=1.51
+ $X2=11.365 $Y2=1.345
r253 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.365
+ $Y=1.51 $X2=11.365 $Y2=1.51
r254 77 79 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.567 $Y=1.035
+ $X2=4.567 $Y2=0.87
r255 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.595
+ $Y=1.035 $X2=4.595 $Y2=1.035
r256 75 79 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.46 $Y=0.69
+ $X2=4.46 $Y2=0.87
r257 73 75 10.0876 $w=3.78e-07 $l=2.15e-07 $layer=LI1_cond $X=4.355 $Y=0.475
+ $X2=4.355 $Y2=0.69
r258 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.265
+ $Y=1.865 $X2=12.265 $Y2=1.865
r259 67 69 35.9702 $w=3.28e-07 $l=1.03e-06 $layer=LI1_cond $X=12.265 $Y=2.895
+ $X2=12.265 $Y2=1.865
r260 65 67 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.1 $Y=2.98
+ $X2=12.265 $Y2=2.895
r261 65 66 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=12.1 $Y=2.98
+ $X2=11.29 $Y2=2.98
r262 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.205 $Y=2.895
+ $X2=11.29 $Y2=2.98
r263 63 83 8.97325 $w=3.04e-07 $l=2.16852e-07 $layer=LI1_cond $X=11.205 $Y=1.675
+ $X2=11.325 $Y2=1.51
r264 63 64 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=11.205 $Y=1.675
+ $X2=11.205 $Y2=2.895
r265 61 83 13.6447 $w=3.04e-07 $l=4.30465e-07 $layer=LI1_cond $X=11.12 $Y=1.17
+ $X2=11.325 $Y2=1.51
r266 61 62 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=11.12 $Y=1.17
+ $X2=10.435 $Y2=1.17
r267 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.35 $Y=1.085
+ $X2=10.435 $Y2=1.17
r268 59 60 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=10.35 $Y=0.435
+ $X2=10.35 $Y2=1.085
r269 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.265 $Y=0.35
+ $X2=10.35 $Y2=0.435
r270 57 58 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=10.265 $Y=0.35
+ $X2=8.555 $Y2=0.35
r271 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.47 $Y=0.435
+ $X2=8.555 $Y2=0.35
r272 55 56 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.47 $Y=0.435
+ $X2=8.47 $Y2=0.705
r273 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.385 $Y=0.79
+ $X2=8.47 $Y2=0.705
r274 53 54 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=8.385 $Y=0.79
+ $X2=7.31 $Y2=0.79
r275 51 90 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.21 $Y=1.215
+ $X2=7.21 $Y2=1.05
r276 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.21
+ $Y=1.215 $X2=7.21 $Y2=1.215
r277 48 54 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=7.177 $Y=0.875
+ $X2=7.31 $Y2=0.79
r278 48 50 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=7.177 $Y=0.875
+ $X2=7.177 $Y2=1.215
r279 46 80 28.7024 $w=2.63e-07 $l=6.6e-07 $layer=LI1_cond $X=4.627 $Y=2.2
+ $X2=4.627 $Y2=1.54
r280 43 80 6.8764 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=4.567 $Y=1.348
+ $X2=4.567 $Y2=1.54
r281 42 77 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=4.567 $Y=1.062
+ $X2=4.567 $Y2=1.035
r282 42 43 8.56101 $w=3.83e-07 $l=2.86e-07 $layer=LI1_cond $X=4.567 $Y=1.062
+ $X2=4.567 $Y2=1.348
r283 38 70 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=12.265 $Y=2.305
+ $X2=12.265 $Y2=1.865
r284 35 38 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=11.93 $Y=2.38
+ $X2=12.265 $Y2=2.38
r285 33 78 53.9022 $w=6.7e-07 $l=6.75e-07 $layer=POLY_cond $X=5.27 $Y=1.205
+ $X2=4.595 $Y2=1.205
r286 33 34 11.9686 $w=6.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.27 $Y=1.205
+ $X2=5.345 $Y2=1.205
r287 30 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.93 $Y=2.455
+ $X2=11.93 $Y2=2.38
r288 30 32 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.93 $Y=2.455
+ $X2=11.93 $Y2=2.74
r289 29 93 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.42 $Y=0.915
+ $X2=11.42 $Y2=1.345
r290 26 90 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.12 $Y=0.73
+ $X2=7.12 $Y2=1.05
r291 23 26 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=7.12 $Y=0.255
+ $X2=7.12 $Y2=0.73
r292 19 21 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=6.4 $Y=3.06
+ $X2=6.4 $Y2=2.105
r293 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.325 $Y=3.135
+ $X2=6.4 $Y2=3.06
r294 17 18 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=6.325 $Y=3.135
+ $X2=5.42 $Y2=3.135
r295 15 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.045 $Y=0.18
+ $X2=7.12 $Y2=0.255
r296 15 16 833.245 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=7.045 $Y=0.18
+ $X2=5.42 $Y2=0.18
r297 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.345 $Y=3.06
+ $X2=5.42 $Y2=3.135
r298 12 14 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=5.345 $Y=3.06
+ $X2=5.345 $Y2=2.155
r299 11 34 56.3093 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.345 $Y=1.54
+ $X2=5.345 $Y2=1.205
r300 11 14 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=5.345 $Y=1.54
+ $X2=5.345 $Y2=2.155
r301 8 34 56.3093 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.345 $Y=0.87
+ $X2=5.345 $Y2=1.205
r302 8 10 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.345 $Y=0.87
+ $X2=5.345 $Y2=0.54
r303 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.345 $Y=0.255
+ $X2=5.42 $Y2=0.18
r304 7 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.345 $Y=0.255
+ $X2=5.345 $Y2=0.54
r305 2 46 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=2.055 $X2=4.58 $Y2=2.2
r306 1 73 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.19
+ $Y=0.25 $X2=4.33 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_1445_324# 1 2 7 9 11 14 18 22 26 27 29 30
+ 34 36 39 40 43 46 47 49
c140 34 0 1.25205e-19 $X=9.77 $Y=1.435
c141 27 0 1.21132e-19 $X=7.94 $Y=1.57
r142 43 44 20.1468 $w=2.18e-07 $l=3.6e-07 $layer=LI1_cond $X=9.41 $Y=1.095
+ $X2=9.77 $Y2=1.095
r143 40 54 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.8 $Y=1.56
+ $X2=10.8 $Y2=1.725
r144 40 53 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.8 $Y=1.56
+ $X2=10.8 $Y2=1.395
r145 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.775
+ $Y=1.56 $X2=10.775 $Y2=1.56
r146 37 47 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.855 $Y=1.58
+ $X2=9.77 $Y2=1.58
r147 37 39 36.5603 $w=2.88e-07 $l=9.2e-07 $layer=LI1_cond $X=9.855 $Y=1.58
+ $X2=10.775 $Y2=1.58
r148 36 46 3.70735 $w=2.5e-07 $l=1.31031e-07 $layer=LI1_cond $X=9.77 $Y=1.915
+ $X2=9.69 $Y2=2.012
r149 35 47 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.77 $Y=1.725
+ $X2=9.77 $Y2=1.58
r150 35 36 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.77 $Y=1.725
+ $X2=9.77 $Y2=1.915
r151 34 47 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.77 $Y=1.435
+ $X2=9.77 $Y2=1.58
r152 33 44 2.19618 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.77 $Y=1.225
+ $X2=9.77 $Y2=1.095
r153 33 34 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.77 $Y=1.225
+ $X2=9.77 $Y2=1.435
r154 29 46 2.76166 $w=1.7e-07 $l=1.71377e-07 $layer=LI1_cond $X=9.525 $Y=2.025
+ $X2=9.69 $Y2=2.012
r155 29 30 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=9.525 $Y=2.025
+ $X2=8.04 $Y2=2.025
r156 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.94
+ $Y=1.57 $X2=7.94 $Y2=1.57
r157 24 30 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.94 $Y=1.94
+ $X2=8.04 $Y2=2.025
r158 24 26 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=7.94 $Y=1.94
+ $X2=7.94 $Y2=1.57
r159 22 54 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=10.915 $Y=2.315
+ $X2=10.915 $Y2=1.725
r160 18 53 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.915 $Y=0.915
+ $X2=10.915 $Y2=1.395
r161 12 27 39.5234 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=7.69 $Y=1.587
+ $X2=7.94 $Y2=1.587
r162 12 49 32.4387 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.69 $Y=1.587
+ $X2=7.615 $Y2=1.587
r163 12 14 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=7.69 $Y=1.405
+ $X2=7.69 $Y2=0.73
r164 11 49 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.375 $Y=1.695
+ $X2=7.615 $Y2=1.695
r165 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.3 $Y=1.77
+ $X2=7.375 $Y2=1.695
r166 7 9 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.3 $Y=1.77 $X2=7.3
+ $Y2=2.105
r167 2 46 300 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=2 $X=8.835
+ $Y=1.895 $X2=9.69 $Y2=2.08
r168 1 43 182 $w=1.7e-07 $l=9.31316e-07 $layer=licon1_NDIFF $count=1 $X=9.195
+ $Y=0.3 $X2=9.41 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%SET_B 3 7 11 13 16 20 22 24 25 28 31 32 35
+ 40 42
c140 35 0 1.21132e-19 $X=8.67 $Y=1.245
c141 32 0 7.66706e-20 $X=13.2 $Y=1.295
c142 24 0 3.07529e-20 $X=13.055 $Y=1.295
c143 20 0 2.27899e-20 $X=13.485 $Y=2.05
r144 40 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.165 $Y=1.51
+ $X2=13.165 $Y2=1.675
r145 40 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.165 $Y=1.51
+ $X2=13.165 $Y2=1.345
r146 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.165
+ $Y=1.51 $X2=13.165 $Y2=1.51
r147 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=1.245
+ $X2=8.67 $Y2=1.41
r148 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=1.245
+ $X2=8.67 $Y2=1.08
r149 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.67
+ $Y=1.245 $X2=8.67 $Y2=1.245
r150 32 41 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=13.165 $Y=1.295
+ $X2=13.165 $Y2=1.51
r151 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=1.295
+ $X2=13.2 $Y2=1.295
r152 28 36 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8.88 $Y=1.245
+ $X2=8.67 $Y2=1.245
r153 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.295
r154 25 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.025 $Y=1.295
+ $X2=8.88 $Y2=1.295
r155 24 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.055 $Y=1.295
+ $X2=13.2 $Y2=1.295
r156 24 25 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=13.055 $Y=1.295
+ $X2=9.025 $Y2=1.295
r157 22 41 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=13.165 $Y=1.665
+ $X2=13.165 $Y2=1.51
r158 18 20 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=13.255 $Y=2.05
+ $X2=13.485 $Y2=2.05
r159 14 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.485 $Y=2.125
+ $X2=13.485 $Y2=2.05
r160 14 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=13.485 $Y=2.125
+ $X2=13.485 $Y2=2.675
r161 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.255 $Y=1.975
+ $X2=13.255 $Y2=2.05
r162 13 43 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=13.255 $Y=1.975
+ $X2=13.255 $Y2=1.675
r163 11 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.105 $Y=0.915
+ $X2=13.105 $Y2=1.345
r164 7 38 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=8.76 $Y=2.315
+ $X2=8.76 $Y2=1.41
r165 3 37 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=8.685 $Y=0.62
+ $X2=8.685 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_1295_379# 1 2 9 11 12 15 19 21 24 25 26
+ 28 29 30 31 37
c129 12 0 1.25205e-19 $X=9.505 $Y=1.66
r130 37 39 4.0283 $w=3.18e-07 $l=1.05e-07 $layer=LI1_cond $X=9.34 $Y=1.57
+ $X2=9.34 $Y2=1.675
r131 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.34
+ $Y=1.57 $X2=9.34 $Y2=1.57
r132 31 34 4.98819 $w=3.33e-07 $l=1.45e-07 $layer=LI1_cond $X=6.697 $Y=1.96
+ $X2=6.697 $Y2=2.105
r133 31 32 2.92411 $w=3.33e-07 $l=8.5e-08 $layer=LI1_cond $X=6.697 $Y=1.96
+ $X2=6.697 $Y2=1.875
r134 29 39 4.40442 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=1.675
+ $X2=9.34 $Y2=1.675
r135 29 30 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=9.175 $Y=1.675
+ $X2=8.39 $Y2=1.675
r136 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.305 $Y=1.59
+ $X2=8.39 $Y2=1.675
r137 27 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.305 $Y=1.225
+ $X2=8.305 $Y2=1.59
r138 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.22 $Y=1.14
+ $X2=8.305 $Y2=1.225
r139 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.22 $Y=1.14
+ $X2=7.66 $Y2=1.14
r140 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.575 $Y=1.225
+ $X2=7.66 $Y2=1.14
r141 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.575 $Y=1.225
+ $X2=7.575 $Y2=1.875
r142 22 31 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.865 $Y=1.96
+ $X2=6.697 $Y2=1.96
r143 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.49 $Y=1.96
+ $X2=7.575 $Y2=1.875
r144 21 22 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=7.49 $Y=1.96
+ $X2=6.865 $Y2=1.96
r145 19 32 38.2402 $w=3.28e-07 $l=1.095e-06 $layer=LI1_cond $X=6.7 $Y=0.78
+ $X2=6.7 $Y2=1.875
r146 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.905 $Y=1.735
+ $X2=9.905 $Y2=2.315
r147 12 38 38.7444 $w=2.79e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.505 $Y=1.66
+ $X2=9.34 $Y2=1.57
r148 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.83 $Y=1.66
+ $X2=9.905 $Y2=1.735
r149 11 12 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=9.83 $Y=1.66
+ $X2=9.505 $Y2=1.66
r150 7 38 38.0072 $w=2.79e-07 $l=2.91033e-07 $layer=POLY_cond $X=9.12 $Y=1.405
+ $X2=9.34 $Y2=1.57
r151 7 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=9.12 $Y=1.405
+ $X2=9.12 $Y2=0.62
r152 2 34 600 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_PDIFF $count=1 $X=6.475
+ $Y=1.895 $X2=6.695 $Y2=2.105
r153 1 19 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=6.48
+ $Y=0.625 $X2=6.7 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_995_66# 1 2 7 11 13 15 18 19 20 24 25 26
+ 28 29 31 32 36 40 44 48 51 52
c122 51 0 1.9702e-19 $X=5.125 $Y=1.51
c123 24 0 4.60649e-20 $X=11.42 $Y=2.56
c124 15 0 4.10494e-20 $X=6.91 $Y=1.77
r125 49 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.835 $Y=1.51
+ $X2=5.835 $Y2=1.42
r126 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.835
+ $Y=1.51 $X2=5.835 $Y2=1.51
r127 46 51 1.39677 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=5.295 $Y=1.51
+ $X2=5.125 $Y2=1.51
r128 46 48 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.295 $Y=1.51
+ $X2=5.835 $Y2=1.51
r129 42 51 5.10169 $w=3.35e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=1.675
+ $X2=5.125 $Y2=1.51
r130 42 44 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=5.125 $Y=1.675
+ $X2=5.125 $Y2=1.98
r131 38 51 5.10169 $w=3.35e-07 $l=1.67481e-07 $layer=LI1_cond $X=5.12 $Y=1.345
+ $X2=5.125 $Y2=1.51
r132 38 40 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=5.12 $Y=1.345
+ $X2=5.12 $Y2=0.54
r133 34 36 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=11.815 $Y=1.385
+ $X2=11.93 $Y2=1.385
r134 29 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.93 $Y=1.31
+ $X2=11.93 $Y2=1.385
r135 29 31 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.93 $Y=1.31
+ $X2=11.93 $Y2=1.025
r136 27 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.815 $Y=1.46
+ $X2=11.815 $Y2=1.385
r137 27 28 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=11.815 $Y=1.46
+ $X2=11.815 $Y2=1.915
r138 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.74 $Y=1.99
+ $X2=11.815 $Y2=1.915
r139 25 26 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=11.74 $Y=1.99
+ $X2=11.495 $Y2=1.99
r140 22 24 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=11.42 $Y=3.075
+ $X2=11.42 $Y2=2.56
r141 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.42 $Y=2.065
+ $X2=11.495 $Y2=1.99
r142 21 24 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.42 $Y=2.065
+ $X2=11.42 $Y2=2.56
r143 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.345 $Y=3.15
+ $X2=11.42 $Y2=3.075
r144 19 20 2235.66 $w=1.5e-07 $l=4.36e-06 $layer=POLY_cond $X=11.345 $Y=3.15
+ $X2=6.985 $Y2=3.15
r145 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.91 $Y=3.075
+ $X2=6.985 $Y2=3.15
r146 16 18 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=6.91 $Y=3.075
+ $X2=6.91 $Y2=2.105
r147 15 33 86.8103 $w=2.02e-07 $l=3.85681e-07 $layer=POLY_cond $X=6.91 $Y=1.77
+ $X2=6.835 $Y2=1.42
r148 15 18 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.91 $Y=1.77
+ $X2=6.91 $Y2=2.105
r149 14 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.48 $Y=1.42
+ $X2=6.405 $Y2=1.42
r150 13 33 9.80621 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.685 $Y=1.42
+ $X2=6.835 $Y2=1.42
r151 13 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=6.685 $Y=1.42
+ $X2=6.48 $Y2=1.42
r152 9 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.405 $Y=1.345
+ $X2=6.405 $Y2=1.42
r153 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.405 $Y=1.345
+ $X2=6.405 $Y2=0.835
r154 8 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6 $Y=1.42 $X2=5.835
+ $Y2=1.42
r155 7 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.33 $Y=1.42
+ $X2=6.405 $Y2=1.42
r156 7 8 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.33 $Y=1.42 $X2=6
+ $Y2=1.42
r157 2 44 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.99
+ $Y=1.835 $X2=5.13 $Y2=1.98
r158 1 40 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.33 $X2=5.12 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_2449_137# 1 2 7 9 10 11 16 20 24 26 29 32
+ 36 37 38 39 40 43 48 51 55 58 59 62 63 65 66 70 74 76
c186 62 0 2.044e-19 $X=15.635 $Y=2.47
c187 48 0 1.44198e-19 $X=13.7 $Y=2.4
c188 29 0 8.21183e-20 $X=16.755 $Y=1.325
c189 24 0 1.28899e-19 $X=15.8 $Y=0.705
r190 76 77 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=15.74 $Y=1.4
+ $X2=15.74 $Y2=1.325
r191 71 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.74 $Y=1.49
+ $X2=15.74 $Y2=1.655
r192 71 76 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=15.74 $Y=1.49
+ $X2=15.74 $Y2=1.4
r193 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.74
+ $Y=1.49 $X2=15.74 $Y2=1.49
r194 67 70 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=15.635 $Y=1.49
+ $X2=15.74 $Y2=1.49
r195 64 65 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=14.062 $Y=1.085
+ $X2=14.062 $Y2=1.255
r196 61 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.635 $Y=1.655
+ $X2=15.635 $Y2=1.49
r197 61 62 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=15.635 $Y=1.655
+ $X2=15.635 $Y2=2.47
r198 60 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.22 $Y=2.555
+ $X2=14.135 $Y2=2.555
r199 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.55 $Y=2.555
+ $X2=15.635 $Y2=2.47
r200 59 60 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=15.55 $Y=2.555
+ $X2=14.22 $Y2=2.555
r201 58 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.135 $Y=2.47
+ $X2=14.135 $Y2=2.555
r202 58 65 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=14.135 $Y=2.47
+ $X2=14.135 $Y2=1.255
r203 55 64 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=14.03 $Y=0.935
+ $X2=14.03 $Y2=1.085
r204 52 63 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.865 $Y=2.555
+ $X2=13.7 $Y2=2.555
r205 51 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.05 $Y=2.555
+ $X2=14.135 $Y2=2.555
r206 51 52 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=14.05 $Y=2.555
+ $X2=13.865 $Y2=2.555
r207 46 63 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.7 $Y=2.47
+ $X2=13.7 $Y2=2.555
r208 46 48 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=13.7 $Y=2.47 $X2=13.7
+ $Y2=2.4
r209 45 48 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=13.7 $Y=2.29
+ $X2=13.7 $Y2=2.4
r210 43 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.805 $Y=2.125
+ $X2=12.805 $Y2=2.29
r211 43 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.805 $Y=2.125
+ $X2=12.805 $Y2=1.96
r212 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.805
+ $Y=2.125 $X2=12.805 $Y2=2.125
r213 40 45 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=13.535 $Y=2.125
+ $X2=13.7 $Y2=2.29
r214 40 42 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=13.535 $Y=2.125
+ $X2=12.805 $Y2=2.125
r215 37 38 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=16.772 $Y=0.78
+ $X2=16.772 $Y2=0.93
r216 36 37 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=16.79 $Y=0.495
+ $X2=16.79 $Y2=0.78
r217 30 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.755 $Y=1.475
+ $X2=16.755 $Y2=1.4
r218 30 32 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=16.755 $Y=1.475
+ $X2=16.755 $Y2=2.155
r219 29 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.755 $Y=1.325
+ $X2=16.755 $Y2=1.4
r220 29 38 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=16.755 $Y=1.325
+ $X2=16.755 $Y2=0.93
r221 27 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.905 $Y=1.4
+ $X2=15.74 $Y2=1.4
r222 26 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.68 $Y=1.4
+ $X2=16.755 $Y2=1.4
r223 26 27 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=16.68 $Y=1.4
+ $X2=15.905 $Y2=1.4
r224 24 77 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.8 $Y=0.705
+ $X2=15.8 $Y2=1.325
r225 20 79 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=15.77 $Y=2.465
+ $X2=15.77 $Y2=1.655
r226 16 75 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=12.745 $Y=2.74
+ $X2=12.745 $Y2=2.29
r227 12 74 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=12.715 $Y=1.46
+ $X2=12.715 $Y2=1.96
r228 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.64 $Y=1.385
+ $X2=12.715 $Y2=1.46
r229 10 11 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=12.64 $Y=1.385
+ $X2=12.395 $Y2=1.385
r230 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.32 $Y=1.31
+ $X2=12.395 $Y2=1.385
r231 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.32 $Y=1.31
+ $X2=12.32 $Y2=1.025
r232 2 48 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.56
+ $Y=2.255 $X2=13.7 $Y2=2.4
r233 1 55 182 $w=1.7e-07 $l=4.36348e-07 $layer=licon1_NDIFF $count=1 $X=13.77
+ $Y=0.595 $X2=13.99 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_2299_119# 1 2 9 13 17 22 27 28 31 32 33
c98 33 0 1.27581e-19 $X=13.705 $Y=1.435
c99 31 0 1.3679e-19 $X=13.705 $Y=1.6
c100 28 0 4.60649e-20 $X=11.675 $Y=2.12
c101 27 0 2.25888e-20 $X=11.635 $Y=2.415
c102 13 0 7.66706e-20 $X=13.915 $Y=2.675
r103 32 35 1.70922 $w=2.82e-07 $l=1e-08 $layer=POLY_cond $X=13.705 $Y=1.6
+ $X2=13.695 $Y2=1.6
r104 31 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.705 $Y=1.6
+ $X2=13.705 $Y2=1.435
r105 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.705
+ $Y=1.6 $X2=13.705 $Y2=1.6
r106 27 28 12.3448 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=11.675 $Y=2.415
+ $X2=11.675 $Y2=2.12
r107 25 28 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=11.795 $Y=1.165
+ $X2=11.795 $Y2=2.12
r108 24 25 11.0799 $w=4.08e-07 $l=2.5e-07 $layer=LI1_cond $X=11.675 $Y=0.915
+ $X2=11.675 $Y2=1.165
r109 22 24 1.26488 $w=4.08e-07 $l=4.5e-08 $layer=LI1_cond $X=11.675 $Y=0.87
+ $X2=11.675 $Y2=0.915
r110 19 33 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=13.625 $Y=1
+ $X2=13.625 $Y2=1.435
r111 18 24 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=11.88 $Y=0.915
+ $X2=11.675 $Y2=0.915
r112 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.54 $Y=0.915
+ $X2=13.625 $Y2=1
r113 17 18 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=13.54 $Y=0.915
+ $X2=11.88 $Y2=0.915
r114 11 32 35.8936 $w=2.82e-07 $l=2.80624e-07 $layer=POLY_cond $X=13.915
+ $Y=1.765 $X2=13.705 $Y2=1.6
r115 11 13 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=13.915 $Y=1.765
+ $X2=13.915 $Y2=2.675
r116 7 35 17.5183 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.695 $Y=1.435
+ $X2=13.695 $Y2=1.6
r117 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=13.695 $Y=1.435
+ $X2=13.695 $Y2=0.915
r118 2 27 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=11.495
+ $Y=2.14 $X2=11.635 $Y2=2.415
r119 1 22 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=11.495
+ $Y=0.595 $X2=11.635 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_1926_21# 1 2 10 11 12 13 14 17 21 26 30
+ 35 40 41 42 43 44 46 50
c122 42 0 1.28899e-19 $X=14.91 $Y=1.08
c123 30 0 1.14e-19 $X=14.565 $Y=1.62
c124 26 0 1.27581e-19 $X=14.285 $Y=0.67
c125 21 0 1.44198e-19 $X=14.275 $Y=2.675
r126 48 50 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=15.075 $Y=0.995
+ $X2=15.075 $Y2=0.495
r127 44 46 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=14.73 $Y=2.125
+ $X2=15.045 $Y2=2.125
r128 42 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.91 $Y=1.08
+ $X2=15.075 $Y2=0.995
r129 42 43 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=14.91 $Y=1.08
+ $X2=14.73 $Y2=1.08
r130 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.565
+ $Y=1.265 $X2=14.565 $Y2=1.265
r131 38 44 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=14.565 $Y=1.96
+ $X2=14.73 $Y2=2.125
r132 38 40 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=14.565 $Y=1.96
+ $X2=14.565 $Y2=1.265
r133 37 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.565 $Y=1.165
+ $X2=14.73 $Y2=1.08
r134 37 40 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=14.565 $Y=1.165
+ $X2=14.565 $Y2=1.265
r135 35 41 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=14.565 $Y=1.25
+ $X2=14.565 $Y2=1.265
r136 32 35 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=14.285 $Y=1.175
+ $X2=14.565 $Y2=1.175
r137 30 41 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=14.565 $Y=1.62
+ $X2=14.565 $Y2=1.265
r138 27 30 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=14.275 $Y=1.695
+ $X2=14.565 $Y2=1.695
r139 24 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.285 $Y=1.1
+ $X2=14.285 $Y2=1.175
r140 24 26 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=14.285 $Y=1.1
+ $X2=14.285 $Y2=0.67
r141 23 26 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=14.285 $Y=0.255
+ $X2=14.285 $Y2=0.67
r142 19 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.275 $Y=1.77
+ $X2=14.275 $Y2=1.695
r143 19 21 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=14.275 $Y=1.77
+ $X2=14.275 $Y2=2.675
r144 15 17 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=10.295 $Y=1.195
+ $X2=10.295 $Y2=2.315
r145 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.22 $Y=1.12
+ $X2=10.295 $Y2=1.195
r146 13 14 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=10.22 $Y=1.12
+ $X2=9.78 $Y2=1.12
r147 11 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.21 $Y=0.18
+ $X2=14.285 $Y2=0.255
r148 11 12 2271.55 $w=1.5e-07 $l=4.43e-06 $layer=POLY_cond $X=14.21 $Y=0.18
+ $X2=9.78 $Y2=0.18
r149 8 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.705 $Y=1.045
+ $X2=9.78 $Y2=1.12
r150 8 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.705 $Y=1.045
+ $X2=9.705 $Y2=0.65
r151 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.705 $Y=0.255
+ $X2=9.78 $Y2=0.18
r152 7 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.705 $Y=0.255
+ $X2=9.705 $Y2=0.65
r153 2 46 600 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=14.905
+ $Y=1.835 $X2=15.045 $Y2=2.125
r154 1 50 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=14.93
+ $Y=0.285 $X2=15.075 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%RESET_B 3 7 9 12 13
c38 12 0 1.35877e-19 $X=15.2 $Y=1.51
r39 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.2 $Y=1.51
+ $X2=15.2 $Y2=1.675
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.2 $Y=1.51
+ $X2=15.2 $Y2=1.345
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.2
+ $Y=1.51 $X2=15.2 $Y2=1.51
r42 9 13 4.96191 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=15.185 $Y=1.665
+ $X2=15.185 $Y2=1.51
r43 7 14 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=15.29 $Y=0.495
+ $X2=15.29 $Y2=1.345
r44 3 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=15.26 $Y=2.155
+ $X2=15.26 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_3279_367# 1 2 9 13 17 21 25 26 28
c53 21 0 1.40041e-19 $X=16.54 $Y=1.98
r54 26 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=17.205 $Y=1.47
+ $X2=17.205 $Y2=1.635
r55 26 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=17.205 $Y=1.47
+ $X2=17.205 $Y2=1.305
r56 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.205
+ $Y=1.47 $X2=17.205 $Y2=1.47
r57 23 28 0.0443336 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=16.705 $Y=1.47
+ $X2=16.58 $Y2=1.47
r58 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=16.705 $Y=1.47
+ $X2=17.205 $Y2=1.47
r59 19 28 6.95506 $w=2.27e-07 $l=1.65e-07 $layer=LI1_cond $X=16.58 $Y=1.635
+ $X2=16.58 $Y2=1.47
r60 19 21 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=16.58 $Y=1.635
+ $X2=16.58 $Y2=1.98
r61 15 28 6.95506 $w=2.27e-07 $l=1.76125e-07 $layer=LI1_cond $X=16.557 $Y=1.305
+ $X2=16.58 $Y2=1.47
r62 15 17 43.8226 $w=2.03e-07 $l=8.1e-07 $layer=LI1_cond $X=16.557 $Y=1.305
+ $X2=16.557 $Y2=0.495
r63 13 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=17.265 $Y=2.465
+ $X2=17.265 $Y2=1.635
r64 9 30 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=17.265 $Y=0.705
+ $X2=17.265 $Y2=1.305
r65 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.395
+ $Y=1.835 $X2=16.54 $Y2=1.98
r66 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=16.43
+ $Y=0.285 $X2=16.575 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_27_474# 1 2 9 11 12 14 15 16 19
c46 16 0 1.17915e-19 $X=1.145 $Y=2.98
r47 17 19 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.93 $Y=2.895
+ $X2=1.93 $Y2=2.515
r48 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.765 $Y=2.98
+ $X2=1.93 $Y2=2.895
r49 15 16 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.765 $Y=2.98
+ $X2=1.145 $Y2=2.98
r50 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.895
+ $X2=1.145 $Y2=2.98
r51 13 14 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.06 $Y=2.235
+ $X2=1.06 $Y2=2.895
r52 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=2.15
+ $X2=1.06 $Y2=2.235
r53 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.975 $Y=2.15
+ $X2=0.365 $Y2=2.15
r54 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=2.235
+ $X2=0.365 $Y2=2.15
r55 7 9 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=2.235 $X2=0.24
+ $Y2=2.515
r56 2 19 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.79
+ $Y=2.37 $X2=1.93 $Y2=2.515
r57 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.37 $X2=0.28 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 61 65 69 74 75 77 78 80 81 83 84 85 87 102 106 121 132 136 143 144 147 150
+ 153 156 159 162
r184 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r185 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r186 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r187 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r188 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r189 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r190 144 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=17.04 $Y2=3.33
r191 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r192 141 162 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.135 $Y=3.33
+ $X2=17.01 $Y2=3.33
r193 141 143 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=17.135 $Y=3.33
+ $X2=17.52 $Y2=3.33
r194 140 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=17.04 $Y2=3.33
r195 140 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=15.6 $Y2=3.33
r196 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r197 137 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.72 $Y=3.33
+ $X2=15.555 $Y2=3.33
r198 137 139 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=15.72 $Y=3.33
+ $X2=16.56 $Y2=3.33
r199 136 162 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.885 $Y=3.33
+ $X2=17.01 $Y2=3.33
r200 136 139 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=16.885 $Y=3.33
+ $X2=16.56 $Y2=3.33
r201 135 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=15.6 $Y2=3.33
r202 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r203 132 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.39 $Y=3.33
+ $X2=15.555 $Y2=3.33
r204 132 134 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=15.39 $Y=3.33
+ $X2=15.12 $Y2=3.33
r205 131 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=15.12 $Y2=3.33
r206 131 157 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.2 $Y2=3.33
r207 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r208 128 156 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.355 $Y=3.33
+ $X2=13.23 $Y2=3.33
r209 128 130 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=13.355 $Y=3.33
+ $X2=14.16 $Y2=3.33
r210 127 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r211 126 127 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r212 124 127 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=12.72 $Y2=3.33
r213 123 126 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=10.8 $Y=3.33
+ $X2=12.72 $Y2=3.33
r214 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r215 121 156 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.105 $Y=3.33
+ $X2=13.23 $Y2=3.33
r216 121 126 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.105 $Y=3.33
+ $X2=12.72 $Y2=3.33
r217 120 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r218 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r219 116 119 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r220 114 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.63 $Y=3.33
+ $X2=8.465 $Y2=3.33
r221 114 116 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.63 $Y=3.33
+ $X2=8.88 $Y2=3.33
r222 113 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r223 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 110 113 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r225 110 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r226 109 112 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r227 109 110 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r228 107 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=3.33
+ $X2=5.635 $Y2=3.33
r229 107 109 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.8 $Y=3.33 $X2=6
+ $Y2=3.33
r230 106 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.3 $Y=3.33
+ $X2=8.465 $Y2=3.33
r231 106 112 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.3 $Y=3.33
+ $X2=7.92 $Y2=3.33
r232 105 151 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r233 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r234 102 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=5.635 $Y2=3.33
r235 102 104 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=4.08 $Y2=3.33
r236 101 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r237 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r238 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r239 97 100 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r240 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r241 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r242 95 148 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.72 $Y2=3.33
r243 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r244 92 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.67 $Y2=3.33
r245 92 94 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=2.16 $Y2=3.33
r246 90 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r247 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r248 87 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.67 $Y2=3.33
r249 87 89 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.24 $Y2=3.33
r250 85 120 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r251 85 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r252 85 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r253 83 130 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=14.325 $Y=3.33
+ $X2=14.16 $Y2=3.33
r254 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.325 $Y=3.33
+ $X2=14.49 $Y2=3.33
r255 82 134 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=14.655 $Y=3.33
+ $X2=15.12 $Y2=3.33
r256 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.655 $Y=3.33
+ $X2=14.49 $Y2=3.33
r257 80 119 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=10.345 $Y=3.33
+ $X2=10.32 $Y2=3.33
r258 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.345 $Y=3.33
+ $X2=10.51 $Y2=3.33
r259 79 123 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.8 $Y2=3.33
r260 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.51 $Y2=3.33
r261 77 100 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.6 $Y2=3.33
r262 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.88 $Y2=3.33
r263 76 104 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=4.08 $Y2=3.33
r264 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.88 $Y2=3.33
r265 74 94 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.16 $Y2=3.33
r266 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.48 $Y2=3.33
r267 73 97 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.64 $Y2=3.33
r268 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.48 $Y2=3.33
r269 69 72 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=17.01 $Y=1.98
+ $X2=17.01 $Y2=2.465
r270 67 162 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=17.01 $Y=3.245
+ $X2=17.01 $Y2=3.33
r271 67 72 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=17.01 $Y=3.245
+ $X2=17.01 $Y2=2.465
r272 63 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.555 $Y=3.245
+ $X2=15.555 $Y2=3.33
r273 63 65 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=15.555 $Y=3.245
+ $X2=15.555 $Y2=2.925
r274 59 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.49 $Y=3.245
+ $X2=14.49 $Y2=3.33
r275 59 61 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=14.49 $Y=3.245
+ $X2=14.49 $Y2=2.925
r276 55 156 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.23 $Y=3.245
+ $X2=13.23 $Y2=3.33
r277 55 57 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=13.23 $Y=3.245
+ $X2=13.23 $Y2=2.79
r278 51 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.51 $Y=3.245
+ $X2=10.51 $Y2=3.33
r279 51 53 41.034 $w=3.28e-07 $l=1.175e-06 $layer=LI1_cond $X=10.51 $Y=3.245
+ $X2=10.51 $Y2=2.07
r280 47 153 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=3.33
r281 47 49 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=2.52
r282 43 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=3.245
+ $X2=5.635 $Y2=3.33
r283 43 45 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=5.635 $Y=3.245
+ $X2=5.635 $Y2=2.84
r284 39 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=3.33
r285 39 41 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=2.39
r286 35 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=3.245
+ $X2=2.48 $Y2=3.33
r287 35 37 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=2.48 $Y=3.245
+ $X2=2.48 $Y2=2.2
r288 31 147 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=3.245
+ $X2=0.67 $Y2=3.33
r289 31 33 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=0.67 $Y=3.245
+ $X2=0.67 $Y2=2.72
r290 10 72 300 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_PDIFF $count=2 $X=16.83
+ $Y=1.835 $X2=17.05 $Y2=2.465
r291 10 69 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=16.83
+ $Y=1.835 $X2=17.05 $Y2=1.98
r292 9 65 600 $w=1.7e-07 $l=1.19495e-06 $layer=licon1_PDIFF $count=1 $X=15.335
+ $Y=1.835 $X2=15.555 $Y2=2.925
r293 8 61 600 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=1 $X=14.35
+ $Y=2.255 $X2=14.49 $Y2=2.925
r294 7 57 600 $w=1.7e-07 $l=5.65243e-07 $layer=licon1_PDIFF $count=1 $X=12.82
+ $Y=2.53 $X2=13.27 $Y2=2.79
r295 6 53 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=10.37
+ $Y=1.895 $X2=10.51 $Y2=2.07
r296 5 49 600 $w=1.7e-07 $l=1.36724e-06 $layer=licon1_PDIFF $count=1 $X=7.375
+ $Y=1.895 $X2=8.465 $Y2=2.52
r297 4 45 600 $w=1.7e-07 $l=1.10729e-06 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.835 $X2=5.635 $Y2=2.84
r298 3 41 600 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=1 $X=3.735
+ $Y=2.055 $X2=3.88 $Y2=2.39
r299 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.34
+ $Y=2.055 $X2=2.48 $Y2=2.2
r300 1 33 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.37 $X2=0.71 $Y2=2.72
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_200_119# 1 2 3 4 15 17 18 21 23 24 26 28
+ 29 32 33 34 36 37 38 40 41 42 44 45 46 47 50 53 54 56
c170 26 0 1.7805e-19 $X=2.085 $Y=1.685
r171 56 58 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.19 $Y=0.835
+ $X2=6.19 $Y2=1.065
r172 54 58 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=6.265 $Y=1.875
+ $X2=6.265 $Y2=1.065
r173 48 50 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.185 $Y=2.325
+ $X2=6.185 $Y2=2.105
r174 47 54 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.185 $Y=2.04
+ $X2=6.185 $Y2=1.875
r175 47 50 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=6.185 $Y=2.04
+ $X2=6.185 $Y2=2.105
r176 45 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.02 $Y=2.41
+ $X2=6.185 $Y2=2.325
r177 45 46 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.02 $Y=2.41
+ $X2=5.29 $Y2=2.41
r178 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.205 $Y=2.495
+ $X2=5.29 $Y2=2.41
r179 43 44 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.205 $Y=2.495
+ $X2=5.205 $Y2=2.895
r180 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.12 $Y=2.98
+ $X2=5.205 $Y2=2.895
r181 41 42 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=5.12 $Y=2.98
+ $X2=4.315 $Y2=2.98
r182 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.23 $Y=2.895
+ $X2=4.315 $Y2=2.98
r183 39 40 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.23 $Y=1.89
+ $X2=4.23 $Y2=2.895
r184 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.145 $Y=1.805
+ $X2=4.23 $Y2=1.89
r185 37 38 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.145 $Y=1.805
+ $X2=3.615 $Y2=1.805
r186 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.53 $Y=1.89
+ $X2=3.615 $Y2=1.805
r187 35 36 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=3.53 $Y=1.89
+ $X2=3.53 $Y2=2.895
r188 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=2.98
+ $X2=3.53 $Y2=2.895
r189 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.445 $Y=2.98
+ $X2=2.915 $Y2=2.98
r190 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.83 $Y=2.895
+ $X2=2.915 $Y2=2.98
r191 31 32 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=2.83 $Y=1.855
+ $X2=2.83 $Y2=2.895
r192 30 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=1.77
+ $X2=2.085 $Y2=1.77
r193 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.745 $Y=1.77
+ $X2=2.83 $Y2=1.855
r194 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.745 $Y=1.77
+ $X2=2.17 $Y2=1.77
r195 27 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=1.855
+ $X2=2.085 $Y2=1.77
r196 27 28 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.085 $Y=1.855
+ $X2=2.085 $Y2=2
r197 26 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=1.685
+ $X2=2.085 $Y2=1.77
r198 25 26 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=2.085 $Y=0.63
+ $X2=2.085 $Y2=1.685
r199 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2 $Y=2.085
+ $X2=2.085 $Y2=2
r200 23 24 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2 $Y=2.085
+ $X2=1.585 $Y2=2.085
r201 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.46 $Y=2.17
+ $X2=1.585 $Y2=2.085
r202 19 21 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=1.46 $Y=2.17
+ $X2=1.46 $Y2=2.53
r203 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2 $Y=0.545
+ $X2=2.085 $Y2=0.63
r204 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2 $Y=0.545 $X2=1.31
+ $Y2=0.545
r205 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.145 $Y=0.63
+ $X2=1.31 $Y2=0.545
r206 13 15 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.145 $Y=0.63
+ $X2=1.145 $Y2=0.805
r207 4 50 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.895 $X2=6.185 $Y2=2.105
r208 3 21 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=2.37 $X2=1.5 $Y2=2.53
r209 2 56 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.045
+ $Y=0.625 $X2=6.19 $Y2=0.835
r210 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.595 $X2=1.145 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%Q_N 1 2 9 13 14 15 16 23 33
c29 33 0 8.21183e-20 $X=16.077 $Y=1.835
r30 21 35 0.389558 $w=3.53e-07 $l=1.2e-08 $layer=LI1_cond $X=16.077 $Y=2.012
+ $X2=16.077 $Y2=2
r31 21 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=16.077 $Y=2.012
+ $X2=16.077 $Y2=2.035
r32 16 30 4.0579 $w=3.53e-07 $l=1.25e-07 $layer=LI1_cond $X=16.077 $Y=2.775
+ $X2=16.077 $Y2=2.9
r33 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=16.077 $Y=2.405
+ $X2=16.077 $Y2=2.775
r34 14 35 0.6168 $w=3.53e-07 $l=1.9e-08 $layer=LI1_cond $X=16.077 $Y=1.981
+ $X2=16.077 $Y2=2
r35 14 33 7.88226 $w=3.53e-07 $l=1.46e-07 $layer=LI1_cond $X=16.077 $Y=1.981
+ $X2=16.077 $Y2=1.835
r36 14 15 11.005 $w=3.53e-07 $l=3.39e-07 $layer=LI1_cond $X=16.077 $Y=2.066
+ $X2=16.077 $Y2=2.405
r37 14 23 1.00636 $w=3.53e-07 $l=3.1e-08 $layer=LI1_cond $X=16.077 $Y=2.066
+ $X2=16.077 $Y2=2.035
r38 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.17 $Y=1.145
+ $X2=16.17 $Y2=1.835
r39 7 13 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=16.052 $Y=0.943
+ $X2=16.052 $Y2=1.145
r40 7 9 14.5976 $w=4.03e-07 $l=5.13e-07 $layer=LI1_cond $X=16.052 $Y=0.943
+ $X2=16.052 $Y2=0.43
r41 2 35 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=15.845
+ $Y=1.835 $X2=15.985 $Y2=2
r42 2 30 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=15.845
+ $Y=1.835 $X2=15.985 $Y2=2.9
r43 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.875
+ $Y=0.285 $X2=16.015 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%Q 1 2 9 14 15 16 17 23 29
r25 21 29 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=17.492 $Y=0.948
+ $X2=17.492 $Y2=0.925
r26 17 31 7.88226 $w=3.53e-07 $l=1.46e-07 $layer=LI1_cond $X=17.492 $Y=0.979
+ $X2=17.492 $Y2=1.125
r27 17 21 1.00636 $w=3.53e-07 $l=3.1e-08 $layer=LI1_cond $X=17.492 $Y=0.979
+ $X2=17.492 $Y2=0.948
r28 17 29 1.00636 $w=3.53e-07 $l=3.1e-08 $layer=LI1_cond $X=17.492 $Y=0.894
+ $X2=17.492 $Y2=0.925
r29 16 17 11.005 $w=3.53e-07 $l=3.39e-07 $layer=LI1_cond $X=17.492 $Y=0.555
+ $X2=17.492 $Y2=0.894
r30 16 23 4.0579 $w=3.53e-07 $l=1.25e-07 $layer=LI1_cond $X=17.492 $Y=0.555
+ $X2=17.492 $Y2=0.43
r31 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=17.585 $Y=1.815
+ $X2=17.585 $Y2=1.125
r32 14 15 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=17.492 $Y=1.98
+ $X2=17.492 $Y2=1.815
r33 7 14 0.389558 $w=3.53e-07 $l=1.2e-08 $layer=LI1_cond $X=17.492 $Y=1.992
+ $X2=17.492 $Y2=1.98
r34 7 9 29.4766 $w=3.53e-07 $l=9.08e-07 $layer=LI1_cond $X=17.492 $Y=1.992
+ $X2=17.492 $Y2=2.9
r35 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=17.34
+ $Y=1.835 $X2=17.48 $Y2=1.98
r36 2 9 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=17.34
+ $Y=1.835 $X2=17.48 $Y2=2.9
r37 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.34
+ $Y=0.285 $X2=17.48 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 52 56 60 66 69 70 72 73 74 76 88 92 97 105 118 119 125 128 131 134 137 140
r173 140 141 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r174 137 138 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r175 135 138 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=12.72 $Y2=0
r176 134 135 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r177 131 132 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r178 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r179 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r180 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r181 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r182 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.52 $Y2=0
r183 116 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=15.6 $Y2=0
r184 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r185 113 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.67 $Y=0
+ $X2=15.545 $Y2=0
r186 113 115 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=15.67 $Y=0
+ $X2=16.56 $Y2=0
r187 112 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=15.6 $Y2=0
r188 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r189 109 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=15.12 $Y2=0
r190 109 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r191 108 111 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=13.2 $Y=0
+ $X2=15.12 $Y2=0
r192 108 109 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r193 106 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=12.81 $Y2=0
r194 106 108 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=13.2 $Y2=0
r195 105 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.42 $Y=0
+ $X2=15.545 $Y2=0
r196 105 111 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=15.42 $Y=0
+ $X2=15.12 $Y2=0
r197 104 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r198 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r199 101 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r200 100 103 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r201 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r202 98 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=8.04 $Y2=0
r203 98 100 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=8.4 $Y2=0
r204 97 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.615 $Y=0
+ $X2=10.74 $Y2=0
r205 97 103 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.615 $Y=0
+ $X2=10.32 $Y2=0
r206 96 132 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r207 96 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r208 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r209 93 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=0
+ $X2=5.63 $Y2=0
r210 93 95 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=6
+ $Y2=0
r211 92 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=0
+ $X2=8.04 $Y2=0
r212 92 95 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=7.875 $Y=0 $X2=6
+ $Y2=0
r213 91 129 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.52 $Y2=0
r214 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r215 88 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=5.63 $Y2=0
r216 88 90 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=4.08 $Y2=0
r217 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r218 87 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r219 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r220 84 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=0
+ $X2=2.515 $Y2=0
r221 84 86 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=3.6
+ $Y2=0
r222 83 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r223 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r224 80 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r225 80 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r226 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r227 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r228 77 122 4.64823 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.242 $Y2=0
r229 77 79 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.72 $Y2=0
r230 76 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0
+ $X2=2.515 $Y2=0
r231 76 82 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.16
+ $Y2=0
r232 74 104 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r233 74 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r234 72 115 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=16.84 $Y=0
+ $X2=16.56 $Y2=0
r235 72 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.84 $Y=0
+ $X2=16.965 $Y2=0
r236 71 118 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=17.09 $Y=0
+ $X2=17.52 $Y2=0
r237 71 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.09 $Y=0
+ $X2=16.965 $Y2=0
r238 69 86 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.6
+ $Y2=0
r239 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.82
+ $Y2=0
r240 68 90 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.985 $Y=0 $X2=4.08
+ $Y2=0
r241 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=3.82
+ $Y2=0
r242 64 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.965 $Y=0.085
+ $X2=16.965 $Y2=0
r243 64 66 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=16.965 $Y=0.085
+ $X2=16.965 $Y2=0.495
r244 60 62 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=15.545 $Y=0.43
+ $X2=15.545 $Y2=0.98
r245 58 140 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.545 $Y=0.085
+ $X2=15.545 $Y2=0
r246 58 60 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=15.545 $Y=0.085
+ $X2=15.545 $Y2=0.43
r247 54 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.81 $Y=0.085
+ $X2=12.81 $Y2=0
r248 54 56 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=12.81 $Y=0.085
+ $X2=12.81 $Y2=0.485
r249 53 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.865 $Y=0
+ $X2=10.74 $Y2=0
r250 52 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.645 $Y=0
+ $X2=12.81 $Y2=0
r251 52 53 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=12.645 $Y=0
+ $X2=10.865 $Y2=0
r252 48 134 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=0.085
+ $X2=10.74 $Y2=0
r253 48 50 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=10.74 $Y=0.085
+ $X2=10.74 $Y2=0.74
r254 44 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=0.085
+ $X2=8.04 $Y2=0
r255 44 46 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.04 $Y=0.085
+ $X2=8.04 $Y2=0.36
r256 40 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.63 $Y=0.085
+ $X2=5.63 $Y2=0
r257 40 42 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.63 $Y=0.085
+ $X2=5.63 $Y2=0.54
r258 36 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=0.085
+ $X2=3.82 $Y2=0
r259 36 38 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=3.82 $Y=0.085
+ $X2=3.82 $Y2=0.46
r260 32 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0
r261 32 34 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0.785
r262 28 122 3.11795 $w=3.3e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.242 $Y2=0
r263 28 30 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.32 $Y2=0.805
r264 9 66 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=16.865
+ $Y=0.285 $X2=17.005 $Y2=0.495
r265 8 62 182 $w=1.7e-07 $l=7.97449e-07 $layer=licon1_NDIFF $count=1 $X=15.365
+ $Y=0.285 $X2=15.585 $Y2=0.98
r266 8 60 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=15.365
+ $Y=0.285 $X2=15.585 $Y2=0.43
r267 7 56 182 $w=1.7e-07 $l=5.56035e-07 $layer=licon1_NDIFF $count=1 $X=12.395
+ $Y=0.815 $X2=12.81 $Y2=0.485
r268 6 50 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=10.555
+ $Y=0.595 $X2=10.7 $Y2=0.74
r269 5 46 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=7.765
+ $Y=0.52 $X2=8.04 $Y2=0.36
r270 4 42 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=5.42
+ $Y=0.33 $X2=5.63 $Y2=0.54
r271 3 38 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.675
+ $Y=0.25 $X2=3.82 $Y2=0.46
r272 2 34 182 $w=1.7e-07 $l=3.88555e-07 $layer=licon1_NDIFF $count=1 $X=2.21
+ $Y=0.595 $X2=2.515 $Y2=0.785
r273 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.595 $X2=0.32 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_1752_60# 1 2 12 14 15
r25 14 15 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.92 $Y=0.745
+ $X2=9.755 $Y2=0.745
r26 12 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.065 $Y=0.7
+ $X2=9.755 $Y2=0.7
r27 10 12 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=8.9 $Y=0.757
+ $X2=9.065 $Y2=0.757
r28 2 14 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=9.78
+ $Y=0.33 $X2=9.92 $Y2=0.705
r29 1 10 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=8.76
+ $Y=0.3 $X2=8.9 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_1%A_2636_119# 1 2 7 11 13
r32 13 16 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=13.4 $Y=0.35
+ $X2=13.4 $Y2=0.485
r33 9 11 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=14.5 $Y=0.435
+ $X2=14.5 $Y2=0.57
r34 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.565 $Y=0.35
+ $X2=13.4 $Y2=0.35
r35 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.335 $Y=0.35
+ $X2=14.5 $Y2=0.435
r36 7 8 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=14.335 $Y=0.35
+ $X2=13.565 $Y2=0.35
r37 2 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=14.36
+ $Y=0.35 $X2=14.5 $Y2=0.57
r38 1 16 182 $w=1.7e-07 $l=2.69444e-07 $layer=licon1_NDIFF $count=1 $X=13.18
+ $Y=0.595 $X2=13.4 $Y2=0.485
.ends

