* File: sky130_fd_sc_lp__a32oi_4.spice
* Created: Fri Aug 28 10:02:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32oi_4.pex.spice"
.subckt sky130_fd_sc_lp__a32oi_4  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B2_M1002_g N_A_28_47#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1002_d N_B2_M1013_g N_A_28_47#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_B2_M1016_g N_A_28_47#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1025 N_VGND_M1016_d N_B2_M1025_g N_A_28_47#_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1010 N_Y_M1010_d N_B1_M1010_g N_A_28_47#_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1023 N_Y_M1010_d N_B1_M1023_g N_A_28_47#_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1024 N_Y_M1024_d N_B1_M1024_g N_A_28_47#_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1038 N_Y_M1024_d N_B1_M1038_g N_A_28_47#_M1038_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A1_M1005_g N_A_840_47#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1014 N_Y_M1005_d N_A1_M1014_g N_A_840_47#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1027 N_Y_M1027_d N_A1_M1027_g N_A_840_47#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1037 N_Y_M1027_d N_A1_M1037_g N_A_840_47#_M1037_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1009 N_A_840_47#_M1037_s N_A2_M1009_g N_A_1267_47#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1028 N_A_840_47#_M1028_d N_A2_M1028_g N_A_1267_47#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1030 N_A_840_47#_M1028_d N_A2_M1030_g N_A_1267_47#_M1030_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1035 N_A_840_47#_M1035_d N_A2_M1035_g N_A_1267_47#_M1030_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A3_M1008_g N_A_1267_47#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A3_M1011_g N_A_1267_47#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1011_d N_A3_M1031_g N_A_1267_47#_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1036 N_VGND_M1036_d N_A3_M1036_g N_A_1267_47#_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_42_367#_M1006_d N_B2_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75009.2 A=0.189 P=2.82 MULT=1
MM1020 N_A_42_367#_M1020_d N_B2_M1020_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75008.7 A=0.189 P=2.82 MULT=1
MM1021 N_A_42_367#_M1020_d N_B2_M1021_g N_Y_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75008.3 A=0.189 P=2.82 MULT=1
MM1032 N_A_42_367#_M1032_d N_B2_M1032_g N_Y_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75007.9 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_42_367#_M1032_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75007.4 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1001_d N_B1_M1015_g N_A_42_367#_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3 SB=75007
+ A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1019_d N_B1_M1019_g N_A_42_367#_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75006.6 A=0.189 P=2.82 MULT=1
MM1033 N_Y_M1019_d N_B1_M1033_g N_A_42_367#_M1033_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2457 PD=1.54 PS=1.65 NRD=0 NRS=8.5892 M=1 R=8.4 SA=75003.2
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_42_367#_M1033_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2457 PD=1.54 PS=1.65 NRD=0 NRS=8.5892 M=1 R=8.4 SA=75003.7
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1003_d N_A1_M1012_g N_A_42_367#_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1034 N_VPWR_M1034_d N_A1_M1034_g N_A_42_367#_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.1764 PD=1.88 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75004.8 A=0.189 P=2.82 MULT=1
MM1039 N_VPWR_M1034_d N_A1_M1039_g N_A_42_367#_M1039_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.1764 PD=1.88 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4 SB=75004
+ A=0.189 P=2.82 MULT=1
MM1004 N_A_42_367#_M1039_s N_A2_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4032 PD=1.54 PS=1.9 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8 SB=75003.6
+ A=0.189 P=2.82 MULT=1
MM1017 N_A_42_367#_M1017_d N_A2_M1017_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4032 PD=1.54 PS=1.9 NRD=0 NRS=0 M=1 R=8.4 SA=75006.6 SB=75002.8
+ A=0.189 P=2.82 MULT=1
MM1022 N_A_42_367#_M1017_d N_A2_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007 SB=75002.3
+ A=0.189 P=2.82 MULT=1
MM1029 N_A_42_367#_M1029_d N_A2_M1029_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.4
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A3_M1000_g N_A_42_367#_M1029_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1000_d N_A3_M1007_g N_A_42_367#_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A3_M1018_g N_A_42_367#_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.7
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1018_d N_A3_M1026_g N_A_42_367#_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75009.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=20.4031 P=25.61
c_133 VPB 0 1.99728e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a32oi_4.pxi.spice"
*
.ends
*
*
