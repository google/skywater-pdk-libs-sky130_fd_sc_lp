* File: sky130_fd_sc_lp__a21boi_1.pxi.spice
* Created: Wed Sep  2 09:19:18 2020
* 
x_PM_SKY130_FD_SC_LP__A21BOI_1%B1_N N_B1_N_c_60_n N_B1_N_M1001_g N_B1_N_c_61_n
+ N_B1_N_c_62_n N_B1_N_M1002_g N_B1_N_c_64_n N_B1_N_c_69_n B1_N B1_N B1_N B1_N
+ N_B1_N_c_66_n PM_SKY130_FD_SC_LP__A21BOI_1%B1_N
x_PM_SKY130_FD_SC_LP__A21BOI_1%A_27_508# N_A_27_508#_M1002_s N_A_27_508#_M1001_s
+ N_A_27_508#_c_100_n N_A_27_508#_M1004_g N_A_27_508#_M1000_g
+ N_A_27_508#_c_103_n N_A_27_508#_c_110_n N_A_27_508#_c_111_n
+ N_A_27_508#_c_112_n N_A_27_508#_c_104_n N_A_27_508#_c_105_n
+ N_A_27_508#_c_106_n N_A_27_508#_c_107_n N_A_27_508#_c_108_n
+ PM_SKY130_FD_SC_LP__A21BOI_1%A_27_508#
x_PM_SKY130_FD_SC_LP__A21BOI_1%A1 N_A1_M1005_g N_A1_M1006_g A1 A1 A1
+ N_A1_c_174_n N_A1_c_175_n PM_SKY130_FD_SC_LP__A21BOI_1%A1
x_PM_SKY130_FD_SC_LP__A21BOI_1%A2 N_A2_M1007_g N_A2_M1003_g A2 N_A2_c_210_n
+ N_A2_c_211_n PM_SKY130_FD_SC_LP__A21BOI_1%A2
x_PM_SKY130_FD_SC_LP__A21BOI_1%VPWR N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_c_232_n
+ N_VPWR_c_233_n VPWR N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n
+ N_VPWR_c_231_n N_VPWR_c_238_n N_VPWR_c_239_n PM_SKY130_FD_SC_LP__A21BOI_1%VPWR
x_PM_SKY130_FD_SC_LP__A21BOI_1%Y N_Y_M1004_d N_Y_M1000_s N_Y_c_268_n N_Y_c_269_n
+ Y Y Y Y Y PM_SKY130_FD_SC_LP__A21BOI_1%Y
x_PM_SKY130_FD_SC_LP__A21BOI_1%A_302_367# N_A_302_367#_M1000_d
+ N_A_302_367#_M1003_d N_A_302_367#_c_305_n N_A_302_367#_c_301_n
+ N_A_302_367#_c_302_n N_A_302_367#_c_303_n
+ PM_SKY130_FD_SC_LP__A21BOI_1%A_302_367#
x_PM_SKY130_FD_SC_LP__A21BOI_1%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_c_326_n
+ N_VGND_c_327_n N_VGND_c_328_n VGND N_VGND_c_329_n N_VGND_c_330_n
+ N_VGND_c_331_n N_VGND_c_332_n PM_SKY130_FD_SC_LP__A21BOI_1%VGND
cc_1 VNB N_B1_N_c_60_n 0.00179801f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.915
cc_2 VNB N_B1_N_c_61_n 0.0318404f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.03
cc_3 VNB N_B1_N_c_62_n 0.0208611f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.03
cc_4 VNB N_B1_N_M1002_g 0.0336845f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.445
cc_5 VNB N_B1_N_c_64_n 0.0185589f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.625
cc_6 VNB B1_N 0.0382451f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_B1_N_c_66_n 0.0304658f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_8 VNB N_A_27_508#_c_100_n 0.0193903f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.03
cc_9 VNB N_A_27_508#_M1004_g 0.0280748f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.445
cc_10 VNB N_A_27_508#_M1000_g 0.00849918f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.625
cc_11 VNB N_A_27_508#_c_103_n 0.0117885f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.99
cc_12 VNB N_A_27_508#_c_104_n 0.00339171f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_13 VNB N_A_27_508#_c_105_n 0.00134123f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=0.925
cc_14 VNB N_A_27_508#_c_106_n 0.0138104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_508#_c_107_n 0.0104285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_508#_c_108_n 0.0251717f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.035
cc_17 VNB N_A1_M1006_g 0.00803106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A1 0.0060088f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.445
cc_19 VNB N_A1_c_174_n 0.0319795f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.625
cc_20 VNB N_A1_c_175_n 0.0177062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_M1003_g 0.0119208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A2 0.0157783f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.03
cc_23 VNB N_A2_c_210_n 0.0375403f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.445
cc_24 VNB N_A2_c_211_n 0.022539f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_25 VNB N_VPWR_c_231_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_268_n 0.0087853f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.03
cc_27 VNB N_Y_c_269_n 0.00283101f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.955
cc_28 VNB Y 0.00263343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_326_n 0.00510685f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.955
cc_30 VNB N_VGND_c_327_n 0.0106846f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.445
cc_31 VNB N_VGND_c_328_n 0.0331498f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_32 VNB N_VGND_c_329_n 0.0303401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_330_n 0.0314948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_VGND_c_331_n 0.00471252f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_35 VNB N_VGND_c_332_n 0.174582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B1_N_c_60_n 0.0174045f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.915
cc_37 VPB N_B1_N_M1001_g 0.0519516f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.75
cc_38 VPB N_B1_N_c_69_n 0.021503f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.99
cc_39 VPB B1_N 0.0207553f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_40 VPB N_A_27_508#_M1000_g 0.0234061f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.625
cc_41 VPB N_A_27_508#_c_110_n 0.0179496f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_42 VPB N_A_27_508#_c_111_n 0.0115444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_27_508#_c_112_n 0.00964557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_27_508#_c_105_n 0.0133945f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=0.925
cc_45 VPB N_A_27_508#_c_108_n 0.0125837f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=2.035
cc_46 VPB N_A1_M1006_g 0.0198705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A2_M1003_g 0.0255526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_232_n 0.00984292f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=0.955
cc_49 VPB N_VPWR_c_233_n 0.00557173f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.105
cc_50 VPB N_VPWR_c_234_n 0.0169178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_235_n 0.0303033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_236_n 0.0177367f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=0.925
cc_53 VPB N_VPWR_c_231_n 0.0554183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_238_n 0.00613202f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.295
cc_55 VPB N_VPWR_c_239_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB Y 0.00385899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_302_367#_c_301_n 0.0142364f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.105
cc_58 VPB N_A_302_367#_c_302_n 0.00669813f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_59 VPB N_A_302_367#_c_303_n 0.0470363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_B1_N_M1002_g N_A_27_508#_M1004_g 0.0171745f $X=0.805 $Y=0.445 $X2=0
+ $Y2=0
cc_61 N_B1_N_M1001_g N_A_27_508#_c_110_n 0.00313661f $X=0.475 $Y=2.75 $X2=0
+ $Y2=0
cc_62 N_B1_N_M1001_g N_A_27_508#_c_111_n 0.0188648f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_63 N_B1_N_c_69_n N_A_27_508#_c_111_n 0.0017256f $X=0.475 $Y=1.99 $X2=0 $Y2=0
cc_64 N_B1_N_c_64_n N_A_27_508#_c_112_n 5.17635e-19 $X=0.27 $Y=1.625 $X2=0 $Y2=0
cc_65 N_B1_N_c_69_n N_A_27_508#_c_112_n 4.48587e-19 $X=0.475 $Y=1.99 $X2=0 $Y2=0
cc_66 B1_N N_A_27_508#_c_112_n 0.0240856f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_B1_N_c_61_n N_A_27_508#_c_104_n 3.75606e-19 $X=0.73 $Y=1.03 $X2=0 $Y2=0
cc_68 N_B1_N_c_64_n N_A_27_508#_c_104_n 0.00409084f $X=0.27 $Y=1.625 $X2=0 $Y2=0
cc_69 N_B1_N_c_60_n N_A_27_508#_c_105_n 0.00409084f $X=0.36 $Y=1.915 $X2=0 $Y2=0
cc_70 N_B1_N_c_69_n N_A_27_508#_c_105_n 0.0117618f $X=0.475 $Y=1.99 $X2=0 $Y2=0
cc_71 N_B1_N_c_61_n N_A_27_508#_c_106_n 2.12993e-19 $X=0.73 $Y=1.03 $X2=0 $Y2=0
cc_72 N_B1_N_c_62_n N_A_27_508#_c_106_n 0.00731346f $X=0.435 $Y=1.03 $X2=0 $Y2=0
cc_73 N_B1_N_M1002_g N_A_27_508#_c_106_n 0.00628184f $X=0.805 $Y=0.445 $X2=0
+ $Y2=0
cc_74 N_B1_N_c_61_n N_A_27_508#_c_107_n 0.00996575f $X=0.73 $Y=1.03 $X2=0 $Y2=0
cc_75 N_B1_N_M1002_g N_A_27_508#_c_107_n 0.0107377f $X=0.805 $Y=0.445 $X2=0
+ $Y2=0
cc_76 B1_N N_A_27_508#_c_107_n 0.066005f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_77 N_B1_N_c_66_n N_A_27_508#_c_107_n 0.00409084f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_78 N_B1_N_c_61_n N_A_27_508#_c_108_n 0.0113482f $X=0.73 $Y=1.03 $X2=0 $Y2=0
cc_79 B1_N N_A_27_508#_c_108_n 3.66534e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_B1_N_c_66_n N_A_27_508#_c_108_n 0.0174071f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_81 N_B1_N_M1001_g N_VPWR_c_232_n 0.0138465f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_82 N_B1_N_M1001_g N_VPWR_c_234_n 0.00383152f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_83 N_B1_N_M1001_g N_VPWR_c_231_n 0.00391732f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_84 N_B1_N_M1001_g Y 0.00537834f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_85 N_B1_N_M1002_g N_VGND_c_326_n 0.00941511f $X=0.805 $Y=0.445 $X2=0 $Y2=0
cc_86 N_B1_N_M1002_g N_VGND_c_329_n 0.00437168f $X=0.805 $Y=0.445 $X2=0 $Y2=0
cc_87 N_B1_N_M1002_g N_VGND_c_332_n 0.00892506f $X=0.805 $Y=0.445 $X2=0 $Y2=0
cc_88 B1_N N_VGND_c_332_n 0.0110936f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A_27_508#_M1000_g N_A1_M1006_g 0.0262982f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_27_508#_M1004_g A1 2.26892e-19 $X=1.33 $Y=0.655 $X2=0 $Y2=0
cc_91 N_A_27_508#_c_103_n N_A1_c_174_n 0.00886879f $X=1.435 $Y=1.42 $X2=0 $Y2=0
cc_92 N_A_27_508#_M1004_g N_A1_c_175_n 0.0160488f $X=1.33 $Y=0.655 $X2=0 $Y2=0
cc_93 N_A_27_508#_M1000_g N_VPWR_c_232_n 0.00308716f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_A_27_508#_c_111_n N_VPWR_c_232_n 0.0255154f $X=0.66 $Y=2.385 $X2=0 $Y2=0
cc_95 N_A_27_508#_c_110_n N_VPWR_c_234_n 0.00864257f $X=0.26 $Y=2.75 $X2=0 $Y2=0
cc_96 N_A_27_508#_M1000_g N_VPWR_c_235_n 0.00585385f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_97 N_A_27_508#_M1000_g N_VPWR_c_231_n 0.0120903f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_98 N_A_27_508#_c_110_n N_VPWR_c_231_n 0.00911154f $X=0.26 $Y=2.75 $X2=0 $Y2=0
cc_99 N_A_27_508#_c_111_n N_VPWR_c_231_n 0.00873716f $X=0.66 $Y=2.385 $X2=0
+ $Y2=0
cc_100 N_A_27_508#_c_100_n N_Y_c_268_n 0.0093004f $X=1.255 $Y=1.42 $X2=0 $Y2=0
cc_101 N_A_27_508#_M1004_g N_Y_c_268_n 0.0127868f $X=1.33 $Y=0.655 $X2=0 $Y2=0
cc_102 N_A_27_508#_M1000_g N_Y_c_268_n 0.00767473f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_27_508#_c_103_n N_Y_c_268_n 0.00784914f $X=1.435 $Y=1.42 $X2=0 $Y2=0
cc_104 N_A_27_508#_c_104_n N_Y_c_268_n 0.0131288f $X=0.792 $Y=1.477 $X2=0 $Y2=0
cc_105 N_A_27_508#_c_107_n N_Y_c_268_n 0.00814406f $X=0.792 $Y=1.345 $X2=0 $Y2=0
cc_106 N_A_27_508#_M1004_g N_Y_c_269_n 0.00268096f $X=1.33 $Y=0.655 $X2=0 $Y2=0
cc_107 N_A_27_508#_c_103_n N_Y_c_269_n 5.15345e-19 $X=1.435 $Y=1.42 $X2=0 $Y2=0
cc_108 N_A_27_508#_c_107_n N_Y_c_269_n 0.00468901f $X=0.792 $Y=1.345 $X2=0 $Y2=0
cc_109 N_A_27_508#_c_100_n Y 0.00366664f $X=1.255 $Y=1.42 $X2=0 $Y2=0
cc_110 N_A_27_508#_M1000_g Y 0.0115925f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_27_508#_c_111_n Y 0.0145391f $X=0.66 $Y=2.385 $X2=0 $Y2=0
cc_112 N_A_27_508#_c_105_n Y 0.0617794f $X=0.84 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A_27_508#_c_108_n Y 0.0013781f $X=0.84 $Y=1.42 $X2=0 $Y2=0
cc_114 N_A_27_508#_M1000_g N_A_302_367#_c_302_n 0.00131456f $X=1.435 $Y=2.465
+ $X2=0 $Y2=0
cc_115 N_A_27_508#_c_100_n N_VGND_c_326_n 7.52731e-19 $X=1.255 $Y=1.42 $X2=0
+ $Y2=0
cc_116 N_A_27_508#_M1004_g N_VGND_c_326_n 0.00385352f $X=1.33 $Y=0.655 $X2=0
+ $Y2=0
cc_117 N_A_27_508#_c_106_n N_VGND_c_326_n 0.0254058f $X=0.745 $Y=0.445 $X2=0
+ $Y2=0
cc_118 N_A_27_508#_c_107_n N_VGND_c_326_n 0.0310328f $X=0.792 $Y=1.345 $X2=0
+ $Y2=0
cc_119 N_A_27_508#_c_108_n N_VGND_c_326_n 0.00334216f $X=0.84 $Y=1.42 $X2=0
+ $Y2=0
cc_120 N_A_27_508#_c_106_n N_VGND_c_329_n 0.0214926f $X=0.745 $Y=0.445 $X2=0
+ $Y2=0
cc_121 N_A_27_508#_M1004_g N_VGND_c_330_n 0.00585385f $X=1.33 $Y=0.655 $X2=0
+ $Y2=0
cc_122 N_A_27_508#_M1002_s N_VGND_c_332_n 0.0021695f $X=0.465 $Y=0.235 $X2=0
+ $Y2=0
cc_123 N_A_27_508#_M1004_g N_VGND_c_332_n 0.0109339f $X=1.33 $Y=0.655 $X2=0
+ $Y2=0
cc_124 N_A_27_508#_c_106_n N_VGND_c_332_n 0.0147683f $X=0.745 $Y=0.445 $X2=0
+ $Y2=0
cc_125 N_A1_M1006_g N_A2_M1003_g 0.0192685f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_126 A1 A2 0.0268329f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A1_c_174_n A2 2.59523e-19 $X=1.915 $Y=1.35 $X2=0 $Y2=0
cc_128 N_A1_c_174_n N_A2_c_210_n 0.0172458f $X=1.915 $Y=1.35 $X2=0 $Y2=0
cc_129 A1 N_A2_c_211_n 0.00762913f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A1_c_175_n N_A2_c_211_n 0.0258804f $X=1.915 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A1_M1006_g N_VPWR_c_233_n 0.00355081f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A1_M1006_g N_VPWR_c_235_n 0.00571722f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A1_M1006_g N_VPWR_c_231_n 0.0105533f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_134 A1 N_Y_c_268_n 0.0256129f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A1_c_174_n N_Y_c_268_n 0.00247551f $X=1.915 $Y=1.35 $X2=0 $Y2=0
cc_136 A1 N_Y_c_269_n 0.0648855f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_137 N_A1_c_175_n N_Y_c_269_n 0.00603145f $X=1.915 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A1_M1006_g N_A_302_367#_c_305_n 0.0144753f $X=1.865 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A1_M1006_g N_A_302_367#_c_301_n 0.0136428f $X=1.865 $Y=2.465 $X2=0
+ $Y2=0
cc_140 A1 N_A_302_367#_c_301_n 4.01007e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_141 A1 N_A_302_367#_c_301_n 0.0341874f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A1_c_174_n N_A_302_367#_c_301_n 9.86927e-19 $X=1.915 $Y=1.35 $X2=0
+ $Y2=0
cc_143 N_A1_M1006_g N_A_302_367#_c_302_n 0.00214002f $X=1.865 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A1_c_174_n N_A_302_367#_c_302_n 0.00193542f $X=1.915 $Y=1.35 $X2=0
+ $Y2=0
cc_145 N_A1_c_175_n N_VGND_c_328_n 0.00190847f $X=1.915 $Y=1.185 $X2=0 $Y2=0
cc_146 A1 N_VGND_c_330_n 0.016074f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_147 N_A1_c_175_n N_VGND_c_330_n 0.00491601f $X=1.915 $Y=1.185 $X2=0 $Y2=0
cc_148 A1 N_VGND_c_332_n 0.0157749f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_149 N_A1_c_175_n N_VGND_c_332_n 0.00887979f $X=1.915 $Y=1.185 $X2=0 $Y2=0
cc_150 A1 A_380_47# 0.0103593f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_151 A1 A_380_47# 7.25904e-19 $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_152 N_A2_M1003_g N_VPWR_c_233_n 0.00362135f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A2_M1003_g N_VPWR_c_236_n 0.00585385f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A2_M1003_g N_VPWR_c_231_n 0.0117391f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A2_M1003_g N_A_302_367#_c_305_n 4.84681e-19 $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A2_M1003_g N_A_302_367#_c_301_n 0.0196654f $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_157 A2 N_A_302_367#_c_301_n 0.0293142f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A2_c_210_n N_A_302_367#_c_301_n 0.00477561f $X=2.51 $Y=1.35 $X2=0 $Y2=0
cc_159 A2 N_VGND_c_328_n 0.024896f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_c_210_n N_VGND_c_328_n 0.00460192f $X=2.51 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A2_c_211_n N_VGND_c_328_n 0.018882f $X=2.497 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A2_c_211_n N_VGND_c_330_n 0.00486043f $X=2.497 $Y=1.185 $X2=0 $Y2=0
cc_163 N_A2_c_211_n N_VGND_c_332_n 0.00870566f $X=2.497 $Y=1.185 $X2=0 $Y2=0
cc_164 N_VPWR_c_231_n N_Y_M1000_s 0.00231748f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_c_232_n Y 0.0272929f $X=0.69 $Y=2.765 $X2=0 $Y2=0
cc_166 N_VPWR_c_235_n Y 0.0163642f $X=1.97 $Y=3.33 $X2=0 $Y2=0
cc_167 N_VPWR_c_231_n Y 0.0100304f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_231_n N_A_302_367#_M1000_d 0.0027574f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_169 N_VPWR_c_231_n N_A_302_367#_M1003_d 0.00215158f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_235_n N_A_302_367#_c_305_n 0.0157299f $X=1.97 $Y=3.33 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_231_n N_A_302_367#_c_305_n 0.0104992f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_172 N_VPWR_M1006_d N_A_302_367#_c_301_n 0.00284866f $X=1.94 $Y=1.835 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_233_n N_A_302_367#_c_301_n 0.0216414f $X=2.135 $Y=2.11 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_236_n N_A_302_367#_c_303_n 0.0194077f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_231_n N_A_302_367#_c_303_n 0.0117799f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_Y_c_268_n N_A_302_367#_c_302_n 0.0118754f $X=1.537 $Y=1.21 $X2=0 $Y2=0
cc_177 Y N_A_302_367#_c_302_n 0.0129504f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_178 N_Y_c_268_n N_VGND_c_326_n 0.0107785f $X=1.537 $Y=1.21 $X2=0 $Y2=0
cc_179 N_Y_c_269_n N_VGND_c_330_n 0.0154837f $X=1.575 $Y=0.42 $X2=0 $Y2=0
cc_180 N_Y_M1004_d N_VGND_c_332_n 0.00623705f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_181 N_Y_c_269_n N_VGND_c_332_n 0.00944728f $X=1.575 $Y=0.42 $X2=0 $Y2=0
cc_182 N_VGND_c_332_n A_380_47# 0.00518631f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
