* File: sky130_fd_sc_lp__o41ai_2.pxi.spice
* Created: Wed Sep  2 10:28:20 2020
* 
x_PM_SKY130_FD_SC_LP__O41AI_2%B1 N_B1_M1009_g N_B1_M1018_g N_B1_c_96_n
+ N_B1_M1007_g N_B1_c_97_n N_B1_M1008_g B1 B1 N_B1_c_98_n
+ PM_SKY130_FD_SC_LP__O41AI_2%B1
x_PM_SKY130_FD_SC_LP__O41AI_2%A4 N_A4_M1002_g N_A4_M1015_g N_A4_M1011_g
+ N_A4_M1016_g A4 A4 N_A4_c_141_n PM_SKY130_FD_SC_LP__O41AI_2%A4
x_PM_SKY130_FD_SC_LP__O41AI_2%A3 N_A3_M1001_g N_A3_M1013_g N_A3_M1019_g
+ N_A3_M1014_g A3 N_A3_c_199_n N_A3_c_200_n PM_SKY130_FD_SC_LP__O41AI_2%A3
x_PM_SKY130_FD_SC_LP__O41AI_2%A2 N_A2_M1003_g N_A2_M1012_g N_A2_c_255_n
+ N_A2_M1000_g N_A2_c_252_n N_A2_c_253_n N_A2_c_258_n N_A2_M1006_g A2 A2 A2
+ PM_SKY130_FD_SC_LP__O41AI_2%A2
x_PM_SKY130_FD_SC_LP__O41AI_2%A1 N_A1_c_304_n N_A1_M1005_g N_A1_c_305_n
+ N_A1_c_306_n N_A1_c_307_n N_A1_M1017_g N_A1_M1004_g N_A1_M1010_g A1 A1
+ N_A1_c_311_n PM_SKY130_FD_SC_LP__O41AI_2%A1
x_PM_SKY130_FD_SC_LP__O41AI_2%VPWR N_VPWR_M1009_d N_VPWR_M1018_d N_VPWR_M1004_s
+ N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n N_VPWR_c_350_n VPWR
+ N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_346_n N_VPWR_c_355_n
+ N_VPWR_c_356_n PM_SKY130_FD_SC_LP__O41AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O41AI_2%Y N_Y_M1007_d N_Y_M1009_s N_Y_M1002_s N_Y_c_448_n
+ N_Y_c_421_n N_Y_c_419_n N_Y_c_437_n Y Y N_Y_c_423_n
+ PM_SKY130_FD_SC_LP__O41AI_2%Y
x_PM_SKY130_FD_SC_LP__O41AI_2%A_313_365# N_A_313_365#_M1002_d
+ N_A_313_365#_M1011_d N_A_313_365#_M1019_d N_A_313_365#_c_466_n
+ N_A_313_365#_c_467_n N_A_313_365#_c_472_n N_A_313_365#_c_474_n
+ N_A_313_365#_c_477_n N_A_313_365#_c_478_n N_A_313_365#_c_468_n
+ N_A_313_365#_c_469_n PM_SKY130_FD_SC_LP__O41AI_2%A_313_365#
x_PM_SKY130_FD_SC_LP__O41AI_2%A_615_365# N_A_615_365#_M1013_s
+ N_A_615_365#_M1000_s N_A_615_365#_c_512_n N_A_615_365#_c_511_n
+ N_A_615_365#_c_515_n N_A_615_365#_c_519_n
+ PM_SKY130_FD_SC_LP__O41AI_2%A_615_365#
x_PM_SKY130_FD_SC_LP__O41AI_2%A_808_367# N_A_808_367#_M1000_d
+ N_A_808_367#_M1006_d N_A_808_367#_M1010_d N_A_808_367#_c_538_n
+ N_A_808_367#_c_539_n N_A_808_367#_c_544_n N_A_808_367#_c_558_n
+ N_A_808_367#_c_549_n N_A_808_367#_c_540_n N_A_808_367#_c_541_n
+ N_A_808_367#_c_548_n PM_SKY130_FD_SC_LP__O41AI_2%A_808_367#
x_PM_SKY130_FD_SC_LP__O41AI_2%A_155_47# N_A_155_47#_M1007_s N_A_155_47#_M1008_s
+ N_A_155_47#_M1016_s N_A_155_47#_M1014_s N_A_155_47#_M1012_s
+ N_A_155_47#_M1017_d N_A_155_47#_c_581_n N_A_155_47#_c_587_n
+ N_A_155_47#_c_588_n N_A_155_47#_c_570_n N_A_155_47#_c_571_n
+ N_A_155_47#_c_596_n N_A_155_47#_c_572_n N_A_155_47#_c_639_p
+ N_A_155_47#_c_573_n N_A_155_47#_c_640_p N_A_155_47#_c_574_n
+ N_A_155_47#_c_575_n N_A_155_47#_c_576_n N_A_155_47#_c_577_n
+ N_A_155_47#_c_578_n N_A_155_47#_c_579_n PM_SKY130_FD_SC_LP__O41AI_2%A_155_47#
x_PM_SKY130_FD_SC_LP__O41AI_2%VGND N_VGND_M1015_d N_VGND_M1001_d N_VGND_M1003_d
+ N_VGND_M1005_s N_VGND_c_655_n N_VGND_c_656_n N_VGND_c_657_n N_VGND_c_658_n
+ N_VGND_c_659_n VGND N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n
+ N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ N_VGND_c_668_n PM_SKY130_FD_SC_LP__O41AI_2%VGND
cc_1 VNB N_B1_M1009_g 0.00394253f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_2 VNB N_B1_M1018_g 0.00275124f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.465
cc_3 VNB N_B1_c_96_n 0.166671f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.185
cc_4 VNB N_B1_c_97_n 0.0159413f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=1.185
cc_5 VNB N_B1_c_98_n 0.0329852f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.44
cc_6 VNB N_A4_M1015_g 0.0256685f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.465
cc_7 VNB N_A4_M1016_g 0.0256813f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB A4 0.00195572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A4_c_141_n 0.0465226f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=1.27
cc_10 VNB N_A3_M1001_g 0.0241035f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_11 VNB N_A3_M1014_g 0.0243113f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_A3_c_199_n 0.03549f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.27
cc_13 VNB N_A3_c_200_n 0.00362479f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.27
cc_14 VNB N_A2_M1003_g 0.0236281f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_15 VNB N_A2_M1012_g 0.0237278f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.465
cc_16 VNB N_A2_c_252_n 0.0138857f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=1.185
cc_17 VNB N_A2_c_253_n 0.0345532f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=0.655
cc_18 VNB A2 0.01143f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.27
cc_19 VNB N_A1_c_304_n 0.0153131f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.605
cc_20 VNB N_A1_c_305_n 0.0128798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_306_n 0.0081134f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.605
cc_22 VNB N_A1_c_307_n 0.0198106f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.465
cc_23 VNB N_A1_M1004_g 0.00357919f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.655
cc_24 VNB N_A1_M1010_g 0.00399138f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB A1 0.0134036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A1_c_311_n 0.111368f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.27
cc_27 VNB N_VPWR_c_346_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_419_n 6.33024e-19 $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.1
cc_29 VNB Y 0.00360516f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.27
cc_30 VNB N_A_155_47#_c_570_n 0.00518945f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.44
cc_31 VNB N_A_155_47#_c_571_n 0.00276554f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.27
cc_32 VNB N_A_155_47#_c_572_n 0.00476487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_155_47#_c_573_n 0.00406958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_155_47#_c_574_n 0.0119533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_155_47#_c_575_n 0.0282223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_155_47#_c_576_n 0.0239774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_155_47#_c_577_n 0.00216703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_155_47#_c_578_n 0.00323033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_155_47#_c_579_n 0.00132773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_655_n 0.00504245f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_41 VNB N_VGND_c_656_n 0.0165128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_657_n 0.00222241f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.1
cc_43 VNB N_VGND_c_658_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.44
cc_44 VNB N_VGND_c_659_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.27
cc_45 VNB N_VGND_c_660_n 0.0573907f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.27
cc_46 VNB N_VGND_c_661_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_662_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_663_n 0.032943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_664_n 0.357174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_665_n 0.00634562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_666_n 0.00525267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_667_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_668_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VPB N_B1_M1009_g 0.0272332f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_55 VPB N_B1_M1018_g 0.0226885f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_56 VPB N_A4_M1002_g 0.0224494f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_57 VPB N_A4_M1011_g 0.0205011f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.655
cc_58 VPB A4 0.00834398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A4_c_141_n 0.0154185f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.27
cc_60 VPB N_A3_M1013_g 0.0207829f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_61 VPB N_A3_M1019_g 0.023738f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.655
cc_62 VPB N_A3_c_199_n 0.012919f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.27
cc_63 VPB N_A3_c_200_n 0.00301075f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.27
cc_64 VPB N_A2_c_255_n 0.021561f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.185
cc_65 VPB N_A2_c_252_n 0.00697467f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.185
cc_66 VPB N_A2_c_253_n 0.0216976f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=0.655
cc_67 VPB N_A2_c_258_n 0.0162141f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=0.655
cc_68 VPB A2 0.0115649f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.27
cc_69 VPB N_A1_M1004_g 0.0199119f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.655
cc_70 VPB N_A1_M1010_g 0.0254689f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_71 VPB A1 0.0122785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_347_n 0.0125708f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.655
cc_73 VPB N_VPWR_c_348_n 0.0571186f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.185
cc_74 VPB N_VPWR_c_349_n 0.0125151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_350_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.44
cc_76 VPB N_VPWR_c_351_n 0.0146078f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.27
cc_77 VPB N_VPWR_c_352_n 0.0937402f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.27
cc_78 VPB N_VPWR_c_353_n 0.018399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_346_n 0.0616014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_355_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_356_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_Y_c_421_n 0.00345305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB Y 0.0100379f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.27
cc_84 VPB N_Y_c_423_n 0.00222393f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.27
cc_85 VPB N_A_313_365#_c_466_n 0.00191946f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.655
cc_86 VPB N_A_313_365#_c_467_n 0.00783226f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.185
cc_87 VPB N_A_313_365#_c_468_n 0.0031496f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.27
cc_88 VPB N_A_313_365#_c_469_n 0.00605419f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.44
cc_89 VPB N_A_615_365#_c_511_n 0.0109112f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.655
cc_90 VPB N_A_808_367#_c_538_n 0.00176898f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.655
cc_91 VPB N_A_808_367#_c_539_n 0.00605419f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.185
cc_92 VPB N_A_808_367#_c_540_n 0.00744325f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.27
cc_93 VPB N_A_808_367#_c_541_n 0.0373194f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.44
cc_94 N_B1_c_97_n N_A4_M1015_g 0.023674f $X=1.545 $Y=1.185 $X2=0 $Y2=0
cc_95 N_B1_c_96_n N_A4_c_141_n 0.0176787f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_96 N_B1_M1009_g N_VPWR_c_348_n 0.00773581f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B1_c_96_n N_VPWR_c_348_n 0.00298442f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_98 N_B1_c_98_n N_VPWR_c_348_n 0.0176849f $X=0.9 $Y=1.44 $X2=0 $Y2=0
cc_99 N_B1_M1009_g N_VPWR_c_349_n 7.53524e-19 $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B1_M1018_g N_VPWR_c_349_n 0.0166682f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B1_c_96_n N_VPWR_c_349_n 4.30846e-19 $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_102 N_B1_M1009_g N_VPWR_c_351_n 0.00585385f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_103 N_B1_M1018_g N_VPWR_c_351_n 0.00486043f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_104 N_B1_M1009_g N_VPWR_c_346_n 0.0114853f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_105 N_B1_M1018_g N_VPWR_c_346_n 0.00824727f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_106 N_B1_M1009_g N_Y_c_421_n 0.00382917f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_107 N_B1_c_96_n N_Y_c_421_n 0.00287509f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_108 N_B1_c_98_n N_Y_c_421_n 0.0183183f $X=0.9 $Y=1.44 $X2=0 $Y2=0
cc_109 N_B1_c_96_n N_Y_c_419_n 0.0123743f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_110 N_B1_c_97_n N_Y_c_419_n 0.00801196f $X=1.545 $Y=1.185 $X2=0 $Y2=0
cc_111 N_B1_c_98_n N_Y_c_419_n 0.0231815f $X=0.9 $Y=1.44 $X2=0 $Y2=0
cc_112 N_B1_M1018_g Y 0.00394238f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B1_c_96_n Y 0.0343554f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_114 N_B1_c_98_n Y 0.0159144f $X=0.9 $Y=1.44 $X2=0 $Y2=0
cc_115 N_B1_M1018_g N_Y_c_423_n 0.0156437f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B1_c_96_n N_Y_c_423_n 0.00860101f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_117 N_B1_c_98_n N_Y_c_423_n 0.0165228f $X=0.9 $Y=1.44 $X2=0 $Y2=0
cc_118 N_B1_M1018_g N_A_313_365#_c_467_n 0.00134386f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_B1_c_96_n N_A_313_365#_c_467_n 4.07348e-19 $X=1.115 $Y=1.185 $X2=0
+ $Y2=0
cc_120 N_B1_c_98_n N_A_155_47#_M1007_s 0.002287f $X=0.9 $Y=1.44 $X2=-0.19
+ $Y2=-0.245
cc_121 N_B1_c_96_n N_A_155_47#_c_581_n 0.0105205f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_122 N_B1_c_97_n N_A_155_47#_c_581_n 0.0118089f $X=1.545 $Y=1.185 $X2=0 $Y2=0
cc_123 N_B1_c_97_n N_A_155_47#_c_571_n 7.54217e-19 $X=1.545 $Y=1.185 $X2=0 $Y2=0
cc_124 N_B1_c_96_n N_A_155_47#_c_576_n 0.00755406f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_125 N_B1_c_97_n N_A_155_47#_c_576_n 4.47146e-19 $X=1.545 $Y=1.185 $X2=0 $Y2=0
cc_126 N_B1_c_98_n N_A_155_47#_c_576_n 0.0235187f $X=0.9 $Y=1.44 $X2=0 $Y2=0
cc_127 N_B1_c_96_n N_VGND_c_660_n 0.00357842f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_128 N_B1_c_97_n N_VGND_c_660_n 0.00357877f $X=1.545 $Y=1.185 $X2=0 $Y2=0
cc_129 N_B1_c_96_n N_VGND_c_664_n 0.00665087f $X=1.115 $Y=1.185 $X2=0 $Y2=0
cc_130 N_B1_c_97_n N_VGND_c_664_n 0.00537654f $X=1.545 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A4_M1016_g N_A3_M1001_g 0.0239727f $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_132 N_A4_M1011_g N_A3_M1013_g 0.0256726f $X=2.335 $Y=2.455 $X2=0 $Y2=0
cc_133 A4 N_A3_M1013_g 0.00560484f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_134 A4 N_A3_M1019_g 5.6651e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_135 A4 N_A3_c_199_n 0.0221114f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A4_c_141_n N_A3_c_199_n 0.0215642f $X=2.57 $Y=1.5 $X2=0 $Y2=0
cc_137 A4 N_A3_c_200_n 0.0336602f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A4_M1002_g N_VPWR_c_349_n 0.00221807f $X=1.905 $Y=2.455 $X2=0 $Y2=0
cc_139 N_A4_M1002_g N_VPWR_c_352_n 0.00351226f $X=1.905 $Y=2.455 $X2=0 $Y2=0
cc_140 N_A4_M1011_g N_VPWR_c_352_n 0.00351226f $X=2.335 $Y=2.455 $X2=0 $Y2=0
cc_141 N_A4_M1002_g N_VPWR_c_346_n 0.00660267f $X=1.905 $Y=2.455 $X2=0 $Y2=0
cc_142 N_A4_M1011_g N_VPWR_c_346_n 0.00580191f $X=2.335 $Y=2.455 $X2=0 $Y2=0
cc_143 N_A4_M1015_g N_Y_c_419_n 0.00106275f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_144 N_A4_M1002_g N_Y_c_437_n 0.0149162f $X=1.905 $Y=2.455 $X2=0 $Y2=0
cc_145 N_A4_M1011_g N_Y_c_437_n 0.0107905f $X=2.335 $Y=2.455 $X2=0 $Y2=0
cc_146 N_A4_c_141_n N_Y_c_437_n 4.25969e-19 $X=2.57 $Y=1.5 $X2=0 $Y2=0
cc_147 N_A4_M1002_g Y 0.0162386f $X=1.905 $Y=2.455 $X2=0 $Y2=0
cc_148 N_A4_M1011_g Y 0.00579146f $X=2.335 $Y=2.455 $X2=0 $Y2=0
cc_149 A4 Y 0.0352957f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A4_c_141_n Y 0.0289135f $X=2.57 $Y=1.5 $X2=0 $Y2=0
cc_151 N_A4_M1002_g N_A_313_365#_c_472_n 0.011776f $X=1.905 $Y=2.455 $X2=0 $Y2=0
cc_152 N_A4_M1011_g N_A_313_365#_c_472_n 0.0147352f $X=2.335 $Y=2.455 $X2=0
+ $Y2=0
cc_153 N_A4_M1011_g N_A_313_365#_c_474_n 0.00186658f $X=2.335 $Y=2.455 $X2=0
+ $Y2=0
cc_154 A4 N_A_313_365#_c_474_n 0.0290942f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A4_c_141_n N_A_313_365#_c_474_n 0.00129777f $X=2.57 $Y=1.5 $X2=0 $Y2=0
cc_156 N_A4_M1011_g N_A_313_365#_c_477_n 0.0114482f $X=2.335 $Y=2.455 $X2=0
+ $Y2=0
cc_157 A4 N_A_313_365#_c_478_n 0.0246057f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A4_M1015_g N_A_155_47#_c_587_n 0.00199195f $X=1.975 $Y=0.655 $X2=0
+ $Y2=0
cc_159 N_A4_M1015_g N_A_155_47#_c_588_n 0.0087504f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_160 N_A4_M1016_g N_A_155_47#_c_588_n 8.42526e-19 $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A4_M1015_g N_A_155_47#_c_570_n 0.0119714f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A4_M1016_g N_A_155_47#_c_570_n 0.0119714f $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_163 A4 N_A_155_47#_c_570_n 0.0121205f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A4_c_141_n N_A_155_47#_c_570_n 0.00868481f $X=2.57 $Y=1.5 $X2=0 $Y2=0
cc_165 N_A4_M1015_g N_A_155_47#_c_571_n 0.00159668f $X=1.975 $Y=0.655 $X2=0
+ $Y2=0
cc_166 N_A4_c_141_n N_A_155_47#_c_571_n 0.00190679f $X=2.57 $Y=1.5 $X2=0 $Y2=0
cc_167 N_A4_M1015_g N_A_155_47#_c_596_n 8.841e-19 $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A4_M1016_g N_A_155_47#_c_596_n 0.0109782f $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_169 A4 N_A_155_47#_c_572_n 0.0236048f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A4_M1016_g N_A_155_47#_c_577_n 0.00179341f $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_171 A4 N_A_155_47#_c_577_n 0.0246648f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A4_c_141_n N_A_155_47#_c_577_n 0.0016307f $X=2.57 $Y=1.5 $X2=0 $Y2=0
cc_173 N_A4_M1015_g N_VGND_c_655_n 0.00687992f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A4_M1016_g N_VGND_c_655_n 0.00745117f $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_175 N_A4_M1016_g N_VGND_c_656_n 0.0054895f $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_176 N_A4_M1016_g N_VGND_c_657_n 6.74436e-19 $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A4_M1015_g N_VGND_c_660_n 0.00547432f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A4_M1015_g N_VGND_c_664_n 0.0102728f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A4_M1016_g N_VGND_c_664_n 0.0103509f $X=2.57 $Y=0.655 $X2=0 $Y2=0
cc_180 N_A3_M1014_g N_A2_M1003_g 0.0233922f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_181 N_A3_c_199_n N_A2_M1003_g 0.0213744f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_182 N_A3_c_200_n N_A2_M1003_g 0.00301323f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_183 N_A3_M1019_g N_A2_c_253_n 0.00203626f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_184 N_A3_c_199_n A2 2.77318e-19 $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_185 N_A3_c_200_n A2 0.0350573f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_186 N_A3_M1013_g N_VPWR_c_352_n 0.00537804f $X=3 $Y=2.455 $X2=0 $Y2=0
cc_187 N_A3_M1019_g N_VPWR_c_352_n 0.00351191f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_188 N_A3_M1013_g N_VPWR_c_346_n 0.0104252f $X=3 $Y=2.455 $X2=0 $Y2=0
cc_189 N_A3_M1019_g N_VPWR_c_346_n 0.00660265f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_190 N_A3_M1013_g N_Y_c_437_n 4.40564e-19 $X=3 $Y=2.455 $X2=0 $Y2=0
cc_191 N_A3_M1013_g Y 5.37592e-19 $X=3 $Y=2.455 $X2=0 $Y2=0
cc_192 N_A3_M1013_g N_A_313_365#_c_472_n 0.0019819f $X=3 $Y=2.455 $X2=0 $Y2=0
cc_193 N_A3_M1013_g N_A_313_365#_c_477_n 0.0114074f $X=3 $Y=2.455 $X2=0 $Y2=0
cc_194 N_A3_M1013_g N_A_313_365#_c_478_n 0.0150738f $X=3 $Y=2.455 $X2=0 $Y2=0
cc_195 N_A3_M1019_g N_A_313_365#_c_478_n 0.0132014f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_196 N_A3_c_199_n N_A_313_365#_c_478_n 0.00359459f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_197 N_A3_c_200_n N_A_313_365#_c_478_n 0.0106171f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_198 N_A3_c_199_n N_A_313_365#_c_468_n 5.09104e-19 $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_199 N_A3_c_200_n N_A_313_365#_c_468_n 0.0179716f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_200 N_A3_M1013_g N_A_615_365#_c_512_n 0.00940873f $X=3 $Y=2.455 $X2=0 $Y2=0
cc_201 N_A3_M1019_g N_A_615_365#_c_512_n 0.0144635f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_202 N_A3_M1019_g N_A_615_365#_c_511_n 0.0125325f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_203 N_A3_M1013_g N_A_615_365#_c_515_n 0.00213152f $X=3 $Y=2.455 $X2=0 $Y2=0
cc_204 N_A3_M1019_g N_A_615_365#_c_515_n 5.84237e-19 $X=3.43 $Y=2.455 $X2=0
+ $Y2=0
cc_205 N_A3_M1001_g N_A_155_47#_c_572_n 0.014152f $X=3 $Y=0.655 $X2=0 $Y2=0
cc_206 N_A3_M1014_g N_A_155_47#_c_572_n 0.0143775f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_207 N_A3_c_199_n N_A_155_47#_c_572_n 0.00526658f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_208 N_A3_c_200_n N_A_155_47#_c_572_n 0.013545f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_209 N_A3_c_199_n N_A_155_47#_c_578_n 5.14458e-19 $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_210 N_A3_c_200_n N_A_155_47#_c_578_n 0.0167987f $X=3.47 $Y=1.5 $X2=0 $Y2=0
cc_211 N_A3_M1001_g N_VGND_c_656_n 0.00564095f $X=3 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A3_M1001_g N_VGND_c_657_n 0.00856384f $X=3 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A3_M1014_g N_VGND_c_657_n 0.00169872f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A3_M1014_g N_VGND_c_658_n 6.27404e-19 $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_215 N_A3_M1014_g N_VGND_c_661_n 0.00585385f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_216 N_A3_M1001_g N_VGND_c_664_n 0.00950825f $X=3 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A3_M1014_g N_VGND_c_664_n 0.0107095f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A2_M1012_g N_A1_c_304_n 0.0244183f $X=4.35 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A2_c_252_n N_A1_c_306_n 0.00986734f $X=4.735 $Y=1.65 $X2=0 $Y2=0
cc_220 A2 N_A1_c_306_n 0.00957467f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_221 N_A2_c_258_n N_A1_M1004_g 0.01114f $X=4.81 $Y=1.725 $X2=0 $Y2=0
cc_222 A2 A1 0.0375512f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_223 N_A2_c_252_n N_A1_c_311_n 0.01114f $X=4.735 $Y=1.65 $X2=0 $Y2=0
cc_224 A2 N_A1_c_311_n 0.00939155f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_225 N_A2_c_258_n N_VPWR_c_350_n 0.00132281f $X=4.81 $Y=1.725 $X2=0 $Y2=0
cc_226 N_A2_c_255_n N_VPWR_c_352_n 0.00357842f $X=4.38 $Y=1.725 $X2=0 $Y2=0
cc_227 N_A2_c_258_n N_VPWR_c_352_n 0.00547432f $X=4.81 $Y=1.725 $X2=0 $Y2=0
cc_228 N_A2_c_255_n N_VPWR_c_346_n 0.00675085f $X=4.38 $Y=1.725 $X2=0 $Y2=0
cc_229 N_A2_c_258_n N_VPWR_c_346_n 0.00990114f $X=4.81 $Y=1.725 $X2=0 $Y2=0
cc_230 N_A2_c_255_n N_A_615_365#_c_511_n 0.0131508f $X=4.38 $Y=1.725 $X2=0 $Y2=0
cc_231 N_A2_c_258_n N_A_615_365#_c_511_n 0.00193114f $X=4.81 $Y=1.725 $X2=0
+ $Y2=0
cc_232 N_A2_c_255_n N_A_615_365#_c_519_n 0.0144635f $X=4.38 $Y=1.725 $X2=0 $Y2=0
cc_233 N_A2_c_258_n N_A_615_365#_c_519_n 0.00858643f $X=4.81 $Y=1.725 $X2=0
+ $Y2=0
cc_234 N_A2_c_253_n N_A_808_367#_c_538_n 0.00187379f $X=4.455 $Y=1.65 $X2=0
+ $Y2=0
cc_235 A2 N_A_808_367#_c_538_n 0.0224541f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_236 N_A2_c_255_n N_A_808_367#_c_544_n 0.0122595f $X=4.38 $Y=1.725 $X2=0 $Y2=0
cc_237 N_A2_c_252_n N_A_808_367#_c_544_n 6.66393e-19 $X=4.735 $Y=1.65 $X2=0
+ $Y2=0
cc_238 N_A2_c_258_n N_A_808_367#_c_544_n 0.0121892f $X=4.81 $Y=1.725 $X2=0 $Y2=0
cc_239 A2 N_A_808_367#_c_544_n 0.0437342f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_240 A2 N_A_808_367#_c_548_n 0.0156741f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_241 N_A2_M1003_g N_A_155_47#_c_573_n 0.0157317f $X=3.92 $Y=0.655 $X2=0 $Y2=0
cc_242 N_A2_M1012_g N_A_155_47#_c_573_n 0.0133082f $X=4.35 $Y=0.655 $X2=0 $Y2=0
cc_243 N_A2_c_253_n N_A_155_47#_c_573_n 8.61545e-19 $X=4.455 $Y=1.65 $X2=0 $Y2=0
cc_244 A2 N_A_155_47#_c_573_n 0.0418472f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A2_c_252_n N_A_155_47#_c_574_n 3.31476e-19 $X=4.735 $Y=1.65 $X2=0 $Y2=0
cc_246 A2 N_A_155_47#_c_574_n 0.0388938f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A2_c_252_n N_A_155_47#_c_579_n 8.80911e-19 $X=4.735 $Y=1.65 $X2=0 $Y2=0
cc_248 A2 N_A_155_47#_c_579_n 0.0170873f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_249 N_A2_M1003_g N_VGND_c_658_n 0.0101678f $X=3.92 $Y=0.655 $X2=0 $Y2=0
cc_250 N_A2_M1012_g N_VGND_c_658_n 0.010076f $X=4.35 $Y=0.655 $X2=0 $Y2=0
cc_251 N_A2_M1012_g N_VGND_c_659_n 6.11179e-19 $X=4.35 $Y=0.655 $X2=0 $Y2=0
cc_252 N_A2_M1003_g N_VGND_c_661_n 0.00486043f $X=3.92 $Y=0.655 $X2=0 $Y2=0
cc_253 N_A2_M1012_g N_VGND_c_662_n 0.00486043f $X=4.35 $Y=0.655 $X2=0 $Y2=0
cc_254 N_A2_M1003_g N_VGND_c_664_n 0.0082726f $X=3.92 $Y=0.655 $X2=0 $Y2=0
cc_255 N_A2_M1012_g N_VGND_c_664_n 0.0082726f $X=4.35 $Y=0.655 $X2=0 $Y2=0
cc_256 N_A1_M1004_g N_VPWR_c_350_n 0.0160917f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A1_M1010_g N_VPWR_c_350_n 0.0167889f $X=5.67 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A1_M1004_g N_VPWR_c_352_n 0.00486043f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A1_M1010_g N_VPWR_c_353_n 0.00486043f $X=5.67 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A1_M1004_g N_VPWR_c_346_n 0.0082726f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A1_M1010_g N_VPWR_c_346_n 0.00925813f $X=5.67 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A1_M1004_g N_A_808_367#_c_549_n 0.0168101f $X=5.24 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A1_M1010_g N_A_808_367#_c_549_n 0.0122595f $X=5.67 $Y=2.465 $X2=0 $Y2=0
cc_264 A1 N_A_808_367#_c_549_n 0.0307003f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_265 N_A1_c_311_n N_A_808_367#_c_549_n 4.72037e-19 $X=5.67 $Y=1.385 $X2=0
+ $Y2=0
cc_266 A1 N_A_808_367#_c_540_n 0.0224548f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_267 N_A1_c_311_n N_A_808_367#_c_540_n 0.00136403f $X=5.67 $Y=1.385 $X2=0
+ $Y2=0
cc_268 N_A1_c_304_n N_A_155_47#_c_574_n 0.0126001f $X=4.78 $Y=1.185 $X2=0 $Y2=0
cc_269 N_A1_c_305_n N_A_155_47#_c_574_n 0.00229041f $X=5.135 $Y=1.26 $X2=0 $Y2=0
cc_270 N_A1_c_307_n N_A_155_47#_c_574_n 0.0180633f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_271 A1 N_A_155_47#_c_574_n 0.0246215f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_272 N_A1_c_311_n N_A_155_47#_c_574_n 0.0108004f $X=5.67 $Y=1.385 $X2=0 $Y2=0
cc_273 N_A1_c_304_n N_VGND_c_658_n 6.11179e-19 $X=4.78 $Y=1.185 $X2=0 $Y2=0
cc_274 N_A1_c_304_n N_VGND_c_659_n 0.010076f $X=4.78 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A1_c_307_n N_VGND_c_659_n 0.0119789f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A1_c_304_n N_VGND_c_662_n 0.00486043f $X=4.78 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A1_c_307_n N_VGND_c_663_n 0.00486043f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_278 N_A1_c_304_n N_VGND_c_664_n 0.0082726f $X=4.78 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A1_c_307_n N_VGND_c_664_n 0.00954696f $X=5.21 $Y=1.185 $X2=0 $Y2=0
cc_280 N_VPWR_c_346_n N_Y_M1009_s 0.00432284f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_281 N_VPWR_c_346_n N_Y_M1002_s 0.00225186f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_282 N_VPWR_c_351_n N_Y_c_448_n 0.0135169f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_346_n N_Y_c_448_n 0.00847534f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_284 N_VPWR_c_348_n N_Y_c_421_n 0.00166817f $X=0.31 $Y=1.98 $X2=0 $Y2=0
cc_285 N_VPWR_M1018_d Y 7.90388e-19 $X=1.03 $Y=1.835 $X2=0 $Y2=0
cc_286 N_VPWR_M1018_d N_Y_c_423_n 0.00161445f $X=1.03 $Y=1.835 $X2=0 $Y2=0
cc_287 N_VPWR_c_349_n N_Y_c_423_n 0.0226604f $X=1.17 $Y=2.13 $X2=0 $Y2=0
cc_288 N_VPWR_c_346_n N_A_313_365#_M1002_d 0.00212303f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_289 N_VPWR_c_346_n N_A_313_365#_M1011_d 0.00709847f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_290 N_VPWR_c_346_n N_A_313_365#_M1019_d 0.00213122f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_291 N_VPWR_c_349_n N_A_313_365#_c_466_n 0.0147176f $X=1.17 $Y=2.13 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_352_n N_A_313_365#_c_466_n 0.0179183f $X=5.29 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_346_n N_A_313_365#_c_466_n 0.0101082f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_294 N_VPWR_c_349_n N_A_313_365#_c_467_n 0.0642548f $X=1.17 $Y=2.13 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_352_n N_A_313_365#_c_472_n 0.062587f $X=5.29 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_c_346_n N_A_313_365#_c_472_n 0.0386766f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_297 N_VPWR_c_346_n N_A_615_365#_M1013_s 0.00223559f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_298 N_VPWR_c_346_n N_A_615_365#_M1000_s 0.00223559f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_299 N_VPWR_c_352_n N_A_615_365#_c_511_n 0.0821667f $X=5.29 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_346_n N_A_615_365#_c_511_n 0.0507876f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_301 N_VPWR_c_352_n N_A_615_365#_c_515_n 0.01906f $X=5.29 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_c_346_n N_A_615_365#_c_515_n 0.0124545f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_c_346_n N_A_808_367#_M1000_d 0.0021598f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_304 N_VPWR_c_346_n N_A_808_367#_M1006_d 0.00536646f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_305 N_VPWR_c_346_n N_A_808_367#_M1010_d 0.00371702f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_306 N_VPWR_c_352_n N_A_808_367#_c_558_n 0.0124525f $X=5.29 $Y=3.33 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_346_n N_A_808_367#_c_558_n 0.00730901f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_M1004_s N_A_808_367#_c_549_n 0.00335998f $X=5.315 $Y=1.835 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_350_n N_A_808_367#_c_549_n 0.0170777f $X=5.455 $Y=2.365 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_353_n N_A_808_367#_c_541_n 0.0178111f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_311 N_VPWR_c_346_n N_A_808_367#_c_541_n 0.0100304f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_312 Y N_A_313_365#_M1002_d 0.00252154f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_313 Y N_A_313_365#_c_467_n 0.021928f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_314 N_Y_M1002_s N_A_313_365#_c_472_n 0.00337224f $X=1.98 $Y=1.825 $X2=0 $Y2=0
cc_315 N_Y_c_437_n N_A_313_365#_c_472_n 0.0153017f $X=2.12 $Y=1.95 $X2=0 $Y2=0
cc_316 N_Y_c_437_n N_A_313_365#_c_474_n 0.0113112f $X=2.12 $Y=1.95 $X2=0 $Y2=0
cc_317 N_Y_c_437_n N_A_313_365#_c_477_n 0.0390852f $X=2.12 $Y=1.95 $X2=0 $Y2=0
cc_318 N_Y_M1007_d N_A_155_47#_c_581_n 0.00332344f $X=1.19 $Y=0.235 $X2=0 $Y2=0
cc_319 N_Y_c_419_n N_A_155_47#_c_581_n 0.0135951f $X=1.33 $Y=0.76 $X2=0 $Y2=0
cc_320 Y N_A_155_47#_c_570_n 0.0276124f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_321 N_Y_c_419_n N_A_155_47#_c_571_n 0.0102912f $X=1.33 $Y=0.76 $X2=0 $Y2=0
cc_322 Y N_A_155_47#_c_571_n 0.024225f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_323 N_Y_M1007_d N_VGND_c_664_n 0.00225186f $X=1.19 $Y=0.235 $X2=0 $Y2=0
cc_324 N_A_313_365#_c_478_n N_A_615_365#_M1013_s 0.00351994f $X=3.55 $Y=2.005
+ $X2=-0.19 $Y2=1.655
cc_325 N_A_313_365#_c_472_n N_A_615_365#_c_512_n 6.69721e-19 $X=2.51 $Y=2.985
+ $X2=0 $Y2=0
cc_326 N_A_313_365#_c_477_n N_A_615_365#_c_512_n 0.0418638f $X=2.675 $Y=2.46
+ $X2=0 $Y2=0
cc_327 N_A_313_365#_c_478_n N_A_615_365#_c_512_n 0.0170777f $X=3.55 $Y=2.005
+ $X2=0 $Y2=0
cc_328 N_A_313_365#_M1019_d N_A_615_365#_c_511_n 0.00495471f $X=3.505 $Y=1.825
+ $X2=0 $Y2=0
cc_329 N_A_313_365#_c_469_n N_A_615_365#_c_511_n 0.0189128f $X=3.645 $Y=2.57
+ $X2=0 $Y2=0
cc_330 N_A_313_365#_c_472_n N_A_615_365#_c_515_n 0.0126067f $X=2.51 $Y=2.985
+ $X2=0 $Y2=0
cc_331 N_A_313_365#_c_468_n N_A_808_367#_c_538_n 0.0147157f $X=3.68 $Y=2.09
+ $X2=0 $Y2=0
cc_332 N_A_313_365#_c_469_n N_A_808_367#_c_539_n 0.0478316f $X=3.645 $Y=2.57
+ $X2=0 $Y2=0
cc_333 N_A_615_365#_c_511_n N_A_808_367#_M1000_d 0.00495471f $X=4.43 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_334 N_A_615_365#_c_511_n N_A_808_367#_c_539_n 0.0189128f $X=4.43 $Y=2.99
+ $X2=0 $Y2=0
cc_335 N_A_615_365#_M1000_s N_A_808_367#_c_544_n 0.00331217f $X=4.455 $Y=1.835
+ $X2=0 $Y2=0
cc_336 N_A_615_365#_c_519_n N_A_808_367#_c_544_n 0.0170777f $X=4.595 $Y=2.365
+ $X2=0 $Y2=0
cc_337 N_A_155_47#_c_570_n N_VGND_M1015_d 0.004138f $X=2.62 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_338 N_A_155_47#_c_572_n N_VGND_M1001_d 0.00240242f $X=3.57 $Y=1.08 $X2=0
+ $Y2=0
cc_339 N_A_155_47#_c_573_n N_VGND_M1003_d 0.00176461f $X=4.47 $Y=1.08 $X2=0
+ $Y2=0
cc_340 N_A_155_47#_c_574_n N_VGND_M1005_s 0.00176461f $X=5.34 $Y=1.08 $X2=0
+ $Y2=0
cc_341 N_A_155_47#_c_570_n N_VGND_c_655_n 0.0261974f $X=2.62 $Y=1.08 $X2=0 $Y2=0
cc_342 N_A_155_47#_c_596_n N_VGND_c_655_n 0.0401245f $X=2.785 $Y=0.42 $X2=0
+ $Y2=0
cc_343 N_A_155_47#_c_596_n N_VGND_c_656_n 0.0163977f $X=2.785 $Y=0.42 $X2=0
+ $Y2=0
cc_344 N_A_155_47#_c_572_n N_VGND_c_657_n 0.0186496f $X=3.57 $Y=1.08 $X2=0 $Y2=0
cc_345 N_A_155_47#_c_573_n N_VGND_c_658_n 0.0170777f $X=4.47 $Y=1.08 $X2=0 $Y2=0
cc_346 N_A_155_47#_c_574_n N_VGND_c_659_n 0.0170777f $X=5.34 $Y=1.08 $X2=0 $Y2=0
cc_347 N_A_155_47#_c_581_n N_VGND_c_660_n 0.0326395f $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_348 N_A_155_47#_c_587_n N_VGND_c_660_n 0.0161465f $X=1.79 $Y=0.425 $X2=0
+ $Y2=0
cc_349 N_A_155_47#_c_576_n N_VGND_c_660_n 0.0209897f $X=0.9 $Y=0.39 $X2=0 $Y2=0
cc_350 N_A_155_47#_c_639_p N_VGND_c_661_n 0.0138717f $X=3.705 $Y=0.42 $X2=0
+ $Y2=0
cc_351 N_A_155_47#_c_640_p N_VGND_c_662_n 0.0124525f $X=4.565 $Y=0.42 $X2=0
+ $Y2=0
cc_352 N_A_155_47#_c_575_n N_VGND_c_663_n 0.0188625f $X=5.445 $Y=0.42 $X2=0
+ $Y2=0
cc_353 N_A_155_47#_M1007_s N_VGND_c_664_n 0.00215158f $X=0.775 $Y=0.235 $X2=0
+ $Y2=0
cc_354 N_A_155_47#_M1008_s N_VGND_c_664_n 0.00223561f $X=1.62 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_A_155_47#_M1016_s N_VGND_c_664_n 0.00310528f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_A_155_47#_M1014_s N_VGND_c_664_n 0.00397496f $X=3.565 $Y=0.235 $X2=0
+ $Y2=0
cc_357 N_A_155_47#_M1012_s N_VGND_c_664_n 0.00536646f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_358 N_A_155_47#_M1017_d N_VGND_c_664_n 0.00423245f $X=5.285 $Y=0.235 $X2=0
+ $Y2=0
cc_359 N_A_155_47#_c_581_n N_VGND_c_664_n 0.0208532f $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_360 N_A_155_47#_c_587_n N_VGND_c_664_n 0.0103094f $X=1.79 $Y=0.425 $X2=0
+ $Y2=0
cc_361 N_A_155_47#_c_596_n N_VGND_c_664_n 0.010625f $X=2.785 $Y=0.42 $X2=0 $Y2=0
cc_362 N_A_155_47#_c_639_p N_VGND_c_664_n 0.00886411f $X=3.705 $Y=0.42 $X2=0
+ $Y2=0
cc_363 N_A_155_47#_c_640_p N_VGND_c_664_n 0.00730901f $X=4.565 $Y=0.42 $X2=0
+ $Y2=0
cc_364 N_A_155_47#_c_575_n N_VGND_c_664_n 0.0104139f $X=5.445 $Y=0.42 $X2=0
+ $Y2=0
cc_365 N_A_155_47#_c_576_n N_VGND_c_664_n 0.0125952f $X=0.9 $Y=0.39 $X2=0 $Y2=0
