* File: sky130_fd_sc_lp__busdriver2_20.spice
* Created: Fri Aug 28 10:13:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__busdriver2_20.pex.spice"
.subckt sky130_fd_sc_lp__busdriver2_20  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_TE_B_M1020_g N_A_114_47#_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_TE_B_M1024_g N_A_114_47#_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1877 AS=0.1176 PD=1.3 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1024_d N_A_114_47#_M1010_g N_A_286_367#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1877 AS=0.23305 PD=1.3 PS=1.48 NRD=11.424 NRS=17.136 M=1 R=5.6
+ SA=75001.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1043 N_VGND_M1043_d N_A_114_47#_M1043_g N_A_286_367#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.365 AS=0.23305 PD=2.68 PS=1.48 NRD=17.136 NRS=17.136 M=1 R=5.6
+ SA=75001.9 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A_114_47#_M1003_g N_A_584_47#_M1003_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75012.5 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1003_d N_A_114_47#_M1011_g N_A_584_47#_M1011_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.0896 PD=1 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75011.9 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_A_114_47#_M1015_g N_A_584_47#_M1011_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75011.5 A=0.096 P=1.58 MULT=1
MM1016 N_VGND_M1015_d N_A_114_47#_M1016_g N_A_584_47#_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75011.1 A=0.096 P=1.58 MULT=1
MM1035 N_VGND_M1035_d N_A_114_47#_M1035_g N_A_584_47#_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.0896 PD=1 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002
+ SB=75010.7 A=0.096 P=1.58 MULT=1
MM1039 N_VGND_M1035_d N_A_114_47#_M1039_g N_A_584_47#_M1039_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.0896 PD=1 PS=0.92 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75002.5 SB=75010.2 A=0.096 P=1.58 MULT=1
MM1044 N_VGND_M1044_d N_A_114_47#_M1044_g N_A_584_47#_M1039_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1408 AS=0.0896 PD=1.08 PS=0.92 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75002.9 SB=75009.7 A=0.096 P=1.58 MULT=1
MM1045 N_VGND_M1044_d N_A_114_47#_M1045_g N_A_584_47#_M1045_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1408 AS=0.0896 PD=1.08 PS=0.92 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75003.5 SB=75009.1 A=0.096 P=1.58 MULT=1
MM1047 N_VGND_M1047_d N_A_114_47#_M1047_g N_A_584_47#_M1045_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004
+ SB=75008.7 A=0.096 P=1.58 MULT=1
MM1051 N_VGND_M1047_d N_A_114_47#_M1051_g N_A_584_47#_M1051_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.4 SB=75008.3 A=0.096 P=1.58 MULT=1
MM1057 N_VGND_M1057_d N_A_114_47#_M1057_g N_A_584_47#_M1051_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.8 SB=75007.8 A=0.096 P=1.58 MULT=1
MM1066 N_VGND_M1057_d N_A_114_47#_M1066_g N_A_584_47#_M1066_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75005.3 SB=75007.4 A=0.096 P=1.58 MULT=1
MM1070 N_VGND_M1070_d N_A_114_47#_M1070_g N_A_584_47#_M1066_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75005.7 SB=75007 A=0.096 P=1.58 MULT=1
MM1080 N_VGND_M1070_d N_A_114_47#_M1080_g N_A_584_47#_M1080_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75006.1 SB=75006.5 A=0.096 P=1.58 MULT=1
MM1017 N_A_584_47#_M1080_s N_A_1909_21#_M1017_g N_Z_M1017_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1152 PD=0.92 PS=1 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75006.5 SB=75006.1 A=0.096 P=1.58 MULT=1
MM1021 N_A_584_47#_M1021_d N_A_1909_21#_M1021_g N_Z_M1017_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.1152 PD=1 PS=1 NRD=14.988 NRS=0 M=1 R=4.26667 SA=75007.1
+ SB=75005.6 A=0.096 P=1.58 MULT=1
MM1027 N_A_584_47#_M1021_d N_A_1909_21#_M1027_g N_Z_M1027_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.1152 PD=1 PS=1 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75007.6
+ SB=75005.1 A=0.096 P=1.58 MULT=1
MM1031 N_A_584_47#_M1031_d N_A_1909_21#_M1031_g N_Z_M1027_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1152 PD=0.92 PS=1 NRD=0 NRS=0 M=1 R=4.26667 SA=75008.1
+ SB=75004.6 A=0.096 P=1.58 MULT=1
MM1033 N_A_584_47#_M1031_d N_A_1909_21#_M1033_g N_Z_M1033_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75008.5 SB=75004.2 A=0.096 P=1.58 MULT=1
MM1036 N_A_584_47#_M1036_d N_A_1909_21#_M1036_g N_Z_M1033_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75008.9 SB=75003.7 A=0.096 P=1.58 MULT=1
MM1048 N_A_584_47#_M1036_d N_A_1909_21#_M1048_g N_Z_M1048_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75009.4 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1053 N_A_584_47#_M1053_d N_A_1909_21#_M1053_g N_Z_M1048_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75009.8 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1059 N_A_584_47#_M1053_d N_A_1909_21#_M1059_g N_Z_M1059_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75010.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1060 N_A_584_47#_M1060_d N_A_1909_21#_M1060_g N_Z_M1059_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75010.7 SB=75002 A=0.096 P=1.58 MULT=1
MM1067 N_A_584_47#_M1060_d N_A_1909_21#_M1067_g N_Z_M1067_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75011.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1073 N_A_584_47#_M1073_d N_A_1909_21#_M1073_g N_Z_M1067_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75011.5 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1081 N_A_584_47#_M1073_d N_A_1909_21#_M1081_g N_Z_M1081_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75011.9 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1086 N_A_584_47#_M1086_d N_A_1909_21#_M1086_g N_Z_M1081_s VNB NSHORT L=0.15
+ W=0.64 AD=0.2336 AS=0.0896 PD=2.01 PS=0.92 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75012.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1028 N_A_1909_21#_M1028_d N_A_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1491 AS=0.2436 PD=1.195 PS=2.26 NRD=10.704 NRS=0.708 M=1 R=5.6 SA=75000.2
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1029 N_A_1909_21#_M1028_d N_A_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1491 AS=0.1848 PD=1.195 PS=1.28 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.7
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1082 N_A_1909_21#_M1082_d N_A_M1082_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1848 PD=1.12 PS=1.28 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1083 N_A_1909_21#_M1082_d N_A_M1083_g N_VGND_M1083_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3066 PD=1.12 PS=2.41 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.7
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_TE_B_M1004_g N_A_114_47#_M1004_s VPB PSHORT L=0.15
+ W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75011 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_TE_B_M1007_g N_A_114_47#_M1004_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75010.5 A=0.189 P=2.82 MULT=1
MM1049 N_A_286_367#_M1049_d N_A_114_47#_M1049_g N_VPWR_M1007_d VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75010.1 A=0.189 P=2.82 MULT=1
MM1054 N_A_286_367#_M1049_d N_A_114_47#_M1054_g N_VPWR_M1054_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75009.7 A=0.189 P=2.82 MULT=1
MM1068 N_A_286_367#_M1068_d N_A_114_47#_M1068_g N_VPWR_M1054_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75009.3 A=0.189 P=2.82 MULT=1
MM1071 N_A_286_367#_M1068_d N_A_114_47#_M1071_g N_VPWR_M1071_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75008.8 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1071_s N_A_286_367#_M1001_g N_A_630_367#_M1001_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75008.4 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_286_367#_M1005_g N_A_630_367#_M1001_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.2 SB=75008 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1005_d N_A_286_367#_M1012_g N_A_630_367#_M1012_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.6 SB=75007.5 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A_286_367#_M1018_g N_A_630_367#_M1012_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75007.1 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1018_d N_A_286_367#_M1019_g N_A_630_367#_M1019_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.5 SB=75006.7 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_286_367#_M1022_g N_A_630_367#_M1019_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.9 SB=75006.2 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1022_d N_A_286_367#_M1037_g N_A_630_367#_M1037_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75005.4 SB=75005.8 A=0.189 P=2.82 MULT=1
MM1040 N_VPWR_M1040_d N_A_286_367#_M1040_g N_A_630_367#_M1037_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75005.8 SB=75005.4 A=0.189 P=2.82 MULT=1
MM1041 N_VPWR_M1040_d N_A_286_367#_M1041_g N_A_630_367#_M1041_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75006.2 SB=75005 A=0.189 P=2.82 MULT=1
MM1055 N_VPWR_M1055_d N_A_286_367#_M1055_g N_A_630_367#_M1041_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75006.7 SB=75004.5 A=0.189 P=2.82 MULT=1
MM1058 N_VPWR_M1055_d N_A_286_367#_M1058_g N_A_630_367#_M1058_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75007.1 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1061 N_VPWR_M1061_d N_A_286_367#_M1061_g N_A_630_367#_M1058_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.189 AS=0.1764 PD=1.56 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75007.5 SB=75003.7 A=0.189 P=2.82 MULT=1
MM1064 N_VPWR_M1061_d N_A_286_367#_M1064_g N_A_630_367#_M1064_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.189 AS=0.1764 PD=1.56 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75008 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1065 N_VPWR_M1065_d N_A_286_367#_M1065_g N_A_630_367#_M1064_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75008.4 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1069 N_VPWR_M1065_d N_A_286_367#_M1069_g N_A_630_367#_M1069_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75008.8 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1074 N_VPWR_M1074_d N_A_286_367#_M1074_g N_A_630_367#_M1069_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75009.3 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1077 N_VPWR_M1074_d N_A_286_367#_M1077_g N_A_630_367#_M1077_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75009.7 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1084 N_VPWR_M1084_d N_A_286_367#_M1084_g N_A_630_367#_M1077_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75010.1 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1087 N_VPWR_M1084_d N_A_286_367#_M1087_g N_A_630_367#_M1087_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75010.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1089 N_VPWR_M1089_d N_A_286_367#_M1089_g N_A_630_367#_M1087_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75011 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_Z_M1000_d N_A_1909_21#_M1000_g N_A_630_367#_M1000_s VPB PSHORT L=0.15
+ W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75008.4 A=0.189 P=2.82 MULT=1
MM1002 N_Z_M1002_d N_A_1909_21#_M1002_g N_A_630_367#_M1000_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75007.9 A=0.189 P=2.82 MULT=1
MM1006 N_Z_M1002_d N_A_1909_21#_M1006_g N_A_630_367#_M1006_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75007.5 A=0.189 P=2.82 MULT=1
MM1008 N_Z_M1008_d N_A_1909_21#_M1008_g N_A_630_367#_M1006_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75007.1 A=0.189 P=2.82 MULT=1
MM1013 N_Z_M1008_d N_A_1909_21#_M1013_g N_A_630_367#_M1013_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75006.7 A=0.189 P=2.82 MULT=1
MM1023 N_Z_M1023_d N_A_1909_21#_M1023_g N_A_630_367#_M1013_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1025 N_Z_M1023_d N_A_1909_21#_M1025_g N_A_630_367#_M1025_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75005.8 A=0.189 P=2.82 MULT=1
MM1026 N_Z_M1026_d N_A_1909_21#_M1026_g N_A_630_367#_M1025_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75005.4 A=0.189 P=2.82 MULT=1
MM1030 N_Z_M1026_d N_A_1909_21#_M1030_g N_A_630_367#_M1030_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1032 N_Z_M1032_d N_A_1909_21#_M1032_g N_A_630_367#_M1030_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1038 N_Z_M1032_d N_A_1909_21#_M1038_g N_A_630_367#_M1038_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1042 N_Z_M1042_d N_A_1909_21#_M1042_g N_A_630_367#_M1038_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1046 N_Z_M1042_d N_A_1909_21#_M1046_g N_A_630_367#_M1046_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1050 N_Z_M1050_d N_A_1909_21#_M1050_g N_A_630_367#_M1046_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1056 N_Z_M1050_d N_A_1909_21#_M1056_g N_A_630_367#_M1056_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1062 N_Z_M1062_d N_A_1909_21#_M1062_g N_A_630_367#_M1056_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.7
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1063 N_Z_M1062_d N_A_1909_21#_M1063_g N_A_630_367#_M1063_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1075 N_Z_M1075_d N_A_1909_21#_M1075_g N_A_630_367#_M1063_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1078 N_Z_M1075_d N_A_1909_21#_M1078_g N_A_630_367#_M1078_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1088 N_Z_M1088_d N_A_1909_21#_M1088_g N_A_630_367#_M1078_s VPB PSHORT L=0.15
+ W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_A_1909_21#_M1009_s VPB PSHORT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_1909_21#_M1009_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1034 N_VPWR_M1014_d N_A_M1034_g N_A_1909_21#_M1034_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1052 N_VPWR_M1052_d N_A_M1052_g N_A_1909_21#_M1034_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1072 N_VPWR_M1052_d N_A_M1072_g N_A_1909_21#_M1072_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1076 N_VPWR_M1076_d N_A_M1076_g N_A_1909_21#_M1072_s VPB PSHORT L=0.15 W=1.26
+ AD=0.19215 AS=0.1764 PD=1.565 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1079 N_VPWR_M1076_d N_A_M1079_g N_A_1909_21#_M1079_s VPB PSHORT L=0.15 W=1.26
+ AD=0.19215 AS=0.1764 PD=1.565 PS=1.54 NRD=3.9006 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1085 N_VPWR_M1085_d N_A_M1085_g N_A_1909_21#_M1079_s VPB PSHORT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX90_noxref VNB VPB NWDIODE A=50.1266 P=55.03
c_388 VPB 0 1.47022e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__busdriver2_20.pxi.spice"
*
.ends
*
*
