* File: sky130_fd_sc_lp__a2111oi_1.pex.spice
* Created: Wed Sep  2 09:16:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111OI_1%D1 3 7 9 10 11 12 21 22
r32 20 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.62 $Y=1.51 $X2=0.71
+ $Y2=1.51
r33 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.51 $X2=0.62 $Y2=1.51
r34 17 20 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.525 $Y=1.51
+ $X2=0.62 $Y2=1.51
r35 11 12 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.695 $Y=2.405
+ $X2=0.695 $Y2=2.775
r36 10 11 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.695 $Y=2.035
+ $X2=0.695 $Y2=2.405
r37 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.695 $Y=1.665
+ $X2=0.695 $Y2=2.035
r38 9 21 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=0.695 $Y=1.665
+ $X2=0.695 $Y2=1.51
r39 5 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.71 $Y=1.675
+ $X2=0.71 $Y2=1.51
r40 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.71 $Y=1.675 $X2=0.71
+ $Y2=2.465
r41 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.345
+ $X2=0.525 $Y2=1.51
r42 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.525 $Y=1.345
+ $X2=0.525 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%C1 3 7 9 10 11 12 13 20
r38 20 23 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.375
+ $X2=1.175 $Y2=1.54
r39 20 22 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.375
+ $X2=1.175 $Y2=1.21
r40 12 13 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=2.405
+ $X2=1.17 $Y2=2.775
r41 11 12 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=2.035
+ $X2=1.17 $Y2=2.405
r42 10 11 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=2.035
r43 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.295
+ $X2=1.17 $Y2=1.665
r44 9 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.375 $X2=1.19 $Y2=1.375
r45 7 23 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.19 $Y=2.465
+ $X2=1.19 $Y2=1.54
r46 3 22 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.07 $Y=0.655
+ $X2=1.07 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%B1 3 5 7 8 15
r32 13 15 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.73 $Y=1.355
+ $X2=1.85 $Y2=1.355
r33 10 13 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.64 $Y=1.355 $X2=1.73
+ $Y2=1.355
r34 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.355 $X2=1.73 $Y2=1.355
r35 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.19
+ $X2=1.85 $Y2=1.355
r36 5 7 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.85 $Y=1.19 $X2=1.85
+ $Y2=0.655
r37 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.64 $Y=1.52
+ $X2=1.64 $Y2=1.355
r38 1 3 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.64 $Y=1.52 $X2=1.64
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%A1 3 5 7 8 9 17
r32 15 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.33 $Y=1.35 $X2=2.42
+ $Y2=1.35
r33 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.35 $X2=2.33 $Y2=1.35
r34 12 15 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.21 $Y=1.35
+ $X2=2.33 $Y2=1.35
r35 9 16 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.64 $Y=1.35 $X2=2.33
+ $Y2=1.35
r36 8 16 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.35 $X2=2.33
+ $Y2=1.35
r37 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.185
+ $X2=2.42 $Y2=1.35
r38 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.42 $Y=1.185 $X2=2.42
+ $Y2=0.655
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.515
+ $X2=2.21 $Y2=1.35
r40 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.21 $Y=1.515 $X2=2.21
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%A2 1 3 6 8 13
r24 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.355 $X2=2.99 $Y2=1.355
r25 10 13 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.78 $Y=1.355
+ $X2=2.99 $Y2=1.355
r26 8 14 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.355
+ $X2=2.99 $Y2=1.355
r27 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=1.52
+ $X2=2.78 $Y2=1.355
r28 4 6 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=2.78 $Y=1.52 $X2=2.78
+ $Y2=2.465
r29 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=1.19
+ $X2=2.78 $Y2=1.355
r30 1 3 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.78 $Y=1.19 $X2=2.78
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%Y 1 2 3 12 16 17 18 19 20 21 37 46 50
r43 49 50 10.894 $w=7.58e-07 $l=1.6e-07 $layer=LI1_cond $X=2.13 $Y=0.635
+ $X2=1.97 $Y2=0.635
r44 46 47 6.07829 $w=2.81e-07 $l=1.4e-07 $layer=LI1_cond $X=0.8 $Y=0.93 $X2=0.8
+ $Y2=1.07
r45 44 46 0.130249 $w=2.81e-07 $l=3e-09 $layer=LI1_cond $X=0.8 $Y=0.927 $X2=0.8
+ $Y2=0.93
r46 30 44 3.52958 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0.927
+ $X2=0.8 $Y2=0.927
r47 20 21 7.55418 $w=7.58e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.635
+ $X2=2.64 $Y2=0.635
r48 20 49 0.472136 $w=7.58e-07 $l=3e-08 $layer=LI1_cond $X=2.16 $Y=0.635
+ $X2=2.13 $Y2=0.635
r49 19 50 18.3792 $w=1.73e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=0.927
+ $X2=1.97 $Y2=0.927
r50 18 19 30.4208 $w=1.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.927
+ $X2=1.68 $Y2=0.927
r51 18 30 14.8935 $w=1.73e-07 $l=2.35e-07 $layer=LI1_cond $X=1.2 $Y=0.927
+ $X2=0.965 $Y2=0.927
r52 17 47 3.67734 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=1.07
+ $X2=0.8 $Y2=1.07
r53 17 44 0.0868327 $w=2.81e-07 $l=2e-09 $layer=LI1_cond $X=0.8 $Y=0.925 $X2=0.8
+ $Y2=0.927
r54 17 37 11.4308 $w=4.98e-07 $l=4.2e-07 $layer=LI1_cond $X=0.8 $Y=0.84 $X2=0.8
+ $Y2=0.42
r55 16 17 15.5683 $w=1.93e-07 $l=2.7e-07 $layer=LI1_cond $X=0.365 $Y=1.07
+ $X2=0.635 $Y2=1.07
r56 12 14 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=0.24 $Y=1.98
+ $X2=0.24 $Y2=2.91
r57 10 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.155
+ $X2=0.365 $Y2=1.07
r58 10 12 38.0306 $w=2.48e-07 $l=8.25e-07 $layer=LI1_cond $X=0.24 $Y=1.155
+ $X2=0.24 $Y2=1.98
r59 3 14 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=2.91
r60 3 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=1.98
r61 2 49 91 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=2 $X=1.925
+ $Y=0.235 $X2=2.13 $Y2=0.42
r62 1 46 182 $w=1.7e-07 $l=7.88686e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.8 $Y2=0.93
r63 1 37 182 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.8 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%A_343_367# 1 2 9 13 14 17
r22 17 19 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.025 $Y=1.98
+ $X2=3.025 $Y2=2.91
r23 15 17 2.34757 $w=2.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.025 $Y=1.925
+ $X2=3.025 $Y2=1.98
r24 13 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.89 $Y=1.84
+ $X2=3.025 $Y2=1.925
r25 13 14 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.89 $Y=1.84
+ $X2=2.095 $Y2=1.84
r26 9 11 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=1.93 $Y=1.98 $X2=1.93
+ $Y2=2.91
r27 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.93 $Y=1.925
+ $X2=2.095 $Y2=1.84
r28 7 9 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.93 $Y=1.925 $X2=1.93
+ $Y2=1.98
r29 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.835 $X2=2.995 $Y2=2.91
r30 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.835 $X2=2.995 $Y2=1.98
r31 1 11 400 $w=1.7e-07 $l=1.1776e-06 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.835 $X2=1.93 $Y2=2.91
r32 1 9 400 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.835 $X2=1.93 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%VPWR 1 6 11 12 13 23 24
r35 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 16 20 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 13 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 13 17 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 11 20 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 11 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.49 $Y2=3.33
r44 10 23 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 10 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=2.49 $Y2=3.33
r46 6 9 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.49 $Y=2.19 $X2=2.49
+ $Y2=2.95
r47 4 12 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=3.245 $X2=2.49
+ $Y2=3.33
r48 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=2.95
r49 1 9 400 $w=1.7e-07 $l=1.21318e-06 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.49 $Y2=2.95
r50 1 6 400 $w=1.7e-07 $l=4.4587e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.49 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_1%VGND 1 2 3 10 12 14 16 18 20 22 41
r38 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 29 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r40 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 26 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r42 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 23 25 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=2.64
+ $Y2=0
r44 22 40 4.0325 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=3.127
+ $Y2=0
r45 22 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=2.64
+ $Y2=0
r46 20 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r47 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r48 16 40 3.21557 $w=2.65e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.027 $Y=0.085
+ $X2=3.127 $Y2=0
r49 16 18 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=3.027 $Y=0.085
+ $X2=3.027 $Y2=0.38
r50 15 28 4.68787 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.232
+ $Y2=0
r51 14 37 6.47501 $w=6.63e-07 $l=3.6e-07 $layer=LI1_cond $X=1.467 $Y=0 $X2=1.467
+ $Y2=0.36
r52 14 23 8.98481 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=1.467 $Y=0 $X2=1.8
+ $Y2=0
r53 14 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 14 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.465
+ $Y2=0
r56 10 28 3.0783 $w=3.3e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.232 $Y2=0
r57 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.3 $Y2=0.36
r58 3 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.855
+ $Y=0.235 $X2=2.995 $Y2=0.38
r59 2 37 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.145
+ $Y=0.235 $X2=1.285 $Y2=0.36
r60 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.3 $Y2=0.36
.ends

