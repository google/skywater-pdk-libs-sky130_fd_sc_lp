* File: sky130_fd_sc_lp__a2bb2o_lp.pxi.spice
* Created: Fri Aug 28 09:56:07 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%B2 N_B2_M1008_g N_B2_M1009_g N_B2_c_100_n
+ N_B2_c_105_n B2 B2 N_B2_c_102_n PM_SKY130_FD_SC_LP__A2BB2O_LP%B2
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%B1 N_B1_M1007_g N_B1_c_135_n N_B1_M1002_g
+ N_B1_c_140_n B1 B1 N_B1_c_137_n PM_SKY130_FD_SC_LP__A2BB2O_LP%B1
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%A_284_31# N_A_284_31#_M1013_d
+ N_A_284_31#_M1015_d N_A_284_31#_c_179_n N_A_284_31#_M1012_g
+ N_A_284_31#_c_180_n N_A_284_31#_c_181_n N_A_284_31#_c_182_n
+ N_A_284_31#_M1005_g N_A_284_31#_c_183_n N_A_284_31#_M1014_g
+ N_A_284_31#_c_192_n N_A_284_31#_c_184_n N_A_284_31#_c_185_n
+ N_A_284_31#_c_186_n N_A_284_31#_c_193_n N_A_284_31#_c_194_n
+ N_A_284_31#_c_211_p N_A_284_31#_c_187_n N_A_284_31#_c_196_n
+ N_A_284_31#_c_188_n N_A_284_31#_c_197_n N_A_284_31#_c_189_n
+ PM_SKY130_FD_SC_LP__A2BB2O_LP%A_284_31#
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%A_63_57# N_A_63_57#_M1009_s N_A_63_57#_M1014_d
+ N_A_63_57#_M1005_d N_A_63_57#_c_291_n N_A_63_57#_c_292_n N_A_63_57#_M1010_g
+ N_A_63_57#_M1003_g N_A_63_57#_M1011_g N_A_63_57#_c_296_n N_A_63_57#_c_297_n
+ N_A_63_57#_c_298_n N_A_63_57#_c_299_n N_A_63_57#_c_300_n N_A_63_57#_c_301_n
+ N_A_63_57#_c_302_n N_A_63_57#_c_306_n N_A_63_57#_c_303_n N_A_63_57#_c_304_n
+ PM_SKY130_FD_SC_LP__A2BB2O_LP%A_63_57#
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%A1_N N_A1_N_M1000_g N_A1_N_M1006_g
+ N_A1_N_M1013_g N_A1_N_c_388_n N_A1_N_c_389_n A1_N A1_N A1_N N_A1_N_c_391_n
+ PM_SKY130_FD_SC_LP__A2BB2O_LP%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%A2_N N_A2_N_c_429_n N_A2_N_M1015_g
+ N_A2_N_M1001_g N_A2_N_M1004_g A2_N A2_N PM_SKY130_FD_SC_LP__A2BB2O_LP%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%A_43_408# N_A_43_408#_M1008_s
+ N_A_43_408#_M1002_d N_A_43_408#_c_460_n N_A_43_408#_c_461_n
+ N_A_43_408#_c_462_n N_A_43_408#_c_463_n N_A_43_408#_c_464_n
+ PM_SKY130_FD_SC_LP__A2BB2O_LP%A_43_408#
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%VPWR N_VPWR_M1008_d N_VPWR_M1003_d
+ N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n VPWR
+ N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_493_n N_VPWR_c_501_n
+ PM_SKY130_FD_SC_LP__A2BB2O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%X N_X_M1010_s N_X_M1003_s N_X_c_538_n
+ N_X_c_539_n X PM_SKY130_FD_SC_LP__A2BB2O_LP%X
x_PM_SKY130_FD_SC_LP__A2BB2O_LP%VGND N_VGND_M1007_d N_VGND_M1011_d
+ N_VGND_M1004_d N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n N_VGND_c_573_n
+ N_VGND_c_574_n N_VGND_c_575_n VGND N_VGND_c_576_n N_VGND_c_577_n
+ N_VGND_c_578_n N_VGND_c_579_n PM_SKY130_FD_SC_LP__A2BB2O_LP%VGND
cc_1 VNB N_B2_M1009_g 0.044572f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.495
cc_2 VNB N_B2_c_100_n 0.023992f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.675
cc_3 VNB B2 0.0338014f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_B2_c_102_n 0.0170897f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.335
cc_5 VNB N_B1_M1007_g 0.0378774f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.54
cc_6 VNB N_B1_c_135_n 0.0225316f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.495
cc_7 VNB B1 0.00195292f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.84
cc_8 VNB N_B1_c_137_n 0.0187949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_284_31#_c_179_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.495
cc_10 VNB N_A_284_31#_c_180_n 0.00690297f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.17
cc_11 VNB N_A_284_31#_c_181_n 0.00893405f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.675
cc_12 VNB N_A_284_31#_c_182_n 0.0206175f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VNB N_A_284_31#_c_183_n 0.0175316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_284_31#_c_184_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.505
cc_15 VNB N_A_284_31#_c_185_n 0.00425489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_284_31#_c_186_n 0.0136769f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.505
cc_17 VNB N_A_284_31#_c_187_n 0.013833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_284_31#_c_188_n 0.00559537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_284_31#_c_189_n 0.0104933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_63_57#_c_291_n 0.0179504f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.17
cc_21 VNB N_A_63_57#_c_292_n 0.0164086f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.675
cc_22 VNB N_A_63_57#_M1010_g 0.0247981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_63_57#_M1003_g 0.0365373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_63_57#_M1011_g 0.0202881f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.335
cc_25 VNB N_A_63_57#_c_296_n 0.0200691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_63_57#_c_297_n 0.0238089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_63_57#_c_298_n 0.0234418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_63_57#_c_299_n 0.0100362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_63_57#_c_300_n 0.00818263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_63_57#_c_301_n 0.0200553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_63_57#_c_302_n 0.00177279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_63_57#_c_303_n 0.0367723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_63_57#_c_304_n 0.00116729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_N_M1000_g 0.029697f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.54
cc_35 VNB N_A1_N_M1013_g 0.0302333f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.675
cc_36 VNB N_A1_N_c_388_n 0.0191909f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_37 VNB N_A1_N_c_389_n 7.4711e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB A1_N 0.00696332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A1_N_c_391_n 0.0242634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A2_N_c_429_n 0.0652618f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.84
cc_41 VNB N_A2_N_M1001_g 0.0269352f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.495
cc_42 VNB N_A2_N_M1004_g 0.0368478f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.675
cc_43 VNB A2_N 0.0280389f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_44 VNB N_VPWR_c_493_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_538_n 0.0125801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_X_c_539_n 0.00900679f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.17
cc_47 VNB N_VGND_c_570_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.84
cc_48 VNB N_VGND_c_571_n 0.0133063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_572_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_573_n 0.0305954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_574_n 0.0506406f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.335
cc_52 VNB N_VGND_c_575_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.505
cc_53 VNB N_VGND_c_576_n 0.0338812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_577_n 0.0368355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_578_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_579_n 0.324687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VPB N_B2_M1008_g 0.0365844f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.54
cc_58 VPB N_B2_c_100_n 0.00142899f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.675
cc_59 VPB N_B2_c_105_n 0.0144588f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.84
cc_60 VPB B2 0.0152727f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_61 VPB N_B1_c_135_n 5.13749e-19 $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.495
cc_62 VPB N_B1_M1002_g 0.0284536f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.335
cc_63 VPB N_B1_c_140_n 0.0158835f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.675
cc_64 VPB B1 7.45523e-19 $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.84
cc_65 VPB N_A_284_31#_c_182_n 9.119e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_66 VPB N_A_284_31#_M1005_g 0.0340727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_284_31#_c_192_n 0.0168564f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.335
cc_68 VPB N_A_284_31#_c_193_n 0.00186372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_284_31#_c_194_n 0.0151227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_284_31#_c_187_n 0.00231366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_284_31#_c_196_n 0.00158259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_284_31#_c_197_n 0.0472272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_63_57#_M1003_g 0.0483504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_63_57#_c_306_n 0.010799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_63_57#_c_303_n 0.00972198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_63_57#_c_304_n 0.00222653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A1_N_M1006_g 0.0286248f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.495
cc_78 VPB N_A1_N_c_389_n 0.0191349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB A1_N 0.00357979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A2_N_c_429_n 0.0272239f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.84
cc_81 VPB N_A2_N_M1015_g 0.0409917f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.54
cc_82 VPB A2_N 0.0175928f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_83 VPB N_A_43_408#_c_460_n 0.00978367f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.495
cc_84 VPB N_A_43_408#_c_461_n 0.0353469f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.335
cc_85 VPB N_A_43_408#_c_462_n 0.00645794f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.675
cc_86 VPB N_A_43_408#_c_463_n 0.0103066f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_87 VPB N_A_43_408#_c_464_n 0.00254768f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_88 VPB N_VPWR_c_494_n 0.0019051f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.335
cc_89 VPB N_VPWR_c_495_n 0.00726456f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_90 VPB N_VPWR_c_496_n 0.0215329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_497_n 0.00503999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_498_n 0.0622194f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.505
cc_93 VPB N_VPWR_c_499_n 0.0464059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_493_n 0.0900866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_501_n 0.00631622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_X_c_538_n 0.00692012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB X 0.0131963f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_98 N_B2_M1009_g N_B1_M1007_g 0.0223199f $X=0.675 $Y=0.495 $X2=0 $Y2=0
cc_99 N_B2_c_100_n N_B1_c_135_n 0.0223199f $X=0.585 $Y=1.675 $X2=0 $Y2=0
cc_100 N_B2_M1008_g N_B1_M1002_g 0.030269f $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_101 N_B2_c_105_n N_B1_c_140_n 0.0223199f $X=0.585 $Y=1.84 $X2=0 $Y2=0
cc_102 B2 B1 0.0540818f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B2_c_102_n B1 6.90539e-19 $X=0.585 $Y=1.335 $X2=0 $Y2=0
cc_104 B2 N_B1_c_137_n 0.00463625f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B2_c_102_n N_B1_c_137_n 0.0223199f $X=0.585 $Y=1.335 $X2=0 $Y2=0
cc_106 N_B2_M1009_g N_A_63_57#_c_297_n 0.0129f $X=0.675 $Y=0.495 $X2=0 $Y2=0
cc_107 N_B2_M1009_g N_A_63_57#_c_298_n 0.00826241f $X=0.675 $Y=0.495 $X2=0 $Y2=0
cc_108 B2 N_A_63_57#_c_298_n 0.0158633f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B2_M1009_g N_A_63_57#_c_299_n 0.00420809f $X=0.675 $Y=0.495 $X2=0 $Y2=0
cc_110 B2 N_A_63_57#_c_299_n 0.0284747f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B2_c_102_n N_A_63_57#_c_299_n 0.0048437f $X=0.585 $Y=1.335 $X2=0 $Y2=0
cc_112 N_B2_M1008_g N_A_43_408#_c_460_n 0.00114325f $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_113 N_B2_c_105_n N_A_43_408#_c_460_n 0.00213543f $X=0.585 $Y=1.84 $X2=0 $Y2=0
cc_114 B2 N_A_43_408#_c_460_n 0.028933f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B2_M1008_g N_A_43_408#_c_461_n 0.0157595f $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_116 N_B2_M1008_g N_A_43_408#_c_462_n 0.0178604f $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_117 B2 N_A_43_408#_c_462_n 0.0230943f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B2_M1008_g N_A_43_408#_c_464_n 8.93705e-19 $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_119 N_B2_M1008_g N_VPWR_c_494_n 0.0174741f $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_120 N_B2_M1008_g N_VPWR_c_496_n 0.00762416f $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_121 N_B2_M1008_g N_VPWR_c_493_n 0.0140677f $X=0.625 $Y=2.54 $X2=0 $Y2=0
cc_122 N_B2_M1009_g N_VGND_c_570_n 0.00189174f $X=0.675 $Y=0.495 $X2=0 $Y2=0
cc_123 N_B2_M1009_g N_VGND_c_576_n 0.00502664f $X=0.675 $Y=0.495 $X2=0 $Y2=0
cc_124 N_B2_M1009_g N_VGND_c_579_n 0.00643675f $X=0.675 $Y=0.495 $X2=0 $Y2=0
cc_125 N_B1_M1007_g N_A_284_31#_c_179_n 0.0199179f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_126 N_B1_c_135_n N_A_284_31#_c_182_n 0.0116663f $X=1.167 $Y=1.663 $X2=0 $Y2=0
cc_127 N_B1_M1002_g N_A_284_31#_M1005_g 0.014813f $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_128 N_B1_c_140_n N_A_284_31#_c_192_n 0.0116663f $X=1.167 $Y=1.84 $X2=0 $Y2=0
cc_129 B1 N_A_284_31#_c_185_n 0.0362729f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B1_c_137_n N_A_284_31#_c_185_n 0.00121792f $X=1.18 $Y=1.335 $X2=0 $Y2=0
cc_131 B1 N_A_284_31#_c_186_n 0.00250411f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_c_137_n N_A_284_31#_c_186_n 0.0116663f $X=1.18 $Y=1.335 $X2=0 $Y2=0
cc_133 N_B1_M1002_g N_A_284_31#_c_193_n 9.59722e-19 $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_134 N_B1_c_135_n N_A_284_31#_c_196_n 0.00121792f $X=1.167 $Y=1.663 $X2=0
+ $Y2=0
cc_135 N_B1_M1007_g N_A_284_31#_c_189_n 0.0014213f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_136 N_B1_M1007_g N_A_63_57#_c_297_n 0.00195075f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_137 N_B1_M1007_g N_A_63_57#_c_298_n 0.0128937f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_138 B1 N_A_63_57#_c_298_n 0.0245995f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_139 N_B1_c_137_n N_A_63_57#_c_298_n 0.00140226f $X=1.18 $Y=1.335 $X2=0 $Y2=0
cc_140 N_B1_M1002_g N_A_43_408#_c_461_n 8.93705e-19 $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_141 N_B1_M1002_g N_A_43_408#_c_462_n 0.0178513f $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_142 N_B1_c_140_n N_A_43_408#_c_462_n 0.00116377f $X=1.167 $Y=1.84 $X2=0 $Y2=0
cc_143 B1 N_A_43_408#_c_462_n 0.0173841f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_144 N_B1_M1002_g N_A_43_408#_c_463_n 9.98113e-19 $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_145 N_B1_c_140_n N_A_43_408#_c_463_n 4.97464e-19 $X=1.167 $Y=1.84 $X2=0 $Y2=0
cc_146 B1 N_A_43_408#_c_463_n 0.00747547f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B1_M1002_g N_A_43_408#_c_464_n 0.0155857f $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_148 N_B1_M1002_g N_VPWR_c_494_n 0.0163971f $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_149 N_B1_M1002_g N_VPWR_c_498_n 0.00762416f $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_150 N_B1_M1002_g N_VPWR_c_493_n 0.013463f $X=1.155 $Y=2.54 $X2=0 $Y2=0
cc_151 N_B1_M1007_g N_VGND_c_570_n 0.0108215f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_152 N_B1_M1007_g N_VGND_c_576_n 0.00445056f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_153 N_B1_M1007_g N_VGND_c_579_n 0.00426841f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_154 N_A_284_31#_c_193_n N_A_63_57#_M1005_d 0.00955878f $X=1.85 $Y=2.495 $X2=0
+ $Y2=0
cc_155 N_A_284_31#_c_194_n N_A_63_57#_M1005_d 0.0227733f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_156 N_A_284_31#_c_211_p N_A_63_57#_M1005_d 7.93348e-19 $X=1.935 $Y=2.58 $X2=0
+ $Y2=0
cc_157 N_A_284_31#_c_189_n N_A_63_57#_c_292_n 0.0183106f $X=1.757 $Y=1.17 $X2=0
+ $Y2=0
cc_158 N_A_284_31#_c_194_n N_A_63_57#_M1003_g 0.0225979f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_159 N_A_284_31#_c_180_n N_A_63_57#_c_298_n 0.00790839f $X=1.78 $Y=0.855 $X2=0
+ $Y2=0
cc_160 N_A_284_31#_c_181_n N_A_63_57#_c_298_n 0.00834857f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_161 N_A_284_31#_c_184_n N_A_63_57#_c_298_n 0.00411533f $X=1.855 $Y=0.855
+ $X2=0 $Y2=0
cc_162 N_A_284_31#_c_185_n N_A_63_57#_c_298_n 0.0227416f $X=1.765 $Y=1.335 $X2=0
+ $Y2=0
cc_163 N_A_284_31#_c_186_n N_A_63_57#_c_298_n 8.8427e-19 $X=1.765 $Y=1.335 $X2=0
+ $Y2=0
cc_164 N_A_284_31#_c_189_n N_A_63_57#_c_298_n 0.00242022f $X=1.757 $Y=1.17 $X2=0
+ $Y2=0
cc_165 N_A_284_31#_c_179_n N_A_63_57#_c_300_n 0.00171786f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_166 N_A_284_31#_c_183_n N_A_63_57#_c_300_n 0.0110761f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_167 N_A_284_31#_c_184_n N_A_63_57#_c_300_n 0.00262536f $X=1.855 $Y=0.855
+ $X2=0 $Y2=0
cc_168 N_A_284_31#_c_184_n N_A_63_57#_c_301_n 0.00256035f $X=1.855 $Y=0.855
+ $X2=0 $Y2=0
cc_169 N_A_284_31#_c_185_n N_A_63_57#_c_301_n 0.00335618f $X=1.765 $Y=1.335
+ $X2=0 $Y2=0
cc_170 N_A_284_31#_c_189_n N_A_63_57#_c_301_n 0.00611099f $X=1.757 $Y=1.17 $X2=0
+ $Y2=0
cc_171 N_A_284_31#_c_185_n N_A_63_57#_c_302_n 0.0296754f $X=1.765 $Y=1.335 $X2=0
+ $Y2=0
cc_172 N_A_284_31#_c_186_n N_A_63_57#_c_302_n 9.9186e-19 $X=1.765 $Y=1.335 $X2=0
+ $Y2=0
cc_173 N_A_284_31#_M1005_g N_A_63_57#_c_306_n 0.00279f $X=1.71 $Y=2.54 $X2=0
+ $Y2=0
cc_174 N_A_284_31#_c_192_n N_A_63_57#_c_306_n 9.9186e-19 $X=1.757 $Y=1.84 $X2=0
+ $Y2=0
cc_175 N_A_284_31#_c_193_n N_A_63_57#_c_306_n 0.0296754f $X=1.85 $Y=2.495 $X2=0
+ $Y2=0
cc_176 N_A_284_31#_c_194_n N_A_63_57#_c_306_n 0.0267445f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_177 N_A_284_31#_c_185_n N_A_63_57#_c_303_n 0.00148926f $X=1.765 $Y=1.335
+ $X2=0 $Y2=0
cc_178 N_A_284_31#_c_186_n N_A_63_57#_c_303_n 0.0183106f $X=1.765 $Y=1.335 $X2=0
+ $Y2=0
cc_179 N_A_284_31#_c_182_n N_A_63_57#_c_304_n 9.9186e-19 $X=1.757 $Y=1.668 $X2=0
+ $Y2=0
cc_180 N_A_284_31#_c_196_n N_A_63_57#_c_304_n 0.0296754f $X=1.767 $Y=1.84 $X2=0
+ $Y2=0
cc_181 N_A_284_31#_c_188_n N_A1_N_M1000_g 0.00125204f $X=4.21 $Y=0.58 $X2=0
+ $Y2=0
cc_182 N_A_284_31#_c_194_n N_A1_N_M1006_g 0.021248f $X=4.095 $Y=2.58 $X2=0 $Y2=0
cc_183 N_A_284_31#_c_197_n N_A1_N_M1006_g 0.0126697f $X=4.43 $Y=2.58 $X2=0 $Y2=0
cc_184 N_A_284_31#_c_187_n N_A1_N_M1013_g 0.0108049f $X=4.18 $Y=2.025 $X2=0
+ $Y2=0
cc_185 N_A_284_31#_c_188_n N_A1_N_M1013_g 0.0095073f $X=4.21 $Y=0.58 $X2=0 $Y2=0
cc_186 N_A_284_31#_c_194_n N_A1_N_c_389_n 4.6718e-19 $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_187 N_A_284_31#_c_194_n A1_N 0.0158221f $X=4.095 $Y=2.58 $X2=0 $Y2=0
cc_188 N_A_284_31#_c_187_n A1_N 0.0562845f $X=4.18 $Y=2.025 $X2=0 $Y2=0
cc_189 N_A_284_31#_c_197_n A1_N 0.00908753f $X=4.43 $Y=2.58 $X2=0 $Y2=0
cc_190 N_A_284_31#_c_187_n N_A1_N_c_391_n 0.00507185f $X=4.18 $Y=2.025 $X2=0
+ $Y2=0
cc_191 N_A_284_31#_c_187_n N_A2_N_c_429_n 0.0106575f $X=4.18 $Y=2.025 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_284_31#_c_188_n N_A2_N_c_429_n 0.00160257f $X=4.21 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_284_31#_c_197_n N_A2_N_c_429_n 0.0079208f $X=4.43 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_284_31#_c_187_n N_A2_N_M1015_g 0.0101294f $X=4.18 $Y=2.025 $X2=0
+ $Y2=0
cc_195 N_A_284_31#_c_197_n N_A2_N_M1015_g 0.0454772f $X=4.43 $Y=2.58 $X2=0 $Y2=0
cc_196 N_A_284_31#_c_187_n N_A2_N_M1001_g 0.00574025f $X=4.18 $Y=2.025 $X2=0
+ $Y2=0
cc_197 N_A_284_31#_c_188_n N_A2_N_M1001_g 0.00957398f $X=4.21 $Y=0.58 $X2=0
+ $Y2=0
cc_198 N_A_284_31#_c_188_n N_A2_N_M1004_g 0.00125204f $X=4.21 $Y=0.58 $X2=0
+ $Y2=0
cc_199 N_A_284_31#_c_187_n A2_N 0.050495f $X=4.18 $Y=2.025 $X2=0 $Y2=0
cc_200 N_A_284_31#_c_197_n A2_N 0.0215025f $X=4.43 $Y=2.58 $X2=0 $Y2=0
cc_201 N_A_284_31#_M1005_g N_A_43_408#_c_463_n 2.0617e-19 $X=1.71 $Y=2.54 $X2=0
+ $Y2=0
cc_202 N_A_284_31#_c_193_n N_A_43_408#_c_463_n 0.0130523f $X=1.85 $Y=2.495 $X2=0
+ $Y2=0
cc_203 N_A_284_31#_M1005_g N_A_43_408#_c_464_n 5.70954e-19 $X=1.71 $Y=2.54 $X2=0
+ $Y2=0
cc_204 N_A_284_31#_c_193_n N_A_43_408#_c_464_n 0.021988f $X=1.85 $Y=2.495 $X2=0
+ $Y2=0
cc_205 N_A_284_31#_c_211_p N_A_43_408#_c_464_n 0.0136579f $X=1.935 $Y=2.58 $X2=0
+ $Y2=0
cc_206 N_A_284_31#_c_194_n N_VPWR_M1003_d 0.0122579f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_207 N_A_284_31#_M1005_g N_VPWR_c_494_n 8.03539e-19 $X=1.71 $Y=2.54 $X2=0
+ $Y2=0
cc_208 N_A_284_31#_c_194_n N_VPWR_c_495_n 0.0250819f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_209 N_A_284_31#_c_197_n N_VPWR_c_495_n 0.00356577f $X=4.43 $Y=2.58 $X2=0
+ $Y2=0
cc_210 N_A_284_31#_M1005_g N_VPWR_c_498_n 0.00817297f $X=1.71 $Y=2.54 $X2=0
+ $Y2=0
cc_211 N_A_284_31#_c_194_n N_VPWR_c_498_n 0.0220375f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_212 N_A_284_31#_c_211_p N_VPWR_c_498_n 0.00245843f $X=1.935 $Y=2.58 $X2=0
+ $Y2=0
cc_213 N_A_284_31#_c_194_n N_VPWR_c_499_n 0.00592116f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_214 N_A_284_31#_c_197_n N_VPWR_c_499_n 0.0355167f $X=4.43 $Y=2.58 $X2=0 $Y2=0
cc_215 N_A_284_31#_M1005_g N_VPWR_c_493_n 0.0152375f $X=1.71 $Y=2.54 $X2=0 $Y2=0
cc_216 N_A_284_31#_c_194_n N_VPWR_c_493_n 0.0500443f $X=4.095 $Y=2.58 $X2=0
+ $Y2=0
cc_217 N_A_284_31#_c_211_p N_VPWR_c_493_n 0.00467785f $X=1.935 $Y=2.58 $X2=0
+ $Y2=0
cc_218 N_A_284_31#_c_197_n N_VPWR_c_493_n 0.0232048f $X=4.43 $Y=2.58 $X2=0 $Y2=0
cc_219 N_A_284_31#_c_194_n N_X_M1003_s 0.00750686f $X=4.095 $Y=2.58 $X2=0 $Y2=0
cc_220 N_A_284_31#_c_183_n N_X_c_539_n 0.00108567f $X=1.855 $Y=0.78 $X2=0 $Y2=0
cc_221 N_A_284_31#_c_194_n X 0.0324736f $X=4.095 $Y=2.58 $X2=0 $Y2=0
cc_222 N_A_284_31#_c_194_n A_794_409# 0.00376324f $X=4.095 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_284_31#_c_197_n A_794_409# 0.00666053f $X=4.43 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_224 N_A_284_31#_c_179_n N_VGND_c_570_n 0.0105659f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_225 N_A_284_31#_c_183_n N_VGND_c_570_n 0.00188065f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_226 N_A_284_31#_c_188_n N_VGND_c_571_n 0.0153904f $X=4.21 $Y=0.58 $X2=0 $Y2=0
cc_227 N_A_284_31#_c_188_n N_VGND_c_573_n 0.0153904f $X=4.21 $Y=0.58 $X2=0 $Y2=0
cc_228 N_A_284_31#_c_179_n N_VGND_c_574_n 0.00445056f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_229 N_A_284_31#_c_180_n N_VGND_c_574_n 4.57848e-19 $X=1.78 $Y=0.855 $X2=0
+ $Y2=0
cc_230 N_A_284_31#_c_183_n N_VGND_c_574_n 0.00502664f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_231 N_A_284_31#_c_188_n N_VGND_c_577_n 0.0143041f $X=4.21 $Y=0.58 $X2=0 $Y2=0
cc_232 N_A_284_31#_c_179_n N_VGND_c_579_n 0.00418511f $X=1.495 $Y=0.78 $X2=0
+ $Y2=0
cc_233 N_A_284_31#_c_180_n N_VGND_c_579_n 6.33118e-19 $X=1.78 $Y=0.855 $X2=0
+ $Y2=0
cc_234 N_A_284_31#_c_183_n N_VGND_c_579_n 0.00650918f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_235 N_A_284_31#_c_188_n N_VGND_c_579_n 0.011808f $X=4.21 $Y=0.58 $X2=0 $Y2=0
cc_236 N_A_63_57#_M1011_g N_A1_N_M1000_g 0.0188003f $X=3.205 $Y=0.58 $X2=0 $Y2=0
cc_237 N_A_63_57#_M1003_g N_A1_N_M1006_g 0.0361464f $X=3.155 $Y=2.545 $X2=0
+ $Y2=0
cc_238 N_A_63_57#_c_296_n N_A1_N_c_388_n 0.0188003f $X=3.205 $Y=1.065 $X2=0
+ $Y2=0
cc_239 N_A_63_57#_M1003_g A1_N 0.0105161f $X=3.155 $Y=2.545 $X2=0 $Y2=0
cc_240 N_A_63_57#_M1003_g N_A1_N_c_391_n 0.0188003f $X=3.155 $Y=2.545 $X2=0
+ $Y2=0
cc_241 N_A_63_57#_M1003_g N_VPWR_c_495_n 0.00477272f $X=3.155 $Y=2.545 $X2=0
+ $Y2=0
cc_242 N_A_63_57#_M1003_g N_VPWR_c_498_n 0.00648402f $X=3.155 $Y=2.545 $X2=0
+ $Y2=0
cc_243 N_A_63_57#_M1003_g N_VPWR_c_493_n 0.00955866f $X=3.155 $Y=2.545 $X2=0
+ $Y2=0
cc_244 N_A_63_57#_c_291_n N_X_c_538_n 0.00753966f $X=2.77 $Y=1.065 $X2=0 $Y2=0
cc_245 N_A_63_57#_M1010_g N_X_c_538_n 0.00649965f $X=2.845 $Y=0.58 $X2=0 $Y2=0
cc_246 N_A_63_57#_M1003_g N_X_c_538_n 0.013824f $X=3.155 $Y=2.545 $X2=0 $Y2=0
cc_247 N_A_63_57#_c_296_n N_X_c_538_n 0.00928512f $X=3.205 $Y=1.065 $X2=0 $Y2=0
cc_248 N_A_63_57#_c_300_n N_X_c_538_n 3.66942e-19 $X=2.07 $Y=0.495 $X2=0 $Y2=0
cc_249 N_A_63_57#_c_301_n N_X_c_538_n 0.0214462f $X=2.307 $Y=1.182 $X2=0 $Y2=0
cc_250 N_A_63_57#_c_302_n N_X_c_538_n 0.034746f $X=2.307 $Y=1.468 $X2=0 $Y2=0
cc_251 N_A_63_57#_c_306_n N_X_c_538_n 0.0163809f $X=2.28 $Y=2.185 $X2=0 $Y2=0
cc_252 N_A_63_57#_c_303_n N_X_c_538_n 0.00447843f $X=2.335 $Y=1.155 $X2=0 $Y2=0
cc_253 N_A_63_57#_c_291_n N_X_c_539_n 0.00752545f $X=2.77 $Y=1.065 $X2=0 $Y2=0
cc_254 N_A_63_57#_c_292_n N_X_c_539_n 2.53927e-19 $X=2.5 $Y=1.065 $X2=0 $Y2=0
cc_255 N_A_63_57#_M1010_g N_X_c_539_n 0.0107588f $X=2.845 $Y=0.58 $X2=0 $Y2=0
cc_256 N_A_63_57#_M1011_g N_X_c_539_n 0.00238321f $X=3.205 $Y=0.58 $X2=0 $Y2=0
cc_257 N_A_63_57#_c_300_n N_X_c_539_n 0.0313782f $X=2.07 $Y=0.495 $X2=0 $Y2=0
cc_258 N_A_63_57#_c_301_n N_X_c_539_n 0.00281209f $X=2.307 $Y=1.182 $X2=0 $Y2=0
cc_259 N_A_63_57#_M1003_g X 0.0263437f $X=3.155 $Y=2.545 $X2=0 $Y2=0
cc_260 N_A_63_57#_c_306_n X 0.0277307f $X=2.28 $Y=2.185 $X2=0 $Y2=0
cc_261 N_A_63_57#_c_297_n N_VGND_c_570_n 0.0118803f $X=0.46 $Y=0.495 $X2=0 $Y2=0
cc_262 N_A_63_57#_c_298_n N_VGND_c_570_n 0.0199879f $X=1.905 $Y=0.905 $X2=0
+ $Y2=0
cc_263 N_A_63_57#_c_300_n N_VGND_c_570_n 0.0125465f $X=2.07 $Y=0.495 $X2=0 $Y2=0
cc_264 N_A_63_57#_M1010_g N_VGND_c_571_n 0.00178084f $X=2.845 $Y=0.58 $X2=0
+ $Y2=0
cc_265 N_A_63_57#_M1011_g N_VGND_c_571_n 0.0126434f $X=3.205 $Y=0.58 $X2=0 $Y2=0
cc_266 N_A_63_57#_M1010_g N_VGND_c_574_n 0.00371957f $X=2.845 $Y=0.58 $X2=0
+ $Y2=0
cc_267 N_A_63_57#_M1011_g N_VGND_c_574_n 0.00383152f $X=3.205 $Y=0.58 $X2=0
+ $Y2=0
cc_268 N_A_63_57#_c_300_n N_VGND_c_574_n 0.0220321f $X=2.07 $Y=0.495 $X2=0 $Y2=0
cc_269 N_A_63_57#_c_297_n N_VGND_c_576_n 0.0220321f $X=0.46 $Y=0.495 $X2=0 $Y2=0
cc_270 N_A_63_57#_M1010_g N_VGND_c_579_n 0.00623738f $X=2.845 $Y=0.58 $X2=0
+ $Y2=0
cc_271 N_A_63_57#_M1011_g N_VGND_c_579_n 0.00756787f $X=3.205 $Y=0.58 $X2=0
+ $Y2=0
cc_272 N_A_63_57#_c_297_n N_VGND_c_579_n 0.0125808f $X=0.46 $Y=0.495 $X2=0 $Y2=0
cc_273 N_A_63_57#_c_298_n N_VGND_c_579_n 0.0301961f $X=1.905 $Y=0.905 $X2=0
+ $Y2=0
cc_274 N_A_63_57#_c_300_n N_VGND_c_579_n 0.0125808f $X=2.07 $Y=0.495 $X2=0 $Y2=0
cc_275 N_A_63_57#_c_301_n N_VGND_c_579_n 0.00200643f $X=2.307 $Y=1.182 $X2=0
+ $Y2=0
cc_276 N_A1_N_M1013_g N_A2_N_c_429_n 0.0112008f $X=3.995 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_277 A1_N N_A2_N_c_429_n 5.32904e-19 $X=3.515 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_278 N_A1_N_c_391_n N_A2_N_c_429_n 0.0504671f $X=3.725 $Y=1.345 $X2=-0.19
+ $Y2=-0.245
cc_279 N_A1_N_c_389_n N_A2_N_M1015_g 0.0429039f $X=3.765 $Y=1.85 $X2=0 $Y2=0
cc_280 N_A1_N_M1013_g N_A2_N_M1001_g 0.0196091f $X=3.995 $Y=0.58 $X2=0 $Y2=0
cc_281 A1_N N_VPWR_M1003_d 0.00412521f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_282 N_A1_N_M1006_g N_VPWR_c_495_n 0.00451729f $X=3.845 $Y=2.545 $X2=0 $Y2=0
cc_283 N_A1_N_M1006_g N_VPWR_c_499_n 0.00648402f $X=3.845 $Y=2.545 $X2=0 $Y2=0
cc_284 N_A1_N_M1006_g N_VPWR_c_493_n 0.00859277f $X=3.845 $Y=2.545 $X2=0 $Y2=0
cc_285 A1_N N_X_c_538_n 0.0234778f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_286 N_A1_N_M1006_g X 9.20641e-19 $X=3.845 $Y=2.545 $X2=0 $Y2=0
cc_287 A1_N X 0.0142796f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_288 N_A1_N_M1000_g N_VGND_c_571_n 0.012388f $X=3.635 $Y=0.58 $X2=0 $Y2=0
cc_289 N_A1_N_M1013_g N_VGND_c_571_n 0.00182089f $X=3.995 $Y=0.58 $X2=0 $Y2=0
cc_290 A1_N N_VGND_c_571_n 0.00511426f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_291 N_A1_N_M1000_g N_VGND_c_577_n 0.00383152f $X=3.635 $Y=0.58 $X2=0 $Y2=0
cc_292 N_A1_N_M1013_g N_VGND_c_577_n 0.00434272f $X=3.995 $Y=0.58 $X2=0 $Y2=0
cc_293 N_A1_N_M1000_g N_VGND_c_579_n 0.00756787f $X=3.635 $Y=0.58 $X2=0 $Y2=0
cc_294 N_A1_N_M1013_g N_VGND_c_579_n 0.00820615f $X=3.995 $Y=0.58 $X2=0 $Y2=0
cc_295 N_A2_N_M1015_g N_VPWR_c_499_n 0.00568409f $X=4.335 $Y=2.545 $X2=0 $Y2=0
cc_296 N_A2_N_M1015_g N_VPWR_c_493_n 0.00849632f $X=4.335 $Y=2.545 $X2=0 $Y2=0
cc_297 N_A2_N_M1001_g N_VGND_c_573_n 0.00182089f $X=4.425 $Y=0.58 $X2=0 $Y2=0
cc_298 N_A2_N_M1004_g N_VGND_c_573_n 0.0138626f $X=4.785 $Y=0.58 $X2=0 $Y2=0
cc_299 A2_N N_VGND_c_573_n 0.0197853f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_300 N_A2_N_M1001_g N_VGND_c_577_n 0.00434272f $X=4.425 $Y=0.58 $X2=0 $Y2=0
cc_301 N_A2_N_M1004_g N_VGND_c_577_n 0.00383152f $X=4.785 $Y=0.58 $X2=0 $Y2=0
cc_302 N_A2_N_M1001_g N_VGND_c_579_n 0.00820615f $X=4.425 $Y=0.58 $X2=0 $Y2=0
cc_303 N_A2_N_M1004_g N_VGND_c_579_n 0.00756787f $X=4.785 $Y=0.58 $X2=0 $Y2=0
cc_304 N_A_43_408#_c_462_n N_VPWR_M1008_d 0.00180746f $X=1.255 $Y=2.105
+ $X2=-0.19 $Y2=1.655
cc_305 N_A_43_408#_c_461_n N_VPWR_c_494_n 0.0454646f $X=0.36 $Y=2.895 $X2=0
+ $Y2=0
cc_306 N_A_43_408#_c_462_n N_VPWR_c_494_n 0.0163515f $X=1.255 $Y=2.105 $X2=0
+ $Y2=0
cc_307 N_A_43_408#_c_464_n N_VPWR_c_494_n 0.0454646f $X=1.42 $Y=2.895 $X2=0
+ $Y2=0
cc_308 N_A_43_408#_c_461_n N_VPWR_c_496_n 0.021393f $X=0.36 $Y=2.895 $X2=0 $Y2=0
cc_309 N_A_43_408#_c_464_n N_VPWR_c_498_n 0.021393f $X=1.42 $Y=2.895 $X2=0 $Y2=0
cc_310 N_A_43_408#_c_461_n N_VPWR_c_493_n 0.0125495f $X=0.36 $Y=2.895 $X2=0
+ $Y2=0
cc_311 N_A_43_408#_c_464_n N_VPWR_c_493_n 0.0125495f $X=1.42 $Y=2.895 $X2=0
+ $Y2=0
cc_312 N_X_c_539_n N_VGND_c_571_n 0.0173472f $X=2.63 $Y=0.58 $X2=0 $Y2=0
cc_313 N_X_c_539_n N_VGND_c_574_n 0.0165886f $X=2.63 $Y=0.58 $X2=0 $Y2=0
cc_314 N_X_c_539_n N_VGND_c_579_n 0.0136626f $X=2.63 $Y=0.58 $X2=0 $Y2=0
