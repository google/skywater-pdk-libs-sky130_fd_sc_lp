* File: sky130_fd_sc_lp__a311oi_0.pxi.spice
* Created: Fri Aug 28 09:58:07 2020
* 
x_PM_SKY130_FD_SC_LP__A311OI_0%A3 N_A3_c_80_n N_A3_M1000_g N_A3_c_73_n
+ N_A3_M1006_g N_A3_c_74_n N_A3_c_75_n N_A3_c_76_n N_A3_c_77_n N_A3_c_83_n A3 A3
+ A3 N_A3_c_79_n PM_SKY130_FD_SC_LP__A311OI_0%A3
x_PM_SKY130_FD_SC_LP__A311OI_0%A2 N_A2_M1005_g N_A2_M1007_g N_A2_c_117_n
+ N_A2_c_121_n A2 A2 A2 A2 N_A2_c_119_n PM_SKY130_FD_SC_LP__A311OI_0%A2
x_PM_SKY130_FD_SC_LP__A311OI_0%A1 N_A1_M1003_g N_A1_M1001_g N_A1_c_166_n
+ N_A1_c_170_n A1 A1 N_A1_c_168_n PM_SKY130_FD_SC_LP__A311OI_0%A1
x_PM_SKY130_FD_SC_LP__A311OI_0%B1 N_B1_M1009_g N_B1_c_206_n N_B1_M1002_g
+ N_B1_c_207_n N_B1_c_208_n N_B1_c_209_n B1 B1 B1 B1 N_B1_c_211_n N_B1_c_212_n
+ B1 PM_SKY130_FD_SC_LP__A311OI_0%B1
x_PM_SKY130_FD_SC_LP__A311OI_0%C1 N_C1_M1008_g N_C1_c_268_n N_C1_M1004_g C1 C1
+ C1 N_C1_c_266_n PM_SKY130_FD_SC_LP__A311OI_0%C1
x_PM_SKY130_FD_SC_LP__A311OI_0%VPWR N_VPWR_M1000_s N_VPWR_M1005_d N_VPWR_c_301_n
+ N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n
+ VPWR N_VPWR_c_307_n N_VPWR_c_300_n PM_SKY130_FD_SC_LP__A311OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A311OI_0%A_158_473# N_A_158_473#_M1000_d
+ N_A_158_473#_M1001_d N_A_158_473#_c_337_n N_A_158_473#_c_338_n
+ N_A_158_473#_c_339_n N_A_158_473#_c_340_n
+ PM_SKY130_FD_SC_LP__A311OI_0%A_158_473#
x_PM_SKY130_FD_SC_LP__A311OI_0%Y N_Y_M1003_d N_Y_M1004_d N_Y_M1008_d N_Y_c_369_n
+ N_Y_c_370_n N_Y_c_371_n Y Y Y Y Y Y N_Y_c_373_n Y N_Y_c_376_n
+ PM_SKY130_FD_SC_LP__A311OI_0%Y
x_PM_SKY130_FD_SC_LP__A311OI_0%VGND N_VGND_M1006_s N_VGND_M1009_d N_VGND_c_416_n
+ VGND N_VGND_c_417_n N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n
+ PM_SKY130_FD_SC_LP__A311OI_0%VGND
cc_1 VNB N_A3_c_73_n 0.0207672f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=0.765
cc_2 VNB N_A3_c_74_n 0.0102254f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.08
cc_3 VNB N_A3_c_75_n 0.0330084f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.585
cc_4 VNB N_A3_c_76_n 0.00683607f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.75
cc_5 VNB N_A3_c_77_n 0.0256971f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=0.84
cc_6 VNB A3 0.0168178f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_7 VNB N_A3_c_79_n 0.0220367f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.245
cc_8 VNB N_A2_M1007_g 0.0299817f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.685
cc_9 VNB N_A2_c_117_n 0.021023f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=0.445
cc_10 VNB A2 0.0109275f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.08
cc_11 VNB N_A2_c_119_n 0.0176554f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.14
cc_12 VNB N_A1_M1003_g 0.0358685f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.75
cc_13 VNB N_A1_c_166_n 0.0206298f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=0.445
cc_14 VNB A1 0.00522051f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.08
cc_15 VNB N_A1_c_168_n 0.0153291f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=0.84
cc_16 VNB N_B1_c_206_n 0.0196277f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.685
cc_17 VNB N_B1_c_207_n 0.0189755f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.245
cc_18 VNB N_B1_c_208_n 0.0177555f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.08
cc_19 VNB N_B1_c_209_n 0.00715825f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.585
cc_20 VNB B1 0.00502275f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.75
cc_21 VNB N_B1_c_211_n 0.0194892f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_B1_c_212_n 0.0113361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_M1004_g 0.064698f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=0.765
cc_24 VNB C1 0.00856794f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.75
cc_25 VNB N_C1_c_266_n 0.0217755f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.14
cc_26 VNB N_VPWR_c_300_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_369_n 7.61769e-19 $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.245
cc_28 VNB N_Y_c_370_n 0.0130218f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.585
cc_29 VNB N_Y_c_371_n 0.00553875f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.75
cc_30 VNB Y 0.0119098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_373_n 0.0223403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Y 0.0389375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_416_n 0.0391629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_417_n 0.0192503f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.08
cc_35 VNB N_VGND_c_418_n 0.18884f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.585
cc_36 VNB N_VGND_c_419_n 0.0339997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_420_n 0.0185716f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.245
cc_38 VPB N_A3_c_80_n 0.0243779f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.065
cc_39 VPB N_A3_M1000_g 0.024699f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.685
cc_40 VPB N_A3_c_76_n 0.0149595f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.75
cc_41 VPB N_A3_c_83_n 0.0198997f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.14
cc_42 VPB A3 0.00782849f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_43 VPB N_A2_M1005_g 0.039607f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.75
cc_44 VPB N_A2_c_121_n 0.0153267f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.245
cc_45 VPB A2 0.00248914f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.08
cc_46 VPB N_A1_M1001_g 0.0405956f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.685
cc_47 VPB N_A1_c_170_n 0.0152651f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.245
cc_48 VPB A1 0.00278257f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.08
cc_49 VPB N_B1_M1002_g 0.042182f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=0.445
cc_50 VPB N_B1_c_209_n 0.0140127f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.585
cc_51 VPB B1 2.39217e-19 $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.75
cc_52 VPB B1 0.002735f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.84
cc_53 VPB B1 0.00364093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_C1_M1008_g 0.0279067f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.75
cc_55 VPB N_C1_c_268_n 0.0649545f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.685
cc_56 VPB C1 0.00567879f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.75
cc_57 VPB N_C1_c_266_n 3.74584e-19 $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.14
cc_58 VPB N_VPWR_c_301_n 0.0388455f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=0.765
cc_59 VPB N_VPWR_c_302_n 0.00980637f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.08
cc_60 VPB N_VPWR_c_303_n 0.0128037f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.84
cc_61 VPB N_VPWR_c_304_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_305_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_306_n 0.00516749f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.14
cc_64 VPB N_VPWR_c_307_n 0.051682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_300_n 0.0738011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_158_473#_c_337_n 0.00638732f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=0.765
cc_67 VPB N_A_158_473#_c_338_n 0.0157105f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=0.445
cc_68 VPB N_A_158_473#_c_339_n 0.00768119f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.245
cc_69 VPB N_A_158_473#_c_340_n 0.00528328f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.75
cc_70 VPB Y 0.0368714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_Y_c_376_n 0.0517483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 N_A3_c_80_n N_A2_M1005_g 0.00837221f $X=0.615 $Y=2.065 $X2=0 $Y2=0
cc_73 N_A3_c_83_n N_A2_M1005_g 0.0168753f $X=0.715 $Y=2.14 $X2=0 $Y2=0
cc_74 A3 N_A2_M1005_g 2.3298e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_75 N_A3_c_73_n N_A2_M1007_g 0.0496031f $X=0.825 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A3_c_74_n N_A2_M1007_g 0.00612985f $X=0.525 $Y=1.08 $X2=0 $Y2=0
cc_77 A3 N_A2_M1007_g 8.85689e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A3_c_75_n N_A2_c_117_n 0.0115875f $X=0.525 $Y=1.585 $X2=0 $Y2=0
cc_79 N_A3_c_76_n N_A2_c_121_n 0.0115875f $X=0.525 $Y=1.75 $X2=0 $Y2=0
cc_80 N_A3_c_73_n A2 0.00636537f $X=0.825 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A3_c_74_n A2 6.47233e-19 $X=0.525 $Y=1.08 $X2=0 $Y2=0
cc_82 A3 A2 0.0843905f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_83 N_A3_c_79_n A2 5.70401e-19 $X=0.525 $Y=1.245 $X2=0 $Y2=0
cc_84 A3 N_A2_c_119_n 0.00483511f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_85 N_A3_c_79_n N_A2_c_119_n 0.0115875f $X=0.525 $Y=1.245 $X2=0 $Y2=0
cc_86 N_A3_M1000_g N_VPWR_c_301_n 0.00382124f $X=0.715 $Y=2.685 $X2=0 $Y2=0
cc_87 N_A3_c_76_n N_VPWR_c_301_n 0.00304217f $X=0.525 $Y=1.75 $X2=0 $Y2=0
cc_88 N_A3_c_83_n N_VPWR_c_301_n 0.00298966f $X=0.715 $Y=2.14 $X2=0 $Y2=0
cc_89 A3 N_VPWR_c_301_n 0.00764735f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A3_M1000_g N_VPWR_c_305_n 0.00499542f $X=0.715 $Y=2.685 $X2=0 $Y2=0
cc_91 N_A3_M1000_g N_VPWR_c_300_n 0.0101368f $X=0.715 $Y=2.685 $X2=0 $Y2=0
cc_92 N_A3_c_83_n N_A_158_473#_c_337_n 0.00516196f $X=0.715 $Y=2.14 $X2=0 $Y2=0
cc_93 N_A3_c_80_n N_A_158_473#_c_339_n 0.00183931f $X=0.615 $Y=2.065 $X2=0 $Y2=0
cc_94 N_A3_c_83_n N_A_158_473#_c_339_n 0.00374343f $X=0.715 $Y=2.14 $X2=0 $Y2=0
cc_95 A3 N_A_158_473#_c_339_n 0.00365421f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A3_c_73_n N_VGND_c_416_n 0.0125489f $X=0.825 $Y=0.765 $X2=0 $Y2=0
cc_97 N_A3_c_77_n N_VGND_c_416_n 0.00519378f $X=0.825 $Y=0.84 $X2=0 $Y2=0
cc_98 A3 N_VGND_c_416_n 0.0261182f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_99 N_A3_c_79_n N_VGND_c_416_n 0.00322843f $X=0.525 $Y=1.245 $X2=0 $Y2=0
cc_100 N_A3_c_73_n N_VGND_c_418_n 0.00617572f $X=0.825 $Y=0.765 $X2=0 $Y2=0
cc_101 A3 N_VGND_c_418_n 0.00340638f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 N_A3_c_73_n N_VGND_c_419_n 0.00292692f $X=0.825 $Y=0.765 $X2=0 $Y2=0
cc_103 N_A2_M1007_g N_A1_M1003_g 0.0262613f $X=1.185 $Y=0.445 $X2=0 $Y2=0
cc_104 A2 N_A1_M1003_g 0.0109607f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A2_M1005_g N_A1_M1001_g 0.0296933f $X=1.145 $Y=2.685 $X2=0 $Y2=0
cc_106 N_A2_c_117_n N_A1_c_166_n 0.0262613f $X=1.095 $Y=1.66 $X2=0 $Y2=0
cc_107 N_A2_c_121_n N_A1_c_170_n 0.0262613f $X=1.095 $Y=1.825 $X2=0 $Y2=0
cc_108 A2 A1 0.0526746f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_109 N_A2_c_119_n A1 7.28384e-19 $X=1.095 $Y=1.32 $X2=0 $Y2=0
cc_110 N_A2_c_119_n N_A1_c_168_n 0.0262613f $X=1.095 $Y=1.32 $X2=0 $Y2=0
cc_111 A2 B1 0.00249568f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A2_M1005_g N_VPWR_c_302_n 0.00180033f $X=1.145 $Y=2.685 $X2=0 $Y2=0
cc_113 N_A2_M1005_g N_VPWR_c_305_n 0.00499542f $X=1.145 $Y=2.685 $X2=0 $Y2=0
cc_114 N_A2_M1005_g N_VPWR_c_300_n 0.00972572f $X=1.145 $Y=2.685 $X2=0 $Y2=0
cc_115 N_A2_M1005_g N_A_158_473#_c_337_n 0.00277344f $X=1.145 $Y=2.685 $X2=0
+ $Y2=0
cc_116 N_A2_M1005_g N_A_158_473#_c_338_n 0.014865f $X=1.145 $Y=2.685 $X2=0 $Y2=0
cc_117 N_A2_c_121_n N_A_158_473#_c_338_n 3.4139e-19 $X=1.095 $Y=1.825 $X2=0
+ $Y2=0
cc_118 A2 N_A_158_473#_c_338_n 0.0190805f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A2_c_121_n N_A_158_473#_c_339_n 0.00422643f $X=1.095 $Y=1.825 $X2=0
+ $Y2=0
cc_120 A2 N_A_158_473#_c_339_n 0.00418278f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A2_M1007_g N_Y_c_369_n 9.26281e-19 $X=1.185 $Y=0.445 $X2=0 $Y2=0
cc_122 A2 N_Y_c_369_n 0.0106859f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_123 A2 N_Y_c_371_n 0.00974696f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_124 N_A2_M1007_g N_VGND_c_416_n 0.00220693f $X=1.185 $Y=0.445 $X2=0 $Y2=0
cc_125 A2 N_VGND_c_416_n 0.0133785f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_126 N_A2_M1007_g N_VGND_c_418_n 0.00520479f $X=1.185 $Y=0.445 $X2=0 $Y2=0
cc_127 A2 N_VGND_c_418_n 0.010109f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A2_M1007_g N_VGND_c_419_n 0.00386151f $X=1.185 $Y=0.445 $X2=0 $Y2=0
cc_129 A2 N_VGND_c_419_n 0.00880201f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_130 A2 A_180_47# 0.00308008f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_131 N_A1_c_166_n N_B1_c_206_n 0.0144408f $X=1.635 $Y=1.66 $X2=0 $Y2=0
cc_132 N_A1_M1001_g N_B1_M1002_g 0.0278464f $X=1.575 $Y=2.685 $X2=0 $Y2=0
cc_133 N_A1_M1003_g N_B1_c_207_n 0.016967f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A1_c_170_n N_B1_c_209_n 0.0144408f $X=1.635 $Y=1.825 $X2=0 $Y2=0
cc_135 N_A1_M1003_g B1 7.13989e-19 $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_136 A1 B1 0.0557917f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A1_c_168_n B1 0.00104926f $X=1.635 $Y=1.32 $X2=0 $Y2=0
cc_138 N_A1_M1001_g B1 6.93262e-19 $X=1.575 $Y=2.685 $X2=0 $Y2=0
cc_139 N_A1_c_166_n B1 0.00104926f $X=1.635 $Y=1.66 $X2=0 $Y2=0
cc_140 N_A1_M1001_g B1 0.00105206f $X=1.575 $Y=2.685 $X2=0 $Y2=0
cc_141 A1 N_B1_c_211_n 0.00210778f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A1_c_168_n N_B1_c_211_n 0.0144408f $X=1.635 $Y=1.32 $X2=0 $Y2=0
cc_143 N_A1_M1003_g N_B1_c_212_n 0.00764376f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A1_M1001_g N_VPWR_c_302_n 0.00317497f $X=1.575 $Y=2.685 $X2=0 $Y2=0
cc_145 N_A1_M1001_g N_VPWR_c_307_n 0.00498026f $X=1.575 $Y=2.685 $X2=0 $Y2=0
cc_146 N_A1_M1001_g N_VPWR_c_300_n 0.00977287f $X=1.575 $Y=2.685 $X2=0 $Y2=0
cc_147 N_A1_M1001_g N_A_158_473#_c_338_n 0.0149555f $X=1.575 $Y=2.685 $X2=0
+ $Y2=0
cc_148 N_A1_c_170_n N_A_158_473#_c_338_n 0.00189898f $X=1.635 $Y=1.825 $X2=0
+ $Y2=0
cc_149 A1 N_A_158_473#_c_338_n 0.0262525f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A1_M1001_g N_A_158_473#_c_340_n 0.00288959f $X=1.575 $Y=2.685 $X2=0
+ $Y2=0
cc_151 N_A1_M1003_g N_Y_c_369_n 0.00748948f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_152 N_A1_M1003_g N_Y_c_371_n 0.0047158f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_153 A1 N_Y_c_371_n 0.0147971f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A1_c_168_n N_Y_c_371_n 0.0013258f $X=1.635 $Y=1.32 $X2=0 $Y2=0
cc_155 N_A1_M1003_g N_VGND_c_418_n 0.010028f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A1_M1003_g N_VGND_c_419_n 0.0054978f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_157 N_B1_M1002_g N_C1_c_268_n 0.0742794f $X=2.085 $Y=2.685 $X2=0 $Y2=0
cc_158 N_B1_c_209_n N_C1_c_268_n 0.0109571f $X=2.205 $Y=1.745 $X2=0 $Y2=0
cc_159 B1 N_C1_c_268_n 8.15594e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_160 B1 N_C1_c_268_n 0.00675938f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_161 N_B1_c_207_n N_C1_M1004_g 0.00618139f $X=2.075 $Y=0.765 $X2=0 $Y2=0
cc_162 N_B1_c_208_n N_C1_M1004_g 0.00831307f $X=2.075 $Y=0.915 $X2=0 $Y2=0
cc_163 B1 N_C1_M1004_g 5.63258e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_164 N_B1_c_211_n N_C1_M1004_g 0.0153281f $X=2.235 $Y=1.24 $X2=0 $Y2=0
cc_165 N_B1_M1002_g C1 8.17721e-19 $X=2.085 $Y=2.685 $X2=0 $Y2=0
cc_166 B1 C1 0.083736f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_167 N_B1_c_211_n C1 0.00467677f $X=2.235 $Y=1.24 $X2=0 $Y2=0
cc_168 N_B1_c_206_n N_C1_c_266_n 0.00874777f $X=2.205 $Y=1.55 $X2=0 $Y2=0
cc_169 N_B1_M1002_g N_VPWR_c_307_n 0.00412169f $X=2.085 $Y=2.685 $X2=0 $Y2=0
cc_170 B1 N_VPWR_c_307_n 0.00383984f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_171 N_B1_M1002_g N_VPWR_c_300_n 0.00687092f $X=2.085 $Y=2.685 $X2=0 $Y2=0
cc_172 B1 N_VPWR_c_300_n 0.00699727f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_173 N_B1_M1002_g N_A_158_473#_c_338_n 0.00136906f $X=2.085 $Y=2.685 $X2=0
+ $Y2=0
cc_174 B1 N_A_158_473#_c_338_n 0.0140872f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_175 N_B1_M1002_g N_A_158_473#_c_340_n 0.00803822f $X=2.085 $Y=2.685 $X2=0
+ $Y2=0
cc_176 B1 N_A_158_473#_c_340_n 0.0360869f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_177 B1 A_432_473# 0.00182346f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_178 N_B1_c_207_n N_Y_c_369_n 0.00235045f $X=2.075 $Y=0.765 $X2=0 $Y2=0
cc_179 N_B1_c_207_n N_Y_c_370_n 0.00495811f $X=2.075 $Y=0.765 $X2=0 $Y2=0
cc_180 N_B1_c_208_n N_Y_c_370_n 0.0152105f $X=2.075 $Y=0.915 $X2=0 $Y2=0
cc_181 B1 N_Y_c_370_n 0.0254415f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_B1_c_211_n N_Y_c_370_n 0.00401956f $X=2.235 $Y=1.24 $X2=0 $Y2=0
cc_183 N_B1_M1002_g N_Y_c_376_n 0.00130303f $X=2.085 $Y=2.685 $X2=0 $Y2=0
cc_184 B1 N_Y_c_376_n 0.0136295f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_185 N_B1_c_207_n N_VGND_c_418_n 0.00669395f $X=2.075 $Y=0.765 $X2=0 $Y2=0
cc_186 N_B1_c_207_n N_VGND_c_419_n 0.00322084f $X=2.075 $Y=0.765 $X2=0 $Y2=0
cc_187 N_B1_c_207_n N_VGND_c_420_n 0.00386763f $X=2.075 $Y=0.765 $X2=0 $Y2=0
cc_188 N_B1_c_208_n N_VGND_c_420_n 7.96729e-19 $X=2.075 $Y=0.915 $X2=0 $Y2=0
cc_189 N_C1_M1008_g N_VPWR_c_307_n 0.00468046f $X=2.445 $Y=2.685 $X2=0 $Y2=0
cc_190 N_C1_M1008_g N_VPWR_c_300_n 0.00942216f $X=2.445 $Y=2.685 $X2=0 $Y2=0
cc_191 N_C1_M1004_g N_Y_c_370_n 0.015198f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_192 C1 N_Y_c_370_n 0.0239332f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_193 N_C1_c_266_n N_Y_c_370_n 3.23136e-19 $X=2.775 $Y=1.63 $X2=0 $Y2=0
cc_194 N_C1_c_266_n Y 0.00443407f $X=2.775 $Y=1.63 $X2=0 $Y2=0
cc_195 N_C1_M1004_g N_Y_c_373_n 0.00391786f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_196 N_C1_M1008_g Y 0.00439775f $X=2.445 $Y=2.685 $X2=0 $Y2=0
cc_197 N_C1_M1004_g Y 0.0103281f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_198 C1 Y 0.0829584f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_199 N_C1_c_266_n Y 0.0189175f $X=2.775 $Y=1.63 $X2=0 $Y2=0
cc_200 N_C1_M1008_g N_Y_c_376_n 0.0112563f $X=2.445 $Y=2.685 $X2=0 $Y2=0
cc_201 N_C1_c_268_n N_Y_c_376_n 0.00881107f $X=2.805 $Y=1.985 $X2=0 $Y2=0
cc_202 C1 N_Y_c_376_n 0.0337241f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_203 N_C1_M1004_g N_VGND_c_417_n 0.00439206f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_204 N_C1_M1004_g N_VGND_c_418_n 0.00770382f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_205 N_C1_M1004_g N_VGND_c_420_n 0.00382939f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_206 N_VPWR_c_301_n N_A_158_473#_c_337_n 0.00226893f $X=0.5 $Y=2.52 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_302_n N_A_158_473#_c_337_n 0.00305856f $X=1.36 $Y=2.51 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_305_n N_A_158_473#_c_337_n 0.0140356f $X=1.23 $Y=3.33 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_300_n N_A_158_473#_c_337_n 0.00977851f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_302_n N_A_158_473#_c_338_n 0.0226354f $X=1.36 $Y=2.51 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_302_n N_A_158_473#_c_340_n 0.0288554f $X=1.36 $Y=2.51 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_307_n N_A_158_473#_c_340_n 0.0121316f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_300_n N_A_158_473#_c_340_n 0.00845197f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_307_n N_Y_c_376_n 0.0421119f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_215 N_VPWR_c_300_n N_Y_c_376_n 0.02942f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_216 N_A_158_473#_c_340_n N_Y_c_376_n 0.0107427f $X=1.79 $Y=2.51 $X2=0 $Y2=0
cc_217 N_Y_c_370_n N_VGND_c_417_n 0.00224537f $X=2.855 $Y=0.82 $X2=0 $Y2=0
cc_218 N_Y_c_373_n N_VGND_c_417_n 0.0239678f $X=2.99 $Y=0.445 $X2=0 $Y2=0
cc_219 N_Y_M1003_d N_VGND_c_418_n 0.00254596f $X=1.62 $Y=0.235 $X2=0 $Y2=0
cc_220 N_Y_M1004_d N_VGND_c_418_n 0.00218596f $X=2.85 $Y=0.235 $X2=0 $Y2=0
cc_221 N_Y_c_369_n N_VGND_c_418_n 0.012253f $X=1.775 $Y=0.445 $X2=0 $Y2=0
cc_222 N_Y_c_370_n N_VGND_c_418_n 0.0100926f $X=2.855 $Y=0.82 $X2=0 $Y2=0
cc_223 N_Y_c_373_n N_VGND_c_418_n 0.0160374f $X=2.99 $Y=0.445 $X2=0 $Y2=0
cc_224 N_Y_c_369_n N_VGND_c_419_n 0.0163523f $X=1.775 $Y=0.445 $X2=0 $Y2=0
cc_225 N_Y_c_370_n N_VGND_c_419_n 0.00158057f $X=2.855 $Y=0.82 $X2=0 $Y2=0
cc_226 N_Y_c_370_n N_VGND_c_420_n 0.0432076f $X=2.855 $Y=0.82 $X2=0 $Y2=0
cc_227 N_VGND_c_418_n A_180_47# 0.00562002f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_228 N_VGND_c_418_n A_252_47# 0.00715371f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
