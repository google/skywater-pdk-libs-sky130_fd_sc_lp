* File: sky130_fd_sc_lp__a31oi_m.spice
* Created: Fri Aug 28 10:00:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a31oi_m  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1006 A_189_82# N_A3_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1004 A_261_82# N_A2_M1004_g A_189_82# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A1_M1005_g A_261_82# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=0.99 PS=0.63 NRD=77.136 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75000.9
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1197 PD=1.37 PS=0.99 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_169_500#_M1007_d N_A3_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_169_500#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_A_169_500#_M1000_d N_A1_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_169_500#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
c_31 VNB 0 1.64292e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a31oi_m.pxi.spice"
*
.ends
*
*
