* File: sky130_fd_sc_lp__nor3_4.pxi.spice
* Created: Wed Sep  2 10:09:11 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3_4%A N_A_c_90_n N_A_M1001_g N_A_M1006_g N_A_c_92_n
+ N_A_M1009_g N_A_M1010_g N_A_c_94_n N_A_M1017_g N_A_M1018_g N_A_c_96_n
+ N_A_M1019_g N_A_M1020_g A A A A N_A_c_99_n PM_SKY130_FD_SC_LP__NOR3_4%A
x_PM_SKY130_FD_SC_LP__NOR3_4%B N_B_c_163_n N_B_M1008_g N_B_M1000_g N_B_c_165_n
+ N_B_M1015_g N_B_M1002_g N_B_c_167_n N_B_M1022_g N_B_M1003_g N_B_M1023_g
+ N_B_M1016_g N_B_c_170_n N_B_c_171_n N_B_c_172_n B B B N_B_c_174_n N_B_c_175_n
+ N_B_c_176_n PM_SKY130_FD_SC_LP__NOR3_4%B
x_PM_SKY130_FD_SC_LP__NOR3_4%C N_C_M1005_g N_C_M1004_g N_C_M1007_g N_C_M1011_g
+ N_C_M1012_g N_C_M1013_g N_C_M1014_g N_C_M1021_g N_C_c_311_n C C N_C_c_292_n
+ N_C_c_293_n C N_C_c_300_n PM_SKY130_FD_SC_LP__NOR3_4%C
x_PM_SKY130_FD_SC_LP__NOR3_4%A_29_367# N_A_29_367#_M1006_d N_A_29_367#_M1010_d
+ N_A_29_367#_M1020_d N_A_29_367#_M1002_s N_A_29_367#_M1016_s
+ N_A_29_367#_c_383_n N_A_29_367#_c_384_n N_A_29_367#_c_385_n
+ N_A_29_367#_c_430_p N_A_29_367#_c_386_n N_A_29_367#_c_431_p
+ N_A_29_367#_c_387_n N_A_29_367#_c_409_n N_A_29_367#_c_410_n
+ N_A_29_367#_c_412_n N_A_29_367#_c_388_n N_A_29_367#_c_389_n
+ N_A_29_367#_c_390_n N_A_29_367#_c_391_n PM_SKY130_FD_SC_LP__NOR3_4%A_29_367#
x_PM_SKY130_FD_SC_LP__NOR3_4%VPWR N_VPWR_M1006_s N_VPWR_M1018_s N_VPWR_c_461_n
+ N_VPWR_c_462_n VPWR N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n
+ N_VPWR_c_460_n N_VPWR_c_467_n N_VPWR_c_468_n PM_SKY130_FD_SC_LP__NOR3_4%VPWR
x_PM_SKY130_FD_SC_LP__NOR3_4%A_456_367# N_A_456_367#_M1000_d
+ N_A_456_367#_M1003_d N_A_456_367#_M1011_d N_A_456_367#_M1021_d
+ N_A_456_367#_c_528_n N_A_456_367#_c_530_n N_A_456_367#_c_533_n
+ PM_SKY130_FD_SC_LP__NOR3_4%A_456_367#
x_PM_SKY130_FD_SC_LP__NOR3_4%Y N_Y_M1001_s N_Y_M1017_s N_Y_M1008_d N_Y_M1022_d
+ N_Y_M1007_s N_Y_M1014_s N_Y_M1004_s N_Y_M1013_s N_Y_c_678_p N_Y_c_564_n
+ N_Y_c_568_n N_Y_c_672_p N_Y_c_570_n N_Y_c_673_p N_Y_c_577_n N_Y_c_581_n
+ N_Y_c_583_n N_Y_c_584_n N_Y_c_623_n N_Y_c_585_n N_Y_c_561_n N_Y_c_590_n
+ N_Y_c_559_n N_Y_c_560_n N_Y_c_572_n N_Y_c_598_n N_Y_c_600_n N_Y_c_602_n
+ N_Y_c_563_n N_Y_c_604_n Y N_Y_c_608_n Y N_Y_c_610_n
+ PM_SKY130_FD_SC_LP__NOR3_4%Y
x_PM_SKY130_FD_SC_LP__NOR3_4%VGND N_VGND_M1001_d N_VGND_M1009_d N_VGND_M1019_d
+ N_VGND_M1015_s N_VGND_M1005_d N_VGND_M1012_d N_VGND_M1023_s N_VGND_c_703_n
+ N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n N_VGND_c_708_n
+ N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n N_VGND_c_712_n N_VGND_c_713_n
+ N_VGND_c_714_n N_VGND_c_715_n N_VGND_c_716_n N_VGND_c_717_n VGND
+ N_VGND_c_718_n N_VGND_c_719_n N_VGND_c_720_n N_VGND_c_721_n N_VGND_c_722_n
+ N_VGND_c_723_n PM_SKY130_FD_SC_LP__NOR3_4%VGND
cc_1 VNB N_A_c_90_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.185
cc_2 VNB N_A_M1006_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_3 VNB N_A_c_92_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.185
cc_4 VNB N_A_M1010_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_5 VNB N_A_c_94_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.185
cc_6 VNB N_A_M1018_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.465
cc_7 VNB N_A_c_96_n 0.016201f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.185
cc_8 VNB N_A_M1020_g 0.00730538f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.465
cc_9 VNB A 0.0161101f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_10 VNB N_A_c_99_n 0.100541f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.35
cc_11 VNB N_B_c_163_n 0.016201f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.185
cc_12 VNB N_B_M1000_g 0.00730538f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_13 VNB N_B_c_165_n 0.0161751f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.185
cc_14 VNB N_B_M1002_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_15 VNB N_B_c_167_n 0.0157973f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.185
cc_16 VNB N_B_M1003_g 0.00728229f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.465
cc_17 VNB N_B_M1016_g 0.00804023f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.465
cc_18 VNB N_B_c_170_n 0.0273803f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_B_c_171_n 0.00248724f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_20 VNB N_B_c_172_n 0.0343045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB B 0.00393724f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.35
cc_22 VNB N_B_c_174_n 0.0540397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_175_n 0.0196625f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.362
cc_24 VNB N_B_c_176_n 0.00783686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C_M1005_g 0.0230925f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.655
cc_26 VNB N_C_M1007_g 0.0228834f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.515
cc_27 VNB N_C_M1012_g 0.0229013f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.465
cc_28 VNB N_C_M1014_g 0.0226582f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.465
cc_29 VNB N_C_c_292_n 0.0646467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_c_293_n 0.00238501f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.362
cc_31 VNB N_VPWR_c_460_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_559_n 0.0090884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_560_n 0.0342429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_703_n 0.0113208f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.185
cc_35 VNB N_VGND_c_704_n 0.0357294f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.655
cc_36 VNB N_VGND_c_705_n 3.14366e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_706_n 3.14366e-19 $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_38 VNB N_VGND_c_707_n 0.00383093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_708_n 0.003699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_709_n 0.003699f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=1.35
cc_41 VNB N_VGND_c_710_n 0.0121548f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=1.35
cc_42 VNB N_VGND_c_711_n 0.0168434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_712_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_713_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.362
cc_45 VNB N_VGND_c_714_n 0.0139823f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.362
cc_46 VNB N_VGND_c_715_n 0.00439335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_716_n 0.0166684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_717_n 0.00362088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_718_n 0.0146078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_719_n 0.0166684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_720_n 0.0166684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_721_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_722_n 0.00362088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_723_n 0.288211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_A_M1006_g 0.0246191f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_56 VPB N_A_M1010_g 0.0184959f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_57 VPB N_A_M1018_g 0.0184959f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=2.465
cc_58 VPB N_A_M1020_g 0.018645f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.465
cc_59 VPB N_B_M1000_g 0.0188441f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_60 VPB N_B_M1002_g 0.018695f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_61 VPB N_B_M1003_g 0.0195977f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=2.465
cc_62 VPB N_B_M1016_g 0.0237102f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.465
cc_63 VPB N_C_M1004_g 0.0181868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_C_M1011_g 0.0180109f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.185
cc_65 VPB N_C_M1013_g 0.0186072f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=0.655
cc_66 VPB N_C_M1021_g 0.0188097f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_67 VPB N_C_c_292_n 0.0118182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_C_c_293_n 0.00428453f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.362
cc_69 VPB N_C_c_300_n 0.00258364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_29_367#_c_383_n 0.0454116f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.515
cc_71 VPB N_A_29_367#_c_384_n 0.00304088f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.185
cc_72 VPB N_A_29_367#_c_385_n 0.00942555f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=0.655
cc_73 VPB N_A_29_367#_c_386_n 0.0035011f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_74 VPB N_A_29_367#_c_387_n 0.00514361f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.35
cc_75 VPB N_A_29_367#_c_388_n 0.0226976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_29_367#_c_389_n 0.00151965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_29_367#_c_390_n 0.00279443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_29_367#_c_391_n 0.0135273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_461_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.655
cc_80 VPB N_VPWR_c_462_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.185
cc_81 VPB N_VPWR_c_463_n 0.0156941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_464_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.465
cc_83 VPB N_VPWR_c_465_n 0.0968411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_460_n 0.0475628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_467_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.35
cc_86 VPB N_VPWR_c_468_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_Y_c_561_n 0.0184505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_Y_c_560_n 0.00800939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_Y_c_563_n 0.00226953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 N_A_c_96_n N_B_c_163_n 0.0247847f $X=1.775 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_91 N_A_M1020_g N_B_M1000_g 0.0247847f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_92 A B 0.0270138f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A_c_99_n B 0.00120533f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_94 A N_B_c_174_n 3.11896e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_95 N_A_c_99_n N_B_c_174_n 0.0247847f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_96 N_A_M1006_g N_A_29_367#_c_384_n 0.0150503f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_M1010_g N_A_29_367#_c_384_n 0.0139931f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_98 A N_A_29_367#_c_384_n 0.0448317f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A_c_99_n N_A_29_367#_c_384_n 0.00320667f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_100 A N_A_29_367#_c_385_n 0.020289f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A_c_99_n N_A_29_367#_c_385_n 0.00472787f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_102 N_A_M1018_g N_A_29_367#_c_386_n 0.0139931f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_M1020_g N_A_29_367#_c_386_n 0.0139577f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_104 A N_A_29_367#_c_386_n 0.0417745f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A_c_99_n N_A_29_367#_c_386_n 0.00221311f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_106 A N_A_29_367#_c_389_n 0.0146616f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A_c_99_n N_A_29_367#_c_389_n 0.00230628f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_108 N_A_M1006_g N_VPWR_c_461_n 0.016151f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_M1010_g N_VPWR_c_461_n 0.0141762f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_M1018_g N_VPWR_c_461_n 7.24342e-19 $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_M1010_g N_VPWR_c_462_n 7.24342e-19 $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_M1018_g N_VPWR_c_462_n 0.0141762f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_M1020_g N_VPWR_c_462_n 0.0153689f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_M1006_g N_VPWR_c_463_n 0.00486043f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_M1010_g N_VPWR_c_464_n 0.00486043f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_M1018_g N_VPWR_c_464_n 0.00486043f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_M1020_g N_VPWR_c_465_n 0.00486043f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_M1006_g N_VPWR_c_460_n 0.00918921f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_M1010_g N_VPWR_c_460_n 0.00824727f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_M1018_g N_VPWR_c_460_n 0.00824727f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_M1020_g N_VPWR_c_460_n 0.0082726f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_c_92_n N_Y_c_564_n 0.0122595f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_123 N_A_c_94_n N_Y_c_564_n 0.0122129f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_124 A N_Y_c_564_n 0.0409662f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A_c_99_n N_Y_c_564_n 0.00230884f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_126 A N_Y_c_568_n 0.0156448f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A_c_99_n N_Y_c_568_n 0.00240082f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_128 N_A_c_96_n N_Y_c_570_n 0.0122129f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_129 A N_Y_c_570_n 0.0122788f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 A N_Y_c_572_n 0.0145274f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A_c_99_n N_Y_c_572_n 0.00240082f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_132 N_A_c_90_n N_VGND_c_704_n 0.00554367f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_133 A N_VGND_c_704_n 0.022474f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A_c_99_n N_VGND_c_704_n 0.00569459f $X=1.775 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A_c_90_n N_VGND_c_705_n 5.88023e-19 $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_136 N_A_c_92_n N_VGND_c_705_n 0.0105794f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_137 N_A_c_94_n N_VGND_c_705_n 0.0105101f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A_c_96_n N_VGND_c_705_n 5.75816e-19 $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_139 N_A_c_94_n N_VGND_c_706_n 5.75816e-19 $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_140 N_A_c_96_n N_VGND_c_706_n 0.0104353f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A_c_94_n N_VGND_c_712_n 0.00486043f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_142 N_A_c_96_n N_VGND_c_712_n 0.00486043f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_143 N_A_c_90_n N_VGND_c_718_n 0.00585385f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_144 N_A_c_92_n N_VGND_c_718_n 0.00486043f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_145 N_A_c_90_n N_VGND_c_723_n 0.0114507f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_146 N_A_c_92_n N_VGND_c_723_n 0.00824727f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_147 N_A_c_94_n N_VGND_c_723_n 0.00824727f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_148 N_A_c_96_n N_VGND_c_723_n 0.00824727f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_149 N_B_c_167_n N_C_M1005_g 0.0299592f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_150 N_B_c_170_n N_C_M1005_g 0.0105063f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_151 N_B_c_176_n N_C_M1005_g 0.00480804f $X=3.25 $Y=1.295 $X2=0 $Y2=0
cc_152 N_B_M1003_g N_C_M1004_g 0.0299592f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_153 N_B_c_170_n N_C_M1007_g 0.0105529f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B_c_170_n N_C_M1012_g 0.0105063f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B_c_170_n N_C_M1014_g 0.0111764f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B_c_171_n N_C_M1014_g 0.00177586f $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B_c_172_n N_C_M1014_g 0.021852f $X=5.235 $Y=1.35 $X2=0 $Y2=0
cc_158 N_B_c_175_n N_C_M1014_g 0.0157557f $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_159 N_B_M1016_g N_C_c_311_n 6.6398e-19 $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B_c_171_n N_C_c_311_n 0.0049224f $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B_c_172_n N_C_c_311_n 3.00603e-19 $X=5.235 $Y=1.35 $X2=0 $Y2=0
cc_162 N_B_M1016_g N_C_c_292_n 0.0613657f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B_c_170_n N_C_c_292_n 0.00730626f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B_c_174_n N_C_c_292_n 0.0299592f $X=3.065 $Y=1.35 $X2=0 $Y2=0
cc_165 N_B_c_176_n N_C_c_292_n 3.89844e-19 $X=3.25 $Y=1.295 $X2=0 $Y2=0
cc_166 N_B_c_170_n N_C_c_293_n 0.0986812f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_167 N_B_c_174_n N_C_c_293_n 0.00149393f $X=3.065 $Y=1.35 $X2=0 $Y2=0
cc_168 N_B_c_176_n N_C_c_293_n 0.00873714f $X=3.25 $Y=1.295 $X2=0 $Y2=0
cc_169 N_B_M1000_g N_A_29_367#_c_387_n 0.0139104f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_170 N_B_M1002_g N_A_29_367#_c_387_n 0.0139459f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B_M1003_g N_A_29_367#_c_387_n 0.00503056f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_172 B N_A_29_367#_c_387_n 0.0649672f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_B_c_174_n N_A_29_367#_c_387_n 0.00451939f $X=3.065 $Y=1.35 $X2=0 $Y2=0
cc_174 N_B_M1003_g N_A_29_367#_c_409_n 0.00790018f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B_M1003_g N_A_29_367#_c_410_n 0.0111487f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_176 N_B_M1016_g N_A_29_367#_c_410_n 0.0111541f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_177 N_B_M1003_g N_A_29_367#_c_412_n 7.4145e-19 $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B_M1016_g N_A_29_367#_c_388_n 0.0065754f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_179 B N_A_29_367#_c_390_n 0.00528506f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_180 N_B_M1016_g N_A_29_367#_c_391_n 0.00342571f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B_M1000_g N_VPWR_c_462_n 0.00136666f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B_M1000_g N_VPWR_c_465_n 0.00547432f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B_M1002_g N_VPWR_c_465_n 0.00357842f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B_M1003_g N_VPWR_c_465_n 0.00357877f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B_M1016_g N_VPWR_c_465_n 0.00579312f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B_M1000_g N_VPWR_c_460_n 0.00990114f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_187 N_B_M1002_g N_VPWR_c_460_n 0.00535118f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B_M1003_g N_VPWR_c_460_n 0.00544922f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B_M1016_g N_VPWR_c_460_n 0.00739704f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B_M1000_g N_A_456_367#_c_528_n 0.0044463f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B_M1002_g N_A_456_367#_c_528_n 0.00129013f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_B_M1000_g N_A_456_367#_c_530_n 0.00677888f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_B_M1002_g N_A_456_367#_c_530_n 0.00822059f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_B_M1003_g N_A_456_367#_c_530_n 8.318e-19 $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_195 N_B_M1002_g N_A_456_367#_c_533_n 0.016523f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_196 N_B_M1003_g N_A_456_367#_c_533_n 0.0142675f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_197 N_B_c_171_n N_Y_M1014_s 7.71934e-19 $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B_c_163_n N_Y_c_570_n 0.0122129f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_199 B N_Y_c_570_n 0.0187291f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_200 N_B_c_167_n N_Y_c_577_n 0.00904331f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_201 B N_Y_c_577_n 0.00630165f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_202 N_B_c_174_n N_Y_c_577_n 7.26385e-19 $X=3.065 $Y=1.35 $X2=0 $Y2=0
cc_203 N_B_c_176_n N_Y_c_577_n 0.00555369f $X=3.25 $Y=1.295 $X2=0 $Y2=0
cc_204 N_B_c_165_n N_Y_c_581_n 5.27972e-19 $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_205 N_B_c_167_n N_Y_c_581_n 0.00628569f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_206 N_B_c_170_n N_Y_c_583_n 0.0320248f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_207 N_B_M1003_g N_Y_c_584_n 6.39431e-19 $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B_c_170_n N_Y_c_585_n 0.0320248f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_209 N_B_M1016_g N_Y_c_561_n 0.0135862f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B_c_170_n N_Y_c_561_n 0.00908185f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B_c_171_n N_Y_c_561_n 0.0124284f $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B_c_172_n N_Y_c_561_n 0.00299653f $X=5.235 $Y=1.35 $X2=0 $Y2=0
cc_213 N_B_c_175_n N_Y_c_590_n 0.0107173f $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_214 N_B_c_171_n N_Y_c_559_n 0.0103103f $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_215 N_B_c_172_n N_Y_c_559_n 0.00207146f $X=5.235 $Y=1.35 $X2=0 $Y2=0
cc_216 N_B_c_175_n N_Y_c_559_n 0.0104144f $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_217 N_B_M1016_g N_Y_c_560_n 0.00980518f $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B_c_171_n N_Y_c_560_n 0.032913f $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_219 N_B_c_172_n N_Y_c_560_n 0.00803689f $X=5.235 $Y=1.35 $X2=0 $Y2=0
cc_220 N_B_c_175_n N_Y_c_560_n 0.00658586f $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_221 B N_Y_c_598_n 0.0156448f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_222 N_B_c_174_n N_Y_c_598_n 0.00240082f $X=3.065 $Y=1.35 $X2=0 $Y2=0
cc_223 N_B_c_167_n N_Y_c_600_n 7.26734e-19 $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_224 N_B_c_176_n N_Y_c_600_n 0.0214902f $X=3.25 $Y=1.295 $X2=0 $Y2=0
cc_225 N_B_c_170_n N_Y_c_602_n 0.02078f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_226 N_B_M1016_g N_Y_c_563_n 9.1042e-19 $X=5.215 $Y=2.465 $X2=0 $Y2=0
cc_227 N_B_c_170_n N_Y_c_604_n 0.0159147f $X=5.07 $Y=1.16 $X2=0 $Y2=0
cc_228 N_B_c_171_n N_Y_c_604_n 0.00521351f $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_229 N_B_c_172_n N_Y_c_604_n 2.69864e-19 $X=5.235 $Y=1.35 $X2=0 $Y2=0
cc_230 N_B_c_175_n N_Y_c_604_n 7.25739e-19 $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_231 N_B_c_165_n N_Y_c_608_n 0.0100534f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_232 B N_Y_c_608_n 0.0212055f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_233 N_B_c_165_n N_Y_c_610_n 0.00316375f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_234 N_B_c_167_n N_Y_c_610_n 0.00418471f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_235 N_B_c_174_n N_Y_c_610_n 0.00152361f $X=3.065 $Y=1.35 $X2=0 $Y2=0
cc_236 N_B_c_171_n N_VGND_M1023_s 4.37347e-19 $X=5.2 $Y=1.16 $X2=0 $Y2=0
cc_237 N_B_c_163_n N_VGND_c_706_n 0.0105046f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_238 N_B_c_165_n N_VGND_c_706_n 5.88023e-19 $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_239 N_B_c_165_n N_VGND_c_707_n 0.001584f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_240 N_B_c_167_n N_VGND_c_707_n 0.00155791f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_241 N_B_c_175_n N_VGND_c_711_n 0.00327088f $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_242 N_B_c_163_n N_VGND_c_714_n 0.00486043f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_243 N_B_c_165_n N_VGND_c_714_n 0.00437852f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_244 N_B_c_167_n N_VGND_c_716_n 0.00426006f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_245 N_B_c_175_n N_VGND_c_720_n 0.00426006f $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_246 N_B_c_163_n N_VGND_c_723_n 0.00824727f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_247 N_B_c_165_n N_VGND_c_723_n 0.00583712f $X=2.635 $Y=1.185 $X2=0 $Y2=0
cc_248 N_B_c_167_n N_VGND_c_723_n 0.00583081f $X=3.065 $Y=1.185 $X2=0 $Y2=0
cc_249 N_B_c_175_n N_VGND_c_723_n 0.00682322f $X=5.235 $Y=1.185 $X2=0 $Y2=0
cc_250 N_C_M1004_g N_A_29_367#_c_387_n 5.99201e-19 $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_251 N_C_c_293_n N_A_29_367#_c_387_n 0.002467f $X=4.06 $Y=1.59 $X2=0 $Y2=0
cc_252 N_C_M1004_g N_A_29_367#_c_409_n 0.00177214f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_253 N_C_M1004_g N_A_29_367#_c_410_n 0.0120798f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_254 N_C_M1011_g N_A_29_367#_c_410_n 0.0105473f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_255 N_C_M1013_g N_A_29_367#_c_410_n 0.0105327f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_256 N_C_M1021_g N_A_29_367#_c_410_n 0.011272f $X=4.785 $Y=2.465 $X2=0 $Y2=0
cc_257 N_C_c_293_n N_A_29_367#_c_410_n 0.00336556f $X=4.06 $Y=1.59 $X2=0 $Y2=0
cc_258 N_C_M1021_g N_A_29_367#_c_391_n 0.00166413f $X=4.785 $Y=2.465 $X2=0 $Y2=0
cc_259 N_C_M1004_g N_VPWR_c_465_n 0.00357877f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_260 N_C_M1011_g N_VPWR_c_465_n 0.00357877f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_261 N_C_M1013_g N_VPWR_c_465_n 0.00357877f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_262 N_C_M1021_g N_VPWR_c_465_n 0.00357877f $X=4.785 $Y=2.465 $X2=0 $Y2=0
cc_263 N_C_M1004_g N_VPWR_c_460_n 0.00544922f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_264 N_C_M1011_g N_VPWR_c_460_n 0.00542194f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_265 N_C_M1013_g N_VPWR_c_460_n 0.00542194f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_266 N_C_M1021_g N_VPWR_c_460_n 0.00544922f $X=4.785 $Y=2.465 $X2=0 $Y2=0
cc_267 N_C_M1004_g N_A_456_367#_c_533_n 0.0142686f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_268 N_C_M1011_g N_A_456_367#_c_533_n 0.0142794f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_269 N_C_M1013_g N_A_456_367#_c_533_n 0.0141544f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_270 N_C_M1021_g N_A_456_367#_c_533_n 0.0141823f $X=4.785 $Y=2.465 $X2=0 $Y2=0
cc_271 N_C_M1005_g N_Y_c_581_n 0.00617717f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_272 N_C_M1007_g N_Y_c_581_n 5.19723e-19 $X=3.925 $Y=0.655 $X2=0 $Y2=0
cc_273 N_C_M1005_g N_Y_c_583_n 0.00885653f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_274 N_C_M1007_g N_Y_c_583_n 0.00885653f $X=3.925 $Y=0.655 $X2=0 $Y2=0
cc_275 N_C_M1004_g N_Y_c_584_n 0.00447929f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_276 N_C_M1011_g N_Y_c_584_n 0.00978764f $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_277 N_C_M1013_g N_Y_c_584_n 0.0103391f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_278 N_C_c_311_n N_Y_c_584_n 0.00679094f $X=4.605 $Y=1.51 $X2=0 $Y2=0
cc_279 N_C_c_292_n N_Y_c_584_n 0.00113868f $X=4.785 $Y=1.51 $X2=0 $Y2=0
cc_280 N_C_c_293_n N_Y_c_584_n 0.0468496f $X=4.06 $Y=1.59 $X2=0 $Y2=0
cc_281 N_C_M1005_g N_Y_c_623_n 5.19723e-19 $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_282 N_C_M1007_g N_Y_c_623_n 0.00617717f $X=3.925 $Y=0.655 $X2=0 $Y2=0
cc_283 N_C_M1012_g N_Y_c_623_n 0.00617717f $X=4.355 $Y=0.655 $X2=0 $Y2=0
cc_284 N_C_M1014_g N_Y_c_623_n 5.19723e-19 $X=4.785 $Y=0.655 $X2=0 $Y2=0
cc_285 N_C_M1012_g N_Y_c_585_n 0.00885653f $X=4.355 $Y=0.655 $X2=0 $Y2=0
cc_286 N_C_M1014_g N_Y_c_585_n 0.00885653f $X=4.785 $Y=0.655 $X2=0 $Y2=0
cc_287 N_C_M1021_g N_Y_c_561_n 0.0101437f $X=4.785 $Y=2.465 $X2=0 $Y2=0
cc_288 N_C_c_311_n N_Y_c_561_n 0.00242874f $X=4.605 $Y=1.51 $X2=0 $Y2=0
cc_289 N_C_M1012_g N_Y_c_590_n 5.19723e-19 $X=4.355 $Y=0.655 $X2=0 $Y2=0
cc_290 N_C_M1014_g N_Y_c_590_n 0.00617717f $X=4.785 $Y=0.655 $X2=0 $Y2=0
cc_291 N_C_M1005_g N_Y_c_600_n 7.26734e-19 $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_292 N_C_M1007_g N_Y_c_602_n 7.26734e-19 $X=3.925 $Y=0.655 $X2=0 $Y2=0
cc_293 N_C_M1012_g N_Y_c_602_n 7.26734e-19 $X=4.355 $Y=0.655 $X2=0 $Y2=0
cc_294 N_C_M1011_g N_Y_c_563_n 6.89398e-19 $X=3.925 $Y=2.465 $X2=0 $Y2=0
cc_295 N_C_M1013_g N_Y_c_563_n 0.00422108f $X=4.355 $Y=2.465 $X2=0 $Y2=0
cc_296 N_C_M1021_g N_Y_c_563_n 0.00488726f $X=4.785 $Y=2.465 $X2=0 $Y2=0
cc_297 N_C_c_311_n N_Y_c_563_n 0.0252874f $X=4.605 $Y=1.51 $X2=0 $Y2=0
cc_298 N_C_c_292_n N_Y_c_563_n 0.00236448f $X=4.785 $Y=1.51 $X2=0 $Y2=0
cc_299 N_C_M1014_g N_Y_c_604_n 7.26734e-19 $X=4.785 $Y=0.655 $X2=0 $Y2=0
cc_300 N_C_M1005_g N_VGND_c_708_n 0.00153274f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_301 N_C_M1007_g N_VGND_c_708_n 0.00153274f $X=3.925 $Y=0.655 $X2=0 $Y2=0
cc_302 N_C_M1012_g N_VGND_c_709_n 0.00153274f $X=4.355 $Y=0.655 $X2=0 $Y2=0
cc_303 N_C_M1014_g N_VGND_c_709_n 0.00153274f $X=4.785 $Y=0.655 $X2=0 $Y2=0
cc_304 N_C_M1005_g N_VGND_c_716_n 0.00426006f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_305 N_C_M1007_g N_VGND_c_719_n 0.00426006f $X=3.925 $Y=0.655 $X2=0 $Y2=0
cc_306 N_C_M1012_g N_VGND_c_719_n 0.00426006f $X=4.355 $Y=0.655 $X2=0 $Y2=0
cc_307 N_C_M1014_g N_VGND_c_720_n 0.00426006f $X=4.785 $Y=0.655 $X2=0 $Y2=0
cc_308 N_C_M1005_g N_VGND_c_723_n 0.00583081f $X=3.495 $Y=0.655 $X2=0 $Y2=0
cc_309 N_C_M1007_g N_VGND_c_723_n 0.00580548f $X=3.925 $Y=0.655 $X2=0 $Y2=0
cc_310 N_C_M1012_g N_VGND_c_723_n 0.00580548f $X=4.355 $Y=0.655 $X2=0 $Y2=0
cc_311 N_C_M1014_g N_VGND_c_723_n 0.00583081f $X=4.785 $Y=0.655 $X2=0 $Y2=0
cc_312 N_A_29_367#_c_384_n N_VPWR_M1006_s 0.00201607f $X=1.035 $Y=1.79 $X2=-0.19
+ $Y2=1.655
cc_313 N_A_29_367#_c_386_n N_VPWR_M1018_s 0.00201607f $X=1.895 $Y=1.79 $X2=0
+ $Y2=0
cc_314 N_A_29_367#_c_384_n N_VPWR_c_461_n 0.013593f $X=1.035 $Y=1.79 $X2=0 $Y2=0
cc_315 N_A_29_367#_c_386_n N_VPWR_c_462_n 0.013593f $X=1.895 $Y=1.79 $X2=0 $Y2=0
cc_316 N_A_29_367#_c_383_n N_VPWR_c_463_n 0.0178111f $X=0.27 $Y=1.98 $X2=0 $Y2=0
cc_317 N_A_29_367#_c_430_p N_VPWR_c_464_n 0.0124525f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_318 N_A_29_367#_c_431_p N_VPWR_c_465_n 0.0124525f $X=1.99 $Y=1.98 $X2=0 $Y2=0
cc_319 N_A_29_367#_c_388_n N_VPWR_c_465_n 0.0210895f $X=5.45 $Y=2.95 $X2=0 $Y2=0
cc_320 N_A_29_367#_M1006_d N_VPWR_c_460_n 0.00371702f $X=0.145 $Y=1.835 $X2=0
+ $Y2=0
cc_321 N_A_29_367#_M1010_d N_VPWR_c_460_n 0.00536646f $X=0.99 $Y=1.835 $X2=0
+ $Y2=0
cc_322 N_A_29_367#_M1020_d N_VPWR_c_460_n 0.00536646f $X=1.85 $Y=1.835 $X2=0
+ $Y2=0
cc_323 N_A_29_367#_M1002_s N_VPWR_c_460_n 0.00225186f $X=2.71 $Y=1.835 $X2=0
+ $Y2=0
cc_324 N_A_29_367#_M1016_s N_VPWR_c_460_n 0.00231914f $X=5.29 $Y=1.835 $X2=0
+ $Y2=0
cc_325 N_A_29_367#_c_383_n N_VPWR_c_460_n 0.0100304f $X=0.27 $Y=1.98 $X2=0 $Y2=0
cc_326 N_A_29_367#_c_430_p N_VPWR_c_460_n 0.00730901f $X=1.13 $Y=1.98 $X2=0
+ $Y2=0
cc_327 N_A_29_367#_c_431_p N_VPWR_c_460_n 0.00730901f $X=1.99 $Y=1.98 $X2=0
+ $Y2=0
cc_328 N_A_29_367#_c_410_n N_VPWR_c_460_n 0.00810645f $X=5.285 $Y=2.41 $X2=0
+ $Y2=0
cc_329 N_A_29_367#_c_388_n N_VPWR_c_460_n 0.0126604f $X=5.45 $Y=2.95 $X2=0 $Y2=0
cc_330 N_A_29_367#_c_387_n N_A_456_367#_M1000_d 0.00180746f $X=2.755 $Y=1.79
+ $X2=-0.19 $Y2=1.655
cc_331 N_A_29_367#_c_410_n N_A_456_367#_M1003_d 0.00811934f $X=5.285 $Y=2.41
+ $X2=0 $Y2=0
cc_332 N_A_29_367#_c_410_n N_A_456_367#_M1011_d 0.00347487f $X=5.285 $Y=2.41
+ $X2=0 $Y2=0
cc_333 N_A_29_367#_c_410_n N_A_456_367#_M1021_d 0.00423283f $X=5.285 $Y=2.41
+ $X2=0 $Y2=0
cc_334 N_A_29_367#_c_387_n N_A_456_367#_c_530_n 0.0163515f $X=2.755 $Y=1.79
+ $X2=0 $Y2=0
cc_335 N_A_29_367#_M1002_s N_A_456_367#_c_533_n 0.00345623f $X=2.71 $Y=1.835
+ $X2=0 $Y2=0
cc_336 N_A_29_367#_c_410_n N_A_456_367#_c_533_n 0.108609f $X=5.285 $Y=2.41 $X2=0
+ $Y2=0
cc_337 N_A_29_367#_c_412_n N_A_456_367#_c_533_n 0.0151462f $X=3.015 $Y=2.41
+ $X2=0 $Y2=0
cc_338 N_A_29_367#_c_410_n N_Y_M1004_s 0.00347487f $X=5.285 $Y=2.41 $X2=0 $Y2=0
cc_339 N_A_29_367#_c_410_n N_Y_M1013_s 0.00347088f $X=5.285 $Y=2.41 $X2=0 $Y2=0
cc_340 N_A_29_367#_c_390_n N_Y_c_570_n 0.00371455f $X=1.99 $Y=1.79 $X2=0 $Y2=0
cc_341 N_A_29_367#_c_409_n N_Y_c_584_n 0.00671999f $X=2.85 $Y=1.98 $X2=0 $Y2=0
cc_342 N_A_29_367#_c_410_n N_Y_c_584_n 0.045264f $X=5.285 $Y=2.41 $X2=0 $Y2=0
cc_343 N_A_29_367#_M1016_s N_Y_c_561_n 0.00330762f $X=5.29 $Y=1.835 $X2=0 $Y2=0
cc_344 N_A_29_367#_c_410_n N_Y_c_561_n 0.0177445f $X=5.285 $Y=2.41 $X2=0 $Y2=0
cc_345 N_A_29_367#_c_391_n N_Y_c_561_n 0.0230903f $X=5.45 $Y=2.24 $X2=0 $Y2=0
cc_346 N_A_29_367#_c_410_n N_Y_c_563_n 0.0161558f $X=5.285 $Y=2.41 $X2=0 $Y2=0
cc_347 N_VPWR_c_460_n N_A_456_367#_M1000_d 0.00223559f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_348 N_VPWR_c_460_n N_A_456_367#_M1003_d 0.00225186f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_460_n N_A_456_367#_M1011_d 0.00225186f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_460_n N_A_456_367#_M1021_d 0.00248137f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_465_n N_A_456_367#_c_528_n 0.01906f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_352 N_VPWR_c_460_n N_A_456_367#_c_528_n 0.0124545f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_465_n N_A_456_367#_c_533_n 0.146853f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPWR_c_460_n N_A_456_367#_c_533_n 0.0926003f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_460_n N_Y_M1004_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_356 N_VPWR_c_460_n N_Y_M1013_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_357 N_A_456_367#_c_533_n N_Y_M1004_s 0.00346062f $X=5 $Y=2.84 $X2=0 $Y2=0
cc_358 N_A_456_367#_c_533_n N_Y_M1013_s 0.00346062f $X=5 $Y=2.84 $X2=2.635
+ $Y2=1.185
cc_359 N_A_456_367#_M1011_d N_Y_c_584_n 0.00336444f $X=4 $Y=1.835 $X2=2.635
+ $Y2=1.35
cc_360 N_A_456_367#_M1021_d N_Y_c_561_n 0.00244731f $X=4.86 $Y=1.835 $X2=2.16
+ $Y2=1.362
cc_361 N_Y_c_564_n N_VGND_M1009_d 0.00329816f $X=1.465 $Y=0.955 $X2=0 $Y2=0
cc_362 N_Y_c_570_n N_VGND_M1019_d 0.00470293f $X=2.325 $Y=0.955 $X2=0 $Y2=0
cc_363 N_Y_c_577_n N_VGND_M1015_s 0.00154697f $X=3.115 $Y=0.81 $X2=0 $Y2=0
cc_364 N_Y_c_610_n N_VGND_M1015_s 0.00386499f $X=2.865 $Y=0.882 $X2=0 $Y2=0
cc_365 N_Y_c_583_n N_VGND_M1005_d 0.0033934f $X=3.975 $Y=0.81 $X2=0 $Y2=0
cc_366 N_Y_c_585_n N_VGND_M1012_d 0.0033934f $X=4.835 $Y=0.81 $X2=0 $Y2=0
cc_367 N_Y_c_559_n N_VGND_M1023_s 0.00740918f $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_368 N_Y_c_560_n N_VGND_M1023_s 0.00264016f $X=5.585 $Y=1.815 $X2=0 $Y2=0
cc_369 N_Y_c_564_n N_VGND_c_705_n 0.0170777f $X=1.465 $Y=0.955 $X2=0 $Y2=0
cc_370 N_Y_c_570_n N_VGND_c_706_n 0.0170777f $X=2.325 $Y=0.955 $X2=0 $Y2=0
cc_371 N_Y_c_610_n N_VGND_c_707_n 0.0132711f $X=2.865 $Y=0.882 $X2=0 $Y2=0
cc_372 N_Y_c_583_n N_VGND_c_708_n 0.0129852f $X=3.975 $Y=0.81 $X2=0 $Y2=0
cc_373 N_Y_c_585_n N_VGND_c_709_n 0.0129852f $X=4.835 $Y=0.81 $X2=0 $Y2=0
cc_374 N_Y_c_559_n N_VGND_c_710_n 0.00127671f $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_375 N_Y_c_559_n N_VGND_c_711_n 0.0201899f $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_376 N_Y_c_672_p N_VGND_c_712_n 0.0124525f $X=1.56 $Y=0.42 $X2=0 $Y2=0
cc_377 N_Y_c_673_p N_VGND_c_714_n 0.0135169f $X=2.42 $Y=0.42 $X2=0 $Y2=0
cc_378 N_Y_c_608_n N_VGND_c_714_n 0.0022105f $X=2.708 $Y=0.882 $X2=0 $Y2=0
cc_379 N_Y_c_577_n N_VGND_c_716_n 0.00200585f $X=3.115 $Y=0.81 $X2=0 $Y2=0
cc_380 N_Y_c_581_n N_VGND_c_716_n 0.0188581f $X=3.28 $Y=0.42 $X2=0 $Y2=0
cc_381 N_Y_c_583_n N_VGND_c_716_n 0.00200585f $X=3.975 $Y=0.81 $X2=0 $Y2=0
cc_382 N_Y_c_678_p N_VGND_c_718_n 0.0135169f $X=0.7 $Y=0.42 $X2=0 $Y2=0
cc_383 N_Y_c_583_n N_VGND_c_719_n 0.00200585f $X=3.975 $Y=0.81 $X2=0 $Y2=0
cc_384 N_Y_c_623_n N_VGND_c_719_n 0.0188581f $X=4.14 $Y=0.42 $X2=0 $Y2=0
cc_385 N_Y_c_585_n N_VGND_c_719_n 0.00200585f $X=4.835 $Y=0.81 $X2=0 $Y2=0
cc_386 N_Y_c_585_n N_VGND_c_720_n 0.00200585f $X=4.835 $Y=0.81 $X2=0 $Y2=0
cc_387 N_Y_c_590_n N_VGND_c_720_n 0.0188581f $X=5 $Y=0.42 $X2=0 $Y2=0
cc_388 N_Y_c_559_n N_VGND_c_720_n 0.00200585f $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_389 N_Y_M1001_s N_VGND_c_723_n 0.00432284f $X=0.56 $Y=0.235 $X2=0 $Y2=0
cc_390 N_Y_M1017_s N_VGND_c_723_n 0.00536646f $X=1.42 $Y=0.235 $X2=0 $Y2=0
cc_391 N_Y_M1008_d N_VGND_c_723_n 0.00386173f $X=2.28 $Y=0.235 $X2=0 $Y2=0
cc_392 N_Y_M1022_d N_VGND_c_723_n 0.00223559f $X=3.14 $Y=0.235 $X2=0 $Y2=0
cc_393 N_Y_M1007_s N_VGND_c_723_n 0.00223559f $X=4 $Y=0.235 $X2=0 $Y2=0
cc_394 N_Y_M1014_s N_VGND_c_723_n 0.00223559f $X=4.86 $Y=0.235 $X2=0 $Y2=0
cc_395 N_Y_c_678_p N_VGND_c_723_n 0.00847534f $X=0.7 $Y=0.42 $X2=0 $Y2=0
cc_396 N_Y_c_672_p N_VGND_c_723_n 0.00730901f $X=1.56 $Y=0.42 $X2=0 $Y2=0
cc_397 N_Y_c_673_p N_VGND_c_723_n 0.00847534f $X=2.42 $Y=0.42 $X2=0 $Y2=0
cc_398 N_Y_c_577_n N_VGND_c_723_n 0.0038586f $X=3.115 $Y=0.81 $X2=0 $Y2=0
cc_399 N_Y_c_581_n N_VGND_c_723_n 0.0123659f $X=3.28 $Y=0.42 $X2=0 $Y2=0
cc_400 N_Y_c_583_n N_VGND_c_723_n 0.00843758f $X=3.975 $Y=0.81 $X2=0 $Y2=0
cc_401 N_Y_c_623_n N_VGND_c_723_n 0.0123659f $X=4.14 $Y=0.42 $X2=0 $Y2=0
cc_402 N_Y_c_585_n N_VGND_c_723_n 0.00843758f $X=4.835 $Y=0.81 $X2=0 $Y2=0
cc_403 N_Y_c_590_n N_VGND_c_723_n 0.0123659f $X=5 $Y=0.42 $X2=0 $Y2=0
cc_404 N_Y_c_559_n N_VGND_c_723_n 0.00706673f $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_405 N_Y_c_608_n N_VGND_c_723_n 0.00377901f $X=2.708 $Y=0.882 $X2=0 $Y2=0
cc_406 N_Y_c_610_n N_VGND_c_723_n 9.04234e-19 $X=2.865 $Y=0.882 $X2=0 $Y2=0
