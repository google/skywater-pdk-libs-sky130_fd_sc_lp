* File: sky130_fd_sc_lp__nor2_1.pex.spice
* Created: Wed Sep  2 10:07:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_1%A 3 6 8 9 13 15
r22 13 16 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.46
+ $X2=0.382 $Y2=1.625
r23 13 15 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.46
+ $X2=0.382 $Y2=1.295
r24 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.46 $X2=0.35 $Y2=1.46
r25 9 14 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.46
r26 8 14 5.43295 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.46
r27 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=1.625
r28 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.505 $Y=0.765
+ $X2=0.505 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_1%B 3 5 7 8 9 16
r25 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.46 $X2=1.07 $Y2=1.46
r26 14 16 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.935 $Y=1.46
+ $X2=1.07 $Y2=1.46
r27 12 14 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.895 $Y=1.46
+ $X2=0.935 $Y2=1.46
r28 9 17 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.46
r29 8 17 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=1.295
+ $X2=1.17 $Y2=1.46
r30 5 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.295
+ $X2=0.935 $Y2=1.46
r31 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=1.295
+ $X2=0.935 $Y2=0.765
r32 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.625
+ $X2=0.895 $Y2=1.46
r33 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.895 $Y=1.625
+ $X2=0.895 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_1%VPWR 1 4 6 10 14 15
r17 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r18 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r19 12 18 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r20 12 14 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r21 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r22 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 6 9 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.29 $Y=2.005
+ $X2=0.29 $Y2=2.95
r24 4 18 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.227 $Y2=3.33
r25 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.95
r26 1 9 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.95
r27 1 6 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_1%Y 1 2 7 8 9 10 11 12 13 41
c21 41 0 5.39665e-20 $X=1.11 $Y=2.005
c22 7 0 1.39483e-20 $X=0.72 $Y=0.555
r23 41 42 8.20685 $w=6.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.95 $Y=2.005
+ $X2=0.95 $Y2=1.92
r24 13 38 2.48416 $w=6.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.95 $Y=2.775
+ $X2=0.95 $Y2=2.91
r25 12 13 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.95 $Y=2.405
+ $X2=0.95 $Y2=2.775
r26 12 32 2.94419 $w=6.48e-07 $l=1.6e-07 $layer=LI1_cond $X=0.95 $Y=2.405
+ $X2=0.95 $Y2=2.245
r27 11 32 3.86425 $w=6.48e-07 $l=2.1e-07 $layer=LI1_cond $X=0.95 $Y=2.035
+ $X2=0.95 $Y2=2.245
r28 11 41 0.552036 $w=6.48e-07 $l=3e-08 $layer=LI1_cond $X=0.95 $Y=2.035
+ $X2=0.95 $Y2=2.005
r29 10 42 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=1.92
r30 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.665
r31 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=0.925 $X2=0.72
+ $Y2=1.295
r32 7 8 25.3923 $w=1.88e-07 $l=4.35e-07 $layer=LI1_cond $X=0.72 $Y=0.49 $X2=0.72
+ $Y2=0.925
r33 2 41 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.835 $X2=1.11 $Y2=2.005
r34 2 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.835 $X2=1.11 $Y2=2.91
r35 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.345 $X2=0.72 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_1%VGND 1 2 7 9 11 13 15 17 27
r22 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r23 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 18 23 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r25 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r26 17 26 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.212
+ $Y2=0
r27 17 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r28 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r29 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r30 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 11 26 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.212 $Y2=0
r32 11 13 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.49
r33 7 23 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r34 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.29 $Y2=0.49
r35 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.345 $X2=1.15 $Y2=0.49
r36 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.345 $X2=0.29 $Y2=0.49
.ends

