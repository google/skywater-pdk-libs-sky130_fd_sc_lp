* File: sky130_fd_sc_lp__inv_4.pxi.spice
* Created: Fri Aug 28 10:38:20 2020
* 
x_PM_SKY130_FD_SC_LP__INV_4%A N_A_c_41_n N_A_M1000_g N_A_M1003_g N_A_c_43_n
+ N_A_M1001_g N_A_M1004_g N_A_c_45_n N_A_M1002_g N_A_M1006_g N_A_c_47_n
+ N_A_M1005_g N_A_M1007_g A A A A N_A_c_50_n PM_SKY130_FD_SC_LP__INV_4%A
x_PM_SKY130_FD_SC_LP__INV_4%VPWR N_VPWR_M1003_d N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_c_108_n N_VPWR_c_109_n N_VPWR_c_110_n N_VPWR_c_111_n N_VPWR_c_112_n
+ N_VPWR_c_113_n N_VPWR_c_114_n VPWR N_VPWR_c_115_n N_VPWR_c_107_n
+ PM_SKY130_FD_SC_LP__INV_4%VPWR
x_PM_SKY130_FD_SC_LP__INV_4%Y N_Y_M1000_d N_Y_M1002_d N_Y_M1003_s N_Y_M1006_s
+ N_Y_c_175_n N_Y_c_191_p N_Y_c_149_n N_Y_c_153_n N_Y_c_144_n N_Y_c_145_n
+ N_Y_c_180_n N_Y_c_192_p N_Y_c_162_n N_Y_c_146_n N_Y_c_147_n N_Y_c_168_n Y Y Y
+ N_Y_c_143_n PM_SKY130_FD_SC_LP__INV_4%Y
x_PM_SKY130_FD_SC_LP__INV_4%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1005_s
+ N_VGND_c_199_n N_VGND_c_200_n N_VGND_c_201_n N_VGND_c_202_n N_VGND_c_203_n
+ N_VGND_c_204_n N_VGND_c_205_n VGND N_VGND_c_206_n N_VGND_c_207_n
+ PM_SKY130_FD_SC_LP__INV_4%VGND
cc_1 VNB N_A_c_41_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.185
cc_2 VNB N_A_M1003_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_3 VNB N_A_c_43_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.185
cc_4 VNB N_A_M1004_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_5 VNB N_A_c_45_n 0.0162035f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.185
cc_6 VNB N_A_M1006_g 0.00706662f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=2.465
cc_7 VNB N_A_c_47_n 0.0193934f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.185
cc_8 VNB N_A_M1007_g 0.00775814f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.465
cc_9 VNB A 0.0163646f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_10 VNB N_A_c_50_n 0.106575f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.35
cc_11 VNB N_VPWR_c_107_n 0.103974f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.35
cc_12 VNB Y 0.0331739f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.35
cc_13 VNB N_Y_c_143_n 0.0129811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_199_n 0.0110651f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.655
cc_15 VNB N_VGND_c_200_n 0.0356924f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_16 VNB N_VGND_c_201_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.655
cc_17 VNB N_VGND_c_202_n 0.0158498f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.515
cc_18 VNB N_VGND_c_203_n 0.0215697f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=2.465
cc_19 VNB N_VGND_c_204_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=0.655
cc_20 VNB N_VGND_c_205_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=0.655
cc_21 VNB N_VGND_c_206_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_22 VNB N_VGND_c_207_n 0.149821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VPB N_A_M1003_g 0.0272503f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_24 VPB N_A_M1004_g 0.0191131f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_25 VPB N_A_M1006_g 0.0190939f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=2.465
cc_26 VPB N_A_M1007_g 0.0234365f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=2.465
cc_27 VPB N_VPWR_c_108_n 0.010943f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.655
cc_28 VPB N_VPWR_c_109_n 0.0561597f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_29 VPB N_VPWR_c_110_n 0.00399476f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.515
cc_30 VPB N_VPWR_c_111_n 0.015824f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=1.185
cc_31 VPB N_VPWR_c_112_n 0.0431603f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=0.655
cc_32 VPB N_VPWR_c_113_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_33 VPB N_VPWR_c_114_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_34 VPB N_VPWR_c_115_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.35
cc_35 VPB N_VPWR_c_107_n 0.049953f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.35
cc_36 VPB N_Y_c_144_n 0.00266319f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=1.515
cc_37 VPB N_Y_c_145_n 0.00350303f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=2.465
cc_38 VPB N_Y_c_146_n 0.0210875f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.35
cc_39 VPB N_Y_c_147_n 0.00247054f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.35
cc_40 VPB Y 0.0056227f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.35
cc_41 N_A_M1003_g N_VPWR_c_109_n 0.00767615f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_42 A N_VPWR_c_109_n 0.0160645f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_43 N_A_c_50_n N_VPWR_c_109_n 0.00505774f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_44 N_A_M1004_g N_VPWR_c_110_n 0.00163834f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_45 N_A_M1006_g N_VPWR_c_110_n 0.0016166f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_46 N_A_M1007_g N_VPWR_c_112_n 0.00344465f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_47 N_A_M1003_g N_VPWR_c_113_n 0.00585385f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_48 N_A_M1004_g N_VPWR_c_113_n 0.00585385f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_49 N_A_M1006_g N_VPWR_c_115_n 0.00585385f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_50 N_A_M1007_g N_VPWR_c_115_n 0.00585385f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_51 N_A_M1003_g N_VPWR_c_107_n 0.0114734f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_52 N_A_M1004_g N_VPWR_c_107_n 0.0105224f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A_M1006_g N_VPWR_c_107_n 0.0105361f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_M1007_g N_VPWR_c_107_n 0.0115723f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A_c_43_n N_Y_c_149_n 0.0129934f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_56 N_A_c_45_n N_Y_c_149_n 0.0129469f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_57 A N_Y_c_149_n 0.0383711f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A_c_50_n N_Y_c_149_n 0.00230884f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_59 A N_Y_c_153_n 0.0171348f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A_c_50_n N_Y_c_153_n 0.00240082f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_Y_c_144_n 0.014207f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A_M1006_g N_Y_c_144_n 0.014313f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_63 A N_Y_c_144_n 0.0331355f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A_c_50_n N_Y_c_144_n 0.00213862f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_Y_c_145_n 0.00219544f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_66 A N_Y_c_145_n 0.0171881f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_c_50_n N_Y_c_145_n 0.00224327f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_68 N_A_c_47_n N_Y_c_162_n 0.0128601f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_69 A N_Y_c_162_n 0.0111091f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_M1007_g N_Y_c_146_n 0.0160651f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_71 A N_Y_c_146_n 0.00862873f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_72 A N_Y_c_147_n 0.0171881f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_c_50_n N_Y_c_147_n 0.00224327f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_74 A N_Y_c_168_n 0.0171348f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_50_n N_Y_c_168_n 0.00240082f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_76 N_A_c_47_n Y 0.00628625f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_77 A Y 0.0240168f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_c_50_n Y 0.0107799f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_79 N_A_c_41_n N_VGND_c_200_n 0.00555149f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_80 A N_VGND_c_200_n 0.0222878f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_c_50_n N_VGND_c_200_n 0.00559057f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_82 N_A_c_43_n N_VGND_c_201_n 0.00211454f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_83 N_A_c_45_n N_VGND_c_201_n 0.00211454f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_84 N_A_c_47_n N_VGND_c_203_n 0.00492463f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_85 N_A_c_41_n N_VGND_c_204_n 0.00585385f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_86 N_A_c_43_n N_VGND_c_204_n 0.00585385f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_87 N_A_c_45_n N_VGND_c_206_n 0.00585385f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_88 N_A_c_47_n N_VGND_c_206_n 0.00585385f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_89 N_A_c_41_n N_VGND_c_207_n 0.0114597f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_90 N_A_c_43_n N_VGND_c_207_n 0.0106297f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A_c_45_n N_VGND_c_207_n 0.0106297f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A_c_47_n N_VGND_c_207_n 0.00734271f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_93 N_VPWR_c_107_n N_Y_M1003_s 0.0027574f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_94 N_VPWR_c_107_n N_Y_M1006_s 0.0027574f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_95 N_VPWR_c_113_n N_Y_c_175_n 0.0151136f $X=0.995 $Y=3.33 $X2=0 $Y2=0
cc_96 N_VPWR_c_107_n N_Y_c_175_n 0.0102248f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_97 N_VPWR_M1004_d N_Y_c_144_n 0.00176461f $X=0.985 $Y=1.835 $X2=0 $Y2=0
cc_98 N_VPWR_c_110_n N_Y_c_144_n 0.0135055f $X=1.125 $Y=2.26 $X2=0 $Y2=0
cc_99 N_VPWR_c_109_n N_Y_c_145_n 0.00166417f $X=0.265 $Y=1.98 $X2=0 $Y2=0
cc_100 N_VPWR_c_115_n N_Y_c_180_n 0.0151136f $X=1.855 $Y=3.33 $X2=0 $Y2=0
cc_101 N_VPWR_c_107_n N_Y_c_180_n 0.0102248f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_102 N_VPWR_M1007_d N_Y_c_146_n 0.00266094f $X=1.845 $Y=1.835 $X2=0 $Y2=0
cc_103 N_VPWR_c_112_n N_Y_c_146_n 0.0212886f $X=1.985 $Y=2.26 $X2=0 $Y2=0
cc_104 N_Y_c_149_n N_VGND_M1001_s 0.00329816f $X=1.425 $Y=0.955 $X2=0 $Y2=0
cc_105 N_Y_c_162_n N_VGND_M1005_s 0.00603322f $X=2.025 $Y=0.94 $X2=0 $Y2=0
cc_106 Y N_VGND_M1005_s 5.78869e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_107 N_Y_c_143_n N_VGND_M1005_s 0.00186881f $X=2.162 $Y=1.04 $X2=0 $Y2=0
cc_108 N_Y_c_149_n N_VGND_c_201_n 0.0135055f $X=1.425 $Y=0.955 $X2=0 $Y2=0
cc_109 N_Y_c_162_n N_VGND_c_203_n 0.00985756f $X=2.025 $Y=0.94 $X2=0 $Y2=0
cc_110 N_Y_c_143_n N_VGND_c_203_n 0.0110452f $X=2.162 $Y=1.04 $X2=0 $Y2=0
cc_111 N_Y_c_191_p N_VGND_c_204_n 0.0149362f $X=0.695 $Y=0.42 $X2=0 $Y2=0
cc_112 N_Y_c_192_p N_VGND_c_206_n 0.0149362f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_113 N_Y_M1000_d N_VGND_c_207_n 0.00293134f $X=0.555 $Y=0.235 $X2=0 $Y2=0
cc_114 N_Y_M1002_d N_VGND_c_207_n 0.00263512f $X=1.415 $Y=0.235 $X2=0 $Y2=0
cc_115 N_Y_c_191_p N_VGND_c_207_n 0.0100304f $X=0.695 $Y=0.42 $X2=0 $Y2=0
cc_116 N_Y_c_192_p N_VGND_c_207_n 0.0100304f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_117 N_Y_c_162_n N_VGND_c_207_n 0.00534191f $X=2.025 $Y=0.94 $X2=0 $Y2=0
cc_118 N_Y_c_143_n N_VGND_c_207_n 0.00640524f $X=2.162 $Y=1.04 $X2=0 $Y2=0
