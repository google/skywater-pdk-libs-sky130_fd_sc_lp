* File: sky130_fd_sc_lp__o221ai_2.pex.spice
* Created: Fri Aug 28 11:08:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221AI_2%C1 1 3 6 8 10 13 15 16 24
r40 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.485 $Y=1.46
+ $X2=0.915 $Y2=1.46
r41 20 23 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.485 $Y2=1.46
r42 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.46 $X2=0.27 $Y2=1.46
r43 16 21 8.91512 $w=2.63e-07 $l=2.05e-07 $layer=LI1_cond $X=0.222 $Y=1.665
+ $X2=0.222 $Y2=1.46
r44 15 21 7.17559 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.222 $Y=1.295
+ $X2=0.222 $Y2=1.46
r45 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.625
+ $X2=0.915 $Y2=1.46
r46 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.915 $Y=1.625
+ $X2=0.915 $Y2=2.465
r47 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.295
+ $X2=0.915 $Y2=1.46
r48 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.915 $Y=1.295
+ $X2=0.915 $Y2=0.765
r49 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.625
+ $X2=0.485 $Y2=1.46
r50 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.485 $Y=1.625
+ $X2=0.485 $Y2=2.465
r51 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.295
+ $X2=0.485 $Y2=1.46
r52 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.485 $Y=1.295
+ $X2=0.485 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%B1 5 9 13 17 19 20 23 24 26 27 31
c96 23 0 9.34296e-20 $X=3.305 $Y=1.51
c97 13 0 5.57328e-20 $X=3.225 $Y=2.465
r98 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.855
+ $Y=1.51 $X2=1.855 $Y2=1.51
r99 27 32 8.92326 $w=4.17e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=1.65
+ $X2=1.855 $Y2=1.65
r100 26 32 5.1199 $w=4.17e-07 $l=1.75e-07 $layer=LI1_cond $X=1.68 $Y=1.65
+ $X2=1.855 $Y2=1.65
r101 24 35 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.51
+ $X2=3.275 $Y2=1.675
r102 24 34 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.51
+ $X2=3.275 $Y2=1.345
r103 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.305
+ $Y=1.51 $X2=3.305 $Y2=1.51
r104 21 23 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.305 $Y=1.705
+ $X2=3.305 $Y2=1.51
r105 20 27 8.94133 $w=4.17e-07 $l=2.13834e-07 $layer=LI1_cond $X=2.315 $Y=1.79
+ $X2=2.16 $Y2=1.65
r106 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.14 $Y=1.79
+ $X2=3.305 $Y2=1.705
r107 19 20 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.14 $Y=1.79
+ $X2=2.315 $Y2=1.79
r108 17 34 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.395 $Y=0.745
+ $X2=3.395 $Y2=1.345
r109 13 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.225 $Y=2.465
+ $X2=3.225 $Y2=1.675
r110 7 31 37.0704 $w=1.5e-07 $l=1.83916e-07 $layer=POLY_cond $X=1.865 $Y=1.675
+ $X2=1.905 $Y2=1.51
r111 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.865 $Y=1.675
+ $X2=1.865 $Y2=2.465
r112 3 31 37.0704 $w=1.5e-07 $l=1.83916e-07 $layer=POLY_cond $X=1.865 $Y=1.345
+ $X2=1.905 $Y2=1.51
r113 3 5 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.865 $Y=1.345 $X2=1.865
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%B2 1 3 6 8 10 13 15 22
c56 1 0 6.7205e-20 $X=2.365 $Y=1.275
r57 20 22 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.44
+ $X2=2.795 $Y2=1.44
r58 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.44 $X2=2.67 $Y2=1.44
r59 17 20 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.365 $Y=1.44
+ $X2=2.67 $Y2=1.44
r60 15 21 4.77441 $w=3.48e-07 $l=1.45e-07 $layer=LI1_cond $X=2.66 $Y=1.295
+ $X2=2.66 $Y2=1.44
r61 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.605
+ $X2=2.795 $Y2=1.44
r62 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.795 $Y=1.605
+ $X2=2.795 $Y2=2.465
r63 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.275
+ $X2=2.795 $Y2=1.44
r64 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.795 $Y=1.275
+ $X2=2.795 $Y2=0.745
r65 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.605
+ $X2=2.365 $Y2=1.44
r66 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.365 $Y=1.605
+ $X2=2.365 $Y2=2.465
r67 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.275
+ $X2=2.365 $Y2=1.44
r68 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.365 $Y=1.275
+ $X2=2.365 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%A1 3 7 9 11 14 18 19 21 22 23 24 35 38 45
c85 19 0 1.62328e-19 $X=3.845 $Y=1.51
c86 18 0 5.57328e-20 $X=3.845 $Y=1.51
c87 7 0 9.34296e-20 $X=3.895 $Y=2.465
r88 38 45 1.06379 $w=3.23e-07 $l=3e-08 $layer=LI1_cond $X=5.507 $Y=1.695
+ $X2=5.507 $Y2=1.665
r89 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.44 $X2=5.49 $Y2=1.44
r90 33 35 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=5.265 $Y=1.44
+ $X2=5.49 $Y2=1.44
r91 31 33 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.195 $Y=1.44
+ $X2=5.265 $Y2=1.44
r92 24 38 2.70504 $w=3.25e-07 $l=9e-08 $layer=LI1_cond $X=5.507 $Y=1.785
+ $X2=5.507 $Y2=1.695
r93 24 45 0.992874 $w=3.23e-07 $l=2.8e-08 $layer=LI1_cond $X=5.507 $Y=1.637
+ $X2=5.507 $Y2=1.665
r94 24 36 6.98558 $w=3.23e-07 $l=1.97e-07 $layer=LI1_cond $X=5.507 $Y=1.637
+ $X2=5.507 $Y2=1.44
r95 23 36 5.14167 $w=3.23e-07 $l=1.45e-07 $layer=LI1_cond $X=5.507 $Y=1.295
+ $X2=5.507 $Y2=1.44
r96 21 24 4.86908 $w=1.8e-07 $l=1.62e-07 $layer=LI1_cond $X=5.345 $Y=1.785
+ $X2=5.507 $Y2=1.785
r97 21 22 81.9495 $w=1.78e-07 $l=1.33e-06 $layer=LI1_cond $X=5.345 $Y=1.785
+ $X2=4.015 $Y2=1.785
r98 19 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.51
+ $X2=3.845 $Y2=1.675
r99 19 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.51
+ $X2=3.845 $Y2=1.345
r100 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.51 $X2=3.845 $Y2=1.51
r101 16 22 7.65203 $w=1.8e-07 $l=2.08192e-07 $layer=LI1_cond $X=3.847 $Y=1.695
+ $X2=4.015 $Y2=1.785
r102 16 18 6.36424 $w=3.33e-07 $l=1.85e-07 $layer=LI1_cond $X=3.847 $Y=1.695
+ $X2=3.847 $Y2=1.51
r103 12 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.605
+ $X2=5.265 $Y2=1.44
r104 12 14 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.265 $Y=1.605
+ $X2=5.265 $Y2=2.465
r105 9 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.195 $Y=1.275
+ $X2=5.195 $Y2=1.44
r106 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.195 $Y=1.275
+ $X2=5.195 $Y2=0.745
r107 7 30 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.895 $Y=2.465
+ $X2=3.895 $Y2=1.675
r108 3 29 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.825 $Y=0.745
+ $X2=3.825 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%A2 1 3 6 8 10 13 15 16 29
r55 27 29 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.745 $Y=1.44
+ $X2=4.835 $Y2=1.44
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=1.44 $X2=4.745 $Y2=1.44
r57 25 27 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.725 $Y=1.44
+ $X2=4.745 $Y2=1.44
r58 24 25 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=4.405 $Y=1.44
+ $X2=4.725 $Y2=1.44
r59 22 24 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.385 $Y=1.44
+ $X2=4.405 $Y2=1.44
r60 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.385
+ $Y=1.44 $X2=4.385 $Y2=1.44
r61 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.295 $Y=1.44
+ $X2=4.385 $Y2=1.44
r62 16 28 10.7927 $w=3.13e-07 $l=2.95e-07 $layer=LI1_cond $X=5.04 $Y=1.367
+ $X2=4.745 $Y2=1.367
r63 15 28 6.76832 $w=3.13e-07 $l=1.85e-07 $layer=LI1_cond $X=4.56 $Y=1.367
+ $X2=4.745 $Y2=1.367
r64 15 23 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=4.56 $Y=1.367
+ $X2=4.385 $Y2=1.367
r65 11 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.605
+ $X2=4.835 $Y2=1.44
r66 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.835 $Y=1.605
+ $X2=4.835 $Y2=2.465
r67 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.725 $Y=1.275
+ $X2=4.725 $Y2=1.44
r68 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.725 $Y=1.275
+ $X2=4.725 $Y2=0.745
r69 4 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.605
+ $X2=4.405 $Y2=1.44
r70 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.405 $Y=1.605
+ $X2=4.405 $Y2=2.465
r71 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.275
+ $X2=4.295 $Y2=1.44
r72 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.295 $Y=1.275
+ $X2=4.295 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%VPWR 1 2 3 4 13 15 21 25 27 29 33 35 40 48
+ 60 63 67
r78 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r81 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r82 55 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 52 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r86 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=5.04
+ $Y2=3.33
r87 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 49 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=3.56 $Y2=3.33
r89 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 48 66 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.537 $Y2=3.33
r91 48 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.04 $Y2=3.33
r92 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r93 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 44 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r96 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 41 60 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.39 $Y2=3.33
r98 41 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.56 $Y2=3.33
r100 40 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 39 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 39 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 36 57 4.11164 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r105 36 38 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 35 60 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.39 $Y2=3.33
r107 35 38 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 33 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 33 44 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 29 32 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=5.48 $Y=2.13
+ $X2=5.48 $Y2=2.95
r111 27 66 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.537 $Y2=3.33
r112 27 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.48 $Y2=2.95
r113 23 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=3.33
r114 23 25 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.51
r115 19 60 3.24638 $w=8.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=3.33
r116 19 21 10.8365 $w=8.48e-07 $l=7.55e-07 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=2.49
r117 15 18 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=0.235 $Y=2.085
+ $X2=0.235 $Y2=2.95
r118 13 57 3.10058 $w=2.6e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.182 $Y2=3.33
r119 13 18 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.235 $Y2=2.95
r120 4 32 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.34
+ $Y=1.835 $X2=5.48 $Y2=2.95
r121 4 29 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=5.34
+ $Y=1.835 $X2=5.48 $Y2=2.13
r122 3 25 300 $w=1.7e-07 $l=7.94434e-07 $layer=licon1_PDIFF $count=2 $X=3.3
+ $Y=1.835 $X2=3.56 $Y2=2.51
r123 2 21 150 $w=1.7e-07 $l=9.31612e-07 $layer=licon1_PDIFF $count=4 $X=0.99
+ $Y=1.835 $X2=1.65 $Y2=2.49
r124 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.95
r125 1 15 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%Y 1 2 3 4 15 17 18 21 26 28 29 30 31 32 33
+ 41
r65 32 33 15.4822 $w=3.94e-07 $l=5e-07 $layer=LI1_cond $X=0.7 $Y=2.015 $X2=1.2
+ $Y2=2.015
r66 32 49 1.08376 $w=3.94e-07 $l=3.5e-08 $layer=LI1_cond $X=0.7 $Y=2.015
+ $X2=0.665 $Y2=2.015
r67 32 39 1.77687 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=0.7 $Y=2.015 $X2=0.7
+ $Y2=1.815
r68 31 39 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.7 $Y=1.665 $X2=0.7
+ $Y2=1.815
r69 30 31 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=1.295 $X2=0.7
+ $Y2=1.665
r70 29 30 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=0.925 $X2=0.7
+ $Y2=1.295
r71 29 41 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.7 $Y=0.925
+ $X2=0.7 $Y2=0.68
r72 22 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=2.13
+ $X2=2.58 $Y2=2.13
r73 21 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=2.13
+ $X2=4.62 $Y2=2.13
r74 21 22 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=4.455 $Y=2.13
+ $X2=2.745 $Y2=2.13
r75 18 33 8.19978 $w=3.94e-07 $l=1.83712e-07 $layer=LI1_cond $X=1.335 $Y=2.13
+ $X2=1.2 $Y2=2.015
r76 17 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=2.13
+ $X2=2.58 $Y2=2.13
r77 17 18 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=2.415 $Y=2.13
+ $X2=1.335 $Y2=2.13
r78 13 49 3.17004 $w=2.6e-07 $l=2e-07 $layer=LI1_cond $X=0.665 $Y=2.215
+ $X2=0.665 $Y2=2.015
r79 13 15 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.665 $Y=2.215
+ $X2=0.665 $Y2=2.435
r80 4 28 300 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=2 $X=4.48
+ $Y=1.835 $X2=4.62 $Y2=2.13
r81 3 26 300 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=2 $X=2.44
+ $Y=1.835 $X2=2.58 $Y2=2.13
r82 2 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=1.98
r83 2 15 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.435
r84 1 41 91 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.345 $X2=0.7 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%A_388_367# 1 2 9 11 12 15
r20 13 15 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=3.045 $Y=2.905
+ $X2=3.045 $Y2=2.55
r21 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.915 $Y=2.99
+ $X2=3.045 $Y2=2.905
r22 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.915 $Y=2.99
+ $X2=2.245 $Y2=2.99
r23 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.115 $Y=2.905
+ $X2=2.245 $Y2=2.99
r24 7 9 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=2.115 $Y=2.905
+ $X2=2.115 $Y2=2.55
r25 2 15 300 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=2 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=2.55
r26 1 9 300 $w=1.7e-07 $l=7.97716e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=1.835 $X2=2.115 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%A_794_367# 1 2 9 11 12 13 15
r17 13 18 3.31928 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=5.05 $Y=2.895 $X2=5.05
+ $Y2=2.985
r18 13 15 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=5.05 $Y=2.895
+ $X2=5.05 $Y2=2.21
r19 11 18 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.955 $Y=2.985
+ $X2=5.05 $Y2=2.985
r20 11 12 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.955 $Y=2.985
+ $X2=4.285 $Y2=2.985
r21 7 12 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=4.155 $Y=2.895
+ $X2=4.285 $Y2=2.985
r22 7 9 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=4.155 $Y=2.895
+ $X2=4.155 $Y2=2.55
r23 2 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.835 $X2=5.05 $Y2=2.91
r24 2 15 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.835 $X2=5.05 $Y2=2.21
r25 1 9 300 $w=1.7e-07 $l=8.17634e-07 $layer=licon1_PDIFF $count=2 $X=3.97
+ $Y=1.835 $X2=4.19 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%A_29_69# 1 2 3 4 15 17 18 22 23 24 25 28 34
c56 23 0 6.7205e-20 $X=1.985 $Y=1.17
r57 34 35 7.40618 $w=4.53e-07 $l=2.75e-07 $layer=LI1_cond $X=3.105 $Y=0.68
+ $X2=3.105 $Y2=0.955
r58 30 31 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.15 $Y=0.955
+ $X2=2.15 $Y2=1.17
r59 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.15 $Y=0.68
+ $X2=2.15 $Y2=0.955
r60 26 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0.955
+ $X2=2.15 $Y2=0.955
r61 25 35 6.54142 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.865 $Y=0.955
+ $X2=3.105 $Y2=0.955
r62 25 26 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.865 $Y=0.955
+ $X2=2.315 $Y2=0.955
r63 23 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=1.17
+ $X2=2.15 $Y2=1.17
r64 23 24 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.985 $Y=1.17
+ $X2=1.235 $Y2=1.17
r65 20 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.14 $Y=1.085
+ $X2=1.235 $Y2=1.17
r66 20 22 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=1.14 $Y=1.085
+ $X2=1.14 $Y2=0.49
r67 19 22 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=1.14 $Y=0.425
+ $X2=1.14 $Y2=0.49
r68 17 19 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.14 $Y2=0.425
r69 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.365 $Y2=0.34
r70 13 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.365 $Y2=0.34
r71 13 15 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.235 $Y2=0.49
r72 4 34 91 $w=1.7e-07 $l=4.2758e-07 $layer=licon1_NDIFF $count=2 $X=2.87
+ $Y=0.325 $X2=3.03 $Y2=0.68
r73 3 28 91 $w=1.7e-07 $l=4.47856e-07 $layer=licon1_NDIFF $count=2 $X=1.94
+ $Y=0.325 $X2=2.15 $Y2=0.68
r74 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.99
+ $Y=0.345 $X2=1.13 $Y2=0.49
r75 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.345 $X2=0.27 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%A_305_65# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 40 42 44 46
c70 33 0 1.62328e-19 $X=3.715 $Y=0.955
r71 40 48 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=0.87
+ $X2=5.435 $Y2=0.955
r72 40 42 16.4635 $w=2.78e-07 $l=4e-07 $layer=LI1_cond $X=5.435 $Y=0.87
+ $X2=5.435 $Y2=0.47
r73 39 46 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.625 $Y=0.955
+ $X2=4.51 $Y2=0.955
r74 38 48 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.295 $Y=0.955
+ $X2=5.435 $Y2=0.955
r75 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=0.955
+ $X2=4.625 $Y2=0.955
r76 34 46 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=0.87
+ $X2=4.51 $Y2=0.955
r77 34 36 20.0425 $w=2.28e-07 $l=4e-07 $layer=LI1_cond $X=4.51 $Y=0.87 $X2=4.51
+ $Y2=0.47
r78 32 46 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.395 $Y=0.955
+ $X2=4.51 $Y2=0.955
r79 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.395 $Y=0.955
+ $X2=3.715 $Y2=0.955
r80 29 33 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.615 $Y=0.87
+ $X2=3.715 $Y2=0.955
r81 29 31 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=3.615 $Y=0.87
+ $X2=3.615 $Y2=0.47
r82 28 31 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=3.615 $Y=0.425
+ $X2=3.615 $Y2=0.47
r83 27 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.695 $Y=0.34
+ $X2=2.59 $Y2=0.34
r84 26 28 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.515 $Y=0.34
+ $X2=3.615 $Y2=0.425
r85 26 27 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.515 $Y=0.34
+ $X2=2.695 $Y2=0.34
r86 22 44 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.425
+ $X2=2.59 $Y2=0.34
r87 22 24 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=2.59 $Y=0.425
+ $X2=2.59 $Y2=0.535
r88 20 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.485 $Y=0.34
+ $X2=2.59 $Y2=0.34
r89 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.485 $Y=0.34
+ $X2=1.815 $Y2=0.34
r90 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.65 $Y=0.425
+ $X2=1.815 $Y2=0.34
r91 16 18 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.65 $Y=0.425
+ $X2=1.65 $Y2=0.47
r92 5 48 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=5.27
+ $Y=0.325 $X2=5.41 $Y2=0.955
r93 5 42 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.27
+ $Y=0.325 $X2=5.41 $Y2=0.47
r94 4 46 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.325 $X2=4.51 $Y2=0.955
r95 4 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.325 $X2=4.51 $Y2=0.47
r96 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.47
+ $Y=0.325 $X2=3.61 $Y2=0.47
r97 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.325 $X2=2.58 $Y2=0.535
r98 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.325 $X2=1.65 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_2%VGND 1 2 9 13 15 17 25 32 33 36 39
r59 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r60 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r63 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=4.96
+ $Y2=0
r64 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=5.52
+ $Y2=0
r65 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r66 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r67 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r68 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.06
+ $Y2=0
r69 26 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.56
+ $Y2=0
r70 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.96
+ $Y2=0
r71 25 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.56
+ $Y2=0
r72 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r73 23 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r74 19 23 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r75 19 20 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r76 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.06
+ $Y2=0
r77 17 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=3.6
+ $Y2=0
r78 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r79 15 20 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.24
+ $Y2=0
r80 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r81 11 13 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.575
r82 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=0.085 $X2=4.06
+ $Y2=0
r83 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.06 $Y=0.085 $X2=4.06
+ $Y2=0.575
r84 2 13 182 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_NDIFF $count=1 $X=4.8
+ $Y=0.325 $X2=4.96 $Y2=0.575
r85 1 9 182 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.325 $X2=4.06 $Y2=0.575
.ends

