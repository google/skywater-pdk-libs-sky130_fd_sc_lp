* File: sky130_fd_sc_lp__o31ai_1.pxi.spice
* Created: Wed Sep  2 10:25:13 2020
* 
x_PM_SKY130_FD_SC_LP__O31AI_1%A1 N_A1_M1004_g N_A1_M1007_g A1 A1 N_A1_c_50_n
+ PM_SKY130_FD_SC_LP__O31AI_1%A1
x_PM_SKY130_FD_SC_LP__O31AI_1%A2 N_A2_M1006_g N_A2_M1005_g A2 A2 A2 A2
+ N_A2_c_73_n N_A2_c_74_n PM_SKY130_FD_SC_LP__O31AI_1%A2
x_PM_SKY130_FD_SC_LP__O31AI_1%A3 N_A3_M1002_g N_A3_M1003_g A3 A3 N_A3_c_116_n
+ PM_SKY130_FD_SC_LP__O31AI_1%A3
x_PM_SKY130_FD_SC_LP__O31AI_1%B1 N_B1_M1000_g N_B1_M1001_g N_B1_c_150_n B1
+ N_B1_c_151_n N_B1_c_152_n PM_SKY130_FD_SC_LP__O31AI_1%B1
x_PM_SKY130_FD_SC_LP__O31AI_1%VPWR N_VPWR_M1007_s N_VPWR_M1000_d N_VPWR_c_179_n
+ N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_182_n N_VPWR_c_183_n VPWR
+ N_VPWR_c_184_n N_VPWR_c_178_n PM_SKY130_FD_SC_LP__O31AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O31AI_1%Y N_Y_M1001_d N_Y_M1002_d N_Y_c_213_n N_Y_c_214_n
+ N_Y_c_215_n Y Y Y PM_SKY130_FD_SC_LP__O31AI_1%Y
x_PM_SKY130_FD_SC_LP__O31AI_1%VGND N_VGND_M1004_s N_VGND_M1005_d N_VGND_c_250_n
+ N_VGND_c_251_n VGND N_VGND_c_252_n N_VGND_c_253_n N_VGND_c_254_n
+ N_VGND_c_255_n PM_SKY130_FD_SC_LP__O31AI_1%VGND
x_PM_SKY130_FD_SC_LP__O31AI_1%A_110_47# N_A_110_47#_M1004_d N_A_110_47#_M1003_d
+ N_A_110_47#_c_308_n N_A_110_47#_c_292_n N_A_110_47#_c_301_n
+ N_A_110_47#_c_290_n PM_SKY130_FD_SC_LP__O31AI_1%A_110_47#
cc_1 VNB N_A1_M1004_g 0.0234223f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A1_M1007_g 0.00606695f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB A1 0.020304f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_50_n 0.0477491f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_5 VNB N_A2_M1005_g 0.0286148f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_6 VNB N_A2_c_73_n 0.0243737f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_7 VNB N_A2_c_74_n 0.00482117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A3_M1003_g 0.0282725f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_9 VNB A3 0.00242367f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A3_c_116_n 0.0350928f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_11 VNB N_B1_M1000_g 0.00161591f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_12 VNB N_B1_M1001_g 0.0290784f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_13 VNB N_B1_c_150_n 0.0110156f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_B1_c_151_n 0.0610027f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_15 VNB N_B1_c_152_n 0.0122438f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_16 VNB N_VPWR_c_178_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_213_n 0.0152384f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_18 VNB N_Y_c_214_n 0.00199942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_215_n 0.0296037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.00458121f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_21 VNB N_VGND_c_250_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_22 VNB N_VGND_c_251_n 0.0339261f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_VGND_c_252_n 0.034895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_253_n 0.17746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_254_n 0.0120212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_255_n 0.0124232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_110_47#_c_290_n 0.00249699f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_28 VPB N_A1_M1007_g 0.0238758f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_29 VPB A1 0.00751527f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_A2_M1006_g 0.0182297f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_31 VPB A2 0.00127568f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_32 VPB N_A2_c_73_n 0.00694058f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.295
cc_33 VPB N_A2_c_74_n 0.00652963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A3_M1002_g 0.0224959f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_35 VPB A3 0.00763759f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_36 VPB N_A3_c_116_n 0.0129854f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.375
cc_37 VPB N_B1_M1000_g 0.0287944f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_38 VPB N_B1_c_152_n 0.0148751f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.375
cc_39 VPB N_VPWR_c_179_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_40 VPB N_VPWR_c_180_n 0.0483776f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_41 VPB N_VPWR_c_181_n 0.0494394f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.375
cc_42 VPB N_VPWR_c_182_n 0.0454035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_183_n 0.00497181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_184_n 0.0129628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_178_n 0.0539931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB Y 0.00124246f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.375
cc_47 N_A1_M1007_g N_A2_M1006_g 0.0559127f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_48 N_A1_M1004_g N_A2_M1005_g 0.0234466f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_49 A1 N_A2_M1005_g 6.21404e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A1_M1007_g A2 0.00598368f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_51 N_A1_c_50_n N_A2_c_73_n 0.0559127f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_52 A1 N_A2_c_74_n 0.0335205f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_53 N_A1_c_50_n N_A2_c_74_n 0.00313912f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_54 N_A1_M1007_g N_VPWR_c_180_n 0.0230031f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_55 A1 N_VPWR_c_180_n 0.0246891f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A1_c_50_n N_VPWR_c_180_n 0.00131059f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_57 N_A1_M1007_g N_VPWR_c_182_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A1_M1007_g N_VPWR_c_178_n 0.00818711f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A1_M1004_g N_VGND_c_251_n 0.0173839f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_60 A1 N_VGND_c_251_n 0.0234206f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A1_c_50_n N_VGND_c_251_n 0.00213281f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_62 N_A1_M1004_g N_VGND_c_253_n 0.0082726f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_63 N_A1_M1004_g N_VGND_c_254_n 0.00486043f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_64 N_A1_M1004_g N_VGND_c_255_n 5.5187e-19 $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_65 N_A1_M1004_g N_A_110_47#_c_290_n 0.00101801f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_66 N_A2_M1006_g N_A3_M1002_g 0.0409859f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_67 A2 N_A3_M1002_g 0.00108129f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_68 N_A2_c_74_n N_A3_M1002_g 2.22431e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_69 N_A2_M1005_g N_A3_M1003_g 0.0138014f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_70 N_A2_c_73_n N_A3_c_116_n 0.020484f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_71 N_A2_c_74_n N_A3_c_116_n 2.84569e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_72 N_A2_M1006_g N_VPWR_c_180_n 0.00230539f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A2_M1006_g N_VPWR_c_182_n 0.00432378f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_74 A2 N_VPWR_c_182_n 0.0106998f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_75 N_A2_M1006_g N_VPWR_c_178_n 0.00709482f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_76 A2 N_VPWR_c_178_n 0.00961964f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_77 A2 A_110_367# 0.00111772f $X=0.635 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_78 N_A2_M1005_g N_Y_c_214_n 0.00393793f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_79 N_A2_M1006_g Y 0.0113017f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A2_M1005_g Y 0.00319154f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_81 A2 Y 0.0937009f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_82 N_A2_c_73_n Y 0.00400417f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_83 N_A2_c_74_n Y 0.0314596f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_84 N_A2_M1005_g N_VGND_c_251_n 6.85633e-19 $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_85 N_A2_M1005_g N_VGND_c_253_n 0.0039364f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_86 N_A2_M1005_g N_VGND_c_254_n 0.00332739f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_87 N_A2_M1005_g N_VGND_c_255_n 0.00866626f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_88 N_A2_M1005_g N_A_110_47#_c_292_n 0.0114816f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_89 N_A2_c_73_n N_A_110_47#_c_292_n 0.00227002f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_90 N_A2_c_74_n N_A_110_47#_c_292_n 0.0044014f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_91 N_A2_M1005_g N_A_110_47#_c_290_n 0.0105495f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_92 N_A2_c_73_n N_A_110_47#_c_290_n 0.00178872f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_93 N_A2_c_74_n N_A_110_47#_c_290_n 0.0169468f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_94 N_A3_M1002_g N_B1_M1000_g 0.00687701f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_95 A3 N_B1_M1000_g 0.0118649f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A3_M1003_g N_B1_M1001_g 0.0289889f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_97 N_A3_M1003_g N_B1_c_150_n 0.00241277f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_98 A3 N_B1_c_150_n 0.00884832f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A3_c_116_n N_B1_c_150_n 0.0197193f $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_100 A3 N_B1_c_151_n 0.00370329f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_101 A3 N_B1_c_152_n 0.0310999f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A3_M1002_g N_VPWR_c_182_n 0.00357668f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A3_M1002_g N_VPWR_c_178_n 0.0062997f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A3_M1003_g N_Y_c_213_n 0.011787f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_105 A3 N_Y_c_213_n 0.0555888f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_106 N_A3_c_116_n N_Y_c_213_n 0.0112829f $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_107 N_A3_M1002_g Y 0.0499951f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A3_M1003_g Y 0.0029961f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_109 A3 Y 0.0720425f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A3_c_116_n Y 0.0132091f $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_111 N_A3_M1003_g N_VGND_c_252_n 0.00360664f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_112 N_A3_M1003_g N_VGND_c_253_n 0.00449768f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_113 N_A3_M1003_g N_VGND_c_255_n 0.00942768f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_114 N_A3_M1003_g N_A_110_47#_c_292_n 0.0134675f $X=1.675 $Y=0.655 $X2=0 $Y2=0
cc_115 N_A3_c_116_n N_A_110_47#_c_292_n 4.30568e-19 $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_116 N_B1_M1000_g N_VPWR_c_181_n 0.00623768f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B1_c_151_n N_VPWR_c_181_n 0.00606277f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_118 N_B1_c_152_n N_VPWR_c_181_n 0.0100035f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_119 N_B1_M1000_g N_VPWR_c_182_n 0.0054895f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_M1000_g N_VPWR_c_178_n 0.0115226f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_121 N_B1_M1001_g N_Y_c_213_n 0.0151733f $X=2.175 $Y=0.655 $X2=0 $Y2=0
cc_122 N_B1_c_150_n N_Y_c_213_n 4.3418e-19 $X=2.167 $Y=1.46 $X2=0 $Y2=0
cc_123 N_B1_c_151_n N_Y_c_213_n 0.0113823f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_124 N_B1_c_152_n N_Y_c_213_n 0.011027f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_125 N_B1_M1000_g Y 0.0152337f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_M1001_g N_VGND_c_252_n 0.00549284f $X=2.175 $Y=0.655 $X2=0 $Y2=0
cc_127 N_B1_M1001_g N_VGND_c_253_n 0.0111876f $X=2.175 $Y=0.655 $X2=0 $Y2=0
cc_128 N_B1_M1001_g N_VGND_c_255_n 0.00105494f $X=2.175 $Y=0.655 $X2=0 $Y2=0
cc_129 N_B1_M1001_g N_A_110_47#_c_292_n 0.00214984f $X=2.175 $Y=0.655 $X2=0
+ $Y2=0
cc_130 N_B1_M1001_g N_A_110_47#_c_301_n 0.00477747f $X=2.175 $Y=0.655 $X2=0
+ $Y2=0
cc_131 N_VPWR_c_178_n A_110_367# 0.00333371f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_132 N_VPWR_c_178_n A_182_367# 0.00770351f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_133 N_VPWR_c_178_n N_Y_M1002_d 0.00518284f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_134 N_VPWR_c_180_n Y 0.00253549f $X=0.26 $Y=2.005 $X2=0 $Y2=0
cc_135 N_VPWR_c_182_n Y 0.0686999f $X=2.28 $Y=3.33 $X2=0 $Y2=0
cc_136 N_VPWR_c_178_n Y 0.0405789f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_137 A_182_367# Y 0.0226826f $X=0.91 $Y=1.835 $X2=2.41 $Y2=2.085
cc_138 N_Y_c_213_n N_VGND_M1005_d 0.00219492f $X=2.295 $Y=1.12 $X2=0 $Y2=0
cc_139 N_Y_c_214_n N_VGND_M1005_d 0.00272326f $X=1.35 $Y=1.12 $X2=0 $Y2=0
cc_140 N_Y_c_215_n N_VGND_c_252_n 0.0178111f $X=2.39 $Y=0.42 $X2=0 $Y2=0
cc_141 N_Y_M1001_d N_VGND_c_253_n 0.00371702f $X=2.25 $Y=0.235 $X2=0 $Y2=0
cc_142 N_Y_c_215_n N_VGND_c_253_n 0.0100304f $X=2.39 $Y=0.42 $X2=0 $Y2=0
cc_143 N_Y_c_213_n N_A_110_47#_M1003_d 0.00250873f $X=2.295 $Y=1.12 $X2=0 $Y2=0
cc_144 N_Y_c_213_n N_A_110_47#_c_292_n 0.0449987f $X=2.295 $Y=1.12 $X2=0 $Y2=0
cc_145 N_Y_c_214_n N_A_110_47#_c_292_n 0.013831f $X=1.35 $Y=1.12 $X2=0 $Y2=0
cc_146 N_Y_c_214_n N_A_110_47#_c_290_n 0.00300064f $X=1.35 $Y=1.12 $X2=0 $Y2=0
cc_147 N_VGND_c_253_n N_A_110_47#_M1004_d 0.00403327f $X=2.64 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_148 N_VGND_c_253_n N_A_110_47#_M1003_d 0.00300225f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_149 N_VGND_c_253_n N_A_110_47#_c_308_n 0.00691495f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_150 N_VGND_c_254_n N_A_110_47#_c_308_n 0.0120977f $X=0.945 $Y=0.22 $X2=0
+ $Y2=0
cc_151 N_VGND_M1005_d N_A_110_47#_c_292_n 0.0154407f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_152 N_VGND_c_252_n N_A_110_47#_c_292_n 0.00215102f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_153 N_VGND_c_253_n N_A_110_47#_c_292_n 0.00873487f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_154 N_VGND_c_254_n N_A_110_47#_c_292_n 0.00127509f $X=0.945 $Y=0.22 $X2=0
+ $Y2=0
cc_155 N_VGND_c_255_n N_A_110_47#_c_292_n 0.0433128f $X=1.625 $Y=0.22 $X2=0
+ $Y2=0
cc_156 N_VGND_c_252_n N_A_110_47#_c_301_n 0.0192194f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_157 N_VGND_c_253_n N_A_110_47#_c_301_n 0.0124653f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_158 N_VGND_c_253_n N_A_110_47#_c_290_n 0.00207489f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_159 N_VGND_c_254_n N_A_110_47#_c_290_n 8.24701e-19 $X=0.945 $Y=0.22 $X2=0
+ $Y2=0
