* File: sky130_fd_sc_lp__or2b_4.spice
* Created: Fri Aug 28 11:22:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2b_4.pex.spice"
.subckt sky130_fd_sc_lp__or2b_4  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B_N_M1005_g N_A_27_496#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=27.132 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1013 N_A_256_367#_M1013_d N_A_27_496#_M1013_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_256_367#_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1000_d N_A_256_367#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_256_367#_M1004_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1004_d N_A_256_367#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_256_367#_M1012_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_B_N_M1008_g N_A_27_496#_M1008_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_339_367# N_A_27_496#_M1009_g N_A_256_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_339_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=7.8012 NRS=7.8012 M=1 R=8.4 SA=75000.6 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1001_d N_A_256_367#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1764 PD=1.65 PS=1.54 NRD=9.3772 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_256_367#_M1006_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1006_d N_A_256_367#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_256_367#_M1011_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__or2b_4.pxi.spice"
*
.ends
*
*
