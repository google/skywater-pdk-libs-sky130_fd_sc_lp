* File: sky130_fd_sc_lp__dlygate4s50_1.pxi.spice
* Created: Wed Sep  2 09:50:11 2020
* 
x_PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A N_A_M1003_g N_A_M1002_g N_A_c_62_n
+ N_A_c_67_n A A N_A_c_64_n PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A
x_PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A_27_52# N_A_27_52#_M1003_s
+ N_A_27_52#_M1002_s N_A_27_52#_c_95_n N_A_27_52#_c_99_n N_A_27_52#_c_100_n
+ N_A_27_52#_c_101_n N_A_27_52#_c_96_n N_A_27_52#_c_97_n N_A_27_52#_c_115_n
+ N_A_27_52#_M1005_g N_A_27_52#_M1006_g
+ PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A_27_52#
x_PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A_288_52# N_A_288_52#_M1005_d
+ N_A_288_52#_M1006_d N_A_288_52#_M1004_g N_A_288_52#_M1007_g
+ N_A_288_52#_c_148_n N_A_288_52#_c_149_n N_A_288_52#_c_150_n
+ N_A_288_52#_c_151_n N_A_288_52#_c_155_n N_A_288_52#_c_156_n
+ N_A_288_52#_c_152_n PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A_288_52#
x_PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A_405_136# N_A_405_136#_M1004_s
+ N_A_405_136#_M1007_s N_A_405_136#_M1000_g N_A_405_136#_M1001_g
+ N_A_405_136#_c_198_n N_A_405_136#_c_203_n N_A_405_136#_c_199_n
+ N_A_405_136#_c_204_n N_A_405_136#_c_200_n N_A_405_136#_c_205_n
+ N_A_405_136#_c_201_n PM_SKY130_FD_SC_LP__DLYGATE4S50_1%A_405_136#
x_PM_SKY130_FD_SC_LP__DLYGATE4S50_1%VPWR N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_c_253_n N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_256_n VPWR
+ N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_252_n N_VPWR_c_260_n
+ PM_SKY130_FD_SC_LP__DLYGATE4S50_1%VPWR
x_PM_SKY130_FD_SC_LP__DLYGATE4S50_1%X N_X_M1000_d N_X_M1001_d X X X X X X X
+ N_X_c_283_n X X N_X_c_287_n PM_SKY130_FD_SC_LP__DLYGATE4S50_1%X
x_PM_SKY130_FD_SC_LP__DLYGATE4S50_1%VGND N_VGND_M1003_d N_VGND_M1004_d
+ N_VGND_c_304_n N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n VGND
+ N_VGND_c_308_n N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n
+ PM_SKY130_FD_SC_LP__DLYGATE4S50_1%VGND
cc_1 VNB N_A_M1003_g 0.0504374f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.47
cc_2 VNB N_A_c_62_n 0.0239894f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.695
cc_3 VNB A 0.0252844f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_64_n 0.0183476f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_5 VNB N_A_27_52#_c_95_n 0.0205357f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_6 VNB N_A_27_52#_c_96_n 0.0126078f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_7 VNB N_A_27_52#_c_97_n 0.0120797f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_8 VNB N_A_27_52#_M1005_g 0.126387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_288_52#_M1004_g 0.0550099f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_10 VNB N_A_288_52#_c_148_n 0.0177778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_288_52#_c_149_n 0.0225004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_288_52#_c_150_n 0.0415905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_288_52#_c_151_n 0.0105713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_288_52#_c_152_n 0.00394989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_405_136#_M1000_g 0.0268094f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_16 VNB N_A_405_136#_M1001_g 0.00154623f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A_405_136#_c_198_n 0.00170405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_405_136#_c_199_n 0.00313351f $X=-0.19 $Y=-0.245 $X2=0.565
+ $Y2=1.355
cc_19 VNB N_A_405_136#_c_200_n 0.00807403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_405_136#_c_201_n 0.0352273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_252_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB X 0.0283845f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_23 VNB N_X_c_283_n 0.0329417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 0.014713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_304_n 0.00643722f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_26 VNB N_VGND_c_305_n 0.0166487f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_VGND_c_306_n 0.0569179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_307_n 0.00532387f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_29 VNB N_VGND_c_308_n 0.0179296f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_30 VNB N_VGND_c_309_n 0.0191738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_310_n 0.243124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_311_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A_M1002_g 0.0486626f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.545
cc_34 VPB N_A_c_62_n 0.00312906f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.695
cc_35 VPB N_A_c_67_n 0.0183476f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.86
cc_36 VPB A 0.0136529f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_37 VPB N_A_27_52#_c_99_n 0.0220524f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_38 VPB N_A_27_52#_c_100_n 0.0137063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_52#_c_101_n 0.0109405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_52#_M1005_g 0.0978933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_288_52#_M1007_g 0.0586806f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_42 VPB N_A_288_52#_c_150_n 0.00783429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_288_52#_c_155_n 0.0125296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_288_52#_c_156_n 0.0183511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_405_136#_M1001_g 0.0259696f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_46 VPB N_A_405_136#_c_203_n 0.00170405f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_47 VPB N_A_405_136#_c_204_n 0.00164652f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.295
cc_48 VPB N_A_405_136#_c_205_n 0.00724414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_253_n 0.0274612f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_50 VPB N_VPWR_c_254_n 0.0315392f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_51 VPB N_VPWR_c_255_n 0.059762f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_52 VPB N_VPWR_c_256_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_53 VPB N_VPWR_c_257_n 0.0188373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_258_n 0.0190092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_252_n 0.111796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_260_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB X 0.00847673f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_58 VPB X 0.0492827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_X_c_287_n 0.0147304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_A_M1003_g N_A_27_52#_c_95_n 0.00955537f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_A_27_52#_c_99_n 0.00631563f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_62 N_A_M1002_g N_A_27_52#_c_100_n 0.0136775f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_63 N_A_c_67_n N_A_27_52#_c_100_n 0.00124917f $X=0.565 $Y=1.86 $X2=0 $Y2=0
cc_64 A N_A_27_52#_c_100_n 0.0257186f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_M1002_g N_A_27_52#_c_101_n 0.00349519f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_66 A N_A_27_52#_c_101_n 0.0280303f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_M1003_g N_A_27_52#_c_96_n 0.0108306f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_68 A N_A_27_52#_c_96_n 0.0251942f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_64_n N_A_27_52#_c_96_n 0.00126146f $X=0.565 $Y=1.355 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_A_27_52#_c_97_n 0.00435937f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_71 A N_A_27_52#_c_97_n 0.028939f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_A_27_52#_c_115_n 9.16519e-19 $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_73 N_A_M1002_g N_A_27_52#_c_115_n 9.16519e-19 $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_74 A N_A_27_52#_c_115_n 0.0394358f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_64_n N_A_27_52#_c_115_n 0.00220941f $X=0.565 $Y=1.355 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_A_27_52#_M1005_g 0.02206f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_77 N_A_M1002_g N_A_27_52#_M1005_g 0.0247334f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_78 A N_A_27_52#_M1005_g 0.00257785f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_c_64_n N_A_27_52#_M1005_g 0.0423481f $X=0.565 $Y=1.355 $X2=0 $Y2=0
cc_80 N_A_M1002_g N_VPWR_c_253_n 0.0039417f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_81 N_A_M1002_g N_VPWR_c_257_n 0.00442668f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_VPWR_c_252_n 0.0048347f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_83 N_A_M1003_g N_VGND_c_304_n 0.00327868f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_84 N_A_M1003_g N_VGND_c_308_n 0.00547602f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_VGND_c_310_n 0.00700251f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_86 N_A_27_52#_c_96_n N_A_288_52#_c_148_n 0.0164122f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_87 N_A_27_52#_c_115_n N_A_288_52#_c_148_n 0.0281345f $X=1.14 $Y=1.085 $X2=0
+ $Y2=0
cc_88 N_A_27_52#_M1005_g N_A_288_52#_c_148_n 0.022787f $X=1.19 $Y=0.47 $X2=0
+ $Y2=0
cc_89 N_A_27_52#_M1005_g N_A_288_52#_c_150_n 0.00405527f $X=1.19 $Y=0.47 $X2=0
+ $Y2=0
cc_90 N_A_27_52#_M1005_g N_A_288_52#_c_151_n 0.00947283f $X=1.19 $Y=0.47 $X2=0
+ $Y2=0
cc_91 N_A_27_52#_M1005_g N_A_288_52#_c_155_n 0.0096967f $X=1.19 $Y=0.47 $X2=0
+ $Y2=0
cc_92 N_A_27_52#_c_100_n N_A_288_52#_c_156_n 0.0143606f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_93 N_A_27_52#_c_115_n N_A_288_52#_c_156_n 0.0289074f $X=1.14 $Y=1.085 $X2=0
+ $Y2=0
cc_94 N_A_27_52#_M1005_g N_A_288_52#_c_156_n 0.022555f $X=1.19 $Y=0.47 $X2=0
+ $Y2=0
cc_95 N_A_27_52#_c_115_n N_A_288_52#_c_152_n 0.0227663f $X=1.14 $Y=1.085 $X2=0
+ $Y2=0
cc_96 N_A_27_52#_M1005_g N_A_288_52#_c_152_n 0.00411974f $X=1.19 $Y=0.47 $X2=0
+ $Y2=0
cc_97 N_A_27_52#_c_100_n N_VPWR_c_253_n 0.0243234f $X=0.975 $Y=2.117 $X2=0 $Y2=0
cc_98 N_A_27_52#_M1005_g N_VPWR_c_253_n 0.00683765f $X=1.19 $Y=0.47 $X2=0 $Y2=0
cc_99 N_A_27_52#_M1005_g N_VPWR_c_255_n 0.0145897f $X=1.19 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A_27_52#_c_99_n N_VPWR_c_257_n 0.00572829f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_101 N_A_27_52#_c_99_n N_VPWR_c_252_n 0.00940928f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_102 N_A_27_52#_M1005_g N_VPWR_c_252_n 0.0161157f $X=1.19 $Y=0.47 $X2=0 $Y2=0
cc_103 N_A_27_52#_c_96_n N_VGND_c_304_n 0.0244282f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_104 N_A_27_52#_M1005_g N_VGND_c_304_n 0.00342898f $X=1.19 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A_27_52#_M1005_g N_VGND_c_306_n 0.0183371f $X=1.19 $Y=0.47 $X2=0 $Y2=0
cc_106 N_A_27_52#_c_95_n N_VGND_c_308_n 0.0152237f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_107 N_A_27_52#_c_95_n N_VGND_c_310_n 0.0118277f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A_27_52#_c_96_n N_VGND_c_310_n 0.018948f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_109 N_A_27_52#_M1005_g N_VGND_c_310_n 0.0218268f $X=1.19 $Y=0.47 $X2=0 $Y2=0
cc_110 N_A_288_52#_M1004_g N_A_405_136#_M1000_g 0.0191704f $X=2.54 $Y=0.89 $X2=0
+ $Y2=0
cc_111 N_A_288_52#_c_150_n N_A_405_136#_M1001_g 0.0212525f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_112 N_A_288_52#_M1004_g N_A_405_136#_c_198_n 0.0352295f $X=2.54 $Y=0.89 $X2=0
+ $Y2=0
cc_113 N_A_288_52#_c_149_n N_A_405_136#_c_198_n 0.0277592f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_114 N_A_288_52#_M1007_g N_A_405_136#_c_203_n 0.0348505f $X=2.54 $Y=2.045
+ $X2=0 $Y2=0
cc_115 N_A_288_52#_c_149_n N_A_405_136#_c_203_n 0.0277592f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_116 N_A_288_52#_M1004_g N_A_405_136#_c_199_n 0.0060691f $X=2.54 $Y=0.89 $X2=0
+ $Y2=0
cc_117 N_A_288_52#_c_149_n N_A_405_136#_c_199_n 0.0203279f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_118 N_A_288_52#_c_149_n N_A_405_136#_c_204_n 0.00234001f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_119 N_A_288_52#_c_150_n N_A_405_136#_c_204_n 0.00462892f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_120 N_A_288_52#_M1004_g N_A_405_136#_c_200_n 0.019051f $X=2.54 $Y=0.89 $X2=0
+ $Y2=0
cc_121 N_A_288_52#_c_148_n N_A_405_136#_c_200_n 0.0304038f $X=1.597 $Y=1.385
+ $X2=0 $Y2=0
cc_122 N_A_288_52#_c_149_n N_A_405_136#_c_200_n 0.0291548f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_123 N_A_288_52#_c_150_n N_A_405_136#_c_200_n 0.00532229f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_124 N_A_288_52#_M1007_g N_A_405_136#_c_205_n 0.0137851f $X=2.54 $Y=2.045
+ $X2=0 $Y2=0
cc_125 N_A_288_52#_c_149_n N_A_405_136#_c_205_n 0.0284046f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_126 N_A_288_52#_c_150_n N_A_405_136#_c_205_n 0.00514979f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_127 N_A_288_52#_c_156_n N_A_405_136#_c_205_n 0.021975f $X=1.567 $Y=2.395
+ $X2=0 $Y2=0
cc_128 N_A_288_52#_M1004_g N_A_405_136#_c_201_n 0.0215925f $X=2.54 $Y=0.89 $X2=0
+ $Y2=0
cc_129 N_A_288_52#_c_149_n N_A_405_136#_c_201_n 2.28029e-19 $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_130 N_A_288_52#_M1007_g N_VPWR_c_254_n 0.00452277f $X=2.54 $Y=2.045 $X2=0
+ $Y2=0
cc_131 N_A_288_52#_c_155_n N_VPWR_c_255_n 0.0056234f $X=1.58 $Y=2.56 $X2=0 $Y2=0
cc_132 N_A_288_52#_c_155_n N_VPWR_c_252_n 0.00929046f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_133 N_A_288_52#_M1004_g N_VGND_c_305_n 0.00524017f $X=2.54 $Y=0.89 $X2=0
+ $Y2=0
cc_134 N_A_288_52#_M1004_g N_VGND_c_306_n 0.012617f $X=2.54 $Y=0.89 $X2=0 $Y2=0
cc_135 N_A_288_52#_c_151_n N_VGND_c_306_n 0.0145253f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_136 N_A_288_52#_M1004_g N_VGND_c_310_n 0.0151498f $X=2.54 $Y=0.89 $X2=0 $Y2=0
cc_137 N_A_288_52#_c_151_n N_VGND_c_310_n 0.0113149f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_138 N_A_405_136#_c_203_n N_VPWR_M1007_d 0.00246287f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_139 N_A_405_136#_M1001_g N_VPWR_c_254_n 0.016516f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_405_136#_c_203_n N_VPWR_c_254_n 0.0217748f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_141 N_A_405_136#_c_201_n N_VPWR_c_254_n 3.8937e-19 $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_142 N_A_405_136#_M1001_g N_VPWR_c_258_n 0.00486043f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_405_136#_M1001_g N_VPWR_c_252_n 0.00930006f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_405_136#_M1000_g X 0.00260428f $X=3.205 $Y=0.68 $X2=0 $Y2=0
cc_145 N_A_405_136#_M1001_g X 0.00292053f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_405_136#_c_199_n X 0.0327253f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_147 N_A_405_136#_c_204_n X 0.00710015f $X=3.032 $Y=1.825 $X2=0 $Y2=0
cc_148 N_A_405_136#_c_201_n X 0.00794767f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_149 N_A_405_136#_M1000_g N_X_c_283_n 0.00337221f $X=3.205 $Y=0.68 $X2=0 $Y2=0
cc_150 N_A_405_136#_c_199_n X 0.00398111f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_151 N_A_405_136#_M1001_g N_X_c_287_n 0.00335846f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_405_136#_c_203_n N_X_c_287_n 0.00755038f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_153 N_A_405_136#_c_204_n N_X_c_287_n 7.53353e-19 $X=3.032 $Y=1.825 $X2=0
+ $Y2=0
cc_154 N_A_405_136#_c_198_n N_VGND_M1004_d 6.59072e-19 $X=2.91 $Y=1.13 $X2=0
+ $Y2=0
cc_155 N_A_405_136#_c_199_n N_VGND_M1004_d 0.0018038f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_156 N_A_405_136#_M1000_g N_VGND_c_305_n 0.012902f $X=3.205 $Y=0.68 $X2=0
+ $Y2=0
cc_157 N_A_405_136#_c_198_n N_VGND_c_305_n 0.00508911f $X=2.91 $Y=1.13 $X2=0
+ $Y2=0
cc_158 N_A_405_136#_c_199_n N_VGND_c_305_n 0.0166857f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_159 N_A_405_136#_c_201_n N_VGND_c_305_n 4.81801e-19 $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_160 N_A_405_136#_c_200_n N_VGND_c_306_n 0.00527907f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_161 N_A_405_136#_M1000_g N_VGND_c_309_n 0.00465098f $X=3.205 $Y=0.68 $X2=0
+ $Y2=0
cc_162 N_A_405_136#_M1000_g N_VGND_c_310_n 0.0091589f $X=3.205 $Y=0.68 $X2=0
+ $Y2=0
cc_163 N_A_405_136#_c_200_n N_VGND_c_310_n 0.0100519f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_252_n N_X_M1001_d 0.00371702f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_c_258_n X 0.0289225f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VPWR_c_252_n X 0.0160565f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_167 N_X_c_283_n N_VGND_c_305_n 0.0234362f $X=3.42 $Y=0.42 $X2=0 $Y2=0
cc_168 N_X_c_283_n N_VGND_c_309_n 0.0296066f $X=3.42 $Y=0.42 $X2=0 $Y2=0
cc_169 N_X_c_283_n N_VGND_c_310_n 0.0160565f $X=3.42 $Y=0.42 $X2=0 $Y2=0
