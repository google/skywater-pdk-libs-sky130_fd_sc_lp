# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__iso1n_lp2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__iso1n_lp2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.165000 2.755000 1.495000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.515000 0.835000 1.845000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.525000 3.715000 0.985000 ;
        RECT 3.385000 2.025000 3.715000 3.065000 ;
        RECT 3.435000 0.985000 3.715000 2.025000 ;
    END
  END X
  PIN KAGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.755000 0.265000 3.075000 0.435000 ;
        RECT 0.755000 0.435000 1.385000 0.985000 ;
        RECT 2.445000 0.435000 3.075000 0.985000 ;
      LAYER mcon ;
        RECT 0.805000 0.470000 0.975000 0.640000 ;
        RECT 1.165000 0.470000 1.335000 0.640000 ;
        RECT 2.495000 0.470000 2.665000 0.640000 ;
        RECT 2.855000 0.470000 3.025000 0.640000 ;
      LAYER met1 ;
        RECT 0.070000 0.440000 3.770000 0.670000 ;
    END
  END KAGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.840000 3.415000 ;
        RECT 0.905000 2.025000 1.235000 3.245000 ;
        RECT 2.855000 2.025000 3.185000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.525000 0.445000 1.165000 ;
      RECT 0.115000 1.165000 1.500000 1.335000 ;
      RECT 0.115000 1.335000 0.285000 2.025000 ;
      RECT 0.115000 2.025000 0.625000 3.065000 ;
      RECT 1.170000 1.335000 1.500000 1.835000 ;
      RECT 1.695000 0.615000 2.055000 0.985000 ;
      RECT 1.695000 0.985000 1.865000 1.675000 ;
      RECT 1.695000 1.675000 3.265000 1.845000 ;
      RECT 1.695000 1.845000 2.295000 3.065000 ;
      RECT 2.935000 1.175000 3.265000 1.675000 ;
  END
END sky130_fd_sc_lp__iso1n_lp2
