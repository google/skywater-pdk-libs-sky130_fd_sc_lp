* File: sky130_fd_sc_lp__or3b_2.pex.spice
* Created: Wed Sep  2 10:31:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3B_2%C_N 3 5 7 8 12 13
c24 5 0 3.8122e-20 $X=0.67 $Y=1.725
c25 3 0 2.76376e-19 $X=0.505 $Y=0.865
r26 11 13 15.8553 $w=3.04e-07 $l=1e-07 $layer=POLY_cond $X=0.405 $Y=1.535
+ $X2=0.505 $Y2=1.535
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.51 $X2=0.405 $Y2=1.51
r28 8 12 5.51168 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.577
+ $X2=0.405 $Y2=1.577
r29 5 13 26.1612 $w=3.04e-07 $l=2.59711e-07 $layer=POLY_cond $X=0.67 $Y=1.725
+ $X2=0.505 $Y2=1.535
r30 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.67 $Y=1.725 $X2=0.67
+ $Y2=2.045
r31 1 13 19.2802 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.505 $Y=1.345
+ $X2=0.505 $Y2=1.535
r32 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.505 $Y=1.345
+ $X2=0.505 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_2%A_195_21# 1 2 3 10 12 15 17 19 22 26 27 29 30
+ 33 35 39 43 45 47
c103 39 0 5.72872e-20 $X=3.1 $Y=0.445
c104 27 0 1.13875e-19 $X=1.535 $Y=1.355
c105 22 0 1.25272e-20 $X=1.625 $Y=2.465
r106 49 50 46.0973 $w=2.98e-07 $l=2.85e-07 $layer=POLY_cond $X=1.195 $Y=1.352
+ $X2=1.48 $Y2=1.352
r107 45 46 16.4231 $w=2.08e-07 $l=2.8e-07 $layer=LI1_cond $X=2.207 $Y=0.87
+ $X2=2.207 $Y2=1.15
r108 41 47 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=0.955
+ $X2=3.125 $Y2=0.87
r109 41 43 48.5672 $w=2.78e-07 $l=1.18e-06 $layer=LI1_cond $X=3.125 $Y=0.955
+ $X2=3.125 $Y2=2.135
r110 37 47 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=0.785
+ $X2=3.125 $Y2=0.87
r111 37 39 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.125 $Y=0.785
+ $X2=3.125 $Y2=0.445
r112 36 45 1.9209 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=2.315 $Y=0.87
+ $X2=2.207 $Y2=0.87
r113 35 47 3.18746 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.985 $Y=0.87
+ $X2=3.125 $Y2=0.87
r114 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.985 $Y=0.87
+ $X2=2.315 $Y2=0.87
r115 31 45 4.82326 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.207 $Y=0.785
+ $X2=2.207 $Y2=0.87
r116 31 33 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.207 $Y=0.785
+ $X2=2.207 $Y2=0.445
r117 29 46 1.9209 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.1 $Y=1.15
+ $X2=2.207 $Y2=1.15
r118 29 30 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.1 $Y=1.15
+ $X2=1.72 $Y2=1.15
r119 27 52 14.557 $w=2.98e-07 $l=9e-08 $layer=POLY_cond $X=1.535 $Y=1.352
+ $X2=1.625 $Y2=1.352
r120 27 50 8.89597 $w=2.98e-07 $l=5.5e-08 $layer=POLY_cond $X=1.535 $Y=1.352
+ $X2=1.48 $Y2=1.352
r121 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.535
+ $Y=1.355 $X2=1.535 $Y2=1.355
r122 24 30 17.0466 $w=9.7e-08 $l=1.77482e-07 $layer=LI1_cond $X=1.58 $Y=1.235
+ $X2=1.72 $Y2=1.15
r123 24 26 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=1.58 $Y=1.235
+ $X2=1.58 $Y2=1.355
r124 20 52 18.8112 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=1.625 $Y=1.52
+ $X2=1.625 $Y2=1.352
r125 20 22 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.625 $Y=1.52
+ $X2=1.625 $Y2=2.465
r126 17 50 18.8112 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=1.48 $Y=1.185
+ $X2=1.48 $Y2=1.352
r127 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.48 $Y=1.185
+ $X2=1.48 $Y2=0.655
r128 13 49 18.8112 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=1.195 $Y=1.52
+ $X2=1.195 $Y2=1.352
r129 13 15 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.195 $Y=1.52
+ $X2=1.195 $Y2=2.465
r130 10 49 23.453 $w=2.98e-07 $l=2.28263e-07 $layer=POLY_cond $X=1.05 $Y=1.185
+ $X2=1.195 $Y2=1.352
r131 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.05 $Y=1.185
+ $X2=1.05 $Y2=0.655
r132 3 43 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.925 $X2=3.1 $Y2=2.135
r133 2 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.445
r134 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.235 $X2=2.22 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_2%A 3 7 9 10 14 15
c43 15 0 1.13875e-19 $X=2.075 $Y=1.51
c44 7 0 8.78014e-20 $X=2.165 $Y=2.135
c45 3 0 3.66459e-20 $X=2.005 $Y=0.445
r46 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.51
+ $X2=2.075 $Y2=1.675
r47 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.51
+ $X2=2.075 $Y2=1.345
r48 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.075
+ $Y=1.51 $X2=2.075 $Y2=1.51
r49 9 10 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.107 $Y=1.665
+ $X2=2.107 $Y2=2.035
r50 9 15 4.52224 $w=3.93e-07 $l=1.55e-07 $layer=LI1_cond $X=2.107 $Y=1.665
+ $X2=2.107 $Y2=1.51
r51 7 17 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.165 $Y=2.135
+ $X2=2.165 $Y2=1.675
r52 3 16 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.005 $Y=0.445
+ $X2=2.005 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_2%B 1 3 8 12 14 15 16 21 23
c46 14 0 9.29714e-20 $X=2.64 $Y=1.295
c47 12 0 5.72872e-20 $X=2.525 $Y=0.84
r48 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.29
+ $X2=2.615 $Y2=1.455
r49 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.29
+ $X2=2.615 $Y2=1.125
r50 15 16 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=1.665
+ $X2=2.645 $Y2=2.035
r51 14 15 12.7108 $w=3.38e-07 $l=3.75e-07 $layer=LI1_cond $X=2.645 $Y=1.29
+ $X2=2.645 $Y2=1.665
r52 14 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=1.29 $X2=2.615 $Y2=1.29
r53 10 12 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.435 $Y=0.84
+ $X2=2.525 $Y2=0.84
r54 8 24 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.525 $Y=2.135
+ $X2=2.525 $Y2=1.455
r55 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.525 $Y=0.915
+ $X2=2.525 $Y2=0.84
r56 4 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.525 $Y=0.915
+ $X2=2.525 $Y2=1.125
r57 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=0.765
+ $X2=2.435 $Y2=0.84
r58 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.435 $Y=0.765
+ $X2=2.435 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_2%A_33_131# 1 2 7 9 13 15 18 22 26 28 29 31 32
+ 36 43 46
c85 36 0 8.78014e-20 $X=2.65 $Y=2.88
c86 31 0 1.25272e-20 $X=0.84 $Y=1.92
r87 42 43 8.10674 $w=5.38e-07 $l=9e-08 $layer=LI1_cond $X=0.84 $Y=2.19 $X2=0.93
+ $Y2=2.19
r88 40 42 8.5276 $w=5.38e-07 $l=3.85e-07 $layer=LI1_cond $X=0.455 $Y=2.19
+ $X2=0.84 $Y2=2.19
r89 37 46 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=2.65 $Y=2.88
+ $X2=2.885 $Y2=2.88
r90 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=2.88 $X2=2.65 $Y2=2.88
r91 34 36 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.65 $Y=2.46
+ $X2=2.65 $Y2=2.88
r92 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.485 $Y=2.375
+ $X2=2.65 $Y2=2.46
r93 32 43 101.449 $w=1.68e-07 $l=1.555e-06 $layer=LI1_cond $X=2.485 $Y=2.375
+ $X2=0.93 $Y2=2.375
r94 31 42 7.28118 $w=1.8e-07 $l=2.7e-07 $layer=LI1_cond $X=0.84 $Y=1.92 $X2=0.84
+ $Y2=2.19
r95 30 31 42.2071 $w=1.78e-07 $l=6.85e-07 $layer=LI1_cond $X=0.84 $Y=1.235
+ $X2=0.84 $Y2=1.92
r96 28 30 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.75 $Y=1.15
+ $X2=0.84 $Y2=1.235
r97 28 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.75 $Y=1.15
+ $X2=0.385 $Y2=1.15
r98 24 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.255 $Y=1.065
+ $X2=0.385 $Y2=1.15
r99 24 26 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=0.255 $Y=1.065
+ $X2=0.255 $Y2=0.865
r100 20 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.885 $Y=1.74
+ $X2=3.095 $Y2=1.74
r101 16 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.885 $Y=0.84
+ $X2=3.095 $Y2=0.84
r102 15 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.095 $Y=1.665
+ $X2=3.095 $Y2=1.74
r103 14 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.095 $Y=0.915
+ $X2=3.095 $Y2=0.84
r104 14 15 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.095 $Y=0.915
+ $X2=3.095 $Y2=1.665
r105 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=2.715
+ $X2=2.885 $Y2=2.88
r106 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.885 $Y=2.715
+ $X2=2.885 $Y2=2.135
r107 10 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=1.815
+ $X2=2.885 $Y2=1.74
r108 10 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.885 $Y=1.815
+ $X2=2.885 $Y2=2.135
r109 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=0.765
+ $X2=2.885 $Y2=0.84
r110 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.885 $Y=0.765
+ $X2=2.885 $Y2=0.445
r111 2 40 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.835 $X2=0.455 $Y2=2.055
r112 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.655 $X2=0.29 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_2%VPWR 1 2 9 11 15 17 18 19 30 31 34
r33 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r34 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r36 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=1.84 $Y2=3.33
r38 25 27 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 19 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 19 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 19 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 17 22 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 17 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.98 $Y2=3.33
r45 13 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=3.245
+ $X2=1.84 $Y2=3.33
r46 13 15 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.84 $Y=3.245
+ $X2=1.84 $Y2=2.765
r47 12 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=0.98 $Y2=3.33
r48 11 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=1.84 $Y2=3.33
r49 11 12 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=1.145 $Y2=3.33
r50 7 18 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.98 $Y=3.245 $X2=0.98
+ $Y2=3.33
r51 7 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.98 $Y=3.245 $X2=0.98
+ $Y2=2.765
r52 2 15 600 $w=1.7e-07 $l=9.97547e-07 $layer=licon1_PDIFF $count=1 $X=1.7
+ $Y=1.835 $X2=1.84 $Y2=2.765
r53 1 9 600 $w=1.7e-07 $l=1.04089e-06 $layer=licon1_PDIFF $count=1 $X=0.745
+ $Y=1.835 $X2=0.98 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_2%X 1 2 8 11 13 14 21 29
c31 21 0 1.3868e-19 $X=1.265 $Y=0.42
c32 11 0 3.8122e-20 $X=1.41 $Y=1.98
c33 8 0 1.74342e-19 $X=1.185 $Y=1.815
r34 19 29 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=1.23 $Y=0.88
+ $X2=1.23 $Y2=0.925
r35 14 29 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=1.23 $Y=0.945
+ $X2=1.23 $Y2=0.925
r36 14 19 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=1.23 $Y=0.86 $X2=1.23
+ $Y2=0.88
r37 13 14 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.23 $Y=0.555
+ $X2=1.23 $Y2=0.86
r38 13 21 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=1.23 $Y=0.555
+ $X2=1.23 $Y2=0.42
r39 8 14 29.9161 $w=3.23e-07 $l=8.05e-07 $layer=LI1_cond $X=1.185 $Y=1.815
+ $X2=1.185 $Y2=1.01
r40 8 11 8.50163 $w=3.03e-07 $l=2.25e-07 $layer=LI1_cond $X=1.185 $Y=1.967
+ $X2=1.41 $Y2=1.967
r41 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.27
+ $Y=1.835 $X2=1.41 $Y2=1.98
r42 1 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.235 $X2=1.265 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_2%VGND 1 2 3 12 18 22 24 26 31 36 43 44 47 50
+ 53
r56 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r57 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 44 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r59 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r60 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.65
+ $Y2=0
r61 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=3.12
+ $Y2=0
r62 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r63 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r64 37 50 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.73
+ $Y2=0
r65 37 39 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.16
+ $Y2=0
r66 36 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.485 $Y=0 $X2=2.65
+ $Y2=0
r67 36 39 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.485 $Y=0 $X2=2.16
+ $Y2=0
r68 35 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r69 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r70 32 47 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.742
+ $Y2=0
r71 32 34 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.2
+ $Y2=0
r72 31 50 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.73
+ $Y2=0
r73 31 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.2
+ $Y2=0
r74 29 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r75 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r76 26 47 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.742
+ $Y2=0
r77 26 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r78 24 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r79 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r80 24 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r81 20 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0
r82 20 22 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0.445
r83 16 50 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.085 $X2=1.73
+ $Y2=0
r84 16 18 8.49927 $w=3.98e-07 $l=2.95e-07 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0.38
r85 12 14 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=0.742 $Y=0.38
+ $X2=0.742 $Y2=0.81
r86 10 47 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0
r87 10 12 9.06588 $w=3.73e-07 $l=2.95e-07 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0.38
r88 3 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.235 $X2=2.65 $Y2=0.445
r89 2 18 91 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=2 $X=1.555
+ $Y=0.235 $X2=1.79 $Y2=0.38
r90 1 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.655 $X2=0.72 $Y2=0.81
r91 1 12 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.655 $X2=0.815 $Y2=0.38
.ends

