* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxbp_lp D GATE VGND VNB VPB VPWR Q Q_N
X0 a_112_481# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VPWR a_798_47# a_1152_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_469_47# a_350_111# a_567_475# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_567_475# a_350_111# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_798_47# a_350_111# a_900_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_798_47# a_1133_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_27_111# D a_112_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 Q a_969_407# a_1403_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_1133_47# a_798_47# a_969_407# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_469_47# a_350_111# a_556_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_969_407# a_1597_361# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_1597_361# a_969_407# a_1662_131# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_720_47# a_469_47# a_798_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_114_111# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_1662_131# a_1863_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_1863_367# a_1662_131# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_27_111# D a_114_111# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 Q a_969_407# a_1418_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VGND a_27_111# a_720_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_927_519# a_969_407# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_900_47# a_969_407# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_741_475# a_350_111# a_798_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_1152_361# a_798_47# a_969_407# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VGND GATE a_272_111# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_1860_53# a_1662_131# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 VGND a_969_407# a_1584_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR GATE a_278_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1418_361# a_969_407# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VPWR a_27_111# a_741_475# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_1403_47# a_969_407# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 a_798_47# a_469_47# a_927_519# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_272_111# GATE a_350_111# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_556_47# a_350_111# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1584_131# a_969_407# a_1662_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_278_481# GATE a_350_111# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 VGND a_1662_131# a_1860_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
