* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor3_1 A B C VGND VNB VPB VPWR X
X0 a_355_451# B a_1090_373# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_1090_373# a_754_367# a_354_109# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_354_109# B a_1090_373# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 X a_81_259# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND a_871_373# a_1090_373# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_81_259# a_244_137# a_354_109# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 VPWR a_871_373# a_1090_373# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_871_373# a_754_367# a_354_109# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 X a_81_259# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_355_451# C a_81_259# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 VPWR B a_754_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_871_373# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_871_373# a_754_367# a_355_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_354_109# C a_81_259# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 a_871_373# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_354_109# B a_871_373# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VGND C a_244_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR C a_244_137# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_81_259# a_244_137# a_355_451# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_1090_373# a_754_367# a_355_451# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_355_451# B a_871_373# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 VGND B a_754_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
