* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o211a_0 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_80_21# A2 a_340_485# VPB phighvt w=640000u l=150000u
+  ad=3.744e+11p pd=3.73e+06u as=1.344e+11p ps=1.7e+06u
M1001 a_257_47# A2 VGND VNB nshort w=420000u l=150000u
+  ad=2.415e+11p pd=2.83e+06u as=2.331e+11p ps=2.79e+06u
M1002 a_340_485# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=4.096e+11p ps=3.84e+06u
M1003 VGND a_80_21# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 a_520_47# B1 a_257_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 VPWR a_80_21# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.872e+11p ps=2.49e+06u
M1006 a_80_21# C1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A1 a_257_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_80_21# C1 a_520_47# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 VPWR B1 a_80_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
