* File: sky130_fd_sc_lp__fa_0.pex.spice
* Created: Fri Aug 28 10:34:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FA_0%A 3 7 10 11 13 16 18 21 22 23 26 29 30 34 39 40
+ 41 43 44 49 51 52 53 61 62
c174 62 0 1.57483e-19 $X=2.785 $Y=1.665
c175 49 0 1.06385e-19 $X=0.955 $Y=1.86
c176 43 0 8.33712e-20 $X=6.665 $Y=1.555
r177 61 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.665
+ $X2=2.785 $Y2=1.83
r178 61 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.665
+ $X2=2.785 $Y2=1.5
r179 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=1.665 $X2=2.785 $Y2=1.665
r180 53 62 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.695
+ $X2=2.785 $Y2=1.695
r181 52 53 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.695
+ $X2=2.64 $Y2=1.695
r182 51 52 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.695
+ $X2=2.16 $Y2=1.695
r183 49 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.86
+ $X2=0.955 $Y2=2.025
r184 49 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.86
+ $X2=0.955 $Y2=1.695
r185 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=1.86 $X2=0.955 $Y2=1.86
r186 45 51 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=1.695
+ $X2=1.68 $Y2=1.695
r187 44 48 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=1.695
+ $X2=0.995 $Y2=1.86
r188 44 45 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.695
+ $X2=1.12 $Y2=1.695
r189 42 43 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.665 $Y=1.405
+ $X2=6.665 $Y2=1.555
r190 39 43 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=6.66 $Y=2.495 $X2=6.66
+ $Y2=1.555
r191 37 39 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.66 $Y=3.075
+ $X2=6.66 $Y2=2.495
r192 34 42 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=6.64 $Y=0.515
+ $X2=6.64 $Y2=1.405
r193 31 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.865 $Y=3.15
+ $X2=4.79 $Y2=3.15
r194 30 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.585 $Y=3.15
+ $X2=6.66 $Y2=3.075
r195 30 31 881.957 $w=1.5e-07 $l=1.72e-06 $layer=POLY_cond $X=6.585 $Y=3.15
+ $X2=4.865 $Y2=3.15
r196 26 29 866.574 $w=1.5e-07 $l=1.69e-06 $layer=POLY_cond $X=4.79 $Y=0.805
+ $X2=4.79 $Y2=2.495
r197 24 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=3.075
+ $X2=4.79 $Y2=3.15
r198 24 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.79 $Y=3.075
+ $X2=4.79 $Y2=2.495
r199 22 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.715 $Y=3.15
+ $X2=4.79 $Y2=3.15
r200 22 23 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=4.715 $Y=3.15
+ $X2=3.415 $Y2=3.15
r201 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.34 $Y=3.075
+ $X2=3.415 $Y2=3.15
r202 20 21 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.34 $Y=2.55
+ $X2=3.34 $Y2=3.075
r203 19 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.92 $Y=2.475
+ $X2=2.845 $Y2=2.475
r204 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.265 $Y=2.475
+ $X2=3.34 $Y2=2.55
r205 18 19 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=3.265 $Y=2.475
+ $X2=2.92 $Y2=2.475
r206 16 63 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.855 $Y=0.805
+ $X2=2.855 $Y2=1.5
r207 11 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.845 $Y=2.55
+ $X2=2.845 $Y2=2.475
r208 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.845 $Y=2.55
+ $X2=2.845 $Y2=2.87
r209 10 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.845 $Y=2.4
+ $X2=2.845 $Y2=2.475
r210 10 64 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.845 $Y=2.4
+ $X2=2.845 $Y2=1.83
r211 7 58 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.045 $Y=0.805
+ $X2=1.045 $Y2=1.695
r212 3 59 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=1.015 $Y=2.87
+ $X2=1.015 $Y2=2.025
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%B 3 7 11 16 20 24 28 30 32 34 35 36 39 43 44 48
+ 49 53 54 55 63
c165 36 0 1.06385e-19 $X=3.13 $Y=2.155
c166 35 0 1.57483e-19 $X=2.32 $Y=1.275
c167 30 0 9.29792e-20 $X=6.12 $Y=2.125
c168 28 0 9.10247e-20 $X=6.12 $Y=0.805
c169 3 0 3.61849e-20 $X=1.405 $Y=0.805
r170 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.21
+ $Y=1.96 $X2=6.21 $Y2=1.96
r171 55 70 1.58771 $w=5.63e-07 $l=7.5e-08 $layer=LI1_cond $X=6.292 $Y=2.035
+ $X2=6.292 $Y2=1.96
r172 54 78 2.39216 $w=4.48e-07 $l=9e-08 $layer=LI1_cond $X=6.35 $Y=1.665
+ $X2=6.35 $Y2=1.755
r173 53 54 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.665
r174 48 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.31 $Y=1.84
+ $X2=4.31 $Y2=2.005
r175 48 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.31 $Y=1.84
+ $X2=4.31 $Y2=1.675
r176 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.31
+ $Y=1.84 $X2=4.31 $Y2=1.84
r177 45 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=1.84
+ $X2=3.215 $Y2=1.84
r178 45 47 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.3 $Y=1.84
+ $X2=4.31 $Y2=1.84
r179 44 70 2.54034 $w=5.63e-07 $l=1.2e-07 $layer=LI1_cond $X=6.292 $Y=1.84
+ $X2=6.292 $Y2=1.96
r180 44 78 2.32906 $w=5.63e-07 $l=8.5e-08 $layer=LI1_cond $X=6.292 $Y=1.84
+ $X2=6.292 $Y2=1.755
r181 44 47 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=6.01 $Y=1.84
+ $X2=4.31 $Y2=1.84
r182 43 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=2.235
+ $X2=2.395 $Y2=2.4
r183 43 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=2.235
+ $X2=2.395 $Y2=2.07
r184 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=2.235 $X2=2.395 $Y2=2.235
r185 39 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=2.155
+ $X2=1.495 $Y2=2.32
r186 39 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=2.155
+ $X2=1.495 $Y2=1.99
r187 38 42 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=1.495 $Y=2.155
+ $X2=2.395 $Y2=2.155
r188 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=2.155 $X2=1.495 $Y2=2.155
r189 36 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.215 $Y=2.155
+ $X2=3.215 $Y2=1.84
r190 36 42 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=3.13 $Y=2.155
+ $X2=2.395 $Y2=2.155
r191 35 63 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.335 $Y=1.275
+ $X2=2.335 $Y2=2.07
r192 34 35 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.32 $Y=1.125
+ $X2=2.32 $Y2=1.275
r193 30 69 38.8824 $w=2.71e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.12 $Y=2.125
+ $X2=6.21 $Y2=1.96
r194 30 32 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.12 $Y=2.125
+ $X2=6.12 $Y2=2.495
r195 26 69 76.233 $w=2.71e-07 $l=4.17582e-07 $layer=POLY_cond $X=6.12 $Y=1.585
+ $X2=6.21 $Y2=1.96
r196 26 28 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.12 $Y=1.585
+ $X2=6.12 $Y2=0.805
r197 24 67 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=4.26 $Y=2.495
+ $X2=4.26 $Y2=2.005
r198 20 66 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=4.26 $Y=0.805
+ $X2=4.26 $Y2=1.675
r199 16 64 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.375 $Y=2.87 $X2=2.375
+ $Y2=2.4
r200 11 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.305 $Y=0.805
+ $X2=2.305 $Y2=1.125
r201 7 61 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.405 $Y=2.87
+ $X2=1.405 $Y2=2.32
r202 3 60 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=1.405 $Y=0.805
+ $X2=1.405 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%CIN 3 7 11 15 19 23 25 28 33 34 35 37 44 46
r120 44 55 3.47578 $w=3.51e-07 $l=1e-07 $layer=LI1_cond $X=3.612 $Y=1.375
+ $X2=3.612 $Y2=1.475
r121 44 53 2.08547 $w=3.51e-07 $l=6e-08 $layer=LI1_cond $X=3.612 $Y=1.375
+ $X2=3.612 $Y2=1.315
r122 43 46 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.6 $Y=1.375
+ $X2=3.83 $Y2=1.375
r123 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=1.375 $X2=3.6 $Y2=1.375
r124 37 53 0.695157 $w=3.51e-07 $l=2e-08 $layer=LI1_cond $X=3.612 $Y=1.295
+ $X2=3.612 $Y2=1.315
r125 34 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.67 $Y=1.46
+ $X2=5.67 $Y2=1.625
r126 34 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.67 $Y=1.46
+ $X2=5.67 $Y2=1.295
r127 33 35 7.25604 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.67 $Y=1.44
+ $X2=5.505 $Y2=1.44
r128 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.67
+ $Y=1.46 $X2=5.67 $Y2=1.46
r129 31 55 3.47043 $w=2.2e-07 $l=1.78e-07 $layer=LI1_cond $X=3.79 $Y=1.475
+ $X2=3.612 $Y2=1.475
r130 31 35 89.8382 $w=2.18e-07 $l=1.715e-06 $layer=LI1_cond $X=3.79 $Y=1.475
+ $X2=5.505 $Y2=1.475
r131 28 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.315
+ $X2=1.855 $Y2=1.48
r132 28 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.315
+ $X2=1.855 $Y2=1.15
r133 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.315 $X2=1.855 $Y2=1.315
r134 25 53 4.99104 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.435 $Y=1.315
+ $X2=3.612 $Y2=1.315
r135 25 27 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=3.435 $Y=1.315
+ $X2=1.855 $Y2=1.315
r136 23 50 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.73 $Y=2.495
+ $X2=5.73 $Y2=1.625
r137 19 49 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.65 $Y=0.805
+ $X2=5.65 $Y2=1.295
r138 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.54
+ $X2=3.83 $Y2=1.375
r139 13 15 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=3.83 $Y=1.54
+ $X2=3.83 $Y2=2.495
r140 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.21
+ $X2=3.83 $Y2=1.375
r141 9 11 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.83 $Y=1.21
+ $X2=3.83 $Y2=0.805
r142 7 41 712.745 $w=1.5e-07 $l=1.39e-06 $layer=POLY_cond $X=1.945 $Y=2.87
+ $X2=1.945 $Y2=1.48
r143 3 40 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.835 $Y=0.805
+ $X2=1.835 $Y2=1.15
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%A_80_225# 1 2 9 14 15 16 20 23 26 28 29 31 32
+ 34 35 37 40 41 45 50
c130 41 0 3.61849e-20 $X=0.597 $Y=1.21
c131 20 0 1.50979e-19 $X=5.22 $Y=0.805
r132 47 50 8.13695 $w=3.28e-07 $l=2.33e-07 $layer=LI1_cond $X=1.387 $Y=0.805
+ $X2=1.62 $Y2=0.805
r133 45 54 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.29
+ $X2=0.577 $Y2=1.455
r134 45 53 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.29
+ $X2=0.577 $Y2=1.125
r135 44 46 9.2829 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.597 $Y=1.29
+ $X2=0.597 $Y2=1.455
r136 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.29 $X2=0.59 $Y2=1.29
r137 41 44 4.32816 $w=2.03e-07 $l=8e-08 $layer=LI1_cond $X=0.597 $Y=1.21
+ $X2=0.597 $Y2=1.29
r138 39 47 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=1.387 $Y=0.97
+ $X2=1.387 $Y2=0.805
r139 39 40 6.7407 $w=2.63e-07 $l=1.55e-07 $layer=LI1_cond $X=1.387 $Y=0.97
+ $X2=1.387 $Y2=1.125
r140 35 37 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.23 $Y=2.87
+ $X2=1.685 $Y2=2.87
r141 34 35 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.145 $Y=2.705
+ $X2=1.23 $Y2=2.87
r142 33 34 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.145 $Y=2.365
+ $X2=1.145 $Y2=2.705
r143 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.28
+ $X2=1.145 $Y2=2.365
r144 31 32 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.06 $Y=2.28
+ $X2=0.7 $Y2=2.28
r145 30 41 1.83547 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=0.7 $Y=1.21
+ $X2=0.597 $Y2=1.21
r146 29 40 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=1.255 $Y=1.21
+ $X2=1.387 $Y2=1.125
r147 29 30 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.255 $Y=1.21
+ $X2=0.7 $Y2=1.21
r148 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.615 $Y=2.195
+ $X2=0.7 $Y2=2.28
r149 28 46 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.615 $Y=2.195
+ $X2=0.615 $Y2=1.455
r150 25 26 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.205 $Y=1.125
+ $X2=5.205 $Y2=1.275
r151 23 26 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=5.22 $Y=2.495
+ $X2=5.22 $Y2=1.275
r152 20 25 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.22 $Y=0.805
+ $X2=5.22 $Y2=1.125
r153 17 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.22 $Y=0.255
+ $X2=5.22 $Y2=0.805
r154 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.145 $Y=0.18
+ $X2=5.22 $Y2=0.255
r155 15 16 2284.37 $w=1.5e-07 $l=4.455e-06 $layer=POLY_cond $X=5.145 $Y=0.18
+ $X2=0.69 $Y2=0.18
r156 14 53 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.615 $Y=0.805
+ $X2=0.615 $Y2=1.125
r157 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.615 $Y=0.255
+ $X2=0.69 $Y2=0.18
r158 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.615 $Y=0.255
+ $X2=0.615 $Y2=0.805
r159 9 54 669.16 $w=1.5e-07 $l=1.305e-06 $layer=POLY_cond $X=0.475 $Y=2.76
+ $X2=0.475 $Y2=1.455
r160 2 37 600 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=2.66 $X2=1.685 $Y2=2.87
r161 1 50 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.595 $X2=1.62 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%A_1059_119# 1 2 9 12 14 16 21 23 27 32 34 36 37
+ 40
c74 36 0 8.33712e-20 $X=7.09 $Y=1.03
c75 23 0 1.50979e-19 $X=5.435 $Y=0.795
c76 21 0 2.1277e-19 $X=6.85 $Y=2.295
c77 14 0 9.29792e-20 $X=6.428 $Y=0.927
r78 37 41 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=7.102 $Y=1.03
+ $X2=7.102 $Y2=1.195
r79 37 40 51.3804 $w=3.55e-07 $l=1.95e-07 $layer=POLY_cond $X=7.102 $Y=1.03
+ $X2=7.102 $Y2=0.835
r80 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.09
+ $Y=1.03 $X2=7.09 $Y2=1.03
r81 33 36 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=6.85 $Y=1.022
+ $X2=7.09 $Y2=1.022
r82 33 34 6.47515 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=6.85 $Y=1.022
+ $X2=6.745 $Y2=1.022
r83 32 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.52 $Y=0.935
+ $X2=6.745 $Y2=0.935
r84 27 30 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.48 $Y=2.38 $X2=5.48
+ $Y2=2.5
r85 23 25 5.2456 $w=2.88e-07 $l=1.32e-07 $layer=LI1_cond $X=5.455 $Y=0.795
+ $X2=5.455 $Y2=0.927
r86 20 33 3.64154 $w=2.1e-07 $l=1.73e-07 $layer=LI1_cond $X=6.85 $Y=1.195
+ $X2=6.85 $Y2=1.022
r87 20 21 58.0952 $w=2.08e-07 $l=1.1e-06 $layer=LI1_cond $X=6.85 $Y=1.195
+ $X2=6.85 $Y2=2.295
r88 17 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=2.38
+ $X2=5.48 $Y2=2.38
r89 16 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.745 $Y=2.38
+ $X2=6.85 $Y2=2.295
r90 16 17 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=6.745 $Y=2.38
+ $X2=5.645 $Y2=2.38
r91 15 25 3.38853 $w=1.85e-07 $l=1.45e-07 $layer=LI1_cond $X=5.6 $Y=0.927
+ $X2=5.455 $Y2=0.927
r92 14 32 5.60801 $w=1.83e-07 $l=9.2e-08 $layer=LI1_cond $X=6.428 $Y=0.927
+ $X2=6.52 $Y2=0.927
r93 14 15 49.6393 $w=1.83e-07 $l=8.28e-07 $layer=LI1_cond $X=6.428 $Y=0.927
+ $X2=5.6 $Y2=0.927
r94 12 41 723 $w=1.5e-07 $l=1.41e-06 $layer=POLY_cond $X=7.205 $Y=2.605
+ $X2=7.205 $Y2=1.195
r95 9 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.07 $Y=0.515
+ $X2=7.07 $Y2=0.835
r96 2 30 600 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_PDIFF $count=1 $X=5.295
+ $Y=2.285 $X2=5.48 $Y2=2.5
r97 1 23 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.595 $X2=5.435 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%COUT 1 2 13 17 19 20 21 22
r17 21 22 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.205 $Y=2.035
+ $X2=0.205 $Y2=2.405
r18 20 21 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.205 $Y=1.665
+ $X2=0.205 $Y2=2.035
r19 19 20 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.205 $Y=1.295
+ $X2=0.205 $Y2=1.665
r20 18 22 4.56175 $w=2.38e-07 $l=9.5e-08 $layer=LI1_cond $X=0.205 $Y=2.5
+ $X2=0.205 $Y2=2.405
r21 17 18 3.89276 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=2.585
+ $X2=0.255 $Y2=2.5
r22 10 19 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.205 $Y=0.955
+ $X2=0.205 $Y2=1.295
r23 9 13 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.205 $Y=0.79
+ $X2=0.4 $Y2=0.79
r24 9 10 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.205 $Y=0.79
+ $X2=0.205 $Y2=0.955
r25 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.44 $X2=0.26 $Y2=2.585
r26 1 13 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.595 $X2=0.4 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%VPWR 1 2 3 4 5 18 22 26 30 34 36 38 43 51 56 61
+ 71 72 75 78 81 84 87
c94 5 0 1.21745e-19 $X=6.735 $Y=2.285
r95 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r96 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r98 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 72 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r101 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r102 69 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.135 $Y=3.33
+ $X2=6.97 $Y2=3.33
r103 69 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.135 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r105 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 65 68 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r107 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r108 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r109 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 62 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.69 $Y=3.33
+ $X2=4.525 $Y2=3.33
r111 62 64 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.69 $Y=3.33
+ $X2=5.04 $Y2=3.33
r112 61 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.97 $Y2=3.33
r113 61 67 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 60 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 57 81 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.607 $Y2=3.33
r117 57 59 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=4.08 $Y2=3.33
r118 56 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.36 $Y=3.33
+ $X2=4.525 $Y2=3.33
r119 56 59 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r120 55 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 55 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r123 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.61 $Y2=3.33
r124 52 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 51 81 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=3.607 $Y2=3.33
r126 51 54 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=3.12 $Y2=3.33
r127 50 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 47 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r132 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 44 75 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.742 $Y2=3.33
r134 44 46 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 43 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.61 $Y2=3.33
r136 43 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 41 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 38 75 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.742 $Y2=3.33
r140 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r141 36 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r142 36 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 32 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=3.245
+ $X2=6.97 $Y2=3.33
r144 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.97 $Y=3.245
+ $X2=6.97 $Y2=2.745
r145 28 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=3.245
+ $X2=4.525 $Y2=3.33
r146 28 30 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=4.525 $Y=3.245
+ $X2=4.525 $Y2=2.54
r147 24 81 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.607 $Y=3.245
+ $X2=3.607 $Y2=3.33
r148 24 26 31.6398 $w=2.73e-07 $l=7.55e-07 $layer=LI1_cond $X=3.607 $Y=3.245
+ $X2=3.607 $Y2=2.49
r149 20 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=3.245
+ $X2=2.61 $Y2=3.33
r150 20 22 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.61 $Y=3.245
+ $X2=2.61 $Y2=2.93
r151 16 75 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=3.33
r152 16 18 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=2.825
r153 5 34 600 $w=1.7e-07 $l=5.6542e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=2.285 $X2=6.97 $Y2=2.745
r154 4 30 600 $w=1.7e-07 $l=3.36861e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=2.285 $X2=4.525 $Y2=2.54
r155 3 26 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=2.285 $X2=3.615 $Y2=2.49
r156 2 22 600 $w=1.7e-07 $l=3.40734e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=2.66 $X2=2.61 $Y2=2.93
r157 1 18 600 $w=1.7e-07 $l=4.72546e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.44 $X2=0.745 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%A_404_532# 1 2 9 11 12 15
r28 13 15 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=3.085 $Y=2.66
+ $X2=3.085 $Y2=2.87
r29 11 13 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.945 $Y=2.575
+ $X2=3.085 $Y2=2.66
r30 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=2.575
+ $X2=2.275 $Y2=2.575
r31 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.135 $Y=2.66
+ $X2=2.275 $Y2=2.575
r32 7 9 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=2.135 $Y=2.66
+ $X2=2.135 $Y2=2.87
r33 2 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=2.66 $X2=3.06 $Y2=2.87
r34 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.02
+ $Y=2.66 $X2=2.16 $Y2=2.87
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%A_781_457# 1 2 9 11 12 15
r29 13 15 9.5026 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=5.002 $Y=2.265
+ $X2=5.002 $Y2=2.5
r30 11 13 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=4.86 $Y=2.18
+ $X2=5.002 $Y2=2.265
r31 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.86 $Y=2.18
+ $X2=4.19 $Y2=2.18
r32 7 12 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=4.052 $Y=2.265
+ $X2=4.19 $Y2=2.18
r33 7 9 9.84815 $w=2.73e-07 $l=2.35e-07 $layer=LI1_cond $X=4.052 $Y=2.265
+ $X2=4.052 $Y2=2.5
r34 2 15 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=2.285 $X2=5.005 $Y2=2.5
r35 1 9 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=2.285 $X2=4.045 $Y2=2.5
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%SUM 1 2 10 14 16 17 18 19 20 21
r17 20 21 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.45 $Y=2.405
+ $X2=7.45 $Y2=2.775
r18 19 20 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.45 $Y=2.035
+ $X2=7.45 $Y2=2.405
r19 18 19 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.45 $Y=1.665
+ $X2=7.45 $Y2=2.035
r20 16 17 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.47 $Y=0.925
+ $X2=7.47 $Y2=1.295
r21 15 17 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=7.47 $Y=1.405
+ $X2=7.47 $Y2=1.295
r22 14 18 4.57003 $w=2.88e-07 $l=1.15e-07 $layer=LI1_cond $X=7.45 $Y=1.55
+ $X2=7.45 $Y2=1.665
r23 14 15 6.01329 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=7.45 $Y=1.55
+ $X2=7.45 $Y2=1.405
r24 11 16 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=7.47 $Y=0.68
+ $X2=7.47 $Y2=0.925
r25 10 11 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=7.47 $Y=0.515
+ $X2=7.47 $Y2=0.68
r26 8 10 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.285 $Y=0.515
+ $X2=7.47 $Y2=0.515
r27 2 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.28
+ $Y=2.285 $X2=7.42 $Y2=2.43
r28 1 8 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.305 $X2=7.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%VGND 1 2 3 4 5 20 24 28 32 36 39 40 41 43 51 56
+ 69 70 73 76 79 82
r90 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r91 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r92 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r93 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r94 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r95 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r96 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r97 64 67 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r98 64 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r99 63 66 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r100 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r101 61 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.69 $Y=0 $X2=4.525
+ $Y2=0
r102 61 63 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.69 $Y=0 $X2=5.04
+ $Y2=0
r103 60 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r104 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r105 57 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=3.615
+ $Y2=0
r106 57 59 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=4.08
+ $Y2=0
r107 56 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.36 $Y=0 $X2=4.525
+ $Y2=0
r108 56 59 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.36 $Y=0 $X2=4.08
+ $Y2=0
r109 55 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r110 55 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r111 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r112 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.58
+ $Y2=0
r113 52 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.12 $Y2=0
r114 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.615
+ $Y2=0
r115 51 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.12
+ $Y2=0
r116 50 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r117 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r118 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r119 47 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r121 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r122 44 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.83
+ $Y2=0
r123 44 46 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.2
+ $Y2=0
r124 43 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.58
+ $Y2=0
r125 43 49 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.16 $Y2=0
r126 41 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r127 41 80 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r128 39 66 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.69 $Y=0 $X2=6.48
+ $Y2=0
r129 39 40 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.69 $Y=0 $X2=6.837
+ $Y2=0
r130 38 69 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.985 $Y=0
+ $X2=7.44 $Y2=0
r131 38 40 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.985 $Y=0
+ $X2=6.837 $Y2=0
r132 34 40 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.837 $Y=0.085
+ $X2=6.837 $Y2=0
r133 34 36 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=6.837 $Y=0.085
+ $X2=6.837 $Y2=0.515
r134 30 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=0.085
+ $X2=4.525 $Y2=0
r135 30 32 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.525 $Y=0.085
+ $X2=4.525 $Y2=0.74
r136 26 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=0.085
+ $X2=3.615 $Y2=0
r137 26 28 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.615 $Y=0.085
+ $X2=3.615 $Y2=0.795
r138 22 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0
r139 22 24 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0.615
r140 18 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0
r141 18 20 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0.805
r142 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.715
+ $Y=0.305 $X2=6.855 $Y2=0.515
r143 4 32 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.595 $X2=4.525 $Y2=0.74
r144 3 28 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=3.49
+ $Y=0.595 $X2=3.615 $Y2=0.795
r145 2 24 182 $w=1.7e-07 $l=2.09762e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.595 $X2=2.58 $Y2=0.615
r146 1 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.595 $X2=0.83 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%A_382_119# 1 2 7 10 15
r27 15 17 6.12235 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=3.075 $Y=0.805
+ $X2=3.075 $Y2=0.975
r28 10 12 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.08 $Y=0.805
+ $X2=2.08 $Y2=0.975
r29 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0.975
+ $X2=2.08 $Y2=0.975
r30 7 17 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.915 $Y=0.975
+ $X2=3.075 $Y2=0.975
r31 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.915 $Y=0.975
+ $X2=2.245 $Y2=0.975
r32 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.595 $X2=3.07 $Y2=0.805
r33 1 10 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.595 $X2=2.08 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__FA_0%A_781_119# 1 2 9 11 12 15
c26 9 0 8.70569e-20 $X=4.045 $Y=0.795
r27 13 15 9.4665 $w=2.78e-07 $l=2.3e-07 $layer=LI1_cond $X=5 $Y=1.025 $X2=5
+ $Y2=0.795
r28 11 13 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.86 $Y=1.11
+ $X2=5 $Y2=1.025
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.86 $Y=1.11
+ $X2=4.19 $Y2=1.11
r30 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.075 $Y=1.025
+ $X2=4.19 $Y2=1.11
r31 7 9 11.5244 $w=2.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.075 $Y=1.025
+ $X2=4.075 $Y2=0.795
r32 2 15 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.595 $X2=5.005 $Y2=0.795
r33 1 9 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.595 $X2=4.045 $Y2=0.795
.ends

