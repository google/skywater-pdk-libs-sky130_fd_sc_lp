* File: sky130_fd_sc_lp__fahcin_1.pex.spice
* Created: Fri Aug 28 10:35:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A 3 7 9 12 13
c35 12 0 1.59397e-19 $X=0.625 $Y=1.51
r36 12 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.51
+ $X2=0.61 $Y2=1.675
r37 12 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.51
+ $X2=0.61 $Y2=1.345
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.51 $X2=0.625 $Y2=1.51
r39 9 13 5.17764 $w=3.43e-07 $l=1.55e-07 $layer=LI1_cond $X=0.632 $Y=1.665
+ $X2=0.632 $Y2=1.51
r40 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=1.675
r41 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.505 $Y=0.655
+ $X2=0.505 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_29_47# 1 2 3 4 15 19 23 24 27 31 33 37 40
+ 41 42 44 45 46 47 48 51 53 54 58 59 60
c111 58 0 1.74527e-19 $X=1.195 $Y=1.37
c112 41 0 1.59397e-19 $X=1.172 $Y=1.392
r113 60 63 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=2.445 $Y=0.35
+ $X2=2.445 $Y2=0.51
r114 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.195
+ $Y=1.37 $X2=1.195 $Y2=1.37
r115 49 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.59 $Y=2.895
+ $X2=3.59 $Y2=2.53
r116 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=2.98
+ $X2=3.59 $Y2=2.895
r117 47 48 148.096 $w=1.68e-07 $l=2.27e-06 $layer=LI1_cond $X=3.505 $Y=2.98
+ $X2=1.235 $Y2=2.98
r118 45 60 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.32 $Y=0.35
+ $X2=2.445 $Y2=0.35
r119 45 46 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=2.32 $Y=0.35
+ $X2=1.155 $Y2=0.35
r120 44 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.895
+ $X2=1.235 $Y2=2.98
r121 44 59 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.15 $Y=2.895
+ $X2=1.15 $Y2=1.875
r122 42 59 7.70346 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=1.172 $Y=1.688
+ $X2=1.172 $Y2=1.875
r123 41 57 1.7631 $w=3.75e-07 $l=9.53677e-08 $layer=LI1_cond $X=1.172 $Y=1.392
+ $X2=1.257 $Y2=1.37
r124 41 42 9.09662 $w=3.73e-07 $l=2.96e-07 $layer=LI1_cond $X=1.172 $Y=1.392
+ $X2=1.172 $Y2=1.688
r125 39 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=0.435
+ $X2=1.155 $Y2=0.35
r126 39 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.07 $Y=0.435
+ $X2=1.07 $Y2=0.995
r127 38 53 2.87242 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.455 $Y=1.08
+ $X2=0.282 $Y2=1.08
r128 37 57 13.3008 $w=2.66e-07 $l=4.03708e-07 $layer=LI1_cond $X=0.985 $Y=1.08
+ $X2=1.257 $Y2=1.37
r129 37 40 5.48216 $w=2.66e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.985 $Y=1.08
+ $X2=1.07 $Y2=0.995
r130 37 38 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.985 $Y=1.08
+ $X2=0.455 $Y2=1.08
r131 33 35 33.7035 $w=2.63e-07 $l=7.75e-07 $layer=LI1_cond $X=0.242 $Y=2.125
+ $X2=0.242 $Y2=2.9
r132 31 54 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=0.242 $Y=2.092
+ $X2=0.242 $Y2=1.96
r133 31 33 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=0.242 $Y=2.092
+ $X2=0.242 $Y2=2.125
r134 29 53 3.6114 $w=2.57e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.195 $Y=1.165
+ $X2=0.282 $Y2=1.08
r135 29 54 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.195 $Y=1.165
+ $X2=0.195 $Y2=1.96
r136 25 53 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=0.282 $Y=0.995
+ $X2=0.282 $Y2=1.08
r137 25 27 18.8733 $w=3.43e-07 $l=5.65e-07 $layer=LI1_cond $X=0.282 $Y=0.995
+ $X2=0.282 $Y2=0.43
r138 23 58 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.195 $Y=1.71
+ $X2=1.195 $Y2=1.37
r139 23 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.71
+ $X2=1.195 $Y2=1.875
r140 22 58 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.205
+ $X2=1.195 $Y2=1.37
r141 19 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.285 $Y=2.535
+ $X2=1.285 $Y2=1.875
r142 15 22 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.205 $Y=0.755
+ $X2=1.205 $Y2=1.205
r143 4 51 600 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.895 $X2=3.59 $Y2=2.53
r144 3 35 400 $w=1.7e-07 $l=1.13519e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.29 $Y2=2.9
r145 3 33 400 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.29 $Y2=2.125
r146 2 63 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.365 $X2=2.485 $Y2=0.51
r147 1 27 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.29 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_439_47# 1 2 9 13 19 21 23 24 26 28 30 31
+ 34 35 38 39 40 44 45 46 47 52 56 58 64
c180 56 0 1.53495e-19 $X=3.965 $Y=1.285
c181 34 0 1.25487e-19 $X=3.615 $Y=1.54
c182 26 0 1.00898e-19 $X=5.685 $Y=2.445
c183 24 0 1.06994e-19 $X=5.685 $Y=1.595
c184 13 0 1.638e-19 $X=2.285 $Y=2.455
c185 9 0 9.51492e-20 $X=2.27 $Y=0.685
r186 63 65 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.375 $Y=1.54
+ $X2=3.4 $Y2=1.54
r187 63 64 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.375 $Y=1.54
+ $X2=3.3 $Y2=1.54
r188 58 61 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.88 $Y=1.935
+ $X2=4.88 $Y2=2.05
r189 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.545
+ $Y=1.43 $X2=5.545 $Y2=1.43
r190 50 52 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=5.507 $Y=1.85
+ $X2=5.507 $Y2=1.43
r191 49 52 19.4334 $w=2.53e-07 $l=4.3e-07 $layer=LI1_cond $X=5.507 $Y=1
+ $X2=5.507 $Y2=1.43
r192 48 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=1.935
+ $X2=4.88 $Y2=1.935
r193 47 50 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.38 $Y=1.935
+ $X2=5.507 $Y2=1.85
r194 47 48 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.38 $Y=1.935
+ $X2=5.045 $Y2=1.935
r195 45 49 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.38 $Y=0.915
+ $X2=5.507 $Y2=1
r196 45 46 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.38 $Y=0.915
+ $X2=5.045 $Y2=0.915
r197 42 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.88 $Y=0.83
+ $X2=5.045 $Y2=0.915
r198 42 44 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.88 $Y=0.83
+ $X2=4.88 $Y2=0.46
r199 41 44 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=4.88 $Y=0.435
+ $X2=4.88 $Y2=0.46
r200 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.715 $Y=0.35
+ $X2=4.88 $Y2=0.435
r201 39 40 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.715 $Y=0.35
+ $X2=4.05 $Y2=0.35
r202 38 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=1.2
+ $X2=3.965 $Y2=1.285
r203 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.965 $Y=0.435
+ $X2=4.05 $Y2=0.35
r204 37 38 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.965 $Y=0.435
+ $X2=3.965 $Y2=1.2
r205 35 65 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.615 $Y=1.54
+ $X2=3.4 $Y2=1.54
r206 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.54 $X2=3.615 $Y2=1.54
r207 32 56 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.615 $Y=1.285
+ $X2=3.965 $Y2=1.285
r208 32 34 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.615 $Y=1.37
+ $X2=3.615 $Y2=1.54
r209 28 53 68.0619 $w=3.27e-07 $l=4.43959e-07 $layer=POLY_cond $X=5.805 $Y=1.065
+ $X2=5.63 $Y2=1.43
r210 28 30 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.805 $Y=1.065
+ $X2=5.805 $Y2=0.635
r211 24 53 38.5818 $w=3.27e-07 $l=1.90526e-07 $layer=POLY_cond $X=5.685 $Y=1.595
+ $X2=5.63 $Y2=1.43
r212 24 26 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=5.685 $Y=1.595
+ $X2=5.685 $Y2=2.445
r213 21 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.375
+ $X2=3.4 $Y2=1.54
r214 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.4 $Y=1.375
+ $X2=3.4 $Y2=0.945
r215 17 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.705
+ $X2=3.375 $Y2=1.54
r216 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.375 $Y=1.705
+ $X2=3.375 $Y2=2.315
r217 16 31 5.30422 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=2.36 $Y=1.45
+ $X2=2.277 $Y2=1.45
r218 16 64 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.36 $Y=1.45 $X2=3.3
+ $Y2=1.45
r219 11 31 20.4101 $w=1.5e-07 $l=7.88987e-08 $layer=POLY_cond $X=2.285 $Y=1.525
+ $X2=2.277 $Y2=1.45
r220 11 13 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.285 $Y=1.525
+ $X2=2.285 $Y2=2.455
r221 7 31 20.4101 $w=1.5e-07 $l=7.84219e-08 $layer=POLY_cond $X=2.27 $Y=1.375
+ $X2=2.277 $Y2=1.45
r222 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.27 $Y=1.375
+ $X2=2.27 $Y2=0.685
r223 2 61 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=4.735
+ $Y=1.835 $X2=4.88 $Y2=2.05
r224 1 44 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.745
+ $Y=0.315 $X2=4.88 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%B 1 3 6 8 9 10 11 12 14 17 19 21 24 26 29
+ 33 35 38 40 41 42 43
c132 43 0 2.92216e-19 $X=5.04 $Y=1.295
c133 29 0 1.46968e-19 $X=5.095 $Y=0.735
c134 19 0 9.84507e-20 $X=4.51 $Y=2.92
c135 17 0 1.25487e-19 $X=4.095 $Y=0.945
c136 12 0 1.53495e-19 $X=4.065 $Y=2.845
r137 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.825
+ $Y=1.505 $X2=4.825 $Y2=1.505
r138 43 47 5.2481 $w=4.88e-07 $l=2.15e-07 $layer=LI1_cond $X=5.04 $Y=1.425
+ $X2=4.825 $Y2=1.425
r139 41 46 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.02 $Y=1.505
+ $X2=4.825 $Y2=1.505
r140 41 42 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.02 $Y=1.505
+ $X2=5.095 $Y2=1.505
r141 39 46 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=4.67 $Y=1.505
+ $X2=4.825 $Y2=1.505
r142 39 40 5.03009 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=4.67 $Y=1.505
+ $X2=4.59 $Y2=1.505
r143 35 36 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.065 $Y=2.92
+ $X2=4.065 $Y2=3.15
r144 31 42 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.095 $Y=1.67
+ $X2=5.095 $Y2=1.505
r145 31 33 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=5.095 $Y=1.67
+ $X2=5.095 $Y2=2.465
r146 27 42 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.095 $Y=1.34
+ $X2=5.095 $Y2=1.505
r147 27 29 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=5.095 $Y=1.34
+ $X2=5.095 $Y2=0.735
r148 26 40 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=4.595 $Y=1.34
+ $X2=4.59 $Y2=1.505
r149 25 26 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=4.595 $Y=0.255
+ $X2=4.595 $Y2=1.34
r150 23 40 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=4.585 $Y=1.67
+ $X2=4.59 $Y2=1.505
r151 23 24 602.5 $w=1.5e-07 $l=1.175e-06 $layer=POLY_cond $X=4.585 $Y=1.67
+ $X2=4.585 $Y2=2.845
r152 22 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.17 $Y=0.18
+ $X2=4.095 $Y2=0.18
r153 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.52 $Y=0.18
+ $X2=4.595 $Y2=0.255
r154 21 22 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.52 $Y=0.18
+ $X2=4.17 $Y2=0.18
r155 20 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.14 $Y=2.92
+ $X2=4.065 $Y2=2.92
r156 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.51 $Y=2.92
+ $X2=4.585 $Y2=2.845
r157 19 20 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.51 $Y=2.92
+ $X2=4.14 $Y2=2.92
r158 15 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.095 $Y=0.255
+ $X2=4.095 $Y2=0.18
r159 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.095 $Y=0.255
+ $X2=4.095 $Y2=0.945
r160 12 35 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.065 $Y=2.845
+ $X2=4.065 $Y2=2.92
r161 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.065 $Y=2.845
+ $X2=4.065 $Y2=2.315
r162 10 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=3.15
+ $X2=4.065 $Y2=3.15
r163 10 11 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=3.99 $Y=3.15
+ $X2=2.79 $Y2=3.15
r164 8 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.02 $Y=0.18
+ $X2=4.095 $Y2=0.18
r165 8 9 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=4.02 $Y=0.18
+ $X2=2.775 $Y2=0.18
r166 4 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.715 $Y=3.075
+ $X2=2.79 $Y2=3.15
r167 4 6 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.715 $Y=3.075
+ $X2=2.715 $Y2=2.455
r168 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=0.255
+ $X2=2.775 $Y2=0.18
r169 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.7 $Y=0.255 $X2=2.7
+ $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_555_73# 1 2 9 13 18 21 25 29 33 35 38 39
+ 40 42 43 44 47 48 51 52 53 55 58 59 61 64 65 66 68 69 71 72 75 78 79
c252 75 0 1.638e-19 $X=3.045 $Y=2.04
c253 71 0 1.75853e-20 $X=9.61 $Y=0.4
c254 68 0 1.10044e-19 $X=8.84 $Y=1.59
c255 59 0 1.57778e-19 $X=7.515 $Y=1.28
r256 77 78 8.86968 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=7.44 $Y=1.575
+ $X2=7.44 $Y2=1.745
r257 72 88 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.61 $Y=0.4
+ $X2=9.61 $Y2=0.565
r258 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.61
+ $Y=0.4 $X2=9.61 $Y2=0.4
r259 69 71 26.3141 $w=2.98e-07 $l=6.85e-07 $layer=LI1_cond $X=8.925 $Y=0.415
+ $X2=9.61 $Y2=0.415
r260 67 69 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=8.84 $Y=0.565
+ $X2=8.925 $Y2=0.415
r261 67 68 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=8.84 $Y=0.565
+ $X2=8.84 $Y2=1.59
r262 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.755 $Y=1.675
+ $X2=8.84 $Y2=1.59
r263 65 66 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=8.755 $Y=1.675
+ $X2=8.315 $Y2=1.675
r264 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.23 $Y=1.76
+ $X2=8.315 $Y2=1.675
r265 63 64 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=8.23 $Y=1.76
+ $X2=8.23 $Y2=2.895
r266 62 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=2.98
+ $X2=7.35 $Y2=2.98
r267 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.145 $Y=2.98
+ $X2=8.23 $Y2=2.895
r268 61 62 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.145 $Y=2.98
+ $X2=7.435 $Y2=2.98
r269 59 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.515 $Y=1.28
+ $X2=7.515 $Y2=1.115
r270 58 77 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=7.482 $Y=1.28
+ $X2=7.482 $Y2=1.575
r271 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.515
+ $Y=1.28 $X2=7.515 $Y2=1.28
r272 55 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=2.895
+ $X2=7.35 $Y2=2.98
r273 55 78 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=7.35 $Y=2.895
+ $X2=7.35 $Y2=1.745
r274 52 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.265 $Y=2.98
+ $X2=7.35 $Y2=2.98
r275 52 53 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=7.265 $Y=2.98
+ $X2=6.345 $Y2=2.98
r276 51 53 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.255 $Y=2.895
+ $X2=6.345 $Y2=2.98
r277 50 76 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=2.605
+ $X2=6.255 $Y2=2.52
r278 50 51 17.8687 $w=1.78e-07 $l=2.9e-07 $layer=LI1_cond $X=6.255 $Y=2.605
+ $X2=6.255 $Y2=2.895
r279 48 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.62
+ $X2=6.255 $Y2=1.785
r280 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.255
+ $Y=1.62 $X2=6.255 $Y2=1.62
r281 45 76 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=2.435
+ $X2=6.255 $Y2=2.52
r282 45 47 50.2172 $w=1.78e-07 $l=8.15e-07 $layer=LI1_cond $X=6.255 $Y=2.435
+ $X2=6.255 $Y2=1.62
r283 43 76 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.165 $Y=2.52
+ $X2=6.255 $Y2=2.52
r284 43 44 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=6.165 $Y=2.52
+ $X2=4.965 $Y2=2.52
r285 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.88 $Y=2.605
+ $X2=4.965 $Y2=2.52
r286 41 42 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.88 $Y=2.605
+ $X2=4.88 $Y2=2.895
r287 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.795 $Y=2.98
+ $X2=4.88 $Y2=2.895
r288 39 40 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.795 $Y=2.98
+ $X2=4.025 $Y2=2.98
r289 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.94 $Y=2.895
+ $X2=4.025 $Y2=2.98
r290 37 38 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.94 $Y=2.13
+ $X2=3.94 $Y2=2.895
r291 36 75 3.18746 $w=1.7e-07 $l=2.1543e-07 $layer=LI1_cond $X=3.27 $Y=2.045
+ $X2=3.075 $Y2=2.002
r292 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=2.045
+ $X2=3.94 $Y2=2.13
r293 35 36 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.855 $Y=2.045
+ $X2=3.27 $Y2=2.045
r294 31 75 3.351 $w=2.8e-07 $l=1.73491e-07 $layer=LI1_cond $X=3.185 $Y=1.875
+ $X2=3.075 $Y2=2.002
r295 31 33 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=3.185 $Y=1.875
+ $X2=3.185 $Y2=0.78
r296 27 75 3.351 $w=2.8e-07 $l=1.28e-07 $layer=LI1_cond $X=3.075 $Y=2.13
+ $X2=3.075 $Y2=2.002
r297 27 29 12.4109 $w=3.88e-07 $l=4.2e-07 $layer=LI1_cond $X=3.075 $Y=2.13
+ $X2=3.075 $Y2=2.55
r298 23 25 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=9.555 $Y=1.5
+ $X2=9.77 $Y2=1.5
r299 19 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.77 $Y=1.575
+ $X2=9.77 $Y2=1.5
r300 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=9.77 $Y=1.575
+ $X2=9.77 $Y2=2.395
r301 18 88 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.555 $Y=0.995
+ $X2=9.555 $Y2=0.565
r302 16 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.555 $Y=1.425
+ $X2=9.555 $Y2=1.5
r303 16 18 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.555 $Y=1.425
+ $X2=9.555 $Y2=0.995
r304 13 84 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.425 $Y=0.635
+ $X2=7.425 $Y2=1.115
r305 9 82 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.23 $Y=2.365
+ $X2=6.23 $Y2=1.785
r306 2 75 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=2.035 $X2=3.045 $Y2=2.04
r307 2 29 600 $w=1.7e-07 $l=6.29722e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=2.035 $X2=3.045 $Y2=2.55
r308 1 33 91 $w=1.7e-07 $l=5.85128e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.365 $X2=3.185 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_364_73# 1 2 3 4 13 15 16 17 19 20 21 22
+ 24 27 31 35 39 43 47 51 52 53 54 55 56 66 68 71 76 77 87 92
c242 68 0 1.78152e-19 $X=10.32 $Y=1.665
c243 66 0 1.57778e-19 $X=6.96 $Y=1.665
c244 54 0 1.91318e-19 $X=4.225 $Y=1.665
c245 31 0 2.81883e-20 $X=10.255 $Y=0.995
r246 87 88 2.18834 $w=4.46e-07 $l=8e-08 $layer=LI1_cond $X=1.95 $Y=1.492
+ $X2=2.03 $Y2=1.492
r247 76 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.27 $Y=1.65
+ $X2=10.27 $Y2=1.815
r248 76 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.27 $Y=1.65
+ $X2=10.27 $Y2=1.485
r249 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.27
+ $Y=1.65 $X2=10.27 $Y2=1.65
r250 68 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=1.665
+ $X2=10.32 $Y2=1.665
r251 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.665
r252 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.665
+ $X2=4.08 $Y2=1.665
r253 59 87 7.38565 $w=4.46e-07 $l=3.45847e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.95 $Y2=1.492
r254 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.665
r255 56 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=1.665
+ $X2=6.96 $Y2=1.665
r256 55 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.175 $Y=1.665
+ $X2=10.32 $Y2=1.665
r257 55 56 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=10.175 $Y=1.665
+ $X2=7.105 $Y2=1.665
r258 54 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.665
+ $X2=4.08 $Y2=1.665
r259 53 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=1.665
+ $X2=6.96 $Y2=1.665
r260 53 54 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=6.815 $Y=1.665
+ $X2=4.225 $Y2=1.665
r261 52 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=1.665
+ $X2=1.68 $Y2=1.665
r262 51 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r263 51 52 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=1.825 $Y2=1.665
r264 50 66 14.9727 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=6.975 $Y=1.395
+ $X2=6.975 $Y2=1.665
r265 48 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.975 $Y=1.23
+ $X2=6.975 $Y2=1.395
r266 48 71 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.975 $Y=1.23
+ $X2=6.975 $Y2=1.14
r267 47 50 7.89576 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=7.007 $Y=1.23
+ $X2=7.007 $Y2=1.395
r268 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.975
+ $Y=1.23 $X2=6.975 $Y2=1.23
r269 41 92 0.201461 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=4.355 $Y=1.55
+ $X2=4.355 $Y2=1.665
r270 41 43 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=4.355 $Y=1.55
+ $X2=4.355 $Y2=0.78
r271 37 92 0.651381 $w=2.28e-07 $l=1.3e-08 $layer=LI1_cond $X=4.342 $Y=1.665
+ $X2=4.355 $Y2=1.665
r272 37 63 13.1278 $w=2.28e-07 $l=2.62e-07 $layer=LI1_cond $X=4.342 $Y=1.665
+ $X2=4.08 $Y2=1.665
r273 37 39 10.8958 $w=2.73e-07 $l=2.6e-07 $layer=LI1_cond $X=4.342 $Y=1.78
+ $X2=4.342 $Y2=2.04
r274 33 88 4.12496 $w=2.5e-07 $l=2.88e-07 $layer=LI1_cond $X=2.03 $Y=1.78
+ $X2=2.03 $Y2=1.492
r275 33 35 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=2.03 $Y=1.78
+ $X2=2.03 $Y2=2.19
r276 31 78 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=10.255 $Y=0.995
+ $X2=10.255 $Y2=1.485
r277 27 79 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.2 $Y=2.395
+ $X2=10.2 $Y2=1.815
r278 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.45 $Y=1.835
+ $X2=7.45 $Y2=2.365
r279 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.375 $Y=1.76
+ $X2=7.45 $Y2=1.835
r280 20 21 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=7.375 $Y=1.76
+ $X2=7.14 $Y2=1.76
r281 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.065 $Y=1.685
+ $X2=7.14 $Y2=1.76
r282 19 74 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.065 $Y=1.685
+ $X2=7.065 $Y2=1.395
r283 16 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.81 $Y=1.14
+ $X2=6.975 $Y2=1.14
r284 16 17 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.81 $Y=1.14 $X2=6.31
+ $Y2=1.14
r285 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.235 $Y=1.065
+ $X2=6.31 $Y2=1.14
r286 13 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.235 $Y=1.065
+ $X2=6.235 $Y2=0.635
r287 4 39 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.14
+ $Y=1.895 $X2=4.29 $Y2=2.04
r288 3 35 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=2.035 $X2=2.07 $Y2=2.19
r289 2 43 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=4.17
+ $Y=0.625 $X2=4.315 $Y2=0.78
r290 1 87 182 $w=1.7e-07 $l=1.06802e-06 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.365 $X2=1.95 $Y2=1.37
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%CIN 3 5 7 8 10 12 14 15
c64 3 0 1.10044e-19 $X=7.995 $Y=2.445
r65 18 20 50.7821 $w=2.8e-07 $l=2.95e-07 $layer=POLY_cond $X=8.115 $Y=1.322
+ $X2=8.41 $Y2=1.322
r66 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.41
+ $Y=1.245 $X2=8.41 $Y2=1.245
r67 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.01 $Y=1.265
+ $X2=9.01 $Y2=0.735
r68 8 12 37.0107 $w=2.8e-07 $l=2.15e-07 $layer=POLY_cond $X=8.795 $Y=1.322
+ $X2=9.01 $Y2=1.322
r69 8 20 66.275 $w=2.8e-07 $l=3.85e-07 $layer=POLY_cond $X=8.795 $Y=1.322
+ $X2=8.41 $Y2=1.322
r70 8 10 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=8.795 $Y=1.415
+ $X2=8.795 $Y2=2.465
r71 5 18 17.3521 $w=1.5e-07 $l=2.42e-07 $layer=POLY_cond $X=8.115 $Y=1.08
+ $X2=8.115 $Y2=1.322
r72 5 7 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=8.115 $Y=1.08
+ $X2=8.115 $Y2=0.635
r73 1 18 20.6571 $w=2.8e-07 $l=2.97e-07 $layer=POLY_cond $X=7.995 $Y=1.565
+ $X2=8.115 $Y2=1.322
r74 1 3 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=7.995 $Y=1.565
+ $X2=7.995 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_1774_367# 1 2 3 12 16 19 20 27 30 32 33
+ 36 39 40 42 43
c98 43 0 8.91215e-20 $X=11.2 $Y=1.77
c99 36 0 1.0603e-20 $X=9.312 $Y=1.335
r100 43 47 16.4943 $w=2.63e-07 $l=9e-08 $layer=POLY_cond $X=11.2 $Y=1.77
+ $X2=11.29 $Y2=1.77
r101 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.2
+ $Y=1.77 $X2=11.2 $Y2=1.77
r102 38 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.525 $Y=2.9
+ $X2=10.69 $Y2=2.9
r103 38 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.525 $Y=2.9
+ $X2=10.36 $Y2=2.9
r104 33 36 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.205 $Y=1.94
+ $X2=9.205 $Y2=1.335
r105 32 33 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=9.067 $Y=2.105
+ $X2=9.067 $Y2=1.94
r106 29 42 8.00292 $w=3.43e-07 $l=3.1285e-07 $layer=LI1_cond $X=11.425 $Y=2.025
+ $X2=11.2 $Y2=1.815
r107 29 30 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=11.425 $Y=2.025
+ $X2=11.425 $Y2=2.895
r108 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.34 $Y=2.98
+ $X2=11.425 $Y2=2.895
r109 27 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.34 $Y=2.98
+ $X2=10.69 $Y2=2.98
r110 26 35 6.34366 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=9.29 $Y=2.98
+ $X2=9.067 $Y2=2.98
r111 26 39 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=9.29 $Y=2.98
+ $X2=10.36 $Y2=2.98
r112 20 36 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=9.312 $Y=1.143
+ $X2=9.312 $Y2=1.335
r113 20 22 3.2639 $w=3.85e-07 $l=1.03e-07 $layer=LI1_cond $X=9.312 $Y=1.143
+ $X2=9.312 $Y2=1.04
r114 19 35 2.41799 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=9.067 $Y=2.895
+ $X2=9.067 $Y2=2.98
r115 18 32 1.47616 $w=4.43e-07 $l=5.7e-08 $layer=LI1_cond $X=9.067 $Y=2.162
+ $X2=9.067 $Y2=2.105
r116 18 19 18.9829 $w=4.43e-07 $l=7.33e-07 $layer=LI1_cond $X=9.067 $Y=2.162
+ $X2=9.067 $Y2=2.895
r117 14 47 15.8942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.29 $Y=1.935
+ $X2=11.29 $Y2=1.77
r118 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.29 $Y=1.935
+ $X2=11.29 $Y2=2.595
r119 10 43 52.2319 $w=2.63e-07 $l=3.5812e-07 $layer=POLY_cond $X=10.915 $Y=1.605
+ $X2=11.2 $Y2=1.77
r120 10 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.915 $Y=1.605
+ $X2=10.915 $Y2=0.915
r121 3 38 600 $w=1.7e-07 $l=1.04253e-06 $layer=licon1_PDIFF $count=1 $X=10.275
+ $Y=1.975 $X2=10.525 $Y2=2.9
r122 2 35 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=8.87
+ $Y=1.835 $X2=9.01 $Y2=2.9
r123 2 32 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=8.87
+ $Y=1.835 $X2=9.01 $Y2=2.105
r124 1 22 182 $w=1.7e-07 $l=8.42912e-07 $layer=licon1_NDIFF $count=1 $X=9.085
+ $Y=0.315 $X2=9.34 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_1926_135# 1 2 7 9 12 15 17 19 20 21 23 24
+ 25 33 35 43
c97 35 0 8.91215e-20 $X=11.775 $Y=1.34
c98 17 0 1.78152e-19 $X=10.08 $Y=1.135
r99 39 43 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.775 $Y=1.51
+ $X2=11.99 $Y2=1.51
r100 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.775
+ $Y=1.51 $X2=11.775 $Y2=1.51
r101 35 38 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=11.775 $Y=1.34
+ $X2=11.775 $Y2=1.51
r102 30 33 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=9.84 $Y=2.12
+ $X2=9.985 $Y2=2.12
r103 24 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.61 $Y=1.34
+ $X2=11.775 $Y2=1.34
r104 24 25 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=11.61 $Y=1.34
+ $X2=11.135 $Y2=1.34
r105 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.05 $Y=1.255
+ $X2=11.135 $Y2=1.34
r106 22 23 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=11.05 $Y=0.435
+ $X2=11.05 $Y2=1.255
r107 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.965 $Y=0.35
+ $X2=11.05 $Y2=0.435
r108 20 21 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=10.965 $Y=0.35
+ $X2=10.205 $Y2=0.35
r109 17 26 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.08 $Y=1.22
+ $X2=9.84 $Y2=1.22
r110 17 19 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=10.08 $Y=1.135
+ $X2=10.08 $Y2=0.98
r111 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.08 $Y=0.435
+ $X2=10.205 $Y2=0.35
r112 16 19 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=10.08 $Y=0.435
+ $X2=10.08 $Y2=0.98
r113 15 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.84 $Y=2.035
+ $X2=9.84 $Y2=2.12
r114 14 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.84 $Y=1.305
+ $X2=9.84 $Y2=1.22
r115 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.84 $Y=1.305
+ $X2=9.84 $Y2=2.035
r116 10 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.99 $Y=1.675
+ $X2=11.99 $Y2=1.51
r117 10 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.99 $Y=1.675
+ $X2=11.99 $Y2=2.465
r118 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.775 $Y=1.345
+ $X2=11.775 $Y2=1.51
r119 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.775 $Y=1.345
+ $X2=11.775 $Y2=0.815
r120 2 33 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.845
+ $Y=1.975 $X2=9.985 $Y2=2.12
r121 1 19 182 $w=1.7e-07 $l=5.41433e-07 $layer=licon1_NDIFF $count=1 $X=9.63
+ $Y=0.675 $X2=10.04 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%VPWR 1 2 3 4 15 21 25 31 36 37 39 40 41 43
+ 61 67 68 71 74
c108 21 0 9.84507e-20 $X=5.31 $Y=2.95
r109 74 75 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r110 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 68 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r112 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r113 65 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.94 $Y=3.33
+ $X2=11.815 $Y2=3.33
r114 65 67 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=11.94 $Y=3.33
+ $X2=12.24 $Y2=3.33
r115 64 75 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=11.76 $Y2=3.33
r116 63 64 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 61 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.69 $Y=3.33
+ $X2=11.815 $Y2=3.33
r118 61 63 183.326 $w=1.68e-07 $l=2.81e-06 $layer=LI1_cond $X=11.69 $Y=3.33
+ $X2=8.88 $Y2=3.33
r119 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r120 59 60 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r121 56 59 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r122 56 57 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r124 53 54 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 51 54 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r126 51 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 50 53 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r128 50 51 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 48 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 46 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 43 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 43 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 41 60 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=8.4 $Y2=3.33
r136 41 57 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=5.52 $Y2=3.33
r137 39 59 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.495 $Y=3.33
+ $X2=8.4 $Y2=3.33
r138 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.495 $Y=3.33
+ $X2=8.58 $Y2=3.33
r139 38 63 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.665 $Y=3.33
+ $X2=8.88 $Y2=3.33
r140 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=3.33
+ $X2=8.58 $Y2=3.33
r141 36 53 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.145 $Y=3.33
+ $X2=5.04 $Y2=3.33
r142 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=3.33
+ $X2=5.31 $Y2=3.33
r143 35 56 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.475 $Y=3.33
+ $X2=5.52 $Y2=3.33
r144 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.475 $Y=3.33
+ $X2=5.31 $Y2=3.33
r145 31 34 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=11.815 $Y=2.02
+ $X2=11.815 $Y2=2.95
r146 29 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.815 $Y=3.245
+ $X2=11.815 $Y2=3.33
r147 29 34 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=11.815 $Y=3.245
+ $X2=11.815 $Y2=2.95
r148 25 28 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.58 $Y=2.105
+ $X2=8.58 $Y2=2.95
r149 23 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.58 $Y=3.245
+ $X2=8.58 $Y2=3.33
r150 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.58 $Y=3.245
+ $X2=8.58 $Y2=2.95
r151 19 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=3.245
+ $X2=5.31 $Y2=3.33
r152 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.31 $Y=3.245
+ $X2=5.31 $Y2=2.95
r153 15 18 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=0.72 $Y=2.22
+ $X2=0.72 $Y2=2.95
r154 13 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r155 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.95
r156 4 34 400 $w=1.7e-07 $l=1.03999e-06 $layer=licon1_PDIFF $count=1 $X=11.365
+ $Y=2.095 $X2=11.775 $Y2=2.95
r157 4 31 400 $w=1.7e-07 $l=4.45926e-07 $layer=licon1_PDIFF $count=1 $X=11.365
+ $Y=2.095 $X2=11.775 $Y2=2.02
r158 3 28 400 $w=1.7e-07 $l=1.23393e-06 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.945 $X2=8.58 $Y2=2.95
r159 3 25 400 $w=1.7e-07 $l=5.84551e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.945 $X2=8.58 $Y2=2.105
r160 2 21 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.835 $X2=5.31 $Y2=2.95
r161 1 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.95
r162 1 15 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_256_87# 1 2 3 4 15 17 19 20 24 26 27 28
+ 31 34 39
c83 34 0 1.74527e-19 $X=1.42 $Y=0.82
c84 28 0 9.51492e-20 $X=2.92 $Y=0.35
r85 34 36 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=1.46 $Y=0.82
+ $X2=1.46 $Y2=0.94
r86 29 31 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=3.575 $Y=0.435
+ $X2=3.575 $Y2=0.81
r87 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.45 $Y=0.35
+ $X2=3.575 $Y2=0.435
r88 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.45 $Y=0.35
+ $X2=2.92 $Y2=0.35
r89 26 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.835 $Y=0.855
+ $X2=2.835 $Y2=0.94
r90 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.835 $Y=0.435
+ $X2=2.92 $Y2=0.35
r91 25 26 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.835 $Y=0.435
+ $X2=2.835 $Y2=0.855
r92 22 24 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.5 $Y=2.545
+ $X2=2.5 $Y2=2.18
r93 21 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.5 $Y=0.94
+ $X2=2.835 $Y2=0.94
r94 21 24 40.3355 $w=3.28e-07 $l=1.155e-06 $layer=LI1_cond $X=2.5 $Y=1.025
+ $X2=2.5 $Y2=2.18
r95 19 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=2.63
+ $X2=2.5 $Y2=2.545
r96 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.335 $Y=2.63
+ $X2=1.665 $Y2=2.63
r97 18 36 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.585 $Y=0.94
+ $X2=1.46 $Y2=0.94
r98 17 21 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0.94
+ $X2=2.5 $Y2=0.94
r99 17 18 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.335 $Y=0.94
+ $X2=1.585 $Y2=0.94
r100 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.54 $Y=2.545
+ $X2=1.665 $Y2=2.63
r101 13 15 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=1.54 $Y=2.545
+ $X2=1.54 $Y2=2.385
r102 4 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=2.035 $X2=2.5 $Y2=2.18
r103 3 15 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=2.035 $X2=1.5 $Y2=2.385
r104 2 31 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.475
+ $Y=0.625 $X2=3.615 $Y2=0.81
r105 1 34 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.435 $X2=1.42 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_1152_389# 1 2 9 13 15
c30 15 0 1.07712e-19 $X=6 $Y=0.975
c31 13 0 3.92553e-20 $X=5.9 $Y=2.09
r32 13 15 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.9 $Y=2.09
+ $X2=5.9 $Y2=0.975
r33 7 15 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6 $Y=0.79 $X2=6
+ $Y2=0.975
r34 7 9 10.2785 $w=3.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6 $Y=0.79 $X2=6
+ $Y2=0.46
r35 2 13 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.76
+ $Y=1.945 $X2=5.9 $Y2=2.09
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.88
+ $Y=0.315 $X2=6.02 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%COUT 1 2 11 13 14 15 16 31
c38 13 0 1.06994e-19 $X=6.69 $Y=1.96
r39 30 31 2.47332 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.59
+ $X2=6.695 $Y2=0.59
r40 15 16 12.4308 $w=4.43e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=0.662
+ $X2=7.44 $Y2=0.662
r41 15 31 6.86286 $w=4.43e-07 $l=2.65e-07 $layer=LI1_cond $X=6.96 $Y=0.662
+ $X2=6.695 $Y2=0.662
r42 14 30 2.63543 $w=5.88e-07 $l=1.3e-07 $layer=LI1_cond $X=6.48 $Y=0.59
+ $X2=6.61 $Y2=0.59
r43 11 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=2.125
+ $X2=6.69 $Y2=1.96
r44 7 30 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.61 $Y=0.885
+ $X2=6.61 $Y2=0.59
r45 7 13 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=6.61 $Y=0.885
+ $X2=6.61 $Y2=1.96
r46 2 11 300 $w=1.7e-07 $l=4.66396e-07 $layer=licon1_PDIFF $count=2 $X=6.305
+ $Y=1.945 $X2=6.69 $Y2=2.125
r47 1 14 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=6.31
+ $Y=0.315 $X2=6.53 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_1500_63# 1 2 11 16 17 18
r33 17 18 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=7.88 $Y=1.925
+ $X2=7.88 $Y2=0.935
r34 16 17 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.79 $Y=2.09
+ $X2=7.79 $Y2=1.925
r35 9 18 7.30505 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.9 $Y=0.77 $X2=7.9
+ $Y2=0.935
r36 9 11 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.9 $Y=0.77 $X2=7.9
+ $Y2=0.615
r37 2 16 300 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=2 $X=7.525
+ $Y=1.945 $X2=7.78 $Y2=2.09
r38 1 11 182 $w=1.7e-07 $l=5.2915e-07 $layer=licon1_NDIFF $count=1 $X=7.5
+ $Y=0.315 $X2=7.9 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%A_1883_395# 1 2 3 10 14 17 18 24 26
r49 26 28 10.8156 $w=4.23e-07 $l=3.75e-07 $layer=LI1_cond $X=10.7 $Y=2.46
+ $X2=11.075 $Y2=2.46
r50 24 25 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=10.602 $Y=1.14
+ $X2=10.602 $Y2=1.305
r51 18 21 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=9.595 $Y=2.47
+ $X2=9.595 $Y2=2.55
r52 17 26 6.11956 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=10.7 $Y=2.205
+ $X2=10.7 $Y2=2.46
r53 17 25 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=10.7 $Y=2.205 $X2=10.7
+ $Y2=1.305
r54 12 24 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=10.602 $Y=1.123
+ $X2=10.602 $Y2=1.14
r55 12 14 10.8298 $w=3.63e-07 $l=3.43e-07 $layer=LI1_cond $X=10.602 $Y=1.123
+ $X2=10.602 $Y2=0.78
r56 11 18 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.72 $Y=2.47
+ $X2=9.595 $Y2=2.47
r57 10 26 6.9565 $w=4.23e-07 $l=8.9861e-08 $layer=LI1_cond $X=10.615 $Y=2.47
+ $X2=10.7 $Y2=2.46
r58 10 11 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=10.615 $Y=2.47
+ $X2=9.72 $Y2=2.47
r59 3 28 600 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=10.935
+ $Y=2.095 $X2=11.075 $Y2=2.46
r60 2 21 600 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=1 $X=9.415
+ $Y=1.975 $X2=9.555 $Y2=2.55
r61 1 24 182 $w=1.7e-07 $l=5.78619e-07 $layer=licon1_NDIFF $count=1 $X=10.33
+ $Y=0.675 $X2=10.585 $Y2=1.14
r62 1 14 182 $w=1.7e-07 $l=3.02985e-07 $layer=licon1_NDIFF $count=1 $X=10.33
+ $Y=0.675 $X2=10.585 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%SUM 1 2 7 8 9 10 11 12 13 37
r15 13 34 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=12.245 $Y=2.775
+ $X2=12.245 $Y2=2.9
r16 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.245 $Y=2.405
+ $X2=12.245 $Y2=2.775
r17 11 12 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=12.245 $Y=1.98
+ $X2=12.245 $Y2=2.405
r18 10 11 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=12.245 $Y=1.665
+ $X2=12.245 $Y2=1.98
r19 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.245 $Y=1.295
+ $X2=12.245 $Y2=1.665
r20 9 43 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=12.245 $Y=1.295
+ $X2=12.245 $Y2=1.075
r21 8 43 6.83074 $w=5.43e-07 $l=1.5e-07 $layer=LI1_cond $X=12.097 $Y=0.925
+ $X2=12.097 $Y2=1.075
r22 7 8 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=12.097 $Y=0.555
+ $X2=12.097 $Y2=0.925
r23 7 37 0.329196 $w=5.43e-07 $l=1.5e-08 $layer=LI1_cond $X=12.097 $Y=0.555
+ $X2=12.097 $Y2=0.54
r24 2 34 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=12.065
+ $Y=1.835 $X2=12.205 $Y2=2.9
r25 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.065
+ $Y=1.835 $X2=12.205 $Y2=1.98
r26 1 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.85
+ $Y=0.395 $X2=11.99 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCIN_1%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 47
+ 60 61 64 67 70
r113 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r114 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r115 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r116 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r117 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r118 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r119 55 58 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=11.28 $Y2=0
r120 55 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r121 54 57 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.88 $Y=0 $X2=11.28
+ $Y2=0
r122 54 55 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r123 52 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.575 $Y=0 $X2=8.41
+ $Y2=0
r124 52 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.575 $Y=0
+ $X2=8.88 $Y2=0
r125 51 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r126 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r127 48 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.555 $Y=0 $X2=5.39
+ $Y2=0
r128 48 50 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=5.555 $Y=0
+ $X2=7.92 $Y2=0
r129 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=8.41
+ $Y2=0
r130 47 50 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.245 $Y=0
+ $X2=7.92 $Y2=0
r131 46 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r132 45 46 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r133 43 46 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r134 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r135 42 45 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r136 42 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r137 40 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.72
+ $Y2=0
r138 40 42 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=1.2
+ $Y2=0
r139 39 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.39
+ $Y2=0
r140 39 45 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.04 $Y2=0
r141 37 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r142 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r143 34 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.72
+ $Y2=0
r144 34 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0
+ $X2=0.24 $Y2=0
r145 32 51 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=7.92 $Y2=0
r146 32 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=0 $X2=5.52
+ $Y2=0
r147 30 57 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=11.315 $Y=0
+ $X2=11.28 $Y2=0
r148 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.315 $Y=0
+ $X2=11.48 $Y2=0
r149 29 60 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=12.24 $Y2=0
r150 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=11.48 $Y2=0
r151 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.48 $Y=0.085
+ $X2=11.48 $Y2=0
r152 25 27 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.48 $Y=0.085
+ $X2=11.48 $Y2=0.54
r153 21 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0
r154 21 23 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0.595
r155 17 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.39 $Y=0.085
+ $X2=5.39 $Y2=0
r156 17 19 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.39 $Y=0.085
+ $X2=5.39 $Y2=0.47
r157 13 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r158 13 15 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.515
r159 4 27 91 $w=1.7e-07 $l=5.16769e-07 $layer=licon1_NDIFF $count=2 $X=10.99
+ $Y=0.595 $X2=11.48 $Y2=0.54
r160 3 23 182 $w=1.7e-07 $l=3.74166e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.315 $X2=8.41 $Y2=0.595
r161 2 19 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=5.17
+ $Y=0.315 $X2=5.39 $Y2=0.47
r162 1 15 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.235 $X2=0.72 $Y2=0.515
.ends

