* File: sky130_fd_sc_lp__a22o_m.spice
* Created: Wed Sep  2 09:22:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22o_m.pex.spice"
.subckt sky130_fd_sc_lp__a22o_m  VNB VPB A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_85_317#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=17.136 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1007 A_265_125# N_A2_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_85_317#_M1004_d N_A1_M1004_g A_265_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 A_445_125# N_B1_M1009_g N_A_85_317#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75001.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_B2_M1008_g A_445_125# VNB NSHORT L=0.15 W=0.42 AD=0.1764
+ AS=0.0441 PD=1.68 PS=0.63 NRD=44.28 NRS=14.28 M=1 R=2.8 SA=75002 SB=75000.3
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_85_317#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0924 AS=0.1113 PD=0.86 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_265_501#_M1005_d N_A2_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=65.6601 M=1 R=2.8
+ SA=75000.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_85_317#_M1000_d N_B1_M1000_g N_A_265_501#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1129 AS=0.0588 PD=0.97 PS=0.7 NRD=53.9386 NRS=0 M=1 R=2.8
+ SA=75001.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_265_501#_M1006_d N_B2_M1006_g N_A_85_317#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1129 PD=0.7 PS=0.97 NRD=0 NRS=56.2829 M=1 R=2.8
+ SA=75001.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_265_501#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a22o_m.pxi.spice"
*
.ends
*
*
