* File: sky130_fd_sc_lp__busdrivernovlp2_20.spice
* Created: Fri Aug 28 10:13:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__busdrivernovlp2_20.pex.spice"
.subckt sky130_fd_sc_lp__busdrivernovlp2_20  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1041 N_VGND_M1041_d N_TE_B_M1041_g N_A_27_367#_M1041_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1057 A_303_85# N_A_27_367#_M1057_g N_VGND_M1041_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1055 N_A_381_85#_M1055_d N_A_217_367#_M1055_g A_303_85# VNB NSHORT L=0.15
+ W=0.42 AD=0.1912 AS=0.0504 PD=1.8 PS=0.66 NRD=34.284 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1024 N_A_726_47#_M1024_d N_TE_B_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.4662 PD=1.12 PS=2.79 NRD=0 NRS=38.568 M=1 R=5.6
+ SA=75000.5 SB=75002.7 A=0.126 P=1.98 MULT=1
MM1049 N_A_726_47#_M1024_d N_TE_B_M1049_g N_VGND_M1049_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2646 PD=1.12 PS=1.47 NRD=0 NRS=49.992 M=1 R=5.6
+ SA=75000.9 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_726_47#_M1001_d N_A_M1001_g N_VGND_M1049_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2211 AS=0.2646 PD=1.47 PS=1.47 NRD=15 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_A_726_47#_M1001_d N_A_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2211 AS=0.277067 PD=1.47 PS=1.98667 NRD=15 NRS=15 M=1 R=5.6 SA=75002.3
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1018 N_A_1238_47#_M1018_d N_TE_B_M1018_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0735 AS=0.138533 PD=0.77 PS=0.993333 NRD=0 NRS=55.704 M=1 R=2.8
+ SA=75003 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_726_47#_M1011_g N_A_1238_47#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.0735 PD=1.43 PS=0.77 NRD=2.856 NRS=19.992 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_1451_47#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1002_d N_A_M1003_g N_A_1451_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.6
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1020 N_A_217_367#_M1020_d N_A_1238_47#_M1020_g N_A_1451_47#_M1003_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75001.1 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1039 N_A_217_367#_M1020_d N_A_1238_47#_M1039_g N_A_1451_47#_M1039_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1512 AS=0.2604 PD=1.2 PS=2.3 NRD=0 NRS=3.564 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A_726_47#_M1005_g N_Z_M1005_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75005.8 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1005_d N_A_726_47#_M1006_g N_Z_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75005.4 A=0.096 P=1.58 MULT=1
MM1013 N_VGND_M1013_d N_A_726_47#_M1013_g N_Z_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75004.9 A=0.096 P=1.58 MULT=1
MM1021 N_VGND_M1013_d N_A_726_47#_M1021_g N_Z_M1021_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75004.5 A=0.096 P=1.58 MULT=1
MM1029 N_VGND_M1029_d N_A_726_47#_M1029_g N_Z_M1021_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75004.1 A=0.096 P=1.58 MULT=1
MM1034 N_VGND_M1029_d N_A_726_47#_M1034_g N_Z_M1034_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.4
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1040 N_VGND_M1040_d N_A_726_47#_M1040_g N_Z_M1034_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.8
+ SB=75003.2 A=0.096 P=1.58 MULT=1
MM1043 N_VGND_M1040_d N_A_726_47#_M1043_g N_Z_M1043_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.2
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1046 N_VGND_M1046_d N_A_726_47#_M1046_g N_Z_M1043_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.7
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1047 N_VGND_M1046_d N_A_726_47#_M1047_g N_Z_M1047_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.1
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1054 N_VGND_M1054_d N_A_726_47#_M1054_g N_Z_M1047_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.5
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1056 N_VGND_M1054_d N_A_726_47#_M1056_g N_Z_M1056_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.9
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1058 N_VGND_M1058_d N_A_726_47#_M1058_g N_Z_M1056_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.4
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1059 N_VGND_M1058_d N_A_726_47#_M1059_g N_Z_M1059_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1052 N_VPWR_M1052_d N_TE_B_M1052_g N_A_27_367#_M1052_s VPB PSHORT L=0.15
+ W=0.84 AD=0.17304 AS=0.2268 PD=1.312 PS=2.22 NRD=23.443 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1015 N_A_217_367#_M1015_d N_A_27_367#_M1015_g N_VPWR_M1052_d VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.25956 PD=1.54 PS=1.968 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1019 N_A_217_367#_M1015_d N_A_27_367#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.24444 PD=1.54 PS=1.944 NRD=0 NRS=0 M=1 R=8.4 SA=75001
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1035 N_A_381_85#_M1035_d N_A_27_367#_M1035_g N_VPWR_M1019_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.16296 PD=1.12 PS=1.296 NRD=0 NRS=18.7544 M=1 R=5.6
+ SA=75001.4 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1038 N_VPWR_M1038_d N_A_217_367#_M1038_g N_A_381_85#_M1035_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2268 AS=0.1176 PD=2.22 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_658_367#_M1007_d N_A_381_85#_M1007_g N_A_726_47#_M1007_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.3906 AS=0.1764 PD=3.14 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1023 N_A_658_367#_M1023_d N_A_381_85#_M1023_g N_A_726_47#_M1007_s VPB PSHORT
+ L=0.15 W=1.26 AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.7 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_658_367#_M1023_d VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75001.2
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1045 N_VPWR_M1030_d N_A_M1045_g N_A_658_367#_M1045_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.5607 PD=1.54 PS=3.41 NRD=0 NRS=24.9993 M=1 R=8.4 SA=75001.6
+ SB=75000.4 A=0.189 P=2.82 MULT=1
MM1044 A_1260_373# N_TE_B_M1044_g N_VPWR_M1044_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2394 PD=1.08 PS=2.25 NRD=15.2281 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1000 N_A_1238_47#_M1000_d N_A_726_47#_M1000_g A_1260_373# VPB PSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1008 PD=2.25 PS=1.08 NRD=0 NRS=15.2281 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1028 N_A_217_367#_M1028_d N_A_M1028_g N_VPWR_M1028_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75009.8 A=0.189 P=2.82 MULT=1
MM1031 N_A_217_367#_M1028_d N_A_M1031_g N_VPWR_M1031_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.54495 PD=1.54 PS=2.125 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75000.6
+ SB=75009.4 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1031_s N_A_217_367#_M1004_g N_Z_M1004_s VPB PSHORT L=0.15 W=1.26
+ AD=0.54495 AS=0.1764 PD=2.125 PS=1.54 NRD=25.7873 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75008.4 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_217_367#_M1008_g N_Z_M1004_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75007.9 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1008_d N_A_217_367#_M1009_g N_Z_M1009_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75007.5 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A_217_367#_M1012_g N_Z_M1009_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75007.1 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1012_d N_A_217_367#_M1014_g N_Z_M1014_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75006.7 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A_217_367#_M1016_g N_Z_M1014_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1016_d N_A_217_367#_M1017_g N_Z_M1017_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75005.8 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_217_367#_M1022_g N_Z_M1017_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.7
+ SB=75005.4 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1022_d N_A_217_367#_M1025_g N_Z_M1025_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_A_217_367#_M1026_g N_Z_M1025_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.5
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1027 N_VPWR_M1026_d N_A_217_367#_M1027_g N_Z_M1027_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006 SB=75004.1
+ A=0.189 P=2.82 MULT=1
MM1032 N_VPWR_M1032_d N_A_217_367#_M1032_g N_Z_M1027_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.4
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1033 N_VPWR_M1032_d N_A_217_367#_M1033_g N_Z_M1033_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.8
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1036 N_VPWR_M1036_d N_A_217_367#_M1036_g N_Z_M1033_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.2
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1036_d N_A_217_367#_M1037_g N_Z_M1037_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.7
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1042 N_VPWR_M1042_d N_A_217_367#_M1042_g N_Z_M1037_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.1
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1048 N_VPWR_M1042_d N_A_217_367#_M1048_g N_Z_M1048_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.5
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1050 N_VPWR_M1050_d N_A_217_367#_M1050_g N_Z_M1048_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75009 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1051 N_VPWR_M1050_d N_A_217_367#_M1051_g N_Z_M1051_s VPB PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75009.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1053 N_VPWR_M1053_d N_A_217_367#_M1053_g N_Z_M1051_s VPB PSHORT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75009.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX60_noxref VNB VPB NWDIODE A=33.8311 P=40.01
c_212 VNB 0 1.75344e-19 $X=0 $Y=0
c_374 VPB 0 1.99473e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__busdrivernovlp2_20.pxi.spice"
*
.ends
*
*
