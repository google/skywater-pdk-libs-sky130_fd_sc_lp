* File: sky130_fd_sc_lp__o211ai_2.pex.spice
* Created: Fri Aug 28 11:02:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211AI_2%C1 1 3 6 8 10 13 15 16 24
r44 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.44
+ $X2=0.925 $Y2=1.44
r45 20 23 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.28 $Y=1.44
+ $X2=0.495 $Y2=1.44
r46 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.44 $X2=0.28 $Y2=1.44
r47 16 21 7.82051 $w=3.51e-07 $l=2.25e-07 $layer=LI1_cond $X=0.265 $Y=1.665
+ $X2=0.265 $Y2=1.44
r48 15 21 5.03989 $w=3.51e-07 $l=1.45e-07 $layer=LI1_cond $X=0.265 $Y=1.295
+ $X2=0.265 $Y2=1.44
r49 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.605
+ $X2=0.925 $Y2=1.44
r50 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.925 $Y=1.605
+ $X2=0.925 $Y2=2.465
r51 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.275
+ $X2=0.925 $Y2=1.44
r52 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.925 $Y=1.275
+ $X2=0.925 $Y2=0.745
r53 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.605
+ $X2=0.495 $Y2=1.44
r54 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.495 $Y=1.605
+ $X2=0.495 $Y2=2.465
r55 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.275
+ $X2=0.495 $Y2=1.44
r56 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.495 $Y=1.275
+ $X2=0.495 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%B1 1 3 6 8 10 13 15 16 23 24
c52 1 0 4.64396e-20 $X=1.355 $Y=1.275
r53 22 24 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.74 $Y=1.44
+ $X2=1.785 $Y2=1.44
r54 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.74
+ $Y=1.44 $X2=1.74 $Y2=1.44
r55 19 22 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=1.355 $Y=1.44
+ $X2=1.74 $Y2=1.44
r56 16 23 2.19513 $w=3.13e-07 $l=6e-08 $layer=LI1_cond $X=1.68 $Y=1.367 $X2=1.74
+ $Y2=1.367
r57 15 16 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.367 $X2=1.68
+ $Y2=1.367
r58 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.605
+ $X2=1.785 $Y2=1.44
r59 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.785 $Y=1.605
+ $X2=1.785 $Y2=2.465
r60 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.275
+ $X2=1.785 $Y2=1.44
r61 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.785 $Y=1.275
+ $X2=1.785 $Y2=0.745
r62 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.605
+ $X2=1.355 $Y2=1.44
r63 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.355 $Y=1.605
+ $X2=1.355 $Y2=2.465
r64 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.275
+ $X2=1.355 $Y2=1.44
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.355 $Y=1.275
+ $X2=1.355 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%A2 1 3 6 8 10 13 17 20 21 29 30 36
r59 25 27 15.383 $w=4.23e-07 $l=1.35e-07 $layer=POLY_cond $X=2.64 $Y=1.44
+ $X2=2.775 $Y2=1.44
r60 21 36 6.5849 $w=3.93e-07 $l=9.5e-08 $layer=LI1_cond $X=2.64 $Y=1.392
+ $X2=2.735 $Y2=1.392
r61 21 30 2.97593 $w=3.93e-07 $l=1.02e-07 $layer=LI1_cond $X=2.64 $Y=1.392
+ $X2=2.538 $Y2=1.392
r62 21 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=1.375 $X2=2.64 $Y2=1.375
r63 20 30 11.0284 $w=3.93e-07 $l=3.78e-07 $layer=LI1_cond $X=2.16 $Y=1.392
+ $X2=2.538 $Y2=1.392
r64 18 29 10.2553 $w=4.23e-07 $l=9e-08 $layer=POLY_cond $X=3.115 $Y=1.44
+ $X2=3.205 $Y2=1.44
r65 18 27 38.7423 $w=4.23e-07 $l=3.4e-07 $layer=POLY_cond $X=3.115 $Y=1.44
+ $X2=2.775 $Y2=1.44
r66 17 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.115 $Y=1.505
+ $X2=2.735 $Y2=1.505
r67 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.115
+ $Y=1.505 $X2=3.115 $Y2=1.505
r68 11 29 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.205 $Y=1.67
+ $X2=3.205 $Y2=1.44
r69 11 13 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=3.205 $Y=1.67
+ $X2=3.205 $Y2=2.465
r70 8 29 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.205 $Y=1.21
+ $X2=3.205 $Y2=1.44
r71 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.205 $Y=1.21
+ $X2=3.205 $Y2=0.68
r72 4 27 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.775 $Y=1.67
+ $X2=2.775 $Y2=1.44
r73 4 6 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.775 $Y=1.67
+ $X2=2.775 $Y2=2.465
r74 1 27 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.775 $Y=1.21
+ $X2=2.775 $Y2=1.44
r75 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.775 $Y=1.21
+ $X2=2.775 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%A1 1 3 6 8 10 13 20 24 25 29
c43 6 0 7.99068e-20 $X=3.635 $Y=2.465
r44 23 29 15.383 $w=4.23e-07 $l=1.35e-07 $layer=POLY_cond $X=4.2 $Y=1.44
+ $X2=4.065 $Y2=1.44
r45 22 24 6.145 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=1.4 $X2=4.115
+ $Y2=1.4
r46 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.2
+ $Y=1.375 $X2=4.2 $Y2=1.375
r47 20 25 7.7335 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=4.305 $Y=1.4
+ $X2=4.56 $Y2=1.4
r48 20 22 3.18438 $w=3.78e-07 $l=1.05e-07 $layer=LI1_cond $X=4.305 $Y=1.4
+ $X2=4.2 $Y2=1.4
r49 18 29 38.7423 $w=4.23e-07 $l=3.4e-07 $layer=POLY_cond $X=3.725 $Y=1.44
+ $X2=4.065 $Y2=1.44
r50 18 27 10.2553 $w=4.23e-07 $l=9e-08 $layer=POLY_cond $X=3.725 $Y=1.44
+ $X2=3.635 $Y2=1.44
r51 17 24 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.725 $Y=1.505
+ $X2=4.115 $Y2=1.505
r52 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.725
+ $Y=1.505 $X2=3.725 $Y2=1.505
r53 11 29 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.065 $Y=1.67
+ $X2=4.065 $Y2=1.44
r54 11 13 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=4.065 $Y=1.67
+ $X2=4.065 $Y2=2.465
r55 8 29 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.065 $Y=1.21
+ $X2=4.065 $Y2=1.44
r56 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.065 $Y=1.21
+ $X2=4.065 $Y2=0.68
r57 4 27 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.635 $Y=1.67
+ $X2=3.635 $Y2=1.44
r58 4 6 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=3.635 $Y=1.67
+ $X2=3.635 $Y2=2.465
r59 1 27 27.2344 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.635 $Y=1.21
+ $X2=3.635 $Y2=1.44
r60 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.635 $Y=1.21
+ $X2=3.635 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%VPWR 1 2 3 4 13 15 21 27 33 38 39 40 42 47
+ 57 58 64 67
r70 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r72 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r74 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r76 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.165 $Y=3.33 $X2=2
+ $Y2=3.33
r77 52 54 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r78 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r79 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r80 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r81 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.14 $Y2=3.33
r82 48 50 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 47 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=3.33 $X2=2
+ $Y2=3.33
r84 47 50 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r86 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r88 43 61 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r89 43 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r90 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.14 $Y2=3.33
r91 42 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r92 40 55 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r93 40 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 38 54 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.6 $Y2=3.33
r95 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.85 $Y2=3.33
r96 37 57 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=3.85 $Y2=3.33
r98 33 36 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.85 $Y=2.185
+ $X2=3.85 $Y2=2.95
r99 31 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=3.245
+ $X2=3.85 $Y2=3.33
r100 31 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.85 $Y=3.245
+ $X2=3.85 $Y2=2.95
r101 27 30 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2 $Y=2.185 $X2=2
+ $Y2=2.95
r102 25 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=3.33
r103 25 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=2.95
r104 21 24 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.14 $Y=2.185
+ $X2=1.14 $Y2=2.95
r105 19 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r106 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.95
r107 15 18 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.28 $Y=2.005
+ $X2=0.28 $Y2=2.95
r108 13 61 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r109 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.95
r110 4 36 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.835 $X2=3.85 $Y2=2.95
r111 4 33 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.835 $X2=3.85 $Y2=2.185
r112 3 30 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.95
r113 3 27 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.185
r114 2 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.95
r115 2 21 400 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.185
r116 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=2.95
r117 1 15 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%Y 1 2 3 4 13 17 21 25 31 32 33 34 35 36 37
+ 38 48 52
c56 34 0 4.64396e-20 $X=0.72 $Y=1.295
c57 21 0 7.99068e-20 $X=2.825 $Y=1.845
r58 46 52 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.71 $Y=0.98
+ $X2=0.71 $Y2=0.925
r59 38 66 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=0.71 $Y=2.775
+ $X2=0.71 $Y2=2.91
r60 37 38 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.405
+ $X2=0.71 $Y2=2.775
r61 36 37 22.7656 $w=1.88e-07 $l=3.9e-07 $layer=LI1_cond $X=0.71 $Y=2.015
+ $X2=0.71 $Y2=2.405
r62 34 35 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.665
r63 34 69 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.145
r64 33 69 5.78896 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.71 $Y=0.995
+ $X2=0.71 $Y2=1.145
r65 33 46 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.71 $Y=0.995
+ $X2=0.71 $Y2=0.98
r66 33 52 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.71 $Y=0.91
+ $X2=0.71 $Y2=0.925
r67 33 48 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.71 $Y=0.91
+ $X2=0.71 $Y2=0.68
r68 30 36 4.96172 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.93
+ $X2=0.71 $Y2=2.015
r69 30 31 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.71 $Y=1.93
+ $X2=0.745 $Y2=1.845
r70 29 35 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=0.745 $Y=1.76
+ $X2=0.745 $Y2=1.665
r71 29 31 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=1.76
+ $X2=0.745 $Y2=1.845
r72 25 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.99 $Y=1.97
+ $X2=2.99 $Y2=2.65
r73 23 25 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.99 $Y=1.93 $X2=2.99
+ $Y2=1.97
r74 22 32 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.665 $Y=1.845
+ $X2=1.57 $Y2=1.845
r75 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.825 $Y=1.845
+ $X2=2.99 $Y2=1.93
r76 21 22 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.825 $Y=1.845
+ $X2=1.665 $Y2=1.845
r77 17 19 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.57 $Y=1.98
+ $X2=1.57 $Y2=2.91
r78 15 32 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=1.93
+ $X2=1.57 $Y2=1.845
r79 15 17 2.91866 $w=1.88e-07 $l=5e-08 $layer=LI1_cond $X=1.57 $Y=1.93 $X2=1.57
+ $Y2=1.98
r80 14 31 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.875 $Y=1.845
+ $X2=0.745 $Y2=1.845
r81 13 32 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.475 $Y=1.845
+ $X2=1.57 $Y2=1.845
r82 13 14 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.475 $Y=1.845
+ $X2=0.875 $Y2=1.845
r83 4 27 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.835 $X2=2.99 $Y2=2.65
r84 4 25 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.835 $X2=2.99 $Y2=1.97
r85 3 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.91
r86 3 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=1.98
r87 2 66 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.91
r88 2 36 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=0.57 $Y=1.835
+ $X2=0.71 $Y2=2.015
r89 1 48 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.325 $X2=0.71 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%A_487_367# 1 2 3 12 14 15 17 20 21 24
r36 24 26 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=4.315 $Y=1.98
+ $X2=4.315 $Y2=2.91
r37 22 24 2.21624 $w=2.58e-07 $l=5e-08 $layer=LI1_cond $X=4.315 $Y=1.93
+ $X2=4.315 $Y2=1.98
r38 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.185 $Y=1.845
+ $X2=4.315 $Y2=1.93
r39 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.185 $Y=1.845
+ $X2=3.515 $Y2=1.845
r40 17 29 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.905
+ $X2=3.42 $Y2=2.99
r41 17 19 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=3.42 $Y=2.905
+ $X2=3.42 $Y2=1.98
r42 16 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.42 $Y=1.93
+ $X2=3.515 $Y2=1.845
r43 16 19 2.91866 $w=1.88e-07 $l=5e-08 $layer=LI1_cond $X=3.42 $Y=1.93 $X2=3.42
+ $Y2=1.98
r44 14 29 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.325 $Y=2.99
+ $X2=3.42 $Y2=2.99
r45 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.325 $Y=2.99
+ $X2=2.655 $Y2=2.99
r46 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.525 $Y=2.905
+ $X2=2.655 $Y2=2.99
r47 10 12 28.3678 $w=2.58e-07 $l=6.4e-07 $layer=LI1_cond $X=2.525 $Y=2.905
+ $X2=2.525 $Y2=2.265
r48 3 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.14
+ $Y=1.835 $X2=4.28 $Y2=2.91
r49 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.14
+ $Y=1.835 $X2=4.28 $Y2=1.98
r50 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.42 $Y2=2.91
r51 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.42 $Y2=1.98
r52 1 12 300 $w=1.7e-07 $l=4.88518e-07 $layer=licon1_PDIFF $count=2 $X=2.435
+ $Y=1.835 $X2=2.56 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%A_31_65# 1 2 3 12 14 15 18 22 25
r28 20 25 3.70046 $w=2.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.235 $Y=0.45
+ $X2=1.14 $Y2=0.45
r29 20 22 22.6056 $w=3.88e-07 $l=7.65e-07 $layer=LI1_cond $X=1.235 $Y=0.45 $X2=2
+ $Y2=0.45
r30 16 25 2.76953 $w=1.9e-07 $l=1.95e-07 $layer=LI1_cond $X=1.14 $Y=0.645
+ $X2=1.14 $Y2=0.45
r31 16 18 13.4258 $w=1.88e-07 $l=2.3e-07 $layer=LI1_cond $X=1.14 $Y=0.645
+ $X2=1.14 $Y2=0.875
r32 14 25 3.70046 $w=2.8e-07 $l=1.50167e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.14 $Y2=0.45
r33 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.375 $Y2=0.34
r34 10 15 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.375 $Y2=0.34
r35 10 12 1.85214 $w=2.78e-07 $l=4.5e-08 $layer=LI1_cond $X=0.235 $Y=0.425
+ $X2=0.235 $Y2=0.47
r36 3 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.325 $X2=2 $Y2=0.48
r37 2 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.325 $X2=1.14 $Y2=0.47
r38 2 18 182 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.325 $X2=1.14 $Y2=0.875
r39 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.325 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%A_286_65# 1 2 3 10 16 18 22 26
r47 26 27 13.9239 $w=1.84e-07 $l=2.1e-07 $layer=LI1_cond $X=2.99 $Y=0.955
+ $X2=2.99 $Y2=1.165
r48 20 22 38.5263 $w=1.88e-07 $l=6.6e-07 $layer=LI1_cond $X=3.85 $Y=1.08
+ $X2=3.85 $Y2=0.42
r49 19 27 1.1945 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.085 $Y=1.165
+ $X2=2.99 $Y2=1.165
r50 18 20 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.755 $Y=1.165
+ $X2=3.85 $Y2=1.08
r51 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.755 $Y=1.165
+ $X2=3.085 $Y2=1.165
r52 14 16 23.0574 $w=1.88e-07 $l=3.95e-07 $layer=LI1_cond $X=2.99 $Y=0.815
+ $X2=2.99 $Y2=0.42
r53 10 26 2.32065 $w=1.84e-07 $l=3.5e-08 $layer=LI1_cond $X=2.99 $Y=0.92
+ $X2=2.99 $Y2=0.955
r54 10 14 6.74211 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.92
+ $X2=2.99 $Y2=0.815
r55 10 12 69.9784 $w=2.08e-07 $l=1.325e-06 $layer=LI1_cond $X=2.895 $Y=0.92
+ $X2=1.57 $Y2=0.92
r56 3 22 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.26 $X2=3.85 $Y2=0.42
r57 2 26 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.26 $X2=2.99 $Y2=0.955
r58 2 16 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.26 $X2=2.99 $Y2=0.42
r59 1 12 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.325 $X2=1.57 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_2%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r60 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r61 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r62 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r63 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r64 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r65 41 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r66 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r67 38 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.56
+ $Y2=0
r68 38 40 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=3.12
+ $Y2=0
r69 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r70 33 37 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r71 32 36 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r72 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.56
+ $Y2=0
r74 30 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.16
+ $Y2=0
r75 28 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r76 28 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r77 26 43 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.08
+ $Y2=0
r78 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.28
+ $Y2=0
r79 25 46 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.56
+ $Y2=0
r80 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.28
+ $Y2=0
r81 23 40 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.12
+ $Y2=0
r82 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r83 22 43 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=4.08
+ $Y2=0
r84 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r85 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0
r86 18 20 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0.405
r87 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r88 14 16 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.405
r89 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r90 10 12 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.52
r91 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.26 $X2=4.28 $Y2=0.405
r92 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.28
+ $Y=0.26 $X2=3.42 $Y2=0.405
r93 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.26 $X2=2.56 $Y2=0.52
.ends

