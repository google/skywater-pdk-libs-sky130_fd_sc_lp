# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a311oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a311oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.210000 5.695000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 1.210000 3.810000 1.435000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 1.840000 1.435000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.865000 1.210000 7.700000 1.435000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.910000 1.210000 9.995000 1.435000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.335200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.995000 0.655000 4.355000 0.870000 ;
        RECT 3.995000 0.870000 9.655000 1.040000 ;
        RECT 3.995000 1.040000 4.175000 1.605000 ;
        RECT 3.995000 1.605000 9.265000 1.775000 ;
        RECT 4.950000 0.655000 5.210000 0.870000 ;
        RECT 5.805000 0.255000 6.045000 0.870000 ;
        RECT 6.715000 0.255000 6.950000 0.870000 ;
        RECT 7.620000 0.255000 7.865000 0.870000 ;
        RECT 8.175000 1.775000 8.365000 2.735000 ;
        RECT 8.535000 0.255000 8.725000 0.870000 ;
        RECT 9.035000 1.775000 9.265000 2.735000 ;
        RECT 9.395000 0.255000 9.655000 0.870000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.095000  0.255000  0.355000 0.870000 ;
      RECT 0.095000  0.870000  3.825000 1.040000 ;
      RECT 0.165000  1.815000  0.495000 3.245000 ;
      RECT 0.525000  0.085000  0.855000 0.700000 ;
      RECT 0.665000  1.605000  3.505000 1.775000 ;
      RECT 0.665000  1.775000  0.855000 3.075000 ;
      RECT 1.025000  0.255000  1.215000 0.870000 ;
      RECT 1.025000  1.945000  1.355000 3.245000 ;
      RECT 1.385000  0.085000  1.715000 0.700000 ;
      RECT 1.525000  1.775000  1.715000 3.075000 ;
      RECT 1.885000  0.255000  2.115000 0.870000 ;
      RECT 1.885000  1.945000  2.215000 3.245000 ;
      RECT 2.285000  0.255000  5.635000 0.445000 ;
      RECT 2.285000  0.445000  2.540000 0.700000 ;
      RECT 2.385000  1.775000  2.575000 3.075000 ;
      RECT 2.710000  0.665000  2.965000 0.870000 ;
      RECT 2.745000  1.945000  3.075000 3.245000 ;
      RECT 3.135000  0.445000  5.635000 0.485000 ;
      RECT 3.135000  0.485000  3.400000 0.700000 ;
      RECT 3.245000  1.775000  3.505000 1.945000 ;
      RECT 3.245000  1.945000  7.505000 2.115000 ;
      RECT 3.245000  2.115000  3.490000 3.075000 ;
      RECT 3.570000  0.665000  3.825000 0.870000 ;
      RECT 3.660000  2.285000  3.990000 3.245000 ;
      RECT 4.160000  2.115000  4.405000 3.075000 ;
      RECT 4.525000  0.485000  4.780000 0.700000 ;
      RECT 4.575000  2.285000  4.905000 3.245000 ;
      RECT 5.075000  2.115000  5.265000 3.075000 ;
      RECT 5.380000  0.485000  5.635000 0.700000 ;
      RECT 5.435000  2.285000  5.765000 3.245000 ;
      RECT 5.955000  2.285000  6.285000 2.905000 ;
      RECT 5.955000  2.905000  9.725000 3.075000 ;
      RECT 6.215000  0.085000  6.545000 0.700000 ;
      RECT 6.455000  2.115000  6.645000 2.735000 ;
      RECT 6.815000  2.285000  7.145000 2.905000 ;
      RECT 7.120000  0.085000  7.450000 0.700000 ;
      RECT 7.315000  2.115000  7.505000 2.735000 ;
      RECT 7.675000  1.945000  8.005000 2.905000 ;
      RECT 8.035000  0.085000  8.365000 0.700000 ;
      RECT 8.535000  1.945000  8.865000 2.905000 ;
      RECT 8.895000  0.085000  9.225000 0.700000 ;
      RECT 9.435000  1.815000  9.725000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__a311oi_4
END LIBRARY
