# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xnor2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__xnor2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.430000 0.715000 2.095000 ;
        RECT 0.085000 2.095000 0.570000 2.245000 ;
        RECT 0.545000 0.255000 1.340000 0.515000 ;
        RECT 0.545000 0.515000 0.715000 1.430000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.305000 1.425000 2.455000 1.895000 ;
        RECT 1.305000 1.895000 1.570000 2.095000 ;
        RECT 1.595000 1.220000 2.455000 1.425000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.303300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.270000 2.405000 3.270000 2.575000 ;
        RECT 2.270000 2.575000 2.600000 3.025000 ;
        RECT 2.750000 0.345000 3.270000 1.380000 ;
        RECT 3.100000 1.380000 3.270000 2.405000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.095000  0.085000 0.375000 1.260000 ;
      RECT 0.260000  2.415000 0.570000 3.245000 ;
      RECT 0.740000  2.265000 2.100000 2.435000 ;
      RECT 0.740000  2.435000 0.990000 3.065000 ;
      RECT 0.885000  0.930000 1.215000 1.260000 ;
      RECT 0.885000  1.260000 1.125000 2.265000 ;
      RECT 1.160000  2.605000 1.790000 3.245000 ;
      RECT 1.510000  0.345000 1.755000 0.845000 ;
      RECT 1.510000  0.845000 2.580000 1.035000 ;
      RECT 1.925000  0.085000 2.180000 0.675000 ;
      RECT 1.930000  2.065000 2.930000 2.235000 ;
      RECT 1.930000  2.235000 2.100000 2.265000 ;
      RECT 2.350000  0.345000 2.580000 0.845000 ;
      RECT 2.670000  1.565000 2.930000 2.065000 ;
      RECT 2.770000  2.745000 3.060000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__xnor2_0
END LIBRARY
