* File: sky130_fd_sc_lp__bufkapwr_4.spice
* Created: Fri Aug 28 10:11:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__bufkapwr_4.pex.spice"
.subckt sky130_fd_sc_lp__bufkapwr_4  VNB VPB A KAPWR X VGND VPWR
* 
* VGND	VGND
* X	X
* KAPWR	KAPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.1113 PD=0.755 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.07035 PD=0.7 PS=0.755 NRD=0 NRS=15.708 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1001_d N_A_27_47#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_27_47#_M1005_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1007 N_X_M1005_d N_A_27_47#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1218 PD=0.7 PS=1.42 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_KAPWR_M1009_d N_A_M1009_g N_A_27_47#_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2079 AS=0.3339 PD=1.59 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1000 N_KAPWR_M1009_d N_A_27_47#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2079 AS=0.1764 PD=1.59 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1003 N_KAPWR_M1003_d N_A_27_47#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_KAPWR_M1003_d N_A_27_47#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1008 N_KAPWR_M1008_d N_A_27_47#_M1008_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.378 AS=0.1764 PD=3.12 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__bufkapwr_4.pxi.spice"
*
.ends
*
*
