* File: sky130_fd_sc_lp__or2_lp.pxi.spice
* Created: Wed Sep  2 10:29:27 2020
* 
x_PM_SKY130_FD_SC_LP__OR2_LP%A N_A_M1004_g N_A_M1006_g N_A_M1001_g N_A_c_58_n
+ N_A_c_62_n A A A N_A_c_60_n PM_SKY130_FD_SC_LP__OR2_LP%A
x_PM_SKY130_FD_SC_LP__OR2_LP%B N_B_M1000_g N_B_c_91_n N_B_c_92_n N_B_c_93_n
+ N_B_M1002_g N_B_c_94_n N_B_M1008_g N_B_c_95_n B B B B N_B_c_97_n
+ PM_SKY130_FD_SC_LP__OR2_LP%B
x_PM_SKY130_FD_SC_LP__OR2_LP%A_196_114# N_A_196_114#_M1001_d
+ N_A_196_114#_M1000_d N_A_196_114#_M1009_g N_A_196_114#_M1005_g
+ N_A_196_114#_M1007_g N_A_196_114#_M1003_g N_A_196_114#_c_144_n
+ N_A_196_114#_c_151_n N_A_196_114#_c_152_n N_A_196_114#_c_145_n
+ N_A_196_114#_c_146_n N_A_196_114#_c_153_n N_A_196_114#_c_147_n
+ PM_SKY130_FD_SC_LP__OR2_LP%A_196_114#
x_PM_SKY130_FD_SC_LP__OR2_LP%VPWR N_VPWR_M1006_s N_VPWR_M1009_s N_VPWR_c_222_n
+ N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n
+ VPWR N_VPWR_c_228_n N_VPWR_c_221_n PM_SKY130_FD_SC_LP__OR2_LP%VPWR
x_PM_SKY130_FD_SC_LP__OR2_LP%X N_X_M1003_d N_X_M1007_d N_X_c_253_n X X X X X X
+ N_X_c_256_n PM_SKY130_FD_SC_LP__OR2_LP%X
x_PM_SKY130_FD_SC_LP__OR2_LP%VGND N_VGND_M1004_s N_VGND_M1008_d N_VGND_c_278_n
+ N_VGND_c_279_n N_VGND_c_280_n VGND N_VGND_c_281_n N_VGND_c_282_n
+ N_VGND_c_283_n N_VGND_c_284_n PM_SKY130_FD_SC_LP__OR2_LP%VGND
cc_1 VNB N_A_M1004_g 0.0267007f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.78
cc_2 VNB N_A_M1001_g 0.0203608f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.78
cc_3 VNB N_A_c_58_n 0.0278551f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.255
cc_4 VNB A 0.0306425f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_c_60_n 0.0283224f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.345
cc_6 VNB N_B_c_91_n 0.00951992f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.85
cc_7 VNB N_B_c_92_n 0.00619137f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.55
cc_8 VNB N_B_c_93_n 0.0154644f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.55
cc_9 VNB N_B_c_94_n 0.0152295f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.78
cc_10 VNB N_B_c_95_n 0.018598f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.255
cc_11 VNB B 0.0146309f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.85
cc_12 VNB N_B_c_97_n 0.0256817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_196_114#_M1005_g 0.0453872f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.255
cc_14 VNB N_A_196_114#_M1003_g 0.0485654f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_A_196_114#_c_144_n 0.00774921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_196_114#_c_145_n 0.00392246f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.345
cc_17 VNB N_A_196_114#_c_146_n 0.00612987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_196_114#_c_147_n 0.0175596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_221_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_253_n 0.0222321f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.78
cc_21 VNB X 0.033027f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.255
cc_22 VNB X 0.00653926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_256_n 0.00240475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_278_n 0.0128547f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.55
cc_25 VNB N_VGND_c_279_n 0.0466398f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.18
cc_26 VNB N_VGND_c_280_n 0.0286048f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.255
cc_27 VNB N_VGND_c_281_n 0.0437284f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.255
cc_28 VNB N_VGND_c_282_n 0.0343054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_283_n 0.245073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_284_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.345
cc_31 VPB N_A_M1006_g 0.0441527f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.55
cc_32 VPB N_A_c_62_n 0.0175467f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.85
cc_33 VPB A 0.0403144f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB N_A_c_60_n 0.00218109f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.345
cc_35 VPB N_B_M1000_g 0.0477921f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.78
cc_36 VPB N_B_c_91_n 0.0260194f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.85
cc_37 VPB N_B_c_92_n 0.00392357f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.55
cc_38 VPB B 0.00494183f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.85
cc_39 VPB N_A_196_114#_M1009_g 0.022993f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.18
cc_40 VPB N_A_196_114#_M1007_g 0.0248666f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.255
cc_41 VPB N_A_196_114#_c_144_n 0.0107071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_196_114#_c_151_n 0.00983191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_196_114#_c_152_n 0.0256611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_196_114#_c_153_n 0.00305473f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.345
cc_45 VPB N_A_196_114#_c_147_n 0.100729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_222_n 0.0462489f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.18
cc_47 VPB N_VPWR_c_223_n 0.0244777f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.255
cc_48 VPB N_VPWR_c_224_n 0.0121672f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.33
cc_49 VPB N_VPWR_c_225_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.255
cc_50 VPB N_VPWR_c_226_n 0.0323113f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.685
cc_51 VPB N_VPWR_c_227_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.85
cc_52 VPB N_VPWR_c_228_n 0.0390971f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_221_n 0.101943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB X 0.0386634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB X 0.0327986f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.33
cc_56 N_A_c_62_n N_B_M1000_g 0.0321625f $X=0.605 $Y=1.85 $X2=0 $Y2=0
cc_57 A N_B_c_92_n 0.00422067f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A_c_60_n N_B_c_92_n 0.0321625f $X=0.605 $Y=1.345 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_B_c_93_n 0.00909856f $X=0.905 $Y=0.78 $X2=0 $Y2=0
cc_60 N_A_c_58_n N_B_c_95_n 0.00909856f $X=0.905 $Y=1.255 $X2=0 $Y2=0
cc_61 N_A_c_60_n N_B_c_97_n 0.00191582f $X=0.605 $Y=1.345 $X2=0 $Y2=0
cc_62 N_A_M1001_g N_A_196_114#_c_144_n 0.00641868f $X=0.905 $Y=0.78 $X2=0 $Y2=0
cc_63 A N_A_196_114#_c_144_n 0.0516922f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A_c_60_n N_A_196_114#_c_144_n 0.00170713f $X=0.605 $Y=1.345 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_A_196_114#_c_151_n 0.00164966f $X=0.695 $Y=2.55 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_A_196_114#_c_146_n 0.00130204f $X=0.515 $Y=0.78 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_A_196_114#_c_146_n 0.00988314f $X=0.905 $Y=0.78 $X2=0 $Y2=0
cc_68 N_A_M1006_g N_A_196_114#_c_153_n 6.21071e-19 $X=0.695 $Y=2.55 $X2=0 $Y2=0
cc_69 A N_A_196_114#_c_153_n 0.0036782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_M1006_g N_VPWR_c_222_n 0.0139578f $X=0.695 $Y=2.55 $X2=0 $Y2=0
cc_71 N_A_c_62_n N_VPWR_c_222_n 7.3727e-19 $X=0.605 $Y=1.85 $X2=0 $Y2=0
cc_72 A N_VPWR_c_222_n 0.0305155f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_M1006_g N_VPWR_c_226_n 0.00370277f $X=0.695 $Y=2.55 $X2=0 $Y2=0
cc_74 N_A_M1006_g N_VPWR_c_221_n 0.00407315f $X=0.695 $Y=2.55 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_VGND_c_279_n 0.0141166f $X=0.515 $Y=0.78 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_VGND_c_279_n 0.0018473f $X=0.905 $Y=0.78 $X2=0 $Y2=0
cc_77 A N_VGND_c_279_n 0.0305157f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_VGND_c_281_n 0.00370277f $X=0.515 $Y=0.78 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_VGND_c_281_n 0.00428184f $X=0.905 $Y=0.78 $X2=0 $Y2=0
cc_80 N_A_M1004_g N_VGND_c_283_n 0.00407315f $X=0.515 $Y=0.78 $X2=0 $Y2=0
cc_81 N_A_M1001_g N_VGND_c_283_n 0.00484898f $X=0.905 $Y=0.78 $X2=0 $Y2=0
cc_82 N_B_c_94_n N_A_196_114#_M1005_g 0.00889596f $X=1.695 $Y=1.1 $X2=0 $Y2=0
cc_83 N_B_c_95_n N_A_196_114#_M1005_g 0.00976407f $X=1.695 $Y=1.175 $X2=0 $Y2=0
cc_84 B N_A_196_114#_M1005_g 0.0107061f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_85 N_B_M1000_g N_A_196_114#_c_144_n 0.00977495f $X=1.085 $Y=2.55 $X2=0 $Y2=0
cc_86 N_B_c_91_n N_A_196_114#_c_144_n 0.00949559f $X=1.455 $Y=1.695 $X2=0 $Y2=0
cc_87 N_B_c_92_n N_A_196_114#_c_144_n 0.00319796f $X=1.16 $Y=1.695 $X2=0 $Y2=0
cc_88 N_B_c_93_n N_A_196_114#_c_144_n 0.00152618f $X=1.335 $Y=1.1 $X2=0 $Y2=0
cc_89 N_B_c_95_n N_A_196_114#_c_144_n 0.00384023f $X=1.695 $Y=1.175 $X2=0 $Y2=0
cc_90 N_B_c_97_n N_A_196_114#_c_144_n 0.00201753f $X=1.62 $Y=1.265 $X2=0 $Y2=0
cc_91 N_B_M1000_g N_A_196_114#_c_151_n 0.0124882f $X=1.085 $Y=2.55 $X2=0 $Y2=0
cc_92 N_B_c_91_n N_A_196_114#_c_152_n 0.00192301f $X=1.455 $Y=1.695 $X2=0 $Y2=0
cc_93 B N_A_196_114#_c_152_n 0.0182598f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_94 B N_A_196_114#_c_145_n 0.0120291f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_95 N_B_c_97_n N_A_196_114#_c_145_n 2.23408e-19 $X=1.62 $Y=1.265 $X2=0 $Y2=0
cc_96 N_B_c_92_n N_A_196_114#_c_146_n 0.00306257f $X=1.16 $Y=1.695 $X2=0 $Y2=0
cc_97 N_B_c_93_n N_A_196_114#_c_146_n 0.00576325f $X=1.335 $Y=1.1 $X2=0 $Y2=0
cc_98 N_B_c_94_n N_A_196_114#_c_146_n 4.22319e-19 $X=1.695 $Y=1.1 $X2=0 $Y2=0
cc_99 B N_A_196_114#_c_146_n 0.0756613f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_100 N_B_M1000_g N_A_196_114#_c_153_n 0.00721486f $X=1.085 $Y=2.55 $X2=0 $Y2=0
cc_101 N_B_c_91_n N_A_196_114#_c_153_n 0.00601177f $X=1.455 $Y=1.695 $X2=0 $Y2=0
cc_102 B N_A_196_114#_c_153_n 5.54311e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_103 B N_A_196_114#_c_147_n 0.00146615f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_104 N_B_c_97_n N_A_196_114#_c_147_n 0.0101832f $X=1.62 $Y=1.265 $X2=0 $Y2=0
cc_105 N_B_M1000_g N_VPWR_c_222_n 0.0018343f $X=1.085 $Y=2.55 $X2=0 $Y2=0
cc_106 N_B_M1000_g N_VPWR_c_223_n 0.00343201f $X=1.085 $Y=2.55 $X2=0 $Y2=0
cc_107 N_B_M1000_g N_VPWR_c_226_n 0.00413742f $X=1.085 $Y=2.55 $X2=0 $Y2=0
cc_108 N_B_M1000_g N_VPWR_c_221_n 0.00484898f $X=1.085 $Y=2.55 $X2=0 $Y2=0
cc_109 N_B_c_94_n N_VGND_c_280_n 0.0022178f $X=1.695 $Y=1.1 $X2=0 $Y2=0
cc_110 B N_VGND_c_280_n 0.0292763f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_111 N_B_c_93_n N_VGND_c_281_n 0.00428184f $X=1.335 $Y=1.1 $X2=0 $Y2=0
cc_112 N_B_c_94_n N_VGND_c_281_n 7.53855e-19 $X=1.695 $Y=1.1 $X2=0 $Y2=0
cc_113 B N_VGND_c_281_n 0.0106551f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_114 N_B_c_93_n N_VGND_c_283_n 0.00484898f $X=1.335 $Y=1.1 $X2=0 $Y2=0
cc_115 B N_VGND_c_283_n 0.0116385f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_116 N_A_196_114#_c_151_n N_VPWR_c_222_n 0.0151773f $X=1.3 $Y=2.55 $X2=0 $Y2=0
cc_117 N_A_196_114#_M1009_g N_VPWR_c_223_n 0.0137423f $X=2.1 $Y=2.66 $X2=0 $Y2=0
cc_118 N_A_196_114#_M1007_g N_VPWR_c_223_n 0.00180376f $X=2.46 $Y=2.66 $X2=0
+ $Y2=0
cc_119 N_A_196_114#_c_151_n N_VPWR_c_223_n 0.0220739f $X=1.3 $Y=2.55 $X2=0 $Y2=0
cc_120 N_A_196_114#_c_152_n N_VPWR_c_223_n 0.0276676f $X=2.025 $Y=2.175 $X2=0
+ $Y2=0
cc_121 N_A_196_114#_c_151_n N_VPWR_c_226_n 0.00840064f $X=1.3 $Y=2.55 $X2=0
+ $Y2=0
cc_122 N_A_196_114#_M1009_g N_VPWR_c_228_n 0.00426961f $X=2.1 $Y=2.66 $X2=0
+ $Y2=0
cc_123 N_A_196_114#_M1007_g N_VPWR_c_228_n 0.00491683f $X=2.46 $Y=2.66 $X2=0
+ $Y2=0
cc_124 N_A_196_114#_M1009_g N_VPWR_c_221_n 0.00434697f $X=2.1 $Y=2.66 $X2=0
+ $Y2=0
cc_125 N_A_196_114#_M1007_g N_VPWR_c_221_n 0.00517496f $X=2.46 $Y=2.66 $X2=0
+ $Y2=0
cc_126 N_A_196_114#_c_151_n N_VPWR_c_221_n 0.0111899f $X=1.3 $Y=2.55 $X2=0 $Y2=0
cc_127 N_A_196_114#_M1005_g N_X_c_253_n 0.00213669f $X=2.345 $Y=0.78 $X2=0 $Y2=0
cc_128 N_A_196_114#_M1003_g N_X_c_253_n 0.00939721f $X=2.735 $Y=0.78 $X2=0 $Y2=0
cc_129 N_A_196_114#_M1005_g X 0.0119205f $X=2.345 $Y=0.78 $X2=0 $Y2=0
cc_130 N_A_196_114#_M1003_g X 0.0213771f $X=2.735 $Y=0.78 $X2=0 $Y2=0
cc_131 N_A_196_114#_M1009_g X 8.09475e-19 $X=2.1 $Y=2.66 $X2=0 $Y2=0
cc_132 N_A_196_114#_M1007_g X 0.00696891f $X=2.46 $Y=2.66 $X2=0 $Y2=0
cc_133 N_A_196_114#_M1003_g X 0.00222268f $X=2.735 $Y=0.78 $X2=0 $Y2=0
cc_134 N_A_196_114#_c_152_n X 0.0143663f $X=2.025 $Y=2.175 $X2=0 $Y2=0
cc_135 N_A_196_114#_c_145_n X 0.0398153f $X=2.19 $Y=1.755 $X2=0 $Y2=0
cc_136 N_A_196_114#_c_147_n X 0.049652f $X=2.735 $Y=1.925 $X2=0 $Y2=0
cc_137 N_A_196_114#_M1009_g X 0.00124449f $X=2.1 $Y=2.66 $X2=0 $Y2=0
cc_138 N_A_196_114#_M1007_g X 0.00996625f $X=2.46 $Y=2.66 $X2=0 $Y2=0
cc_139 N_A_196_114#_M1003_g N_X_c_256_n 0.00661078f $X=2.735 $Y=0.78 $X2=0 $Y2=0
cc_140 N_A_196_114#_c_146_n N_VGND_c_279_n 0.0145731f $X=1.12 $Y=0.78 $X2=0
+ $Y2=0
cc_141 N_A_196_114#_M1005_g N_VGND_c_280_n 0.0134474f $X=2.345 $Y=0.78 $X2=0
+ $Y2=0
cc_142 N_A_196_114#_M1003_g N_VGND_c_280_n 0.0018473f $X=2.735 $Y=0.78 $X2=0
+ $Y2=0
cc_143 N_A_196_114#_c_145_n N_VGND_c_280_n 0.00929697f $X=2.19 $Y=1.755 $X2=0
+ $Y2=0
cc_144 N_A_196_114#_c_147_n N_VGND_c_280_n 0.00154893f $X=2.735 $Y=1.925 $X2=0
+ $Y2=0
cc_145 N_A_196_114#_c_146_n N_VGND_c_281_n 0.00779082f $X=1.12 $Y=0.78 $X2=0
+ $Y2=0
cc_146 N_A_196_114#_M1005_g N_VGND_c_282_n 0.00370277f $X=2.345 $Y=0.78 $X2=0
+ $Y2=0
cc_147 N_A_196_114#_M1003_g N_VGND_c_282_n 0.00428184f $X=2.735 $Y=0.78 $X2=0
+ $Y2=0
cc_148 N_A_196_114#_M1005_g N_VGND_c_283_n 0.00407315f $X=2.345 $Y=0.78 $X2=0
+ $Y2=0
cc_149 N_A_196_114#_M1003_g N_VGND_c_283_n 0.00484898f $X=2.735 $Y=0.78 $X2=0
+ $Y2=0
cc_150 N_A_196_114#_c_146_n N_VGND_c_283_n 0.0104511f $X=1.12 $Y=0.78 $X2=0
+ $Y2=0
cc_151 N_VPWR_c_223_n X 0.0162933f $X=1.885 $Y=2.66 $X2=0 $Y2=0
cc_152 N_VPWR_c_228_n X 0.0235675f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_153 N_VPWR_c_221_n X 0.0251781f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_154 N_X_c_253_n N_VGND_c_280_n 0.0145731f $X=2.95 $Y=0.78 $X2=0 $Y2=0
cc_155 N_X_c_253_n N_VGND_c_282_n 0.00784587f $X=2.95 $Y=0.78 $X2=0 $Y2=0
cc_156 N_X_c_253_n N_VGND_c_283_n 0.0104774f $X=2.95 $Y=0.78 $X2=0 $Y2=0
