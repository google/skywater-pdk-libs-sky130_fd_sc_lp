* File: sky130_fd_sc_lp__bufbuf_8.pxi.spice
* Created: Wed Sep  2 09:35:35 2020
* 
x_PM_SKY130_FD_SC_LP__BUFBUF_8%A_117_265# N_A_117_265#_M1004_d
+ N_A_117_265#_M1018_d N_A_117_265#_M1000_d N_A_117_265#_M1025_d
+ N_A_117_265#_M1002_g N_A_117_265#_M1001_g N_A_117_265#_M1009_g
+ N_A_117_265#_M1003_g N_A_117_265#_M1012_g N_A_117_265#_M1006_g
+ N_A_117_265#_M1013_g N_A_117_265#_M1008_g N_A_117_265#_M1017_g
+ N_A_117_265#_M1015_g N_A_117_265#_M1020_g N_A_117_265#_M1016_g
+ N_A_117_265#_M1022_g N_A_117_265#_M1021_g N_A_117_265#_M1024_g
+ N_A_117_265#_M1023_g N_A_117_265#_c_137_n N_A_117_265#_c_138_n
+ N_A_117_265#_c_139_n N_A_117_265#_c_140_n N_A_117_265#_c_141_n
+ N_A_117_265#_c_258_p N_A_117_265#_c_156_n N_A_117_265#_c_194_p
+ N_A_117_265#_c_213_p N_A_117_265#_c_313_p N_A_117_265#_c_142_n
+ N_A_117_265#_c_157_n N_A_117_265#_c_158_n N_A_117_265#_c_143_n
+ N_A_117_265#_c_144_n N_A_117_265#_c_159_n N_A_117_265#_c_145_n
+ PM_SKY130_FD_SC_LP__BUFBUF_8%A_117_265#
x_PM_SKY130_FD_SC_LP__BUFBUF_8%A_837_23# N_A_837_23#_M1007_s N_A_837_23#_M1019_s
+ N_A_837_23#_M1004_g N_A_837_23#_M1000_g N_A_837_23#_M1010_g
+ N_A_837_23#_M1014_g N_A_837_23#_M1018_g N_A_837_23#_M1025_g
+ N_A_837_23#_c_329_n N_A_837_23#_c_330_n N_A_837_23#_c_331_n
+ N_A_837_23#_c_339_n N_A_837_23#_c_340_n N_A_837_23#_c_332_n
+ N_A_837_23#_c_333_n N_A_837_23#_c_334_n PM_SKY130_FD_SC_LP__BUFBUF_8%A_837_23#
x_PM_SKY130_FD_SC_LP__BUFBUF_8%A_1217_23# N_A_1217_23#_M1005_d
+ N_A_1217_23#_M1011_d N_A_1217_23#_M1007_g N_A_1217_23#_M1019_g
+ N_A_1217_23#_c_429_n N_A_1217_23#_c_415_n N_A_1217_23#_c_416_n
+ N_A_1217_23#_c_417_n N_A_1217_23#_c_436_n N_A_1217_23#_c_455_p
+ N_A_1217_23#_c_422_n N_A_1217_23#_c_418_n N_A_1217_23#_c_448_p
+ N_A_1217_23#_c_419_n PM_SKY130_FD_SC_LP__BUFBUF_8%A_1217_23#
x_PM_SKY130_FD_SC_LP__BUFBUF_8%A N_A_M1005_g N_A_M1011_g A N_A_c_474_n
+ N_A_c_475_n PM_SKY130_FD_SC_LP__BUFBUF_8%A
x_PM_SKY130_FD_SC_LP__BUFBUF_8%VPWR N_VPWR_M1001_s N_VPWR_M1003_s N_VPWR_M1008_s
+ N_VPWR_M1016_s N_VPWR_M1023_s N_VPWR_M1014_s N_VPWR_M1019_d N_VPWR_c_502_n
+ N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n
+ N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n
+ N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_515_n VPWR N_VPWR_c_516_n
+ N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_501_n N_VPWR_c_521_n
+ N_VPWR_c_522_n N_VPWR_c_523_n N_VPWR_c_524_n PM_SKY130_FD_SC_LP__BUFBUF_8%VPWR
x_PM_SKY130_FD_SC_LP__BUFBUF_8%X N_X_M1002_s N_X_M1012_s N_X_M1017_s N_X_M1022_s
+ N_X_M1001_d N_X_M1006_d N_X_M1015_d N_X_M1021_d N_X_c_607_n N_X_c_616_n
+ N_X_c_617_n N_X_c_682_n N_X_c_706_p N_X_c_608_n N_X_c_618_n N_X_c_686_n
+ N_X_c_703_p N_X_c_609_n N_X_c_619_n N_X_c_690_n N_X_c_707_p N_X_c_610_n
+ N_X_c_620_n N_X_c_694_n N_X_c_708_p N_X_c_621_n N_X_c_611_n N_X_c_622_n
+ N_X_c_612_n N_X_c_623_n N_X_c_613_n X X N_X_c_614_n X
+ PM_SKY130_FD_SC_LP__BUFBUF_8%X
x_PM_SKY130_FD_SC_LP__BUFBUF_8%VGND N_VGND_M1002_d N_VGND_M1009_d N_VGND_M1013_d
+ N_VGND_M1020_d N_VGND_M1024_d N_VGND_M1010_s N_VGND_M1007_d N_VGND_c_717_n
+ N_VGND_c_718_n N_VGND_c_719_n N_VGND_c_720_n N_VGND_c_721_n N_VGND_c_722_n
+ N_VGND_c_723_n N_VGND_c_724_n N_VGND_c_725_n N_VGND_c_726_n N_VGND_c_727_n
+ N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n VGND N_VGND_c_731_n
+ N_VGND_c_732_n N_VGND_c_733_n N_VGND_c_734_n N_VGND_c_735_n N_VGND_c_736_n
+ N_VGND_c_737_n N_VGND_c_738_n N_VGND_c_739_n PM_SKY130_FD_SC_LP__BUFBUF_8%VGND
cc_1 VNB N_A_117_265#_M1002_g 0.0261659f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.665
cc_2 VNB N_A_117_265#_M1009_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.665
cc_3 VNB N_A_117_265#_M1012_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=0.665
cc_4 VNB N_A_117_265#_M1013_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=0.665
cc_5 VNB N_A_117_265#_M1017_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.665
cc_6 VNB N_A_117_265#_M1020_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.665
cc_7 VNB N_A_117_265#_M1022_g 0.0213881f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=0.665
cc_8 VNB N_A_117_265#_M1024_g 0.0222095f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.665
cc_9 VNB N_A_117_265#_c_137_n 0.00180021f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=1.49
cc_10 VNB N_A_117_265#_c_138_n 0.153471f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.49
cc_11 VNB N_A_117_265#_c_139_n 0.00162357f $X=-0.19 $Y=-0.245 $X2=3.92 $Y2=1.395
cc_12 VNB N_A_117_265#_c_140_n 6.66824e-19 $X=-0.19 $Y=-0.245 $X2=3.92 $Y2=1.755
cc_13 VNB N_A_117_265#_c_141_n 0.00256213f $X=-0.19 $Y=-0.245 $X2=4.36 $Y2=1.14
cc_14 VNB N_A_117_265#_c_142_n 0.00660339f $X=-0.19 $Y=-0.245 $X2=5.24 $Y2=1.14
cc_15 VNB N_A_117_265#_c_143_n 0.00888512f $X=-0.19 $Y=-0.245 $X2=5.335
+ $Y2=0.455
cc_16 VNB N_A_117_265#_c_144_n 0.00117784f $X=-0.19 $Y=-0.245 $X2=3.92 $Y2=1.49
cc_17 VNB N_A_117_265#_c_145_n 0.00163095f $X=-0.19 $Y=-0.245 $X2=4.465 $Y2=1.14
cc_18 VNB N_A_837_23#_M1004_g 0.0221777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_837_23#_M1010_g 0.0213937f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.655
cc_20 VNB N_A_837_23#_M1018_g 0.0273834f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.655
cc_21 VNB N_A_837_23#_c_329_n 0.00119513f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=0.665
cc_22 VNB N_A_837_23#_c_330_n 0.0510334f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=0.665
cc_23 VNB N_A_837_23#_c_331_n 0.0118771f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.655
cc_24 VNB N_A_837_23#_c_332_n 0.00116062f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.465
cc_25 VNB N_A_837_23#_c_333_n 4.38724e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_837_23#_c_334_n 0.0443276f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.325
cc_27 VNB N_A_1217_23#_M1019_g 0.00651157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_1217_23#_c_415_n 0.0367739f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.465
cc_29 VNB N_A_1217_23#_c_416_n 8.46216e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_1217_23#_c_417_n 0.0170073f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.325
cc_31 VNB N_A_1217_23#_c_418_n 0.0188262f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.325
cc_32 VNB N_A_1217_23#_c_419_n 0.0210931f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.655
cc_33 VNB N_A_M1005_g 0.0320091f $X=-0.19 $Y=-0.245 $X2=4.335 $Y2=1.835
cc_34 VNB N_A_c_474_n 0.0332723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_c_475_n 0.0112128f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.325
cc_36 VNB N_VPWR_c_501_n 0.302998f $X=-0.19 $Y=-0.245 $X2=5.21 $Y2=1.84
cc_37 VNB N_X_c_607_n 0.00426803f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.655
cc_38 VNB N_X_c_608_n 0.00304705f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=0.665
cc_39 VNB N_X_c_609_n 0.00304705f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.325
cc_40 VNB N_X_c_610_n 0.005522f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=2.465
cc_41 VNB N_X_c_611_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.49
cc_42 VNB N_X_c_612_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=3.92 $Y2=1.225
cc_43 VNB N_X_c_613_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=3.92 $Y2=1.585
cc_44 VNB N_X_c_614_n 0.0216863f $X=-0.19 $Y=-0.245 $X2=4.472 $Y2=1.925
cc_45 VNB X 0.0247579f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=2.05
cc_46 VNB N_VGND_c_717_n 0.028153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_718_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_719_n 0.0131884f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=0.665
cc_49 VNB N_VGND_c_720_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.465
cc_50 VNB N_VGND_c_721_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=0.665
cc_51 VNB N_VGND_c_722_n 4.77201e-19 $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=2.465
cc_52 VNB N_VGND_c_723_n 6.14598e-19 $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.665
cc_53 VNB N_VGND_c_724_n 0.0158701f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.465
cc_54 VNB N_VGND_c_725_n 0.014713f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.665
cc_55 VNB N_VGND_c_726_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_727_n 0.0131884f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.655
cc_57 VNB N_VGND_c_728_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=2.465
cc_58 VNB N_VGND_c_729_n 0.0302792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_730_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=1.325
cc_60 VNB N_VGND_c_731_n 0.0131884f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.665
cc_61 VNB N_VGND_c_732_n 0.0131884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_733_n 0.0136491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_734_n 0.0217702f $X=-0.19 $Y=-0.245 $X2=4.335 $Y2=1.84
cc_64 VNB N_VGND_c_735_n 0.382206f $X=-0.19 $Y=-0.245 $X2=4.005 $Y2=1.84
cc_65 VNB N_VGND_c_736_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=2.05
cc_66 VNB N_VGND_c_737_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_738_n 0.0048588f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=0.455
cc_68 VNB N_VGND_c_739_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=4.57 $Y2=1.14
cc_69 VPB N_A_117_265#_M1001_g 0.0235615f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=2.465
cc_70 VPB N_A_117_265#_M1003_g 0.0190623f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=2.465
cc_71 VPB N_A_117_265#_M1006_g 0.0190623f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=2.465
cc_72 VPB N_A_117_265#_M1008_g 0.0190623f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=2.465
cc_73 VPB N_A_117_265#_M1015_g 0.0190623f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=2.465
cc_74 VPB N_A_117_265#_M1016_g 0.0190623f $X=-0.19 $Y=1.655 $X2=2.925 $Y2=2.465
cc_75 VPB N_A_117_265#_M1021_g 0.0190376f $X=-0.19 $Y=1.655 $X2=3.355 $Y2=2.465
cc_76 VPB N_A_117_265#_M1023_g 0.0193192f $X=-0.19 $Y=1.655 $X2=3.785 $Y2=2.465
cc_77 VPB N_A_117_265#_c_138_n 0.0223314f $X=-0.19 $Y=1.655 $X2=3.81 $Y2=1.49
cc_78 VPB N_A_117_265#_c_140_n 9.56747e-19 $X=-0.19 $Y=1.655 $X2=3.92 $Y2=1.755
cc_79 VPB N_A_117_265#_c_156_n 0.00234165f $X=-0.19 $Y=1.655 $X2=4.335 $Y2=1.84
cc_80 VPB N_A_117_265#_c_157_n 0.00621042f $X=-0.19 $Y=1.655 $X2=5.21 $Y2=1.84
cc_81 VPB N_A_117_265#_c_158_n 0.0145824f $X=-0.19 $Y=1.655 $X2=5.335 $Y2=2.05
cc_82 VPB N_A_117_265#_c_159_n 0.00224133f $X=-0.19 $Y=1.655 $X2=4.472 $Y2=1.84
cc_83 VPB N_A_837_23#_M1000_g 0.0197585f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.325
cc_84 VPB N_A_837_23#_M1014_g 0.0190431f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.325
cc_85 VPB N_A_837_23#_M1025_g 0.0242637f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.325
cc_86 VPB N_A_837_23#_c_330_n 0.0254777f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=0.665
cc_87 VPB N_A_837_23#_c_339_n 0.00329534f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=1.325
cc_88 VPB N_A_837_23#_c_340_n 0.00964986f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=0.665
cc_89 VPB N_A_837_23#_c_333_n 0.0030419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_837_23#_c_334_n 0.00467327f $X=-0.19 $Y=1.655 $X2=2.925 $Y2=1.325
cc_91 VPB N_A_1217_23#_M1019_g 0.0248447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_1217_23#_c_416_n 0.0014624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_1217_23#_c_422_n 0.0133501f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.655
cc_94 VPB N_A_M1011_g 0.0285806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_c_474_n 0.00687124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_c_475_n 0.0070564f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.325
cc_97 VPB N_VPWR_c_502_n 0.0418465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_503_n 0.00400996f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=0.665
cc_99 VPB N_VPWR_c_504_n 0.0166024f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=2.465
cc_100 VPB N_VPWR_c_505_n 0.00400996f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=0.665
cc_101 VPB N_VPWR_c_506_n 0.00396563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_507_n 0.00215653f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=2.465
cc_103 VPB N_VPWR_c_508_n 0.00463375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_509_n 0.0230442f $X=-0.19 $Y=1.655 $X2=3.355 $Y2=0.665
cc_105 VPB N_VPWR_c_510_n 0.014713f $X=-0.19 $Y=1.655 $X2=3.355 $Y2=1.655
cc_106 VPB N_VPWR_c_511_n 0.00564836f $X=-0.19 $Y=1.655 $X2=3.355 $Y2=2.465
cc_107 VPB N_VPWR_c_512_n 0.0166024f $X=-0.19 $Y=1.655 $X2=3.355 $Y2=2.465
cc_108 VPB N_VPWR_c_513_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_514_n 0.0169258f $X=-0.19 $Y=1.655 $X2=3.785 $Y2=0.665
cc_110 VPB N_VPWR_c_515_n 0.00497514f $X=-0.19 $Y=1.655 $X2=3.785 $Y2=0.665
cc_111 VPB N_VPWR_c_516_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_517_n 0.0147711f $X=-0.19 $Y=1.655 $X2=3.92 $Y2=1.395
cc_113 VPB N_VPWR_c_518_n 0.0333204f $X=-0.19 $Y=1.655 $X2=4.475 $Y2=2.05
cc_114 VPB N_VPWR_c_519_n 0.0218729f $X=-0.19 $Y=1.655 $X2=4.57 $Y2=1.14
cc_115 VPB N_VPWR_c_501_n 0.089887f $X=-0.19 $Y=1.655 $X2=5.21 $Y2=1.84
cc_116 VPB N_VPWR_c_521_n 0.00497514f $X=-0.19 $Y=1.655 $X2=5.355 $Y2=2.05
cc_117 VPB N_VPWR_c_522_n 0.00497514f $X=-0.19 $Y=1.655 $X2=5.335 $Y2=2.84
cc_118 VPB N_VPWR_c_523_n 0.00510842f $X=-0.19 $Y=1.655 $X2=5.37 $Y2=0.455
cc_119 VPB N_VPWR_c_524_n 0.00510842f $X=-0.19 $Y=1.655 $X2=3.92 $Y2=1.49
cc_120 VPB N_X_c_616_n 0.00351027f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=2.465
cc_121 VPB N_X_c_617_n 0.0216377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_X_c_618_n 0.00240399f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=1.655
cc_123 VPB N_X_c_619_n 0.00240399f $X=-0.19 $Y=1.655 $X2=2.925 $Y2=0.665
cc_124 VPB N_X_c_620_n 0.0047539f $X=-0.19 $Y=1.655 $X2=3.785 $Y2=1.325
cc_125 VPB N_X_c_621_n 0.00210048f $X=-0.19 $Y=1.655 $X2=3.81 $Y2=1.49
cc_126 VPB N_X_c_622_n 0.00210048f $X=-0.19 $Y=1.655 $X2=3.81 $Y2=1.49
cc_127 VPB N_X_c_623_n 0.00210048f $X=-0.19 $Y=1.655 $X2=3.92 $Y2=1.395
cc_128 VPB X 0.00597596f $X=-0.19 $Y=1.655 $X2=4.475 $Y2=2.05
cc_129 N_A_117_265#_M1024_g N_A_837_23#_M1004_g 0.0180966f $X=3.785 $Y=0.665
+ $X2=0 $Y2=0
cc_130 N_A_117_265#_c_139_n N_A_837_23#_M1004_g 0.00350436f $X=3.92 $Y=1.395
+ $X2=0 $Y2=0
cc_131 N_A_117_265#_c_141_n N_A_837_23#_M1004_g 0.0148344f $X=4.36 $Y=1.14 $X2=0
+ $Y2=0
cc_132 N_A_117_265#_M1023_g N_A_837_23#_M1000_g 0.018608f $X=3.785 $Y=2.465
+ $X2=0 $Y2=0
cc_133 N_A_117_265#_c_156_n N_A_837_23#_M1000_g 0.0131985f $X=4.335 $Y=1.84
+ $X2=0 $Y2=0
cc_134 N_A_117_265#_c_159_n N_A_837_23#_M1000_g 0.0011944f $X=4.472 $Y=1.84
+ $X2=0 $Y2=0
cc_135 N_A_117_265#_c_142_n N_A_837_23#_M1010_g 0.014127f $X=5.24 $Y=1.14 $X2=0
+ $Y2=0
cc_136 N_A_117_265#_c_157_n N_A_837_23#_M1014_g 0.0141989f $X=5.21 $Y=1.84 $X2=0
+ $Y2=0
cc_137 N_A_117_265#_c_142_n N_A_837_23#_M1018_g 0.015399f $X=5.24 $Y=1.14 $X2=0
+ $Y2=0
cc_138 N_A_117_265#_c_157_n N_A_837_23#_M1025_g 0.0150166f $X=5.21 $Y=1.84 $X2=0
+ $Y2=0
cc_139 N_A_117_265#_c_138_n N_A_837_23#_c_329_n 2.17684e-19 $X=3.81 $Y=1.49
+ $X2=0 $Y2=0
cc_140 N_A_117_265#_c_141_n N_A_837_23#_c_329_n 0.0120203f $X=4.36 $Y=1.14 $X2=0
+ $Y2=0
cc_141 N_A_117_265#_c_156_n N_A_837_23#_c_329_n 0.0102209f $X=4.335 $Y=1.84
+ $X2=0 $Y2=0
cc_142 N_A_117_265#_c_142_n N_A_837_23#_c_329_n 0.0682115f $X=5.24 $Y=1.14 $X2=0
+ $Y2=0
cc_143 N_A_117_265#_c_157_n N_A_837_23#_c_329_n 0.0656013f $X=5.21 $Y=1.84 $X2=0
+ $Y2=0
cc_144 N_A_117_265#_c_144_n N_A_837_23#_c_329_n 0.0160482f $X=3.92 $Y=1.49 $X2=0
+ $Y2=0
cc_145 N_A_117_265#_c_159_n N_A_837_23#_c_329_n 0.0223524f $X=4.472 $Y=1.84
+ $X2=0 $Y2=0
cc_146 N_A_117_265#_c_145_n N_A_837_23#_c_329_n 0.0170684f $X=4.465 $Y=1.14
+ $X2=0 $Y2=0
cc_147 N_A_117_265#_c_142_n N_A_837_23#_c_330_n 0.00766569f $X=5.24 $Y=1.14
+ $X2=0 $Y2=0
cc_148 N_A_117_265#_c_157_n N_A_837_23#_c_330_n 0.00769592f $X=5.21 $Y=1.84
+ $X2=0 $Y2=0
cc_149 N_A_117_265#_c_142_n N_A_837_23#_c_331_n 0.0109849f $X=5.24 $Y=1.14 $X2=0
+ $Y2=0
cc_150 N_A_117_265#_c_143_n N_A_837_23#_c_331_n 0.0370206f $X=5.335 $Y=0.455
+ $X2=0 $Y2=0
cc_151 N_A_117_265#_c_158_n N_A_837_23#_c_339_n 0.0446617f $X=5.335 $Y=2.05
+ $X2=0 $Y2=0
cc_152 N_A_117_265#_c_157_n N_A_837_23#_c_333_n 0.00897907f $X=5.21 $Y=1.84
+ $X2=0 $Y2=0
cc_153 N_A_117_265#_c_138_n N_A_837_23#_c_334_n 0.0217948f $X=3.81 $Y=1.49 $X2=0
+ $Y2=0
cc_154 N_A_117_265#_c_140_n N_A_837_23#_c_334_n 0.00350436f $X=3.92 $Y=1.755
+ $X2=0 $Y2=0
cc_155 N_A_117_265#_c_142_n N_A_837_23#_c_334_n 0.00243542f $X=5.24 $Y=1.14
+ $X2=0 $Y2=0
cc_156 N_A_117_265#_c_157_n N_A_837_23#_c_334_n 0.00243542f $X=5.21 $Y=1.84
+ $X2=0 $Y2=0
cc_157 N_A_117_265#_c_144_n N_A_837_23#_c_334_n 7.20588e-19 $X=3.92 $Y=1.49
+ $X2=0 $Y2=0
cc_158 N_A_117_265#_c_159_n N_A_837_23#_c_334_n 0.00253619f $X=4.472 $Y=1.84
+ $X2=0 $Y2=0
cc_159 N_A_117_265#_c_145_n N_A_837_23#_c_334_n 0.00253619f $X=4.465 $Y=1.14
+ $X2=0 $Y2=0
cc_160 N_A_117_265#_c_158_n N_A_1217_23#_M1019_g 0.00725096f $X=5.335 $Y=2.05
+ $X2=0 $Y2=0
cc_161 N_A_117_265#_c_143_n N_A_1217_23#_c_419_n 0.00411175f $X=5.335 $Y=0.455
+ $X2=0 $Y2=0
cc_162 N_A_117_265#_c_156_n N_VPWR_M1023_s 0.00129688f $X=4.335 $Y=1.84 $X2=0
+ $Y2=0
cc_163 N_A_117_265#_c_194_p N_VPWR_M1023_s 9.73829e-19 $X=4.005 $Y=1.84 $X2=0
+ $Y2=0
cc_164 N_A_117_265#_c_157_n N_VPWR_M1014_s 0.00176461f $X=5.21 $Y=1.84 $X2=0
+ $Y2=0
cc_165 N_A_117_265#_M1001_g N_VPWR_c_502_n 0.00343774f $X=0.775 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_117_265#_M1003_g N_VPWR_c_503_n 0.0016342f $X=1.205 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_117_265#_M1006_g N_VPWR_c_503_n 0.0016342f $X=1.635 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_117_265#_M1006_g N_VPWR_c_504_n 0.00585385f $X=1.635 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_117_265#_M1008_g N_VPWR_c_504_n 0.00585385f $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_117_265#_M1008_g N_VPWR_c_505_n 0.0016342f $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_117_265#_M1015_g N_VPWR_c_505_n 0.0016342f $X=2.495 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_117_265#_M1016_g N_VPWR_c_506_n 0.0016342f $X=2.925 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_117_265#_M1021_g N_VPWR_c_506_n 0.00158567f $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_174 N_A_117_265#_M1021_g N_VPWR_c_507_n 7.77579e-19 $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_117_265#_M1023_g N_VPWR_c_507_n 0.0142387f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_117_265#_c_138_n N_VPWR_c_507_n 3.98642e-19 $X=3.81 $Y=1.49 $X2=0
+ $Y2=0
cc_177 N_A_117_265#_c_156_n N_VPWR_c_507_n 0.00997062f $X=4.335 $Y=1.84 $X2=0
+ $Y2=0
cc_178 N_A_117_265#_c_194_p N_VPWR_c_507_n 0.00992353f $X=4.005 $Y=1.84 $X2=0
+ $Y2=0
cc_179 N_A_117_265#_c_157_n N_VPWR_c_508_n 0.0135055f $X=5.21 $Y=1.84 $X2=0
+ $Y2=0
cc_180 N_A_117_265#_M1001_g N_VPWR_c_512_n 0.00585385f $X=0.775 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_117_265#_M1003_g N_VPWR_c_512_n 0.00585385f $X=1.205 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_117_265#_c_213_p N_VPWR_c_514_n 0.0154684f $X=4.475 $Y=2.05 $X2=0
+ $Y2=0
cc_183 N_A_117_265#_M1015_g N_VPWR_c_516_n 0.00585385f $X=2.495 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_117_265#_M1016_g N_VPWR_c_516_n 0.00585385f $X=2.925 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_117_265#_M1021_g N_VPWR_c_517_n 0.00585385f $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_117_265#_M1023_g N_VPWR_c_517_n 0.00486043f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_117_265#_c_158_n N_VPWR_c_518_n 0.0188755f $X=5.335 $Y=2.05 $X2=0
+ $Y2=0
cc_188 N_A_117_265#_M1000_d N_VPWR_c_501_n 0.00245236f $X=4.335 $Y=1.835 $X2=0
+ $Y2=0
cc_189 N_A_117_265#_M1025_d N_VPWR_c_501_n 0.00271622f $X=5.195 $Y=1.835 $X2=0
+ $Y2=0
cc_190 N_A_117_265#_M1001_g N_VPWR_c_501_n 0.0117494f $X=0.775 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_117_265#_M1003_g N_VPWR_c_501_n 0.0106302f $X=1.205 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_A_117_265#_M1006_g N_VPWR_c_501_n 0.0106302f $X=1.635 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A_117_265#_M1008_g N_VPWR_c_501_n 0.0106302f $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A_117_265#_M1015_g N_VPWR_c_501_n 0.0106302f $X=2.495 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_117_265#_M1016_g N_VPWR_c_501_n 0.0106302f $X=2.925 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A_117_265#_M1021_g N_VPWR_c_501_n 0.0106302f $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A_117_265#_M1023_g N_VPWR_c_501_n 0.00835506f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_117_265#_c_213_p N_VPWR_c_501_n 0.0106136f $X=4.475 $Y=2.05 $X2=0
+ $Y2=0
cc_199 N_A_117_265#_c_158_n N_VPWR_c_501_n 0.0111968f $X=5.335 $Y=2.05 $X2=0
+ $Y2=0
cc_200 N_A_117_265#_M1002_g N_X_c_607_n 0.0160451f $X=0.775 $Y=0.665 $X2=0 $Y2=0
cc_201 N_A_117_265#_c_137_n N_X_c_607_n 0.0217546f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_202 N_A_117_265#_c_138_n N_X_c_607_n 0.00280073f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_203 N_A_117_265#_M1001_g N_X_c_616_n 0.016117f $X=0.775 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A_117_265#_c_137_n N_X_c_616_n 0.0192302f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_205 N_A_117_265#_c_138_n N_X_c_616_n 0.00280073f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_206 N_A_117_265#_M1009_g N_X_c_608_n 0.014127f $X=1.205 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A_117_265#_M1012_g N_X_c_608_n 0.014127f $X=1.635 $Y=0.665 $X2=0 $Y2=0
cc_208 N_A_117_265#_c_137_n N_X_c_608_n 0.0471185f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_209 N_A_117_265#_c_138_n N_X_c_608_n 0.00243542f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_210 N_A_117_265#_M1003_g N_X_c_618_n 0.0141989f $X=1.205 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_117_265#_M1006_g N_X_c_618_n 0.0141989f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_117_265#_c_137_n N_X_c_618_n 0.0420697f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_213 N_A_117_265#_c_138_n N_X_c_618_n 0.00243542f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_214 N_A_117_265#_M1013_g N_X_c_609_n 0.014127f $X=2.065 $Y=0.665 $X2=0 $Y2=0
cc_215 N_A_117_265#_M1017_g N_X_c_609_n 0.014127f $X=2.495 $Y=0.665 $X2=0 $Y2=0
cc_216 N_A_117_265#_c_137_n N_X_c_609_n 0.0471185f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_217 N_A_117_265#_c_138_n N_X_c_609_n 0.00243542f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_218 N_A_117_265#_M1008_g N_X_c_619_n 0.0141989f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A_117_265#_M1015_g N_X_c_619_n 0.0141989f $X=2.495 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A_117_265#_c_137_n N_X_c_619_n 0.0420697f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_221 N_A_117_265#_c_138_n N_X_c_619_n 0.00243542f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_222 N_A_117_265#_M1020_g N_X_c_610_n 0.0140805f $X=2.925 $Y=0.665 $X2=0 $Y2=0
cc_223 N_A_117_265#_M1022_g N_X_c_610_n 0.0137149f $X=3.355 $Y=0.665 $X2=0 $Y2=0
cc_224 N_A_117_265#_M1024_g N_X_c_610_n 0.00121251f $X=3.785 $Y=0.665 $X2=0
+ $Y2=0
cc_225 N_A_117_265#_c_137_n N_X_c_610_n 0.0625611f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_226 N_A_117_265#_c_138_n N_X_c_610_n 0.00497162f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_227 N_A_117_265#_c_258_p N_X_c_610_n 0.0137028f $X=4.005 $Y=1.14 $X2=0 $Y2=0
cc_228 N_A_117_265#_M1016_g N_X_c_620_n 0.0141523f $X=2.925 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A_117_265#_M1021_g N_X_c_620_n 0.013934f $X=3.355 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_117_265#_M1023_g N_X_c_620_n 7.40393e-19 $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_231 N_A_117_265#_c_137_n N_X_c_620_n 0.0603575f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_232 N_A_117_265#_c_138_n N_X_c_620_n 0.00497162f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_233 N_A_117_265#_c_194_p N_X_c_620_n 0.0108938f $X=4.005 $Y=1.84 $X2=0 $Y2=0
cc_234 N_A_117_265#_c_137_n N_X_c_621_n 0.021133f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_235 N_A_117_265#_c_138_n N_X_c_621_n 0.00253619f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_236 N_A_117_265#_c_137_n N_X_c_611_n 0.0154426f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_237 N_A_117_265#_c_138_n N_X_c_611_n 0.00253619f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_238 N_A_117_265#_c_137_n N_X_c_622_n 0.021133f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_239 N_A_117_265#_c_138_n N_X_c_622_n 0.00253619f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_240 N_A_117_265#_c_137_n N_X_c_612_n 0.0154426f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_241 N_A_117_265#_c_138_n N_X_c_612_n 0.00253619f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_242 N_A_117_265#_c_137_n N_X_c_623_n 0.021133f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_243 N_A_117_265#_c_138_n N_X_c_623_n 0.00253619f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_244 N_A_117_265#_c_137_n N_X_c_613_n 0.0154426f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_245 N_A_117_265#_c_138_n N_X_c_613_n 0.00253619f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_246 N_A_117_265#_M1002_g X 0.00320084f $X=0.775 $Y=0.665 $X2=0 $Y2=0
cc_247 N_A_117_265#_M1001_g X 0.00320084f $X=0.775 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A_117_265#_c_137_n X 0.0150718f $X=3.835 $Y=1.49 $X2=0 $Y2=0
cc_249 N_A_117_265#_c_138_n X 0.00757048f $X=3.81 $Y=1.49 $X2=0 $Y2=0
cc_250 N_A_117_265#_c_141_n N_VGND_M1024_d 0.00129688f $X=4.36 $Y=1.14 $X2=0
+ $Y2=0
cc_251 N_A_117_265#_c_258_p N_VGND_M1024_d 9.73829e-19 $X=4.005 $Y=1.14 $X2=0
+ $Y2=0
cc_252 N_A_117_265#_c_142_n N_VGND_M1010_s 0.00176461f $X=5.24 $Y=1.14 $X2=0
+ $Y2=0
cc_253 N_A_117_265#_M1002_g N_VGND_c_717_n 0.0118775f $X=0.775 $Y=0.665 $X2=0
+ $Y2=0
cc_254 N_A_117_265#_M1009_g N_VGND_c_717_n 6.60038e-19 $X=1.205 $Y=0.665 $X2=0
+ $Y2=0
cc_255 N_A_117_265#_M1002_g N_VGND_c_718_n 6.60038e-19 $X=0.775 $Y=0.665 $X2=0
+ $Y2=0
cc_256 N_A_117_265#_M1009_g N_VGND_c_718_n 0.010814f $X=1.205 $Y=0.665 $X2=0
+ $Y2=0
cc_257 N_A_117_265#_M1012_g N_VGND_c_718_n 0.010814f $X=1.635 $Y=0.665 $X2=0
+ $Y2=0
cc_258 N_A_117_265#_M1013_g N_VGND_c_718_n 6.60038e-19 $X=2.065 $Y=0.665 $X2=0
+ $Y2=0
cc_259 N_A_117_265#_M1012_g N_VGND_c_719_n 0.00477554f $X=1.635 $Y=0.665 $X2=0
+ $Y2=0
cc_260 N_A_117_265#_M1013_g N_VGND_c_719_n 0.00477554f $X=2.065 $Y=0.665 $X2=0
+ $Y2=0
cc_261 N_A_117_265#_M1012_g N_VGND_c_720_n 6.60038e-19 $X=1.635 $Y=0.665 $X2=0
+ $Y2=0
cc_262 N_A_117_265#_M1013_g N_VGND_c_720_n 0.010814f $X=2.065 $Y=0.665 $X2=0
+ $Y2=0
cc_263 N_A_117_265#_M1017_g N_VGND_c_720_n 0.010814f $X=2.495 $Y=0.665 $X2=0
+ $Y2=0
cc_264 N_A_117_265#_M1020_g N_VGND_c_720_n 6.60038e-19 $X=2.925 $Y=0.665 $X2=0
+ $Y2=0
cc_265 N_A_117_265#_M1017_g N_VGND_c_721_n 6.60038e-19 $X=2.495 $Y=0.665 $X2=0
+ $Y2=0
cc_266 N_A_117_265#_M1020_g N_VGND_c_721_n 0.010814f $X=2.925 $Y=0.665 $X2=0
+ $Y2=0
cc_267 N_A_117_265#_M1022_g N_VGND_c_721_n 0.010814f $X=3.355 $Y=0.665 $X2=0
+ $Y2=0
cc_268 N_A_117_265#_M1024_g N_VGND_c_721_n 6.60038e-19 $X=3.785 $Y=0.665 $X2=0
+ $Y2=0
cc_269 N_A_117_265#_M1022_g N_VGND_c_722_n 6.61235e-19 $X=3.355 $Y=0.665 $X2=0
+ $Y2=0
cc_270 N_A_117_265#_M1024_g N_VGND_c_722_n 0.0109705f $X=3.785 $Y=0.665 $X2=0
+ $Y2=0
cc_271 N_A_117_265#_c_138_n N_VGND_c_722_n 3.98642e-19 $X=3.81 $Y=1.49 $X2=0
+ $Y2=0
cc_272 N_A_117_265#_c_141_n N_VGND_c_722_n 0.0102332f $X=4.36 $Y=1.14 $X2=0
+ $Y2=0
cc_273 N_A_117_265#_c_258_p N_VGND_c_722_n 0.00992353f $X=4.005 $Y=1.14 $X2=0
+ $Y2=0
cc_274 N_A_117_265#_c_142_n N_VGND_c_723_n 0.0170777f $X=5.24 $Y=1.14 $X2=0
+ $Y2=0
cc_275 N_A_117_265#_M1002_g N_VGND_c_727_n 0.00477554f $X=0.775 $Y=0.665 $X2=0
+ $Y2=0
cc_276 N_A_117_265#_M1009_g N_VGND_c_727_n 0.00477554f $X=1.205 $Y=0.665 $X2=0
+ $Y2=0
cc_277 N_A_117_265#_c_143_n N_VGND_c_729_n 0.0145405f $X=5.335 $Y=0.455 $X2=0
+ $Y2=0
cc_278 N_A_117_265#_M1017_g N_VGND_c_731_n 0.00477554f $X=2.495 $Y=0.665 $X2=0
+ $Y2=0
cc_279 N_A_117_265#_M1020_g N_VGND_c_731_n 0.00477554f $X=2.925 $Y=0.665 $X2=0
+ $Y2=0
cc_280 N_A_117_265#_M1022_g N_VGND_c_732_n 0.00477554f $X=3.355 $Y=0.665 $X2=0
+ $Y2=0
cc_281 N_A_117_265#_M1024_g N_VGND_c_732_n 0.00477554f $X=3.785 $Y=0.665 $X2=0
+ $Y2=0
cc_282 N_A_117_265#_c_313_p N_VGND_c_733_n 0.0107575f $X=4.475 $Y=0.455 $X2=0
+ $Y2=0
cc_283 N_A_117_265#_M1004_d N_VGND_c_735_n 0.00476883f $X=4.335 $Y=0.245 $X2=0
+ $Y2=0
cc_284 N_A_117_265#_M1018_d N_VGND_c_735_n 0.00374439f $X=5.195 $Y=0.245 $X2=0
+ $Y2=0
cc_285 N_A_117_265#_M1002_g N_VGND_c_735_n 0.0083043f $X=0.775 $Y=0.665 $X2=0
+ $Y2=0
cc_286 N_A_117_265#_M1009_g N_VGND_c_735_n 0.0083043f $X=1.205 $Y=0.665 $X2=0
+ $Y2=0
cc_287 N_A_117_265#_M1012_g N_VGND_c_735_n 0.0083043f $X=1.635 $Y=0.665 $X2=0
+ $Y2=0
cc_288 N_A_117_265#_M1013_g N_VGND_c_735_n 0.0083043f $X=2.065 $Y=0.665 $X2=0
+ $Y2=0
cc_289 N_A_117_265#_M1017_g N_VGND_c_735_n 0.0083043f $X=2.495 $Y=0.665 $X2=0
+ $Y2=0
cc_290 N_A_117_265#_M1020_g N_VGND_c_735_n 0.0083043f $X=2.925 $Y=0.665 $X2=0
+ $Y2=0
cc_291 N_A_117_265#_M1022_g N_VGND_c_735_n 0.0083043f $X=3.355 $Y=0.665 $X2=0
+ $Y2=0
cc_292 N_A_117_265#_M1024_g N_VGND_c_735_n 0.0083043f $X=3.785 $Y=0.665 $X2=0
+ $Y2=0
cc_293 N_A_117_265#_c_313_p N_VGND_c_735_n 0.00794711f $X=4.475 $Y=0.455 $X2=0
+ $Y2=0
cc_294 N_A_117_265#_c_143_n N_VGND_c_735_n 0.00985747f $X=5.335 $Y=0.455 $X2=0
+ $Y2=0
cc_295 N_A_837_23#_c_330_n N_A_1217_23#_M1019_g 0.00610168f $X=5.71 $Y=1.49
+ $X2=0 $Y2=0
cc_296 N_A_837_23#_c_339_n N_A_1217_23#_M1019_g 4.39703e-19 $X=5.955 $Y=1.93
+ $X2=0 $Y2=0
cc_297 N_A_837_23#_c_332_n N_A_1217_23#_M1019_g 4.67154e-19 $X=5.89 $Y=1.49
+ $X2=0 $Y2=0
cc_298 N_A_837_23#_c_333_n N_A_1217_23#_M1019_g 0.00387294f $X=5.955 $Y=1.815
+ $X2=0 $Y2=0
cc_299 N_A_837_23#_c_331_n N_A_1217_23#_c_429_n 0.0120985f $X=5.925 $Y=0.6 $X2=0
+ $Y2=0
cc_300 N_A_837_23#_c_332_n N_A_1217_23#_c_429_n 0.0107215f $X=5.89 $Y=1.49 $X2=0
+ $Y2=0
cc_301 N_A_837_23#_c_330_n N_A_1217_23#_c_415_n 0.0124746f $X=5.71 $Y=1.49 $X2=0
+ $Y2=0
cc_302 N_A_837_23#_c_332_n N_A_1217_23#_c_415_n 9.96272e-19 $X=5.89 $Y=1.49
+ $X2=0 $Y2=0
cc_303 N_A_837_23#_c_339_n N_A_1217_23#_c_416_n 0.004536f $X=5.955 $Y=1.93 $X2=0
+ $Y2=0
cc_304 N_A_837_23#_c_332_n N_A_1217_23#_c_416_n 0.00400662f $X=5.89 $Y=1.49
+ $X2=0 $Y2=0
cc_305 N_A_837_23#_c_333_n N_A_1217_23#_c_416_n 0.0137256f $X=5.955 $Y=1.815
+ $X2=0 $Y2=0
cc_306 N_A_837_23#_c_331_n N_A_1217_23#_c_436_n 0.0139413f $X=5.925 $Y=0.6 $X2=0
+ $Y2=0
cc_307 N_A_837_23#_c_331_n N_A_1217_23#_c_419_n 0.0114909f $X=5.925 $Y=0.6 $X2=0
+ $Y2=0
cc_308 N_A_837_23#_M1000_g N_VPWR_c_507_n 0.00171522f $X=4.26 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_837_23#_M1014_g N_VPWR_c_508_n 0.00163259f $X=4.69 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A_837_23#_M1025_g N_VPWR_c_508_n 0.00312749f $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_837_23#_M1000_g N_VPWR_c_514_n 0.00585385f $X=4.26 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A_837_23#_M1014_g N_VPWR_c_514_n 0.00585385f $X=4.69 $Y=2.465 $X2=0
+ $Y2=0
cc_313 N_A_837_23#_M1025_g N_VPWR_c_518_n 0.00585385f $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_A_837_23#_c_340_n N_VPWR_c_518_n 0.00599726f $X=5.985 $Y=1.98 $X2=0
+ $Y2=0
cc_315 N_A_837_23#_M1019_s N_VPWR_c_501_n 0.00448802f $X=5.86 $Y=1.835 $X2=0
+ $Y2=0
cc_316 N_A_837_23#_M1000_g N_VPWR_c_501_n 0.0107878f $X=4.26 $Y=2.465 $X2=0
+ $Y2=0
cc_317 N_A_837_23#_M1014_g N_VPWR_c_501_n 0.0106439f $X=4.69 $Y=2.465 $X2=0
+ $Y2=0
cc_318 N_A_837_23#_M1025_g N_VPWR_c_501_n 0.0120162f $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_319 N_A_837_23#_c_340_n N_VPWR_c_501_n 0.00759383f $X=5.985 $Y=1.98 $X2=0
+ $Y2=0
cc_320 N_A_837_23#_M1004_g N_VGND_c_722_n 0.00918433f $X=4.26 $Y=0.665 $X2=0
+ $Y2=0
cc_321 N_A_837_23#_M1010_g N_VGND_c_722_n 6.37194e-19 $X=4.69 $Y=0.665 $X2=0
+ $Y2=0
cc_322 N_A_837_23#_M1004_g N_VGND_c_723_n 6.68496e-19 $X=4.26 $Y=0.665 $X2=0
+ $Y2=0
cc_323 N_A_837_23#_M1010_g N_VGND_c_723_n 0.0108688f $X=4.69 $Y=0.665 $X2=0
+ $Y2=0
cc_324 N_A_837_23#_M1018_g N_VGND_c_723_n 0.013405f $X=5.12 $Y=0.665 $X2=0 $Y2=0
cc_325 N_A_837_23#_c_331_n N_VGND_c_724_n 0.0321795f $X=5.925 $Y=0.6 $X2=0 $Y2=0
cc_326 N_A_837_23#_M1018_g N_VGND_c_729_n 0.00477554f $X=5.12 $Y=0.665 $X2=0
+ $Y2=0
cc_327 N_A_837_23#_c_331_n N_VGND_c_729_n 0.00832758f $X=5.925 $Y=0.6 $X2=0
+ $Y2=0
cc_328 N_A_837_23#_M1004_g N_VGND_c_733_n 0.00554242f $X=4.26 $Y=0.665 $X2=0
+ $Y2=0
cc_329 N_A_837_23#_M1010_g N_VGND_c_733_n 0.00477554f $X=4.69 $Y=0.665 $X2=0
+ $Y2=0
cc_330 N_A_837_23#_M1007_s N_VGND_c_735_n 0.00481424f $X=5.8 $Y=0.245 $X2=0
+ $Y2=0
cc_331 N_A_837_23#_M1004_g N_VGND_c_735_n 0.00954162f $X=4.26 $Y=0.665 $X2=0
+ $Y2=0
cc_332 N_A_837_23#_M1010_g N_VGND_c_735_n 0.0083043f $X=4.69 $Y=0.665 $X2=0
+ $Y2=0
cc_333 N_A_837_23#_M1018_g N_VGND_c_735_n 0.00960399f $X=5.12 $Y=0.665 $X2=0
+ $Y2=0
cc_334 N_A_837_23#_c_331_n N_VGND_c_735_n 0.00902581f $X=5.925 $Y=0.6 $X2=0
+ $Y2=0
cc_335 N_A_1217_23#_c_429_n N_A_M1005_g 7.91722e-19 $X=6.275 $Y=1.36 $X2=0 $Y2=0
cc_336 N_A_1217_23#_c_415_n N_A_M1005_g 0.0211689f $X=6.275 $Y=1.36 $X2=0 $Y2=0
cc_337 N_A_1217_23#_c_417_n N_A_M1005_g 0.0152966f $X=6.775 $Y=1.15 $X2=0 $Y2=0
cc_338 N_A_1217_23#_c_418_n N_A_M1005_g 0.00688485f $X=6.94 $Y=0.875 $X2=0 $Y2=0
cc_339 N_A_1217_23#_c_419_n N_A_M1005_g 0.0103363f $X=6.262 $Y=1.195 $X2=0 $Y2=0
cc_340 N_A_1217_23#_c_422_n N_A_M1011_g 0.0162967f $X=6.94 $Y=2.06 $X2=0 $Y2=0
cc_341 N_A_1217_23#_M1019_g N_A_c_474_n 0.0262383f $X=6.2 $Y=2.465 $X2=0 $Y2=0
cc_342 N_A_1217_23#_c_416_n N_A_c_474_n 0.00521339f $X=6.34 $Y=1.925 $X2=0 $Y2=0
cc_343 N_A_1217_23#_c_417_n N_A_c_474_n 0.00463857f $X=6.775 $Y=1.15 $X2=0 $Y2=0
cc_344 N_A_1217_23#_c_422_n N_A_c_474_n 9.46187e-19 $X=6.94 $Y=2.06 $X2=0 $Y2=0
cc_345 N_A_1217_23#_c_448_p N_A_c_474_n 7.91722e-19 $X=6.315 $Y=1.525 $X2=0
+ $Y2=0
cc_346 N_A_1217_23#_M1019_g N_A_c_475_n 2.31571e-19 $X=6.2 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A_1217_23#_c_415_n N_A_c_475_n 4.23032e-19 $X=6.275 $Y=1.36 $X2=0 $Y2=0
cc_348 N_A_1217_23#_c_417_n N_A_c_475_n 0.0369939f $X=6.775 $Y=1.15 $X2=0 $Y2=0
cc_349 N_A_1217_23#_c_422_n N_A_c_475_n 0.0337563f $X=6.94 $Y=2.06 $X2=0 $Y2=0
cc_350 N_A_1217_23#_c_448_p N_A_c_475_n 0.0229154f $X=6.315 $Y=1.525 $X2=0 $Y2=0
cc_351 N_A_1217_23#_c_416_n N_VPWR_M1019_d 0.00108321f $X=6.34 $Y=1.925 $X2=0
+ $Y2=0
cc_352 N_A_1217_23#_c_455_p N_VPWR_M1019_d 0.00118409f $X=6.44 $Y=2.062 $X2=0
+ $Y2=0
cc_353 N_A_1217_23#_c_422_n N_VPWR_M1019_d 0.00842854f $X=6.94 $Y=2.06 $X2=0
+ $Y2=0
cc_354 N_A_1217_23#_M1019_g N_VPWR_c_509_n 0.0235546f $X=6.2 $Y=2.465 $X2=0
+ $Y2=0
cc_355 N_A_1217_23#_c_455_p N_VPWR_c_509_n 0.0116817f $X=6.44 $Y=2.062 $X2=0
+ $Y2=0
cc_356 N_A_1217_23#_c_422_n N_VPWR_c_509_n 0.0116482f $X=6.94 $Y=2.06 $X2=0
+ $Y2=0
cc_357 N_A_1217_23#_M1019_g N_VPWR_c_518_n 0.00486043f $X=6.2 $Y=2.465 $X2=0
+ $Y2=0
cc_358 N_A_1217_23#_M1019_g N_VPWR_c_501_n 0.00975473f $X=6.2 $Y=2.465 $X2=0
+ $Y2=0
cc_359 N_A_1217_23#_c_417_n N_VGND_M1007_d 0.00310216f $X=6.775 $Y=1.15 $X2=0
+ $Y2=0
cc_360 N_A_1217_23#_c_436_n N_VGND_M1007_d 0.0016378f $X=6.44 $Y=1.15 $X2=0
+ $Y2=0
cc_361 N_A_1217_23#_c_415_n N_VGND_c_724_n 0.00104341f $X=6.275 $Y=1.36 $X2=0
+ $Y2=0
cc_362 N_A_1217_23#_c_417_n N_VGND_c_724_n 0.00801802f $X=6.775 $Y=1.15 $X2=0
+ $Y2=0
cc_363 N_A_1217_23#_c_436_n N_VGND_c_724_n 0.0152745f $X=6.44 $Y=1.15 $X2=0
+ $Y2=0
cc_364 N_A_1217_23#_c_418_n N_VGND_c_724_n 0.0139248f $X=6.94 $Y=0.875 $X2=0
+ $Y2=0
cc_365 N_A_1217_23#_c_419_n N_VGND_c_724_n 0.0196188f $X=6.262 $Y=1.195 $X2=0
+ $Y2=0
cc_366 N_A_1217_23#_c_419_n N_VGND_c_729_n 0.00477554f $X=6.262 $Y=1.195 $X2=0
+ $Y2=0
cc_367 N_A_1217_23#_c_418_n N_VGND_c_734_n 0.00536063f $X=6.94 $Y=0.875 $X2=0
+ $Y2=0
cc_368 N_A_1217_23#_c_418_n N_VGND_c_735_n 0.00962526f $X=6.94 $Y=0.875 $X2=0
+ $Y2=0
cc_369 N_A_1217_23#_c_419_n N_VGND_c_735_n 0.00960399f $X=6.262 $Y=1.195 $X2=0
+ $Y2=0
cc_370 N_A_M1011_g N_VPWR_c_509_n 0.00652757f $X=6.725 $Y=2.155 $X2=0 $Y2=0
cc_371 N_A_M1011_g N_VPWR_c_519_n 0.00312414f $X=6.725 $Y=2.155 $X2=0 $Y2=0
cc_372 N_A_M1011_g N_VPWR_c_501_n 0.00410284f $X=6.725 $Y=2.155 $X2=0 $Y2=0
cc_373 N_A_M1005_g N_VGND_c_724_n 0.00559556f $X=6.725 $Y=0.875 $X2=0 $Y2=0
cc_374 N_A_M1005_g N_VGND_c_734_n 0.00380885f $X=6.725 $Y=0.875 $X2=0 $Y2=0
cc_375 N_A_M1005_g N_VGND_c_735_n 0.00458517f $X=6.725 $Y=0.875 $X2=0 $Y2=0
cc_376 N_VPWR_c_501_n N_X_M1001_d 0.003017f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPWR_c_501_n N_X_M1006_d 0.003017f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_378 N_VPWR_c_501_n N_X_M1015_d 0.003017f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_379 N_VPWR_c_501_n N_X_M1021_d 0.00423456f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_M1001_s N_X_c_616_n 0.00299978f $X=0.415 $Y=1.835 $X2=0 $Y2=0
cc_381 N_VPWR_c_502_n N_X_c_616_n 0.0185481f $X=0.56 $Y=2.27 $X2=0 $Y2=0
cc_382 N_VPWR_c_502_n N_X_c_617_n 7.64598e-19 $X=0.56 $Y=2.27 $X2=0 $Y2=0
cc_383 N_VPWR_c_512_n N_X_c_682_n 0.0149362f $X=1.29 $Y=3.33 $X2=0 $Y2=0
cc_384 N_VPWR_c_501_n N_X_c_682_n 0.0100304f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_M1003_s N_X_c_618_n 0.00180746f $X=1.28 $Y=1.835 $X2=0 $Y2=0
cc_386 N_VPWR_c_503_n N_X_c_618_n 0.0129403f $X=1.42 $Y=2.27 $X2=0 $Y2=0
cc_387 N_VPWR_c_504_n N_X_c_686_n 0.0149362f $X=2.15 $Y=3.33 $X2=0 $Y2=0
cc_388 N_VPWR_c_501_n N_X_c_686_n 0.0100304f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_389 N_VPWR_M1008_s N_X_c_619_n 0.00180746f $X=2.14 $Y=1.835 $X2=0 $Y2=0
cc_390 N_VPWR_c_505_n N_X_c_619_n 0.0129403f $X=2.28 $Y=2.27 $X2=0 $Y2=0
cc_391 N_VPWR_c_516_n N_X_c_690_n 0.0149362f $X=3.01 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_c_501_n N_X_c_690_n 0.0100304f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_M1016_s N_X_c_620_n 0.00180746f $X=3 $Y=1.835 $X2=0 $Y2=0
cc_394 N_VPWR_c_506_n N_X_c_620_n 0.0129403f $X=3.14 $Y=2.27 $X2=0 $Y2=0
cc_395 N_VPWR_c_517_n N_X_c_694_n 0.0136943f $X=3.835 $Y=3.33 $X2=0 $Y2=0
cc_396 N_VPWR_c_501_n N_X_c_694_n 0.00866972f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_397 N_X_c_607_n N_VGND_M1002_d 0.00234752f $X=0.895 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_398 N_X_c_608_n N_VGND_M1009_d 0.00176461f $X=1.755 $Y=1.14 $X2=0 $Y2=0
cc_399 N_X_c_609_n N_VGND_M1013_d 0.00176461f $X=2.615 $Y=1.14 $X2=0 $Y2=0
cc_400 N_X_c_610_n N_VGND_M1020_d 0.00176461f $X=3.475 $Y=1.14 $X2=0 $Y2=0
cc_401 N_X_c_607_n N_VGND_c_717_n 0.0212047f $X=0.895 $Y=1.14 $X2=0 $Y2=0
cc_402 N_X_c_614_n N_VGND_c_717_n 8.43278e-19 $X=0.245 $Y=1.225 $X2=0 $Y2=0
cc_403 N_X_c_608_n N_VGND_c_718_n 0.0170777f $X=1.755 $Y=1.14 $X2=0 $Y2=0
cc_404 N_X_c_703_p N_VGND_c_719_n 0.0101681f $X=1.85 $Y=0.455 $X2=0 $Y2=0
cc_405 N_X_c_609_n N_VGND_c_720_n 0.0170777f $X=2.615 $Y=1.14 $X2=0 $Y2=0
cc_406 N_X_c_610_n N_VGND_c_721_n 0.0170777f $X=3.475 $Y=1.14 $X2=0 $Y2=0
cc_407 N_X_c_706_p N_VGND_c_727_n 0.0101681f $X=0.99 $Y=0.455 $X2=0 $Y2=0
cc_408 N_X_c_707_p N_VGND_c_731_n 0.0101681f $X=2.71 $Y=0.455 $X2=0 $Y2=0
cc_409 N_X_c_708_p N_VGND_c_732_n 0.0101681f $X=3.57 $Y=0.455 $X2=0 $Y2=0
cc_410 N_X_M1002_s N_VGND_c_735_n 0.00546338f $X=0.85 $Y=0.245 $X2=0 $Y2=0
cc_411 N_X_M1012_s N_VGND_c_735_n 0.00546338f $X=1.71 $Y=0.245 $X2=0 $Y2=0
cc_412 N_X_M1017_s N_VGND_c_735_n 0.00546338f $X=2.57 $Y=0.245 $X2=0 $Y2=0
cc_413 N_X_M1022_s N_VGND_c_735_n 0.00546338f $X=3.43 $Y=0.245 $X2=0 $Y2=0
cc_414 N_X_c_706_p N_VGND_c_735_n 0.00718296f $X=0.99 $Y=0.455 $X2=0 $Y2=0
cc_415 N_X_c_703_p N_VGND_c_735_n 0.00718296f $X=1.85 $Y=0.455 $X2=0 $Y2=0
cc_416 N_X_c_707_p N_VGND_c_735_n 0.00718296f $X=2.71 $Y=0.455 $X2=0 $Y2=0
cc_417 N_X_c_708_p N_VGND_c_735_n 0.00718296f $X=3.57 $Y=0.455 $X2=0 $Y2=0
