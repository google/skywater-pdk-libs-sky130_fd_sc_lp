* File: sky130_fd_sc_lp__clkbuflp_2.pex.spice
* Created: Wed Sep  2 09:39:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_2%A 1 3 6 8 10 11 12 19
r39 19 20 17.2143 $w=3.22e-07 $l=1.15e-07 $layer=POLY_cond $X=0.72 $Y=0.94
+ $X2=0.835 $Y2=0.94
r40 17 19 5.98758 $w=3.22e-07 $l=4e-08 $layer=POLY_cond $X=0.68 $Y=0.94 $X2=0.72
+ $Y2=0.94
r41 15 17 30.6863 $w=3.22e-07 $l=2.05e-07 $layer=POLY_cond $X=0.475 $Y=0.94
+ $X2=0.68 $Y2=0.94
r42 11 12 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=0.68 $Y=0.94 $X2=1.2
+ $Y2=0.94
r43 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=0.94 $X2=0.68 $Y2=0.94
r44 8 20 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=0.775
+ $X2=0.835 $Y2=0.94
r45 8 10 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.835 $Y=0.775
+ $X2=0.835 $Y2=0.445
r46 4 19 8.77827 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.105
+ $X2=0.72 $Y2=0.94
r47 4 6 367.711 $w=2.5e-07 $l=1.48e-06 $layer=POLY_cond $X=0.72 $Y=1.105
+ $X2=0.72 $Y2=2.585
r48 1 15 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.775
+ $X2=0.475 $Y2=0.94
r49 1 3 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.475 $Y=0.775
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_2%A_27_47# 1 2 9 13 17 21 25 29 33 37 43 46
+ 56
r75 55 56 61.0986 $w=3.4e-07 $l=3.6e-07 $layer=POLY_cond $X=2.055 $Y=1.375
+ $X2=2.415 $Y2=1.375
r76 54 55 46.6725 $w=3.4e-07 $l=2.75e-07 $layer=POLY_cond $X=1.78 $Y=1.375
+ $X2=2.055 $Y2=1.375
r77 53 54 26.3063 $w=3.4e-07 $l=1.55e-07 $layer=POLY_cond $X=1.625 $Y=1.375
+ $X2=1.78 $Y2=1.375
r78 52 53 61.0986 $w=3.4e-07 $l=3.6e-07 $layer=POLY_cond $X=1.265 $Y=1.375
+ $X2=1.625 $Y2=1.375
r79 51 52 2.54577 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=1.25 $Y=1.375
+ $X2=1.265 $Y2=1.375
r80 46 48 11.0966 $w=5.23e-07 $l=4.15e-07 $layer=LI1_cond $X=0.357 $Y=1.405
+ $X2=0.357 $Y2=1.82
r81 46 47 5.55122 $w=5.23e-07 $l=1.3e-07 $layer=LI1_cond $X=0.357 $Y=1.405
+ $X2=0.357 $Y2=1.275
r82 44 51 5.09155 $w=3.4e-07 $l=3e-08 $layer=POLY_cond $X=1.22 $Y=1.375 $X2=1.25
+ $Y2=1.375
r83 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.38 $X2=1.22 $Y2=1.38
r84 41 46 4.85815 $w=2.6e-07 $l=2.63e-07 $layer=LI1_cond $X=0.62 $Y=1.405
+ $X2=0.357 $Y2=1.405
r85 41 43 26.5948 $w=2.58e-07 $l=6e-07 $layer=LI1_cond $X=0.62 $Y=1.405 $X2=1.22
+ $Y2=1.405
r86 37 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.455 $Y=2.23
+ $X2=0.455 $Y2=2.91
r87 37 48 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.455 $Y=2.23
+ $X2=0.455 $Y2=1.82
r88 33 47 34.3675 $w=2.78e-07 $l=8.35e-07 $layer=LI1_cond $X=0.235 $Y=0.44
+ $X2=0.235 $Y2=1.275
r89 27 56 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.415 $Y=1.205
+ $X2=2.415 $Y2=1.375
r90 27 29 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.415 $Y=1.205
+ $X2=2.415 $Y2=0.445
r91 23 55 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.055 $Y=1.205
+ $X2=2.055 $Y2=1.375
r92 23 25 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.055 $Y=1.205
+ $X2=2.055 $Y2=0.445
r93 19 54 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.78 $Y=1.545
+ $X2=1.78 $Y2=1.375
r94 19 21 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.78 $Y=1.545
+ $X2=1.78 $Y2=2.585
r95 15 53 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.625 $Y=1.205
+ $X2=1.625 $Y2=1.375
r96 15 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.625 $Y=1.205
+ $X2=1.625 $Y2=0.445
r97 11 52 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.265 $Y=1.205
+ $X2=1.265 $Y2=1.375
r98 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.265 $Y=1.205
+ $X2=1.265 $Y2=0.445
r99 7 51 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.25 $Y=1.545
+ $X2=1.25 $Y2=1.375
r100 7 9 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.25 $Y=1.545
+ $X2=1.25 $Y2=2.585
r101 2 39 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=2.085 $X2=0.455 $Y2=2.91
r102 2 37 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=2.085 $X2=0.455 $Y2=2.23
r103 1 33 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_2%VPWR 1 2 9 15 20 21 22 28 34 35 38
r33 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 32 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=3.33
+ $X2=2.045 $Y2=3.33
r37 32 34 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.21 $Y=3.33 $X2=3.12
+ $Y2=3.33
r38 28 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=3.33
+ $X2=2.045 $Y2=3.33
r39 28 30 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=3.33 $X2=1.68
+ $Y2=3.33
r40 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 22 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 20 25 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=0.72
+ $Y2=3.33
r45 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.985 $Y2=3.33
r46 19 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=0.985 $Y2=3.33
r48 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.045 $Y=2.23
+ $X2=2.045 $Y2=2.91
r49 13 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=3.245
+ $X2=2.045 $Y2=3.33
r50 13 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.045 $Y=3.245
+ $X2=2.045 $Y2=2.91
r51 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.985 $Y=2.23
+ $X2=0.985 $Y2=2.91
r52 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=3.245
+ $X2=0.985 $Y2=3.33
r53 7 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.985 $Y=3.245
+ $X2=0.985 $Y2=2.91
r54 2 18 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.085 $X2=2.045 $Y2=2.91
r55 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.085 $X2=2.045 $Y2=2.23
r56 1 12 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.845
+ $Y=2.085 $X2=0.985 $Y2=2.91
r57 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.845
+ $Y=2.085 $X2=0.985 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_2%X 1 2 9 13 14 15 16 33 46
r32 46 49 0.669135 $w=7.13e-07 $l=4e-08 $layer=LI1_cond $X=1.912 $Y=1.665
+ $X2=1.912 $Y2=1.705
r33 16 50 6.81426 $w=9.48e-07 $l=1.48e-07 $layer=LI1_cond $X=1.795 $Y=1.727
+ $X2=1.795 $Y2=1.875
r34 16 49 1.05701 $w=9.48e-07 $l=2.2e-08 $layer=LI1_cond $X=1.795 $Y=1.727
+ $X2=1.795 $Y2=1.705
r35 16 46 0.384752 $w=7.13e-07 $l=2.3e-08 $layer=LI1_cond $X=1.912 $Y=1.642
+ $X2=1.912 $Y2=1.665
r36 15 16 5.80474 $w=7.13e-07 $l=3.47e-07 $layer=LI1_cond $X=1.912 $Y=1.295
+ $X2=1.912 $Y2=1.642
r37 14 15 6.1895 $w=7.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.912 $Y=0.925
+ $X2=1.912 $Y2=1.295
r38 13 14 6.1895 $w=7.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.912 $Y=0.555
+ $X2=1.912 $Y2=0.925
r39 13 33 1.92376 $w=7.13e-07 $l=1.15e-07 $layer=LI1_cond $X=1.912 $Y=0.555
+ $X2=1.912 $Y2=0.44
r40 9 11 21.7684 $w=3.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.5 $Y=2.23 $X2=1.5
+ $Y2=2.91
r41 9 50 11.3644 $w=3.58e-07 $l=3.55e-07 $layer=LI1_cond $X=1.5 $Y=2.23 $X2=1.5
+ $Y2=1.875
r42 2 11 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.375
+ $Y=2.085 $X2=1.515 $Y2=2.91
r43 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.375
+ $Y=2.085 $X2=1.515 $Y2=2.23
r44 1 33 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=1.84 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_2%VGND 1 2 9 13 15 17 22 29 30 33 36
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r44 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.63
+ $Y2=0
r46 27 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.12
+ $Y2=0
r47 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r48 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=0 $X2=1.05
+ $Y2=0
r50 23 25 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=1.215 $Y=0 $X2=2.16
+ $Y2=0
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.63
+ $Y2=0
r52 22 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.16
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r54 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.05
+ $Y2=0
r56 17 19 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.72
+ $Y2=0
r57 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 15 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r60 11 13 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.44
r61 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.085 $X2=1.05
+ $Y2=0
r62 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.05 $Y=0.085
+ $X2=1.05 $Y2=0.44
r63 2 13 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.235 $X2=2.63 $Y2=0.44
r64 1 9 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.44
.ends

