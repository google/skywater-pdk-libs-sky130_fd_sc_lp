* File: sky130_fd_sc_lp__nor4b_2.pex.spice
* Created: Wed Sep  2 10:11:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4B_2%D_N 3 5 7 8 13
r27 13 14 8.55161 $w=3.1e-07 $l=5.5e-08 $layer=POLY_cond $X=0.475 $Y=1.35
+ $X2=0.53 $Y2=1.35
r28 11 13 31.8742 $w=3.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.35
+ $X2=0.475 $Y2=1.35
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.35 $X2=0.27 $Y2=1.35
r30 5 14 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.185
+ $X2=0.53 $Y2=1.35
r31 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.53 $Y=1.185 $X2=0.53
+ $Y2=0.865
r32 1 13 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=1.35
r33 1 3 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%C 1 3 6 10 13 15 16 19 25 30 31 32 35
c89 32 0 3.33133e-20 $X=2.795 $Y=1.185
c90 31 0 3.38577e-19 $X=2.795 $Y=1.35
c91 30 0 7.14239e-20 $X=2.795 $Y=1.35
r92 30 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.35
+ $X2=2.795 $Y2=1.515
r93 30 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.35
+ $X2=2.795 $Y2=1.185
r94 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.35 $X2=2.795 $Y2=1.35
r95 25 31 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.64 $Y=1.3
+ $X2=2.795 $Y2=1.3
r96 25 35 8.38288 $w=4.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=1.3 $X2=2.49
+ $Y2=1.3
r97 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.35 $X2=0.98 $Y2=1.35
r98 19 22 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=0.965 $Y=1.17
+ $X2=0.965 $Y2=1.35
r99 18 19 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.065 $Y=1.17 $X2=0.965
+ $Y2=1.17
r100 18 35 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=1.065 $Y=1.17
+ $X2=2.49 $Y2=1.17
r101 15 23 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.41 $Y=1.35
+ $X2=0.98 $Y2=1.35
r102 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.35
+ $X2=1.485 $Y2=1.35
r103 13 33 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.775 $Y=2.465
+ $X2=2.775 $Y2=1.515
r104 10 32 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.775 $Y=0.655
+ $X2=2.775 $Y2=1.185
r105 4 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.515
+ $X2=1.485 $Y2=1.35
r106 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.485 $Y=1.515
+ $X2=1.485 $Y2=2.465
r107 1 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.485 $Y2=1.35
r108 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.485 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%A_27_535# 1 2 9 13 17 21 25 27 32 33 34 35
+ 37 50
c86 37 0 7.14239e-20 $X=2.155 $Y=1.51
r87 38 50 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.155 $Y=1.51
+ $X2=2.345 $Y2=1.51
r88 38 47 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=2.155 $Y=1.51
+ $X2=1.915 $Y2=1.51
r89 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.155
+ $Y=1.51 $X2=2.155 $Y2=1.51
r90 35 45 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.33 $Y=1.53
+ $X2=1.33 $Y2=1.78
r91 35 37 39.0823 $w=2.08e-07 $l=7.4e-07 $layer=LI1_cond $X=1.415 $Y=1.53
+ $X2=2.155 $Y2=1.53
r92 34 42 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.78
+ $X2=0.61 $Y2=1.78
r93 33 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=1.78
+ $X2=1.33 $Y2=1.78
r94 33 34 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.245 $Y=1.78
+ $X2=0.695 $Y2=1.78
r95 32 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.695
+ $X2=0.61 $Y2=1.78
r96 31 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.61 $Y=1.005
+ $X2=0.61 $Y2=1.695
r97 27 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.525 $Y=0.9
+ $X2=0.61 $Y2=1.005
r98 27 29 11.0909 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=0.525 $Y=0.9
+ $X2=0.315 $Y2=0.9
r99 23 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.225 $Y=1.78
+ $X2=0.61 $Y2=1.78
r100 23 25 45.2112 $w=2.58e-07 $l=1.02e-06 $layer=LI1_cond $X=0.225 $Y=1.865
+ $X2=0.225 $Y2=2.885
r101 19 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.345 $Y=1.675
+ $X2=2.345 $Y2=1.51
r102 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.345 $Y=1.675
+ $X2=2.345 $Y2=2.465
r103 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.345 $Y=1.345
+ $X2=2.345 $Y2=1.51
r104 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.345 $Y=1.345
+ $X2=2.345 $Y2=0.655
r105 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.675
+ $X2=1.915 $Y2=1.51
r106 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.915 $Y=1.675
+ $X2=1.915 $Y2=2.465
r107 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.345
+ $X2=1.915 $Y2=1.51
r108 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.915 $Y=1.345
+ $X2=1.915 $Y2=0.655
r109 2 25 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.885
r110 1 29 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.655 $X2=0.315 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%B 3 7 9 11 14 16 19 24 25 32 37 40
c79 32 0 2.22562e-19 $X=3.515 $Y=1.51
c80 19 0 1.92271e-19 $X=3.495 $Y=1.51
c81 7 0 1.93207e-19 $X=3.515 $Y=0.655
c82 3 0 1.61991e-19 $X=3.285 $Y=2.465
r83 34 37 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.805 $Y=1.35
+ $X2=4.98 $Y2=1.35
r84 25 40 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=1.7
+ $X2=5.005 $Y2=1.615
r85 25 40 0.545894 $w=3.78e-07 $l=1.8e-08 $layer=LI1_cond $X=5.005 $Y=1.597
+ $X2=5.005 $Y2=1.615
r86 24 25 9.15889 $w=3.78e-07 $l=3.02e-07 $layer=LI1_cond $X=5.005 $Y=1.295
+ $X2=5.005 $Y2=1.597
r87 24 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.98
+ $Y=1.35 $X2=4.98 $Y2=1.35
r88 20 32 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.495 $Y=1.51
+ $X2=3.515 $Y2=1.51
r89 20 29 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.495 $Y=1.51
+ $X2=3.285 $Y2=1.51
r90 19 22 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=3.53 $Y=1.51 $X2=3.53
+ $Y2=1.7
r91 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.495
+ $Y=1.51 $X2=3.495 $Y2=1.51
r92 17 22 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.66 $Y=1.7 $X2=3.53
+ $Y2=1.7
r93 16 25 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.815 $Y=1.7
+ $X2=5.005 $Y2=1.7
r94 16 17 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=4.815 $Y=1.7
+ $X2=3.66 $Y2=1.7
r95 12 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.515
+ $X2=4.805 $Y2=1.35
r96 12 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.805 $Y=1.515
+ $X2=4.805 $Y2=2.465
r97 9 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.185
+ $X2=4.805 $Y2=1.35
r98 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.805 $Y=1.185
+ $X2=4.805 $Y2=0.655
r99 5 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.345
+ $X2=3.515 $Y2=1.51
r100 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.515 $Y=1.345
+ $X2=3.515 $Y2=0.655
r101 1 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.675
+ $X2=3.285 $Y2=1.51
r102 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.285 $Y=1.675
+ $X2=3.285 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%A 1 3 6 8 10 13 15 16 24
c51 6 0 4.32342e-19 $X=3.945 $Y=2.465
r52 22 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.285 $Y=1.35
+ $X2=4.375 $Y2=1.35
r53 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.285
+ $Y=1.35 $X2=4.285 $Y2=1.35
r54 19 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.945 $Y=1.35
+ $X2=4.285 $Y2=1.35
r55 16 23 13.486 $w=2.33e-07 $l=2.75e-07 $layer=LI1_cond $X=4.56 $Y=1.327
+ $X2=4.285 $Y2=1.327
r56 15 23 10.0532 $w=2.33e-07 $l=2.05e-07 $layer=LI1_cond $X=4.08 $Y=1.327
+ $X2=4.285 $Y2=1.327
r57 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.515
+ $X2=4.375 $Y2=1.35
r58 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.375 $Y=1.515
+ $X2=4.375 $Y2=2.465
r59 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.185
+ $X2=4.375 $Y2=1.35
r60 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.375 $Y=1.185
+ $X2=4.375 $Y2=0.655
r61 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.515
+ $X2=3.945 $Y2=1.35
r62 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.945 $Y=1.515
+ $X2=3.945 $Y2=2.465
r63 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.185
+ $X2=3.945 $Y2=1.35
r64 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.945 $Y=1.185
+ $X2=3.945 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%VPWR 1 2 9 11 16 17 19 24 33 37 44
c64 11 0 1.61991e-19 $X=4.935 $Y=2.56
r65 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r66 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r68 31 44 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=2.88 $Y2=3.33
r69 30 31 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r70 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 27 30 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 27 28 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 25 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r74 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 24 36 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=5.107 $Y2=3.33
r76 24 30 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r79 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r80 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 17 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.88 $Y2=3.33
r82 17 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r83 16 36 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.065 $Y=3.245
+ $X2=5.107 $Y2=3.33
r84 15 16 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=5.065 $Y=2.665
+ $X2=5.065 $Y2=3.245
r85 11 15 6.91731 $w=2.1e-07 $l=1.74786e-07 $layer=LI1_cond $X=4.935 $Y=2.56
+ $X2=5.065 $Y2=2.665
r86 11 13 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=4.935 $Y=2.56
+ $X2=4.16 $Y2=2.56
r87 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r88 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.885
r89 2 13 600 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=2.56
r90 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.675 $X2=0.69 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%A_229_367# 1 2 3 12 14 18 24 27 32 35 36
c58 36 0 7.71915e-20 $X=3.815 $Y=2.16
c59 18 0 1.52478e-19 $X=3.07 $Y=2.6
r60 35 36 8.76268 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=3.645 $Y=2.16
+ $X2=3.815 $Y2=2.16
r61 32 34 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.07 $Y=2.23
+ $X2=3.07 $Y2=2.4
r62 29 30 3.15992 $w=3.08e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=2.4 $X2=1.26
+ $Y2=2.485
r63 27 29 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=1.26 $Y=2.2 $X2=1.26
+ $Y2=2.4
r64 24 36 49.5962 $w=2.78e-07 $l=1.205e-06 $layer=LI1_cond $X=5.02 $Y=2.145
+ $X2=3.815 $Y2=2.145
r65 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=2.23
+ $X2=3.07 $Y2=2.23
r66 21 35 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.235 $Y=2.23
+ $X2=3.645 $Y2=2.23
r67 16 34 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=2.485
+ $X2=3.07 $Y2=2.4
r68 16 18 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.07 $Y=2.485
+ $X2=3.07 $Y2=2.6
r69 15 29 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.415 $Y=2.4
+ $X2=1.26 $Y2=2.4
r70 14 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=2.4
+ $X2=3.07 $Y2=2.4
r71 14 15 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=2.905 $Y=2.4
+ $X2=1.415 $Y2=2.4
r72 12 30 16.0586 $w=3.03e-07 $l=4.25e-07 $layer=LI1_cond $X=1.257 $Y=2.91
+ $X2=1.257 $Y2=2.485
r73 3 24 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.835 $X2=5.02 $Y2=2.17
r74 2 32 600 $w=1.7e-07 $l=4.92874e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.835 $X2=3.07 $Y2=2.23
r75 2 18 300 $w=1.7e-07 $l=8.68058e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=1.835 $X2=3.07 $Y2=2.6
r76 1 27 400 $w=1.7e-07 $l=4.22907e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.835 $X2=1.27 $Y2=2.2
r77 1 12 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.835 $X2=1.27 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%A_312_367# 1 2 11
r14 8 11 27.9183 $w=3.53e-07 $l=8.6e-07 $layer=LI1_cond $X=1.7 $Y=2.832 $X2=2.56
+ $Y2=2.832
r15 2 11 600 $w=1.7e-07 $l=1.05268e-06 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=2.82
r16 1 8 600 $w=1.7e-07 $l=1.05268e-06 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.835 $X2=1.7 $Y2=2.82
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%Y 1 2 3 4 5 16 18 20 24 26 28 31 34 36 37 40
+ 45 48 49 50 55 64 66
c94 31 0 1.20906e-19 $X=3.145 $Y=1.805
r95 55 64 2.54215 $w=3.38e-07 $l=7.5e-08 $layer=LI1_cond $X=2.565 $Y=1.975
+ $X2=2.64 $Y2=1.975
r96 50 66 5.92976 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=2.645 $Y=1.975
+ $X2=2.735 $Y2=1.975
r97 50 64 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=1.975
+ $X2=2.64 $Y2=1.975
r98 50 55 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.56 $Y=1.975
+ $X2=2.565 $Y2=1.975
r99 49 50 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=2.13 $Y=1.975
+ $X2=2.56 $Y2=1.975
r100 48 49 15.2529 $w=3.38e-07 $l=4.5e-07 $layer=LI1_cond $X=1.68 $Y=1.975
+ $X2=2.13 $Y2=1.975
r101 46 47 16.4865 $w=4.07e-07 $l=5.5e-07 $layer=LI1_cond $X=3.145 $Y=0.96
+ $X2=3.695 $Y2=0.96
r102 38 40 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=4.59 $Y=0.87
+ $X2=4.59 $Y2=0.43
r103 37 47 8.13703 $w=4.07e-07 $l=1.32476e-07 $layer=LI1_cond $X=3.825 $Y=0.955
+ $X2=3.695 $Y2=0.96
r104 36 38 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.495 $Y=0.955
+ $X2=4.59 $Y2=0.87
r105 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.495 $Y=0.955
+ $X2=3.825 $Y2=0.955
r106 32 47 3.35936 $w=2.6e-07 $l=2.15e-07 $layer=LI1_cond $X=3.695 $Y=0.745
+ $X2=3.695 $Y2=0.96
r107 32 34 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=3.695 $Y=0.745
+ $X2=3.695 $Y2=0.42
r108 30 46 5.88399 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.145 $Y=1.175
+ $X2=3.145 $Y2=0.96
r109 30 31 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.145 $Y=1.175
+ $X2=3.145 $Y2=1.805
r110 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=1.89
+ $X2=3.145 $Y2=1.805
r111 28 66 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.06 $Y=1.89
+ $X2=2.735 $Y2=1.89
r112 27 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.725 $Y=0.83
+ $X2=2.595 $Y2=0.83
r113 26 46 6.78813 $w=4.07e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.06 $Y=0.83
+ $X2=3.145 $Y2=0.96
r114 26 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.06 $Y=0.83
+ $X2=2.725 $Y2=0.83
r115 22 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.745
+ $X2=2.595 $Y2=0.83
r116 22 24 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=2.595 $Y=0.745
+ $X2=2.595 $Y2=0.42
r117 21 43 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.795 $Y=0.83
+ $X2=1.665 $Y2=0.83
r118 20 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.465 $Y=0.83
+ $X2=2.595 $Y2=0.83
r119 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.465 $Y=0.83
+ $X2=1.795 $Y2=0.83
r120 16 43 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.745
+ $X2=1.665 $Y2=0.83
r121 16 18 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=1.665 $Y=0.745
+ $X2=1.665 $Y2=0.42
r122 5 49 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.835 $X2=2.13 $Y2=1.98
r123 4 40 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=4.45
+ $Y=0.235 $X2=4.59 $Y2=0.43
r124 3 34 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.59
+ $Y=0.235 $X2=3.73 $Y2=0.42
r125 2 45 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.235 $X2=2.56 $Y2=0.83
r126 2 24 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.235 $X2=2.56 $Y2=0.42
r127 1 43 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.83
r128 1 18 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%A_672_367# 1 2 7 9 13
r24 11 16 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=3.77 $Y=2.955
+ $X2=3.605 $Y2=2.955
r25 11 13 39.3751 $w=2.38e-07 $l=8.2e-07 $layer=LI1_cond $X=3.77 $Y=2.955
+ $X2=4.59 $Y2=2.955
r26 7 16 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=3.605 $Y=2.835
+ $X2=3.605 $Y2=2.955
r27 7 9 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.605 $Y=2.835
+ $X2=3.605 $Y2=2.57
r28 2 13 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.45
+ $Y=1.835 $X2=4.59 $Y2=2.95
r29 1 16 600 $w=1.7e-07 $l=1.23142e-06 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.605 $Y2=2.95
r30 1 9 600 $w=1.7e-07 $l=8.48705e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.605 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_2%VGND 1 2 3 4 5 18 24 28 32 34 36 38 40 45 50
+ 55 60 66 69 72 75 79 87
r86 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r87 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r88 73 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.88
+ $Y2=0
r89 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r90 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r91 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 64 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r93 64 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r94 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r95 61 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.16
+ $Y2=0
r96 61 63 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.56
+ $Y2=0
r97 60 78 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=5.067
+ $Y2=0
r98 60 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=4.56
+ $Y2=0
r99 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r100 59 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r101 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r102 56 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.15
+ $Y2=0
r103 56 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.6
+ $Y2=0
r104 55 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.16
+ $Y2=0
r105 55 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.6
+ $Y2=0
r106 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.13
+ $Y2=0
r107 51 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.64
+ $Y2=0
r108 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=3.15
+ $Y2=0
r109 50 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.64
+ $Y2=0
r110 49 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r111 49 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r112 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r113 46 66 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.115
+ $Y2=0
r114 46 48 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=0
+ $X2=1.68 $Y2=0
r115 45 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=2.13
+ $Y2=0
r116 45 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=0
+ $X2=1.68 $Y2=0
r117 43 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r118 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r119 40 66 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.115
+ $Y2=0
r120 40 42 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.865 $Y=0
+ $X2=0.72 $Y2=0
r121 38 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.88 $Y2=0
r122 38 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r123 38 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r124 34 78 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=5.02 $Y=0.085
+ $X2=5.067 $Y2=0
r125 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.02 $Y=0.085
+ $X2=5.02 $Y2=0.38
r126 30 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=0.085
+ $X2=4.16 $Y2=0
r127 30 32 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.16 $Y=0.085
+ $X2=4.16 $Y2=0.575
r128 26 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=0.085
+ $X2=3.15 $Y2=0
r129 26 28 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.15 $Y=0.085
+ $X2=3.15 $Y2=0.45
r130 22 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0
r131 22 24 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0.45
r132 18 20 10.7647 $w=4.98e-07 $l=4.5e-07 $layer=LI1_cond $X=1.115 $Y=0.38
+ $X2=1.115 $Y2=0.83
r133 16 66 2.07448 $w=5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r134 16 18 7.05686 $w=4.98e-07 $l=2.95e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.38
r135 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.88
+ $Y=0.235 $X2=5.02 $Y2=0.38
r136 4 32 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.16 $Y2=0.575
r137 3 28 182 $w=1.7e-07 $l=3.93065e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.235 $X2=3.15 $Y2=0.45
r138 2 24 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.235 $X2=2.13 $Y2=0.45
r139 1 20 182 $w=1.7e-07 $l=5.04975e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.655 $X2=1.03 $Y2=0.83
r140 1 18 182 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.655 $X2=1.19 $Y2=0.38
.ends

