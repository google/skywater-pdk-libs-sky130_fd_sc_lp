* File: sky130_fd_sc_lp__o211ai_m.pxi.spice
* Created: Wed Sep  2 10:14:58 2020
* 
x_PM_SKY130_FD_SC_LP__O211AI_M%A1 N_A1_M1007_g N_A1_M1000_g N_A1_c_58_n
+ N_A1_c_62_n A1 A1 A1 A1 N_A1_c_60_n PM_SKY130_FD_SC_LP__O211AI_M%A1
x_PM_SKY130_FD_SC_LP__O211AI_M%A2 N_A2_M1002_g N_A2_M1004_g N_A2_c_91_n
+ N_A2_c_92_n A2 N_A2_c_94_n PM_SKY130_FD_SC_LP__O211AI_M%A2
x_PM_SKY130_FD_SC_LP__O211AI_M%B1 N_B1_M1005_g N_B1_M1003_g N_B1_c_134_n
+ N_B1_c_135_n B1 N_B1_c_132_n PM_SKY130_FD_SC_LP__O211AI_M%B1
x_PM_SKY130_FD_SC_LP__O211AI_M%C1 N_C1_c_176_n N_C1_M1006_g N_C1_M1001_g C1
+ N_C1_c_179_n PM_SKY130_FD_SC_LP__O211AI_M%C1
x_PM_SKY130_FD_SC_LP__O211AI_M%VPWR N_VPWR_M1000_s N_VPWR_M1003_d N_VPWR_c_210_n
+ N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_213_n VPWR N_VPWR_c_214_n
+ N_VPWR_c_215_n N_VPWR_c_209_n N_VPWR_c_217_n PM_SKY130_FD_SC_LP__O211AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O211AI_M%Y N_Y_M1006_d N_Y_M1004_d N_Y_M1001_d N_Y_c_257_n
+ N_Y_c_252_n N_Y_c_253_n N_Y_c_247_n N_Y_c_248_n N_Y_c_249_n N_Y_c_250_n
+ N_Y_c_254_n Y Y Y Y Y PM_SKY130_FD_SC_LP__O211AI_M%Y
x_PM_SKY130_FD_SC_LP__O211AI_M%A_29_47# N_A_29_47#_M1007_s N_A_29_47#_M1002_d
+ N_A_29_47#_c_314_n N_A_29_47#_c_315_n N_A_29_47#_c_316_n N_A_29_47#_c_325_n
+ PM_SKY130_FD_SC_LP__O211AI_M%A_29_47#
x_PM_SKY130_FD_SC_LP__O211AI_M%VGND N_VGND_M1007_d N_VGND_c_340_n VGND
+ N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n N_VGND_c_344_n
+ PM_SKY130_FD_SC_LP__O211AI_M%VGND
cc_1 VNB N_A1_M1007_g 0.0610873f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.445
cc_2 VNB N_A1_c_58_n 0.0178258f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.475
cc_3 VNB A1 0.0200286f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_60_n 0.014792f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.49
cc_5 VNB N_A2_M1002_g 0.0241948f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.445
cc_6 VNB N_A2_M1004_g 0.00272325f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.885
cc_7 VNB N_A2_c_91_n 0.0187158f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.475
cc_8 VNB N_A2_c_92_n 0.0201542f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.92
cc_9 VNB A2 0.0177014f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_10 VNB N_A2_c_94_n 0.0147303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_M1005_g 0.0624334f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.445
cc_12 VNB N_B1_c_132_n 0.0081233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C1_c_176_n 0.0213169f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.325
cc_14 VNB N_C1_M1001_g 0.0383229f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.885
cc_15 VNB C1 0.00939502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_c_179_n 0.053116f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.475
cc_17 VNB N_VPWR_c_209_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_247_n 0.0108932f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_Y_c_248_n 0.0131112f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB N_Y_c_249_n 0.00364419f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_21 VNB N_Y_c_250_n 0.00201845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.0120222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_29_47#_c_314_n 4.12885e-19 $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.475
cc_24 VNB N_A_29_47#_c_315_n 0.0153763f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.475
cc_25 VNB N_A_29_47#_c_316_n 0.00951254f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.92
cc_26 VNB N_VGND_c_340_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.885
cc_27 VNB N_VGND_c_341_n 0.0163548f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.325
cc_28 VNB N_VGND_c_342_n 0.0423134f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_29 VNB N_VGND_c_343_n 0.154644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_344_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_A1_M1000_g 0.0534677f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.885
cc_32 VPB N_A1_c_62_n 0.0384831f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.92
cc_33 VPB A1 0.0443735f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB N_A1_c_60_n 0.0165534f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.49
cc_35 VPB N_A2_M1004_g 0.0622385f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.885
cc_36 VPB N_B1_M1003_g 0.0298274f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.885
cc_37 VPB N_B1_c_134_n 0.0187158f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.475
cc_38 VPB N_B1_c_135_n 0.014967f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.92
cc_39 VPB B1 0.0116523f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.845
cc_40 VPB N_B1_c_132_n 0.00814006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_C1_M1001_g 0.0758773f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.885
cc_42 VPB N_VPWR_c_210_n 0.01277f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.475
cc_43 VPB N_VPWR_c_211_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.845
cc_44 VPB N_VPWR_c_212_n 0.0112126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_213_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_46 VPB N_VPWR_c_214_n 0.0243979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_215_n 0.0160358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_209_n 0.0495773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_217_n 0.00436274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_Y_c_252_n 0.00850348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_Y_c_253_n 0.00928935f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.92
cc_52 VPB N_Y_c_254_n 0.00781329f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.295
cc_53 VPB Y 0.0328522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB Y 4.12885e-19 $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.665
cc_55 N_A1_M1007_g N_A2_M1002_g 0.0190584f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_56 N_A1_c_62_n N_A2_M1004_g 0.0862219f $X=0.665 $Y=1.92 $X2=0 $Y2=0
cc_57 A1 N_A2_M1004_g 0.00176296f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A1_c_60_n N_A2_M1004_g 0.00804067f $X=0.385 $Y=1.49 $X2=0 $Y2=0
cc_59 N_A1_c_58_n N_A2_c_91_n 0.016712f $X=0.39 $Y=1.475 $X2=0 $Y2=0
cc_60 A1 N_A2_c_91_n 3.4658e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 A1 N_A2_c_92_n 4.78123e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A1_c_60_n N_A2_c_92_n 0.00817153f $X=0.385 $Y=1.49 $X2=0 $Y2=0
cc_63 N_A1_M1007_g A2 0.00221453f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_64 A1 A2 0.0154082f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A1_M1007_g N_A2_c_94_n 0.016712f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A1_M1000_g N_VPWR_c_210_n 0.0113246f $X=0.665 $Y=2.885 $X2=0 $Y2=0
cc_67 A1 N_VPWR_c_210_n 0.00865755f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A1_M1000_g N_VPWR_c_214_n 0.00486043f $X=0.665 $Y=2.885 $X2=0 $Y2=0
cc_69 N_A1_M1000_g N_VPWR_c_209_n 0.00818711f $X=0.665 $Y=2.885 $X2=0 $Y2=0
cc_70 A1 N_VPWR_c_209_n 0.00612305f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A1_M1007_g N_A_29_47#_c_314_n 3.64605e-19 $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A1_M1007_g N_A_29_47#_c_315_n 0.0163081f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_73 A1 N_A_29_47#_c_315_n 0.00405873f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A1_c_58_n N_A_29_47#_c_316_n 8.48361e-19 $X=0.39 $Y=1.475 $X2=0 $Y2=0
cc_75 A1 N_A_29_47#_c_316_n 0.0110656f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A1_M1007_g N_VGND_c_340_n 0.00998194f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A1_M1007_g N_VGND_c_341_n 0.00414412f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_78 N_A1_M1007_g N_VGND_c_343_n 0.0058521f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A2_M1002_g N_B1_M1005_g 0.0219875f $X=0.955 $Y=0.445 $X2=0 $Y2=0
cc_80 A2 N_B1_M1005_g 0.00530725f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A2_c_94_n N_B1_M1005_g 0.0208367f $X=0.935 $Y=1.1 $X2=0 $Y2=0
cc_82 N_A2_M1004_g N_B1_M1003_g 0.0275303f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_83 N_A2_c_92_n N_B1_c_134_n 0.0208367f $X=0.935 $Y=1.605 $X2=0 $Y2=0
cc_84 N_A2_M1004_g N_B1_c_135_n 0.0208367f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_85 N_A2_M1004_g B1 0.00336917f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_86 N_A2_c_91_n N_B1_c_132_n 0.0208367f $X=0.935 $Y=1.44 $X2=0 $Y2=0
cc_87 N_A2_M1004_g N_VPWR_c_210_n 0.00207709f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_88 N_A2_M1004_g N_VPWR_c_211_n 0.00148579f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_89 N_A2_M1004_g N_VPWR_c_214_n 0.00585385f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_90 N_A2_M1004_g N_VPWR_c_209_n 0.0108402f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_91 N_A2_M1004_g N_Y_c_257_n 2.1266e-19 $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_92 N_A2_M1004_g N_Y_c_253_n 0.00551383f $X=1.025 $Y=2.885 $X2=0 $Y2=0
cc_93 A2 N_Y_c_247_n 0.0124773f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 A2 N_Y_c_249_n 0.0130953f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 A2 Y 0.00442066f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A2_M1002_g N_A_29_47#_c_315_n 0.0116442f $X=0.955 $Y=0.445 $X2=0 $Y2=0
cc_97 A2 N_A_29_47#_c_315_n 0.03917f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_98 N_A2_c_94_n N_A_29_47#_c_315_n 0.00515085f $X=0.935 $Y=1.1 $X2=0 $Y2=0
cc_99 N_A2_M1002_g N_A_29_47#_c_325_n 2.1266e-19 $X=0.955 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A2_M1002_g N_VGND_c_340_n 0.00741705f $X=0.955 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A2_M1002_g N_VGND_c_342_n 0.00414412f $X=0.955 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A2_M1002_g N_VGND_c_343_n 0.00486498f $X=0.955 $Y=0.445 $X2=0 $Y2=0
cc_103 N_B1_M1005_g N_C1_c_176_n 0.0484827f $X=1.385 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_104 N_B1_M1003_g N_C1_M1001_g 0.0224633f $X=1.455 $Y=2.885 $X2=0 $Y2=0
cc_105 B1 N_C1_M1001_g 0.00330273f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_106 N_B1_c_132_n N_C1_M1001_g 0.0401351f $X=1.475 $Y=1.79 $X2=0 $Y2=0
cc_107 N_B1_M1005_g N_C1_c_179_n 0.0183974f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B1_M1003_g N_VPWR_c_211_n 0.00740843f $X=1.455 $Y=2.885 $X2=0 $Y2=0
cc_109 N_B1_M1003_g N_VPWR_c_214_n 0.00414412f $X=1.455 $Y=2.885 $X2=0 $Y2=0
cc_110 N_B1_M1003_g N_VPWR_c_209_n 0.00486498f $X=1.455 $Y=2.885 $X2=0 $Y2=0
cc_111 N_B1_M1003_g N_Y_c_257_n 2.1266e-19 $X=1.455 $Y=2.885 $X2=0 $Y2=0
cc_112 N_B1_M1003_g N_Y_c_252_n 0.0122727f $X=1.455 $Y=2.885 $X2=0 $Y2=0
cc_113 N_B1_c_135_n N_Y_c_252_n 0.00381935f $X=1.475 $Y=2.295 $X2=0 $Y2=0
cc_114 B1 N_Y_c_252_n 0.0224396f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_115 N_B1_c_135_n N_Y_c_253_n 9.65395e-19 $X=1.475 $Y=2.295 $X2=0 $Y2=0
cc_116 B1 N_Y_c_253_n 0.00204221f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_117 N_B1_M1005_g N_Y_c_247_n 0.00736205f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_118 B1 N_Y_c_248_n 0.00480633f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_119 N_B1_M1005_g N_Y_c_249_n 0.0017889f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_120 B1 N_Y_c_249_n 0.00897632f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_121 N_B1_c_132_n N_Y_c_249_n 0.00370524f $X=1.475 $Y=1.79 $X2=0 $Y2=0
cc_122 N_B1_M1005_g N_Y_c_250_n 0.00111799f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B1_M1005_g Y 0.00101703f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_124 N_B1_M1003_g Y 0.00100823f $X=1.455 $Y=2.885 $X2=0 $Y2=0
cc_125 N_B1_c_134_n Y 2.15931e-19 $X=1.475 $Y=2.13 $X2=0 $Y2=0
cc_126 N_B1_c_135_n Y 4.64927e-19 $X=1.475 $Y=2.295 $X2=0 $Y2=0
cc_127 B1 Y 0.0393967f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_128 N_B1_c_132_n Y 6.80858e-19 $X=1.475 $Y=1.79 $X2=0 $Y2=0
cc_129 N_B1_M1005_g N_A_29_47#_c_315_n 0.00163086f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_130 N_B1_M1005_g N_VGND_c_340_n 0.00146097f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_131 N_B1_M1005_g N_VGND_c_342_n 0.00585385f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_132 N_B1_M1005_g N_VGND_c_343_n 0.0108402f $X=1.385 $Y=0.445 $X2=0 $Y2=0
cc_133 N_C1_M1001_g N_VPWR_c_211_n 0.00998194f $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_134 N_C1_M1001_g N_VPWR_c_215_n 0.00414359f $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_135 N_C1_M1001_g N_VPWR_c_209_n 0.00584114f $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_136 N_C1_M1001_g N_Y_c_252_n 0.00994076f $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_137 N_C1_c_176_n N_Y_c_247_n 0.00512909f $X=1.745 $Y=0.765 $X2=0 $Y2=0
cc_138 C1 N_Y_c_247_n 0.012684f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_139 N_C1_c_179_n N_Y_c_247_n 0.00429105f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_140 N_C1_M1001_g N_Y_c_248_n 0.0137536f $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_141 C1 N_Y_c_248_n 0.0190454f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_142 N_C1_c_179_n N_Y_c_248_n 0.00748624f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_143 N_C1_c_176_n N_Y_c_250_n 0.0113884f $X=1.745 $Y=0.765 $X2=0 $Y2=0
cc_144 C1 N_Y_c_250_n 0.0151733f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_145 N_C1_c_179_n N_Y_c_250_n 0.00674175f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_146 N_C1_M1001_g N_Y_c_254_n 0.00545025f $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_147 N_C1_M1001_g Y 0.040278f $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_148 C1 Y 0.00448395f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_149 N_C1_c_179_n Y 0.0012715f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_150 N_C1_M1001_g Y 3.64605e-19 $X=1.925 $Y=2.885 $X2=0 $Y2=0
cc_151 N_C1_c_176_n N_VGND_c_342_n 0.00373071f $X=1.745 $Y=0.765 $X2=0 $Y2=0
cc_152 N_C1_c_179_n N_VGND_c_342_n 0.00218039f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_153 N_C1_c_176_n N_VGND_c_343_n 0.00643757f $X=1.745 $Y=0.765 $X2=0 $Y2=0
cc_154 C1 N_VGND_c_343_n 0.0060984f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_155 N_C1_c_179_n N_VGND_c_343_n 0.00272466f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_156 N_VPWR_c_209_n A_148_535# 0.00899413f $X=2.16 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_157 N_VPWR_c_209_n N_Y_M1004_d 0.00369956f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_158 N_VPWR_c_209_n N_Y_M1001_d 0.00308519f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_214_n N_Y_c_257_n 0.0081737f $X=1.525 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_209_n N_Y_c_257_n 0.00762225f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_161 N_VPWR_c_211_n N_Y_c_252_n 0.0194898f $X=1.69 $Y=2.95 $X2=0 $Y2=0
cc_162 N_VPWR_c_214_n N_Y_c_252_n 0.002793f $X=1.525 $Y=3.33 $X2=0 $Y2=0
cc_163 N_VPWR_c_215_n N_Y_c_252_n 0.0013569f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_c_209_n N_Y_c_252_n 0.00783924f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_c_215_n N_Y_c_254_n 0.00158832f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VPWR_c_209_n N_Y_c_254_n 0.00238794f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_167 N_VPWR_c_215_n Y 0.00877924f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_209_n Y 0.00770513f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_169 N_Y_c_247_n N_A_29_47#_c_315_n 0.0117746f $X=1.585 $Y=1.195 $X2=0 $Y2=0
cc_170 N_Y_c_247_n N_A_29_47#_c_325_n 2.82212e-19 $X=1.585 $Y=1.195 $X2=0 $Y2=0
cc_171 N_Y_c_250_n N_A_29_47#_c_325_n 2.07669e-19 $X=1.96 $Y=0.495 $X2=0 $Y2=0
cc_172 N_Y_c_250_n N_VGND_c_342_n 0.0223833f $X=1.96 $Y=0.495 $X2=0 $Y2=0
cc_173 N_Y_M1006_d N_VGND_c_343_n 0.00234714f $X=1.82 $Y=0.235 $X2=0 $Y2=0
cc_174 N_Y_c_250_n N_VGND_c_343_n 0.019907f $X=1.96 $Y=0.495 $X2=0 $Y2=0
cc_175 N_Y_c_250_n A_292_47# 0.00107385f $X=1.96 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_176 N_A_29_47#_c_315_n N_VGND_c_340_n 0.0194898f $X=1.065 $Y=0.75 $X2=0 $Y2=0
cc_177 N_A_29_47#_c_314_n N_VGND_c_341_n 0.0085932f $X=0.27 $Y=0.51 $X2=0 $Y2=0
cc_178 N_A_29_47#_c_315_n N_VGND_c_341_n 0.002793f $X=1.065 $Y=0.75 $X2=0 $Y2=0
cc_179 N_A_29_47#_c_315_n N_VGND_c_342_n 0.002793f $X=1.065 $Y=0.75 $X2=0 $Y2=0
cc_180 N_A_29_47#_c_325_n N_VGND_c_342_n 0.0081737f $X=1.17 $Y=0.51 $X2=0 $Y2=0
cc_181 N_A_29_47#_M1007_s N_VGND_c_343_n 0.0030857f $X=0.145 $Y=0.235 $X2=0
+ $Y2=0
cc_182 N_A_29_47#_M1002_d N_VGND_c_343_n 0.00369956f $X=1.03 $Y=0.235 $X2=0
+ $Y2=0
cc_183 N_A_29_47#_c_314_n N_VGND_c_343_n 0.00762225f $X=0.27 $Y=0.51 $X2=0 $Y2=0
cc_184 N_A_29_47#_c_315_n N_VGND_c_343_n 0.0100753f $X=1.065 $Y=0.75 $X2=0 $Y2=0
cc_185 N_A_29_47#_c_325_n N_VGND_c_343_n 0.00762225f $X=1.17 $Y=0.51 $X2=0 $Y2=0
cc_186 N_VGND_c_343_n A_292_47# 0.00310179f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
