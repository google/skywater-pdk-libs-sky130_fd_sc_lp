* File: sky130_fd_sc_lp__sdfrtp_lp2.spice
* Created: Fri Aug 28 11:28:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrtp_lp2.pex.spice"
.subckt sky130_fd_sc_lp__sdfrtp_lp2  VNB VPB D SCE SCD CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* SCE	SCE
* D	D
* VPB	VPB
* VNB	VNB
MM1000 noxref_24 N_A_81_194#_M1000_g N_noxref_23_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.22145 PD=0.66 PS=2.04 NRD=18.564 NRS=134.928 M=1 R=2.8
+ SA=75000.3 SB=75003 A=0.063 P=1.14 MULT=1
MM1043 N_A_116_419#_M1043_d N_D_M1043_g noxref_24 VNB NSHORT L=0.15 W=0.42
+ AD=0.101825 AS=0.0504 PD=0.925 PS=0.66 NRD=24.276 NRS=18.564 M=1 R=2.8
+ SA=75000.7 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1010 noxref_25 N_SCE_M1010_g N_A_116_419#_M1043_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.101825 PD=0.66 PS=0.925 NRD=18.564 NRS=24.276 M=1 R=2.8
+ SA=75001.3 SB=75002 A=0.063 P=1.14 MULT=1
MM1044 N_noxref_23_M1044_d N_SCD_M1044_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_RESET_B_M1011_g N_noxref_23_M1044_d VNB NSHORT L=0.15
+ W=0.42 AD=0.227 AS=0.0588 PD=1.405 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1025 A_697_119# N_SCE_M1025_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.227 PD=0.63 PS=1.405 NRD=14.28 NRS=135.708 M=1 R=2.8 SA=75002.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_81_194#_M1013_d N_SCE_M1013_g A_697_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_959_119# N_CLK_M1015_g N_A_876_119#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_CLK_M1032_g A_959_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1127 AS=0.0441 PD=1 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1029 A_1149_119# N_A_876_119#_M1029_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1127 PD=0.63 PS=1 NRD=14.28 NRS=24.276 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1038 N_A_1147_408#_M1038_d N_A_876_119#_M1038_g A_1149_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_1432_119#_M1014_d N_A_876_119#_M1014_g N_A_116_419#_M1014_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.10395 AS=0.1197 PD=0.915 PS=1.41 NRD=0 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1008 A_1561_119# N_A_1147_408#_M1008_g N_A_1432_119#_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0462 AS=0.10395 PD=0.64 PS=0.915 NRD=15.708 NRS=61.428 M=1 R=2.8
+ SA=75000.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1026 A_1635_119# N_A_1605_93#_M1026_g A_1561_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1411 AS=0.0462 PD=1.155 PS=0.64 NRD=80.268 NRS=15.708 M=1 R=2.8
+ SA=75001.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_RESET_B_M1021_g A_1635_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.150287 AS=0.1411 PD=1.17 PS=1.155 NRD=24.276 NRS=80.268 M=1 R=2.8
+ SA=75000.9 SB=75004 A=0.063 P=1.14 MULT=1
MM1022 A_1900_47# N_A_1432_119#_M1022_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.150287 PD=0.66 PS=1.17 NRD=18.564 NRS=57.132 M=1 R=2.8
+ SA=75001.1 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1033 N_A_1605_93#_M1033_d N_A_1432_119#_M1033_g A_1900_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75004 A=0.063 P=1.14 MULT=1
MM1039 N_A_2092_47#_M1039_d N_A_1147_408#_M1039_g N_A_1605_93#_M1033_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.29085 AS=0.0882 PD=1.805 PS=0.84 NRD=307.14 NRS=0
+ M=1 R=2.8 SA=75002.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1020 A_2399_47# N_A_876_119#_M1020_g N_A_2092_47#_M1039_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.29085 PD=0.81 PS=1.805 NRD=39.996 NRS=8.568 M=1 R=2.8
+ SA=75003.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_A_2435_296#_M1034_g A_2399_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0819 PD=1.04 PS=0.81 NRD=35.712 NRS=39.996 M=1 R=2.8 SA=75004.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 A_2661_47# N_RESET_B_M1012_g N_VGND_M1034_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1302 PD=0.66 PS=1.04 NRD=18.564 NRS=61.428 M=1 R=2.8 SA=75004.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_A_2435_296#_M1027_d N_A_2092_47#_M1027_g A_2661_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75005.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 A_2950_90# N_A_2092_47#_M1035_g N_A_2863_90#_M1035_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_2092_47#_M1017_g A_2950_90# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1040 A_3108_90# N_A_2863_90#_M1040_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1036 N_Q_M1036_d N_A_2863_90#_M1036_g A_3108_90# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_223_419# N_D_M1001_g N_A_116_419#_M1001_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1018 N_VPWR_M1018_d N_SCE_M1018_g A_223_419# VPB PHIGHVT L=0.25 W=1 AD=0.17
+ AS=0.12 PD=1.34 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1041 A_439_419# N_SCD_M1041_g N_VPWR_M1018_d VPB PHIGHVT L=0.25 W=1 AD=0.135
+ AS=0.17 PD=1.27 PS=1.34 NRD=15.7403 NRS=11.8003 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1030 N_A_116_419#_M1030_d N_A_81_194#_M1030_g A_439_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=15.7403 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_RESET_B_M1009_g N_A_116_419#_M1030_d VPB PHIGHVT L=0.25
+ W=1 AD=0.1825 AS=0.14 PD=1.365 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1023 N_A_81_194#_M1023_d N_SCE_M1023_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1825 PD=2.57 PS=1.365 NRD=0 NRS=16.7253 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1031 N_VPWR_M1031_d N_CLK_M1031_g N_A_876_119#_M1031_s VPB PHIGHVT L=0.25 W=1
+ AD=0.255 AS=0.285 PD=1.51 PS=2.57 NRD=45.2903 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1016 N_A_1147_408#_M1016_d N_A_876_119#_M1016_g N_VPWR_M1031_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.265 AS=0.255 PD=2.53 PS=1.51 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1019 N_A_1432_119#_M1019_d N_A_1147_408#_M1019_g N_A_116_419#_M1019_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.215 AS=0.3895 PD=1.43 PS=2.82 NRD=0 NRS=28.565 M=1 R=4
+ SA=125000 SB=125002 A=0.25 P=2.5 MULT=1
MM1042 A_1633_347# N_A_876_119#_M1042_g N_A_1432_119#_M1019_d VPB PHIGHVT L=0.25
+ W=1 AD=0.105 AS=0.215 PD=1.21 PS=1.43 NRD=9.8303 NRS=29.5303 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1045 N_VPWR_M1045_d N_A_1605_93#_M1045_g A_1633_347# VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1024 N_A_1432_119#_M1024_d N_RESET_B_M1024_g N_VPWR_M1045_d VPB PHIGHVT L=0.25
+ W=1 AD=0.43 AS=0.14 PD=2.86 PS=1.28 NRD=28.5453 NRS=0 M=1 R=4 SA=125002
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1006 N_A_1605_93#_M1006_d N_A_1432_119#_M1006_g N_VPWR_M1006_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.18 AS=0.285 PD=1.36 PS=2.57 NRD=15.7403 NRS=0 M=1 R=4
+ SA=125000 SB=125003 A=0.25 P=2.5 MULT=1
MM1002 N_A_2092_47#_M1002_d N_A_876_119#_M1002_g N_A_1605_93#_M1006_d VPB
+ PHIGHVT L=0.25 W=1 AD=0.27655 AS=0.18 PD=1.83 PS=1.36 NRD=15.7403 NRS=0 M=1
+ R=4 SA=125001 SB=125002 A=0.25 P=2.5 MULT=1
MM1037 A_2387_419# N_A_1147_408#_M1037_g N_A_2092_47#_M1002_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.27655 PD=1.24 PS=1.83 NRD=12.7853 NRS=15.7403 M=1 R=4
+ SA=125001 SB=125002 A=0.25 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_A_2435_296#_M1003_g A_2387_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.4225 AS=0.12 PD=1.845 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1028 N_A_2435_296#_M1028_d N_RESET_B_M1028_g N_VPWR_M1003_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.4225 PD=1.28 PS=1.845 NRD=0 NRS=111.285 M=1 R=4 SA=125003
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_2092_47#_M1004_g N_A_2435_296#_M1028_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_A_2092_47#_M1005_g N_A_2863_90#_M1005_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1007 N_Q_M1007_d N_A_2863_90#_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX46_noxref VNB VPB NWDIODE A=31.8065 P=37.39
c_281 VPB 0 2.64776e-19 $X=0 $Y=3.085
c_2300 A_1635_119# 0 1.52796e-19 $X=8.175 $Y=0.595
*
.include "sky130_fd_sc_lp__sdfrtp_lp2.pxi.spice"
*
.ends
*
*
