* File: sky130_fd_sc_lp__o41ai_1.pxi.spice
* Created: Wed Sep  2 10:28:11 2020
* 
x_PM_SKY130_FD_SC_LP__O41AI_1%B1 N_B1_M1004_g N_B1_M1005_g N_B1_c_62_n
+ N_B1_c_63_n B1 N_B1_c_64_n PM_SKY130_FD_SC_LP__O41AI_1%B1
x_PM_SKY130_FD_SC_LP__O41AI_1%A4 N_A4_M1003_g N_A4_M1008_g A4 N_A4_c_99_n
+ N_A4_c_100_n PM_SKY130_FD_SC_LP__O41AI_1%A4
x_PM_SKY130_FD_SC_LP__O41AI_1%A3 N_A3_M1009_g N_A3_M1006_g A3 A3 A3 A3
+ N_A3_c_137_n N_A3_c_140_n PM_SKY130_FD_SC_LP__O41AI_1%A3
x_PM_SKY130_FD_SC_LP__O41AI_1%A2 N_A2_M1000_g N_A2_M1002_g A2 A2 A2 A2
+ N_A2_c_171_n N_A2_c_172_n PM_SKY130_FD_SC_LP__O41AI_1%A2
x_PM_SKY130_FD_SC_LP__O41AI_1%A1 N_A1_M1007_g N_A1_c_212_n N_A1_M1001_g A1 A1
+ N_A1_c_214_n PM_SKY130_FD_SC_LP__O41AI_1%A1
x_PM_SKY130_FD_SC_LP__O41AI_1%VPWR N_VPWR_M1005_s N_VPWR_M1007_d N_VPWR_c_240_n
+ N_VPWR_c_241_n N_VPWR_c_242_n N_VPWR_c_243_n N_VPWR_c_244_n N_VPWR_c_245_n
+ N_VPWR_c_246_n N_VPWR_c_247_n N_VPWR_c_248_n VPWR N_VPWR_c_239_n
+ PM_SKY130_FD_SC_LP__O41AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O41AI_1%Y N_Y_M1004_s N_Y_M1005_d N_Y_c_284_n N_Y_c_285_n
+ N_Y_c_295_n N_Y_c_286_n N_Y_c_299_n N_Y_c_287_n Y Y
+ PM_SKY130_FD_SC_LP__O41AI_1%Y
x_PM_SKY130_FD_SC_LP__O41AI_1%A_156_49# N_A_156_49#_M1004_d N_A_156_49#_M1006_d
+ N_A_156_49#_M1001_d N_A_156_49#_c_366_p N_A_156_49#_c_335_n
+ N_A_156_49#_c_330_n N_A_156_49#_c_331_n N_A_156_49#_c_347_n
+ N_A_156_49#_c_332_n N_A_156_49#_c_333_n N_A_156_49#_c_361_n
+ N_A_156_49#_c_334_n PM_SKY130_FD_SC_LP__O41AI_1%A_156_49#
x_PM_SKY130_FD_SC_LP__O41AI_1%VGND N_VGND_M1003_d N_VGND_M1000_d N_VGND_c_375_n
+ N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n
+ VGND N_VGND_c_381_n N_VGND_c_382_n PM_SKY130_FD_SC_LP__O41AI_1%VGND
cc_1 VNB N_B1_M1004_g 0.0265875f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_2 VNB N_B1_M1005_g 0.00140588f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_3 VNB N_B1_c_62_n 0.0631146f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_4 VNB N_B1_c_63_n 0.00892181f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.46
cc_5 VNB N_B1_c_64_n 0.00133231f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_6 VNB N_A4_M1003_g 0.0251639f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_7 VNB N_A4_c_99_n 0.0238903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A4_c_100_n 0.00349935f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_9 VNB N_A3_M1006_g 0.0242505f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_10 VNB N_A3_c_137_n 0.0256238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_M1000_g 0.0258652f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_12 VNB N_A2_c_171_n 0.0240668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_172_n 0.0018225f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_14 VNB N_A1_M1007_g 0.00617342f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_15 VNB N_A1_c_212_n 0.0241591f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.625
cc_16 VNB A1 0.0270004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_214_n 0.056972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_239_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_284_n 0.0559865f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_20 VNB N_Y_c_285_n 0.00512794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_286_n 0.00312589f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_22 VNB N_Y_c_287_n 0.0011565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_156_49#_c_330_n 0.00727168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_156_49#_c_331_n 0.00293128f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_25 VNB N_A_156_49#_c_332_n 0.016709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_156_49#_c_333_n 0.0240525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_156_49#_c_334_n 0.00776206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_375_n 6.31895e-19 $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_29 VNB N_VGND_c_376_n 0.00527698f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_30 VNB N_VGND_c_377_n 0.0343089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_378_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_32 VNB N_VGND_c_379_n 0.0159489f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_33 VNB N_VGND_c_380_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_381_n 0.0235955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_382_n 0.197622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B1_M1005_g 0.0247258f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.465
cc_37 VPB N_B1_c_64_n 0.0125667f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_38 VPB N_A4_M1008_g 0.0184253f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.465
cc_39 VPB N_A4_c_99_n 0.00604703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A4_c_100_n 0.00403622f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_41 VPB N_A3_M1009_g 0.0187087f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.665
cc_42 VPB N_A3_c_137_n 0.00647694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A3_c_140_n 9.91125e-19 $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.665
cc_44 VPB N_A2_M1002_g 0.0197733f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.465
cc_45 VPB N_A2_c_171_n 0.00635559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A2_c_172_n 0.00280287f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.665
cc_47 VPB N_A1_M1007_g 0.0256895f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.665
cc_48 VPB A1 0.0146462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_240_n 0.0157682f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.46
cc_50 VPB N_VPWR_c_241_n 0.024835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_242_n 0.0487765f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_52 VPB N_VPWR_c_243_n 0.00756884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_244_n 0.0120081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_245_n 0.00592961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_246_n 0.0115308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_247_n 0.053391f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_248_n 0.00564109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_239_n 0.0612855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_Y_c_287_n 0.00134343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_B1_M1004_g N_A4_M1003_g 0.0159512f $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_61 N_B1_M1005_g N_A4_M1008_g 0.0248894f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_62 N_B1_c_63_n N_A4_c_99_n 0.0204739f $X=0.705 $Y=1.46 $X2=0 $Y2=0
cc_63 N_B1_M1005_g N_A4_c_100_n 2.95813e-19 $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_64 N_B1_c_63_n N_A4_c_100_n 2.84307e-19 $X=0.705 $Y=1.46 $X2=0 $Y2=0
cc_65 N_B1_M1005_g N_VPWR_c_240_n 0.00203034f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_66 N_B1_c_62_n N_VPWR_c_240_n 0.00489383f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_67 N_B1_c_64_n N_VPWR_c_240_n 0.0123768f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_68 N_B1_M1005_g N_VPWR_c_241_n 0.0156237f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_69 N_B1_M1005_g N_VPWR_c_243_n 0.00576034f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_70 N_B1_M1005_g N_VPWR_c_247_n 0.00329941f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_71 N_B1_M1005_g N_VPWR_c_239_n 0.00621015f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_72 N_B1_M1004_g N_Y_c_284_n 0.0232088f $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_73 N_B1_c_62_n N_Y_c_284_n 0.016623f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_74 N_B1_c_64_n N_Y_c_284_n 0.026848f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_75 N_B1_M1004_g N_Y_c_285_n 0.00327281f $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_76 N_B1_c_62_n N_Y_c_285_n 0.0020886f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_77 N_B1_c_63_n N_Y_c_285_n 0.00145124f $X=0.705 $Y=1.46 $X2=0 $Y2=0
cc_78 N_B1_M1005_g N_Y_c_295_n 0.0078023f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_79 N_B1_c_62_n N_Y_c_286_n 0.00328001f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_80 N_B1_c_63_n N_Y_c_286_n 0.0082896f $X=0.705 $Y=1.46 $X2=0 $Y2=0
cc_81 N_B1_c_64_n N_Y_c_286_n 0.0103421f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_82 N_B1_M1005_g N_Y_c_299_n 0.00833149f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_83 N_B1_M1005_g N_Y_c_287_n 0.0122852f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_84 N_B1_c_63_n N_Y_c_287_n 0.00314786f $X=0.705 $Y=1.46 $X2=0 $Y2=0
cc_85 N_B1_c_64_n N_Y_c_287_n 0.0119309f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_86 N_B1_M1004_g N_A_156_49#_c_335_n 8.68324e-19 $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_87 N_B1_M1004_g N_A_156_49#_c_331_n 8.15239e-19 $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_88 N_B1_M1004_g N_VGND_c_375_n 9.86076e-19 $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_89 N_B1_M1004_g N_VGND_c_377_n 0.00567689f $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_90 N_B1_M1004_g N_VGND_c_382_n 0.011931f $X=0.705 $Y=0.665 $X2=0 $Y2=0
cc_91 N_A4_M1008_g N_A3_M1009_g 0.055106f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A4_M1003_g N_A3_M1006_g 0.0227449f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_93 N_A4_c_99_n N_A3_c_137_n 0.055106f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_94 N_A4_c_100_n N_A3_c_137_n 0.0037331f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_95 N_A4_M1008_g N_A3_c_140_n 0.00415135f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A4_c_99_n N_A3_c_140_n 4.09673e-19 $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_97 N_A4_c_100_n N_A3_c_140_n 0.0277709f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_98 N_A4_M1008_g N_VPWR_c_243_n 0.00119488f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A4_M1008_g N_VPWR_c_247_n 0.00585385f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A4_M1008_g N_VPWR_c_239_n 0.0109726f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A4_M1003_g N_Y_c_284_n 9.39668e-19 $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_102 N_A4_M1003_g N_Y_c_285_n 0.00255463f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_103 N_A4_c_99_n N_Y_c_286_n 0.00109306f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A4_c_100_n N_Y_c_286_n 0.0130455f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A4_c_99_n N_Y_c_299_n 0.00365618f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_106 N_A4_c_100_n N_Y_c_299_n 0.00596726f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_107 N_A4_M1008_g N_Y_c_287_n 0.0014647f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A4_c_99_n N_Y_c_287_n 9.92202e-19 $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A4_c_100_n N_Y_c_287_n 0.020145f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_110 N_A4_M1003_g N_A_156_49#_c_330_n 0.014674f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_111 N_A4_c_99_n N_A_156_49#_c_330_n 2.43608e-19 $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_112 N_A4_c_100_n N_A_156_49#_c_330_n 0.0168491f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A4_c_99_n N_A_156_49#_c_331_n 0.00410629f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_114 N_A4_c_100_n N_A_156_49#_c_331_n 0.00552785f $X=1.155 $Y=1.51 $X2=0 $Y2=0
cc_115 N_A4_M1003_g N_VGND_c_375_n 0.00952815f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_116 N_A4_M1003_g N_VGND_c_377_n 0.00554242f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_117 N_A4_M1003_g N_VGND_c_382_n 0.0097429f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_118 N_A3_M1006_g N_A2_M1000_g 0.0217579f $X=1.685 $Y=0.665 $X2=0 $Y2=0
cc_119 N_A3_M1009_g N_A2_M1002_g 0.0463739f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A3_c_140_n N_A2_M1002_g 0.00448739f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_121 N_A3_c_137_n N_A2_c_171_n 0.0215729f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_122 N_A3_c_140_n N_A2_c_171_n 2.88395e-19 $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_123 N_A3_M1009_g N_A2_c_172_n 0.00121245f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A3_c_137_n N_A2_c_172_n 0.00142573f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A3_c_140_n N_A2_c_172_n 0.0786783f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_126 N_A3_M1009_g N_VPWR_c_247_n 0.00380992f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A3_c_140_n N_VPWR_c_247_n 0.0120634f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A3_M1009_g N_VPWR_c_239_n 0.00560506f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A3_c_140_n N_VPWR_c_239_n 0.0112808f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A3_c_140_n N_Y_c_287_n 0.00450668f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A3_c_140_n A_336_367# 0.011279f $X=1.695 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_132 N_A3_M1006_g N_A_156_49#_c_330_n 0.0139306f $X=1.685 $Y=0.665 $X2=0 $Y2=0
cc_133 N_A3_c_137_n N_A_156_49#_c_330_n 0.00324294f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A3_c_140_n N_A_156_49#_c_330_n 0.0157617f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A3_c_137_n N_A_156_49#_c_334_n 0.00137126f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_136 N_A3_c_140_n N_A_156_49#_c_334_n 0.00360051f $X=1.695 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A3_M1006_g N_VGND_c_375_n 0.0103237f $X=1.685 $Y=0.665 $X2=0 $Y2=0
cc_138 N_A3_M1006_g N_VGND_c_379_n 0.00477554f $X=1.685 $Y=0.665 $X2=0 $Y2=0
cc_139 N_A3_M1006_g N_VGND_c_382_n 0.0083544f $X=1.685 $Y=0.665 $X2=0 $Y2=0
cc_140 N_A2_M1002_g N_A1_M1007_g 0.0418446f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A2_c_172_n N_A1_M1007_g 0.0134457f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_142 N_A2_M1000_g N_A1_c_212_n 0.0269469f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_143 N_A2_M1000_g A1 4.73389e-19 $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_144 N_A2_c_171_n A1 5.72294e-19 $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A2_c_172_n A1 0.0113653f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_146 N_A2_M1000_g N_A1_c_214_n 0.00508057f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_147 N_A2_c_171_n N_A1_c_214_n 0.021735f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_148 N_A2_c_172_n N_A1_c_214_n 0.00102653f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A2_M1002_g N_VPWR_c_242_n 0.00254586f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A2_c_172_n N_VPWR_c_242_n 0.0538401f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A2_M1002_g N_VPWR_c_247_n 0.0037962f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A2_c_172_n N_VPWR_c_247_n 0.0129487f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_153 N_A2_M1002_g N_VPWR_c_239_n 0.00607065f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A2_c_172_n N_VPWR_c_239_n 0.0127399f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A2_c_172_n A_444_367# 0.013998f $X=2.235 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_156 N_A2_M1000_g N_A_156_49#_c_347_n 0.00907968f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_157 N_A2_M1000_g N_A_156_49#_c_332_n 0.017185f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_158 N_A2_c_171_n N_A_156_49#_c_332_n 0.00429673f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A2_c_172_n N_A_156_49#_c_332_n 0.0190054f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A2_M1000_g N_A_156_49#_c_333_n 6.22624e-19 $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_161 N_A2_M1000_g N_A_156_49#_c_334_n 0.00180647f $X=2.145 $Y=0.665 $X2=0
+ $Y2=0
cc_162 N_A2_c_172_n N_A_156_49#_c_334_n 0.00371555f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A2_M1000_g N_VGND_c_375_n 6.60715e-19 $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_164 N_A2_M1000_g N_VGND_c_376_n 0.0045014f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_165 N_A2_M1000_g N_VGND_c_379_n 0.00554241f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_166 N_A2_M1000_g N_VGND_c_382_n 0.0105709f $X=2.145 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A1_M1007_g N_VPWR_c_242_n 0.0330202f $X=2.685 $Y=2.465 $X2=0 $Y2=0
cc_168 A1 N_VPWR_c_242_n 0.0140416f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_169 N_A1_c_214_n N_VPWR_c_242_n 0.00490531f $X=2.99 $Y=1.375 $X2=0 $Y2=0
cc_170 N_A1_M1007_g N_VPWR_c_247_n 0.00329941f $X=2.685 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A1_M1007_g N_VPWR_c_239_n 0.00621015f $X=2.685 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A1_c_212_n N_A_156_49#_c_347_n 6.11959e-19 $X=2.705 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A1_c_212_n N_A_156_49#_c_332_n 0.0272608f $X=2.705 $Y=1.21 $X2=0 $Y2=0
cc_174 A1 N_A_156_49#_c_332_n 0.0154542f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A1_c_214_n N_A_156_49#_c_332_n 0.00665908f $X=2.99 $Y=1.375 $X2=0 $Y2=0
cc_176 N_A1_c_212_n N_A_156_49#_c_333_n 0.0114533f $X=2.705 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A1_c_212_n N_VGND_c_376_n 0.00577032f $X=2.705 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A1_c_212_n N_VGND_c_381_n 0.00539298f $X=2.705 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A1_c_212_n N_VGND_c_382_n 0.0111955f $X=2.705 $Y=1.21 $X2=0 $Y2=0
cc_180 N_VPWR_c_239_n N_Y_M1005_d 0.00635978f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_240_n N_Y_c_295_n 0.00857317f $X=0.475 $Y=2.09 $X2=0 $Y2=0
cc_182 N_VPWR_c_243_n N_Y_c_295_n 0.0572577f $X=0.49 $Y=2.505 $X2=0 $Y2=0
cc_183 N_VPWR_c_247_n N_Y_c_295_n 0.0191767f $X=2.695 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_239_n N_Y_c_295_n 0.0115856f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_c_240_n N_Y_c_287_n 0.0188506f $X=0.475 $Y=2.09 $X2=0 $Y2=0
cc_186 N_VPWR_c_239_n A_264_367# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_187 N_VPWR_c_239_n A_336_367# 0.00922383f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_188 N_VPWR_c_239_n A_444_367# 0.0106195f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_189 N_Y_c_284_n N_A_156_49#_c_335_n 0.0068948f $X=0.71 $Y=1.195 $X2=0 $Y2=0
cc_190 N_Y_c_284_n N_A_156_49#_c_331_n 0.0121466f $X=0.71 $Y=1.195 $X2=0 $Y2=0
cc_191 N_Y_c_286_n N_A_156_49#_c_361_n 0.00296877f $X=0.815 $Y=1.43 $X2=0 $Y2=0
cc_192 N_Y_c_284_n N_VGND_c_377_n 0.0370279f $X=0.71 $Y=1.195 $X2=0 $Y2=0
cc_193 N_Y_M1004_s N_VGND_c_382_n 0.00212301f $X=0.365 $Y=0.245 $X2=0 $Y2=0
cc_194 N_Y_c_284_n N_VGND_c_382_n 0.0212867f $X=0.71 $Y=1.195 $X2=0 $Y2=0
cc_195 N_A_156_49#_c_330_n N_VGND_M1003_d 0.00197722f $X=1.805 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_156_49#_c_332_n N_VGND_M1000_d 0.00379592f $X=2.583 $Y=1.022 $X2=0
+ $Y2=0
cc_197 N_A_156_49#_c_330_n N_VGND_c_375_n 0.0171814f $X=1.805 $Y=1.09 $X2=0
+ $Y2=0
cc_198 N_A_156_49#_c_332_n N_VGND_c_376_n 0.0250691f $X=2.583 $Y=1.022 $X2=0
+ $Y2=0
cc_199 N_A_156_49#_c_366_p N_VGND_c_377_n 0.020821f $X=0.97 $Y=0.4 $X2=0 $Y2=0
cc_200 N_A_156_49#_c_347_n N_VGND_c_379_n 0.0171157f $X=1.9 $Y=0.42 $X2=0 $Y2=0
cc_201 N_A_156_49#_c_333_n N_VGND_c_381_n 0.0210467f $X=2.92 $Y=0.39 $X2=0 $Y2=0
cc_202 N_A_156_49#_M1004_d N_VGND_c_382_n 0.00477913f $X=0.78 $Y=0.245 $X2=0
+ $Y2=0
cc_203 N_A_156_49#_M1006_d N_VGND_c_382_n 0.00404228f $X=1.76 $Y=0.245 $X2=0
+ $Y2=0
cc_204 N_A_156_49#_M1001_d N_VGND_c_382_n 0.00212301f $X=2.78 $Y=0.245 $X2=0
+ $Y2=0
cc_205 N_A_156_49#_c_366_p N_VGND_c_382_n 0.0127317f $X=0.97 $Y=0.4 $X2=0 $Y2=0
cc_206 N_A_156_49#_c_347_n N_VGND_c_382_n 0.0106708f $X=1.9 $Y=0.42 $X2=0 $Y2=0
cc_207 N_A_156_49#_c_333_n N_VGND_c_382_n 0.0125689f $X=2.92 $Y=0.39 $X2=0 $Y2=0
