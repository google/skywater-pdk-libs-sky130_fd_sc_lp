* File: sky130_fd_sc_lp__o311a_2.pex.spice
* Created: Wed Sep  2 10:23:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311A_2%A_85_21# 1 2 3 10 12 15 17 19 22 26 27 29 30
+ 31 33 35 38 41 45 49 52
r114 56 57 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.93 $Y=1.35
+ $X2=0.965 $Y2=1.35
r115 55 56 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=0.535 $Y=1.35
+ $X2=0.93 $Y2=1.35
r116 53 55 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.5 $Y=1.35
+ $X2=0.535 $Y2=1.35
r117 50 52 22.5665 $w=1.73e-07 $l=3.2e-07 $layer=LI1_cond $X=3.58 $Y=2.01
+ $X2=3.9 $Y2=2.01
r118 45 52 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=3.935 $Y=2.91
+ $X2=3.935 $Y2=2.1
r119 39 49 2.63236 $w=3.65e-07 $l=3.05e-07 $layer=LI1_cond $X=3.79 $Y=1.005
+ $X2=3.485 $Y2=1.005
r120 39 41 12.9575 $w=5.38e-07 $l=5.85e-07 $layer=LI1_cond $X=3.79 $Y=1.005
+ $X2=3.79 $Y2=0.42
r121 38 50 0.136533 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=3.58 $Y=1.92 $X2=3.58
+ $Y2=2.01
r122 37 49 2.63236 $w=3.65e-07 $l=2.1225e-07 $layer=LI1_cond $X=3.58 $Y=1.175
+ $X2=3.485 $Y2=1.005
r123 37 38 43.488 $w=1.88e-07 $l=7.45e-07 $layer=LI1_cond $X=3.58 $Y=1.175
+ $X2=3.58 $Y2=1.92
r124 36 48 3.99943 $w=1.8e-07 $l=1.2e-07 $layer=LI1_cond $X=3.135 $Y=2.01
+ $X2=3.015 $Y2=2.01
r125 35 50 6.43889 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.485 $Y=2.01
+ $X2=3.58 $Y2=2.01
r126 35 36 21.5657 $w=1.78e-07 $l=3.5e-07 $layer=LI1_cond $X=3.485 $Y=2.01
+ $X2=3.135 $Y2=2.01
r127 31 48 2.99957 $w=2.4e-07 $l=9e-08 $layer=LI1_cond $X=3.015 $Y=2.1 $X2=3.015
+ $Y2=2.01
r128 31 33 38.895 $w=2.38e-07 $l=8.1e-07 $layer=LI1_cond $X=3.015 $Y=2.1
+ $X2=3.015 $Y2=2.91
r129 29 49 4.19346 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=1.09
+ $X2=3.485 $Y2=1.005
r130 29 30 146.791 $w=1.68e-07 $l=2.25e-06 $layer=LI1_cond $X=3.485 $Y=1.09
+ $X2=1.235 $Y2=1.09
r131 27 57 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.07 $Y=1.35
+ $X2=0.965 $Y2=1.35
r132 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.35 $X2=1.07 $Y2=1.35
r133 24 30 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.107 $Y=1.175
+ $X2=1.235 $Y2=1.09
r134 24 26 7.90892 $w=2.53e-07 $l=1.75e-07 $layer=LI1_cond $X=1.107 $Y=1.175
+ $X2=1.107 $Y2=1.35
r135 20 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=1.35
r136 20 22 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=2.465
r137 17 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=1.35
r138 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=0.655
r139 13 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.515
+ $X2=0.535 $Y2=1.35
r140 13 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.535 $Y=1.515
+ $X2=0.535 $Y2=2.465
r141 10 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.185
+ $X2=0.5 $Y2=1.35
r142 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.5 $Y=1.185
+ $X2=0.5 $Y2=0.655
r143 3 52 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.76
+ $Y=1.835 $X2=3.9 $Y2=2.095
r144 3 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.76
+ $Y=1.835 $X2=3.9 $Y2=2.91
r145 2 48 400 $w=1.7e-07 $l=4.3229e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.835 $X2=3 $Y2=2.085
r146 2 33 400 $w=1.7e-07 $l=1.22678e-06 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.835 $X2=3 $Y2=2.91
r147 1 41 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.755
+ $Y=0.235 $X2=3.895 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%A1 3 7 9 10 11 12 19 36
r39 23 36 2.91812 $w=2.35e-07 $l=1.7e-07 $layer=LI1_cond $X=1.712 $Y=1.685
+ $X2=1.712 $Y2=1.515
r40 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.51
+ $X2=1.61 $Y2=1.675
r41 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.51
+ $X2=1.61 $Y2=1.345
r42 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.51 $X2=1.61 $Y2=1.51
r43 11 12 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.712 $Y=2.405
+ $X2=1.712 $Y2=2.775
r44 10 11 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.712 $Y=2.035
+ $X2=1.712 $Y2=2.405
r45 9 36 1.08465 $w=3.38e-07 $l=3.2e-08 $layer=LI1_cond $X=1.68 $Y=1.515
+ $X2=1.712 $Y2=1.515
r46 9 20 2.37268 $w=3.38e-07 $l=7e-08 $layer=LI1_cond $X=1.68 $Y=1.515 $X2=1.61
+ $Y2=1.515
r47 9 10 15.5948 $w=2.33e-07 $l=3.18e-07 $layer=LI1_cond $X=1.712 $Y=1.717
+ $X2=1.712 $Y2=2.035
r48 9 23 1.56928 $w=2.33e-07 $l=3.2e-08 $layer=LI1_cond $X=1.712 $Y=1.717
+ $X2=1.712 $Y2=1.685
r49 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.7 $Y=2.465 $X2=1.7
+ $Y2=1.675
r50 3 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.7 $Y=0.655 $X2=1.7
+ $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%A2 1 3 7 9 10 11 12 19
r35 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.51 $X2=2.15 $Y2=1.51
r36 11 12 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.152 $Y=2.405
+ $X2=2.152 $Y2=2.775
r37 10 11 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.152 $Y=2.035
+ $X2=2.152 $Y2=2.405
r38 9 10 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.152 $Y=1.665
+ $X2=2.152 $Y2=2.035
r39 9 19 5.85668 $w=3.03e-07 $l=1.55e-07 $layer=LI1_cond $X=2.152 $Y=1.665
+ $X2=2.152 $Y2=1.51
r40 5 18 42.2564 $w=3.29e-07 $l=2.28583e-07 $layer=POLY_cond $X=2.235 $Y=1.32
+ $X2=2.15 $Y2=1.51
r41 5 7 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.235 $Y=1.32
+ $X2=2.235 $Y2=0.655
r42 1 18 38.5938 $w=3.29e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.06 $Y=1.675
+ $X2=2.15 $Y2=1.51
r43 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.06 $Y=1.675 $X2=2.06
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%A3 3 7 9 10 11 12 19 20 36
c38 20 0 1.54763e-19 $X=2.69 $Y=1.51
r39 36 37 3.17508 $w=3.33e-07 $l=7e-08 $layer=LI1_cond $X=2.642 $Y=1.665
+ $X2=2.642 $Y2=1.735
r40 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.51
+ $X2=2.69 $Y2=1.675
r41 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.51
+ $X2=2.69 $Y2=1.345
r42 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.51 $X2=2.69 $Y2=1.51
r43 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.6 $Y=2.405 $X2=2.6
+ $Y2=2.775
r44 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.6 $Y=2.035 $X2=2.6
+ $Y2=2.405
r45 9 36 0.27521 $w=3.33e-07 $l=8e-09 $layer=LI1_cond $X=2.642 $Y=1.657
+ $X2=2.642 $Y2=1.665
r46 9 20 5.05699 $w=3.33e-07 $l=1.47e-07 $layer=LI1_cond $X=2.642 $Y=1.657
+ $X2=2.642 $Y2=1.51
r47 9 10 13.5066 $w=2.48e-07 $l=2.93e-07 $layer=LI1_cond $X=2.6 $Y=1.742 $X2=2.6
+ $Y2=2.035
r48 9 37 0.322684 $w=2.48e-07 $l=7e-09 $layer=LI1_cond $X=2.6 $Y=1.742 $X2=2.6
+ $Y2=1.735
r49 7 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.78 $Y=0.655
+ $X2=2.78 $Y2=1.345
r50 3 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.6 $Y=2.465 $X2=2.6
+ $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%B1 3 7 9 12 13
c36 3 0 1.54763e-19 $X=3.255 $Y=2.465
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.51
+ $X2=3.23 $Y2=1.675
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.51
+ $X2=3.23 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.23
+ $Y=1.51 $X2=3.23 $Y2=1.51
r40 9 13 5.3322 $w=3.33e-07 $l=1.55e-07 $layer=LI1_cond $X=3.147 $Y=1.665
+ $X2=3.147 $Y2=1.51
r41 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.32 $Y=0.655
+ $X2=3.32 $Y2=1.345
r42 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.255 $Y=2.465
+ $X2=3.255 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%C1 3 7 10 11 14 15
r27 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.46 $X2=4.01 $Y2=1.46
r28 11 15 6.05771 $w=3.88e-07 $l=2.05e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=1.46
r29 9 14 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.76 $Y=1.46 $X2=4.01
+ $Y2=1.46
r30 9 10 5.03009 $w=3.3e-07 $l=2.29783e-07 $layer=POLY_cond $X=3.76 $Y=1.46
+ $X2=3.605 $Y2=1.295
r31 5 10 37.0704 $w=1.5e-07 $l=3.67831e-07 $layer=POLY_cond $X=3.685 $Y=1.625
+ $X2=3.605 $Y2=1.295
r32 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.685 $Y=1.625
+ $X2=3.685 $Y2=2.465
r33 1 10 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.68 $Y=1.295
+ $X2=3.605 $Y2=1.295
r34 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.68 $Y=1.295 $X2=3.68
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%VPWR 1 2 3 10 12 16 20 26 29 30 31 41 42 48
r57 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 36 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 35 38 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r65 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 33 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.29 $Y2=3.33
r67 33 35 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 31 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 31 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 29 38 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=3.12 $Y2=3.33
r71 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=3.47 $Y2=3.33
r72 28 41 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.635 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=3.33
+ $X2=3.47 $Y2=3.33
r74 24 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=3.245
+ $X2=3.47 $Y2=3.33
r75 24 26 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.47 $Y=3.245
+ $X2=3.47 $Y2=2.375
r76 20 23 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.29 $Y=2.02
+ $X2=1.29 $Y2=2.95
r77 18 48 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=3.245
+ $X2=1.29 $Y2=3.33
r78 18 23 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.29 $Y=3.245
+ $X2=1.29 $Y2=2.95
r79 17 45 4.1267 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r80 16 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.29 $Y2=3.33
r81 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.425 $Y2=3.33
r82 12 15 41.4026 $w=2.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.29 $Y=1.98
+ $X2=0.29 $Y2=2.95
r83 10 45 3.15799 $w=2.7e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.212 $Y2=3.33
r84 10 15 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.95
r85 3 26 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=3.33
+ $Y=1.835 $X2=3.47 $Y2=2.375
r86 2 23 400 $w=1.7e-07 $l=1.24717e-06 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.835 $X2=1.32 $Y2=2.95
r87 2 20 400 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.835 $X2=1.32 $Y2=2.02
r88 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.32 $Y2=2.95
r89 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.32 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%X 1 2 7 8 9 10 11 12 13 24 34
r24 34 47 1.60806 $w=2.13e-07 $l=3e-08 $layer=LI1_cond $X=0.702 $Y=1.665
+ $X2=0.702 $Y2=1.695
r25 13 44 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=0.755 $Y=2.775
+ $X2=0.755 $Y2=2.91
r26 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=2.405
+ $X2=0.755 $Y2=2.775
r27 11 12 15.3059 $w=3.18e-07 $l=4.25e-07 $layer=LI1_cond $X=0.755 $Y=1.98
+ $X2=0.755 $Y2=2.405
r28 11 35 4.50173 $w=3.18e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=1.98
+ $X2=0.755 $Y2=1.855
r29 10 35 4.78984 $w=3.18e-07 $l=1.33e-07 $layer=LI1_cond $X=0.755 $Y=1.722
+ $X2=0.755 $Y2=1.855
r30 10 47 2.21774 $w=3.18e-07 $l=2.7e-08 $layer=LI1_cond $X=0.755 $Y=1.722
+ $X2=0.755 $Y2=1.695
r31 10 34 1.50086 $w=2.13e-07 $l=2.8e-08 $layer=LI1_cond $X=0.702 $Y=1.637
+ $X2=0.702 $Y2=1.665
r32 9 10 18.3319 $w=2.13e-07 $l=3.42e-07 $layer=LI1_cond $X=0.702 $Y=1.295
+ $X2=0.702 $Y2=1.637
r33 8 9 19.8327 $w=2.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.702 $Y=0.925
+ $X2=0.702 $Y2=1.295
r34 7 8 19.8327 $w=2.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.702 $Y=0.555
+ $X2=0.702 $Y2=0.925
r35 7 24 7.23627 $w=2.13e-07 $l=1.35e-07 $layer=LI1_cond $X=0.702 $Y=0.555
+ $X2=0.702 $Y2=0.42
r36 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.835 $X2=0.75 $Y2=2.91
r37 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.835 $X2=0.75 $Y2=1.98
r38 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r56 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r57 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r58 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 37 47 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=2.64
+ $Y2=0
r60 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.51
+ $Y2=0
r62 34 36 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.675 $Y=0
+ $X2=4.08 $Y2=0
r63 30 43 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.315
+ $Y2=0
r64 30 32 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=2.16
+ $Y2=0
r65 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.51
+ $Y2=0
r66 29 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.16
+ $Y2=0
r67 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r68 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r69 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r70 25 40 4.49694 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r71 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r72 24 43 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.315
+ $Y2=0
r73 24 27 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.72
+ $Y2=0
r74 22 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r75 22 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r76 22 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r77 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0
r78 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0.37
r79 14 43 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=0.085
+ $X2=1.315 $Y2=0
r80 14 16 4.90928 $w=6.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.315 $Y=0.085
+ $X2=1.315 $Y2=0.36
r81 10 40 3.0613 $w=3.05e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.272 $Y=0.085
+ $X2=0.212 $Y2=0
r82 10 12 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.272 $Y=0.085
+ $X2=0.272 $Y2=0.38
r83 3 20 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.235 $X2=2.51 $Y2=0.37
r84 2 16 45.5 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=4 $X=1.005
+ $Y=0.235 $X2=1.485 $Y2=0.36
r85 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_2%A_355_47# 1 2 7 9 11 13 15
r18 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=0.665 $X2=3.05
+ $Y2=0.75
r19 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.05 $Y=0.665
+ $X2=3.05 $Y2=0.37
r20 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=0.75
+ $X2=1.985 $Y2=0.75
r21 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=0.75
+ $X2=3.05 $Y2=0.75
r22 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.885 $Y=0.75
+ $X2=2.15 $Y2=0.75
r23 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.665
+ $X2=1.985 $Y2=0.75
r24 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.985 $Y=0.665
+ $X2=1.985 $Y2=0.37
r25 2 20 182 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.235 $X2=3.05 $Y2=0.75
r26 2 15 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.235 $X2=3.05 $Y2=0.37
r27 1 18 182 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.235 $X2=1.985 $Y2=0.75
r28 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.235 $X2=1.985 $Y2=0.37
.ends

