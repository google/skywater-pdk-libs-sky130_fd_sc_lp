* File: sky130_fd_sc_lp__dlrtn_1.pxi.spice
* Created: Fri Aug 28 10:26:27 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTN_1%D N_D_M1018_g N_D_c_129_n N_D_M1008_g N_D_c_131_n
+ D D D D N_D_c_133_n N_D_c_134_n PM_SKY130_FD_SC_LP__DLRTN_1%D
x_PM_SKY130_FD_SC_LP__DLRTN_1%GATE_N N_GATE_N_c_167_n N_GATE_N_c_172_n
+ N_GATE_N_M1011_g N_GATE_N_c_168_n N_GATE_N_M1002_g N_GATE_N_c_169_n GATE_N
+ GATE_N GATE_N PM_SKY130_FD_SC_LP__DLRTN_1%GATE_N
x_PM_SKY130_FD_SC_LP__DLRTN_1%A_47_47# N_A_47_47#_M1018_s N_A_47_47#_M1008_s
+ N_A_47_47#_M1012_g N_A_47_47#_M1004_g N_A_47_47#_c_212_n N_A_47_47#_c_216_n
+ N_A_47_47#_c_217_n N_A_47_47#_c_230_n N_A_47_47#_c_218_n N_A_47_47#_c_219_n
+ N_A_47_47#_c_220_n N_A_47_47#_c_239_p N_A_47_47#_c_221_n N_A_47_47#_c_222_n
+ N_A_47_47#_c_213_n N_A_47_47#_c_224_n PM_SKY130_FD_SC_LP__DLRTN_1%A_47_47#
x_PM_SKY130_FD_SC_LP__DLRTN_1%A_387_385# N_A_387_385#_M1009_s
+ N_A_387_385#_M1001_s N_A_387_385#_M1003_g N_A_387_385#_M1006_g
+ N_A_387_385#_c_308_n N_A_387_385#_c_318_n N_A_387_385#_c_309_n
+ N_A_387_385#_c_310_n N_A_387_385#_c_311_n N_A_387_385#_c_312_n
+ N_A_387_385#_c_313_n N_A_387_385#_c_314_n N_A_387_385#_c_315_n
+ N_A_387_385#_c_320_n N_A_387_385#_c_343_p N_A_387_385#_c_316_n
+ PM_SKY130_FD_SC_LP__DLRTN_1%A_387_385#
x_PM_SKY130_FD_SC_LP__DLRTN_1%A_270_465# N_A_270_465#_M1002_d
+ N_A_270_465#_M1011_d N_A_270_465#_c_407_n N_A_270_465#_c_408_n
+ N_A_270_465#_c_409_n N_A_270_465#_c_410_n N_A_270_465#_M1009_g
+ N_A_270_465#_M1001_g N_A_270_465#_c_411_n N_A_270_465#_M1015_g
+ N_A_270_465#_c_413_n N_A_270_465#_M1016_g N_A_270_465#_c_415_n
+ N_A_270_465#_c_416_n N_A_270_465#_c_421_n N_A_270_465#_c_417_n
+ PM_SKY130_FD_SC_LP__DLRTN_1%A_270_465#
x_PM_SKY130_FD_SC_LP__DLRTN_1%A_820_99# N_A_820_99#_M1013_s N_A_820_99#_M1000_d
+ N_A_820_99#_M1019_g N_A_820_99#_M1014_g N_A_820_99#_M1010_g
+ N_A_820_99#_M1017_g N_A_820_99#_c_512_n N_A_820_99#_c_522_n
+ N_A_820_99#_c_523_n N_A_820_99#_c_513_n N_A_820_99#_c_536_p
+ N_A_820_99#_c_566_p N_A_820_99#_c_514_n N_A_820_99#_c_515_n
+ N_A_820_99#_c_516_n N_A_820_99#_c_517_n N_A_820_99#_c_518_n
+ N_A_820_99#_c_527_n N_A_820_99#_c_540_p PM_SKY130_FD_SC_LP__DLRTN_1%A_820_99#
x_PM_SKY130_FD_SC_LP__DLRTN_1%A_670_125# N_A_670_125#_M1015_d
+ N_A_670_125#_M1003_d N_A_670_125#_M1000_g N_A_670_125#_c_626_n
+ N_A_670_125#_M1013_g N_A_670_125#_c_635_n N_A_670_125#_c_645_n
+ N_A_670_125#_c_627_n N_A_670_125#_c_628_n N_A_670_125#_c_633_n
+ N_A_670_125#_c_629_n N_A_670_125#_c_630_n N_A_670_125#_c_631_n
+ PM_SKY130_FD_SC_LP__DLRTN_1%A_670_125#
x_PM_SKY130_FD_SC_LP__DLRTN_1%RESET_B N_RESET_B_M1005_g N_RESET_B_M1007_g
+ RESET_B RESET_B RESET_B RESET_B N_RESET_B_c_718_n N_RESET_B_c_719_n
+ PM_SKY130_FD_SC_LP__DLRTN_1%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTN_1%VPWR N_VPWR_M1008_d N_VPWR_M1001_d N_VPWR_M1014_d
+ N_VPWR_M1007_d N_VPWR_c_759_n N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_762_n
+ N_VPWR_c_763_n N_VPWR_c_764_n N_VPWR_c_765_n VPWR N_VPWR_c_766_n
+ N_VPWR_c_767_n N_VPWR_c_768_n N_VPWR_c_758_n N_VPWR_c_770_n N_VPWR_c_771_n
+ N_VPWR_c_772_n PM_SKY130_FD_SC_LP__DLRTN_1%VPWR
x_PM_SKY130_FD_SC_LP__DLRTN_1%Q N_Q_M1010_d N_Q_M1017_d N_Q_c_845_n Q Q Q Q Q Q
+ N_Q_c_844_n PM_SKY130_FD_SC_LP__DLRTN_1%Q
x_PM_SKY130_FD_SC_LP__DLRTN_1%VGND N_VGND_M1018_d N_VGND_M1009_d N_VGND_M1019_d
+ N_VGND_M1005_d N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n
+ N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n VGND
+ N_VGND_c_878_n N_VGND_c_879_n N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n
+ N_VGND_c_883_n PM_SKY130_FD_SC_LP__DLRTN_1%VGND
cc_1 VNB N_D_c_129_n 0.0234373f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.248
cc_2 VNB N_D_M1008_g 0.0122079f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.645
cc_3 VNB N_D_c_131_n 0.0229354f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.435
cc_4 VNB D 0.00269226f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_D_c_133_n 0.0218461f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.93
cc_6 VNB N_D_c_134_n 0.0208505f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.765
cc_7 VNB N_GATE_N_c_167_n 0.0313622f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.445
cc_8 VNB N_GATE_N_c_168_n 0.019891f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.435
cc_9 VNB N_GATE_N_c_169_n 0.0175544f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_10 VNB GATE_N 0.010837f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_A_47_47#_M1012_g 0.0233204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_47_47#_c_212_n 0.0649261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_47_47#_c_213_n 0.0258868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_387_385#_c_308_n 0.00152832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_387_385#_c_309_n 0.015342f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.765
cc_16 VNB N_A_387_385#_c_310_n 0.00205317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_387_385#_c_311_n 0.00244775f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.925
cc_18 VNB N_A_387_385#_c_312_n 0.00747861f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_19 VNB N_A_387_385#_c_313_n 0.040823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_387_385#_c_314_n 0.0107628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_387_385#_c_315_n 0.00471887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_387_385#_c_316_n 0.013342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_270_465#_c_407_n 0.0507294f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.645
cc_24 VNB N_A_270_465#_c_408_n 0.100933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_270_465#_c_409_n 0.0104045f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.435
cc_26 VNB N_A_270_465#_c_410_n 0.0157988f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_27 VNB N_A_270_465#_c_411_n 0.0191698f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.93
cc_28 VNB N_A_270_465#_M1015_g 0.0245497f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.93
cc_29 VNB N_A_270_465#_c_413_n 0.0317407f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.765
cc_30 VNB N_A_270_465#_M1016_g 0.00723459f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.925
cc_31 VNB N_A_270_465#_c_415_n 0.00968786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_270_465#_c_416_n 0.00504028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_270_465#_c_417_n 0.0884684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_820_99#_M1019_g 0.0361883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_820_99#_M1010_g 0.0297018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_820_99#_c_512_n 0.00672907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_820_99#_c_513_n 0.00345932f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_38 VNB N_A_820_99#_c_514_n 0.00107129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_820_99#_c_515_n 0.0290307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_820_99#_c_516_n 0.00168047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_820_99#_c_517_n 0.0170945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_820_99#_c_518_n 0.00589895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_670_125#_M1000_g 0.00791515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_670_125#_c_626_n 0.0181934f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_45 VNB N_A_670_125#_c_627_n 0.0314809f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.765
cc_46 VNB N_A_670_125#_c_628_n 0.00231246f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.925
cc_47 VNB N_A_670_125#_c_629_n 0.00342886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_670_125#_c_630_n 0.00117957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_670_125#_c_631_n 0.0507061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_M1007_g 0.00724144f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.435
cc_51 VNB RESET_B 0.0019867f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.645
cc_52 VNB N_RESET_B_c_718_n 0.0332538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_RESET_B_c_719_n 0.0162467f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.93
cc_54 VNB N_VPWR_c_758_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB Q 0.0187234f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_56 VNB Q 0.0299703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Q_c_844_n 0.0295031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_870_n 0.00501021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_871_n 0.0091586f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.93
cc_60 VNB N_VGND_c_872_n 0.0166246f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.555
cc_61 VNB N_VGND_c_873_n 0.0055721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_874_n 0.0362891f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_63 VNB N_VGND_c_875_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_876_n 0.0287045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_877_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_878_n 0.0298668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_879_n 0.0334976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_880_n 0.0223734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_881_n 0.358235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_882_n 0.00420608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_883_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_D_M1008_g 0.053648f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.645
cc_73 VPB D 0.00359562f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_74 VPB N_GATE_N_c_167_n 8.49495e-19 $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.445
cc_75 VPB N_GATE_N_c_172_n 0.0805383f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.445
cc_76 VPB GATE_N 0.00470789f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_77 VPB N_A_47_47#_M1004_g 0.0382299f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_78 VPB N_A_47_47#_c_212_n 0.0264057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_47_47#_c_216_n 0.0267258f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.93
cc_80 VPB N_A_47_47#_c_217_n 0.007554f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.555
cc_81 VPB N_A_47_47#_c_218_n 0.0159931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_47_47#_c_219_n 0.00128839f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.295
cc_83 VPB N_A_47_47#_c_220_n 0.00373348f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_84 VPB N_A_47_47#_c_221_n 0.00239166f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_47_47#_c_222_n 0.00481838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_47_47#_c_213_n 0.00741181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_47_47#_c_224_n 0.00805403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_387_385#_M1003_g 0.0229307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_387_385#_c_318_n 0.00576894f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.93
cc_90 VPB N_A_387_385#_c_315_n 0.00219115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_387_385#_c_320_n 0.0313812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_270_465#_M1001_g 0.0227417f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_270_465#_M1016_g 0.0383862f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.925
cc_94 VPB N_A_270_465#_c_415_n 0.0109429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_270_465#_c_421_n 0.00685209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_270_465#_c_417_n 0.0720361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_820_99#_M1014_g 0.0210687f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_98 VPB N_A_820_99#_M1017_g 0.024492f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.93
cc_99 VPB N_A_820_99#_c_512_n 0.0190866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_820_99#_c_522_n 0.0182854f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.925
cc_101 VPB N_A_820_99#_c_523_n 0.00968538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_820_99#_c_514_n 0.00147968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_820_99#_c_515_n 0.00859372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_820_99#_c_516_n 0.00318324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_820_99#_c_527_n 9.14999e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_670_125#_M1000_g 0.0226007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_670_125#_c_633_n 0.00598245f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_108 VPB N_A_670_125#_c_629_n 0.00427426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_RESET_B_M1007_g 0.0206274f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.435
cc_110 VPB RESET_B 0.00119034f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.645
cc_111 VPB N_VPWR_c_759_n 0.00850036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_760_n 0.0168777f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.93
cc_113 VPB N_VPWR_c_761_n 0.00292979f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.555
cc_114 VPB N_VPWR_c_762_n 0.0238595f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.925
cc_115 VPB N_VPWR_c_763_n 0.00505807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_764_n 0.0180046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_765_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_766_n 0.0432895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_767_n 0.0435739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_768_n 0.0237917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_758_n 0.108197f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_770_n 0.0258405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_771_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_772_n 0.0118963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_Q_c_845_n 0.0196162f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.435
cc_126 VPB Q 0.053005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 N_D_c_129_n N_GATE_N_c_167_n 0.0209066f $X=0.687 $Y=1.248 $X2=0 $Y2=0
cc_128 N_D_M1008_g N_GATE_N_c_167_n 0.00580494f $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_129 D N_GATE_N_c_167_n 6.82779e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_130 N_D_M1008_g N_GATE_N_c_172_n 0.0324702f $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_131 D N_GATE_N_c_172_n 0.00229783f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_132 D N_GATE_N_c_168_n 0.00286746f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_133 N_D_c_134_n N_GATE_N_c_168_n 0.00787502f $X=0.687 $Y=0.765 $X2=0 $Y2=0
cc_134 D N_GATE_N_c_169_n 8.14617e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_135 N_D_c_133_n N_GATE_N_c_169_n 0.0209066f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_136 N_D_M1008_g GATE_N 9.26449e-19 $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_137 D GATE_N 0.0926576f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_138 N_D_c_133_n GATE_N 0.00410908f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_139 D N_A_47_47#_c_212_n 0.110193f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_140 N_D_c_134_n N_A_47_47#_c_212_n 0.0402948f $X=0.687 $Y=0.765 $X2=0 $Y2=0
cc_141 N_D_M1008_g N_A_47_47#_c_216_n 4.69023e-19 $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_142 N_D_M1008_g N_A_47_47#_c_217_n 0.0208687f $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_143 D N_A_47_47#_c_217_n 0.0156797f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_144 N_D_M1008_g N_A_47_47#_c_230_n 0.00166975f $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_145 N_D_M1008_g N_VPWR_c_759_n 0.00404132f $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_146 N_D_M1008_g N_VPWR_c_758_n 0.00927489f $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_147 N_D_M1008_g N_VPWR_c_770_n 0.00465548f $X=0.575 $Y=2.645 $X2=0 $Y2=0
cc_148 D N_VGND_M1018_d 0.00417427f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_149 D N_VGND_c_870_n 0.0171752f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_150 N_D_c_134_n N_VGND_c_870_n 0.00432284f $X=0.687 $Y=0.765 $X2=0 $Y2=0
cc_151 D N_VGND_c_878_n 0.00631205f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_152 N_D_c_133_n N_VGND_c_878_n 0.00159997f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_153 N_D_c_134_n N_VGND_c_878_n 0.00552764f $X=0.687 $Y=0.765 $X2=0 $Y2=0
cc_154 D N_VGND_c_881_n 0.00672091f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_155 N_D_c_133_n N_VGND_c_881_n 0.00161114f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_156 N_D_c_134_n N_VGND_c_881_n 0.0117986f $X=0.687 $Y=0.765 $X2=0 $Y2=0
cc_157 N_GATE_N_c_172_n N_A_47_47#_c_217_n 0.014528f $X=1.275 $Y=2.215 $X2=0
+ $Y2=0
cc_158 GATE_N N_A_47_47#_c_217_n 0.0207563f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_159 N_GATE_N_c_172_n N_A_47_47#_c_230_n 0.0128978f $X=1.275 $Y=2.215 $X2=0
+ $Y2=0
cc_160 N_GATE_N_c_172_n N_A_47_47#_c_218_n 0.0119547f $X=1.275 $Y=2.215 $X2=0
+ $Y2=0
cc_161 N_GATE_N_c_172_n N_A_47_47#_c_219_n 0.00292372f $X=1.275 $Y=2.215 $X2=0
+ $Y2=0
cc_162 N_GATE_N_c_172_n N_A_47_47#_c_220_n 0.00258806f $X=1.275 $Y=2.215 $X2=0
+ $Y2=0
cc_163 N_GATE_N_c_167_n N_A_270_465#_c_407_n 0.00348267f $X=1.16 $Y=1.675 $X2=0
+ $Y2=0
cc_164 N_GATE_N_c_169_n N_A_270_465#_c_407_n 0.00701624f $X=1.285 $Y=0.84 $X2=0
+ $Y2=0
cc_165 N_GATE_N_c_168_n N_A_270_465#_c_409_n 0.00701624f $X=1.285 $Y=0.765 $X2=0
+ $Y2=0
cc_166 N_GATE_N_c_167_n N_A_270_465#_c_415_n 0.00141936f $X=1.16 $Y=1.675 $X2=0
+ $Y2=0
cc_167 N_GATE_N_c_172_n N_A_270_465#_c_415_n 0.00995905f $X=1.275 $Y=2.215 $X2=0
+ $Y2=0
cc_168 N_GATE_N_c_168_n N_A_270_465#_c_415_n 0.00495694f $X=1.285 $Y=0.765 $X2=0
+ $Y2=0
cc_169 GATE_N N_A_270_465#_c_415_n 0.0941572f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_170 N_GATE_N_c_172_n N_A_270_465#_c_421_n 4.42944e-19 $X=1.275 $Y=2.215 $X2=0
+ $Y2=0
cc_171 N_GATE_N_c_167_n N_A_270_465#_c_417_n 0.043922f $X=1.16 $Y=1.675 $X2=0
+ $Y2=0
cc_172 GATE_N N_A_270_465#_c_417_n 0.00463206f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_173 N_GATE_N_c_172_n N_VPWR_c_759_n 0.00353178f $X=1.275 $Y=2.215 $X2=0 $Y2=0
cc_174 N_GATE_N_c_172_n N_VPWR_c_766_n 0.00293691f $X=1.275 $Y=2.215 $X2=0 $Y2=0
cc_175 N_GATE_N_c_172_n N_VPWR_c_758_n 0.00381813f $X=1.275 $Y=2.215 $X2=0 $Y2=0
cc_176 N_GATE_N_c_168_n N_VGND_c_870_n 0.00356344f $X=1.285 $Y=0.765 $X2=0 $Y2=0
cc_177 N_GATE_N_c_169_n N_VGND_c_870_n 0.00314676f $X=1.285 $Y=0.84 $X2=0 $Y2=0
cc_178 GATE_N N_VGND_c_870_n 0.0148129f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_179 N_GATE_N_c_168_n N_VGND_c_879_n 0.00585385f $X=1.285 $Y=0.765 $X2=0 $Y2=0
cc_180 N_GATE_N_c_168_n N_VGND_c_881_n 0.00822221f $X=1.285 $Y=0.765 $X2=0 $Y2=0
cc_181 GATE_N N_VGND_c_881_n 0.00476953f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_182 N_A_47_47#_c_218_n N_A_387_385#_M1001_s 0.00120072f $X=1.875 $Y=2.9 $X2=0
+ $Y2=0
cc_183 N_A_47_47#_c_220_n N_A_387_385#_M1001_s 0.00624878f $X=1.96 $Y=2.815
+ $X2=0 $Y2=0
cc_184 N_A_47_47#_c_239_p N_A_387_385#_M1001_s 0.0080818f $X=2.66 $Y=2.4 $X2=0
+ $Y2=0
cc_185 N_A_47_47#_c_221_n N_A_387_385#_M1001_s 0.00211295f $X=2.045 $Y=2.4 $X2=0
+ $Y2=0
cc_186 N_A_47_47#_c_239_p N_A_387_385#_M1003_g 5.72527e-19 $X=2.66 $Y=2.4 $X2=0
+ $Y2=0
cc_187 N_A_47_47#_M1012_g N_A_387_385#_c_318_n 3.61442e-19 $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_188 N_A_47_47#_c_239_p N_A_387_385#_c_318_n 0.0161875f $X=2.66 $Y=2.4 $X2=0
+ $Y2=0
cc_189 N_A_47_47#_c_221_n N_A_387_385#_c_318_n 0.0116852f $X=2.045 $Y=2.4 $X2=0
+ $Y2=0
cc_190 N_A_47_47#_c_222_n N_A_387_385#_c_318_n 0.0291278f $X=2.825 $Y=1.52 $X2=0
+ $Y2=0
cc_191 N_A_47_47#_c_213_n N_A_387_385#_c_318_n 0.00101062f $X=2.825 $Y=1.52
+ $X2=0 $Y2=0
cc_192 N_A_47_47#_M1012_g N_A_387_385#_c_309_n 0.00856884f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_193 N_A_47_47#_c_222_n N_A_387_385#_c_309_n 0.0256196f $X=2.825 $Y=1.52 $X2=0
+ $Y2=0
cc_194 N_A_47_47#_c_213_n N_A_387_385#_c_309_n 0.00445034f $X=2.825 $Y=1.52
+ $X2=0 $Y2=0
cc_195 N_A_47_47#_M1012_g N_A_387_385#_c_310_n 0.0130086f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_196 N_A_47_47#_M1012_g N_A_387_385#_c_311_n 6.6765e-19 $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_197 N_A_47_47#_M1012_g N_A_387_385#_c_314_n 0.00360829f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_198 N_A_47_47#_M1012_g N_A_387_385#_c_315_n 0.00806255f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_199 N_A_47_47#_M1004_g N_A_387_385#_c_315_n 9.95958e-19 $X=2.915 $Y=2.555
+ $X2=0 $Y2=0
cc_200 N_A_47_47#_c_222_n N_A_387_385#_c_315_n 0.0410594f $X=2.825 $Y=1.52 $X2=0
+ $Y2=0
cc_201 N_A_47_47#_M1004_g N_A_387_385#_c_320_n 0.073737f $X=2.915 $Y=2.555 $X2=0
+ $Y2=0
cc_202 N_A_47_47#_c_222_n N_A_387_385#_c_320_n 0.0020676f $X=2.825 $Y=1.52 $X2=0
+ $Y2=0
cc_203 N_A_47_47#_c_218_n N_A_270_465#_M1011_d 0.00296578f $X=1.875 $Y=2.9 $X2=0
+ $Y2=0
cc_204 N_A_47_47#_M1012_g N_A_270_465#_c_408_n 0.0087168f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_205 N_A_47_47#_M1012_g N_A_270_465#_c_410_n 0.0185783f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_206 N_A_47_47#_c_218_n N_A_270_465#_M1001_g 0.0035232f $X=1.875 $Y=2.9 $X2=0
+ $Y2=0
cc_207 N_A_47_47#_c_220_n N_A_270_465#_M1001_g 0.00814904f $X=1.96 $Y=2.815
+ $X2=0 $Y2=0
cc_208 N_A_47_47#_c_239_p N_A_270_465#_M1001_g 0.0184092f $X=2.66 $Y=2.4 $X2=0
+ $Y2=0
cc_209 N_A_47_47#_M1012_g N_A_270_465#_c_411_n 0.0120518f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_210 N_A_47_47#_M1012_g N_A_270_465#_M1015_g 0.0482648f $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_211 N_A_47_47#_c_217_n N_A_270_465#_c_415_n 0.00759985f $X=1.065 $Y=2.26
+ $X2=0 $Y2=0
cc_212 N_A_47_47#_c_217_n N_A_270_465#_c_421_n 0.00246742f $X=1.065 $Y=2.26
+ $X2=0 $Y2=0
cc_213 N_A_47_47#_c_218_n N_A_270_465#_c_421_n 0.0218442f $X=1.875 $Y=2.9 $X2=0
+ $Y2=0
cc_214 N_A_47_47#_c_220_n N_A_270_465#_c_421_n 0.0117657f $X=1.96 $Y=2.815 $X2=0
+ $Y2=0
cc_215 N_A_47_47#_c_221_n N_A_270_465#_c_421_n 0.0149366f $X=2.045 $Y=2.4 $X2=0
+ $Y2=0
cc_216 N_A_47_47#_M1004_g N_A_270_465#_c_417_n 0.0292974f $X=2.915 $Y=2.555
+ $X2=0 $Y2=0
cc_217 N_A_47_47#_c_239_p N_A_270_465#_c_417_n 0.00208085f $X=2.66 $Y=2.4 $X2=0
+ $Y2=0
cc_218 N_A_47_47#_c_221_n N_A_270_465#_c_417_n 0.00191283f $X=2.045 $Y=2.4 $X2=0
+ $Y2=0
cc_219 N_A_47_47#_c_222_n N_A_270_465#_c_417_n 0.00988122f $X=2.825 $Y=1.52
+ $X2=0 $Y2=0
cc_220 N_A_47_47#_c_213_n N_A_270_465#_c_417_n 0.0227381f $X=2.825 $Y=1.52 $X2=0
+ $Y2=0
cc_221 N_A_47_47#_M1012_g N_A_670_125#_c_635_n 2.02503e-19 $X=2.915 $Y=0.835
+ $X2=0 $Y2=0
cc_222 N_A_47_47#_M1004_g N_A_670_125#_c_633_n 0.00179252f $X=2.915 $Y=2.555
+ $X2=0 $Y2=0
cc_223 N_A_47_47#_c_239_p N_A_670_125#_c_633_n 0.00777134f $X=2.66 $Y=2.4 $X2=0
+ $Y2=0
cc_224 N_A_47_47#_c_222_n N_A_670_125#_c_633_n 0.00299881f $X=2.825 $Y=1.52
+ $X2=0 $Y2=0
cc_225 N_A_47_47#_M1004_g N_A_670_125#_c_629_n 3.87407e-19 $X=2.915 $Y=2.555
+ $X2=0 $Y2=0
cc_226 N_A_47_47#_c_222_n N_A_670_125#_c_629_n 0.00459713f $X=2.825 $Y=1.52
+ $X2=0 $Y2=0
cc_227 N_A_47_47#_c_217_n N_VPWR_M1008_d 0.00855316f $X=1.065 $Y=2.26 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_47_47#_c_230_n N_VPWR_M1008_d 0.00527728f $X=1.15 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_229 N_A_47_47#_c_219_n N_VPWR_M1008_d 0.00143624f $X=1.235 $Y=2.9 $X2=-0.19
+ $Y2=-0.245
cc_230 N_A_47_47#_c_239_p N_VPWR_M1001_d 0.00702377f $X=2.66 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A_47_47#_c_222_n N_VPWR_M1001_d 9.96038e-19 $X=2.825 $Y=1.52 $X2=0
+ $Y2=0
cc_232 N_A_47_47#_c_216_n N_VPWR_c_759_n 0.00125589f $X=0.36 $Y=2.47 $X2=0 $Y2=0
cc_233 N_A_47_47#_c_217_n N_VPWR_c_759_n 0.015214f $X=1.065 $Y=2.26 $X2=0 $Y2=0
cc_234 N_A_47_47#_c_230_n N_VPWR_c_759_n 0.0221042f $X=1.15 $Y=2.815 $X2=0 $Y2=0
cc_235 N_A_47_47#_c_219_n N_VPWR_c_759_n 0.0140935f $X=1.235 $Y=2.9 $X2=0 $Y2=0
cc_236 N_A_47_47#_M1004_g N_VPWR_c_760_n 0.00370729f $X=2.915 $Y=2.555 $X2=0
+ $Y2=0
cc_237 N_A_47_47#_c_218_n N_VPWR_c_760_n 0.00616379f $X=1.875 $Y=2.9 $X2=0 $Y2=0
cc_238 N_A_47_47#_c_239_p N_VPWR_c_760_n 0.020144f $X=2.66 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A_47_47#_c_218_n N_VPWR_c_766_n 0.0337576f $X=1.875 $Y=2.9 $X2=0 $Y2=0
cc_240 N_A_47_47#_c_219_n N_VPWR_c_766_n 0.00763527f $X=1.235 $Y=2.9 $X2=0 $Y2=0
cc_241 N_A_47_47#_M1004_g N_VPWR_c_767_n 0.00517164f $X=2.915 $Y=2.555 $X2=0
+ $Y2=0
cc_242 N_A_47_47#_M1004_g N_VPWR_c_758_n 0.00519032f $X=2.915 $Y=2.555 $X2=0
+ $Y2=0
cc_243 N_A_47_47#_c_216_n N_VPWR_c_758_n 0.00992777f $X=0.36 $Y=2.47 $X2=0 $Y2=0
cc_244 N_A_47_47#_c_218_n N_VPWR_c_758_n 0.0284471f $X=1.875 $Y=2.9 $X2=0 $Y2=0
cc_245 N_A_47_47#_c_219_n N_VPWR_c_758_n 0.00612903f $X=1.235 $Y=2.9 $X2=0 $Y2=0
cc_246 N_A_47_47#_c_239_p N_VPWR_c_758_n 0.0219985f $X=2.66 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_47_47#_c_216_n N_VPWR_c_770_n 0.0122031f $X=0.36 $Y=2.47 $X2=0 $Y2=0
cc_248 N_A_47_47#_M1012_g N_VGND_c_871_n 0.00357265f $X=2.915 $Y=0.835 $X2=0
+ $Y2=0
cc_249 N_A_47_47#_c_212_n N_VGND_c_878_n 0.0138111f $X=0.36 $Y=0.465 $X2=0 $Y2=0
cc_250 N_A_47_47#_M1018_s N_VGND_c_881_n 0.00377973f $X=0.235 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_47_47#_M1012_g N_VGND_c_881_n 5.38325e-19 $X=2.915 $Y=0.835 $X2=0
+ $Y2=0
cc_252 N_A_47_47#_c_212_n N_VGND_c_881_n 0.00980511f $X=0.36 $Y=0.465 $X2=0
+ $Y2=0
cc_253 N_A_387_385#_c_308_n N_A_270_465#_c_407_n 0.00990191f $X=2.14 $Y=0.85
+ $X2=0 $Y2=0
cc_254 N_A_387_385#_c_343_p N_A_270_465#_c_407_n 6.82956e-19 $X=2.08 $Y=1.18
+ $X2=0 $Y2=0
cc_255 N_A_387_385#_c_308_n N_A_270_465#_c_408_n 0.00398135f $X=2.14 $Y=0.85
+ $X2=0 $Y2=0
cc_256 N_A_387_385#_c_311_n N_A_270_465#_c_408_n 0.00543698f $X=3.145 $Y=0.375
+ $X2=0 $Y2=0
cc_257 N_A_387_385#_c_313_n N_A_270_465#_c_408_n 0.0218994f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_258 N_A_387_385#_c_308_n N_A_270_465#_c_410_n 0.00177837f $X=2.14 $Y=0.85
+ $X2=0 $Y2=0
cc_259 N_A_387_385#_c_309_n N_A_270_465#_c_410_n 0.00876678f $X=2.925 $Y=1.18
+ $X2=0 $Y2=0
cc_260 N_A_387_385#_c_310_n N_A_270_465#_c_410_n 8.3592e-19 $X=3.035 $Y=1.095
+ $X2=0 $Y2=0
cc_261 N_A_387_385#_c_318_n N_A_270_465#_M1001_g 0.00173365f $X=2.08 $Y=2.06
+ $X2=0 $Y2=0
cc_262 N_A_387_385#_c_314_n N_A_270_465#_c_411_n 0.0050303f $X=3.33 $Y=1.265
+ $X2=0 $Y2=0
cc_263 N_A_387_385#_c_315_n N_A_270_465#_c_411_n 0.00900246f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_264 N_A_387_385#_c_320_n N_A_270_465#_c_411_n 0.0205951f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_265 N_A_387_385#_c_316_n N_A_270_465#_c_411_n 0.00103842f $X=3.725 $Y=0.515
+ $X2=0 $Y2=0
cc_266 N_A_387_385#_c_310_n N_A_270_465#_M1015_g 0.00497935f $X=3.035 $Y=1.095
+ $X2=0 $Y2=0
cc_267 N_A_387_385#_c_312_n N_A_270_465#_M1015_g 0.015166f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_268 N_A_387_385#_c_314_n N_A_270_465#_M1015_g 0.00538928f $X=3.33 $Y=1.265
+ $X2=0 $Y2=0
cc_269 N_A_387_385#_c_316_n N_A_270_465#_M1015_g 0.0117965f $X=3.725 $Y=0.515
+ $X2=0 $Y2=0
cc_270 N_A_387_385#_c_314_n N_A_270_465#_c_413_n 4.71716e-19 $X=3.33 $Y=1.265
+ $X2=0 $Y2=0
cc_271 N_A_387_385#_c_315_n N_A_270_465#_c_413_n 0.00513632f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_272 N_A_387_385#_c_316_n N_A_270_465#_c_413_n 0.00972241f $X=3.725 $Y=0.515
+ $X2=0 $Y2=0
cc_273 N_A_387_385#_M1003_g N_A_270_465#_M1016_g 0.0120823f $X=3.275 $Y=2.555
+ $X2=0 $Y2=0
cc_274 N_A_387_385#_c_315_n N_A_270_465#_M1016_g 0.0014707f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_275 N_A_387_385#_c_320_n N_A_270_465#_M1016_g 0.0203599f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_276 N_A_387_385#_c_308_n N_A_270_465#_c_415_n 0.0266922f $X=2.14 $Y=0.85
+ $X2=0 $Y2=0
cc_277 N_A_387_385#_c_318_n N_A_270_465#_c_415_n 0.0564881f $X=2.08 $Y=2.06
+ $X2=0 $Y2=0
cc_278 N_A_387_385#_c_343_p N_A_270_465#_c_415_n 0.0112872f $X=2.08 $Y=1.18
+ $X2=0 $Y2=0
cc_279 N_A_387_385#_c_318_n N_A_270_465#_c_417_n 0.0481927f $X=2.08 $Y=2.06
+ $X2=0 $Y2=0
cc_280 N_A_387_385#_c_309_n N_A_270_465#_c_417_n 0.0135643f $X=2.925 $Y=1.18
+ $X2=0 $Y2=0
cc_281 N_A_387_385#_c_343_p N_A_270_465#_c_417_n 0.00915731f $X=2.08 $Y=1.18
+ $X2=0 $Y2=0
cc_282 N_A_387_385#_c_313_n N_A_820_99#_M1019_g 0.00129738f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_283 N_A_387_385#_c_316_n N_A_820_99#_M1019_g 0.0240821f $X=3.725 $Y=0.515
+ $X2=0 $Y2=0
cc_284 N_A_387_385#_c_312_n N_A_670_125#_c_635_n 0.0301332f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_285 N_A_387_385#_c_313_n N_A_670_125#_c_635_n 0.00147959f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_286 N_A_387_385#_c_314_n N_A_670_125#_c_635_n 0.00790827f $X=3.33 $Y=1.265
+ $X2=0 $Y2=0
cc_287 N_A_387_385#_c_316_n N_A_670_125#_c_635_n 0.00694068f $X=3.725 $Y=0.515
+ $X2=0 $Y2=0
cc_288 N_A_387_385#_c_310_n N_A_670_125#_c_645_n 0.00260574f $X=3.035 $Y=1.095
+ $X2=0 $Y2=0
cc_289 N_A_387_385#_c_316_n N_A_670_125#_c_645_n 0.00329447f $X=3.725 $Y=0.515
+ $X2=0 $Y2=0
cc_290 N_A_387_385#_c_312_n N_A_670_125#_c_627_n 0.00263325f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_291 N_A_387_385#_c_313_n N_A_670_125#_c_627_n 0.0015149f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_292 N_A_387_385#_M1003_g N_A_670_125#_c_633_n 0.00997211f $X=3.275 $Y=2.555
+ $X2=0 $Y2=0
cc_293 N_A_387_385#_c_315_n N_A_670_125#_c_633_n 0.00765302f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_294 N_A_387_385#_c_320_n N_A_670_125#_c_633_n 0.00379559f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_295 N_A_387_385#_M1003_g N_A_670_125#_c_629_n 0.00153148f $X=3.275 $Y=2.555
+ $X2=0 $Y2=0
cc_296 N_A_387_385#_c_314_n N_A_670_125#_c_629_n 0.00241129f $X=3.33 $Y=1.265
+ $X2=0 $Y2=0
cc_297 N_A_387_385#_c_315_n N_A_670_125#_c_629_n 0.0605397f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_298 N_A_387_385#_c_320_n N_A_670_125#_c_629_n 0.00200461f $X=3.365 $Y=1.91
+ $X2=0 $Y2=0
cc_299 N_A_387_385#_c_310_n N_A_670_125#_c_630_n 0.00110084f $X=3.035 $Y=1.095
+ $X2=0 $Y2=0
cc_300 N_A_387_385#_c_314_n N_A_670_125#_c_630_n 0.0126644f $X=3.33 $Y=1.265
+ $X2=0 $Y2=0
cc_301 N_A_387_385#_c_316_n N_A_670_125#_c_630_n 0.00451857f $X=3.725 $Y=0.515
+ $X2=0 $Y2=0
cc_302 N_A_387_385#_M1003_g N_VPWR_c_767_n 0.00508842f $X=3.275 $Y=2.555 $X2=0
+ $Y2=0
cc_303 N_A_387_385#_M1003_g N_VPWR_c_758_n 0.00519032f $X=3.275 $Y=2.555 $X2=0
+ $Y2=0
cc_304 N_A_387_385#_c_309_n N_VGND_c_871_n 0.0243655f $X=2.925 $Y=1.18 $X2=0
+ $Y2=0
cc_305 N_A_387_385#_c_310_n N_VGND_c_871_n 0.0325666f $X=3.035 $Y=1.095 $X2=0
+ $Y2=0
cc_306 N_A_387_385#_c_311_n N_VGND_c_871_n 0.0212305f $X=3.145 $Y=0.375 $X2=0
+ $Y2=0
cc_307 N_A_387_385#_c_312_n N_VGND_c_872_n 0.0120133f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_308 N_A_387_385#_c_313_n N_VGND_c_872_n 0.00337756f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_309 N_A_387_385#_c_316_n N_VGND_c_872_n 9.57027e-19 $X=3.725 $Y=0.515 $X2=0
+ $Y2=0
cc_310 N_A_387_385#_c_311_n N_VGND_c_874_n 0.0149979f $X=3.145 $Y=0.375 $X2=0
+ $Y2=0
cc_311 N_A_387_385#_c_312_n N_VGND_c_874_n 0.0476644f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_312 N_A_387_385#_c_313_n N_VGND_c_874_n 0.00647615f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_313 N_A_387_385#_c_308_n N_VGND_c_879_n 0.00572179f $X=2.14 $Y=0.85 $X2=0
+ $Y2=0
cc_314 N_A_387_385#_c_308_n N_VGND_c_881_n 0.00825693f $X=2.14 $Y=0.85 $X2=0
+ $Y2=0
cc_315 N_A_387_385#_c_311_n N_VGND_c_881_n 0.00754646f $X=3.145 $Y=0.375 $X2=0
+ $Y2=0
cc_316 N_A_387_385#_c_312_n N_VGND_c_881_n 0.0257792f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_317 N_A_387_385#_c_313_n N_VGND_c_881_n 0.00941423f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_318 N_A_270_465#_c_411_n N_A_820_99#_M1019_g 0.0018922f $X=3.275 $Y=1.155
+ $X2=0 $Y2=0
cc_319 N_A_270_465#_c_413_n N_A_820_99#_M1019_g 0.0413027f $X=3.74 $Y=1.46 $X2=0
+ $Y2=0
cc_320 N_A_270_465#_M1016_g N_A_820_99#_c_512_n 0.0413027f $X=3.815 $Y=2.445
+ $X2=0 $Y2=0
cc_321 N_A_270_465#_c_413_n N_A_820_99#_c_516_n 0.00230089f $X=3.74 $Y=1.46
+ $X2=0 $Y2=0
cc_322 N_A_270_465#_M1015_g N_A_670_125#_c_635_n 0.00330952f $X=3.275 $Y=0.835
+ $X2=0 $Y2=0
cc_323 N_A_270_465#_c_413_n N_A_670_125#_c_635_n 0.00372305f $X=3.74 $Y=1.46
+ $X2=0 $Y2=0
cc_324 N_A_270_465#_M1015_g N_A_670_125#_c_645_n 2.62598e-19 $X=3.275 $Y=0.835
+ $X2=0 $Y2=0
cc_325 N_A_270_465#_c_413_n N_A_670_125#_c_627_n 0.00379958f $X=3.74 $Y=1.46
+ $X2=0 $Y2=0
cc_326 N_A_270_465#_M1016_g N_A_670_125#_c_633_n 0.0193825f $X=3.815 $Y=2.445
+ $X2=0 $Y2=0
cc_327 N_A_270_465#_c_411_n N_A_670_125#_c_629_n 5.15196e-19 $X=3.275 $Y=1.155
+ $X2=0 $Y2=0
cc_328 N_A_270_465#_c_413_n N_A_670_125#_c_629_n 0.0103026f $X=3.74 $Y=1.46
+ $X2=0 $Y2=0
cc_329 N_A_270_465#_M1016_g N_A_670_125#_c_629_n 0.017866f $X=3.815 $Y=2.445
+ $X2=0 $Y2=0
cc_330 N_A_270_465#_c_411_n N_A_670_125#_c_630_n 2.73169e-19 $X=3.275 $Y=1.155
+ $X2=0 $Y2=0
cc_331 N_A_270_465#_M1001_g N_VPWR_c_760_n 0.0021075f $X=2.41 $Y=2.555 $X2=0
+ $Y2=0
cc_332 N_A_270_465#_M1001_g N_VPWR_c_766_n 0.00517164f $X=2.41 $Y=2.555 $X2=0
+ $Y2=0
cc_333 N_A_270_465#_M1016_g N_VPWR_c_767_n 0.00260298f $X=3.815 $Y=2.445 $X2=0
+ $Y2=0
cc_334 N_A_270_465#_M1001_g N_VPWR_c_758_n 0.00519032f $X=2.41 $Y=2.555 $X2=0
+ $Y2=0
cc_335 N_A_270_465#_M1016_g N_VPWR_c_758_n 0.00276537f $X=3.815 $Y=2.445 $X2=0
+ $Y2=0
cc_336 N_A_270_465#_c_407_n N_VGND_c_871_n 0.00506056f $X=1.865 $Y=1.155 $X2=0
+ $Y2=0
cc_337 N_A_270_465#_c_408_n N_VGND_c_871_n 0.0255017f $X=3.2 $Y=0.18 $X2=0 $Y2=0
cc_338 N_A_270_465#_c_410_n N_VGND_c_871_n 0.00845289f $X=2.375 $Y=1.155 $X2=0
+ $Y2=0
cc_339 N_A_270_465#_M1015_g N_VGND_c_871_n 9.86783e-19 $X=3.275 $Y=0.835 $X2=0
+ $Y2=0
cc_340 N_A_270_465#_c_408_n N_VGND_c_874_n 0.0154091f $X=3.2 $Y=0.18 $X2=0 $Y2=0
cc_341 N_A_270_465#_c_409_n N_VGND_c_879_n 0.0199199f $X=1.94 $Y=0.18 $X2=0
+ $Y2=0
cc_342 N_A_270_465#_c_416_n N_VGND_c_879_n 0.0160982f $X=1.6 $Y=0.465 $X2=0
+ $Y2=0
cc_343 N_A_270_465#_M1002_d N_VGND_c_881_n 0.00269994f $X=1.36 $Y=0.235 $X2=0
+ $Y2=0
cc_344 N_A_270_465#_c_408_n N_VGND_c_881_n 0.0344474f $X=3.2 $Y=0.18 $X2=0 $Y2=0
cc_345 N_A_270_465#_c_409_n N_VGND_c_881_n 0.00974353f $X=1.94 $Y=0.18 $X2=0
+ $Y2=0
cc_346 N_A_270_465#_c_410_n N_VGND_c_881_n 7.97988e-19 $X=2.375 $Y=1.155 $X2=0
+ $Y2=0
cc_347 N_A_270_465#_c_416_n N_VGND_c_881_n 0.0122742f $X=1.6 $Y=0.465 $X2=0
+ $Y2=0
cc_348 N_A_820_99#_c_523_n N_A_670_125#_M1000_g 0.0127381f $X=5.075 $Y=1.77
+ $X2=0 $Y2=0
cc_349 N_A_820_99#_c_513_n N_A_670_125#_M1000_g 0.00494502f $X=5.165 $Y=1.685
+ $X2=0 $Y2=0
cc_350 N_A_820_99#_c_536_p N_A_670_125#_M1000_g 0.00984148f $X=5.17 $Y=2.3 $X2=0
+ $Y2=0
cc_351 N_A_820_99#_c_516_n N_A_670_125#_M1000_g 0.00129078f $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_352 N_A_820_99#_c_517_n N_A_670_125#_M1000_g 0.00916505f $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_353 N_A_820_99#_c_527_n N_A_670_125#_M1000_g 0.0025012f $X=5.165 $Y=1.77
+ $X2=0 $Y2=0
cc_354 N_A_820_99#_c_540_p N_A_670_125#_M1000_g 0.0101998f $X=5.27 $Y=2.465
+ $X2=0 $Y2=0
cc_355 N_A_820_99#_c_513_n N_A_670_125#_c_626_n 0.0117383f $X=5.165 $Y=1.685
+ $X2=0 $Y2=0
cc_356 N_A_820_99#_c_518_n N_A_670_125#_c_626_n 0.0122939f $X=4.91 $Y=0.43 $X2=0
+ $Y2=0
cc_357 N_A_820_99#_M1019_g N_A_670_125#_c_645_n 6.83666e-19 $X=4.175 $Y=0.835
+ $X2=0 $Y2=0
cc_358 N_A_820_99#_M1013_s N_A_670_125#_c_627_n 0.00145019f $X=4.785 $Y=0.235
+ $X2=0 $Y2=0
cc_359 N_A_820_99#_M1019_g N_A_670_125#_c_627_n 0.0161703f $X=4.175 $Y=0.835
+ $X2=0 $Y2=0
cc_360 N_A_820_99#_c_523_n N_A_670_125#_c_627_n 0.00862788f $X=5.075 $Y=1.77
+ $X2=0 $Y2=0
cc_361 N_A_820_99#_c_513_n N_A_670_125#_c_627_n 0.0134898f $X=5.165 $Y=1.685
+ $X2=0 $Y2=0
cc_362 N_A_820_99#_c_516_n N_A_670_125#_c_627_n 0.0256239f $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_363 N_A_820_99#_c_517_n N_A_670_125#_c_627_n 0.00124654f $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_364 N_A_820_99#_c_518_n N_A_670_125#_c_627_n 0.0127261f $X=4.91 $Y=0.43 $X2=0
+ $Y2=0
cc_365 N_A_820_99#_M1019_g N_A_670_125#_c_628_n 9.70365e-19 $X=4.175 $Y=0.835
+ $X2=0 $Y2=0
cc_366 N_A_820_99#_c_523_n N_A_670_125#_c_628_n 0.019183f $X=5.075 $Y=1.77 $X2=0
+ $Y2=0
cc_367 N_A_820_99#_c_513_n N_A_670_125#_c_628_n 0.0196058f $X=5.165 $Y=1.685
+ $X2=0 $Y2=0
cc_368 N_A_820_99#_c_516_n N_A_670_125#_c_628_n 0.00646041f $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_369 N_A_820_99#_c_517_n N_A_670_125#_c_628_n 3.95101e-19 $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_370 N_A_820_99#_c_512_n N_A_670_125#_c_633_n 0.00239017f $X=4.265 $Y=1.91
+ $X2=0 $Y2=0
cc_371 N_A_820_99#_M1019_g N_A_670_125#_c_629_n 0.00550992f $X=4.175 $Y=0.835
+ $X2=0 $Y2=0
cc_372 N_A_820_99#_c_516_n N_A_670_125#_c_629_n 0.0303091f $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_373 N_A_820_99#_M1019_g N_A_670_125#_c_631_n 0.00714438f $X=4.175 $Y=0.835
+ $X2=0 $Y2=0
cc_374 N_A_820_99#_c_523_n N_A_670_125#_c_631_n 0.00460331f $X=5.075 $Y=1.77
+ $X2=0 $Y2=0
cc_375 N_A_820_99#_c_513_n N_A_670_125#_c_631_n 0.0105709f $X=5.165 $Y=1.685
+ $X2=0 $Y2=0
cc_376 N_A_820_99#_c_516_n N_A_670_125#_c_631_n 4.22693e-19 $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_377 N_A_820_99#_c_517_n N_A_670_125#_c_631_n 0.00633707f $X=4.265 $Y=1.57
+ $X2=0 $Y2=0
cc_378 N_A_820_99#_c_518_n N_A_670_125#_c_631_n 0.00540271f $X=4.91 $Y=0.43
+ $X2=0 $Y2=0
cc_379 N_A_820_99#_c_536_p N_RESET_B_M1007_g 0.00502514f $X=5.17 $Y=2.3 $X2=0
+ $Y2=0
cc_380 N_A_820_99#_c_566_p N_RESET_B_M1007_g 0.0110202f $X=5.95 $Y=2.385 $X2=0
+ $Y2=0
cc_381 N_A_820_99#_c_514_n N_RESET_B_M1007_g 0.00159622f $X=6.115 $Y=1.51 $X2=0
+ $Y2=0
cc_382 N_A_820_99#_c_515_n N_RESET_B_M1007_g 0.0408094f $X=6.115 $Y=1.51 $X2=0
+ $Y2=0
cc_383 N_A_820_99#_c_527_n N_RESET_B_M1007_g 0.00111966f $X=5.165 $Y=1.77 $X2=0
+ $Y2=0
cc_384 N_A_820_99#_M1010_g RESET_B 0.00445543f $X=6.025 $Y=0.655 $X2=0 $Y2=0
cc_385 N_A_820_99#_c_513_n RESET_B 0.0544873f $X=5.165 $Y=1.685 $X2=0 $Y2=0
cc_386 N_A_820_99#_c_536_p RESET_B 0.0201957f $X=5.17 $Y=2.3 $X2=0 $Y2=0
cc_387 N_A_820_99#_c_566_p RESET_B 0.0201332f $X=5.95 $Y=2.385 $X2=0 $Y2=0
cc_388 N_A_820_99#_c_514_n RESET_B 0.0506066f $X=6.115 $Y=1.51 $X2=0 $Y2=0
cc_389 N_A_820_99#_c_515_n RESET_B 0.00441571f $X=6.115 $Y=1.51 $X2=0 $Y2=0
cc_390 N_A_820_99#_c_527_n RESET_B 0.0142558f $X=5.165 $Y=1.77 $X2=0 $Y2=0
cc_391 N_A_820_99#_M1010_g N_RESET_B_c_718_n 0.020219f $X=6.025 $Y=0.655 $X2=0
+ $Y2=0
cc_392 N_A_820_99#_c_514_n N_RESET_B_c_718_n 5.92853e-19 $X=6.115 $Y=1.51 $X2=0
+ $Y2=0
cc_393 N_A_820_99#_M1010_g N_RESET_B_c_719_n 0.018866f $X=6.025 $Y=0.655 $X2=0
+ $Y2=0
cc_394 N_A_820_99#_c_513_n N_RESET_B_c_719_n 0.00546758f $X=5.165 $Y=1.685 $X2=0
+ $Y2=0
cc_395 N_A_820_99#_c_523_n N_VPWR_M1014_d 0.00281272f $X=5.075 $Y=1.77 $X2=0
+ $Y2=0
cc_396 N_A_820_99#_c_566_p N_VPWR_M1007_d 0.0103501f $X=5.95 $Y=2.385 $X2=0
+ $Y2=0
cc_397 N_A_820_99#_M1014_g N_VPWR_c_761_n 0.00554376f $X=4.175 $Y=2.445 $X2=0
+ $Y2=0
cc_398 N_A_820_99#_c_522_n N_VPWR_c_761_n 0.00144589f $X=4.265 $Y=2.075 $X2=0
+ $Y2=0
cc_399 N_A_820_99#_c_523_n N_VPWR_c_761_n 0.0310234f $X=5.075 $Y=1.77 $X2=0
+ $Y2=0
cc_400 N_A_820_99#_c_536_p N_VPWR_c_761_n 0.0201404f $X=5.17 $Y=2.3 $X2=0 $Y2=0
cc_401 N_A_820_99#_c_516_n N_VPWR_c_761_n 0.0126848f $X=4.265 $Y=1.57 $X2=0
+ $Y2=0
cc_402 N_A_820_99#_c_540_p N_VPWR_c_761_n 0.0248948f $X=5.27 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_820_99#_M1014_g N_VPWR_c_762_n 0.00395146f $X=4.175 $Y=2.445 $X2=0
+ $Y2=0
cc_404 N_A_820_99#_c_540_p N_VPWR_c_762_n 0.0388509f $X=5.27 $Y=2.465 $X2=0
+ $Y2=0
cc_405 N_A_820_99#_M1017_g N_VPWR_c_763_n 0.00571734f $X=6.025 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_A_820_99#_c_566_p N_VPWR_c_763_n 0.0219993f $X=5.95 $Y=2.385 $X2=0
+ $Y2=0
cc_407 N_A_820_99#_c_540_p N_VPWR_c_764_n 0.0177611f $X=5.27 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_A_820_99#_M1014_g N_VPWR_c_767_n 0.00389919f $X=4.175 $Y=2.445 $X2=0
+ $Y2=0
cc_409 N_A_820_99#_M1017_g N_VPWR_c_768_n 0.00550964f $X=6.025 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_A_820_99#_M1000_d N_VPWR_c_758_n 0.0023939f $X=5.13 $Y=1.835 $X2=0
+ $Y2=0
cc_411 N_A_820_99#_M1014_g N_VPWR_c_758_n 0.00455831f $X=4.175 $Y=2.445 $X2=0
+ $Y2=0
cc_412 N_A_820_99#_M1017_g N_VPWR_c_758_n 0.00770762f $X=6.025 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A_820_99#_c_566_p N_VPWR_c_758_n 0.0119156f $X=5.95 $Y=2.385 $X2=0
+ $Y2=0
cc_414 N_A_820_99#_c_540_p N_VPWR_c_758_n 0.011311f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_415 N_A_820_99#_c_566_p N_Q_M1017_d 0.00234612f $X=5.95 $Y=2.385 $X2=0 $Y2=0
cc_416 N_A_820_99#_c_514_n N_Q_M1017_d 0.00500356f $X=6.115 $Y=1.51 $X2=0 $Y2=0
cc_417 N_A_820_99#_M1017_g N_Q_c_845_n 0.00403788f $X=6.025 $Y=2.465 $X2=0 $Y2=0
cc_418 N_A_820_99#_c_566_p N_Q_c_845_n 0.00544159f $X=5.95 $Y=2.385 $X2=0 $Y2=0
cc_419 N_A_820_99#_M1010_g Q 0.00435261f $X=6.025 $Y=0.655 $X2=0 $Y2=0
cc_420 N_A_820_99#_c_514_n Q 0.00716064f $X=6.115 $Y=1.51 $X2=0 $Y2=0
cc_421 N_A_820_99#_c_515_n Q 0.00405119f $X=6.115 $Y=1.51 $X2=0 $Y2=0
cc_422 N_A_820_99#_M1010_g Q 0.00534456f $X=6.025 $Y=0.655 $X2=0 $Y2=0
cc_423 N_A_820_99#_M1017_g Q 0.009612f $X=6.025 $Y=2.465 $X2=0 $Y2=0
cc_424 N_A_820_99#_c_566_p Q 0.0145039f $X=5.95 $Y=2.385 $X2=0 $Y2=0
cc_425 N_A_820_99#_c_514_n Q 0.0745562f $X=6.115 $Y=1.51 $X2=0 $Y2=0
cc_426 N_A_820_99#_c_515_n Q 0.0082253f $X=6.115 $Y=1.51 $X2=0 $Y2=0
cc_427 N_A_820_99#_M1010_g N_Q_c_844_n 0.00967557f $X=6.025 $Y=0.655 $X2=0 $Y2=0
cc_428 N_A_820_99#_M1019_g N_VGND_c_872_n 0.0102961f $X=4.175 $Y=0.835 $X2=0
+ $Y2=0
cc_429 N_A_820_99#_c_513_n N_VGND_c_872_n 6.43955e-19 $X=5.165 $Y=1.685 $X2=0
+ $Y2=0
cc_430 N_A_820_99#_c_518_n N_VGND_c_872_n 0.0437911f $X=4.91 $Y=0.43 $X2=0 $Y2=0
cc_431 N_A_820_99#_M1010_g N_VGND_c_873_n 0.00383036f $X=6.025 $Y=0.655 $X2=0
+ $Y2=0
cc_432 N_A_820_99#_M1019_g N_VGND_c_874_n 0.00345209f $X=4.175 $Y=0.835 $X2=0
+ $Y2=0
cc_433 N_A_820_99#_c_518_n N_VGND_c_876_n 0.0215458f $X=4.91 $Y=0.43 $X2=0 $Y2=0
cc_434 N_A_820_99#_M1010_g N_VGND_c_880_n 0.00571722f $X=6.025 $Y=0.655 $X2=0
+ $Y2=0
cc_435 N_A_820_99#_M1013_s N_VGND_c_881_n 0.00220275f $X=4.785 $Y=0.235 $X2=0
+ $Y2=0
cc_436 N_A_820_99#_M1019_g N_VGND_c_881_n 0.00394323f $X=4.175 $Y=0.835 $X2=0
+ $Y2=0
cc_437 N_A_820_99#_M1010_g N_VGND_c_881_n 0.0117608f $X=6.025 $Y=0.655 $X2=0
+ $Y2=0
cc_438 N_A_820_99#_c_518_n N_VGND_c_881_n 0.0181717f $X=4.91 $Y=0.43 $X2=0 $Y2=0
cc_439 N_A_670_125#_M1000_g N_RESET_B_M1007_g 0.023496f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_A_670_125#_c_626_n RESET_B 5.43708e-19 $X=5.125 $Y=1.185 $X2=0 $Y2=0
cc_441 N_A_670_125#_c_631_n RESET_B 8.05787e-19 $X=5.055 $Y=1.35 $X2=0 $Y2=0
cc_442 N_A_670_125#_c_631_n N_RESET_B_c_718_n 0.0607367f $X=5.055 $Y=1.35 $X2=0
+ $Y2=0
cc_443 N_A_670_125#_c_626_n N_RESET_B_c_719_n 0.0372407f $X=5.125 $Y=1.185 $X2=0
+ $Y2=0
cc_444 N_A_670_125#_c_633_n N_VPWR_c_760_n 0.00387406f $X=3.505 $Y=2.38 $X2=0
+ $Y2=0
cc_445 N_A_670_125#_M1000_g N_VPWR_c_761_n 0.00248011f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_A_670_125#_M1000_g N_VPWR_c_762_n 0.00516139f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_670_125#_c_633_n N_VPWR_c_762_n 0.0102062f $X=3.505 $Y=2.38 $X2=0
+ $Y2=0
cc_448 N_A_670_125#_M1000_g N_VPWR_c_764_n 0.00518588f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A_670_125#_c_633_n N_VPWR_c_767_n 0.0146903f $X=3.505 $Y=2.38 $X2=0
+ $Y2=0
cc_450 N_A_670_125#_M1000_g N_VPWR_c_758_n 0.0104042f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_451 N_A_670_125#_c_633_n N_VPWR_c_758_n 0.0158823f $X=3.505 $Y=2.38 $X2=0
+ $Y2=0
cc_452 N_A_670_125#_c_626_n N_VGND_c_872_n 0.00330551f $X=5.125 $Y=1.185 $X2=0
+ $Y2=0
cc_453 N_A_670_125#_c_627_n N_VGND_c_872_n 0.0244345f $X=4.655 $Y=1.15 $X2=0
+ $Y2=0
cc_454 N_A_670_125#_c_626_n N_VGND_c_876_n 0.00371894f $X=5.125 $Y=1.185 $X2=0
+ $Y2=0
cc_455 N_A_670_125#_c_626_n N_VGND_c_881_n 0.00651528f $X=5.125 $Y=1.185 $X2=0
+ $Y2=0
cc_456 RESET_B N_VPWR_M1007_d 0.00412508f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_457 N_RESET_B_M1007_g N_VPWR_c_763_n 0.00268041f $X=5.485 $Y=2.465 $X2=0
+ $Y2=0
cc_458 N_RESET_B_M1007_g N_VPWR_c_764_n 0.00585385f $X=5.485 $Y=2.465 $X2=0
+ $Y2=0
cc_459 N_RESET_B_M1007_g N_VPWR_c_758_n 0.00658858f $X=5.485 $Y=2.465 $X2=0
+ $Y2=0
cc_460 RESET_B Q 0.0117908f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_461 N_RESET_B_c_719_n Q 2.15176e-19 $X=5.575 $Y=1.185 $X2=0 $Y2=0
cc_462 RESET_B Q 0.00746504f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_463 N_RESET_B_c_719_n N_Q_c_844_n 7.04616e-19 $X=5.575 $Y=1.185 $X2=0 $Y2=0
cc_464 RESET_B N_VGND_M1005_d 0.00407639f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_465 RESET_B N_VGND_c_873_n 0.0107347f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_466 N_RESET_B_c_718_n N_VGND_c_873_n 5.24997e-19 $X=5.575 $Y=1.35 $X2=0 $Y2=0
cc_467 N_RESET_B_c_719_n N_VGND_c_873_n 0.00383036f $X=5.575 $Y=1.185 $X2=0
+ $Y2=0
cc_468 N_RESET_B_c_719_n N_VGND_c_876_n 0.00585385f $X=5.575 $Y=1.185 $X2=0
+ $Y2=0
cc_469 RESET_B N_VGND_c_881_n 0.00597407f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_470 N_RESET_B_c_719_n N_VGND_c_881_n 0.00693719f $X=5.575 $Y=1.185 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_758_n N_Q_M1017_d 0.00226663f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_472 N_VPWR_c_768_n N_Q_c_845_n 0.0213515f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_473 N_VPWR_c_758_n N_Q_c_845_n 0.0199201f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_474 N_Q_c_844_n N_VGND_c_880_n 0.0364845f $X=6.26 $Y=0.42 $X2=0 $Y2=0
cc_475 N_Q_M1010_d N_VGND_c_881_n 0.00231914f $X=6.1 $Y=0.235 $X2=0 $Y2=0
cc_476 N_Q_c_844_n N_VGND_c_881_n 0.0209962f $X=6.26 $Y=0.42 $X2=0 $Y2=0
cc_477 N_VGND_c_881_n A_1040_47# 0.00712607f $X=6.48 $Y=0 $X2=-0.19 $Y2=-0.245
