* File: sky130_fd_sc_lp__bufbuf_8.pex.spice
* Created: Wed Sep  2 09:35:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFBUF_8%A_117_265# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 77 84 86 88 89 90 91 92 95 101 103 105 109 115 117 118
+ 119
r197 128 129 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.355 $Y=1.49
+ $X2=3.785 $Y2=1.49
r198 127 128 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.925 $Y=1.49
+ $X2=3.355 $Y2=1.49
r199 126 127 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.495 $Y=1.49
+ $X2=2.925 $Y2=1.49
r200 125 126 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.065 $Y=1.49
+ $X2=2.495 $Y2=1.49
r201 124 125 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.635 $Y=1.49
+ $X2=2.065 $Y2=1.49
r202 123 124 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.205 $Y=1.49
+ $X2=1.635 $Y2=1.49
r203 122 123 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.775 $Y=1.49
+ $X2=1.205 $Y2=1.49
r204 113 115 26.5948 $w=2.58e-07 $l=6e-07 $layer=LI1_cond $X=5.37 $Y=1.055
+ $X2=5.37 $Y2=0.455
r205 109 111 31.3941 $w=2.88e-07 $l=7.9e-07 $layer=LI1_cond $X=5.355 $Y=2.05
+ $X2=5.355 $Y2=2.84
r206 107 109 4.96743 $w=2.88e-07 $l=1.25e-07 $layer=LI1_cond $X=5.355 $Y=1.925
+ $X2=5.355 $Y2=2.05
r207 106 118 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=4.61 $Y=1.84
+ $X2=4.472 $Y2=1.84
r208 105 107 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=5.21 $Y=1.84
+ $X2=5.355 $Y2=1.925
r209 105 106 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.21 $Y=1.84
+ $X2=4.61 $Y2=1.84
r210 104 119 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.57 $Y=1.14
+ $X2=4.465 $Y2=1.14
r211 103 113 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.24 $Y=1.14
+ $X2=5.37 $Y2=1.055
r212 103 104 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.24 $Y=1.14
+ $X2=4.57 $Y2=1.14
r213 99 119 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=1.055
+ $X2=4.465 $Y2=1.14
r214 99 101 31.6883 $w=2.08e-07 $l=6e-07 $layer=LI1_cond $X=4.465 $Y=1.055
+ $X2=4.465 $Y2=0.455
r215 95 97 33.1065 $w=2.73e-07 $l=7.9e-07 $layer=LI1_cond $X=4.472 $Y=2.05
+ $X2=4.472 $Y2=2.84
r216 93 118 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.472 $Y=1.925
+ $X2=4.472 $Y2=1.84
r217 93 95 5.23838 $w=2.73e-07 $l=1.25e-07 $layer=LI1_cond $X=4.472 $Y=1.925
+ $X2=4.472 $Y2=2.05
r218 91 118 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.335 $Y=1.84
+ $X2=4.472 $Y2=1.84
r219 91 92 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.335 $Y=1.84
+ $X2=4.005 $Y2=1.84
r220 89 119 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.36 $Y=1.14
+ $X2=4.465 $Y2=1.14
r221 89 90 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.36 $Y=1.14
+ $X2=4.005 $Y2=1.14
r222 88 92 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=1.755
+ $X2=4.005 $Y2=1.84
r223 87 117 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.92 $Y=1.585
+ $X2=3.92 $Y2=1.49
r224 87 88 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.92 $Y=1.585
+ $X2=3.92 $Y2=1.755
r225 86 117 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.92 $Y=1.395
+ $X2=3.92 $Y2=1.49
r226 85 90 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=1.225
+ $X2=4.005 $Y2=1.14
r227 85 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.92 $Y=1.225
+ $X2=3.92 $Y2=1.395
r228 84 129 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.81 $Y=1.49
+ $X2=3.785 $Y2=1.49
r229 83 84 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=3.81
+ $Y=1.49 $X2=3.81 $Y2=1.49
r230 80 122 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.75 $Y=1.49
+ $X2=0.775 $Y2=1.49
r231 79 83 178.622 $w=1.88e-07 $l=3.06e-06 $layer=LI1_cond $X=0.75 $Y=1.49
+ $X2=3.81 $Y2=1.49
r232 79 80 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=0.75
+ $Y=1.49 $X2=0.75 $Y2=1.49
r233 77 117 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=1.49
+ $X2=3.92 $Y2=1.49
r234 77 83 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=3.835 $Y=1.49
+ $X2=3.81 $Y2=1.49
r235 73 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.655
+ $X2=3.785 $Y2=1.49
r236 73 75 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.785 $Y=1.655
+ $X2=3.785 $Y2=2.465
r237 69 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.325
+ $X2=3.785 $Y2=1.49
r238 69 71 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.785 $Y=1.325
+ $X2=3.785 $Y2=0.665
r239 65 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.655
+ $X2=3.355 $Y2=1.49
r240 65 67 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.355 $Y=1.655
+ $X2=3.355 $Y2=2.465
r241 61 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.325
+ $X2=3.355 $Y2=1.49
r242 61 63 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.355 $Y=1.325
+ $X2=3.355 $Y2=0.665
r243 57 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.655
+ $X2=2.925 $Y2=1.49
r244 57 59 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.925 $Y=1.655
+ $X2=2.925 $Y2=2.465
r245 53 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.325
+ $X2=2.925 $Y2=1.49
r246 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.925 $Y=1.325
+ $X2=2.925 $Y2=0.665
r247 49 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.655
+ $X2=2.495 $Y2=1.49
r248 49 51 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.495 $Y=1.655
+ $X2=2.495 $Y2=2.465
r249 45 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.325
+ $X2=2.495 $Y2=1.49
r250 45 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.495 $Y=1.325
+ $X2=2.495 $Y2=0.665
r251 41 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.655
+ $X2=2.065 $Y2=1.49
r252 41 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.065 $Y=1.655
+ $X2=2.065 $Y2=2.465
r253 37 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.325
+ $X2=2.065 $Y2=1.49
r254 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.065 $Y=1.325
+ $X2=2.065 $Y2=0.665
r255 33 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.655
+ $X2=1.635 $Y2=1.49
r256 33 35 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.635 $Y=1.655
+ $X2=1.635 $Y2=2.465
r257 29 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.325
+ $X2=1.635 $Y2=1.49
r258 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.635 $Y=1.325
+ $X2=1.635 $Y2=0.665
r259 25 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.655
+ $X2=1.205 $Y2=1.49
r260 25 27 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.205 $Y=1.655
+ $X2=1.205 $Y2=2.465
r261 21 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.325
+ $X2=1.205 $Y2=1.49
r262 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.205 $Y=1.325
+ $X2=1.205 $Y2=0.665
r263 17 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.775 $Y=1.655
+ $X2=0.775 $Y2=1.49
r264 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.775 $Y=1.655
+ $X2=0.775 $Y2=2.465
r265 13 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.775 $Y=1.325
+ $X2=0.775 $Y2=1.49
r266 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.775 $Y=1.325
+ $X2=0.775 $Y2=0.665
r267 4 111 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=5.195
+ $Y=1.835 $X2=5.335 $Y2=2.84
r268 4 109 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=5.195
+ $Y=1.835 $X2=5.335 $Y2=2.05
r269 3 97 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.835 $X2=4.475 $Y2=2.84
r270 3 95 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.835 $X2=4.475 $Y2=2.05
r271 2 115 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=5.195
+ $Y=0.245 $X2=5.335 $Y2=0.455
r272 1 101 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=4.335
+ $Y=0.245 $X2=4.475 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_8%A_837_23# 1 2 9 13 17 21 25 29 31 38 41 45
+ 47 51 52 53
c88 38 0 2.74112e-19 $X=5.71 $Y=1.49
r89 59 60 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.69 $Y=1.49
+ $X2=5.12 $Y2=1.49
r90 53 60 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.195 $Y=1.49
+ $X2=5.12 $Y2=1.49
r91 47 49 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.955 $Y=1.98
+ $X2=5.955 $Y2=2.66
r92 45 52 6.33825 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.955 $Y=1.93
+ $X2=5.955 $Y2=1.815
r93 45 47 2.50531 $w=2.28e-07 $l=5e-08 $layer=LI1_cond $X=5.955 $Y=1.93
+ $X2=5.955 $Y2=1.98
r94 43 51 4.56504 $w=2.2e-07 $l=1.13248e-07 $layer=LI1_cond $X=5.93 $Y=1.585
+ $X2=5.89 $Y2=1.49
r95 43 52 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=5.93 $Y=1.585
+ $X2=5.93 $Y2=1.815
r96 39 51 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.89 $Y=1.395
+ $X2=5.89 $Y2=1.49
r97 39 41 35.2382 $w=2.58e-07 $l=7.95e-07 $layer=LI1_cond $X=5.89 $Y=1.395
+ $X2=5.89 $Y2=0.6
r98 38 53 90.0536 $w=3.3e-07 $l=5.15e-07 $layer=POLY_cond $X=5.71 $Y=1.49
+ $X2=5.195 $Y2=1.49
r99 37 38 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.71
+ $Y=1.49 $X2=5.71 $Y2=1.49
r100 34 59 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.35 $Y=1.49
+ $X2=4.69 $Y2=1.49
r101 34 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.35 $Y=1.49 $X2=4.26
+ $Y2=1.49
r102 33 37 79.3876 $w=1.88e-07 $l=1.36e-06 $layer=LI1_cond $X=4.35 $Y=1.49
+ $X2=5.71 $Y2=1.49
r103 33 34 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.35
+ $Y=1.49 $X2=4.35 $Y2=1.49
r104 31 51 1.87542 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=5.76 $Y=1.49
+ $X2=5.89 $Y2=1.49
r105 31 37 2.91866 $w=1.88e-07 $l=5e-08 $layer=LI1_cond $X=5.76 $Y=1.49 $X2=5.71
+ $Y2=1.49
r106 27 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.12 $Y=1.655
+ $X2=5.12 $Y2=1.49
r107 27 29 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.12 $Y=1.655
+ $X2=5.12 $Y2=2.465
r108 23 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.12 $Y=1.325
+ $X2=5.12 $Y2=1.49
r109 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.12 $Y=1.325
+ $X2=5.12 $Y2=0.665
r110 19 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=1.655
+ $X2=4.69 $Y2=1.49
r111 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.69 $Y=1.655
+ $X2=4.69 $Y2=2.465
r112 15 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.69 $Y2=1.49
r113 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.69 $Y2=0.665
r114 11 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.26 $Y=1.655
+ $X2=4.26 $Y2=1.49
r115 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.26 $Y=1.655
+ $X2=4.26 $Y2=2.465
r116 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.26 $Y=1.325
+ $X2=4.26 $Y2=1.49
r117 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.26 $Y=1.325
+ $X2=4.26 $Y2=0.665
r118 2 49 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=5.86
+ $Y=1.835 $X2=5.985 $Y2=2.66
r119 2 47 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.86
+ $Y=1.835 $X2=5.985 $Y2=1.98
r120 1 41 91 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_NDIFF $count=2 $X=5.8
+ $Y=0.245 $X2=5.925 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_8%A_1217_23# 1 2 9 12 17 18 20 21 22 23 25 29
+ 31 33
c59 20 0 1.12004e-19 $X=6.34 $Y=1.925
c60 17 0 1.62107e-19 $X=6.275 $Y=1.36
r61 27 29 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.94 $Y=1.065
+ $X2=6.94 $Y2=0.875
r62 23 25 20.9535 $w=2.73e-07 $l=5e-07 $layer=LI1_cond $X=6.44 $Y=2.062 $X2=6.94
+ $Y2=2.062
r63 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.775 $Y=1.15
+ $X2=6.94 $Y2=1.065
r64 21 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.775 $Y=1.15
+ $X2=6.44 $Y2=1.15
r65 20 23 7.03987 $w=2.75e-07 $l=1.80192e-07 $layer=LI1_cond $X=6.34 $Y=1.925
+ $X2=6.44 $Y2=2.062
r66 20 31 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=6.34 $Y=1.925 $X2=6.34
+ $Y2=1.525
r67 18 34 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=6.262 $Y=1.36
+ $X2=6.262 $Y2=1.525
r68 18 33 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=6.262 $Y=1.36
+ $X2=6.262 $Y2=1.195
r69 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.275
+ $Y=1.36 $X2=6.275 $Y2=1.36
r70 15 31 6.25636 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=1.4
+ $X2=6.315 $Y2=1.525
r71 15 17 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=6.315 $Y=1.4 $X2=6.315
+ $Y2=1.36
r72 14 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.315 $Y=1.235
+ $X2=6.44 $Y2=1.15
r73 14 17 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=1.235
+ $X2=6.315 $Y2=1.36
r74 12 34 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=6.2 $Y=2.465 $X2=6.2
+ $Y2=1.525
r75 9 33 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.16 $Y=0.665
+ $X2=6.16 $Y2=1.195
r76 2 25 600 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.835 $X2=6.94 $Y2=2.06
r77 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.665 $X2=6.94 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_8%A 3 7 9 12 13
r28 12 15 49.7087 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=6.815 $Y=1.49
+ $X2=6.815 $Y2=1.675
r29 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.49
+ $X2=6.815 $Y2=1.325
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.815
+ $Y=1.49 $X2=6.815 $Y2=1.49
r31 9 13 4.50137 $w=4.63e-07 $l=1.75e-07 $layer=LI1_cond $X=6.882 $Y=1.665
+ $X2=6.882 $Y2=1.49
r32 7 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.725 $Y=2.155
+ $X2=6.725 $Y2=1.675
r33 3 14 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.725 $Y=0.875
+ $X2=6.725 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_8%VPWR 1 2 3 4 5 6 7 24 30 34 38 44 50 56 62
+ 65 66 67 68 70 71 72 81 86 95 104 105 108 111 114 117
r106 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r107 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 105 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r112 102 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.415 $Y2=3.33
r113 102 104 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 101 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r115 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r116 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r117 97 100 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r118 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 95 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=3.33
+ $X2=6.415 $Y2=3.33
r120 95 100 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=3.33 $X2=6
+ $Y2=3.33
r121 94 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 94 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r123 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r124 91 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.165 $Y=3.33
+ $X2=4 $Y2=3.33
r125 91 93 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.165 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 87 111 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.27 $Y=3.33
+ $X2=3.14 $Y2=3.33
r127 87 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.27 $Y=3.33
+ $X2=3.6 $Y2=3.33
r128 86 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=3.33
+ $X2=4 $Y2=3.33
r129 86 89 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.835 $Y=3.33
+ $X2=3.6 $Y2=3.33
r130 85 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 85 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r132 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 82 108 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.28 $Y2=3.33
r134 82 84 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 81 111 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=3.14 $Y2=3.33
r136 81 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=2.64 $Y2=3.33
r137 80 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r141 72 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r142 72 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r143 72 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r144 71 97 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.91 $Y=3.33
+ $X2=5.04 $Y2=3.33
r145 70 93 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.78 $Y=3.33
+ $X2=4.56 $Y2=3.33
r146 70 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.78 $Y=3.33
+ $X2=4.91 $Y2=3.33
r147 67 79 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.29 $Y=3.33 $X2=1.2
+ $Y2=3.33
r148 67 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.42 $Y2=3.33
r149 65 75 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.24 $Y2=3.33
r150 65 66 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.542 $Y2=3.33
r151 64 79 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.69 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 64 66 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.69 $Y=3.33
+ $X2=0.542 $Y2=3.33
r153 60 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.415 $Y2=3.33
r154 60 62 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.415 $Y2=2.475
r155 56 59 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=4.91 $Y=2.26
+ $X2=4.91 $Y2=2.94
r156 54 71 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=3.245
+ $X2=4.91 $Y2=3.33
r157 54 59 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=4.91 $Y=3.245
+ $X2=4.91 $Y2=2.94
r158 50 53 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4 $Y=2.23 $X2=4
+ $Y2=2.91
r159 48 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=3.245 $X2=4
+ $Y2=3.33
r160 48 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4 $Y=3.245 $X2=4
+ $Y2=2.91
r161 44 47 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.14 $Y=2.27
+ $X2=3.14 $Y2=2.95
r162 42 111 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=3.33
r163 42 47 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=2.95
r164 38 41 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=2.28 $Y=2.27
+ $X2=2.28 $Y2=2.95
r165 36 108 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=3.33
r166 36 41 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=2.95
r167 35 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.42 $Y2=3.33
r168 34 108 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.28 $Y2=3.33
r169 34 35 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.15 $Y=3.33 $X2=1.55
+ $Y2=3.33
r170 30 33 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.42 $Y=2.27
+ $X2=1.42 $Y2=2.95
r171 28 68 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=3.245
+ $X2=1.42 $Y2=3.33
r172 28 33 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.42 $Y=3.245
+ $X2=1.42 $Y2=2.95
r173 24 27 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.542 $Y=2.27
+ $X2=0.542 $Y2=2.95
r174 22 66 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.542 $Y=3.245
+ $X2=0.542 $Y2=3.33
r175 22 27 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.542 $Y=3.245
+ $X2=0.542 $Y2=2.95
r176 7 62 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.835 $X2=6.415 $Y2=2.475
r177 6 59 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.835 $X2=4.905 $Y2=2.94
r178 6 56 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.835 $X2=4.905 $Y2=2.26
r179 5 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.835 $X2=4 $Y2=2.91
r180 5 50 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.835 $X2=4 $Y2=2.23
r181 4 47 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3
+ $Y=1.835 $X2=3.14 $Y2=2.95
r182 4 44 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=3
+ $Y=1.835 $X2=3.14 $Y2=2.27
r183 3 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.835 $X2=2.28 $Y2=2.95
r184 3 38 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.835 $X2=2.28 $Y2=2.27
r185 2 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=1.835 $X2=1.42 $Y2=2.95
r186 2 30 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=1.835 $X2=1.42 $Y2=2.27
r187 1 27 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.415
+ $Y=1.835 $X2=0.56 $Y2=2.95
r188 1 24 400 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=0.415
+ $Y=1.835 $X2=0.56 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_8%X 1 2 3 4 5 6 7 8 25 27 28 31 37 39 41 45
+ 51 53 55 59 65 67 69 73 79 82 83 84 85 86 87 88 89 93 95
r110 93 95 2.52097 $w=3.18e-07 $l=7e-08 $layer=LI1_cond $X=0.245 $Y=1.225
+ $X2=0.245 $Y2=1.295
r111 88 93 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.14
+ $X2=0.245 $Y2=1.225
r112 88 89 13.073 $w=3.18e-07 $l=3.63e-07 $layer=LI1_cond $X=0.245 $Y=1.302
+ $X2=0.245 $Y2=1.665
r113 88 95 0.252097 $w=3.18e-07 $l=7e-09 $layer=LI1_cond $X=0.245 $Y=1.302
+ $X2=0.245 $Y2=1.295
r114 81 89 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=0.245 $Y=1.755
+ $X2=0.245 $Y2=1.665
r115 77 79 35.0239 $w=1.88e-07 $l=6e-07 $layer=LI1_cond $X=3.57 $Y=1.055
+ $X2=3.57 $Y2=0.455
r116 73 75 40.4636 $w=2.23e-07 $l=7.9e-07 $layer=LI1_cond $X=3.552 $Y=2.05
+ $X2=3.552 $Y2=2.84
r117 71 73 6.40246 $w=2.23e-07 $l=1.25e-07 $layer=LI1_cond $X=3.552 $Y=1.925
+ $X2=3.552 $Y2=2.05
r118 70 86 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.84 $Y=1.84
+ $X2=2.71 $Y2=1.84
r119 69 71 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.44 $Y=1.84
+ $X2=3.552 $Y2=1.925
r120 69 70 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.44 $Y=1.84 $X2=2.84
+ $Y2=1.84
r121 68 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.805 $Y=1.14
+ $X2=2.71 $Y2=1.14
r122 67 77 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.475 $Y=1.14
+ $X2=3.57 $Y2=1.055
r123 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.475 $Y=1.14
+ $X2=2.805 $Y2=1.14
r124 63 87 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=1.055
+ $X2=2.71 $Y2=1.14
r125 63 65 35.0239 $w=1.88e-07 $l=6e-07 $layer=LI1_cond $X=2.71 $Y=1.055
+ $X2=2.71 $Y2=0.455
r126 59 61 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=2.71 $Y=2.05
+ $X2=2.71 $Y2=2.84
r127 57 86 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=1.925
+ $X2=2.71 $Y2=1.84
r128 57 59 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=2.71 $Y=1.925
+ $X2=2.71 $Y2=2.05
r129 56 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.98 $Y=1.84
+ $X2=1.85 $Y2=1.84
r130 55 86 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.58 $Y=1.84
+ $X2=2.71 $Y2=1.84
r131 55 56 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.58 $Y=1.84 $X2=1.98
+ $Y2=1.84
r132 54 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.945 $Y=1.14
+ $X2=1.85 $Y2=1.14
r133 53 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.615 $Y=1.14
+ $X2=2.71 $Y2=1.14
r134 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.615 $Y=1.14
+ $X2=1.945 $Y2=1.14
r135 49 85 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.85 $Y=1.055
+ $X2=1.85 $Y2=1.14
r136 49 51 35.0239 $w=1.88e-07 $l=6e-07 $layer=LI1_cond $X=1.85 $Y=1.055
+ $X2=1.85 $Y2=0.455
r137 45 47 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=1.85 $Y=2.05
+ $X2=1.85 $Y2=2.84
r138 43 84 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.85 $Y=1.925
+ $X2=1.85 $Y2=1.84
r139 43 45 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=1.85 $Y=1.925
+ $X2=1.85 $Y2=2.05
r140 42 82 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.12 $Y=1.84
+ $X2=0.99 $Y2=1.84
r141 41 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.72 $Y=1.84
+ $X2=1.85 $Y2=1.84
r142 41 42 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.72 $Y=1.84 $X2=1.12
+ $Y2=1.84
r143 40 83 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.085 $Y=1.14
+ $X2=0.99 $Y2=1.14
r144 39 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.755 $Y=1.14
+ $X2=1.85 $Y2=1.14
r145 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.755 $Y=1.14
+ $X2=1.085 $Y2=1.14
r146 35 83 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=1.055
+ $X2=0.99 $Y2=1.14
r147 35 37 35.0239 $w=1.88e-07 $l=6e-07 $layer=LI1_cond $X=0.99 $Y=1.055
+ $X2=0.99 $Y2=0.455
r148 31 33 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=0.99 $Y=2.05
+ $X2=0.99 $Y2=2.84
r149 29 82 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=1.925
+ $X2=0.99 $Y2=1.84
r150 29 31 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.99 $Y=1.925
+ $X2=0.99 $Y2=2.05
r151 28 81 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=0.405 $Y=1.84
+ $X2=0.245 $Y2=1.755
r152 27 82 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.86 $Y=1.84
+ $X2=0.99 $Y2=1.84
r153 27 28 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=0.86 $Y=1.84
+ $X2=0.405 $Y2=1.84
r154 26 88 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.405 $Y=1.14
+ $X2=0.245 $Y2=1.14
r155 25 83 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.895 $Y=1.14
+ $X2=0.99 $Y2=1.14
r156 25 26 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=0.895 $Y=1.14
+ $X2=0.405 $Y2=1.14
r157 8 75 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.835 $X2=3.57 $Y2=2.84
r158 8 73 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.835 $X2=3.57 $Y2=2.05
r159 7 61 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.835 $X2=2.71 $Y2=2.84
r160 7 59 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.835 $X2=2.71 $Y2=2.05
r161 6 47 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.835 $X2=1.85 $Y2=2.84
r162 6 45 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.835 $X2=1.85 $Y2=2.05
r163 5 33 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=0.85
+ $Y=1.835 $X2=0.99 $Y2=2.84
r164 5 31 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=0.85
+ $Y=1.835 $X2=0.99 $Y2=2.05
r165 4 79 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.245 $X2=3.57 $Y2=0.455
r166 3 65 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.245 $X2=2.71 $Y2=0.455
r167 2 51 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=1.71
+ $Y=0.245 $X2=1.85 $Y2=0.455
r168 1 37 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=0.85
+ $Y=0.245 $X2=0.99 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__BUFBUF_8%VGND 1 2 3 4 5 6 7 24 28 30 34 38 42 46 50
+ 55 56 57 58 60 61 62 71 76 81 91 92 95 98 101 104
r118 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r119 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r120 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r121 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r122 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r123 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r124 89 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r125 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r126 86 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=0
+ $X2=4.905 $Y2=0
r127 86 88 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=5.07 $Y=0 $X2=6
+ $Y2=0
r128 85 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r129 85 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r130 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r131 82 101 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=4.19 $Y=0
+ $X2=4.012 $Y2=0
r132 82 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.56
+ $Y2=0
r133 81 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=0
+ $X2=4.905 $Y2=0
r134 81 84 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.56
+ $Y2=0
r135 77 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.14
+ $Y2=0
r136 77 79 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.6
+ $Y2=0
r137 76 101 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.835 $Y=0
+ $X2=4.012 $Y2=0
r138 76 79 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.835 $Y=0 $X2=3.6
+ $Y2=0
r139 75 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r140 75 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r141 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r142 72 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r143 72 74 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.64 $Y2=0
r144 71 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.14
+ $Y2=0
r145 71 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=2.64 $Y2=0
r146 70 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r147 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r148 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r149 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r150 62 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r151 62 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r152 62 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r153 60 88 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.21 $Y=0 $X2=6
+ $Y2=0
r154 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.21 $Y=0 $X2=6.375
+ $Y2=0
r155 59 91 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6.54 $Y=0 $X2=6.96
+ $Y2=0
r156 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.54 $Y=0 $X2=6.375
+ $Y2=0
r157 57 69 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.2
+ $Y2=0
r158 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.42
+ $Y2=0
r159 55 65 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.24 $Y2=0
r160 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.56
+ $Y2=0
r161 54 69 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=1.2
+ $Y2=0
r162 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.56
+ $Y2=0
r163 50 52 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=6.375 $Y=0.39
+ $X2=6.375 $Y2=0.785
r164 48 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0
r165 48 50 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0.39
r166 44 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=0.085
+ $X2=4.905 $Y2=0
r167 44 46 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.905 $Y=0.085
+ $X2=4.905 $Y2=0.415
r168 40 101 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.012 $Y=0.085
+ $X2=4.012 $Y2=0
r169 40 42 10.7129 $w=3.53e-07 $l=3.3e-07 $layer=LI1_cond $X=4.012 $Y=0.085
+ $X2=4.012 $Y2=0.415
r170 36 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r171 36 38 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.415
r172 32 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r173 32 34 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.415
r174 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.42
+ $Y2=0
r175 30 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r176 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=1.585 $Y2=0
r177 26 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=0.085
+ $X2=1.42 $Y2=0
r178 26 28 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.42 $Y=0.085
+ $X2=1.42 $Y2=0.415
r179 22 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0
r180 22 24 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0.415
r181 7 52 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.245 $X2=6.375 $Y2=0.785
r182 7 50 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.245 $X2=6.375 $Y2=0.39
r183 6 46 91 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=2 $X=4.765
+ $Y=0.245 $X2=4.905 $Y2=0.415
r184 5 42 91 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.245 $X2=4.025 $Y2=0.415
r185 4 38 91 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=2 $X=3
+ $Y=0.245 $X2=3.14 $Y2=0.415
r186 3 34 91 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=2 $X=2.14
+ $Y=0.245 $X2=2.28 $Y2=0.415
r187 2 28 91 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=2 $X=1.28
+ $Y=0.245 $X2=1.42 $Y2=0.415
r188 1 24 91 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=2 $X=0.435
+ $Y=0.245 $X2=0.56 $Y2=0.415
.ends

