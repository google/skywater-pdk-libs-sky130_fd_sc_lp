* File: sky130_fd_sc_lp__o311ai_2.spice
* Created: Wed Sep  2 10:23:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311ai_2.pex.spice"
.subckt sky130_fd_sc_lp__o311ai_2  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A1_M1018_g N_A_35_47#_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1018_d N_A1_M1019_g N_A_35_47#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_35_47#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1006_d N_A2_M1017_g N_A_35_47#_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.136 M=1 R=5.6 SA=75001.5
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1002 N_A_35_47#_M1017_s N_A3_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.2604 PD=1.16 PS=1.46 NRD=3.564 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1014 N_A_35_47#_M1014_d N_A3_M1014_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75002.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1000 N_A_35_47#_M1014_d N_B1_M1000_g N_A_710_47#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_35_47#_M1009_d N_B1_M1009_g N_A_710_47#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_710_47#_M1008_d N_C1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_A_710_47#_M1008_d N_C1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_35_367#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1004_d N_A1_M1012_g N_A_35_367#_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_A_290_367#_M1003_d N_A2_M1003_g N_A_35_367#_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_290_367#_M1003_d N_A2_M1015_g N_A_35_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_290_367#_M1005_d N_A3_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1016 N_A_290_367#_M1005_d N_A3_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1016_s N_B1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4158 PD=1.54 PS=1.92 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1013 N_Y_M1013_d N_B1_M1013_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4158 PD=1.54 PS=1.92 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_C1_M1001_g N_Y_M1013_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1001_d N_C1_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__o311ai_2.pxi.spice"
*
.ends
*
*
