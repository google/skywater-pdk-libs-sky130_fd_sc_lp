* File: sky130_fd_sc_lp__ha_m.pex.spice
* Created: Wed Sep  2 09:54:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__HA_M%A_80_60# 1 2 9 12 13 14 17 21 22 24 25 27 28 31
+ 32 34 39 41
r81 36 39 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.06 $Y=0.51
+ $X2=1.215 $Y2=0.51
r82 32 34 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=1.85 $Y=2.465
+ $X2=1.96 $Y2=2.465
r83 31 32 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.765 $Y=2.36
+ $X2=1.85 $Y2=2.465
r84 30 31 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.765 $Y=2.12
+ $X2=1.765 $Y2=2.36
r85 29 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.035
+ $X2=1.06 $Y2=2.035
r86 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.765 $Y2=2.12
r87 28 29 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.145 $Y2=2.035
r88 27 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=1.95 $X2=1.06
+ $Y2=2.035
r89 26 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0.675
+ $X2=1.06 $Y2=0.51
r90 26 27 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=1.06 $Y=0.675
+ $X2=1.06 $Y2=1.95
r91 24 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=2.035
+ $X2=1.06 $Y2=2.035
r92 24 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.975 $Y=2.035
+ $X2=0.775 $Y2=2.035
r93 22 43 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.627 $Y=1.615
+ $X2=0.627 $Y2=1.45
r94 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.615 $X2=0.69 $Y2=1.615
r95 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=1.95
+ $X2=0.775 $Y2=2.035
r96 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=1.95
+ $X2=0.69 $Y2=1.615
r97 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.14 $Y=2.12
+ $X2=1.14 $Y2=2.53
r98 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.065 $Y=2.045
+ $X2=1.14 $Y2=2.12
r99 13 14 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.065 $Y=2.045
+ $X2=0.855 $Y2=2.045
r100 12 14 36.9868 $w=1.5e-07 $l=2.62838e-07 $layer=POLY_cond $X=0.627 $Y=1.97
+ $X2=0.855 $Y2=2.045
r101 11 22 7.57836 $w=4.55e-07 $l=6.2e-08 $layer=POLY_cond $X=0.627 $Y=1.677
+ $X2=0.627 $Y2=1.615
r102 11 12 35.8139 $w=4.55e-07 $l=2.93e-07 $layer=POLY_cond $X=0.627 $Y=1.677
+ $X2=0.627 $Y2=1.97
r103 9 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.475 $Y=0.64
+ $X2=0.475 $Y2=1.45
r104 2 34 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=2.32 $X2=1.96 $Y2=2.465
r105 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.215 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%A_249_212# 1 2 9 12 15 17 21 24 27 28 31 35 36
+ 38 39 41 43 46 53 54 59
c120 38 0 1.70003e-19 $X=2.61 $Y=1.645
c121 31 0 9.8052e-20 $X=1.745 $Y=2.11
r122 52 54 15.1258 $w=3.18e-07 $l=4.2e-07 $layer=LI1_cond $X=3.215 $Y=0.955
+ $X2=3.635 $Y2=0.955
r123 52 53 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=0.955
+ $X2=3.05 $Y2=0.955
r124 49 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.635 $Y=2.94
+ $X2=3.8 $Y2=2.94
r125 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.635
+ $Y=2.94 $X2=3.635 $Y2=2.94
r126 46 48 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=3.635 $Y=2.29
+ $X2=3.635 $Y2=2.94
r127 44 54 0.527965 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=3.635 $Y=1.115
+ $X2=3.635 $Y2=0.955
r128 44 46 41.034 $w=3.28e-07 $l=1.175e-06 $layer=LI1_cond $X=3.635 $Y=1.115
+ $X2=3.635 $Y2=2.29
r129 43 53 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.78 $Y=1.03
+ $X2=3.05 $Y2=1.03
r130 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.695 $Y=1.115
+ $X2=2.78 $Y2=1.03
r131 40 41 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.695 $Y=1.115
+ $X2=2.695 $Y2=1.56
r132 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=1.645
+ $X2=2.695 $Y2=1.56
r133 38 39 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.61 $Y=1.645
+ $X2=1.495 $Y2=1.645
r134 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.41
+ $Y=1.225 $X2=1.41 $Y2=1.225
r135 33 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.41 $Y=1.56
+ $X2=1.495 $Y2=1.645
r136 33 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.41 $Y=1.56
+ $X2=1.41 $Y2=1.225
r137 29 31 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.5 $Y=2.11
+ $X2=1.745 $Y2=2.11
r138 27 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.41 $Y=1.565
+ $X2=1.41 $Y2=1.225
r139 27 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.565
+ $X2=1.41 $Y2=1.73
r140 26 36 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.06
+ $X2=1.41 $Y2=1.225
r141 21 24 712.745 $w=1.5e-07 $l=1.39e-06 $layer=POLY_cond $X=4.315 $Y=0.835
+ $X2=4.315 $Y2=2.225
r142 19 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.315 $Y=2.805
+ $X2=4.315 $Y2=2.225
r143 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.24 $Y=2.88
+ $X2=4.315 $Y2=2.805
r144 17 59 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.24 $Y=2.88
+ $X2=3.8 $Y2=2.88
r145 13 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.745 $Y=2.185
+ $X2=1.745 $Y2=2.11
r146 13 15 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.745 $Y=2.185
+ $X2=1.745 $Y2=2.53
r147 12 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.5 $Y=2.035
+ $X2=1.5 $Y2=2.11
r148 12 28 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.5 $Y=2.035
+ $X2=1.5 $Y2=1.73
r149 9 26 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.43 $Y=0.445
+ $X2=1.43 $Y2=1.06
r150 2 46 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.015 $X2=3.575 $Y2=2.29
r151 1 52 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.625 $X2=3.215 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%B 3 5 7 9 11 14 17 20 22 23 24 29 31 34
c81 29 0 1.9418e-19 $X=3.125 $Y=1.91
c82 24 0 9.8052e-20 $X=2.96 $Y=2.015
r83 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.38 $X2=3.125 $Y2=1.38
r84 29 34 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=3.125 $Y=1.91
+ $X2=3.125 $Y2=2.015
r85 29 31 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.125 $Y=1.91
+ $X2=3.125 $Y2=1.38
r86 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.195
+ $Y=1.995 $X2=2.195 $Y2=1.995
r87 24 34 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=2.015
+ $X2=3.125 $Y2=2.015
r88 24 26 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=2.96 $Y=2.015
+ $X2=2.195 $Y2=2.015
r89 22 32 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.45 $Y=1.38
+ $X2=3.125 $Y2=1.38
r90 22 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.45 $Y=1.38
+ $X2=3.525 $Y2=1.38
r91 18 20 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.265 $Y=1.83
+ $X2=3.525 $Y2=1.83
r92 17 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.525 $Y=1.755
+ $X2=3.525 $Y2=1.83
r93 16 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.545
+ $X2=3.525 $Y2=1.38
r94 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.525 $Y=1.545
+ $X2=3.525 $Y2=1.755
r95 12 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.215
+ $X2=3.525 $Y2=1.38
r96 12 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=3.525 $Y=1.215
+ $X2=3.525 $Y2=0.835
r97 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.905
+ $X2=3.265 $Y2=1.83
r98 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.265 $Y=1.905
+ $X2=3.265 $Y2=2.225
r99 5 27 38.6446 $w=3.36e-07 $l=2.10286e-07 $layer=POLY_cond $X=2.175 $Y=2.16
+ $X2=2.072 $Y2=1.995
r100 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.175 $Y=2.16
+ $X2=2.175 $Y2=2.53
r101 1 27 65.1833 $w=3.36e-07 $l=4.43509e-07 $layer=POLY_cond $X=1.86 $Y=1.645
+ $X2=2.072 $Y2=1.995
r102 1 3 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=1.86 $Y=1.645
+ $X2=1.86 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%A 1 3 4 6 8 11 12 13 16 18 20 25
c67 4 0 2.97734e-19 $X=2.865 $Y=0.84
r68 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.345
+ $Y=1.215 $X2=2.345 $Y2=1.215
r69 20 25 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.16 $Y=1.215
+ $X2=2.345 $Y2=1.215
r70 16 18 712.745 $w=1.5e-07 $l=1.39e-06 $layer=POLY_cond $X=3.885 $Y=0.835
+ $X2=3.885 $Y2=2.225
r71 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.885 $Y=0.255
+ $X2=3.885 $Y2=0.835
r72 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.81 $Y=0.18
+ $X2=3.885 $Y2=0.255
r73 12 13 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=3.81 $Y=0.18
+ $X2=3.015 $Y2=0.18
r74 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.94 $Y=0.255
+ $X2=3.015 $Y2=0.18
r75 10 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.94 $Y=0.255
+ $X2=2.94 $Y2=0.765
r76 6 24 42.5185 $w=3.03e-07 $l=2.73998e-07 $layer=POLY_cond $X=2.645 $Y=1.405
+ $X2=2.45 $Y2=1.215
r77 6 8 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.645 $Y=1.405
+ $X2=2.645 $Y2=2.53
r78 5 24 59.6535 $w=3.03e-07 $l=3.75e-07 $layer=POLY_cond $X=2.45 $Y=0.84
+ $X2=2.45 $Y2=1.215
r79 4 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.865 $Y=0.84
+ $X2=2.94 $Y2=0.765
r80 4 5 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.865 $Y=0.84 $X2=2.525
+ $Y2=0.84
r81 1 5 24.2248 $w=3.03e-07 $l=7.5e-08 $layer=POLY_cond $X=2.45 $Y=0.765
+ $X2=2.45 $Y2=0.84
r82 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.45 $Y=0.765 $X2=2.45
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%SUM 1 2 9 11 12 13 14 15 16 17
r25 16 17 3.88743 $w=5e-07 $l=1.94743e-07 $layer=LI1_cond $X=0.24 $Y=2.49
+ $X2=0.26 $Y2=2.675
r26 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.035
+ $X2=0.26 $Y2=2.405
r27 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r28 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r29 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.925
+ $X2=0.26 $Y2=1.295
r30 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.555
+ $X2=0.26 $Y2=0.925
r31 7 17 3.1289 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.675
+ $X2=0.26 $Y2=2.675
r32 7 9 15.5736 $w=3.68e-07 $l=5e-07 $layer=LI1_cond $X=0.425 $Y=2.675 $X2=0.925
+ $Y2=2.675
r33 2 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.8
+ $Y=2.32 $X2=0.925 $Y2=2.595
r34 1 11 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.43 $X2=0.26 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%VPWR 1 2 3 12 16 20 23 24 26 27 28 43 49 50 53
r60 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 50 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r63 47 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.09 $Y2=3.33
r64 47 49 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r65 46 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r67 43 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.995 $Y=3.33
+ $X2=4.09 $Y2=3.33
r68 43 45 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.995 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 42 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r70 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r72 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 36 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r75 32 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 31 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r77 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r78 28 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r79 28 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r80 26 41 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=3.33 $X2=2.64
+ $Y2=3.33
r81 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=3.33
+ $X2=2.955 $Y2=3.33
r82 25 45 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=3.6
+ $Y2=3.33
r83 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.955 $Y2=3.33
r84 23 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.27 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.375 $Y2=3.33
r86 22 38 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.48 $Y=3.33 $X2=1.68
+ $Y2=3.33
r87 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.48 $Y=3.33
+ $X2=1.375 $Y2=3.33
r88 18 53 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=3.245
+ $X2=4.09 $Y2=3.33
r89 18 20 55.7464 $w=1.88e-07 $l=9.55e-07 $layer=LI1_cond $X=4.09 $Y=3.245
+ $X2=4.09 $Y2=2.29
r90 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=3.33
r91 14 16 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=2.595
r92 10 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=3.245
+ $X2=1.375 $Y2=3.33
r93 10 12 34.329 $w=2.08e-07 $l=6.5e-07 $layer=LI1_cond $X=1.375 $Y=3.245
+ $X2=1.375 $Y2=2.595
r94 3 20 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=2.015 $X2=4.1 $Y2=2.29
r95 2 16 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=2.32 $X2=2.955 $Y2=2.595
r96 1 12 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=2.32 $X2=1.375 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%COUT 1 2 7 8 9 10 11 12 13
r12 12 13 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=4.535 $Y=2.405
+ $X2=4.535 $Y2=2.775
r13 12 35 12.834 $w=2.18e-07 $l=2.45e-07 $layer=LI1_cond $X=4.535 $Y=2.405
+ $X2=4.535 $Y2=2.16
r14 11 35 6.54797 $w=2.18e-07 $l=1.25e-07 $layer=LI1_cond $X=4.535 $Y=2.035
+ $X2=4.535 $Y2=2.16
r15 10 11 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=4.535 $Y=1.665
+ $X2=4.535 $Y2=2.035
r16 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=4.535 $Y=1.295
+ $X2=4.535 $Y2=1.665
r17 8 9 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=4.535 $Y=0.925
+ $X2=4.535 $Y2=1.295
r18 8 25 8.11948 $w=2.18e-07 $l=1.55e-07 $layer=LI1_cond $X=4.535 $Y=0.925
+ $X2=4.535 $Y2=0.77
r19 7 25 11.2625 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=4.535 $Y=0.555
+ $X2=4.535 $Y2=0.77
r20 2 35 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=2.015 $X2=4.53 $Y2=2.16
r21 1 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.625 $X2=4.53 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%VGND 1 2 3 12 16 18 20 25 30 40 41 44 48 54
c53 41 0 1.27732e-19 $X=4.56 $Y=0
r54 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r55 48 51 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=2.155
+ $Y2=0.33
r56 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r57 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r59 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r60 38 54 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.09
+ $Y2=0
r61 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.56
+ $Y2=0
r62 37 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r63 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r64 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r65 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r66 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r67 31 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.155
+ $Y2=0
r68 31 33 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.64
+ $Y2=0
r69 30 54 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.09
+ $Y2=0
r70 30 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.6
+ $Y2=0
r71 29 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r72 29 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r73 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 26 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.7
+ $Y2=0
r75 26 28 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.68
+ $Y2=0
r76 25 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=0 $X2=2.155
+ $Y2=0
r77 25 28 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.99 $Y=0 $X2=1.68
+ $Y2=0
r78 23 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r79 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r80 20 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.7
+ $Y2=0
r81 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r82 18 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r83 18 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r84 14 54 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0
r85 14 16 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0.77
r86 10 44 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r87 10 12 28.6029 $w=1.88e-07 $l=4.9e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.575
r88 3 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.96
+ $Y=0.625 $X2=4.1 $Y2=0.77
r89 2 51 182 $w=1.7e-07 $l=2.63249e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.235 $X2=2.155 $Y2=0.33
r90 1 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.43 $X2=0.69 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__HA_M%A_301_47# 1 2 7 10 15
r28 15 17 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=2.665 $Y=0.51
+ $X2=2.665 $Y2=0.68
r29 10 12 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=1.645 $Y=0.51
+ $X2=1.645 $Y2=0.68
r30 8 12 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.75 $Y=0.68 $X2=1.645
+ $Y2=0.68
r31 7 17 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.56 $Y=0.68 $X2=2.665
+ $Y2=0.68
r32 7 8 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.56 $Y=0.68 $X2=1.75
+ $Y2=0.68
r33 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.665 $Y2=0.51
r34 1 10 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.645 $Y2=0.51
.ends

