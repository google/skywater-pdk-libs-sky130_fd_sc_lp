# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxbp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxbp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.570000 1.180000 0.900000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.585900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.560000 0.265000 6.890000 0.925000 ;
        RECT 6.560000 0.925000 8.035000 1.095000 ;
        RECT 6.635000 1.785000 8.035000 1.955000 ;
        RECT 6.635000 1.955000 6.965000 3.065000 ;
        RECT 7.805000 1.095000 8.035000 1.785000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.579600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.635000 0.265000 9.980000 3.065000 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.525000 1.390000 2.195000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 0.905000  0.085000  1.155000 0.995000 ;
        RECT 3.145000  0.085000  3.475000 0.645000 ;
        RECT 5.210000  0.085000  5.540000 1.095000 ;
        RECT 7.350000  0.085000  7.680000 0.745000 ;
        RECT 8.845000  0.085000  9.175000 1.125000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 0.895000 2.735000  1.225000 3.245000 ;
        RECT 3.250000 2.375000  3.580000 3.245000 ;
        RECT 5.305000 2.545000  5.635000 3.245000 ;
        RECT 7.425000 2.135000  7.755000 3.245000 ;
        RECT 8.860000 1.815000  9.190000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105000 0.535000 0.445000 0.995000 ;
      RECT 0.105000 0.995000 0.275000 2.385000 ;
      RECT 0.105000 2.385000 1.575000 2.555000 ;
      RECT 0.105000 2.555000 0.435000 3.065000 ;
      RECT 1.375000 0.265000 2.655000 0.435000 ;
      RECT 1.375000 0.435000 1.545000 1.175000 ;
      RECT 1.375000 1.175000 1.740000 1.345000 ;
      RECT 1.405000 2.555000 1.575000 2.895000 ;
      RECT 1.405000 2.895000 3.070000 3.065000 ;
      RECT 1.570000 1.345000 1.740000 2.035000 ;
      RECT 1.570000 2.035000 2.710000 2.205000 ;
      RECT 1.725000 0.615000 2.090000 0.995000 ;
      RECT 1.920000 0.995000 2.090000 1.525000 ;
      RECT 1.920000 1.525000 2.960000 1.845000 ;
      RECT 1.920000 1.845000 2.170000 1.855000 ;
      RECT 2.325000 0.435000 2.655000 0.825000 ;
      RECT 2.325000 0.825000 4.140000 0.995000 ;
      RECT 2.380000 2.205000 2.710000 2.715000 ;
      RECT 2.630000 1.175000 2.960000 1.335000 ;
      RECT 2.630000 1.335000 4.520000 1.505000 ;
      RECT 2.630000 1.505000 2.960000 1.525000 ;
      RECT 2.900000 2.025000 3.735000 2.195000 ;
      RECT 2.900000 2.195000 3.070000 2.895000 ;
      RECT 3.405000 1.865000 3.735000 2.025000 ;
      RECT 3.810000 0.995000 4.140000 1.155000 ;
      RECT 3.945000 1.505000 4.275000 2.165000 ;
      RECT 4.045000 0.295000 5.030000 0.645000 ;
      RECT 4.070000 2.575000 4.625000 2.745000 ;
      RECT 4.070000 2.745000 4.400000 3.035000 ;
      RECT 4.350000 0.825000 4.680000 1.155000 ;
      RECT 4.350000 1.155000 4.520000 1.335000 ;
      RECT 4.455000 1.685000 5.030000 1.855000 ;
      RECT 4.455000 1.855000 4.625000 2.575000 ;
      RECT 4.845000 2.035000 6.425000 2.365000 ;
      RECT 4.860000 0.645000 5.030000 1.275000 ;
      RECT 4.860000 1.275000 5.970000 1.605000 ;
      RECT 4.860000 1.605000 5.030000 1.685000 ;
      RECT 6.000000 0.265000 6.330000 1.095000 ;
      RECT 6.095000 1.785000 6.425000 2.035000 ;
      RECT 6.095000 2.365000 6.425000 3.065000 ;
      RECT 6.160000 1.095000 6.330000 1.275000 ;
      RECT 6.160000 1.275000 7.625000 1.605000 ;
      RECT 6.160000 1.605000 6.425000 1.785000 ;
      RECT 8.285000 0.635000 8.615000 1.305000 ;
      RECT 8.285000 1.305000 9.455000 1.635000 ;
      RECT 8.285000 1.635000 8.650000 2.465000 ;
  END
END sky130_fd_sc_lp__dlxbp_lp
