* File: sky130_fd_sc_lp__o311a_m.pex.spice
* Created: Fri Aug 28 11:14:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311A_M%A1 2 7 11 12 13 14 15 16 17 22 24
r44 22 24 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.032 $Y=1.32
+ $X2=1.032 $Y2=1.155
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.02
+ $Y=1.32 $X2=1.02 $Y2=1.32
r46 17 23 8.77972 $w=4.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.87 $Y=1.665
+ $X2=0.87 $Y2=1.32
r47 16 23 0.636212 $w=4.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=1.32
r48 15 16 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.87 $Y=0.925
+ $X2=0.87 $Y2=1.295
r49 14 24 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.135 $Y=0.915
+ $X2=1.135 $Y2=1.155
r50 13 14 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.155 $Y=0.765
+ $X2=1.155 $Y2=0.915
r51 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.175 $Y=0.445
+ $X2=1.175 $Y2=0.765
r52 7 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.135 $Y=2.195
+ $X2=1.135 $Y2=1.825
r53 2 12 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=1.032 $Y=1.648
+ $X2=1.032 $Y2=1.825
r54 1 22 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=1.032 $Y=1.332
+ $X2=1.032 $Y2=1.32
r55 1 2 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=1.032 $Y=1.332
+ $X2=1.032 $Y2=1.648
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%A2 3 7 11 12 13 14 15 16 22
c42 11 0 1.4009e-19 $X=1.585 $Y=1.66
r43 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.585
+ $Y=1.32 $X2=1.585 $Y2=1.32
r44 15 16 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.632 $Y=2.035
+ $X2=1.632 $Y2=2.405
r45 14 15 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.632 $Y=1.665
+ $X2=1.632 $Y2=2.035
r46 14 23 15.0035 $w=2.63e-07 $l=3.45e-07 $layer=LI1_cond $X=1.632 $Y=1.665
+ $X2=1.632 $Y2=1.32
r47 13 23 1.08721 $w=2.63e-07 $l=2.5e-08 $layer=LI1_cond $X=1.632 $Y=1.295
+ $X2=1.632 $Y2=1.32
r48 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.585 $Y=1.66
+ $X2=1.585 $Y2=1.32
r49 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.66
+ $X2=1.585 $Y2=1.825
r50 10 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.155
+ $X2=1.585 $Y2=1.32
r51 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.605 $Y=0.445
+ $X2=1.605 $Y2=1.155
r52 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.495 $Y=2.195
+ $X2=1.495 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%A_93_153# 1 2 3 13 14 15 16 18 21 26 27 28
+ 31 34 36 37 40 44
c87 16 0 1.1261e-19 $X=0.745 $Y=0.765
r88 41 44 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=3.22 $Y=0.51
+ $X2=3.33 $Y2=0.51
r89 37 48 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.19 $Y=2.94 $X2=2.19
+ $Y2=3.03
r90 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=2.94 $X2=2.19 $Y2=2.94
r91 34 40 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=3.22 $Y=1.765
+ $X2=3.21 $Y2=1.85
r92 33 41 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.22 $Y=0.615
+ $X2=3.22 $Y2=0.51
r93 33 34 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=3.22 $Y=0.615
+ $X2=3.22 $Y2=1.765
r94 29 40 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=1.935
+ $X2=3.21 $Y2=1.85
r95 29 31 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=3.21 $Y=1.935
+ $X2=3.21 $Y2=2.11
r96 27 40 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.115 $Y=1.85
+ $X2=3.21 $Y2=1.85
r97 27 28 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.115 $Y=1.85
+ $X2=2.355 $Y2=1.85
r98 26 36 38.29 $w=2.08e-07 $l=7.25e-07 $layer=LI1_cond $X=2.25 $Y=2.13 $X2=2.25
+ $Y2=2.855
r99 23 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.25 $Y=1.935
+ $X2=2.355 $Y2=1.85
r100 23 26 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=2.25 $Y=1.935
+ $X2=2.25 $Y2=2.13
r101 19 21 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.54 $Y=0.84
+ $X2=0.745 $Y2=0.84
r102 16 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.745 $Y=0.765
+ $X2=0.745 $Y2=0.84
r103 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.745 $Y=0.765
+ $X2=0.745 $Y2=0.445
r104 14 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.025 $Y=3.03
+ $X2=2.19 $Y2=3.03
r105 14 15 723 $w=1.5e-07 $l=1.41e-06 $layer=POLY_cond $X=2.025 $Y=3.03
+ $X2=0.615 $Y2=3.03
r106 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.54 $Y=2.955
+ $X2=0.615 $Y2=3.03
r107 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.54 $Y=2.955
+ $X2=0.54 $Y2=2.195
r108 10 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.54 $Y=0.915
+ $X2=0.54 $Y2=0.84
r109 10 13 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=0.54 $Y=0.915
+ $X2=0.54 $Y2=2.195
r110 3 31 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.985 $X2=3.22 $Y2=2.11
r111 2 26 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=1.985 $X2=2.25 $Y2=2.13
r112 1 44 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.235 $X2=3.33 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%A3 3 7 11 12 13 16 17
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.125
+ $Y=1.16 $X2=2.125 $Y2=1.16
r40 13 17 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.125 $Y=1.295
+ $X2=2.125 $Y2=1.16
r41 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.125 $Y=1.5
+ $X2=2.125 $Y2=1.16
r42 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.125 $Y=1.5
+ $X2=2.125 $Y2=1.665
r43 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.125 $Y=0.995
+ $X2=2.125 $Y2=1.16
r44 7 12 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.035 $Y=2.195
+ $X2=2.035 $Y2=1.665
r45 3 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.035 $Y=0.445
+ $X2=2.035 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%B1 3 7 11 12 13 14 18
r42 13 14 21.0443 $w=1.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.652 $Y=0.925
+ $X2=2.652 $Y2=1.295
r43 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.665
+ $Y=0.96 $X2=2.665 $Y2=0.96
r44 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.665 $Y=1.3
+ $X2=2.665 $Y2=0.96
r45 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.3
+ $X2=2.665 $Y2=1.465
r46 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=0.795
+ $X2=2.665 $Y2=0.96
r47 7 12 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.575 $Y=2.195
+ $X2=2.575 $Y2=1.465
r48 3 10 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.575 $Y=0.445
+ $X2=2.575 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%C1 3 7 9 10 11 12 14 17 18 19 20 21 22 29
r43 21 22 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.585 $Y=2.035
+ $X2=3.585 $Y2=2.405
r44 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.585 $Y=1.665
+ $X2=3.585 $Y2=2.035
r45 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.585 $Y=1.295
+ $X2=3.585 $Y2=1.665
r46 18 19 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.585 $Y=0.925
+ $X2=3.585 $Y2=1.295
r47 18 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.005 $X2=3.57 $Y2=1.005
r48 16 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.005
r49 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.51
r50 15 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.57 $Y=0.99
+ $X2=3.57 $Y2=1.005
r51 14 17 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.48 $Y=1.705
+ $X2=3.48 $Y2=1.51
r52 11 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.405 $Y=0.915
+ $X2=3.57 $Y2=0.99
r53 11 12 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.405 $Y=0.915
+ $X2=3.19 $Y2=0.915
r54 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.405 $Y=1.78
+ $X2=3.48 $Y2=1.705
r55 9 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.405 $Y=1.78
+ $X2=3.08 $Y2=1.78
r56 5 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.115 $Y=0.84
+ $X2=3.19 $Y2=0.915
r57 5 7 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.115 $Y=0.84
+ $X2=3.115 $Y2=0.445
r58 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.005 $Y=1.855
+ $X2=3.08 $Y2=1.78
r59 1 3 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.005 $Y=1.855
+ $X2=3.005 $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%X 1 2 10 11 13 19
c12 19 0 2.08402e-19 $X=0.53 $Y=0.495
r13 13 19 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.24 $Y=0.495
+ $X2=0.53 $Y2=0.495
r14 10 11 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.282 $Y=2.13
+ $X2=0.282 $Y2=1.965
r15 7 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.66 $X2=0.24
+ $Y2=0.495
r16 7 11 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=0.24 $Y=0.66
+ $X2=0.24 $Y2=1.965
r17 2 10 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.985 $X2=0.305 $Y2=2.13
r18 1 19 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=0.405
+ $Y=0.235 $X2=0.53 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%VPWR 1 2 9 13 16 17 18 20 33 34 37
r37 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=0.755 $Y2=3.33
r45 25 27 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.92 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.755 $Y2=3.33
r49 20 22 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 16 30 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.79 $Y2=3.33
r54 15 33 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.79 $Y2=3.33
r56 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=3.33
r57 11 13 50.9654 $w=2.08e-07 $l=9.65e-07 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=2.28
r58 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=3.245
+ $X2=0.755 $Y2=3.33
r59 7 9 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=0.755 $Y=3.245
+ $X2=0.755 $Y2=2.26
r60 2 13 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.985 $X2=2.79 $Y2=2.28
r61 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.985 $X2=0.755 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%VGND 1 2 9 13 16 17 19 20 21 34 35
r52 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r53 32 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r54 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r55 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r58 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r59 21 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r60 21 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r61 19 28 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.68
+ $Y2=0
r62 19 20 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.82
+ $Y2=0
r63 18 31 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=2.16
+ $Y2=0
r64 18 20 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=1.82
+ $Y2=0
r65 16 24 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.72
+ $Y2=0
r66 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.96
+ $Y2=0
r67 15 28 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.68
+ $Y2=0
r68 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.96
+ $Y2=0
r69 11 20 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.82 $Y=0.085
+ $X2=1.82 $Y2=0
r70 11 13 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.82 $Y=0.085
+ $X2=1.82 $Y2=0.38
r71 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0
r72 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0.38
r73 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.68
+ $Y=0.235 $X2=1.82 $Y2=0.38
r74 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.82
+ $Y=0.235 $X2=0.96 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_M%A_250_47# 1 2 9 11 12 15
c29 9 0 9.57924e-20 $X=1.39 $Y=0.51
r30 13 15 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.24 $Y=0.725
+ $X2=2.24 $Y2=0.51
r31 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.145 $Y=0.81
+ $X2=2.24 $Y2=0.725
r32 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.145 $Y=0.81
+ $X2=1.495 $Y2=0.81
r33 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.39 $Y=0.725
+ $X2=1.495 $Y2=0.81
r34 7 9 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.39 $Y=0.725 $X2=1.39
+ $Y2=0.51
r35 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.11
+ $Y=0.235 $X2=2.25 $Y2=0.51
r36 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.25
+ $Y=0.235 $X2=1.39 $Y2=0.51
.ends

