* NGSPICE file created from sky130_fd_sc_lp__dfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
M1000 a_628_119# a_236_463# a_537_119# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.281e+11p ps=1.45e+06u
M1001 a_537_119# a_110_70# a_429_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1002 a_110_70# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=2.5364e+12p ps=1.955e+07u
M1003 Q a_1169_93# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1004 VGND a_1169_93# a_1125_119# VNB nshort w=420000u l=150000u
+  ad=2.0153e+12p pd=1.608e+07u as=9.24e+10p ps=1.28e+06u
M1005 a_1169_93# a_982_369# VGND VNB nshort w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1006 VGND a_670_93# a_628_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_670_93# a_669_499# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.92e+06u
M1008 a_110_70# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 a_670_93# a_537_119# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1010 VPWR a_1169_93# a_1157_453# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.526e+11p ps=1.58e+06u
M1011 VPWR a_1513_137# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1012 VPWR a_1169_93# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Q a_1169_93# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1014 VGND a_1169_93# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_110_70# a_236_463# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1016 a_537_119# a_236_463# a_429_119# VPB phighvt w=420000u l=150000u
+  ad=2.424e+11p pd=2.14e+06u as=1.176e+11p ps=1.4e+06u
M1017 a_669_499# a_110_70# a_537_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1169_93# a_1513_137# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1019 a_1157_453# a_236_463# a_982_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=5.628e+11p ps=3.13e+06u
M1020 Q_N a_1513_137# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1021 VPWR a_1169_93# a_1513_137# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1022 a_670_93# a_537_119# VGND VNB nshort w=640000u l=150000u
+  ad=2.158e+11p pd=2.03e+06u as=0p ps=0u
M1023 a_982_369# a_110_70# a_670_93# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_429_119# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_982_369# a_236_463# a_670_93# VNB nshort w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=0p ps=0u
M1026 a_1125_119# a_110_70# a_982_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_429_119# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_110_70# a_236_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1029 VGND a_1513_137# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1169_93# a_982_369# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1031 Q_N a_1513_137# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

