* File: sky130_fd_sc_lp__invkapwr_2.pxi.spice
* Created: Wed Sep  2 09:56:33 2020
* 
x_PM_SKY130_FD_SC_LP__INVKAPWR_2%A N_A_M1001_g N_A_M1002_g N_A_M1000_g
+ N_A_M1004_g N_A_M1003_g A A N_A_c_32_n N_A_c_33_n
+ PM_SKY130_FD_SC_LP__INVKAPWR_2%A
x_PM_SKY130_FD_SC_LP__INVKAPWR_2%Y N_Y_M1000_d N_Y_M1001_s N_Y_M1002_s
+ N_Y_c_88_n N_Y_c_83_n N_Y_c_84_n N_Y_c_93_n N_Y_c_78_n N_Y_c_85_n N_Y_c_86_n
+ N_Y_c_79_n Y Y N_Y_c_82_n PM_SKY130_FD_SC_LP__INVKAPWR_2%Y
x_PM_SKY130_FD_SC_LP__INVKAPWR_2%KAPWR N_KAPWR_M1001_d N_KAPWR_M1004_d KAPWR
+ N_KAPWR_c_139_n N_KAPWR_c_142_n N_KAPWR_c_133_n KAPWR
+ PM_SKY130_FD_SC_LP__INVKAPWR_2%KAPWR
x_PM_SKY130_FD_SC_LP__INVKAPWR_2%VGND N_VGND_M1000_s N_VGND_M1003_s
+ N_VGND_c_156_n N_VGND_c_157_n N_VGND_c_158_n VGND N_VGND_c_159_n
+ N_VGND_c_160_n N_VGND_c_161_n N_VGND_c_162_n
+ PM_SKY130_FD_SC_LP__INVKAPWR_2%VGND
x_PM_SKY130_FD_SC_LP__INVKAPWR_2%VPWR VPWR N_VPWR_c_180_n VPWR
+ PM_SKY130_FD_SC_LP__INVKAPWR_2%VPWR
cc_1 VNB N_A_M1000_g 0.0525956f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.56
cc_2 VNB N_A_M1003_g 0.0435876f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=0.56
cc_3 VNB N_A_c_32_n 0.0293436f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.46
cc_4 VNB N_A_c_33_n 0.084547f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.485
cc_5 VNB N_Y_c_78_n 0.00149799f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.485
cc_6 VNB N_Y_c_79_n 0.00456845f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.485
cc_7 VNB Y 0.00295631f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.46
cc_8 VNB Y 0.0291489f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.485
cc_9 VNB N_Y_c_82_n 0.0103855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_156_n 0.0256902f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.295
cc_11 VNB N_VGND_c_157_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.56
cc_12 VNB N_VGND_c_158_n 0.0222797f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.675
cc_13 VNB N_VGND_c_159_n 0.0223503f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.295
cc_14 VNB N_VGND_c_160_n 0.0160313f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_15 VNB N_VGND_c_161_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.46
cc_16 VNB N_VGND_c_162_n 0.152942f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.46
cc_17 VNB VPWR 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.675
cc_18 VPB N_A_M1001_g 0.0233545f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_19 VPB N_A_M1002_g 0.0176925f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_20 VPB N_A_M1004_g 0.0223382f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_21 VPB N_A_c_33_n 0.00870531f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.485
cc_22 VPB N_Y_c_83_n 0.00234264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 VPB N_Y_c_84_n 0.0176848f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=1.295
cc_24 VPB N_Y_c_85_n 0.0132482f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.46
cc_25 VPB N_Y_c_86_n 0.00209286f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.485
cc_26 VPB Y 0.00298715f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.485
cc_27 VPB N_KAPWR_c_133_n 0.0310203f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_28 VPB VPWR 0.0438343f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.675
cc_29 VPB N_VPWR_c_180_n 0.0561076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 N_A_M1001_g N_Y_c_88_n 0.0023724f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_31 N_A_M1001_g N_Y_c_83_n 0.0153265f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_32 N_A_M1002_g N_Y_c_83_n 0.0143812f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_33 N_A_c_32_n N_Y_c_83_n 0.0436107f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_34 N_A_c_33_n N_Y_c_83_n 0.002829f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_35 N_A_M1002_g N_Y_c_93_n 8.22659e-19 $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_36 N_A_M1004_g N_Y_c_93_n 8.22659e-19 $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_37 N_A_M1000_g N_Y_c_78_n 0.00189162f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_38 N_A_M1003_g N_Y_c_78_n 0.00180689f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_39 N_A_M1004_g N_Y_c_85_n 0.0159989f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_40 N_A_c_32_n N_Y_c_85_n 0.0110823f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_41 N_A_c_33_n N_Y_c_85_n 0.00322171f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_42 N_A_c_32_n N_Y_c_86_n 0.0219511f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_43 N_A_c_33_n N_Y_c_86_n 0.00314903f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_44 N_A_M1000_g N_Y_c_79_n 0.006617f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_45 N_A_c_32_n N_Y_c_79_n 0.0198419f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_46 N_A_c_33_n N_Y_c_79_n 6.24756e-19 $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_47 N_A_M1003_g Y 0.0152312f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_48 N_A_c_32_n Y 0.00755553f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_49 N_A_M1003_g Y 0.0205853f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_50 N_A_c_32_n Y 0.0267298f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_51 N_A_c_33_n Y 0.00240773f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_52 N_A_M1001_g N_KAPWR_c_133_n 0.00731133f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A_M1002_g N_KAPWR_c_133_n 0.00731133f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_M1004_g N_KAPWR_c_133_n 0.00731133f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A_M1000_g N_VGND_c_156_n 0.00406185f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_56 N_A_c_32_n N_VGND_c_156_n 0.0110952f $X=1.26 $Y=1.46 $X2=0 $Y2=0
cc_57 N_A_c_33_n N_VGND_c_156_n 0.00153298f $X=1.355 $Y=1.485 $X2=0 $Y2=0
cc_58 N_A_M1000_g N_VGND_c_158_n 5.44985e-19 $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_VGND_c_158_n 0.00957799f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_VGND_c_160_n 0.00478016f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_61 N_A_M1003_g N_VGND_c_160_n 0.00396895f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VGND_c_162_n 0.0096052f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_63 N_A_M1003_g N_VGND_c_162_n 0.00397666f $X=1.445 $Y=0.56 $X2=0 $Y2=0
cc_64 N_A_M1001_g VPWR 0.00634705f $X=0.495 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_65 N_A_M1002_g VPWR 0.0053229f $X=0.925 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_66 N_A_M1004_g VPWR 0.00633019f $X=1.355 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_67 N_A_M1001_g N_VPWR_c_180_n 0.00585385f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_M1002_g N_VPWR_c_180_n 0.00585385f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A_M1004_g N_VPWR_c_180_n 0.00585385f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_70 N_Y_c_83_n N_KAPWR_M1001_d 0.00176461f $X=1.01 $Y=1.8 $X2=-0.19 $Y2=-0.245
cc_71 N_Y_c_85_n N_KAPWR_M1004_d 0.00246823f $X=1.595 $Y=1.8 $X2=0 $Y2=0
cc_72 N_Y_c_88_n N_KAPWR_c_139_n 0.0091127f $X=0.28 $Y=2 $X2=0 $Y2=0
cc_73 N_Y_c_83_n N_KAPWR_c_139_n 0.0135055f $X=1.01 $Y=1.8 $X2=0 $Y2=0
cc_74 N_Y_c_93_n N_KAPWR_c_139_n 0.00911549f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_75 N_Y_c_93_n N_KAPWR_c_142_n 0.0091127f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_76 N_Y_c_85_n N_KAPWR_c_142_n 0.0176763f $X=1.595 $Y=1.8 $X2=0 $Y2=0
cc_77 N_Y_M1001_s N_KAPWR_c_133_n 3.61265e-19 $X=0.155 $Y=1.835 $X2=0 $Y2=0
cc_78 N_Y_M1002_s N_KAPWR_c_133_n 7.22529e-19 $X=1 $Y=1.835 $X2=0 $Y2=0
cc_79 N_Y_c_88_n N_KAPWR_c_133_n 0.0313835f $X=0.28 $Y=2 $X2=0 $Y2=0
cc_80 N_Y_c_93_n N_KAPWR_c_133_n 0.0288605f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_81 Y N_VGND_c_158_n 0.00530131f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_82 N_Y_c_82_n N_VGND_c_158_n 0.0165893f $X=1.687 $Y=1.04 $X2=0 $Y2=0
cc_83 N_Y_c_78_n N_VGND_c_160_n 0.00717541f $X=1.23 $Y=0.56 $X2=0 $Y2=0
cc_84 N_Y_c_78_n N_VGND_c_162_n 0.00799322f $X=1.23 $Y=0.56 $X2=0 $Y2=0
cc_85 Y N_VGND_c_162_n 0.00538134f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_86 N_Y_c_82_n N_VGND_c_162_n 6.73317e-19 $X=1.687 $Y=1.04 $X2=0 $Y2=0
cc_87 N_Y_M1001_s VPWR 0.00115465f $X=0.155 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_88 N_Y_M1002_s VPWR 0.0012358f $X=1 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_89 N_Y_c_88_n VPWR 0.0024325f $X=0.28 $Y=2 $X2=-0.19 $Y2=-0.245
cc_90 N_Y_c_93_n VPWR 0.00248057f $X=1.14 $Y=2 $X2=-0.19 $Y2=-0.245
cc_91 N_Y_c_88_n N_VPWR_c_180_n 0.0135826f $X=0.28 $Y=2 $X2=0 $Y2=0
cc_92 N_Y_c_93_n N_VPWR_c_180_n 0.012556f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_93 N_KAPWR_M1001_d VPWR 0.00121489f $X=0.57 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_94 N_KAPWR_M1004_d VPWR 0.00114194f $X=1.43 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_95 N_KAPWR_c_139_n VPWR 0.00242444f $X=0.71 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_96 N_KAPWR_c_142_n VPWR 0.00237745f $X=1.57 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_97 N_KAPWR_c_133_n VPWR 0.185305f $X=1.565 $Y=2.81 $X2=-0.19 $Y2=1.655
cc_98 N_KAPWR_c_139_n N_VPWR_c_180_n 0.0149362f $X=0.71 $Y=2.22 $X2=0 $Y2=0
cc_99 N_KAPWR_c_142_n N_VPWR_c_180_n 0.0161868f $X=1.57 $Y=2.22 $X2=0 $Y2=0
cc_100 N_KAPWR_c_133_n N_VPWR_c_180_n 0.00456099f $X=1.565 $Y=2.81 $X2=0 $Y2=0
