* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y a_44_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_842_67# C a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_324_45# a_44_69# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_324_45# a_217_69# a_842_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_1251_47# C a_842_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_324_45# a_44_69# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR a_217_69# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR a_44_69# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 Y a_44_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_1251_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND D a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_44_69# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_1251_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Y a_217_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR a_217_69# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR a_44_69# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 Y a_217_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 Y a_44_69# a_324_45# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_842_67# a_217_69# a_324_45# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VGND B_N a_217_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VGND D a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 Y a_44_69# a_324_45# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_842_67# C a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 VPWR B_N a_217_69# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_44_69# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 a_842_67# a_217_69# a_324_45# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_324_45# a_217_69# a_842_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 a_1251_47# C a_842_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
