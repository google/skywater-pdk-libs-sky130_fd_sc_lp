# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o21a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.585000 1.425000 3.915000 1.675000 ;
        RECT 3.745000 1.675000 3.915000 2.310000 ;
        RECT 3.745000 2.310000 5.125000 2.500000 ;
        RECT 4.955000 1.425000 5.430000 1.645000 ;
        RECT 4.955000 1.645000 5.125000 2.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.425000 4.775000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.425000 3.185000 1.760000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.695000 1.225000 ;
        RECT 0.085000 1.225000 0.350000 1.755000 ;
        RECT 0.085000 1.755000 2.005000 1.925000 ;
        RECT 0.645000 0.255000 0.835000 1.055000 ;
        RECT 0.965000 1.925000 1.155000 3.075000 ;
        RECT 1.505000 0.255000 1.695000 1.055000 ;
        RECT 1.825000 1.925000 2.005000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.145000  0.085000 0.475000 0.885000 ;
      RECT 0.465000  2.095000 0.795000 3.245000 ;
      RECT 0.520000  1.395000 2.345000 1.585000 ;
      RECT 1.005000  0.085000 1.335000 0.885000 ;
      RECT 1.325000  2.095000 1.655000 3.245000 ;
      RECT 1.865000  0.085000 2.195000 0.905000 ;
      RECT 2.175000  1.075000 4.265000 1.245000 ;
      RECT 2.175000  1.245000 2.345000 1.395000 ;
      RECT 2.175000  1.585000 2.345000 1.930000 ;
      RECT 2.175000  1.930000 2.875000 2.100000 ;
      RECT 2.185000  2.270000 2.515000 3.245000 ;
      RECT 2.415000  0.255000 3.755000 0.425000 ;
      RECT 2.415000  0.425000 2.745000 0.895000 ;
      RECT 2.685000  2.100000 2.875000 3.075000 ;
      RECT 2.915000  0.595000 3.245000 1.075000 ;
      RECT 3.045000  2.805000 3.815000 3.245000 ;
      RECT 3.245000  1.925000 3.575000 2.805000 ;
      RECT 3.425000  0.425000 3.755000 0.735000 ;
      RECT 3.425000  0.735000 4.625000 0.905000 ;
      RECT 3.925000  0.085000 4.265000 0.565000 ;
      RECT 3.995000  2.670000 5.065000 3.000000 ;
      RECT 4.085000  1.245000 4.265000 1.930000 ;
      RECT 4.085000  1.930000 4.695000 2.140000 ;
      RECT 4.435000  0.305000 4.625000 0.735000 ;
      RECT 4.435000  0.905000 4.625000 1.085000 ;
      RECT 4.435000  1.085000 5.555000 1.255000 ;
      RECT 4.795000  0.085000 5.125000 0.915000 ;
      RECT 5.295000  0.305000 5.555000 1.085000 ;
      RECT 5.295000  1.815000 5.555000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__o21a_4
END LIBRARY
