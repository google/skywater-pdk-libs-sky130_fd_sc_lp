* File: sky130_fd_sc_lp__dlxbp_lp2.pxi.spice
* Created: Wed Sep  2 09:48:11 2020
* 
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%D N_D_M1011_g N_D_M1018_g N_D_M1000_g
+ N_D_c_170_n N_D_c_171_n D D N_D_c_173_n PM_SKY130_FD_SC_LP__DLXBP_LP2%D
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%GATE N_GATE_M1005_g N_GATE_M1021_g
+ N_GATE_M1012_g GATE GATE N_GATE_c_208_n PM_SKY130_FD_SC_LP__DLXBP_LP2%GATE
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%A_278_409# N_A_278_409#_M1012_d
+ N_A_278_409#_M1005_d N_A_278_409#_M1003_g N_A_278_409#_M1019_g
+ N_A_278_409#_M1020_g N_A_278_409#_M1009_g N_A_278_409#_M1013_g
+ N_A_278_409#_c_259_n N_A_278_409#_c_260_n N_A_278_409#_c_261_n
+ N_A_278_409#_c_269_n N_A_278_409#_c_262_n N_A_278_409#_c_263_n
+ N_A_278_409#_c_301_p N_A_278_409#_c_264_n N_A_278_409#_c_265_n
+ N_A_278_409#_c_272_n N_A_278_409#_c_266_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP2%A_278_409#
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%A_27_57# N_A_27_57#_M1011_s N_A_27_57#_M1018_s
+ N_A_27_57#_c_387_n N_A_27_57#_M1027_g N_A_27_57#_c_389_n N_A_27_57#_M1006_g
+ N_A_27_57#_c_391_n N_A_27_57#_c_392_n N_A_27_57#_c_393_n N_A_27_57#_c_394_n
+ N_A_27_57#_c_385_n N_A_27_57#_c_395_n N_A_27_57#_c_386_n N_A_27_57#_c_397_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP2%A_27_57#
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%A_461_55# N_A_461_55#_M1003_s
+ N_A_461_55#_M1019_s N_A_461_55#_M1007_g N_A_461_55#_M1016_g
+ N_A_461_55#_c_457_n N_A_461_55#_c_458_n N_A_461_55#_c_459_n
+ N_A_461_55#_c_460_n N_A_461_55#_c_461_n N_A_461_55#_c_462_n
+ N_A_461_55#_c_463_n N_A_461_55#_c_470_n N_A_461_55#_c_464_n
+ N_A_461_55#_c_465_n N_A_461_55#_c_466_n N_A_461_55#_c_467_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP2%A_461_55#
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%A_934_29# N_A_934_29#_M1024_d
+ N_A_934_29#_M1023_d N_A_934_29#_c_555_n N_A_934_29#_M1014_g
+ N_A_934_29#_c_556_n N_A_934_29#_c_557_n N_A_934_29#_c_558_n
+ N_A_934_29#_M1001_g N_A_934_29#_M1002_g N_A_934_29#_c_560_n
+ N_A_934_29#_c_561_n N_A_934_29#_M1025_g N_A_934_29#_M1010_g
+ N_A_934_29#_M1004_g N_A_934_29#_M1026_g N_A_934_29#_M1008_g
+ N_A_934_29#_c_567_n N_A_934_29#_c_577_n N_A_934_29#_c_568_n
+ N_A_934_29#_c_569_n N_A_934_29#_c_570_n N_A_934_29#_c_579_n
+ N_A_934_29#_c_625_p N_A_934_29#_c_571_n N_A_934_29#_c_572_n
+ N_A_934_29#_c_573_n PM_SKY130_FD_SC_LP__DLXBP_LP2%A_934_29#
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%A_784_55# N_A_784_55#_M1007_d
+ N_A_784_55#_M1009_d N_A_784_55#_c_708_n N_A_784_55#_M1022_g
+ N_A_784_55#_c_709_n N_A_784_55#_c_710_n N_A_784_55#_c_711_n
+ N_A_784_55#_M1024_g N_A_784_55#_M1023_g N_A_784_55#_c_713_n
+ N_A_784_55#_c_728_n N_A_784_55#_c_724_n N_A_784_55#_c_725_n
+ N_A_784_55#_c_726_n N_A_784_55#_c_714_n N_A_784_55#_c_715_n
+ N_A_784_55#_c_716_n N_A_784_55#_c_717_n N_A_784_55#_c_718_n
+ N_A_784_55#_c_719_n N_A_784_55#_c_720_n N_A_784_55#_c_721_n
+ N_A_784_55#_c_722_n PM_SKY130_FD_SC_LP__DLXBP_LP2%A_784_55#
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%A_1662_57# N_A_1662_57#_M1008_d
+ N_A_1662_57#_M1026_d N_A_1662_57#_M1015_g N_A_1662_57#_M1028_g
+ N_A_1662_57#_M1017_g N_A_1662_57#_c_823_n N_A_1662_57#_c_829_n
+ N_A_1662_57#_c_824_n N_A_1662_57#_c_825_n N_A_1662_57#_c_826_n
+ N_A_1662_57#_c_827_n PM_SKY130_FD_SC_LP__DLXBP_LP2%A_1662_57#
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%VPWR N_VPWR_M1018_d N_VPWR_M1019_d
+ N_VPWR_M1001_d N_VPWR_M1010_d N_VPWR_M1028_s N_VPWR_c_872_n N_VPWR_c_873_n
+ N_VPWR_c_874_n N_VPWR_c_875_n N_VPWR_c_876_n N_VPWR_c_877_n N_VPWR_c_878_n
+ N_VPWR_c_879_n VPWR N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n
+ N_VPWR_c_883_n N_VPWR_c_871_n N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n
+ N_VPWR_c_888_n PM_SKY130_FD_SC_LP__DLXBP_LP2%VPWR
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%Q N_Q_M1002_s N_Q_M1010_s N_Q_c_963_n Q Q Q Q Q
+ N_Q_c_966_n PM_SKY130_FD_SC_LP__DLXBP_LP2%Q
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%Q_N N_Q_N_M1017_d N_Q_N_M1028_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N Q_N PM_SKY130_FD_SC_LP__DLXBP_LP2%Q_N
x_PM_SKY130_FD_SC_LP__DLXBP_LP2%VGND N_VGND_M1000_d N_VGND_M1020_d
+ N_VGND_M1014_d N_VGND_M1025_d N_VGND_M1015_s N_VGND_c_1017_n N_VGND_c_1018_n
+ N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n
+ N_VGND_c_1023_n N_VGND_c_1024_n VGND N_VGND_c_1025_n N_VGND_c_1026_n
+ N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n
+ N_VGND_c_1031_n N_VGND_c_1032_n N_VGND_c_1033_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP2%VGND
cc_1 VNB N_D_M1011_g 0.035665f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_2 VNB N_D_M1000_g 0.0307794f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_3 VNB N_D_c_170_n 0.017139f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.26
cc_4 VNB N_D_c_171_n 0.010672f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.78
cc_5 VNB D 0.00121962f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_D_c_173_n 0.0257984f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.275
cc_7 VNB N_GATE_M1021_g 0.031794f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.545
cc_8 VNB N_GATE_M1012_g 0.0400864f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_9 VNB GATE 0.00137587f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.26
cc_10 VNB N_GATE_c_208_n 0.0699556f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.275
cc_11 VNB N_A_278_409#_M1003_g 0.0388713f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.11
cc_12 VNB N_A_278_409#_M1019_g 0.00131742f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.26
cc_13 VNB N_A_278_409#_M1020_g 0.0316037f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.78
cc_14 VNB N_A_278_409#_M1013_g 0.059716f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.275
cc_15 VNB N_A_278_409#_c_259_n 0.00174902f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.665
cc_16 VNB N_A_278_409#_c_260_n 0.0188382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_278_409#_c_261_n 0.0024114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_278_409#_c_262_n 0.00773762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_278_409#_c_263_n 0.00323781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_278_409#_c_264_n 0.00739663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_278_409#_c_265_n 0.0189114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_278_409#_c_266_n 0.0402928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_57#_M1006_g 0.0586108f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.26
cc_24 VNB N_A_27_57#_c_385_n 0.0251105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_57#_c_386_n 0.0443842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_461_55#_c_457_n 0.00761141f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.54
cc_27 VNB N_A_461_55#_c_458_n 0.0128079f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_28 VNB N_A_461_55#_c_459_n 0.00743362f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.275
cc_29 VNB N_A_461_55#_c_460_n 0.00186107f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.275
cc_30 VNB N_A_461_55#_c_461_n 0.0309867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_461_55#_c_462_n 0.0043183f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.665
cc_32 VNB N_A_461_55#_c_463_n 0.00772043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_461_55#_c_464_n 0.0188102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_461_55#_c_465_n 0.00804321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_461_55#_c_466_n 0.00984061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_461_55#_c_467_n 0.0178715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_934_29#_c_555_n 0.0175403f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.545
cc_38 VNB N_A_934_29#_c_556_n 0.0350592f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_39 VNB N_A_934_29#_c_557_n 0.00844801f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_40 VNB N_A_934_29#_c_558_n 0.03962f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.26
cc_41 VNB N_A_934_29#_M1002_g 0.0228151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_934_29#_c_560_n 0.00996185f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.275
cc_43 VNB N_A_934_29#_c_561_n 0.0312056f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.275
cc_44 VNB N_A_934_29#_M1025_g 0.0191254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_934_29#_M1010_g 0.0416435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_934_29#_M1004_g 0.0191427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_934_29#_M1026_g 0.0400953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_934_29#_M1008_g 0.0239513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_934_29#_c_567_n 0.0308438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_934_29#_c_568_n 0.0179672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_934_29#_c_569_n 0.00766002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_934_29#_c_570_n 0.00865238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_934_29#_c_571_n 0.0433077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_934_29#_c_572_n 0.00272419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_934_29#_c_573_n 0.0151436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_784_55#_c_708_n 0.0180097f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.545
cc_57 VNB N_A_784_55#_c_709_n 0.00970588f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_58 VNB N_A_784_55#_c_710_n 0.00970563f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_59 VNB N_A_784_55#_c_711_n 0.017515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_784_55#_M1023_g 0.00403873f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_61 VNB N_A_784_55#_c_713_n 0.00626823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_784_55#_c_714_n 0.00580407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_784_55#_c_715_n 0.0102495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_784_55#_c_716_n 0.00323583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_784_55#_c_717_n 0.00316957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_784_55#_c_718_n 0.0213319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_784_55#_c_719_n 5.98074e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_784_55#_c_720_n 0.00242631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_784_55#_c_721_n 0.0337392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_784_55#_c_722_n 0.0141565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1662_57#_M1015_g 0.024094f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.11
cc_72 VNB N_A_1662_57#_M1017_g 0.0260751f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.78
cc_73 VNB N_A_1662_57#_c_823_n 0.0174655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1662_57#_c_824_n 0.00868302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1662_57#_c_825_n 0.00276577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1662_57#_c_826_n 3.00516e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1662_57#_c_827_n 0.0901812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VPWR_c_871_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_Q_c_963_n 0.00631488f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.545
cc_80 VNB Q 0.0077495f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.26
cc_81 VNB Q 0.00435942f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.11
cc_82 VNB N_Q_c_966_n 0.00389826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB Q_N 0.0576865f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.545
cc_84 VNB N_VGND_c_1017_n 0.00420298f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_85 VNB N_VGND_c_1018_n 0.0516021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1019_n 0.00151893f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.275
cc_87 VNB N_VGND_c_1020_n 0.0102717f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.665
cc_88 VNB N_VGND_c_1021_n 0.00934305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1022_n 0.017938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1023_n 0.0587682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1024_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1025_n 0.0271986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1026_n 0.0439496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1027_n 0.0286512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1028_n 0.028795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1029_n 0.578736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1030_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1031_n 0.00485883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1032_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1033_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VPB N_D_M1018_g 0.0403693f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.545
cc_102 VPB N_D_c_171_n 0.0207303f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.78
cc_103 VPB D 0.00544765f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_104 VPB N_GATE_M1005_g 0.0375127f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.495
cc_105 VPB GATE 0.00369843f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.26
cc_106 VPB N_GATE_c_208_n 0.0387988f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.275
cc_107 VPB N_A_278_409#_M1019_g 0.0267382f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.26
cc_108 VPB N_A_278_409#_M1009_g 0.0332158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_278_409#_c_269_n 0.0312688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_278_409#_c_264_n 0.0157585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_278_409#_c_265_n 0.0286621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_278_409#_c_272_n 0.0093578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_27_57#_c_387_n 0.0975314f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.545
cc_114 VPB N_A_27_57#_M1027_g 0.00730077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_27_57#_c_389_n 0.0123826f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.26
cc_116 VPB N_A_27_57#_M1006_g 0.0145961f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.26
cc_117 VPB N_A_27_57#_c_391_n 0.0129495f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_27_57#_c_392_n 0.0122735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_27_57#_c_393_n 8.09409e-19 $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.275
cc_120 VPB N_A_27_57#_c_394_n 0.0654114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_27_57#_c_395_n 0.0139041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_27_57#_c_386_n 0.0178668f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_27_57#_c_397_n 0.0234767f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_461_55#_M1016_g 0.0300348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_461_55#_c_458_n 0.00439235f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_126 VPB N_A_461_55#_c_470_n 0.0181256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_461_55#_c_465_n 0.0129071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_461_55#_c_466_n 0.0230685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_934_29#_M1001_g 0.0292762f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.54
cc_130 VPB N_A_934_29#_M1010_g 0.0303756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_934_29#_M1026_g 0.0282186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_934_29#_c_577_n 0.010732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_934_29#_c_570_n 0.021522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_934_29#_c_579_n 0.0235085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_934_29#_c_571_n 0.00661054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_934_29#_c_572_n 0.00300155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_934_29#_c_573_n 0.0366577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_784_55#_M1023_g 0.0542989f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_139 VPB N_A_784_55#_c_724_n 0.00325539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_784_55#_c_725_n 0.00434674f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.665
cc_141 VPB N_A_784_55#_c_726_n 0.00414135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_784_55#_c_717_n 0.0034024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1662_57#_M1028_g 0.0431808f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.26
cc_144 VPB N_A_1662_57#_c_829_n 0.0148884f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.275
cc_145 VPB N_A_1662_57#_c_824_n 0.0115087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_1662_57#_c_826_n 4.85449e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_1662_57#_c_827_n 0.0191159f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_872_n 0.00561105f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_149 VPB N_VPWR_c_873_n 0.0110955f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.275
cc_150 VPB N_VPWR_c_874_n 0.00983154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_875_n 0.0256426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_876_n 0.0221169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_877_n 0.0197914f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_878_n 0.0215888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_879_n 0.00631318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_880_n 0.0538946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_881_n 0.057433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_882_n 0.0559589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_883_n 0.0254718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_871_n 0.136282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_885_n 0.00449074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_886_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_887_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_888_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB Q 0.0295921f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.11
cc_166 VPB Q_N 0.0220411f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.545
cc_167 VPB Q_N 0.0648075f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.26
cc_168 N_D_M1000_g N_GATE_M1021_g 0.0261883f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_169 N_D_M1018_g N_GATE_c_208_n 0.038296f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_170 N_D_c_170_n N_GATE_c_208_n 0.0414783f $X=0.675 $Y=1.26 $X2=0 $Y2=0
cc_171 D N_GATE_c_208_n 0.00219001f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_172 N_D_M1018_g N_A_278_409#_c_259_n 0.00128705f $X=0.575 $Y=2.545 $X2=0
+ $Y2=0
cc_173 N_D_M1000_g N_A_278_409#_c_259_n 0.00257169f $X=0.855 $Y=0.495 $X2=0
+ $Y2=0
cc_174 N_D_c_170_n N_A_278_409#_c_259_n 0.002136f $X=0.675 $Y=1.26 $X2=0 $Y2=0
cc_175 D N_A_278_409#_c_259_n 0.0252621f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_176 N_D_M1000_g N_A_278_409#_c_261_n 0.00413741f $X=0.855 $Y=0.495 $X2=0
+ $Y2=0
cc_177 N_D_M1018_g N_A_278_409#_c_272_n 0.00171003f $X=0.575 $Y=2.545 $X2=0
+ $Y2=0
cc_178 N_D_M1018_g N_A_27_57#_c_391_n 0.00753306f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_179 N_D_M1018_g N_A_27_57#_c_392_n 0.0217745f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_180 N_D_M1011_g N_A_27_57#_c_385_n 0.0101678f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_181 N_D_M1000_g N_A_27_57#_c_385_n 0.00143555f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_182 N_D_M1018_g N_A_27_57#_c_395_n 0.00577384f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_183 N_D_M1011_g N_A_27_57#_c_386_n 0.0158222f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_184 D N_A_27_57#_c_386_n 0.0414404f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_185 N_D_c_173_n N_A_27_57#_c_386_n 0.0200357f $X=0.67 $Y=1.275 $X2=0 $Y2=0
cc_186 N_D_M1018_g N_A_27_57#_c_397_n 0.00838332f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_187 N_D_M1018_g N_VPWR_c_872_n 0.00408642f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_188 N_D_M1018_g N_VPWR_c_878_n 0.0063172f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_189 N_D_M1018_g N_VPWR_c_871_n 0.0090514f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_190 N_D_M1011_g N_VGND_c_1017_n 0.00189426f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_191 N_D_M1000_g N_VGND_c_1017_n 0.0114298f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_192 N_D_M1011_g N_VGND_c_1025_n 0.00502664f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_193 N_D_M1000_g N_VGND_c_1025_n 0.00445056f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_194 N_D_M1011_g N_VGND_c_1029_n 0.0100616f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_195 N_D_M1000_g N_VGND_c_1029_n 0.00796275f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_196 N_GATE_M1005_g N_A_278_409#_c_259_n 0.0127843f $X=1.265 $Y=2.545 $X2=0
+ $Y2=0
cc_197 N_GATE_M1021_g N_A_278_409#_c_259_n 0.00534827f $X=1.315 $Y=0.495 $X2=0
+ $Y2=0
cc_198 N_GATE_M1012_g N_A_278_409#_c_259_n 0.0011866f $X=1.675 $Y=0.495 $X2=0
+ $Y2=0
cc_199 GATE N_A_278_409#_c_259_n 0.0457028f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_200 N_GATE_c_208_n N_A_278_409#_c_259_n 0.0282074f $X=1.73 $Y=1.34 $X2=0
+ $Y2=0
cc_201 N_GATE_M1021_g N_A_278_409#_c_260_n 0.00156812f $X=1.315 $Y=0.495 $X2=0
+ $Y2=0
cc_202 N_GATE_M1012_g N_A_278_409#_c_260_n 0.0122732f $X=1.675 $Y=0.495 $X2=0
+ $Y2=0
cc_203 GATE N_A_278_409#_c_260_n 0.0259452f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_204 N_GATE_c_208_n N_A_278_409#_c_260_n 0.00233943f $X=1.73 $Y=1.34 $X2=0
+ $Y2=0
cc_205 N_GATE_M1021_g N_A_278_409#_c_261_n 0.0069586f $X=1.315 $Y=0.495 $X2=0
+ $Y2=0
cc_206 GATE N_A_278_409#_c_269_n 0.0094082f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_207 N_GATE_c_208_n N_A_278_409#_c_269_n 0.00119479f $X=1.73 $Y=1.34 $X2=0
+ $Y2=0
cc_208 N_GATE_M1021_g N_A_278_409#_c_262_n 0.0019515f $X=1.315 $Y=0.495 $X2=0
+ $Y2=0
cc_209 N_GATE_M1012_g N_A_278_409#_c_262_n 0.0129546f $X=1.675 $Y=0.495 $X2=0
+ $Y2=0
cc_210 N_GATE_M1005_g N_A_278_409#_c_272_n 0.0151713f $X=1.265 $Y=2.545 $X2=0
+ $Y2=0
cc_211 GATE N_A_278_409#_c_272_n 0.0103542f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_212 N_GATE_c_208_n N_A_278_409#_c_272_n 0.00864712f $X=1.73 $Y=1.34 $X2=0
+ $Y2=0
cc_213 N_GATE_c_208_n N_A_278_409#_c_266_n 0.00369333f $X=1.73 $Y=1.34 $X2=0
+ $Y2=0
cc_214 N_GATE_M1005_g N_A_27_57#_c_392_n 0.0221153f $X=1.265 $Y=2.545 $X2=0
+ $Y2=0
cc_215 N_GATE_M1005_g N_A_27_57#_c_393_n 0.00258788f $X=1.265 $Y=2.545 $X2=0
+ $Y2=0
cc_216 N_GATE_M1005_g N_A_27_57#_c_394_n 0.0105671f $X=1.265 $Y=2.545 $X2=0
+ $Y2=0
cc_217 N_GATE_M1005_g N_A_27_57#_c_395_n 0.00209591f $X=1.265 $Y=2.545 $X2=0
+ $Y2=0
cc_218 N_GATE_M1005_g N_A_27_57#_c_397_n 8.4847e-19 $X=1.265 $Y=2.545 $X2=0
+ $Y2=0
cc_219 N_GATE_M1012_g N_A_461_55#_c_457_n 0.00130312f $X=1.675 $Y=0.495 $X2=0
+ $Y2=0
cc_220 N_GATE_M1012_g N_A_461_55#_c_458_n 0.00423221f $X=1.675 $Y=0.495 $X2=0
+ $Y2=0
cc_221 GATE N_A_461_55#_c_458_n 0.0202139f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_222 N_GATE_c_208_n N_A_461_55#_c_458_n 0.00720351f $X=1.73 $Y=1.34 $X2=0
+ $Y2=0
cc_223 N_GATE_M1012_g N_A_461_55#_c_463_n 7.3292e-19 $X=1.675 $Y=0.495 $X2=0
+ $Y2=0
cc_224 GATE N_A_461_55#_c_470_n 0.00743911f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_225 N_GATE_c_208_n N_A_461_55#_c_470_n 0.00389405f $X=1.73 $Y=1.34 $X2=0
+ $Y2=0
cc_226 N_GATE_M1005_g N_VPWR_c_872_n 0.00442529f $X=1.265 $Y=2.545 $X2=0 $Y2=0
cc_227 N_GATE_M1005_g N_VPWR_c_880_n 0.0063971f $X=1.265 $Y=2.545 $X2=0 $Y2=0
cc_228 N_GATE_M1005_g N_VPWR_c_871_n 0.00887298f $X=1.265 $Y=2.545 $X2=0 $Y2=0
cc_229 N_GATE_M1021_g N_VGND_c_1017_n 0.00304977f $X=1.315 $Y=0.495 $X2=0 $Y2=0
cc_230 N_GATE_c_208_n N_VGND_c_1017_n 0.00197584f $X=1.73 $Y=1.34 $X2=0 $Y2=0
cc_231 N_GATE_M1021_g N_VGND_c_1018_n 0.0053602f $X=1.315 $Y=0.495 $X2=0 $Y2=0
cc_232 N_GATE_M1012_g N_VGND_c_1018_n 0.00502664f $X=1.675 $Y=0.495 $X2=0 $Y2=0
cc_233 N_GATE_M1021_g N_VGND_c_1029_n 0.00561494f $X=1.315 $Y=0.495 $X2=0 $Y2=0
cc_234 N_GATE_M1012_g N_VGND_c_1029_n 0.00651958f $X=1.675 $Y=0.495 $X2=0 $Y2=0
cc_235 N_A_278_409#_M1019_g N_A_27_57#_c_387_n 0.0151533f $X=2.85 $Y=2.195 $X2=0
+ $Y2=0
cc_236 N_A_278_409#_c_269_n N_A_27_57#_M1027_g 0.00454006f $X=2.93 $Y=2.27 $X2=0
+ $Y2=0
cc_237 N_A_278_409#_M1019_g N_A_27_57#_c_389_n 0.0278412f $X=2.85 $Y=2.195 $X2=0
+ $Y2=0
cc_238 N_A_278_409#_M1009_g N_A_27_57#_c_389_n 0.0750005f $X=3.95 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A_278_409#_c_301_p N_A_27_57#_c_389_n 0.00708747f $X=3.015 $Y=2.185
+ $X2=0 $Y2=0
cc_240 N_A_278_409#_c_264_n N_A_27_57#_c_389_n 0.00496808f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_241 N_A_278_409#_M1019_g N_A_27_57#_M1006_g 0.00905664f $X=2.85 $Y=2.195
+ $X2=0 $Y2=0
cc_242 N_A_278_409#_M1020_g N_A_27_57#_M1006_g 0.0437013f $X=3.025 $Y=0.485
+ $X2=0 $Y2=0
cc_243 N_A_278_409#_c_263_n N_A_27_57#_M1006_g 0.0016329f $X=3.015 $Y=1.755
+ $X2=0 $Y2=0
cc_244 N_A_278_409#_c_301_p N_A_27_57#_M1006_g 0.0015212f $X=3.015 $Y=2.185
+ $X2=0 $Y2=0
cc_245 N_A_278_409#_c_264_n N_A_27_57#_M1006_g 0.0241621f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_246 N_A_278_409#_c_265_n N_A_27_57#_M1006_g 0.0167186f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_247 N_A_278_409#_M1005_d N_A_27_57#_c_392_n 0.00722001f $X=1.39 $Y=2.045
+ $X2=0 $Y2=0
cc_248 N_A_278_409#_M1019_g N_A_27_57#_c_392_n 0.00549535f $X=2.85 $Y=2.195
+ $X2=0 $Y2=0
cc_249 N_A_278_409#_c_269_n N_A_27_57#_c_392_n 0.0262234f $X=2.93 $Y=2.27 $X2=0
+ $Y2=0
cc_250 N_A_278_409#_c_272_n N_A_27_57#_c_392_n 0.0484592f $X=1.695 $Y=2.19 $X2=0
+ $Y2=0
cc_251 N_A_278_409#_M1019_g N_A_27_57#_c_393_n 0.00139933f $X=2.85 $Y=2.195
+ $X2=0 $Y2=0
cc_252 N_A_278_409#_M1019_g N_A_27_57#_c_394_n 0.00274403f $X=2.85 $Y=2.195
+ $X2=0 $Y2=0
cc_253 N_A_278_409#_c_269_n N_A_27_57#_c_394_n 0.00143433f $X=2.93 $Y=2.27 $X2=0
+ $Y2=0
cc_254 N_A_278_409#_c_269_n N_A_461_55#_M1019_s 0.0121066f $X=2.93 $Y=2.27 $X2=0
+ $Y2=0
cc_255 N_A_278_409#_M1003_g N_A_461_55#_c_457_n 0.0124039f $X=2.665 $Y=0.485
+ $X2=0 $Y2=0
cc_256 N_A_278_409#_M1020_g N_A_461_55#_c_457_n 0.00190675f $X=3.025 $Y=0.485
+ $X2=0 $Y2=0
cc_257 N_A_278_409#_c_262_n N_A_461_55#_c_457_n 0.0370464f $X=1.89 $Y=0.495
+ $X2=0 $Y2=0
cc_258 N_A_278_409#_M1003_g N_A_461_55#_c_458_n 0.0111545f $X=2.665 $Y=0.485
+ $X2=0 $Y2=0
cc_259 N_A_278_409#_M1019_g N_A_461_55#_c_458_n 0.00386343f $X=2.85 $Y=2.195
+ $X2=0 $Y2=0
cc_260 N_A_278_409#_c_260_n N_A_461_55#_c_458_n 6.52458e-19 $X=1.725 $Y=0.91
+ $X2=0 $Y2=0
cc_261 N_A_278_409#_c_263_n N_A_461_55#_c_458_n 0.0224591f $X=3.015 $Y=1.755
+ $X2=0 $Y2=0
cc_262 N_A_278_409#_M1013_g N_A_461_55#_c_459_n 0.0161328f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_263 N_A_278_409#_c_265_n N_A_461_55#_c_459_n 0.00594474f $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_264 N_A_278_409#_c_264_n N_A_461_55#_c_460_n 0.0215966f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_265 N_A_278_409#_c_265_n N_A_461_55#_c_460_n 0.00110664f $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_266 N_A_278_409#_M1013_g N_A_461_55#_c_461_n 0.021337f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_267 N_A_278_409#_c_264_n N_A_461_55#_c_461_n 0.00301047f $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_268 N_A_278_409#_c_265_n N_A_461_55#_c_461_n 0.0114061f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_269 N_A_278_409#_M1013_g N_A_461_55#_c_462_n 0.0171448f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_270 N_A_278_409#_c_264_n N_A_461_55#_c_462_n 0.00353187f $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_271 N_A_278_409#_c_265_n N_A_461_55#_c_462_n 0.00187393f $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_272 N_A_278_409#_M1003_g N_A_461_55#_c_463_n 0.00501569f $X=2.665 $Y=0.485
+ $X2=0 $Y2=0
cc_273 N_A_278_409#_c_260_n N_A_461_55#_c_463_n 0.0121096f $X=1.725 $Y=0.91
+ $X2=0 $Y2=0
cc_274 N_A_278_409#_c_262_n N_A_461_55#_c_463_n 6.8158e-19 $X=1.89 $Y=0.495
+ $X2=0 $Y2=0
cc_275 N_A_278_409#_M1019_g N_A_461_55#_c_470_n 0.00732296f $X=2.85 $Y=2.195
+ $X2=0 $Y2=0
cc_276 N_A_278_409#_c_269_n N_A_461_55#_c_470_n 0.0301328f $X=2.93 $Y=2.27 $X2=0
+ $Y2=0
cc_277 N_A_278_409#_c_263_n N_A_461_55#_c_470_n 0.00620491f $X=3.015 $Y=1.755
+ $X2=0 $Y2=0
cc_278 N_A_278_409#_c_301_p N_A_461_55#_c_470_n 0.0175175f $X=3.015 $Y=2.185
+ $X2=0 $Y2=0
cc_279 N_A_278_409#_c_266_n N_A_461_55#_c_470_n 0.005925f $X=3.025 $Y=1.33 $X2=0
+ $Y2=0
cc_280 N_A_278_409#_M1003_g N_A_461_55#_c_464_n 0.0115506f $X=2.665 $Y=0.485
+ $X2=0 $Y2=0
cc_281 N_A_278_409#_M1020_g N_A_461_55#_c_464_n 0.0111604f $X=3.025 $Y=0.485
+ $X2=0 $Y2=0
cc_282 N_A_278_409#_c_263_n N_A_461_55#_c_464_n 0.024016f $X=3.015 $Y=1.755
+ $X2=0 $Y2=0
cc_283 N_A_278_409#_c_264_n N_A_461_55#_c_464_n 0.0250608f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_284 N_A_278_409#_c_266_n N_A_461_55#_c_464_n 2.06137e-19 $X=3.025 $Y=1.33
+ $X2=0 $Y2=0
cc_285 N_A_278_409#_M1009_g N_A_461_55#_c_465_n 2.71649e-19 $X=3.95 $Y=2.465
+ $X2=0 $Y2=0
cc_286 N_A_278_409#_c_264_n N_A_461_55#_c_465_n 0.0176617f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_287 N_A_278_409#_c_265_n N_A_461_55#_c_465_n 0.00521414f $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_288 N_A_278_409#_M1009_g N_A_461_55#_c_466_n 0.0216431f $X=3.95 $Y=2.465
+ $X2=0 $Y2=0
cc_289 N_A_278_409#_c_264_n N_A_461_55#_c_466_n 2.37597e-19 $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_290 N_A_278_409#_c_265_n N_A_461_55#_c_466_n 0.0101946f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_291 N_A_278_409#_M1013_g N_A_461_55#_c_467_n 0.0165141f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_292 N_A_278_409#_M1013_g N_A_934_29#_c_555_n 0.0428785f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_293 N_A_278_409#_M1013_g N_A_784_55#_c_728_n 0.0110542f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_294 N_A_278_409#_M1009_g N_A_784_55#_c_724_n 0.00196492f $X=3.95 $Y=2.465
+ $X2=0 $Y2=0
cc_295 N_A_278_409#_M1009_g N_A_784_55#_c_725_n 0.00780962f $X=3.95 $Y=2.465
+ $X2=0 $Y2=0
cc_296 N_A_278_409#_c_264_n N_A_784_55#_c_725_n 0.00186167f $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_297 N_A_278_409#_c_265_n N_A_784_55#_c_725_n 0.0074659f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_298 N_A_278_409#_M1013_g N_A_784_55#_c_714_n 0.0024343f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_299 N_A_278_409#_M1013_g N_A_784_55#_c_716_n 0.00113259f $X=4.355 $Y=0.485
+ $X2=0 $Y2=0
cc_300 N_A_278_409#_c_269_n N_VPWR_M1019_d 0.0032149f $X=2.93 $Y=2.27 $X2=0
+ $Y2=0
cc_301 N_A_278_409#_c_301_p N_VPWR_M1019_d 0.00524546f $X=3.015 $Y=2.185 $X2=0
+ $Y2=0
cc_302 N_A_278_409#_c_264_n N_VPWR_M1019_d 0.00527295f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_303 N_A_278_409#_M1019_g N_VPWR_c_873_n 0.00465843f $X=2.85 $Y=2.195 $X2=0
+ $Y2=0
cc_304 N_A_278_409#_M1009_g N_VPWR_c_873_n 0.00244298f $X=3.95 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_278_409#_c_269_n N_VPWR_c_873_n 0.00587285f $X=2.93 $Y=2.27 $X2=0
+ $Y2=0
cc_306 N_A_278_409#_M1009_g N_VPWR_c_881_n 0.00775913f $X=3.95 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_278_409#_M1019_g N_VPWR_c_871_n 0.00156346f $X=2.85 $Y=2.195 $X2=0
+ $Y2=0
cc_308 N_A_278_409#_M1009_g N_VPWR_c_871_n 0.0152633f $X=3.95 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_278_409#_c_262_n N_VGND_c_1017_n 0.00639517f $X=1.89 $Y=0.495 $X2=0
+ $Y2=0
cc_310 N_A_278_409#_M1003_g N_VGND_c_1018_n 0.00511657f $X=2.665 $Y=0.485 $X2=0
+ $Y2=0
cc_311 N_A_278_409#_M1020_g N_VGND_c_1018_n 0.00452967f $X=3.025 $Y=0.485 $X2=0
+ $Y2=0
cc_312 N_A_278_409#_c_262_n N_VGND_c_1018_n 0.0220321f $X=1.89 $Y=0.495 $X2=0
+ $Y2=0
cc_313 N_A_278_409#_M1003_g N_VGND_c_1019_n 0.00195145f $X=2.665 $Y=0.485 $X2=0
+ $Y2=0
cc_314 N_A_278_409#_M1020_g N_VGND_c_1019_n 0.0108855f $X=3.025 $Y=0.485 $X2=0
+ $Y2=0
cc_315 N_A_278_409#_M1013_g N_VGND_c_1026_n 0.00346579f $X=4.355 $Y=0.485 $X2=0
+ $Y2=0
cc_316 N_A_278_409#_M1003_g N_VGND_c_1029_n 0.00669497f $X=2.665 $Y=0.485 $X2=0
+ $Y2=0
cc_317 N_A_278_409#_M1020_g N_VGND_c_1029_n 0.00421151f $X=3.025 $Y=0.485 $X2=0
+ $Y2=0
cc_318 N_A_278_409#_M1013_g N_VGND_c_1029_n 0.00512297f $X=4.355 $Y=0.485 $X2=0
+ $Y2=0
cc_319 N_A_278_409#_c_260_n N_VGND_c_1029_n 0.0109451f $X=1.725 $Y=0.91 $X2=0
+ $Y2=0
cc_320 N_A_278_409#_c_261_n N_VGND_c_1029_n 0.00498505f $X=1.385 $Y=0.91 $X2=0
+ $Y2=0
cc_321 N_A_278_409#_c_262_n N_VGND_c_1029_n 0.0125808f $X=1.89 $Y=0.495 $X2=0
+ $Y2=0
cc_322 N_A_27_57#_M1006_g N_A_461_55#_c_460_n 0.00104945f $X=3.455 $Y=0.485
+ $X2=0 $Y2=0
cc_323 N_A_27_57#_M1006_g N_A_461_55#_c_461_n 0.0205198f $X=3.455 $Y=0.485 $X2=0
+ $Y2=0
cc_324 N_A_27_57#_M1006_g N_A_461_55#_c_464_n 0.0125143f $X=3.455 $Y=0.485 $X2=0
+ $Y2=0
cc_325 N_A_27_57#_M1006_g N_A_461_55#_c_467_n 0.0360354f $X=3.455 $Y=0.485 $X2=0
+ $Y2=0
cc_326 N_A_27_57#_c_392_n N_VPWR_M1018_d 0.0165839f $X=1.95 $Y=2.62 $X2=-0.19
+ $Y2=-0.245
cc_327 N_A_27_57#_c_392_n N_VPWR_c_872_n 0.0235397f $X=1.95 $Y=2.62 $X2=0 $Y2=0
cc_328 N_A_27_57#_c_397_n N_VPWR_c_872_n 0.00515182f $X=0.295 $Y=2.62 $X2=0
+ $Y2=0
cc_329 N_A_27_57#_c_387_n N_VPWR_c_873_n 0.0226195f $X=3.335 $Y=3.14 $X2=0 $Y2=0
cc_330 N_A_27_57#_M1027_g N_VPWR_c_873_n 0.0142226f $X=3.46 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A_27_57#_c_392_n N_VPWR_c_878_n 0.00430381f $X=1.95 $Y=2.62 $X2=0 $Y2=0
cc_332 N_A_27_57#_c_397_n N_VPWR_c_878_n 0.0240548f $X=0.295 $Y=2.62 $X2=0 $Y2=0
cc_333 N_A_27_57#_c_392_n N_VPWR_c_880_n 0.0144799f $X=1.95 $Y=2.62 $X2=0 $Y2=0
cc_334 N_A_27_57#_c_393_n N_VPWR_c_880_n 0.0206075f $X=2.115 $Y=2.9 $X2=0 $Y2=0
cc_335 N_A_27_57#_c_394_n N_VPWR_c_880_n 0.0337647f $X=2.115 $Y=2.9 $X2=0 $Y2=0
cc_336 N_A_27_57#_c_387_n N_VPWR_c_881_n 0.00860995f $X=3.335 $Y=3.14 $X2=0
+ $Y2=0
cc_337 N_A_27_57#_c_387_n N_VPWR_c_871_n 0.0517061f $X=3.335 $Y=3.14 $X2=0 $Y2=0
cc_338 N_A_27_57#_c_392_n N_VPWR_c_871_n 0.0322043f $X=1.95 $Y=2.62 $X2=0 $Y2=0
cc_339 N_A_27_57#_c_393_n N_VPWR_c_871_n 0.0110969f $X=2.115 $Y=2.9 $X2=0 $Y2=0
cc_340 N_A_27_57#_c_394_n N_VPWR_c_871_n 0.00943448f $X=2.115 $Y=2.9 $X2=0 $Y2=0
cc_341 N_A_27_57#_c_397_n N_VPWR_c_871_n 0.0137416f $X=0.295 $Y=2.62 $X2=0 $Y2=0
cc_342 N_A_27_57#_c_385_n N_VGND_c_1017_n 0.0127138f $X=0.28 $Y=0.495 $X2=0
+ $Y2=0
cc_343 N_A_27_57#_M1006_g N_VGND_c_1019_n 0.0115826f $X=3.455 $Y=0.485 $X2=0
+ $Y2=0
cc_344 N_A_27_57#_c_385_n N_VGND_c_1025_n 0.0217285f $X=0.28 $Y=0.495 $X2=0
+ $Y2=0
cc_345 N_A_27_57#_M1006_g N_VGND_c_1026_n 0.00452967f $X=3.455 $Y=0.485 $X2=0
+ $Y2=0
cc_346 N_A_27_57#_M1006_g N_VGND_c_1029_n 0.00430406f $X=3.455 $Y=0.485 $X2=0
+ $Y2=0
cc_347 N_A_27_57#_c_385_n N_VGND_c_1029_n 0.0125175f $X=0.28 $Y=0.495 $X2=0
+ $Y2=0
cc_348 N_A_461_55#_c_459_n N_A_934_29#_c_557_n 7.78137e-19 $X=4.335 $Y=0.98
+ $X2=0 $Y2=0
cc_349 N_A_461_55#_c_465_n N_A_934_29#_c_557_n 2.29287e-19 $X=4.42 $Y=1.64 $X2=0
+ $Y2=0
cc_350 N_A_461_55#_c_466_n N_A_934_29#_c_557_n 0.00466167f $X=4.805 $Y=1.64
+ $X2=0 $Y2=0
cc_351 N_A_461_55#_M1016_g N_A_934_29#_M1001_g 0.047491f $X=4.765 $Y=2.465 $X2=0
+ $Y2=0
cc_352 N_A_461_55#_c_465_n N_A_934_29#_c_573_n 3.57021e-19 $X=4.42 $Y=1.64 $X2=0
+ $Y2=0
cc_353 N_A_461_55#_c_466_n N_A_934_29#_c_573_n 0.0174432f $X=4.805 $Y=1.64 $X2=0
+ $Y2=0
cc_354 N_A_461_55#_c_459_n N_A_784_55#_c_728_n 0.0348683f $X=4.335 $Y=0.98 $X2=0
+ $Y2=0
cc_355 N_A_461_55#_c_461_n N_A_784_55#_c_728_n 0.00214119f $X=3.905 $Y=0.98
+ $X2=0 $Y2=0
cc_356 N_A_461_55#_M1016_g N_A_784_55#_c_725_n 0.0231812f $X=4.765 $Y=2.465
+ $X2=0 $Y2=0
cc_357 N_A_461_55#_c_465_n N_A_784_55#_c_725_n 0.0078057f $X=4.42 $Y=1.64 $X2=0
+ $Y2=0
cc_358 N_A_461_55#_M1016_g N_A_784_55#_c_726_n 0.0226744f $X=4.765 $Y=2.465
+ $X2=0 $Y2=0
cc_359 N_A_461_55#_c_459_n N_A_784_55#_c_714_n 0.0247041f $X=4.335 $Y=0.98 $X2=0
+ $Y2=0
cc_360 N_A_461_55#_c_465_n N_A_784_55#_c_715_n 0.00755775f $X=4.42 $Y=1.64 $X2=0
+ $Y2=0
cc_361 N_A_461_55#_c_466_n N_A_784_55#_c_715_n 6.48665e-19 $X=4.805 $Y=1.64
+ $X2=0 $Y2=0
cc_362 N_A_461_55#_c_459_n N_A_784_55#_c_716_n 0.00179882f $X=4.335 $Y=0.98
+ $X2=0 $Y2=0
cc_363 N_A_461_55#_c_462_n N_A_784_55#_c_716_n 0.0121277f $X=4.42 $Y=1.475 $X2=0
+ $Y2=0
cc_364 N_A_461_55#_c_465_n N_A_784_55#_c_716_n 0.013796f $X=4.42 $Y=1.64 $X2=0
+ $Y2=0
cc_365 N_A_461_55#_c_466_n N_A_784_55#_c_716_n 8.0922e-19 $X=4.805 $Y=1.64 $X2=0
+ $Y2=0
cc_366 N_A_461_55#_M1016_g N_A_784_55#_c_717_n 0.0197162f $X=4.765 $Y=2.465
+ $X2=0 $Y2=0
cc_367 N_A_461_55#_c_462_n N_A_784_55#_c_717_n 0.00538096f $X=4.42 $Y=1.475
+ $X2=0 $Y2=0
cc_368 N_A_461_55#_c_465_n N_A_784_55#_c_717_n 0.0244649f $X=4.42 $Y=1.64 $X2=0
+ $Y2=0
cc_369 N_A_461_55#_c_466_n N_A_784_55#_c_717_n 0.00190737f $X=4.805 $Y=1.64
+ $X2=0 $Y2=0
cc_370 N_A_461_55#_M1016_g N_VPWR_c_881_n 0.00489539f $X=4.765 $Y=2.465 $X2=0
+ $Y2=0
cc_371 N_A_461_55#_M1016_g N_VPWR_c_871_n 0.00609976f $X=4.765 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_A_461_55#_c_457_n N_VGND_c_1018_n 0.022078f $X=2.45 $Y=0.49 $X2=0 $Y2=0
cc_373 N_A_461_55#_c_457_n N_VGND_c_1019_n 0.0123792f $X=2.45 $Y=0.49 $X2=0
+ $Y2=0
cc_374 N_A_461_55#_c_464_n N_VGND_c_1019_n 0.0200517f $X=3.74 $Y=0.98 $X2=0
+ $Y2=0
cc_375 N_A_461_55#_c_467_n N_VGND_c_1019_n 0.00214415f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_376 N_A_461_55#_c_467_n N_VGND_c_1026_n 0.00545548f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_377 N_A_461_55#_c_457_n N_VGND_c_1029_n 0.0125905f $X=2.45 $Y=0.49 $X2=0
+ $Y2=0
cc_378 N_A_461_55#_c_461_n N_VGND_c_1029_n 0.00195629f $X=3.905 $Y=0.98 $X2=0
+ $Y2=0
cc_379 N_A_461_55#_c_464_n N_VGND_c_1029_n 0.0344617f $X=3.74 $Y=0.98 $X2=0
+ $Y2=0
cc_380 N_A_461_55#_c_467_n N_VGND_c_1029_n 0.00613009f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_381 N_A_934_29#_c_569_n N_A_784_55#_c_708_n 0.00252788f $X=6.31 $Y=0.49 $X2=0
+ $Y2=0
cc_382 N_A_934_29#_c_556_n N_A_784_55#_c_710_n 0.00881671f $X=5.21 $Y=0.845
+ $X2=0 $Y2=0
cc_383 N_A_934_29#_c_573_n N_A_784_55#_c_710_n 0.00243377f $X=5.645 $Y=1.64
+ $X2=0 $Y2=0
cc_384 N_A_934_29#_c_569_n N_A_784_55#_c_711_n 0.0112001f $X=6.31 $Y=0.49 $X2=0
+ $Y2=0
cc_385 N_A_934_29#_c_558_n N_A_784_55#_M1023_g 4.34875e-19 $X=5.285 $Y=1.475
+ $X2=0 $Y2=0
cc_386 N_A_934_29#_M1001_g N_A_784_55#_M1023_g 0.0142852f $X=5.335 $Y=2.465
+ $X2=0 $Y2=0
cc_387 N_A_934_29#_c_577_n N_A_784_55#_M1023_g 0.0183235f $X=6.275 $Y=1.72 $X2=0
+ $Y2=0
cc_388 N_A_934_29#_c_570_n N_A_784_55#_M1023_g 0.0074988f $X=6.44 $Y=1.805 $X2=0
+ $Y2=0
cc_389 N_A_934_29#_c_579_n N_A_784_55#_M1023_g 0.0317972f $X=6.44 $Y=2.11 $X2=0
+ $Y2=0
cc_390 N_A_934_29#_c_571_n N_A_784_55#_M1023_g 0.00453004f $X=6.755 $Y=1.06
+ $X2=0 $Y2=0
cc_391 N_A_934_29#_c_572_n N_A_784_55#_M1023_g 0.00120267f $X=5.645 $Y=1.64
+ $X2=0 $Y2=0
cc_392 N_A_934_29#_c_573_n N_A_784_55#_M1023_g 0.019118f $X=5.645 $Y=1.64 $X2=0
+ $Y2=0
cc_393 N_A_934_29#_c_561_n N_A_784_55#_c_713_n 0.00357855f $X=7.16 $Y=0.97 $X2=0
+ $Y2=0
cc_394 N_A_934_29#_c_568_n N_A_784_55#_c_713_n 0.010523f $X=6.31 $Y=0.775 $X2=0
+ $Y2=0
cc_395 N_A_934_29#_c_555_n N_A_784_55#_c_728_n 0.013914f $X=4.745 $Y=0.77 $X2=0
+ $Y2=0
cc_396 N_A_934_29#_M1001_g N_A_784_55#_c_726_n 0.00637711f $X=5.335 $Y=2.465
+ $X2=0 $Y2=0
cc_397 N_A_934_29#_c_555_n N_A_784_55#_c_714_n 0.00529334f $X=4.745 $Y=0.77
+ $X2=0 $Y2=0
cc_398 N_A_934_29#_c_556_n N_A_784_55#_c_714_n 0.00799955f $X=5.21 $Y=0.845
+ $X2=0 $Y2=0
cc_399 N_A_934_29#_c_557_n N_A_784_55#_c_714_n 0.0051652f $X=4.82 $Y=0.845 $X2=0
+ $Y2=0
cc_400 N_A_934_29#_c_558_n N_A_784_55#_c_714_n 0.00573729f $X=5.285 $Y=1.475
+ $X2=0 $Y2=0
cc_401 N_A_934_29#_c_556_n N_A_784_55#_c_715_n 0.00687778f $X=5.21 $Y=0.845
+ $X2=0 $Y2=0
cc_402 N_A_934_29#_c_558_n N_A_784_55#_c_717_n 0.0110276f $X=5.285 $Y=1.475
+ $X2=0 $Y2=0
cc_403 N_A_934_29#_M1001_g N_A_784_55#_c_717_n 0.0301596f $X=5.335 $Y=2.465
+ $X2=0 $Y2=0
cc_404 N_A_934_29#_c_572_n N_A_784_55#_c_717_n 0.0224548f $X=5.645 $Y=1.64 $X2=0
+ $Y2=0
cc_405 N_A_934_29#_c_573_n N_A_784_55#_c_717_n 0.00910337f $X=5.645 $Y=1.64
+ $X2=0 $Y2=0
cc_406 N_A_934_29#_c_558_n N_A_784_55#_c_718_n 0.00725836f $X=5.285 $Y=1.475
+ $X2=0 $Y2=0
cc_407 N_A_934_29#_c_577_n N_A_784_55#_c_718_n 0.00979f $X=6.275 $Y=1.72 $X2=0
+ $Y2=0
cc_408 N_A_934_29#_c_572_n N_A_784_55#_c_718_n 0.0229991f $X=5.645 $Y=1.64 $X2=0
+ $Y2=0
cc_409 N_A_934_29#_c_573_n N_A_784_55#_c_718_n 0.00701693f $X=5.645 $Y=1.64
+ $X2=0 $Y2=0
cc_410 N_A_934_29#_c_556_n N_A_784_55#_c_719_n 0.00156115f $X=5.21 $Y=0.845
+ $X2=0 $Y2=0
cc_411 N_A_934_29#_c_558_n N_A_784_55#_c_719_n 0.00735642f $X=5.285 $Y=1.475
+ $X2=0 $Y2=0
cc_412 N_A_934_29#_c_558_n N_A_784_55#_c_720_n 8.57445e-19 $X=5.285 $Y=1.475
+ $X2=0 $Y2=0
cc_413 N_A_934_29#_c_577_n N_A_784_55#_c_720_n 0.017489f $X=6.275 $Y=1.72 $X2=0
+ $Y2=0
cc_414 N_A_934_29#_c_568_n N_A_784_55#_c_720_n 0.0164415f $X=6.31 $Y=0.775 $X2=0
+ $Y2=0
cc_415 N_A_934_29#_c_570_n N_A_784_55#_c_720_n 0.00903689f $X=6.44 $Y=1.805
+ $X2=0 $Y2=0
cc_416 N_A_934_29#_c_625_p N_A_784_55#_c_720_n 0.0156384f $X=6.755 $Y=1.06 $X2=0
+ $Y2=0
cc_417 N_A_934_29#_c_571_n N_A_784_55#_c_720_n 0.00108275f $X=6.755 $Y=1.06
+ $X2=0 $Y2=0
cc_418 N_A_934_29#_c_568_n N_A_784_55#_c_721_n 0.00138706f $X=6.31 $Y=0.775
+ $X2=0 $Y2=0
cc_419 N_A_934_29#_c_570_n N_A_784_55#_c_721_n 5.87723e-19 $X=6.44 $Y=1.805
+ $X2=0 $Y2=0
cc_420 N_A_934_29#_c_625_p N_A_784_55#_c_721_n 0.00101176f $X=6.755 $Y=1.06
+ $X2=0 $Y2=0
cc_421 N_A_934_29#_c_571_n N_A_784_55#_c_721_n 0.0171714f $X=6.755 $Y=1.06 $X2=0
+ $Y2=0
cc_422 N_A_934_29#_c_558_n N_A_784_55#_c_722_n 0.00974614f $X=5.285 $Y=1.475
+ $X2=0 $Y2=0
cc_423 N_A_934_29#_c_568_n N_A_784_55#_c_722_n 0.00186868f $X=6.31 $Y=0.775
+ $X2=0 $Y2=0
cc_424 N_A_934_29#_c_625_p N_A_784_55#_c_722_n 0.00101104f $X=6.755 $Y=1.06
+ $X2=0 $Y2=0
cc_425 N_A_934_29#_c_571_n N_A_784_55#_c_722_n 0.00357855f $X=6.755 $Y=1.06
+ $X2=0 $Y2=0
cc_426 N_A_934_29#_M1010_g N_A_1662_57#_c_823_n 0.00233827f $X=7.655 $Y=2.335
+ $X2=0 $Y2=0
cc_427 N_A_934_29#_M1004_g N_A_1662_57#_c_823_n 0.00209968f $X=7.875 $Y=0.495
+ $X2=0 $Y2=0
cc_428 N_A_934_29#_M1026_g N_A_1662_57#_c_823_n 0.0196053f $X=8.185 $Y=2.335
+ $X2=0 $Y2=0
cc_429 N_A_934_29#_M1008_g N_A_1662_57#_c_823_n 0.0152804f $X=8.235 $Y=0.495
+ $X2=0 $Y2=0
cc_430 N_A_934_29#_c_567_n N_A_1662_57#_c_823_n 0.0105303f $X=8.235 $Y=0.97
+ $X2=0 $Y2=0
cc_431 N_A_934_29#_M1010_g N_A_1662_57#_c_829_n 5.13349e-19 $X=7.655 $Y=2.335
+ $X2=0 $Y2=0
cc_432 N_A_934_29#_M1026_g N_A_1662_57#_c_829_n 0.0206848f $X=8.185 $Y=2.335
+ $X2=0 $Y2=0
cc_433 N_A_934_29#_M1026_g N_A_1662_57#_c_825_n 4.25713e-19 $X=8.185 $Y=2.335
+ $X2=0 $Y2=0
cc_434 N_A_934_29#_M1010_g N_A_1662_57#_c_826_n 7.25172e-19 $X=7.655 $Y=2.335
+ $X2=0 $Y2=0
cc_435 N_A_934_29#_M1026_g N_A_1662_57#_c_826_n 0.00693094f $X=8.185 $Y=2.335
+ $X2=0 $Y2=0
cc_436 N_A_934_29#_M1026_g N_A_1662_57#_c_827_n 0.0107927f $X=8.185 $Y=2.335
+ $X2=0 $Y2=0
cc_437 N_A_934_29#_M1001_g N_VPWR_c_874_n 0.00636755f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_438 N_A_934_29#_c_577_n N_VPWR_c_874_n 7.13784e-19 $X=6.275 $Y=1.72 $X2=0
+ $Y2=0
cc_439 N_A_934_29#_c_579_n N_VPWR_c_874_n 0.0362821f $X=6.44 $Y=2.11 $X2=0 $Y2=0
cc_440 N_A_934_29#_c_572_n N_VPWR_c_874_n 0.0241194f $X=5.645 $Y=1.64 $X2=0
+ $Y2=0
cc_441 N_A_934_29#_c_573_n N_VPWR_c_874_n 0.00241669f $X=5.645 $Y=1.64 $X2=0
+ $Y2=0
cc_442 N_A_934_29#_M1010_g N_VPWR_c_875_n 0.0257154f $X=7.655 $Y=2.335 $X2=0
+ $Y2=0
cc_443 N_A_934_29#_M1026_g N_VPWR_c_875_n 0.0266623f $X=8.185 $Y=2.335 $X2=0
+ $Y2=0
cc_444 N_A_934_29#_M1026_g N_VPWR_c_876_n 0.00714707f $X=8.185 $Y=2.335 $X2=0
+ $Y2=0
cc_445 N_A_934_29#_M1026_g N_VPWR_c_877_n 0.00442745f $X=8.185 $Y=2.335 $X2=0
+ $Y2=0
cc_446 N_A_934_29#_M1001_g N_VPWR_c_881_n 0.00661271f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_934_29#_M1010_g N_VPWR_c_882_n 0.00714193f $X=7.655 $Y=2.335 $X2=0
+ $Y2=0
cc_448 N_A_934_29#_c_579_n N_VPWR_c_882_n 0.0148628f $X=6.44 $Y=2.11 $X2=0 $Y2=0
cc_449 N_A_934_29#_M1001_g N_VPWR_c_871_n 0.0115781f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_934_29#_M1010_g N_VPWR_c_871_n 0.00763694f $X=7.655 $Y=2.335 $X2=0
+ $Y2=0
cc_451 N_A_934_29#_M1026_g N_VPWR_c_871_n 0.00763694f $X=8.185 $Y=2.335 $X2=0
+ $Y2=0
cc_452 N_A_934_29#_c_579_n N_VPWR_c_871_n 0.0120349f $X=6.44 $Y=2.11 $X2=0 $Y2=0
cc_453 N_A_934_29#_M1002_g N_Q_c_963_n 0.0115698f $X=7.085 $Y=0.495 $X2=0 $Y2=0
cc_454 N_A_934_29#_c_561_n N_Q_c_963_n 0.00383731f $X=7.16 $Y=0.97 $X2=0 $Y2=0
cc_455 N_A_934_29#_M1025_g N_Q_c_963_n 0.0023972f $X=7.445 $Y=0.495 $X2=0 $Y2=0
cc_456 N_A_934_29#_c_568_n N_Q_c_963_n 0.0129349f $X=6.31 $Y=0.775 $X2=0 $Y2=0
cc_457 N_A_934_29#_c_569_n N_Q_c_963_n 0.0231249f $X=6.31 $Y=0.49 $X2=0 $Y2=0
cc_458 N_A_934_29#_c_560_n Q 0.00844283f $X=7.37 $Y=0.97 $X2=0 $Y2=0
cc_459 N_A_934_29#_M1010_g Q 0.00938698f $X=7.655 $Y=2.335 $X2=0 $Y2=0
cc_460 N_A_934_29#_M1026_g Q 0.00271826f $X=8.185 $Y=2.335 $X2=0 $Y2=0
cc_461 N_A_934_29#_c_570_n Q 0.0128544f $X=6.44 $Y=1.805 $X2=0 $Y2=0
cc_462 N_A_934_29#_c_571_n Q 7.57529e-19 $X=6.755 $Y=1.06 $X2=0 $Y2=0
cc_463 N_A_934_29#_M1010_g Q 0.0368858f $X=7.655 $Y=2.335 $X2=0 $Y2=0
cc_464 N_A_934_29#_M1026_g Q 2.9786e-19 $X=8.185 $Y=2.335 $X2=0 $Y2=0
cc_465 N_A_934_29#_c_570_n Q 0.0130446f $X=6.44 $Y=1.805 $X2=0 $Y2=0
cc_466 N_A_934_29#_c_579_n Q 0.0441897f $X=6.44 $Y=2.11 $X2=0 $Y2=0
cc_467 N_A_934_29#_M1002_g N_Q_c_966_n 0.00774429f $X=7.085 $Y=0.495 $X2=0 $Y2=0
cc_468 N_A_934_29#_c_560_n N_Q_c_966_n 0.0113004f $X=7.37 $Y=0.97 $X2=0 $Y2=0
cc_469 N_A_934_29#_c_561_n N_Q_c_966_n 0.004429f $X=7.16 $Y=0.97 $X2=0 $Y2=0
cc_470 N_A_934_29#_M1025_g N_Q_c_966_n 0.00448731f $X=7.445 $Y=0.495 $X2=0 $Y2=0
cc_471 N_A_934_29#_M1010_g N_Q_c_966_n 0.00293349f $X=7.655 $Y=2.335 $X2=0 $Y2=0
cc_472 N_A_934_29#_c_568_n N_Q_c_966_n 0.00935757f $X=6.31 $Y=0.775 $X2=0 $Y2=0
cc_473 N_A_934_29#_c_569_n N_Q_c_966_n 0.00506326f $X=6.31 $Y=0.49 $X2=0 $Y2=0
cc_474 N_A_934_29#_c_625_p N_Q_c_966_n 0.0335126f $X=6.755 $Y=1.06 $X2=0 $Y2=0
cc_475 N_A_934_29#_c_571_n N_Q_c_966_n 0.00360799f $X=6.755 $Y=1.06 $X2=0 $Y2=0
cc_476 N_A_934_29#_c_555_n N_VGND_c_1020_n 0.00837488f $X=4.745 $Y=0.77 $X2=0
+ $Y2=0
cc_477 N_A_934_29#_c_556_n N_VGND_c_1020_n 0.0101433f $X=5.21 $Y=0.845 $X2=0
+ $Y2=0
cc_478 N_A_934_29#_M1002_g N_VGND_c_1021_n 0.00126149f $X=7.085 $Y=0.495 $X2=0
+ $Y2=0
cc_479 N_A_934_29#_M1025_g N_VGND_c_1021_n 0.0106321f $X=7.445 $Y=0.495 $X2=0
+ $Y2=0
cc_480 N_A_934_29#_M1004_g N_VGND_c_1021_n 0.0134712f $X=7.875 $Y=0.495 $X2=0
+ $Y2=0
cc_481 N_A_934_29#_M1008_g N_VGND_c_1021_n 0.002112f $X=8.235 $Y=0.495 $X2=0
+ $Y2=0
cc_482 N_A_934_29#_c_567_n N_VGND_c_1021_n 0.00483855f $X=8.235 $Y=0.97 $X2=0
+ $Y2=0
cc_483 N_A_934_29#_M1008_g N_VGND_c_1022_n 0.00347989f $X=8.235 $Y=0.495 $X2=0
+ $Y2=0
cc_484 N_A_934_29#_M1002_g N_VGND_c_1023_n 0.00327653f $X=7.085 $Y=0.495 $X2=0
+ $Y2=0
cc_485 N_A_934_29#_M1025_g N_VGND_c_1023_n 0.00445056f $X=7.445 $Y=0.495 $X2=0
+ $Y2=0
cc_486 N_A_934_29#_c_569_n N_VGND_c_1023_n 0.0220321f $X=6.31 $Y=0.49 $X2=0
+ $Y2=0
cc_487 N_A_934_29#_c_555_n N_VGND_c_1026_n 0.00346421f $X=4.745 $Y=0.77 $X2=0
+ $Y2=0
cc_488 N_A_934_29#_c_556_n N_VGND_c_1026_n 0.0028667f $X=5.21 $Y=0.845 $X2=0
+ $Y2=0
cc_489 N_A_934_29#_M1004_g N_VGND_c_1027_n 0.00445056f $X=7.875 $Y=0.495 $X2=0
+ $Y2=0
cc_490 N_A_934_29#_M1008_g N_VGND_c_1027_n 0.00502664f $X=8.235 $Y=0.495 $X2=0
+ $Y2=0
cc_491 N_A_934_29#_c_555_n N_VGND_c_1029_n 0.0059633f $X=4.745 $Y=0.77 $X2=0
+ $Y2=0
cc_492 N_A_934_29#_c_556_n N_VGND_c_1029_n 0.00385076f $X=5.21 $Y=0.845 $X2=0
+ $Y2=0
cc_493 N_A_934_29#_M1002_g N_VGND_c_1029_n 0.00563487f $X=7.085 $Y=0.495 $X2=0
+ $Y2=0
cc_494 N_A_934_29#_M1025_g N_VGND_c_1029_n 0.00796275f $X=7.445 $Y=0.495 $X2=0
+ $Y2=0
cc_495 N_A_934_29#_M1004_g N_VGND_c_1029_n 0.00796275f $X=7.875 $Y=0.495 $X2=0
+ $Y2=0
cc_496 N_A_934_29#_M1008_g N_VGND_c_1029_n 0.010303f $X=8.235 $Y=0.495 $X2=0
+ $Y2=0
cc_497 N_A_934_29#_c_568_n N_VGND_c_1029_n 0.00913902f $X=6.31 $Y=0.775 $X2=0
+ $Y2=0
cc_498 N_A_934_29#_c_569_n N_VGND_c_1029_n 0.0125808f $X=6.31 $Y=0.49 $X2=0
+ $Y2=0
cc_499 N_A_784_55#_M1023_g N_VPWR_c_874_n 0.0144727f $X=6.175 $Y=2.465 $X2=0
+ $Y2=0
cc_500 N_A_784_55#_c_726_n N_VPWR_c_874_n 0.00760059f $X=5.14 $Y=2.9 $X2=0 $Y2=0
cc_501 N_A_784_55#_c_724_n N_VPWR_c_881_n 0.0150262f $X=4.295 $Y=2.815 $X2=0
+ $Y2=0
cc_502 N_A_784_55#_c_726_n N_VPWR_c_881_n 0.0347328f $X=5.14 $Y=2.9 $X2=0 $Y2=0
cc_503 N_A_784_55#_M1023_g N_VPWR_c_882_n 0.00748399f $X=6.175 $Y=2.465 $X2=0
+ $Y2=0
cc_504 N_A_784_55#_M1023_g N_VPWR_c_871_n 0.014492f $X=6.175 $Y=2.465 $X2=0
+ $Y2=0
cc_505 N_A_784_55#_c_724_n N_VPWR_c_871_n 0.0122245f $X=4.295 $Y=2.815 $X2=0
+ $Y2=0
cc_506 N_A_784_55#_c_726_n N_VPWR_c_871_n 0.028733f $X=5.14 $Y=2.9 $X2=0 $Y2=0
cc_507 N_A_784_55#_c_726_n A_978_393# 0.00732587f $X=5.14 $Y=2.9 $X2=-0.19
+ $Y2=-0.245
cc_508 N_A_784_55#_c_717_n A_978_393# 0.0104592f $X=5.225 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_509 N_A_784_55#_c_711_n N_Q_c_963_n 7.06601e-19 $X=6.095 $Y=0.77 $X2=0 $Y2=0
cc_510 N_A_784_55#_c_708_n N_VGND_c_1020_n 0.0175225f $X=5.735 $Y=0.77 $X2=0
+ $Y2=0
cc_511 N_A_784_55#_c_714_n N_VGND_c_1020_n 0.00379276f $X=4.77 $Y=1.125 $X2=0
+ $Y2=0
cc_512 N_A_784_55#_c_715_n N_VGND_c_1020_n 0.00472534f $X=5.14 $Y=1.21 $X2=0
+ $Y2=0
cc_513 N_A_784_55#_c_718_n N_VGND_c_1020_n 0.00226042f $X=6.02 $Y=1.21 $X2=0
+ $Y2=0
cc_514 N_A_784_55#_c_719_n N_VGND_c_1020_n 0.00812704f $X=5.225 $Y=1.21 $X2=0
+ $Y2=0
cc_515 N_A_784_55#_c_708_n N_VGND_c_1023_n 0.00545548f $X=5.735 $Y=0.77 $X2=0
+ $Y2=0
cc_516 N_A_784_55#_c_709_n N_VGND_c_1023_n 4.63617e-19 $X=6.02 $Y=0.845 $X2=0
+ $Y2=0
cc_517 N_A_784_55#_c_711_n N_VGND_c_1023_n 0.00511657f $X=6.095 $Y=0.77 $X2=0
+ $Y2=0
cc_518 N_A_784_55#_c_728_n N_VGND_c_1026_n 0.0340901f $X=4.685 $Y=0.485 $X2=0
+ $Y2=0
cc_519 N_A_784_55#_c_708_n N_VGND_c_1029_n 0.0113884f $X=5.735 $Y=0.77 $X2=0
+ $Y2=0
cc_520 N_A_784_55#_c_709_n N_VGND_c_1029_n 6.36806e-19 $X=6.02 $Y=0.845 $X2=0
+ $Y2=0
cc_521 N_A_784_55#_c_711_n N_VGND_c_1029_n 0.0104992f $X=6.095 $Y=0.77 $X2=0
+ $Y2=0
cc_522 N_A_784_55#_c_728_n N_VGND_c_1029_n 0.0306474f $X=4.685 $Y=0.485 $X2=0
+ $Y2=0
cc_523 N_A_784_55#_c_728_n A_886_55# 0.00603173f $X=4.685 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_524 N_A_1662_57#_c_829_n N_VPWR_c_875_n 0.0685263f $X=8.45 $Y=1.98 $X2=0
+ $Y2=0
cc_525 N_A_1662_57#_c_829_n N_VPWR_c_876_n 0.00963752f $X=8.45 $Y=1.98 $X2=0
+ $Y2=0
cc_526 N_A_1662_57#_M1028_g N_VPWR_c_877_n 0.0250181f $X=9.275 $Y=2.545 $X2=0
+ $Y2=0
cc_527 N_A_1662_57#_c_829_n N_VPWR_c_877_n 0.0559573f $X=8.45 $Y=1.98 $X2=0
+ $Y2=0
cc_528 N_A_1662_57#_c_824_n N_VPWR_c_877_n 0.0207477f $X=8.865 $Y=1.675 $X2=0
+ $Y2=0
cc_529 N_A_1662_57#_c_827_n N_VPWR_c_877_n 0.00211868f $X=9.275 $Y=1.425 $X2=0
+ $Y2=0
cc_530 N_A_1662_57#_M1028_g N_VPWR_c_883_n 0.00767656f $X=9.275 $Y=2.545 $X2=0
+ $Y2=0
cc_531 N_A_1662_57#_M1028_g N_VPWR_c_871_n 0.014159f $X=9.275 $Y=2.545 $X2=0
+ $Y2=0
cc_532 N_A_1662_57#_c_829_n N_VPWR_c_871_n 0.0111417f $X=8.45 $Y=1.98 $X2=0
+ $Y2=0
cc_533 N_A_1662_57#_M1015_g Q_N 0.00219999f $X=9.225 $Y=0.67 $X2=0 $Y2=0
cc_534 N_A_1662_57#_M1017_g Q_N 0.0161322f $X=9.585 $Y=0.67 $X2=0 $Y2=0
cc_535 N_A_1662_57#_c_824_n Q_N 0.00696862f $X=8.865 $Y=1.675 $X2=0 $Y2=0
cc_536 N_A_1662_57#_c_825_n Q_N 0.018805f $X=9.03 $Y=1.255 $X2=0 $Y2=0
cc_537 N_A_1662_57#_c_827_n Q_N 0.0308658f $X=9.275 $Y=1.425 $X2=0 $Y2=0
cc_538 N_A_1662_57#_M1028_g Q_N 0.0209205f $X=9.275 $Y=2.545 $X2=0 $Y2=0
cc_539 N_A_1662_57#_c_823_n N_VGND_c_1021_n 0.0153904f $X=8.45 $Y=0.495 $X2=0
+ $Y2=0
cc_540 N_A_1662_57#_M1015_g N_VGND_c_1022_n 0.0137632f $X=9.225 $Y=0.67 $X2=0
+ $Y2=0
cc_541 N_A_1662_57#_M1017_g N_VGND_c_1022_n 0.00180376f $X=9.585 $Y=0.67 $X2=0
+ $Y2=0
cc_542 N_A_1662_57#_c_823_n N_VGND_c_1022_n 0.0428108f $X=8.45 $Y=0.495 $X2=0
+ $Y2=0
cc_543 N_A_1662_57#_c_825_n N_VGND_c_1022_n 0.0251002f $X=9.03 $Y=1.255 $X2=0
+ $Y2=0
cc_544 N_A_1662_57#_c_827_n N_VGND_c_1022_n 0.00219312f $X=9.275 $Y=1.425 $X2=0
+ $Y2=0
cc_545 N_A_1662_57#_c_823_n N_VGND_c_1027_n 0.0220321f $X=8.45 $Y=0.495 $X2=0
+ $Y2=0
cc_546 N_A_1662_57#_M1015_g N_VGND_c_1028_n 0.00426961f $X=9.225 $Y=0.67 $X2=0
+ $Y2=0
cc_547 N_A_1662_57#_M1017_g N_VGND_c_1028_n 0.00491683f $X=9.585 $Y=0.67 $X2=0
+ $Y2=0
cc_548 N_A_1662_57#_M1015_g N_VGND_c_1029_n 0.00434697f $X=9.225 $Y=0.67 $X2=0
+ $Y2=0
cc_549 N_A_1662_57#_M1017_g N_VGND_c_1029_n 0.00517496f $X=9.585 $Y=0.67 $X2=0
+ $Y2=0
cc_550 N_A_1662_57#_c_823_n N_VGND_c_1029_n 0.0125808f $X=8.45 $Y=0.495 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_875_n Q 0.0726161f $X=7.92 $Y=1.98 $X2=0 $Y2=0
cc_552 N_VPWR_c_882_n Q 0.0147493f $X=7.755 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_871_n Q 0.0157711f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_554 N_VPWR_c_877_n Q_N 0.0714805f $X=9.01 $Y=2.19 $X2=0 $Y2=0
cc_555 N_VPWR_c_883_n Q_N 0.0306496f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_556 N_VPWR_c_871_n Q_N 0.0217118f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_557 N_Q_c_963_n N_VGND_c_1021_n 0.0216684f $X=7.1 $Y=0.43 $X2=0 $Y2=0
cc_558 Q N_VGND_c_1021_n 0.00251427f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_559 N_Q_c_966_n N_VGND_c_1021_n 0.00773457f $X=7.327 $Y=1.18 $X2=0 $Y2=0
cc_560 N_Q_c_963_n N_VGND_c_1023_n 0.0360378f $X=7.1 $Y=0.43 $X2=0 $Y2=0
cc_561 N_Q_c_963_n N_VGND_c_1029_n 0.0208746f $X=7.1 $Y=0.43 $X2=0 $Y2=0
cc_562 N_Q_c_963_n A_1432_57# 0.00292994f $X=7.1 $Y=0.43 $X2=-0.19 $Y2=-0.245
cc_563 N_Q_c_966_n A_1432_57# 9.97329e-19 $X=7.327 $Y=1.18 $X2=-0.19 $Y2=-0.245
cc_564 Q_N N_VGND_c_1022_n 0.0153904f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_565 Q_N N_VGND_c_1028_n 0.0106618f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_566 Q_N N_VGND_c_1029_n 0.0114128f $X=9.755 $Y=0.47 $X2=0 $Y2=0
