* File: sky130_fd_sc_lp__dfxtp_lp.spice
* Created: Wed Sep  2 09:45:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfxtp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dfxtp_lp  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1026 A_112_57# N_CLK_M1026_g N_A_27_57#_M1026_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_CLK_M1020_g A_112_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1028 A_270_57# N_A_27_57#_M1028_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_263_409#_M1000_d N_A_27_57#_M1000_g A_270_57# VNB NSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.0441 PD=1.39 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 A_543_125# N_D_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1176 PD=0.7 PS=1.4 NRD=24.276 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.4
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_629_125#_M1004_d N_D_M1004_g A_543_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.12575 AS=0.0588 PD=1.09 PS=0.7 NRD=24.276 NRS=24.276 M=1 R=2.8 SA=75000.6
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1013 N_A_747_79#_M1013_d N_A_27_57#_M1013_g N_A_629_125#_M1004_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.13125 AS=0.12575 PD=1.275 PS=1.09 NRD=0 NRS=22.848 M=1
+ R=2.8 SA=75000.7 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1024 A_902_125# N_A_263_409#_M1024_g N_A_747_79#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.10815 AS=0.13125 PD=0.935 PS=1.275 NRD=57.852 NRS=99.996 M=1 R=2.8
+ SA=75001 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1005_99#_M1029_g A_902_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.34075 AS=0.10815 PD=2.12 PS=0.935 NRD=216.084 NRS=57.852 M=1 R=2.8
+ SA=75001.7 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1021 A_1355_125# N_A_747_79#_M1021_g N_VGND_M1029_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.34075 PD=0.63 PS=2.12 NRD=14.28 NRS=216.084 M=1 R=2.8
+ SA=75003.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1018 N_A_1005_99#_M1018_d N_A_747_79#_M1018_g A_1355_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.0609 AS=0.0441 PD=0.71 PS=0.63 NRD=1.428 NRS=14.28 M=1 R=2.8
+ SA=75003.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1006 N_A_1429_383#_M1006_d N_A_263_409#_M1006_g N_A_1005_99#_M1018_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.1013 AS=0.0609 PD=1.075 PS=0.71 NRD=53.196 NRS=1.428
+ M=1 R=2.8 SA=75004.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 A_1626_75# N_A_27_57#_M1001_g N_A_1429_383#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1013 PD=0.63 PS=1.075 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_1583_285#_M1002_g A_1626_75# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1012 A_1784_75# N_A_1429_383#_M1012_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_1583_285#_M1014_d N_A_1429_383#_M1014_g A_1784_75# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_2054_92# N_A_1583_285#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_Q_M1025_d N_A_1583_285#_M1025_g A_2054_92# VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0441 PD=1.39 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_CLK_M1003_g N_A_27_57#_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1019 N_A_263_409#_M1019_d N_A_27_57#_M1019_g N_VPWR_M1003_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1022 N_A_629_125#_M1022_d N_D_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.25 W=1
+ AD=0.348225 AS=0.365 PD=1.7 PS=2.73 NRD=26.5753 NRS=15.7403 M=1 R=4 SA=125000
+ SB=125005 A=0.25 P=2.5 MULT=1
MM1010 N_A_747_79#_M1010_d N_A_263_409#_M1010_g N_A_629_125#_M1022_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.24175 AS=0.348225 PD=1.59 PS=1.7 NRD=16.0752 NRS=55.1403 M=1
+ R=4 SA=125001 SB=125004 A=0.25 P=2.5 MULT=1
MM1007 A_962_371# N_A_27_57#_M1007_g N_A_747_79#_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.175625 AS=0.24175 PD=1.475 PS=1.59 NRD=23.7582 NRS=16.0752 M=1 R=4
+ SA=125002 SB=125004 A=0.25 P=2.5 MULT=1
MM1016 N_VPWR_M1016_d N_A_1005_99#_M1016_g A_962_371# VPB PHIGHVT L=0.25 W=1
+ AD=0.41 AS=0.175625 PD=1.82 PS=1.475 NRD=0 NRS=23.7582 M=1 R=4 SA=125002
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1015 N_A_1005_99#_M1015_d N_A_747_79#_M1015_g N_VPWR_M1016_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.25045 AS=0.41 PD=1.65 PS=1.82 NRD=16.0752 NRS=106.36 M=1 R=4
+ SA=125003 SB=125003 A=0.25 P=2.5 MULT=1
MM1008 N_A_1429_383#_M1008_d N_A_27_57#_M1008_g N_A_1005_99#_M1015_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.25045 PD=1.28 PS=1.65 NRD=0 NRS=16.0752 M=1 R=4
+ SA=125003 SB=125002 A=0.25 P=2.5 MULT=1
MM1023 A_1535_383# N_A_263_409#_M1023_g N_A_1429_383#_M1008_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125004
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_A_1583_285#_M1005_g A_1535_383# VPB PHIGHVT L=0.25 W=1
+ AD=0.46 AS=0.12 PD=1.92 PS=1.24 NRD=77.7953 NRS=12.7853 M=1 R=4 SA=125004
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1017 N_A_1583_285#_M1017_d N_A_1429_383#_M1017_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.365 AS=0.46 PD=2.73 PS=1.92 NRD=15.7403 NRS=48.2453 M=1 R=4
+ SA=125006 SB=125000 A=0.25 P=2.5 MULT=1
MM1027 N_Q_M1027_d N_A_1583_285#_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX30_noxref VNB VPB NWDIODE A=21.8989 P=26.83
c_114 VNB 0 1.17622e-19 $X=0 $Y=0
c_192 VPB 0 7.95967e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dfxtp_lp.pxi.spice"
*
.ends
*
*
