* File: sky130_fd_sc_lp__sdfrbp_2.pxi.spice
* Created: Fri Aug 28 11:27:50 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRBP_2%SCE N_SCE_M1014_g N_SCE_c_287_n N_SCE_c_288_n
+ N_SCE_M1021_g N_SCE_c_289_n N_SCE_c_290_n N_SCE_M1004_g N_SCE_M1024_g
+ N_SCE_c_291_n N_SCE_c_292_n N_SCE_c_282_n N_SCE_c_283_n N_SCE_c_284_n SCE SCE
+ N_SCE_c_285_n N_SCE_c_300_p SCE N_SCE_c_286_n PM_SKY130_FD_SC_LP__SDFRBP_2%SCE
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_27_81# N_A_27_81#_M1014_s N_A_27_81#_M1021_s
+ N_A_27_81#_c_368_n N_A_27_81#_c_369_n N_A_27_81#_c_370_n N_A_27_81#_c_371_n
+ N_A_27_81#_M1033_g N_A_27_81#_M1041_g N_A_27_81#_c_372_n N_A_27_81#_c_373_n
+ N_A_27_81#_c_374_n N_A_27_81#_c_375_n N_A_27_81#_c_379_n N_A_27_81#_c_380_n
+ N_A_27_81#_c_381_n N_A_27_81#_c_382_n N_A_27_81#_c_376_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_27_81#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%D N_D_M1009_g N_D_M1035_g D D N_D_c_457_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%D
x_PM_SKY130_FD_SC_LP__SDFRBP_2%SCD N_SCD_M1034_g N_SCD_M1047_g N_SCD_c_501_n
+ N_SCD_c_502_n SCD SCD N_SCD_c_499_n PM_SKY130_FD_SC_LP__SDFRBP_2%SCD
x_PM_SKY130_FD_SC_LP__SDFRBP_2%CLK N_CLK_c_541_n N_CLK_M1019_g N_CLK_c_542_n
+ N_CLK_M1022_g N_CLK_M1042_g CLK CLK N_CLK_c_545_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%CLK
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_934_367# N_A_934_367#_M1013_d
+ N_A_934_367#_M1017_d N_A_934_367#_M1038_g N_A_934_367#_c_594_n
+ N_A_934_367#_M1028_g N_A_934_367#_M1046_g N_A_934_367#_M1032_g
+ N_A_934_367#_c_596_n N_A_934_367#_c_597_n N_A_934_367#_c_598_n
+ N_A_934_367#_c_599_n N_A_934_367#_c_600_n N_A_934_367#_c_615_p
+ N_A_934_367#_c_620_p N_A_934_367#_c_601_n N_A_934_367#_c_602_n
+ N_A_934_367#_c_608_n N_A_934_367#_c_609_n N_A_934_367#_c_603_n
+ N_A_934_367#_c_611_n N_A_934_367#_c_612_n N_A_934_367#_c_604_n
+ N_A_934_367#_c_605_n PM_SKY130_FD_SC_LP__SDFRBP_2%A_934_367#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_1290_365# N_A_1290_365#_M1005_d
+ N_A_1290_365#_M1031_d N_A_1290_365#_M1000_g N_A_1290_365#_M1036_g
+ N_A_1290_365#_c_782_n N_A_1290_365#_c_789_n N_A_1290_365#_c_783_n
+ N_A_1290_365#_c_784_n N_A_1290_365#_c_807_n N_A_1290_365#_c_819_p
+ N_A_1290_365#_c_790_n N_A_1290_365#_c_785_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_1290_365#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%RESET_B N_RESET_B_M1002_g N_RESET_B_M1015_g
+ N_RESET_B_c_859_n N_RESET_B_c_860_n N_RESET_B_c_865_n N_RESET_B_M1018_g
+ N_RESET_B_M1025_g N_RESET_B_M1016_g N_RESET_B_M1012_g N_RESET_B_c_869_n
+ N_RESET_B_c_870_n N_RESET_B_c_871_n N_RESET_B_c_872_n N_RESET_B_c_873_n
+ RESET_B N_RESET_B_c_875_n N_RESET_B_c_876_n N_RESET_B_c_877_n
+ N_RESET_B_c_878_n N_RESET_B_c_879_n PM_SKY130_FD_SC_LP__SDFRBP_2%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_1162_463# N_A_1162_463#_M1043_d
+ N_A_1162_463#_M1038_d N_A_1162_463#_M1018_d N_A_1162_463#_M1005_g
+ N_A_1162_463#_M1031_g N_A_1162_463#_c_1069_n N_A_1162_463#_c_1064_n
+ N_A_1162_463#_c_1095_n N_A_1162_463#_c_1071_n N_A_1162_463#_c_1065_n
+ N_A_1162_463#_c_1083_n N_A_1162_463#_c_1106_n N_A_1162_463#_c_1107_n
+ N_A_1162_463#_c_1066_n N_A_1162_463#_c_1067_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_1162_463#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_759_119# N_A_759_119#_M1019_d
+ N_A_759_119#_M1042_s N_A_759_119#_M1017_g N_A_759_119#_c_1177_n
+ N_A_759_119#_M1013_g N_A_759_119#_c_1178_n N_A_759_119#_c_1179_n
+ N_A_759_119#_M1027_g N_A_759_119#_c_1193_n N_A_759_119#_c_1194_n
+ N_A_759_119#_c_1180_n N_A_759_119#_c_1181_n N_A_759_119#_M1023_g
+ N_A_759_119#_c_1182_n N_A_759_119#_M1043_g N_A_759_119#_c_1196_n
+ N_A_759_119#_M1010_g N_A_759_119#_c_1183_n N_A_759_119#_c_1184_n
+ N_A_759_119#_M1040_g N_A_759_119#_c_1200_n N_A_759_119#_c_1186_n
+ N_A_759_119#_c_1209_n N_A_759_119#_c_1187_n N_A_759_119#_c_1188_n
+ N_A_759_119#_c_1189_n N_A_759_119#_c_1219_n N_A_759_119#_c_1190_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_759_119#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_1923_174# N_A_1923_174#_M1020_d
+ N_A_1923_174#_M1012_d N_A_1923_174#_M1044_g N_A_1923_174#_M1001_g
+ N_A_1923_174#_c_1361_n N_A_1923_174#_c_1362_n N_A_1923_174#_c_1363_n
+ N_A_1923_174#_c_1364_n N_A_1923_174#_c_1365_n N_A_1923_174#_c_1366_n
+ N_A_1923_174#_c_1371_n N_A_1923_174#_c_1372_n N_A_1923_174#_c_1367_n
+ N_A_1923_174#_c_1373_n N_A_1923_174#_c_1368_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_1923_174#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_1770_412# N_A_1770_412#_M1046_d
+ N_A_1770_412#_M1010_d N_A_1770_412#_M1020_g N_A_1770_412#_M1045_g
+ N_A_1770_412#_c_1456_n N_A_1770_412#_M1007_g N_A_1770_412#_M1003_g
+ N_A_1770_412#_c_1459_n N_A_1770_412#_M1039_g N_A_1770_412#_M1037_g
+ N_A_1770_412#_c_1462_n N_A_1770_412#_M1029_g N_A_1770_412#_M1011_g
+ N_A_1770_412#_c_1465_n N_A_1770_412#_c_1466_n N_A_1770_412#_c_1467_n
+ N_A_1770_412#_c_1485_n N_A_1770_412#_c_1490_n N_A_1770_412#_c_1468_n
+ N_A_1770_412#_c_1469_n N_A_1770_412#_c_1470_n N_A_1770_412#_c_1479_n
+ N_A_1770_412#_c_1471_n N_A_1770_412#_c_1481_n N_A_1770_412#_c_1472_n
+ N_A_1770_412#_c_1473_n N_A_1770_412#_c_1474_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_1770_412#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_2516_367# N_A_2516_367#_M1011_d
+ N_A_2516_367#_M1029_d N_A_2516_367#_c_1643_n N_A_2516_367#_M1006_g
+ N_A_2516_367#_M1008_g N_A_2516_367#_c_1645_n N_A_2516_367#_M1030_g
+ N_A_2516_367#_M1026_g N_A_2516_367#_c_1647_n N_A_2516_367#_c_1648_n
+ N_A_2516_367#_c_1649_n N_A_2516_367#_c_1650_n N_A_2516_367#_c_1651_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_2516_367#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%VPWR N_VPWR_M1021_d N_VPWR_M1034_d N_VPWR_M1042_d
+ N_VPWR_M1000_d N_VPWR_M1031_s N_VPWR_M1001_d N_VPWR_M1045_d N_VPWR_M1039_s
+ N_VPWR_M1008_d N_VPWR_M1026_d N_VPWR_c_1702_n N_VPWR_c_1703_n N_VPWR_c_1704_n
+ N_VPWR_c_1705_n N_VPWR_c_1706_n N_VPWR_c_1707_n N_VPWR_c_1708_n
+ N_VPWR_c_1709_n N_VPWR_c_1710_n N_VPWR_c_1711_n N_VPWR_c_1712_n
+ N_VPWR_c_1713_n N_VPWR_c_1714_n N_VPWR_c_1715_n N_VPWR_c_1716_n
+ N_VPWR_c_1717_n VPWR N_VPWR_c_1718_n N_VPWR_c_1719_n N_VPWR_c_1720_n
+ N_VPWR_c_1721_n N_VPWR_c_1722_n N_VPWR_c_1723_n N_VPWR_c_1724_n
+ N_VPWR_c_1725_n N_VPWR_c_1726_n N_VPWR_c_1727_n N_VPWR_c_1728_n
+ N_VPWR_c_1729_n N_VPWR_c_1730_n N_VPWR_c_1701_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%VPWR
x_PM_SKY130_FD_SC_LP__SDFRBP_2%A_359_489# N_A_359_489#_M1035_d
+ N_A_359_489#_M1043_s N_A_359_489#_M1009_d N_A_359_489#_M1002_d
+ N_A_359_489#_M1038_s N_A_359_489#_c_1916_n N_A_359_489#_c_1902_n
+ N_A_359_489#_c_1903_n N_A_359_489#_c_1907_n N_A_359_489#_c_1908_n
+ N_A_359_489#_c_1909_n N_A_359_489#_c_1910_n N_A_359_489#_c_1904_n
+ N_A_359_489#_c_1912_n N_A_359_489#_c_1905_n N_A_359_489#_c_1913_n
+ N_A_359_489#_c_1914_n N_A_359_489#_c_1915_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%A_359_489#
x_PM_SKY130_FD_SC_LP__SDFRBP_2%Q_N N_Q_N_M1003_s N_Q_N_M1007_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_2043_n PM_SKY130_FD_SC_LP__SDFRBP_2%Q_N
x_PM_SKY130_FD_SC_LP__SDFRBP_2%Q N_Q_M1006_s N_Q_M1008_s Q Q Q Q Q Q Q
+ N_Q_c_2065_n PM_SKY130_FD_SC_LP__SDFRBP_2%Q
x_PM_SKY130_FD_SC_LP__SDFRBP_2%VGND N_VGND_M1014_d N_VGND_M1015_d N_VGND_M1022_s
+ N_VGND_M1027_s N_VGND_M1025_d N_VGND_M1044_d N_VGND_M1003_d N_VGND_M1037_d
+ N_VGND_M1006_d N_VGND_M1030_d N_VGND_c_2083_n N_VGND_c_2084_n N_VGND_c_2085_n
+ N_VGND_c_2086_n N_VGND_c_2087_n N_VGND_c_2088_n N_VGND_c_2089_n
+ N_VGND_c_2090_n N_VGND_c_2091_n N_VGND_c_2092_n N_VGND_c_2093_n
+ N_VGND_c_2094_n N_VGND_c_2095_n N_VGND_c_2096_n N_VGND_c_2097_n
+ N_VGND_c_2098_n N_VGND_c_2099_n N_VGND_c_2100_n N_VGND_c_2101_n VGND
+ N_VGND_c_2102_n N_VGND_c_2103_n N_VGND_c_2104_n N_VGND_c_2105_n
+ N_VGND_c_2106_n N_VGND_c_2107_n N_VGND_c_2108_n N_VGND_c_2109_n
+ N_VGND_c_2110_n N_VGND_c_2111_n N_VGND_c_2112_n N_VGND_c_2113_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%VGND
x_PM_SKY130_FD_SC_LP__SDFRBP_2%noxref_25 N_noxref_25_M1033_s N_noxref_25_M1047_d
+ N_noxref_25_c_2245_n N_noxref_25_c_2246_n N_noxref_25_c_2247_n
+ PM_SKY130_FD_SC_LP__SDFRBP_2%noxref_25
cc_1 VNB N_SCE_M1014_g 0.0614052f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.615
cc_2 VNB N_SCE_M1024_g 0.0216341f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.615
cc_3 VNB N_SCE_c_282_n 0.0056018f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.675
cc_4 VNB N_SCE_c_283_n 0.00576046f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_5 VNB N_SCE_c_284_n 0.0353486f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_6 VNB N_SCE_c_285_n 0.0370819f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.68
cc_7 VNB N_SCE_c_286_n 0.0032464f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.68
cc_8 VNB N_A_27_81#_c_368_n 0.0401425f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_9 VNB N_A_27_81#_c_369_n 0.0337086f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_10 VNB N_A_27_81#_c_370_n 0.0163205f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.26
cc_11 VNB N_A_27_81#_c_371_n 0.0157627f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.26
cc_12 VNB N_A_27_81#_c_372_n 0.0194304f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.76
cc_13 VNB N_A_27_81#_c_373_n 0.0201834f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.675
cc_14 VNB N_A_27_81#_c_374_n 0.0120624f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_15 VNB N_A_27_81#_c_375_n 0.0340454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_81#_c_376_n 0.015373f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.68
cc_17 VNB N_D_M1009_g 0.0105071f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.615
cc_18 VNB N_D_M1035_g 0.0289571f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.335
cc_19 VNB D 0.0074374f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_20 VNB N_D_c_457_n 0.0489201f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.615
cc_21 VNB N_SCD_M1047_g 0.0508699f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.335
cc_22 VNB SCD 0.00409677f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.765
cc_23 VNB N_SCD_c_499_n 0.00928164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_CLK_c_541_n 0.0136245f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.515
cc_25 VNB N_CLK_c_542_n 0.0137057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_CLK_M1042_g 0.00279f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_27 VNB CLK 0.0114824f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.765
cc_28 VNB N_CLK_c_545_n 0.0679159f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_29 VNB N_A_934_367#_c_594_n 0.0572274f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.26
cc_30 VNB N_A_934_367#_M1028_g 0.0258274f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.065
cc_31 VNB N_A_934_367#_c_596_n 0.0118624f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_32 VNB N_A_934_367#_c_597_n 0.00139456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_934_367#_c_598_n 0.0227826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_934_367#_c_599_n 0.00343443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_934_367#_c_600_n 0.00108121f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.68
cc_36 VNB N_A_934_367#_c_601_n 0.0072612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_934_367#_c_602_n 0.0322432f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_38 VNB N_A_934_367#_c_603_n 0.0132673f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.68
cc_39 VNB N_A_934_367#_c_604_n 0.0177366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_934_367#_c_605_n 0.0190529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1290_365#_M1036_g 0.0355942f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.765
cc_42 VNB N_A_1290_365#_c_782_n 0.00386583f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.615
cc_43 VNB N_A_1290_365#_c_783_n 0.0216367f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.76
cc_44 VNB N_A_1290_365#_c_784_n 7.24291e-19 $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=1.76
cc_45 VNB N_A_1290_365#_c_785_n 0.00832646f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.58
cc_46 VNB N_RESET_B_M1015_g 0.0524509f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_47 VNB N_RESET_B_c_859_n 0.299094f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_48 VNB N_RESET_B_c_860_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.26
cc_49 VNB N_RESET_B_M1025_g 0.055326f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.615
cc_50 VNB N_RESET_B_M1016_g 0.0471651f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.76
cc_51 VNB N_A_1162_463#_M1005_g 0.0418821f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.335
cc_52 VNB N_A_1162_463#_c_1064_n 0.00534568f $X=-0.19 $Y=-0.245 $X2=2.27
+ $Y2=1.675
cc_53 VNB N_A_1162_463#_c_1065_n 2.34762e-19 $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_54 VNB N_A_1162_463#_c_1066_n 0.02681f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_55 VNB N_A_1162_463#_c_1067_n 0.0107292f $X=-0.19 $Y=-0.245 $X2=2.35
+ $Y2=1.065
cc_56 VNB N_A_759_119#_M1017_g 0.00239128f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_57 VNB N_A_759_119#_c_1177_n 0.0136455f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.26
cc_58 VNB N_A_759_119#_c_1178_n 0.00183601f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=1.065
cc_59 VNB N_A_759_119#_c_1179_n 0.0137372f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.615
cc_60 VNB N_A_759_119#_c_1180_n 0.0588172f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.76
cc_61 VNB N_A_759_119#_c_1181_n 0.06056f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.395
cc_62 VNB N_A_759_119#_c_1182_n 0.0131348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_759_119#_c_1183_n 0.0129655f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.68
cc_64 VNB N_A_759_119#_c_1184_n 0.00283737f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.68
cc_65 VNB N_A_759_119#_M1040_g 0.0529212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_759_119#_c_1186_n 0.00418456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_759_119#_c_1187_n 0.00453346f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.68
cc_68 VNB N_A_759_119#_c_1188_n 0.00110293f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_69 VNB N_A_759_119#_c_1189_n 0.0037708f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.68
cc_70 VNB N_A_759_119#_c_1190_n 0.00303063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1923_174#_M1001_g 0.0226161f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.335
cc_72 VNB N_A_1923_174#_c_1361_n 0.0300565f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.615
cc_73 VNB N_A_1923_174#_c_1362_n 0.00604801f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=2.26
cc_74 VNB N_A_1923_174#_c_1363_n 0.00189158f $X=-0.19 $Y=-0.245 $X2=2.185
+ $Y2=1.76
cc_75 VNB N_A_1923_174#_c_1364_n 0.00758711f $X=-0.19 $Y=-0.245 $X2=2.27
+ $Y2=1.675
cc_76 VNB N_A_1923_174#_c_1365_n 0.00419186f $X=-0.19 $Y=-0.245 $X2=2.35
+ $Y2=1.395
cc_77 VNB N_A_1923_174#_c_1366_n 0.00841306f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_78 VNB N_A_1923_174#_c_1367_n 0.0178508f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=1.68
cc_79 VNB N_A_1923_174#_c_1368_n 0.0175041f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_80 VNB N_A_1770_412#_M1020_g 0.0477722f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.765
cc_81 VNB N_A_1770_412#_c_1456_n 0.0286556f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=1.065
cc_82 VNB N_A_1770_412#_M1007_g 0.00699844f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.26
cc_83 VNB N_A_1770_412#_M1003_g 0.0302611f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.675
cc_84 VNB N_A_1770_412#_c_1459_n 0.00983103f $X=-0.19 $Y=-0.245 $X2=2.35
+ $Y2=1.23
cc_85 VNB N_A_1770_412#_M1039_g 0.00623595f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_86 VNB N_A_1770_412#_M1037_g 0.0273082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1770_412#_c_1462_n 0.0151002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1770_412#_M1029_g 0.00791199f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.68
cc_89 VNB N_A_1770_412#_M1011_g 0.0596174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1770_412#_c_1465_n 0.00270629f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.68
cc_91 VNB N_A_1770_412#_c_1466_n 0.00270629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1770_412#_c_1467_n 0.00647697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1770_412#_c_1468_n 0.00897395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1770_412#_c_1469_n 0.0106006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1770_412#_c_1470_n 0.0017616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1770_412#_c_1471_n 0.00419533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1770_412#_c_1472_n 0.00376919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1770_412#_c_1473_n 0.00198975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1770_412#_c_1474_n 0.0257421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2516_367#_c_1643_n 0.0192445f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=2.335
cc_101 VNB N_A_2516_367#_M1008_g 0.00578998f $X=-0.19 $Y=-0.245 $X2=1.36
+ $Y2=2.335
cc_102 VNB N_A_2516_367#_c_1645_n 0.0211749f $X=-0.19 $Y=-0.245 $X2=1.36
+ $Y2=2.765
cc_103 VNB N_A_2516_367#_M1026_g 0.00753401f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=2.26
cc_104 VNB N_A_2516_367#_c_1647_n 0.0113211f $X=-0.19 $Y=-0.245 $X2=2.27
+ $Y2=1.675
cc_105 VNB N_A_2516_367#_c_1648_n 0.00167746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2516_367#_c_1649_n 0.0161825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2516_367#_c_1650_n 0.00234025f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=1.68
cc_108 VNB N_A_2516_367#_c_1651_n 0.0720285f $X=-0.19 $Y=-0.245 $X2=1.14
+ $Y2=1.68
cc_109 VNB N_VPWR_c_1701_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_359_489#_c_1902_n 0.00861231f $X=-0.19 $Y=-0.245 $X2=2.185
+ $Y2=1.76
cc_111 VNB N_A_359_489#_c_1903_n 0.0143072f $X=-0.19 $Y=-0.245 $X2=2.27
+ $Y2=1.675
cc_112 VNB N_A_359_489#_c_1904_n 0.00533699f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=1.68
cc_113 VNB N_A_359_489#_c_1905_n 0.00990342f $X=-0.19 $Y=-0.245 $X2=1.14
+ $Y2=1.68
cc_114 VNB N_Q_N_c_2043_n 0.00731622f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.395
cc_115 VNB N_Q_c_2065_n 0.00596029f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.395
cc_116 VNB N_VGND_c_2083_n 0.0111582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2084_n 0.00615701f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.68
cc_118 VNB N_VGND_c_2085_n 0.00937698f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.23
cc_119 VNB N_VGND_c_2086_n 0.0101738f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.68
cc_120 VNB N_VGND_c_2087_n 0.00889511f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.68
cc_121 VNB N_VGND_c_2088_n 0.00319234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2089_n 0.0116807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2090_n 0.0161796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2091_n 0.0113072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2092_n 0.0117359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2093_n 0.0456412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2094_n 0.059261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2095_n 0.0034624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2096_n 0.0172836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2097_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2098_n 0.0175989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2099_n 0.00226387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2100_n 0.0541677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2101_n 0.00567616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2102_n 0.017242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2103_n 0.0517562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2104_n 0.0281017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2105_n 0.0167145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2106_n 0.0189835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2107_n 0.0152915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2108_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2109_n 0.00631927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2110_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2111_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2112_n 0.00517589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2113_n 0.714336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_noxref_25_c_2245_n 0.00896647f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=2.335
cc_148 VNB N_noxref_25_c_2246_n 4.58069e-19 $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=2.765
cc_149 VNB N_noxref_25_c_2247_n 0.00225349f $X=-0.19 $Y=-0.245 $X2=1.36
+ $Y2=2.335
cc_150 VPB N_SCE_c_287_n 0.0196369f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.185
cc_151 VPB N_SCE_c_288_n 0.0200361f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.335
cc_152 VPB N_SCE_c_289_n 0.01934f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.26
cc_153 VPB N_SCE_c_290_n 0.0153707f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.335
cc_154 VPB N_SCE_c_291_n 0.00664226f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.26
cc_155 VPB N_SCE_c_292_n 0.0265861f $X=-0.19 $Y=1.655 $X2=2.185 $Y2=1.76
cc_156 VPB N_SCE_c_282_n 4.53481e-19 $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.675
cc_157 VPB N_SCE_c_285_n 0.0430577f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.68
cc_158 VPB N_SCE_c_286_n 4.92123e-19 $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.68
cc_159 VPB N_A_27_81#_M1041_g 0.0203335f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.615
cc_160 VPB N_A_27_81#_c_373_n 0.0198654f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.675
cc_161 VPB N_A_27_81#_c_379_n 0.033126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_27_81#_c_380_n 0.0354348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_27_81#_c_381_n 0.0176942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_27_81#_c_382_n 0.0322204f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.68
cc_165 VPB N_D_M1009_g 0.058038f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.615
cc_166 VPB N_SCD_M1034_g 0.0211976f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.615
cc_167 VPB N_SCD_c_501_n 0.0243259f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.26
cc_168 VPB N_SCD_c_502_n 0.0151558f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.335
cc_169 VPB SCD 0.00902817f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.765
cc_170 VPB N_SCD_c_499_n 0.00953234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_CLK_M1042_g 0.0261201f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.765
cc_172 VPB CLK 0.0071909f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.765
cc_173 VPB N_A_934_367#_M1038_g 0.0445245f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.765
cc_174 VPB N_A_934_367#_M1032_g 0.0221168f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.395
cc_175 VPB N_A_934_367#_c_608_n 0.00211647f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.065
cc_176 VPB N_A_934_367#_c_609_n 0.00163866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_934_367#_c_603_n 0.0103179f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.68
cc_178 VPB N_A_934_367#_c_611_n 0.00926272f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.665
cc_179 VPB N_A_934_367#_c_612_n 0.0347726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_934_367#_c_604_n 0.0184455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_1290_365#_M1000_g 0.0195674f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.765
cc_182 VPB N_A_1290_365#_M1036_g 0.00116044f $X=-0.19 $Y=1.655 $X2=1.36
+ $Y2=2.765
cc_183 VPB N_A_1290_365#_c_782_n 0.00416947f $X=-0.19 $Y=1.655 $X2=2.355
+ $Y2=0.615
cc_184 VPB N_A_1290_365#_c_789_n 0.065528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1290_365#_c_790_n 0.0038176f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.23
cc_186 VPB N_A_1290_365#_c_785_n 0.00749235f $X=-0.19 $Y=1.655 $X2=1.115
+ $Y2=1.58
cc_187 VPB N_RESET_B_M1002_g 0.0310574f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.615
cc_188 VPB N_RESET_B_M1015_g 0.010957f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.765
cc_189 VPB N_RESET_B_c_865_n 0.0164531f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.26
cc_190 VPB N_RESET_B_M1025_g 0.00973488f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.615
cc_191 VPB N_RESET_B_M1016_g 0.0165388f $X=-0.19 $Y=1.655 $X2=2.185 $Y2=1.76
cc_192 VPB N_RESET_B_M1012_g 0.020742f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.23
cc_193 VPB N_RESET_B_c_869_n 0.0112785f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.23
cc_194 VPB N_RESET_B_c_870_n 0.00176516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_RESET_B_c_871_n 0.0245018f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.395
cc_196 VPB N_RESET_B_c_872_n 3.70249e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_197 VPB N_RESET_B_c_873_n 0.00130189f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.68
cc_198 VPB RESET_B 0.00147278f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.68
cc_199 VPB N_RESET_B_c_875_n 0.0516172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_RESET_B_c_876_n 0.00175319f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=1.68
cc_201 VPB N_RESET_B_c_877_n 0.0595127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_RESET_B_c_878_n 0.0382392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_c_879_n 0.00408033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1162_463#_M1031_g 0.0211892f $X=-0.19 $Y=1.655 $X2=2.355
+ $Y2=0.615
cc_205 VPB N_A_1162_463#_c_1069_n 0.00200829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1162_463#_c_1064_n 0.010242f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.675
cc_207 VPB N_A_1162_463#_c_1071_n 0.00926724f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1162_463#_c_1066_n 0.0149645f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.23
cc_209 VPB N_A_759_119#_M1017_g 0.0205557f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.765
cc_210 VPB N_A_759_119#_c_1178_n 0.0807518f $X=-0.19 $Y=1.655 $X2=2.355
+ $Y2=1.065
cc_211 VPB N_A_759_119#_c_1193_n 0.0651644f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.26
cc_212 VPB N_A_759_119#_c_1194_n 0.00989679f $X=-0.19 $Y=1.655 $X2=2.185
+ $Y2=1.76
cc_213 VPB N_A_759_119#_M1023_g 0.0363577f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.23
cc_214 VPB N_A_759_119#_c_1196_n 0.195177f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_215 VPB N_A_759_119#_M1010_g 0.0311795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_759_119#_c_1183_n 0.0230453f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.68
cc_217 VPB N_A_759_119#_c_1184_n 0.00507009f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.68
cc_218 VPB N_A_759_119#_c_1200_n 0.00749069f $X=-0.19 $Y=1.655 $X2=2.35
+ $Y2=1.065
cc_219 VPB N_A_759_119#_c_1188_n 0.00289249f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.665
cc_220 VPB N_A_1923_174#_M1001_g 0.0522999f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.335
cc_221 VPB N_A_1923_174#_c_1365_n 0.00450235f $X=-0.19 $Y=1.655 $X2=2.35
+ $Y2=1.395
cc_222 VPB N_A_1923_174#_c_1371_n 9.01215e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_1923_174#_c_1372_n 0.00316093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1923_174#_c_1373_n 0.00915761f $X=-0.19 $Y=1.655 $X2=1.14
+ $Y2=1.68
cc_225 VPB N_A_1770_412#_M1045_g 0.0502421f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.765
cc_226 VPB N_A_1770_412#_M1007_g 0.0226f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.26
cc_227 VPB N_A_1770_412#_M1039_g 0.022327f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_228 VPB N_A_1770_412#_M1029_g 0.0256385f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.68
cc_229 VPB N_A_1770_412#_c_1479_n 0.00545656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_1770_412#_c_1471_n 0.00381811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_1770_412#_c_1481_n 0.00306534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_1770_412#_c_1473_n 0.00107197f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1770_412#_c_1474_n 0.0200884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_2516_367#_M1008_g 0.023501f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.335
cc_235 VPB N_A_2516_367#_M1026_g 0.0271626f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.26
cc_236 VPB N_A_2516_367#_c_1648_n 0.0155278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1702_n 0.00434601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1703_n 0.00314922f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.68
cc_239 VPB N_VPWR_c_1704_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.23
cc_240 VPB N_VPWR_c_1705_n 0.0085795f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.68
cc_241 VPB N_VPWR_c_1706_n 0.021936f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.68
cc_242 VPB N_VPWR_c_1707_n 0.00819156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1708_n 0.0342255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1709_n 0.0318423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1710_n 0.01171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1711_n 0.0592771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1712_n 0.0355903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1713_n 0.00517888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1714_n 0.0306899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1715_n 0.0043639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1716_n 0.0584272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1717_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1718_n 0.0321584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1719_n 0.020199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1720_n 0.0457563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1721_n 0.0204151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1722_n 0.0155485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1723_n 0.0218935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1724_n 0.0149952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1725_n 0.00383448f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1726_n 0.00330333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1727_n 0.0268252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1728_n 0.00522677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1729_n 0.0061259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1730_n 0.00484208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1701_n 0.109202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_359_489#_c_1903_n 0.00723661f $X=-0.19 $Y=1.655 $X2=2.27
+ $Y2=1.675
cc_268 VPB N_A_359_489#_c_1907_n 0.0154716f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.23
cc_269 VPB N_A_359_489#_c_1908_n 5.11207e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_359_489#_c_1909_n 0.00690391f $X=-0.19 $Y=1.655 $X2=1.115
+ $Y2=1.58
cc_271 VPB N_A_359_489#_c_1910_n 0.00290116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_359_489#_c_1904_n 0.00544118f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=1.68
cc_273 VPB N_A_359_489#_c_1912_n 0.00154424f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.68
cc_274 VPB N_A_359_489#_c_1913_n 0.00651043f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.68
cc_275 VPB N_A_359_489#_c_1914_n 0.00246313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_359_489#_c_1915_n 0.00391196f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.68
cc_277 VPB N_Q_N_c_2043_n 0.00176292f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.395
cc_278 VPB N_Q_c_2065_n 0.00401513f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.395
cc_279 N_SCE_M1014_g N_A_27_81#_c_370_n 0.0267688f $X=0.475 $Y=0.615 $X2=0 $Y2=0
cc_280 N_SCE_M1014_g N_A_27_81#_c_372_n 0.0044975f $X=0.475 $Y=0.615 $X2=0 $Y2=0
cc_281 N_SCE_M1014_g N_A_27_81#_c_373_n 0.0207812f $X=0.475 $Y=0.615 $X2=0 $Y2=0
cc_282 N_SCE_c_287_n N_A_27_81#_c_373_n 0.00483323f $X=0.93 $Y=2.185 $X2=0 $Y2=0
cc_283 N_SCE_c_300_p N_A_27_81#_c_373_n 0.0271102f $X=1.18 $Y=1.68 $X2=0 $Y2=0
cc_284 N_SCE_M1014_g N_A_27_81#_c_374_n 0.0282808f $X=0.475 $Y=0.615 $X2=0 $Y2=0
cc_285 N_SCE_c_285_n N_A_27_81#_c_374_n 0.00893016f $X=1.14 $Y=1.68 $X2=0 $Y2=0
cc_286 N_SCE_c_300_p N_A_27_81#_c_374_n 0.0411154f $X=1.18 $Y=1.68 $X2=0 $Y2=0
cc_287 N_SCE_c_285_n N_A_27_81#_c_375_n 0.0190503f $X=1.14 $Y=1.68 $X2=0 $Y2=0
cc_288 N_SCE_c_300_p N_A_27_81#_c_375_n 0.00150571f $X=1.18 $Y=1.68 $X2=0 $Y2=0
cc_289 N_SCE_c_288_n N_A_27_81#_c_379_n 0.0107013f $X=0.93 $Y=2.335 $X2=0 $Y2=0
cc_290 N_SCE_c_290_n N_A_27_81#_c_379_n 6.67685e-19 $X=1.36 $Y=2.335 $X2=0 $Y2=0
cc_291 N_SCE_c_291_n N_A_27_81#_c_379_n 0.00472195f $X=0.93 $Y=2.26 $X2=0 $Y2=0
cc_292 N_SCE_c_287_n N_A_27_81#_c_380_n 0.0049247f $X=0.93 $Y=2.185 $X2=0 $Y2=0
cc_293 N_SCE_c_291_n N_A_27_81#_c_380_n 0.00187336f $X=0.93 $Y=2.26 $X2=0 $Y2=0
cc_294 N_SCE_c_285_n N_A_27_81#_c_380_n 0.0131931f $X=1.14 $Y=1.68 $X2=0 $Y2=0
cc_295 N_SCE_c_300_p N_A_27_81#_c_380_n 0.0289823f $X=1.18 $Y=1.68 $X2=0 $Y2=0
cc_296 N_SCE_c_287_n N_A_27_81#_c_381_n 0.0052595f $X=0.93 $Y=2.185 $X2=0 $Y2=0
cc_297 N_SCE_c_289_n N_A_27_81#_c_381_n 0.0197389f $X=1.285 $Y=2.26 $X2=0 $Y2=0
cc_298 N_SCE_c_291_n N_A_27_81#_c_381_n 0.00665722f $X=0.93 $Y=2.26 $X2=0 $Y2=0
cc_299 N_SCE_c_292_n N_A_27_81#_c_381_n 0.0124118f $X=2.185 $Y=1.76 $X2=0 $Y2=0
cc_300 N_SCE_c_285_n N_A_27_81#_c_381_n 0.00214308f $X=1.14 $Y=1.68 $X2=0 $Y2=0
cc_301 N_SCE_c_300_p N_A_27_81#_c_381_n 0.0988105f $X=1.18 $Y=1.68 $X2=0 $Y2=0
cc_302 N_SCE_c_292_n N_A_27_81#_c_382_n 0.00665224f $X=2.185 $Y=1.76 $X2=0 $Y2=0
cc_303 N_SCE_c_284_n N_A_27_81#_c_382_n 0.0023135f $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_304 N_SCE_c_287_n N_D_M1009_g 0.00285215f $X=0.93 $Y=2.185 $X2=0 $Y2=0
cc_305 N_SCE_c_289_n N_D_M1009_g 0.0627856f $X=1.285 $Y=2.26 $X2=0 $Y2=0
cc_306 N_SCE_c_292_n N_D_M1009_g 0.0126878f $X=2.185 $Y=1.76 $X2=0 $Y2=0
cc_307 N_SCE_c_282_n N_D_M1009_g 0.00485399f $X=2.27 $Y=1.675 $X2=0 $Y2=0
cc_308 N_SCE_c_285_n N_D_M1009_g 0.0111936f $X=1.14 $Y=1.68 $X2=0 $Y2=0
cc_309 N_SCE_c_286_n N_D_M1009_g 0.0038425f $X=1.345 $Y=1.68 $X2=0 $Y2=0
cc_310 N_SCE_M1024_g N_D_M1035_g 0.0189135f $X=2.355 $Y=0.615 $X2=0 $Y2=0
cc_311 N_SCE_c_283_n N_D_M1035_g 7.16447e-19 $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_312 N_SCE_c_284_n N_D_M1035_g 0.0159518f $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_313 N_SCE_c_292_n D 0.0172089f $X=2.185 $Y=1.76 $X2=0 $Y2=0
cc_314 N_SCE_c_283_n D 0.0140752f $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_315 N_SCE_c_284_n D 6.94216e-19 $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_316 N_SCE_c_292_n N_D_c_457_n 0.00776935f $X=2.185 $Y=1.76 $X2=0 $Y2=0
cc_317 N_SCE_c_282_n N_D_c_457_n 0.00208522f $X=2.27 $Y=1.675 $X2=0 $Y2=0
cc_318 N_SCE_c_283_n N_D_c_457_n 3.30599e-19 $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_319 N_SCE_c_284_n N_D_c_457_n 0.00308223f $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_320 N_SCE_M1024_g N_SCD_M1047_g 0.0337834f $X=2.355 $Y=0.615 $X2=0 $Y2=0
cc_321 N_SCE_c_282_n N_SCD_M1047_g 0.00329469f $X=2.27 $Y=1.675 $X2=0 $Y2=0
cc_322 N_SCE_c_283_n N_SCD_M1047_g 9.4742e-19 $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_323 N_SCE_c_284_n N_SCD_M1047_g 0.020319f $X=2.35 $Y=1.23 $X2=0 $Y2=0
cc_324 N_SCE_c_292_n SCD 0.0148609f $X=2.185 $Y=1.76 $X2=0 $Y2=0
cc_325 N_SCE_c_282_n SCD 0.00857017f $X=2.27 $Y=1.675 $X2=0 $Y2=0
cc_326 N_SCE_c_292_n N_SCD_c_499_n 0.0012705f $X=2.185 $Y=1.76 $X2=0 $Y2=0
cc_327 N_SCE_c_282_n N_SCD_c_499_n 4.64512e-19 $X=2.27 $Y=1.675 $X2=0 $Y2=0
cc_328 N_SCE_c_288_n N_VPWR_c_1702_n 0.00287644f $X=0.93 $Y=2.335 $X2=0 $Y2=0
cc_329 N_SCE_c_289_n N_VPWR_c_1702_n 0.00217652f $X=1.285 $Y=2.26 $X2=0 $Y2=0
cc_330 N_SCE_c_290_n N_VPWR_c_1702_n 0.0150882f $X=1.36 $Y=2.335 $X2=0 $Y2=0
cc_331 N_SCE_c_290_n N_VPWR_c_1712_n 0.00477554f $X=1.36 $Y=2.335 $X2=0 $Y2=0
cc_332 N_SCE_c_288_n N_VPWR_c_1718_n 0.00539298f $X=0.93 $Y=2.335 $X2=0 $Y2=0
cc_333 N_SCE_c_288_n N_VPWR_c_1701_n 0.0110783f $X=0.93 $Y=2.335 $X2=0 $Y2=0
cc_334 N_SCE_c_290_n N_VPWR_c_1701_n 0.00814835f $X=1.36 $Y=2.335 $X2=0 $Y2=0
cc_335 N_SCE_c_292_n N_A_359_489#_c_1916_n 6.62623e-19 $X=2.185 $Y=1.76 $X2=0
+ $Y2=0
cc_336 N_SCE_M1024_g N_A_359_489#_c_1902_n 0.00878302f $X=2.355 $Y=0.615 $X2=0
+ $Y2=0
cc_337 N_SCE_c_283_n N_A_359_489#_c_1902_n 0.0153366f $X=2.35 $Y=1.23 $X2=0
+ $Y2=0
cc_338 N_SCE_c_284_n N_A_359_489#_c_1902_n 0.00208514f $X=2.35 $Y=1.23 $X2=0
+ $Y2=0
cc_339 N_SCE_c_282_n N_A_359_489#_c_1903_n 0.00512949f $X=2.27 $Y=1.675 $X2=0
+ $Y2=0
cc_340 N_SCE_c_283_n N_A_359_489#_c_1903_n 0.00922968f $X=2.35 $Y=1.23 $X2=0
+ $Y2=0
cc_341 N_SCE_c_290_n N_A_359_489#_c_1912_n 0.00171137f $X=1.36 $Y=2.335 $X2=0
+ $Y2=0
cc_342 N_SCE_M1024_g N_A_359_489#_c_1905_n 0.00659604f $X=2.355 $Y=0.615 $X2=0
+ $Y2=0
cc_343 N_SCE_c_283_n N_A_359_489#_c_1905_n 0.00994922f $X=2.35 $Y=1.23 $X2=0
+ $Y2=0
cc_344 N_SCE_c_284_n N_A_359_489#_c_1905_n 0.00237833f $X=2.35 $Y=1.23 $X2=0
+ $Y2=0
cc_345 N_SCE_M1014_g N_VGND_c_2083_n 0.0138018f $X=0.475 $Y=0.615 $X2=0 $Y2=0
cc_346 N_SCE_M1024_g N_VGND_c_2094_n 9.29198e-19 $X=2.355 $Y=0.615 $X2=0 $Y2=0
cc_347 N_SCE_M1014_g N_VGND_c_2102_n 0.0045897f $X=0.475 $Y=0.615 $X2=0 $Y2=0
cc_348 N_SCE_M1014_g N_VGND_c_2113_n 0.0044912f $X=0.475 $Y=0.615 $X2=0 $Y2=0
cc_349 N_SCE_M1024_g N_noxref_25_c_2245_n 0.0111747f $X=2.355 $Y=0.615 $X2=0
+ $Y2=0
cc_350 N_SCE_M1024_g N_noxref_25_c_2247_n 9.61094e-19 $X=2.355 $Y=0.615 $X2=0
+ $Y2=0
cc_351 N_A_27_81#_M1041_g N_D_M1009_g 0.0151019f $X=2.15 $Y=2.765 $X2=0 $Y2=0
cc_352 N_A_27_81#_c_381_n N_D_M1009_g 0.0183983f $X=2.17 $Y=2.11 $X2=0 $Y2=0
cc_353 N_A_27_81#_c_382_n N_D_M1009_g 0.0217775f $X=2.17 $Y=2.11 $X2=0 $Y2=0
cc_354 N_A_27_81#_c_369_n N_D_M1035_g 0.0411497f $X=1.465 $Y=0.22 $X2=0 $Y2=0
cc_355 N_A_27_81#_c_375_n N_D_M1035_g 0.00279222f $X=1.09 $Y=1.1 $X2=0 $Y2=0
cc_356 N_A_27_81#_c_368_n D 4.91366e-19 $X=1.007 $Y=0.935 $X2=0 $Y2=0
cc_357 N_A_27_81#_c_371_n D 0.00436527f $X=1.54 $Y=0.295 $X2=0 $Y2=0
cc_358 N_A_27_81#_c_374_n D 0.0164132f $X=1.09 $Y=1.1 $X2=0 $Y2=0
cc_359 N_A_27_81#_c_375_n D 0.00102379f $X=1.09 $Y=1.1 $X2=0 $Y2=0
cc_360 N_A_27_81#_c_371_n N_D_c_457_n 0.00491941f $X=1.54 $Y=0.295 $X2=0 $Y2=0
cc_361 N_A_27_81#_c_374_n N_D_c_457_n 4.13577e-19 $X=1.09 $Y=1.1 $X2=0 $Y2=0
cc_362 N_A_27_81#_c_375_n N_D_c_457_n 0.0043203f $X=1.09 $Y=1.1 $X2=0 $Y2=0
cc_363 N_A_27_81#_M1041_g N_SCD_M1034_g 0.0370642f $X=2.15 $Y=2.765 $X2=0 $Y2=0
cc_364 N_A_27_81#_c_381_n N_SCD_c_501_n 2.97132e-19 $X=2.17 $Y=2.11 $X2=0 $Y2=0
cc_365 N_A_27_81#_c_382_n N_SCD_c_501_n 0.0212014f $X=2.17 $Y=2.11 $X2=0 $Y2=0
cc_366 N_A_27_81#_c_381_n SCD 0.0188951f $X=2.17 $Y=2.11 $X2=0 $Y2=0
cc_367 N_A_27_81#_c_382_n SCD 0.00261945f $X=2.17 $Y=2.11 $X2=0 $Y2=0
cc_368 N_A_27_81#_c_379_n N_VPWR_c_1702_n 0.0245928f $X=0.715 $Y=2.59 $X2=0
+ $Y2=0
cc_369 N_A_27_81#_c_381_n N_VPWR_c_1702_n 0.0212103f $X=2.17 $Y=2.11 $X2=0 $Y2=0
cc_370 N_A_27_81#_M1041_g N_VPWR_c_1703_n 0.00172486f $X=2.15 $Y=2.765 $X2=0
+ $Y2=0
cc_371 N_A_27_81#_M1041_g N_VPWR_c_1712_n 0.00412022f $X=2.15 $Y=2.765 $X2=0
+ $Y2=0
cc_372 N_A_27_81#_c_379_n N_VPWR_c_1718_n 0.0224804f $X=0.715 $Y=2.59 $X2=0
+ $Y2=0
cc_373 N_A_27_81#_M1021_s N_VPWR_c_1701_n 0.00212301f $X=0.59 $Y=2.445 $X2=0
+ $Y2=0
cc_374 N_A_27_81#_M1041_g N_VPWR_c_1701_n 0.00602177f $X=2.15 $Y=2.765 $X2=0
+ $Y2=0
cc_375 N_A_27_81#_c_379_n N_VPWR_c_1701_n 0.0133464f $X=0.715 $Y=2.59 $X2=0
+ $Y2=0
cc_376 N_A_27_81#_M1041_g N_A_359_489#_c_1916_n 0.00986508f $X=2.15 $Y=2.765
+ $X2=0 $Y2=0
cc_377 N_A_27_81#_c_381_n N_A_359_489#_c_1916_n 0.0141226f $X=2.17 $Y=2.11 $X2=0
+ $Y2=0
cc_378 N_A_27_81#_c_382_n N_A_359_489#_c_1916_n 0.00235362f $X=2.17 $Y=2.11
+ $X2=0 $Y2=0
cc_379 N_A_27_81#_M1041_g N_A_359_489#_c_1912_n 0.00877623f $X=2.15 $Y=2.765
+ $X2=0 $Y2=0
cc_380 N_A_27_81#_c_381_n N_A_359_489#_c_1912_n 0.0211919f $X=2.17 $Y=2.11 $X2=0
+ $Y2=0
cc_381 N_A_27_81#_c_382_n N_A_359_489#_c_1912_n 0.00145791f $X=2.17 $Y=2.11
+ $X2=0 $Y2=0
cc_382 N_A_27_81#_c_370_n N_VGND_c_2083_n 0.0105681f $X=1.125 $Y=0.22 $X2=0
+ $Y2=0
cc_383 N_A_27_81#_c_374_n N_VGND_c_2083_n 0.0257385f $X=1.09 $Y=1.1 $X2=0 $Y2=0
cc_384 N_A_27_81#_c_370_n N_VGND_c_2094_n 0.0187139f $X=1.125 $Y=0.22 $X2=0
+ $Y2=0
cc_385 N_A_27_81#_c_372_n N_VGND_c_2102_n 0.00746314f $X=0.26 $Y=0.63 $X2=0
+ $Y2=0
cc_386 N_A_27_81#_c_369_n N_VGND_c_2113_n 0.0136737f $X=1.465 $Y=0.22 $X2=0
+ $Y2=0
cc_387 N_A_27_81#_c_370_n N_VGND_c_2113_n 0.0157175f $X=1.125 $Y=0.22 $X2=0
+ $Y2=0
cc_388 N_A_27_81#_c_372_n N_VGND_c_2113_n 0.00884402f $X=0.26 $Y=0.63 $X2=0
+ $Y2=0
cc_389 N_A_27_81#_c_369_n N_noxref_25_c_2245_n 0.0017572f $X=1.465 $Y=0.22 $X2=0
+ $Y2=0
cc_390 N_A_27_81#_c_371_n N_noxref_25_c_2245_n 0.0071694f $X=1.54 $Y=0.295 $X2=0
+ $Y2=0
cc_391 N_A_27_81#_c_368_n N_noxref_25_c_2246_n 0.0127855f $X=1.007 $Y=0.935
+ $X2=0 $Y2=0
cc_392 N_A_27_81#_c_369_n N_noxref_25_c_2246_n 0.00736693f $X=1.465 $Y=0.22
+ $X2=0 $Y2=0
cc_393 N_A_27_81#_c_370_n N_noxref_25_c_2246_n 4.88574e-19 $X=1.125 $Y=0.22
+ $X2=0 $Y2=0
cc_394 N_A_27_81#_c_371_n N_noxref_25_c_2246_n 0.00719687f $X=1.54 $Y=0.295
+ $X2=0 $Y2=0
cc_395 N_A_27_81#_c_374_n N_noxref_25_c_2246_n 0.0113779f $X=1.09 $Y=1.1 $X2=0
+ $Y2=0
cc_396 N_A_27_81#_c_375_n N_noxref_25_c_2246_n 0.00250745f $X=1.09 $Y=1.1 $X2=0
+ $Y2=0
cc_397 N_D_M1009_g N_VPWR_c_1702_n 0.00289588f $X=1.72 $Y=2.765 $X2=0 $Y2=0
cc_398 N_D_M1009_g N_VPWR_c_1712_n 0.00539298f $X=1.72 $Y=2.765 $X2=0 $Y2=0
cc_399 N_D_M1009_g N_VPWR_c_1701_n 0.00984182f $X=1.72 $Y=2.765 $X2=0 $Y2=0
cc_400 N_D_M1009_g N_A_359_489#_c_1912_n 0.0105578f $X=1.72 $Y=2.765 $X2=0 $Y2=0
cc_401 N_D_M1035_g N_A_359_489#_c_1905_n 0.00150345f $X=1.9 $Y=0.615 $X2=0 $Y2=0
cc_402 D N_A_359_489#_c_1905_n 0.0101404f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_403 N_D_M1035_g N_VGND_c_2094_n 9.29198e-19 $X=1.9 $Y=0.615 $X2=0 $Y2=0
cc_404 N_D_M1035_g N_noxref_25_c_2245_n 0.0143897f $X=1.9 $Y=0.615 $X2=0 $Y2=0
cc_405 D N_noxref_25_c_2245_n 0.00669514f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_406 N_D_M1035_g N_noxref_25_c_2246_n 0.00107357f $X=1.9 $Y=0.615 $X2=0 $Y2=0
cc_407 N_SCD_M1034_g N_RESET_B_M1002_g 0.0218998f $X=2.62 $Y=2.765 $X2=0 $Y2=0
cc_408 N_SCD_c_502_n N_RESET_B_M1002_g 0.0125361f $X=2.71 $Y=2.275 $X2=0 $Y2=0
cc_409 N_SCD_M1047_g N_RESET_B_M1015_g 0.0486452f $X=2.8 $Y=0.615 $X2=0 $Y2=0
cc_410 N_SCD_c_501_n N_RESET_B_c_875_n 0.0125361f $X=2.71 $Y=2.11 $X2=0 $Y2=0
cc_411 SCD N_RESET_B_c_875_n 3.63672e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_412 N_SCD_M1034_g N_VPWR_c_1703_n 0.00981324f $X=2.62 $Y=2.765 $X2=0 $Y2=0
cc_413 N_SCD_M1034_g N_VPWR_c_1712_n 0.00351296f $X=2.62 $Y=2.765 $X2=0 $Y2=0
cc_414 N_SCD_M1034_g N_VPWR_c_1701_n 0.00434205f $X=2.62 $Y=2.765 $X2=0 $Y2=0
cc_415 N_SCD_M1034_g N_A_359_489#_c_1916_n 0.0141655f $X=2.62 $Y=2.765 $X2=0
+ $Y2=0
cc_416 N_SCD_c_502_n N_A_359_489#_c_1916_n 0.00364809f $X=2.71 $Y=2.275 $X2=0
+ $Y2=0
cc_417 SCD N_A_359_489#_c_1916_n 0.0191084f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_418 N_SCD_M1047_g N_A_359_489#_c_1902_n 0.0142126f $X=2.8 $Y=0.615 $X2=0
+ $Y2=0
cc_419 SCD N_A_359_489#_c_1902_n 0.00911823f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_420 N_SCD_c_499_n N_A_359_489#_c_1902_n 8.50781e-19 $X=2.71 $Y=1.77 $X2=0
+ $Y2=0
cc_421 N_SCD_M1034_g N_A_359_489#_c_1903_n 0.00321899f $X=2.62 $Y=2.765 $X2=0
+ $Y2=0
cc_422 N_SCD_M1047_g N_A_359_489#_c_1903_n 0.0129262f $X=2.8 $Y=0.615 $X2=0
+ $Y2=0
cc_423 SCD N_A_359_489#_c_1903_n 0.0525844f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_424 N_SCD_M1034_g N_A_359_489#_c_1912_n 0.00158635f $X=2.62 $Y=2.765 $X2=0
+ $Y2=0
cc_425 N_SCD_M1047_g N_A_359_489#_c_1905_n 9.65228e-19 $X=2.8 $Y=0.615 $X2=0
+ $Y2=0
cc_426 N_SCD_M1034_g N_A_359_489#_c_1913_n 6.14712e-19 $X=2.62 $Y=2.765 $X2=0
+ $Y2=0
cc_427 N_SCD_M1047_g N_VGND_c_2094_n 9.22791e-19 $X=2.8 $Y=0.615 $X2=0 $Y2=0
cc_428 N_SCD_M1047_g N_noxref_25_c_2245_n 0.00860433f $X=2.8 $Y=0.615 $X2=0
+ $Y2=0
cc_429 N_SCD_M1047_g N_noxref_25_c_2247_n 0.00651957f $X=2.8 $Y=0.615 $X2=0
+ $Y2=0
cc_430 N_CLK_c_542_n N_A_934_367#_c_597_n 9.16491e-19 $X=4.15 $Y=1.09 $X2=0
+ $Y2=0
cc_431 N_CLK_c_541_n N_RESET_B_M1015_g 0.0313802f $X=3.72 $Y=1.09 $X2=0 $Y2=0
cc_432 CLK N_RESET_B_M1015_g 0.00727528f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_433 N_CLK_c_541_n N_RESET_B_c_859_n 0.0104164f $X=3.72 $Y=1.09 $X2=0 $Y2=0
cc_434 N_CLK_c_542_n N_RESET_B_c_859_n 0.0100709f $X=4.15 $Y=1.09 $X2=0 $Y2=0
cc_435 N_CLK_M1042_g N_RESET_B_c_869_n 0.0014525f $X=4.165 $Y=2.465 $X2=0 $Y2=0
cc_436 CLK N_RESET_B_c_869_n 0.00825278f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_437 CLK N_RESET_B_c_870_n 0.00868781f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_438 N_CLK_M1042_g N_RESET_B_c_875_n 0.00551271f $X=4.165 $Y=2.465 $X2=0 $Y2=0
cc_439 CLK N_RESET_B_c_875_n 0.00837137f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_440 N_CLK_c_545_n N_RESET_B_c_875_n 4.73007e-19 $X=4.165 $Y=1.35 $X2=0 $Y2=0
cc_441 N_CLK_M1042_g N_RESET_B_c_876_n 3.94636e-19 $X=4.165 $Y=2.465 $X2=0 $Y2=0
cc_442 CLK N_RESET_B_c_876_n 0.0272562f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_443 N_CLK_M1042_g N_A_759_119#_M1017_g 0.0344039f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_444 N_CLK_c_542_n N_A_759_119#_c_1177_n 0.0145683f $X=4.15 $Y=1.09 $X2=0
+ $Y2=0
cc_445 CLK N_A_759_119#_c_1181_n 3.28545e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_446 N_CLK_c_545_n N_A_759_119#_c_1181_n 0.0396442f $X=4.165 $Y=1.35 $X2=0
+ $Y2=0
cc_447 N_CLK_c_542_n N_A_759_119#_c_1186_n 0.0100171f $X=4.15 $Y=1.09 $X2=0
+ $Y2=0
cc_448 CLK N_A_759_119#_c_1186_n 0.00864121f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_449 N_CLK_c_545_n N_A_759_119#_c_1186_n 7.13623e-19 $X=4.165 $Y=1.35 $X2=0
+ $Y2=0
cc_450 N_CLK_M1042_g N_A_759_119#_c_1209_n 0.00937349f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_451 CLK N_A_759_119#_c_1209_n 0.0038223f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_452 N_CLK_c_542_n N_A_759_119#_c_1187_n 0.00114317f $X=4.15 $Y=1.09 $X2=0
+ $Y2=0
cc_453 CLK N_A_759_119#_c_1187_n 0.00551376f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_454 N_CLK_c_545_n N_A_759_119#_c_1187_n 0.00372673f $X=4.165 $Y=1.35 $X2=0
+ $Y2=0
cc_455 N_CLK_M1042_g N_A_759_119#_c_1188_n 0.00482146f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_456 CLK N_A_759_119#_c_1188_n 0.0110653f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_c_541_n N_A_759_119#_c_1189_n 5.09956e-19 $X=3.72 $Y=1.09 $X2=0
+ $Y2=0
cc_458 CLK N_A_759_119#_c_1189_n 0.0217774f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_459 N_CLK_c_545_n N_A_759_119#_c_1189_n 0.00291001f $X=4.165 $Y=1.35 $X2=0
+ $Y2=0
cc_460 N_CLK_M1042_g N_A_759_119#_c_1219_n 0.00532702f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_461 CLK N_A_759_119#_c_1219_n 0.0161145f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_462 N_CLK_c_545_n N_A_759_119#_c_1219_n 0.00106503f $X=4.165 $Y=1.35 $X2=0
+ $Y2=0
cc_463 CLK N_A_759_119#_c_1190_n 0.0282424f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_464 N_CLK_c_545_n N_A_759_119#_c_1190_n 0.00272106f $X=4.165 $Y=1.35 $X2=0
+ $Y2=0
cc_465 N_CLK_M1042_g N_VPWR_c_1704_n 0.0113322f $X=4.165 $Y=2.465 $X2=0 $Y2=0
cc_466 N_CLK_M1042_g N_VPWR_c_1714_n 0.00358332f $X=4.165 $Y=2.465 $X2=0 $Y2=0
cc_467 N_CLK_M1042_g N_VPWR_c_1701_n 0.00567344f $X=4.165 $Y=2.465 $X2=0 $Y2=0
cc_468 CLK N_A_359_489#_c_1903_n 0.0454064f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_469 N_CLK_M1042_g N_A_359_489#_c_1907_n 0.014627f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_470 N_CLK_M1042_g N_A_359_489#_c_1913_n 0.00816322f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_471 N_CLK_c_541_n N_VGND_c_2084_n 0.00291051f $X=3.72 $Y=1.09 $X2=0 $Y2=0
cc_472 CLK N_VGND_c_2084_n 0.0112098f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_473 N_CLK_c_542_n N_VGND_c_2085_n 0.00268637f $X=4.15 $Y=1.09 $X2=0 $Y2=0
cc_474 N_CLK_c_541_n N_VGND_c_2113_n 9.39239e-19 $X=3.72 $Y=1.09 $X2=0 $Y2=0
cc_475 N_CLK_c_542_n N_VGND_c_2113_n 9.39239e-19 $X=4.15 $Y=1.09 $X2=0 $Y2=0
cc_476 N_A_934_367#_c_615_p N_A_1290_365#_M1005_d 0.0195983f $X=8.67 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_477 N_A_934_367#_c_594_n N_A_1290_365#_M1036_g 0.00120763f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_478 N_A_934_367#_M1028_g N_A_1290_365#_M1036_g 0.0664358f $X=6.67 $Y=0.805
+ $X2=0 $Y2=0
cc_479 N_A_934_367#_c_598_n N_A_1290_365#_M1036_g 0.00533349f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_480 N_A_934_367#_c_600_n N_A_1290_365#_M1036_g 0.00423197f $X=7.335 $Y=0.72
+ $X2=0 $Y2=0
cc_481 N_A_934_367#_c_620_p N_A_1290_365#_M1036_g 0.0021697f $X=7.425 $Y=0.805
+ $X2=0 $Y2=0
cc_482 N_A_934_367#_c_594_n N_A_1290_365#_c_782_n 0.0062266f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_483 N_A_934_367#_M1028_g N_A_1290_365#_c_782_n 0.00312215f $X=6.67 $Y=0.805
+ $X2=0 $Y2=0
cc_484 N_A_934_367#_M1038_g N_A_1290_365#_c_789_n 0.00450248f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_485 N_A_934_367#_c_594_n N_A_1290_365#_c_789_n 0.0175679f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_486 N_A_934_367#_c_598_n N_A_1290_365#_c_783_n 0.0134883f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_487 N_A_934_367#_c_615_p N_A_1290_365#_c_783_n 0.0580688f $X=8.67 $Y=0.805
+ $X2=0 $Y2=0
cc_488 N_A_934_367#_c_620_p N_A_1290_365#_c_783_n 0.0114695f $X=7.425 $Y=0.805
+ $X2=0 $Y2=0
cc_489 N_A_934_367#_M1028_g N_A_1290_365#_c_784_n 0.00808363f $X=6.67 $Y=0.805
+ $X2=0 $Y2=0
cc_490 N_A_934_367#_c_598_n N_A_1290_365#_c_784_n 0.00506646f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_491 N_A_934_367#_c_615_p N_A_1290_365#_c_807_n 0.0203396f $X=8.67 $Y=0.805
+ $X2=0 $Y2=0
cc_492 N_A_934_367#_c_601_n N_A_1290_365#_c_807_n 0.0146055f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_493 N_A_934_367#_c_602_n N_A_1290_365#_c_807_n 0.00151433f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_494 N_A_934_367#_c_601_n N_A_1290_365#_c_785_n 0.0368125f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_495 N_A_934_367#_c_602_n N_A_1290_365#_c_785_n 0.00178362f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_496 N_A_934_367#_c_609_n N_A_1290_365#_c_785_n 0.0163962f $X=9.07 $Y=1.8
+ $X2=0 $Y2=0
cc_497 N_A_934_367#_M1028_g N_RESET_B_c_859_n 0.00880557f $X=6.67 $Y=0.805 $X2=0
+ $Y2=0
cc_498 N_A_934_367#_c_597_n N_RESET_B_c_859_n 0.00497606f $X=4.915 $Y=0.785
+ $X2=0 $Y2=0
cc_499 N_A_934_367#_c_598_n N_RESET_B_c_859_n 0.0259217f $X=7.245 $Y=0.395 $X2=0
+ $Y2=0
cc_500 N_A_934_367#_c_599_n N_RESET_B_c_859_n 0.00410689f $X=5.77 $Y=0.395 $X2=0
+ $Y2=0
cc_501 N_A_934_367#_c_598_n N_RESET_B_M1025_g 0.00783098f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_502 N_A_934_367#_c_600_n N_RESET_B_M1025_g 0.00657266f $X=7.335 $Y=0.72 $X2=0
+ $Y2=0
cc_503 N_A_934_367#_c_615_p N_RESET_B_M1025_g 0.00527029f $X=8.67 $Y=0.805 $X2=0
+ $Y2=0
cc_504 N_A_934_367#_c_620_p N_RESET_B_M1025_g 0.00392911f $X=7.425 $Y=0.805
+ $X2=0 $Y2=0
cc_505 N_A_934_367#_M1017_d N_RESET_B_c_869_n 2.61106e-19 $X=4.67 $Y=1.835 $X2=0
+ $Y2=0
cc_506 N_A_934_367#_c_594_n N_RESET_B_c_869_n 0.00319163f $X=6.42 $Y=1.525 $X2=0
+ $Y2=0
cc_507 N_A_934_367#_c_603_n N_RESET_B_c_869_n 0.0475782f $X=5.535 $Y=1.615 $X2=0
+ $Y2=0
cc_508 N_A_934_367#_c_608_n N_RESET_B_c_871_n 0.00707824f $X=9.275 $Y=1.8 $X2=0
+ $Y2=0
cc_509 N_A_934_367#_c_609_n N_RESET_B_c_871_n 0.0120493f $X=9.07 $Y=1.8 $X2=0
+ $Y2=0
cc_510 N_A_934_367#_c_611_n N_RESET_B_c_871_n 0.0188789f $X=9.435 $Y=1.8 $X2=0
+ $Y2=0
cc_511 N_A_934_367#_c_612_n N_RESET_B_c_871_n 0.00242448f $X=9.44 $Y=2.155 $X2=0
+ $Y2=0
cc_512 N_A_934_367#_c_600_n N_A_1162_463#_M1005_g 8.33316e-19 $X=7.335 $Y=0.72
+ $X2=0 $Y2=0
cc_513 N_A_934_367#_c_615_p N_A_1162_463#_M1005_g 0.0151336f $X=8.67 $Y=0.805
+ $X2=0 $Y2=0
cc_514 N_A_934_367#_c_601_n N_A_1162_463#_M1005_g 0.00157589f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_515 N_A_934_367#_c_602_n N_A_1162_463#_M1005_g 0.00477661f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_516 N_A_934_367#_c_605_n N_A_1162_463#_M1005_g 0.0189426f $X=8.87 $Y=1.09
+ $X2=0 $Y2=0
cc_517 N_A_934_367#_M1038_g N_A_1162_463#_c_1069_n 0.00536908f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_518 N_A_934_367#_c_594_n N_A_1162_463#_c_1069_n 0.00201046f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_519 N_A_934_367#_M1038_g N_A_1162_463#_c_1064_n 0.00146087f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_520 N_A_934_367#_c_594_n N_A_1162_463#_c_1064_n 0.0150823f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_521 N_A_934_367#_M1028_g N_A_1162_463#_c_1064_n 0.00741987f $X=6.67 $Y=0.805
+ $X2=0 $Y2=0
cc_522 N_A_934_367#_c_594_n N_A_1162_463#_c_1083_n 0.0032984f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_523 N_A_934_367#_M1028_g N_A_1162_463#_c_1083_n 0.00578597f $X=6.67 $Y=0.805
+ $X2=0 $Y2=0
cc_524 N_A_934_367#_c_598_n N_A_1162_463#_c_1083_n 0.0201656f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_525 N_A_934_367#_c_600_n N_A_1162_463#_c_1083_n 0.00181535f $X=7.335 $Y=0.72
+ $X2=0 $Y2=0
cc_526 N_A_934_367#_c_620_p N_A_1162_463#_c_1083_n 0.00499642f $X=7.425 $Y=0.805
+ $X2=0 $Y2=0
cc_527 N_A_934_367#_c_602_n N_A_1162_463#_c_1066_n 3.17528e-19 $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_528 N_A_934_367#_c_603_n N_A_759_119#_M1017_g 0.00282708f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_529 N_A_934_367#_c_597_n N_A_759_119#_c_1177_n 0.00688984f $X=4.915 $Y=0.785
+ $X2=0 $Y2=0
cc_530 N_A_934_367#_c_603_n N_A_759_119#_c_1177_n 8.79431e-19 $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_531 N_A_934_367#_M1038_g N_A_759_119#_c_1178_n 0.0193058f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_532 N_A_934_367#_c_603_n N_A_759_119#_c_1178_n 0.0244517f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_533 N_A_934_367#_c_596_n N_A_759_119#_c_1179_n 0.00311645f $X=4.93 $Y=1.05
+ $X2=0 $Y2=0
cc_534 N_A_934_367#_c_597_n N_A_759_119#_c_1179_n 0.00764845f $X=4.915 $Y=0.785
+ $X2=0 $Y2=0
cc_535 N_A_934_367#_c_603_n N_A_759_119#_c_1179_n 0.00723411f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_536 N_A_934_367#_M1038_g N_A_759_119#_c_1193_n 0.0103532f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_537 N_A_934_367#_c_598_n N_A_759_119#_c_1180_n 0.00409015f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_538 N_A_934_367#_c_603_n N_A_759_119#_c_1180_n 0.0258738f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_539 N_A_934_367#_c_604_n N_A_759_119#_c_1180_n 0.0633344f $X=5.81 $Y=1.615
+ $X2=0 $Y2=0
cc_540 N_A_934_367#_c_603_n N_A_759_119#_c_1181_n 0.0408393f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_541 N_A_934_367#_c_604_n N_A_759_119#_c_1181_n 0.0214278f $X=5.81 $Y=1.615
+ $X2=0 $Y2=0
cc_542 N_A_934_367#_M1038_g N_A_759_119#_M1023_g 0.0135072f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_543 N_A_934_367#_c_594_n N_A_759_119#_M1023_g 0.00280988f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_544 N_A_934_367#_M1028_g N_A_759_119#_c_1182_n 0.0174663f $X=6.67 $Y=0.805
+ $X2=0 $Y2=0
cc_545 N_A_934_367#_c_596_n N_A_759_119#_c_1182_n 0.00478106f $X=4.93 $Y=1.05
+ $X2=0 $Y2=0
cc_546 N_A_934_367#_c_598_n N_A_759_119#_c_1182_n 0.00709841f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_547 N_A_934_367#_c_609_n N_A_759_119#_M1010_g 0.00676711f $X=9.07 $Y=1.8
+ $X2=0 $Y2=0
cc_548 N_A_934_367#_c_611_n N_A_759_119#_M1010_g 0.00293206f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_549 N_A_934_367#_c_612_n N_A_759_119#_M1010_g 0.016892f $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_550 N_A_934_367#_c_601_n N_A_759_119#_c_1183_n 0.00689232f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_551 N_A_934_367#_c_608_n N_A_759_119#_c_1183_n 0.011713f $X=9.275 $Y=1.8
+ $X2=0 $Y2=0
cc_552 N_A_934_367#_c_609_n N_A_759_119#_c_1183_n 0.00530766f $X=9.07 $Y=1.8
+ $X2=0 $Y2=0
cc_553 N_A_934_367#_c_611_n N_A_759_119#_c_1183_n 0.00449236f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_554 N_A_934_367#_c_612_n N_A_759_119#_c_1183_n 0.0078491f $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_555 N_A_934_367#_c_601_n N_A_759_119#_c_1184_n 0.00224126f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_556 N_A_934_367#_c_602_n N_A_759_119#_c_1184_n 0.0216823f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_557 N_A_934_367#_c_609_n N_A_759_119#_c_1184_n 0.00133531f $X=9.07 $Y=1.8
+ $X2=0 $Y2=0
cc_558 N_A_934_367#_c_615_p N_A_759_119#_M1040_g 6.42287e-19 $X=8.67 $Y=0.805
+ $X2=0 $Y2=0
cc_559 N_A_934_367#_c_601_n N_A_759_119#_M1040_g 0.00605019f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_560 N_A_934_367#_c_602_n N_A_759_119#_M1040_g 0.0213206f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_561 N_A_934_367#_c_605_n N_A_759_119#_M1040_g 0.0222411f $X=8.87 $Y=1.09
+ $X2=0 $Y2=0
cc_562 N_A_934_367#_c_597_n N_A_759_119#_c_1186_n 0.0105597f $X=4.915 $Y=0.785
+ $X2=0 $Y2=0
cc_563 N_A_934_367#_c_603_n N_A_759_119#_c_1209_n 0.00495768f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_564 N_A_934_367#_c_597_n N_A_759_119#_c_1187_n 4.98226e-19 $X=4.915 $Y=0.785
+ $X2=0 $Y2=0
cc_565 N_A_934_367#_c_603_n N_A_759_119#_c_1187_n 0.0102513f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_566 N_A_934_367#_c_603_n N_A_759_119#_c_1188_n 0.0103659f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_567 N_A_934_367#_c_603_n N_A_759_119#_c_1219_n 0.00286477f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_568 N_A_934_367#_c_603_n N_A_759_119#_c_1190_n 0.0339138f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_569 N_A_934_367#_M1032_g N_A_1923_174#_M1001_g 0.0197349f $X=9.35 $Y=2.69
+ $X2=0 $Y2=0
cc_570 N_A_934_367#_c_611_n N_A_1923_174#_M1001_g 0.0021312f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_571 N_A_934_367#_c_612_n N_A_1923_174#_M1001_g 0.0211427f $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_572 N_A_934_367#_c_615_p N_A_1770_412#_M1046_d 0.00338754f $X=8.67 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_573 N_A_934_367#_M1032_g N_A_1770_412#_c_1485_n 0.00214551f $X=9.35 $Y=2.69
+ $X2=0 $Y2=0
cc_574 N_A_934_367#_c_608_n N_A_1770_412#_c_1485_n 0.00207485f $X=9.275 $Y=1.8
+ $X2=0 $Y2=0
cc_575 N_A_934_367#_c_609_n N_A_1770_412#_c_1485_n 0.0155677f $X=9.07 $Y=1.8
+ $X2=0 $Y2=0
cc_576 N_A_934_367#_c_611_n N_A_1770_412#_c_1485_n 0.0182209f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_577 N_A_934_367#_c_612_n N_A_1770_412#_c_1485_n 9.03822e-19 $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_578 N_A_934_367#_M1032_g N_A_1770_412#_c_1490_n 0.0121679f $X=9.35 $Y=2.69
+ $X2=0 $Y2=0
cc_579 N_A_934_367#_c_608_n N_A_1770_412#_c_1490_n 0.00112603f $X=9.275 $Y=1.8
+ $X2=0 $Y2=0
cc_580 N_A_934_367#_c_611_n N_A_1770_412#_c_1490_n 0.0213289f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_581 N_A_934_367#_c_612_n N_A_1770_412#_c_1490_n 0.00145528f $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_582 N_A_934_367#_c_615_p N_A_1770_412#_c_1468_n 0.0133632f $X=8.67 $Y=0.805
+ $X2=0 $Y2=0
cc_583 N_A_934_367#_c_601_n N_A_1770_412#_c_1468_n 0.0317087f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_584 N_A_934_367#_c_602_n N_A_1770_412#_c_1468_n 7.48445e-19 $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_585 N_A_934_367#_c_605_n N_A_1770_412#_c_1468_n 0.00120386f $X=8.87 $Y=1.09
+ $X2=0 $Y2=0
cc_586 N_A_934_367#_c_611_n N_A_1770_412#_c_1469_n 0.00722534f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_587 N_A_934_367#_c_612_n N_A_1770_412#_c_1469_n 9.23168e-19 $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_588 N_A_934_367#_c_601_n N_A_1770_412#_c_1470_n 0.0150915f $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_589 N_A_934_367#_c_602_n N_A_1770_412#_c_1470_n 2.09021e-19 $X=8.87 $Y=1.255
+ $X2=0 $Y2=0
cc_590 N_A_934_367#_c_608_n N_A_1770_412#_c_1470_n 0.00251706f $X=9.275 $Y=1.8
+ $X2=0 $Y2=0
cc_591 N_A_934_367#_c_611_n N_A_1770_412#_c_1470_n 0.0140949f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_592 N_A_934_367#_c_612_n N_A_1770_412#_c_1470_n 2.72876e-19 $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_593 N_A_934_367#_M1032_g N_A_1770_412#_c_1479_n 0.0013796f $X=9.35 $Y=2.69
+ $X2=0 $Y2=0
cc_594 N_A_934_367#_c_611_n N_A_1770_412#_c_1479_n 0.0380275f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_595 N_A_934_367#_c_612_n N_A_1770_412#_c_1479_n 0.0016233f $X=9.44 $Y=2.155
+ $X2=0 $Y2=0
cc_596 N_A_934_367#_M1032_g N_A_1770_412#_c_1481_n 0.00592655f $X=9.35 $Y=2.69
+ $X2=0 $Y2=0
cc_597 N_A_934_367#_c_608_n N_A_1770_412#_c_1481_n 6.71205e-19 $X=9.275 $Y=1.8
+ $X2=0 $Y2=0
cc_598 N_A_934_367#_c_615_p N_A_1770_412#_c_1472_n 0.00419414f $X=8.67 $Y=0.805
+ $X2=0 $Y2=0
cc_599 N_A_934_367#_c_605_n N_A_1770_412#_c_1472_n 0.0106001f $X=8.87 $Y=1.09
+ $X2=0 $Y2=0
cc_600 N_A_934_367#_c_611_n N_A_1770_412#_c_1473_n 0.00428371f $X=9.435 $Y=1.8
+ $X2=0 $Y2=0
cc_601 N_A_934_367#_M1032_g N_VPWR_c_1720_n 0.00412011f $X=9.35 $Y=2.69 $X2=0
+ $Y2=0
cc_602 N_A_934_367#_M1032_g N_VPWR_c_1727_n 0.00363377f $X=9.35 $Y=2.69 $X2=0
+ $Y2=0
cc_603 N_A_934_367#_M1017_d N_VPWR_c_1701_n 0.00323595f $X=4.67 $Y=1.835 $X2=0
+ $Y2=0
cc_604 N_A_934_367#_M1038_g N_VPWR_c_1701_n 9.39239e-19 $X=5.735 $Y=2.525 $X2=0
+ $Y2=0
cc_605 N_A_934_367#_M1032_g N_VPWR_c_1701_n 0.00526787f $X=9.35 $Y=2.69 $X2=0
+ $Y2=0
cc_606 N_A_934_367#_M1017_d N_A_359_489#_c_1907_n 0.00590858f $X=4.67 $Y=1.835
+ $X2=0 $Y2=0
cc_607 N_A_934_367#_c_603_n N_A_359_489#_c_1907_n 0.0284549f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_608 N_A_934_367#_M1038_g N_A_359_489#_c_1909_n 0.0168153f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_609 N_A_934_367#_c_594_n N_A_359_489#_c_1909_n 0.00364701f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_610 N_A_934_367#_c_603_n N_A_359_489#_c_1909_n 0.0100259f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_611 N_A_934_367#_c_604_n N_A_359_489#_c_1909_n 2.4455e-19 $X=5.81 $Y=1.615
+ $X2=0 $Y2=0
cc_612 N_A_934_367#_c_603_n N_A_359_489#_c_1910_n 0.0271413f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_613 N_A_934_367#_c_604_n N_A_359_489#_c_1910_n 0.00185657f $X=5.81 $Y=1.615
+ $X2=0 $Y2=0
cc_614 N_A_934_367#_c_594_n N_A_359_489#_c_1904_n 0.011781f $X=6.42 $Y=1.525
+ $X2=0 $Y2=0
cc_615 N_A_934_367#_c_596_n N_A_359_489#_c_1904_n 0.0314775f $X=4.93 $Y=1.05
+ $X2=0 $Y2=0
cc_616 N_A_934_367#_c_598_n N_A_359_489#_c_1904_n 0.013115f $X=7.245 $Y=0.395
+ $X2=0 $Y2=0
cc_617 N_A_934_367#_c_603_n N_A_359_489#_c_1904_n 0.0562403f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_618 N_A_934_367#_c_604_n N_A_359_489#_c_1904_n 0.00922181f $X=5.81 $Y=1.615
+ $X2=0 $Y2=0
cc_619 N_A_934_367#_c_603_n N_A_359_489#_c_1914_n 5.1233e-19 $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_620 N_A_934_367#_M1038_g N_A_359_489#_c_1915_n 0.0031255f $X=5.735 $Y=2.525
+ $X2=0 $Y2=0
cc_621 N_A_934_367#_c_603_n N_A_359_489#_c_1915_n 0.00998569f $X=5.535 $Y=1.615
+ $X2=0 $Y2=0
cc_622 N_A_934_367#_c_615_p N_VGND_M1025_d 0.0121283f $X=8.67 $Y=0.805 $X2=0
+ $Y2=0
cc_623 N_A_934_367#_c_596_n N_VGND_c_2086_n 0.0315509f $X=4.93 $Y=1.05 $X2=0
+ $Y2=0
cc_624 N_A_934_367#_c_599_n N_VGND_c_2086_n 0.0143582f $X=5.77 $Y=0.395 $X2=0
+ $Y2=0
cc_625 N_A_934_367#_c_603_n N_VGND_c_2086_n 0.0154417f $X=5.535 $Y=1.615 $X2=0
+ $Y2=0
cc_626 N_A_934_367#_c_598_n N_VGND_c_2087_n 0.0140539f $X=7.245 $Y=0.395 $X2=0
+ $Y2=0
cc_627 N_A_934_367#_c_600_n N_VGND_c_2087_n 0.0051663f $X=7.335 $Y=0.72 $X2=0
+ $Y2=0
cc_628 N_A_934_367#_c_615_p N_VGND_c_2087_n 0.0256243f $X=8.67 $Y=0.805 $X2=0
+ $Y2=0
cc_629 N_A_934_367#_c_597_n N_VGND_c_2098_n 0.005425f $X=4.915 $Y=0.785 $X2=0
+ $Y2=0
cc_630 N_A_934_367#_c_615_p N_VGND_c_2100_n 0.0122049f $X=8.67 $Y=0.805 $X2=0
+ $Y2=0
cc_631 N_A_934_367#_c_605_n N_VGND_c_2100_n 0.00394604f $X=8.87 $Y=1.09 $X2=0
+ $Y2=0
cc_632 N_A_934_367#_c_598_n N_VGND_c_2103_n 0.0797017f $X=7.245 $Y=0.395 $X2=0
+ $Y2=0
cc_633 N_A_934_367#_c_599_n N_VGND_c_2103_n 0.00902328f $X=5.77 $Y=0.395 $X2=0
+ $Y2=0
cc_634 N_A_934_367#_c_615_p N_VGND_c_2103_n 0.00203983f $X=8.67 $Y=0.805 $X2=0
+ $Y2=0
cc_635 N_A_934_367#_c_597_n N_VGND_c_2113_n 0.00854487f $X=4.915 $Y=0.785 $X2=0
+ $Y2=0
cc_636 N_A_934_367#_c_598_n N_VGND_c_2113_n 0.0536088f $X=7.245 $Y=0.395 $X2=0
+ $Y2=0
cc_637 N_A_934_367#_c_599_n N_VGND_c_2113_n 0.00574501f $X=5.77 $Y=0.395 $X2=0
+ $Y2=0
cc_638 N_A_934_367#_c_615_p N_VGND_c_2113_n 0.0360116f $X=8.67 $Y=0.805 $X2=0
+ $Y2=0
cc_639 N_A_934_367#_c_605_n N_VGND_c_2113_n 0.00513096f $X=8.87 $Y=1.09 $X2=0
+ $Y2=0
cc_640 N_A_934_367#_c_600_n A_1421_119# 0.0016103f $X=7.335 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_641 N_A_934_367#_c_620_p A_1421_119# 0.00265301f $X=7.425 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_642 N_A_1290_365#_M1036_g N_RESET_B_c_859_n 0.00880557f $X=7.03 $Y=0.805
+ $X2=0 $Y2=0
cc_643 N_A_1290_365#_M1036_g N_RESET_B_M1025_g 0.0444002f $X=7.03 $Y=0.805 $X2=0
+ $Y2=0
cc_644 N_A_1290_365#_c_783_n N_RESET_B_M1025_g 0.0113305f $X=8.31 $Y=1.147 $X2=0
+ $Y2=0
cc_645 N_A_1290_365#_c_782_n N_RESET_B_c_869_n 0.0129164f $X=6.705 $Y=1.99 $X2=0
+ $Y2=0
cc_646 N_A_1290_365#_c_789_n N_RESET_B_c_869_n 0.0145122f $X=6.705 $Y=1.99 $X2=0
+ $Y2=0
cc_647 N_A_1290_365#_M1031_d N_RESET_B_c_871_n 0.00524882f $X=8.275 $Y=1.895
+ $X2=0 $Y2=0
cc_648 N_A_1290_365#_c_819_p N_RESET_B_c_871_n 0.0202585f $X=8.47 $Y=2.24 $X2=0
+ $Y2=0
cc_649 N_A_1290_365#_c_785_n N_RESET_B_c_871_n 0.0242004f $X=8.47 $Y=2.08 $X2=0
+ $Y2=0
cc_650 N_A_1290_365#_c_789_n N_RESET_B_c_873_n 3.5882e-19 $X=6.705 $Y=1.99 $X2=0
+ $Y2=0
cc_651 N_A_1290_365#_M1000_g N_RESET_B_c_877_n 0.0122779f $X=6.525 $Y=2.525
+ $X2=0 $Y2=0
cc_652 N_A_1290_365#_c_789_n N_RESET_B_c_877_n 0.0545067f $X=6.705 $Y=1.99 $X2=0
+ $Y2=0
cc_653 N_A_1290_365#_c_783_n N_A_1162_463#_M1005_g 0.0136689f $X=8.31 $Y=1.147
+ $X2=0 $Y2=0
cc_654 N_A_1290_365#_c_785_n N_A_1162_463#_M1005_g 0.00436612f $X=8.47 $Y=2.08
+ $X2=0 $Y2=0
cc_655 N_A_1290_365#_c_819_p N_A_1162_463#_M1031_g 0.00848302f $X=8.47 $Y=2.24
+ $X2=0 $Y2=0
cc_656 N_A_1290_365#_c_782_n N_A_1162_463#_c_1064_n 0.0655984f $X=6.705 $Y=1.99
+ $X2=0 $Y2=0
cc_657 N_A_1290_365#_c_789_n N_A_1162_463#_c_1064_n 0.00639347f $X=6.705 $Y=1.99
+ $X2=0 $Y2=0
cc_658 N_A_1290_365#_c_784_n N_A_1162_463#_c_1064_n 0.0139848f $X=6.79 $Y=1.147
+ $X2=0 $Y2=0
cc_659 N_A_1290_365#_M1000_g N_A_1162_463#_c_1095_n 0.00625211f $X=6.525
+ $Y=2.525 $X2=0 $Y2=0
cc_660 N_A_1290_365#_c_782_n N_A_1162_463#_c_1095_n 0.0105354f $X=6.705 $Y=1.99
+ $X2=0 $Y2=0
cc_661 N_A_1290_365#_c_789_n N_A_1162_463#_c_1095_n 0.00686293f $X=6.705 $Y=1.99
+ $X2=0 $Y2=0
cc_662 N_A_1290_365#_M1000_g N_A_1162_463#_c_1071_n 0.00200703f $X=6.525
+ $Y=2.525 $X2=0 $Y2=0
cc_663 N_A_1290_365#_M1036_g N_A_1162_463#_c_1071_n 6.74356e-19 $X=7.03 $Y=0.805
+ $X2=0 $Y2=0
cc_664 N_A_1290_365#_c_782_n N_A_1162_463#_c_1071_n 0.0351578f $X=6.705 $Y=1.99
+ $X2=0 $Y2=0
cc_665 N_A_1290_365#_c_789_n N_A_1162_463#_c_1071_n 0.011867f $X=6.705 $Y=1.99
+ $X2=0 $Y2=0
cc_666 N_A_1290_365#_M1036_g N_A_1162_463#_c_1065_n 0.00860506f $X=7.03 $Y=0.805
+ $X2=0 $Y2=0
cc_667 N_A_1290_365#_c_782_n N_A_1162_463#_c_1065_n 0.0191797f $X=6.705 $Y=1.99
+ $X2=0 $Y2=0
cc_668 N_A_1290_365#_c_783_n N_A_1162_463#_c_1065_n 0.0131832f $X=8.31 $Y=1.147
+ $X2=0 $Y2=0
cc_669 N_A_1290_365#_M1036_g N_A_1162_463#_c_1083_n 7.06276e-19 $X=7.03 $Y=0.805
+ $X2=0 $Y2=0
cc_670 N_A_1290_365#_M1000_g N_A_1162_463#_c_1106_n 0.0116295f $X=6.525 $Y=2.525
+ $X2=0 $Y2=0
cc_671 N_A_1290_365#_c_785_n N_A_1162_463#_c_1107_n 0.0262565f $X=8.47 $Y=2.08
+ $X2=0 $Y2=0
cc_672 N_A_1290_365#_c_783_n N_A_1162_463#_c_1066_n 0.0073032f $X=8.31 $Y=1.147
+ $X2=0 $Y2=0
cc_673 N_A_1290_365#_c_785_n N_A_1162_463#_c_1066_n 0.00848302f $X=8.47 $Y=2.08
+ $X2=0 $Y2=0
cc_674 N_A_1290_365#_c_783_n N_A_1162_463#_c_1067_n 0.0759056f $X=8.31 $Y=1.147
+ $X2=0 $Y2=0
cc_675 N_A_1290_365#_M1000_g N_A_759_119#_M1023_g 0.0421213f $X=6.525 $Y=2.525
+ $X2=0 $Y2=0
cc_676 N_A_1290_365#_M1000_g N_A_759_119#_c_1196_n 0.00991692f $X=6.525 $Y=2.525
+ $X2=0 $Y2=0
cc_677 N_A_1290_365#_c_790_n N_A_759_119#_c_1196_n 0.00678272f $X=8.415 $Y=2.27
+ $X2=0 $Y2=0
cc_678 N_A_1290_365#_c_819_p N_A_759_119#_M1010_g 0.00831176f $X=8.47 $Y=2.24
+ $X2=0 $Y2=0
cc_679 N_A_1290_365#_c_785_n N_A_759_119#_c_1184_n 0.00617069f $X=8.47 $Y=2.08
+ $X2=0 $Y2=0
cc_680 N_A_1290_365#_c_819_p N_A_1770_412#_c_1485_n 0.0285834f $X=8.47 $Y=2.24
+ $X2=0 $Y2=0
cc_681 N_A_1290_365#_c_790_n N_A_1770_412#_c_1481_n 0.0285834f $X=8.415 $Y=2.27
+ $X2=0 $Y2=0
cc_682 N_A_1290_365#_M1000_g N_VPWR_c_1705_n 0.00504141f $X=6.525 $Y=2.525 $X2=0
+ $Y2=0
cc_683 N_A_1290_365#_c_819_p N_VPWR_c_1706_n 0.0270903f $X=8.47 $Y=2.24 $X2=0
+ $Y2=0
cc_684 N_A_1290_365#_c_790_n N_VPWR_c_1720_n 0.0110482f $X=8.415 $Y=2.27 $X2=0
+ $Y2=0
cc_685 N_A_1290_365#_M1000_g N_VPWR_c_1701_n 9.39239e-19 $X=6.525 $Y=2.525 $X2=0
+ $Y2=0
cc_686 N_A_1290_365#_c_790_n N_VPWR_c_1701_n 0.00996136f $X=8.415 $Y=2.27 $X2=0
+ $Y2=0
cc_687 N_RESET_B_c_859_n N_A_1162_463#_M1005_g 0.0227619f $X=7.315 $Y=0.18 $X2=0
+ $Y2=0
cc_688 N_RESET_B_M1025_g N_A_1162_463#_M1031_g 0.00193099f $X=7.39 $Y=0.805
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_871_n N_A_1162_463#_M1031_g 0.0140916f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_873_n N_A_1162_463#_M1031_g 0.00147624f $X=7.44 $Y=2.035
+ $X2=0 $Y2=0
cc_691 N_RESET_B_c_877_n N_A_1162_463#_M1031_g 0.00817172f $X=7.39 $Y=2.03 $X2=0
+ $Y2=0
cc_692 N_RESET_B_c_869_n N_A_1162_463#_c_1069_n 0.0102825f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_869_n N_A_1162_463#_c_1064_n 0.0190173f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_694 N_RESET_B_c_869_n N_A_1162_463#_c_1095_n 0.0116621f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_695 N_RESET_B_c_865_n N_A_1162_463#_c_1071_n 0.016705f $X=7.185 $Y=2.24 $X2=0
+ $Y2=0
cc_696 N_RESET_B_M1025_g N_A_1162_463#_c_1071_n 0.00352375f $X=7.39 $Y=0.805
+ $X2=0 $Y2=0
cc_697 N_RESET_B_c_869_n N_A_1162_463#_c_1071_n 0.0228429f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_698 N_RESET_B_c_872_n N_A_1162_463#_c_1071_n 0.0047582f $X=7.585 $Y=2.035
+ $X2=0 $Y2=0
cc_699 N_RESET_B_c_873_n N_A_1162_463#_c_1071_n 0.0408999f $X=7.44 $Y=2.035
+ $X2=0 $Y2=0
cc_700 N_RESET_B_c_877_n N_A_1162_463#_c_1071_n 0.0132454f $X=7.39 $Y=2.03 $X2=0
+ $Y2=0
cc_701 N_RESET_B_c_865_n N_A_1162_463#_c_1106_n 6.05512e-19 $X=7.185 $Y=2.24
+ $X2=0 $Y2=0
cc_702 N_RESET_B_c_869_n N_A_1162_463#_c_1106_n 0.00271146f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_703 N_RESET_B_M1025_g N_A_1162_463#_c_1107_n 4.41981e-19 $X=7.39 $Y=0.805
+ $X2=0 $Y2=0
cc_704 N_RESET_B_c_871_n N_A_1162_463#_c_1107_n 0.00632872f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_705 N_RESET_B_M1025_g N_A_1162_463#_c_1066_n 0.00914674f $X=7.39 $Y=0.805
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_871_n N_A_1162_463#_c_1066_n 0.00595038f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_707 N_RESET_B_M1025_g N_A_1162_463#_c_1067_n 0.013433f $X=7.39 $Y=0.805 $X2=0
+ $Y2=0
cc_708 N_RESET_B_c_869_n N_A_1162_463#_c_1067_n 0.00665416f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_709 N_RESET_B_c_871_n N_A_1162_463#_c_1067_n 0.0114411f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_710 N_RESET_B_c_872_n N_A_1162_463#_c_1067_n 0.00190431f $X=7.585 $Y=2.035
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_873_n N_A_1162_463#_c_1067_n 0.0202286f $X=7.44 $Y=2.035
+ $X2=0 $Y2=0
cc_712 N_RESET_B_c_877_n N_A_1162_463#_c_1067_n 0.010187f $X=7.39 $Y=2.03 $X2=0
+ $Y2=0
cc_713 N_RESET_B_c_869_n N_A_759_119#_M1042_s 7.58599e-19 $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_869_n N_A_759_119#_M1017_g 0.00426681f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_RESET_B_c_859_n N_A_759_119#_c_1177_n 0.0104164f $X=7.315 $Y=0.18 $X2=0
+ $Y2=0
cc_716 N_RESET_B_c_869_n N_A_759_119#_c_1178_n 0.00218246f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_859_n N_A_759_119#_c_1179_n 0.010259f $X=7.315 $Y=0.18 $X2=0
+ $Y2=0
cc_718 N_RESET_B_c_869_n N_A_759_119#_M1023_g 0.00238159f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_859_n N_A_759_119#_c_1182_n 0.00880557f $X=7.315 $Y=0.18
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_865_n N_A_759_119#_c_1196_n 0.00991634f $X=7.185 $Y=2.24
+ $X2=0 $Y2=0
cc_721 N_RESET_B_c_871_n N_A_759_119#_M1010_g 0.00914494f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_722 N_RESET_B_c_859_n N_A_759_119#_c_1186_n 0.00123232f $X=7.315 $Y=0.18
+ $X2=0 $Y2=0
cc_723 N_RESET_B_c_869_n N_A_759_119#_c_1209_n 0.0200121f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_724 N_RESET_B_c_870_n N_A_759_119#_c_1188_n 2.2421e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_725 N_RESET_B_c_859_n N_A_759_119#_c_1189_n 0.00451754f $X=7.315 $Y=0.18
+ $X2=0 $Y2=0
cc_726 N_RESET_B_M1002_g N_A_759_119#_c_1219_n 0.00255063f $X=3.16 $Y=2.765
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_869_n N_A_759_119#_c_1219_n 0.0117881f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_728 N_RESET_B_c_870_n N_A_759_119#_c_1219_n 0.00243944f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_875_n N_A_759_119#_c_1219_n 8.30166e-19 $X=3.49 $Y=2.035
+ $X2=0 $Y2=0
cc_730 N_RESET_B_c_876_n N_A_759_119#_c_1219_n 0.0193265f $X=3.49 $Y=2.035 $X2=0
+ $Y2=0
cc_731 N_RESET_B_c_869_n N_A_759_119#_c_1190_n 0.00671515f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_732 N_RESET_B_M1012_g N_A_1923_174#_M1001_g 0.0148623f $X=10.515 $Y=2.69
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_871_n N_A_1923_174#_M1001_g 0.00224629f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_734 RESET_B N_A_1923_174#_M1001_g 2.94452e-19 $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_735 N_RESET_B_c_878_n N_A_1923_174#_M1001_g 0.0205471f $X=10.515 $Y=2.155
+ $X2=0 $Y2=0
cc_736 N_RESET_B_c_879_n N_A_1923_174#_M1001_g 0.00183701f $X=10.29 $Y=2.035
+ $X2=0 $Y2=0
cc_737 N_RESET_B_M1016_g N_A_1923_174#_c_1361_n 0.0671928f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_738 N_RESET_B_M1016_g N_A_1923_174#_c_1362_n 0.0042641f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_739 N_RESET_B_M1016_g N_A_1923_174#_c_1363_n 0.0139503f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_740 N_RESET_B_M1016_g N_A_1923_174#_c_1364_n 0.00187525f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_741 N_RESET_B_M1012_g N_A_1923_174#_c_1371_n 3.10874e-19 $X=10.515 $Y=2.69
+ $X2=0 $Y2=0
cc_742 RESET_B N_A_1923_174#_c_1372_n 2.56255e-19 $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_743 N_RESET_B_c_878_n N_A_1923_174#_c_1372_n 0.00557492f $X=10.515 $Y=2.155
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_879_n N_A_1923_174#_c_1372_n 0.0144665f $X=10.29 $Y=2.035
+ $X2=0 $Y2=0
cc_745 RESET_B N_A_1923_174#_c_1373_n 0.00113689f $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_746 N_RESET_B_c_878_n N_A_1923_174#_c_1373_n 0.00100236f $X=10.515 $Y=2.155
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_879_n N_A_1923_174#_c_1373_n 0.013066f $X=10.29 $Y=2.035
+ $X2=0 $Y2=0
cc_748 N_RESET_B_M1016_g N_A_1923_174#_c_1368_n 0.0144142f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_749 N_RESET_B_M1016_g N_A_1770_412#_M1020_g 0.0984829f $X=10.26 $Y=0.55 $X2=0
+ $Y2=0
cc_750 N_RESET_B_M1016_g N_A_1770_412#_M1045_g 0.00520259f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_751 RESET_B N_A_1770_412#_M1045_g 2.79328e-19 $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_752 N_RESET_B_c_878_n N_A_1770_412#_M1045_g 0.0272761f $X=10.515 $Y=2.155
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_879_n N_A_1770_412#_M1045_g 3.86278e-19 $X=10.29 $Y=2.035
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_871_n N_A_1770_412#_c_1485_n 0.0177681f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_755 N_RESET_B_M1012_g N_A_1770_412#_c_1490_n 2.9297e-19 $X=10.515 $Y=2.69
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_871_n N_A_1770_412#_c_1490_n 0.0106114f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_871_n N_A_1770_412#_c_1469_n 0.00799873f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_871_n N_A_1770_412#_c_1470_n 7.86049e-19 $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_759 N_RESET_B_M1016_g N_A_1770_412#_c_1479_n 0.0011681f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_760 N_RESET_B_M1012_g N_A_1770_412#_c_1479_n 8.81388e-19 $X=10.515 $Y=2.69
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_871_n N_A_1770_412#_c_1479_n 0.0235207f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_762 RESET_B N_A_1770_412#_c_1479_n 0.00132301f $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_763 N_RESET_B_c_878_n N_A_1770_412#_c_1479_n 5.35563e-19 $X=10.515 $Y=2.155
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_879_n N_A_1770_412#_c_1479_n 0.0235661f $X=10.29 $Y=2.035
+ $X2=0 $Y2=0
cc_765 N_RESET_B_M1016_g N_A_1770_412#_c_1471_n 0.0148403f $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_871_n N_A_1770_412#_c_1471_n 0.00807134f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_767 RESET_B N_A_1770_412#_c_1471_n 0.00757528f $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_768 N_RESET_B_c_878_n N_A_1770_412#_c_1471_n 0.0031813f $X=10.515 $Y=2.155
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_879_n N_A_1770_412#_c_1471_n 0.0251085f $X=10.29 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_871_n N_A_1770_412#_c_1481_n 0.00123766f $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_771 N_RESET_B_M1016_g N_A_1770_412#_c_1473_n 4.46351e-19 $X=10.26 $Y=0.55
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_871_n N_A_1770_412#_c_1473_n 8.07599e-19 $X=10.145 $Y=2.035
+ $X2=0 $Y2=0
cc_773 N_RESET_B_c_878_n N_A_1770_412#_c_1474_n 0.00343497f $X=10.515 $Y=2.155
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_869_n N_VPWR_M1042_d 0.00285593f $X=7.295 $Y=2.035 $X2=0
+ $Y2=0
cc_775 N_RESET_B_c_871_n N_VPWR_M1031_s 0.00666183f $X=10.145 $Y=2.035 $X2=0
+ $Y2=0
cc_776 N_RESET_B_M1002_g N_VPWR_c_1703_n 0.00523771f $X=3.16 $Y=2.765 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_865_n N_VPWR_c_1705_n 0.00504141f $X=7.185 $Y=2.24 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_869_n N_VPWR_c_1705_n 5.7432e-19 $X=7.295 $Y=2.035 $X2=0
+ $Y2=0
cc_779 N_RESET_B_c_865_n N_VPWR_c_1706_n 0.00538542f $X=7.185 $Y=2.24 $X2=0
+ $Y2=0
cc_780 N_RESET_B_c_871_n N_VPWR_c_1706_n 0.016919f $X=10.145 $Y=2.035 $X2=0
+ $Y2=0
cc_781 N_RESET_B_c_872_n N_VPWR_c_1706_n 3.31316e-19 $X=7.585 $Y=2.035 $X2=0
+ $Y2=0
cc_782 N_RESET_B_c_873_n N_VPWR_c_1706_n 0.00484065f $X=7.44 $Y=2.035 $X2=0
+ $Y2=0
cc_783 N_RESET_B_c_877_n N_VPWR_c_1706_n 0.00205156f $X=7.39 $Y=2.03 $X2=0 $Y2=0
cc_784 N_RESET_B_M1002_g N_VPWR_c_1714_n 0.00411906f $X=3.16 $Y=2.765 $X2=0
+ $Y2=0
cc_785 N_RESET_B_M1012_g N_VPWR_c_1721_n 0.00479724f $X=10.515 $Y=2.69 $X2=0
+ $Y2=0
cc_786 N_RESET_B_M1012_g N_VPWR_c_1727_n 0.0149179f $X=10.515 $Y=2.69 $X2=0
+ $Y2=0
cc_787 N_RESET_B_c_871_n N_VPWR_c_1727_n 9.75304e-19 $X=10.145 $Y=2.035 $X2=0
+ $Y2=0
cc_788 RESET_B N_VPWR_c_1727_n 0.00178525f $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_789 N_RESET_B_c_878_n N_VPWR_c_1727_n 0.00649976f $X=10.515 $Y=2.155 $X2=0
+ $Y2=0
cc_790 N_RESET_B_c_879_n N_VPWR_c_1727_n 0.0184765f $X=10.29 $Y=2.035 $X2=0
+ $Y2=0
cc_791 N_RESET_B_M1002_g N_VPWR_c_1701_n 0.00740422f $X=3.16 $Y=2.765 $X2=0
+ $Y2=0
cc_792 N_RESET_B_c_865_n N_VPWR_c_1701_n 9.39239e-19 $X=7.185 $Y=2.24 $X2=0
+ $Y2=0
cc_793 N_RESET_B_M1012_g N_VPWR_c_1701_n 0.00474109f $X=10.515 $Y=2.69 $X2=0
+ $Y2=0
cc_794 N_RESET_B_M1015_g N_A_359_489#_c_1902_n 0.00262237f $X=3.23 $Y=0.615
+ $X2=0 $Y2=0
cc_795 N_RESET_B_M1002_g N_A_359_489#_c_1903_n 0.0123038f $X=3.16 $Y=2.765 $X2=0
+ $Y2=0
cc_796 N_RESET_B_M1015_g N_A_359_489#_c_1903_n 0.012728f $X=3.23 $Y=0.615 $X2=0
+ $Y2=0
cc_797 N_RESET_B_c_870_n N_A_359_489#_c_1903_n 0.00112914f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_875_n N_A_359_489#_c_1903_n 0.0108103f $X=3.49 $Y=2.035 $X2=0
+ $Y2=0
cc_799 N_RESET_B_c_876_n N_A_359_489#_c_1903_n 0.0181363f $X=3.49 $Y=2.035 $X2=0
+ $Y2=0
cc_800 N_RESET_B_c_869_n N_A_359_489#_c_1907_n 0.0297622f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_801 N_RESET_B_c_870_n N_A_359_489#_c_1907_n 0.00302339f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_802 N_RESET_B_c_875_n N_A_359_489#_c_1907_n 0.00237779f $X=3.49 $Y=2.035
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_876_n N_A_359_489#_c_1907_n 0.00681109f $X=3.49 $Y=2.035
+ $X2=0 $Y2=0
cc_804 N_RESET_B_M1002_g N_A_359_489#_c_1908_n 0.0145424f $X=3.16 $Y=2.765 $X2=0
+ $Y2=0
cc_805 N_RESET_B_c_870_n N_A_359_489#_c_1908_n 6.30115e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_806 N_RESET_B_c_875_n N_A_359_489#_c_1908_n 0.00718486f $X=3.49 $Y=2.035
+ $X2=0 $Y2=0
cc_807 N_RESET_B_c_876_n N_A_359_489#_c_1908_n 0.0109949f $X=3.49 $Y=2.035 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_869_n N_A_359_489#_c_1909_n 0.0301997f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_809 N_RESET_B_c_869_n N_A_359_489#_c_1910_n 0.019911f $X=7.295 $Y=2.035 $X2=0
+ $Y2=0
cc_810 N_RESET_B_M1002_g N_A_359_489#_c_1913_n 0.00644891f $X=3.16 $Y=2.765
+ $X2=0 $Y2=0
cc_811 N_RESET_B_c_869_n N_A_359_489#_c_1914_n 0.00100847f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_812 N_RESET_B_M1015_g N_VGND_c_2084_n 0.00163721f $X=3.23 $Y=0.615 $X2=0
+ $Y2=0
cc_813 N_RESET_B_c_859_n N_VGND_c_2084_n 0.0195255f $X=7.315 $Y=0.18 $X2=0 $Y2=0
cc_814 N_RESET_B_c_859_n N_VGND_c_2085_n 0.0239437f $X=7.315 $Y=0.18 $X2=0 $Y2=0
cc_815 N_RESET_B_c_859_n N_VGND_c_2086_n 0.0162969f $X=7.315 $Y=0.18 $X2=0 $Y2=0
cc_816 N_RESET_B_c_859_n N_VGND_c_2087_n 0.00832272f $X=7.315 $Y=0.18 $X2=0
+ $Y2=0
cc_817 N_RESET_B_M1016_g N_VGND_c_2088_n 0.00998474f $X=10.26 $Y=0.55 $X2=0
+ $Y2=0
cc_818 N_RESET_B_c_860_n N_VGND_c_2094_n 0.00720997f $X=3.305 $Y=0.18 $X2=0
+ $Y2=0
cc_819 N_RESET_B_c_859_n N_VGND_c_2096_n 0.0200455f $X=7.315 $Y=0.18 $X2=0 $Y2=0
cc_820 N_RESET_B_c_859_n N_VGND_c_2098_n 0.0200856f $X=7.315 $Y=0.18 $X2=0 $Y2=0
cc_821 N_RESET_B_c_859_n N_VGND_c_2103_n 0.0459765f $X=7.315 $Y=0.18 $X2=0 $Y2=0
cc_822 N_RESET_B_M1016_g N_VGND_c_2104_n 0.0040395f $X=10.26 $Y=0.55 $X2=0 $Y2=0
cc_823 N_RESET_B_c_859_n N_VGND_c_2113_n 0.098719f $X=7.315 $Y=0.18 $X2=0 $Y2=0
cc_824 N_RESET_B_c_860_n N_VGND_c_2113_n 0.0105672f $X=3.305 $Y=0.18 $X2=0 $Y2=0
cc_825 N_RESET_B_M1016_g N_VGND_c_2113_n 0.0040417f $X=10.26 $Y=0.55 $X2=0 $Y2=0
cc_826 N_RESET_B_M1015_g N_noxref_25_c_2247_n 0.00725814f $X=3.23 $Y=0.615 $X2=0
+ $Y2=0
cc_827 N_A_1162_463#_c_1069_n N_A_759_119#_c_1193_n 0.00328899f $X=6.28 $Y=2.492
+ $X2=0 $Y2=0
cc_828 N_A_1162_463#_c_1064_n N_A_759_119#_c_1180_n 0.00389851f $X=6.365 $Y=2.29
+ $X2=0 $Y2=0
cc_829 N_A_1162_463#_c_1069_n N_A_759_119#_M1023_g 0.0142952f $X=6.28 $Y=2.492
+ $X2=0 $Y2=0
cc_830 N_A_1162_463#_c_1064_n N_A_759_119#_M1023_g 0.00128094f $X=6.365 $Y=2.29
+ $X2=0 $Y2=0
cc_831 N_A_1162_463#_c_1064_n N_A_759_119#_c_1182_n 0.00320468f $X=6.365 $Y=2.29
+ $X2=0 $Y2=0
cc_832 N_A_1162_463#_c_1083_n N_A_759_119#_c_1182_n 0.00324584f $X=6.455
+ $Y=0.775 $X2=0 $Y2=0
cc_833 N_A_1162_463#_M1031_g N_A_759_119#_c_1196_n 0.0104164f $X=8.2 $Y=2.315
+ $X2=0 $Y2=0
cc_834 N_A_1162_463#_c_1095_n N_A_759_119#_c_1196_n 0.00250273f $X=6.96 $Y=2.42
+ $X2=0 $Y2=0
cc_835 N_A_1162_463#_c_1071_n N_A_759_119#_c_1196_n 0.00757414f $X=7.045
+ $Y=2.335 $X2=0 $Y2=0
cc_836 N_A_1162_463#_c_1106_n N_A_759_119#_c_1196_n 0.00217491f $X=6.28 $Y=2.29
+ $X2=0 $Y2=0
cc_837 N_A_1162_463#_M1031_g N_A_759_119#_M1010_g 0.0107715f $X=8.2 $Y=2.315
+ $X2=0 $Y2=0
cc_838 N_A_1162_463#_c_1066_n N_A_759_119#_c_1184_n 0.0107715f $X=8.05 $Y=1.57
+ $X2=0 $Y2=0
cc_839 N_A_1162_463#_c_1095_n N_VPWR_M1000_d 0.00602989f $X=6.96 $Y=2.42 $X2=0
+ $Y2=0
cc_840 N_A_1162_463#_c_1071_n N_VPWR_M1000_d 0.00116866f $X=7.045 $Y=2.335 $X2=0
+ $Y2=0
cc_841 N_A_1162_463#_c_1095_n N_VPWR_c_1705_n 0.0206919f $X=6.96 $Y=2.42 $X2=0
+ $Y2=0
cc_842 N_A_1162_463#_c_1071_n N_VPWR_c_1705_n 0.00657508f $X=7.045 $Y=2.335
+ $X2=0 $Y2=0
cc_843 N_A_1162_463#_c_1106_n N_VPWR_c_1705_n 0.00164807f $X=6.28 $Y=2.29 $X2=0
+ $Y2=0
cc_844 N_A_1162_463#_M1031_g N_VPWR_c_1706_n 0.00578392f $X=8.2 $Y=2.315 $X2=0
+ $Y2=0
cc_845 N_A_1162_463#_c_1071_n N_VPWR_c_1706_n 0.0310743f $X=7.045 $Y=2.335 $X2=0
+ $Y2=0
cc_846 N_A_1162_463#_c_1107_n N_VPWR_c_1706_n 0.0016941f $X=8.05 $Y=1.57 $X2=0
+ $Y2=0
cc_847 N_A_1162_463#_c_1066_n N_VPWR_c_1706_n 0.00271454f $X=8.05 $Y=1.57 $X2=0
+ $Y2=0
cc_848 N_A_1162_463#_c_1067_n N_VPWR_c_1706_n 0.0043187f $X=7.965 $Y=1.57 $X2=0
+ $Y2=0
cc_849 N_A_1162_463#_c_1069_n N_VPWR_c_1716_n 0.00741458f $X=6.28 $Y=2.492 $X2=0
+ $Y2=0
cc_850 N_A_1162_463#_c_1106_n N_VPWR_c_1716_n 0.00377769f $X=6.28 $Y=2.29 $X2=0
+ $Y2=0
cc_851 N_A_1162_463#_c_1071_n N_VPWR_c_1719_n 0.00635448f $X=7.045 $Y=2.335
+ $X2=0 $Y2=0
cc_852 N_A_1162_463#_M1031_g N_VPWR_c_1701_n 9.39239e-19 $X=8.2 $Y=2.315 $X2=0
+ $Y2=0
cc_853 N_A_1162_463#_c_1069_n N_VPWR_c_1701_n 0.0121941f $X=6.28 $Y=2.492 $X2=0
+ $Y2=0
cc_854 N_A_1162_463#_c_1095_n N_VPWR_c_1701_n 0.00593413f $X=6.96 $Y=2.42 $X2=0
+ $Y2=0
cc_855 N_A_1162_463#_c_1071_n N_VPWR_c_1701_n 0.0153f $X=7.045 $Y=2.335 $X2=0
+ $Y2=0
cc_856 N_A_1162_463#_c_1106_n N_VPWR_c_1701_n 0.00619882f $X=6.28 $Y=2.29 $X2=0
+ $Y2=0
cc_857 N_A_1162_463#_c_1069_n N_A_359_489#_c_1909_n 0.0241635f $X=6.28 $Y=2.492
+ $X2=0 $Y2=0
cc_858 N_A_1162_463#_c_1064_n N_A_359_489#_c_1909_n 0.0127113f $X=6.365 $Y=2.29
+ $X2=0 $Y2=0
cc_859 N_A_1162_463#_c_1064_n N_A_359_489#_c_1904_n 0.0719922f $X=6.365 $Y=2.29
+ $X2=0 $Y2=0
cc_860 N_A_1162_463#_c_1069_n N_A_359_489#_c_1915_n 0.0162354f $X=6.28 $Y=2.492
+ $X2=0 $Y2=0
cc_861 N_A_1162_463#_c_1064_n N_A_359_489#_c_1915_n 0.00500153f $X=6.365 $Y=2.29
+ $X2=0 $Y2=0
cc_862 N_A_1162_463#_c_1106_n A_1248_463# 0.00151427f $X=6.28 $Y=2.29 $X2=-0.19
+ $Y2=-0.245
cc_863 N_A_1162_463#_M1005_g N_VGND_c_2087_n 0.00952974f $X=8.1 $Y=0.66 $X2=0
+ $Y2=0
cc_864 N_A_1162_463#_M1005_g N_VGND_c_2100_n 0.00355322f $X=8.1 $Y=0.66 $X2=0
+ $Y2=0
cc_865 N_A_1162_463#_M1005_g N_VGND_c_2113_n 0.00519272f $X=8.1 $Y=0.66 $X2=0
+ $Y2=0
cc_866 N_A_759_119#_M1040_g N_A_1923_174#_M1001_g 0.014558f $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_867 N_A_759_119#_M1040_g N_A_1923_174#_c_1361_n 0.0201128f $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_868 N_A_759_119#_M1040_g N_A_1923_174#_c_1366_n 3.98181e-19 $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_869 N_A_759_119#_M1040_g N_A_1923_174#_c_1368_n 0.0199546f $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_870 N_A_759_119#_M1010_g N_A_1770_412#_c_1485_n 0.00486021f $X=8.775 $Y=2.48
+ $X2=0 $Y2=0
cc_871 N_A_759_119#_c_1183_n N_A_1770_412#_c_1485_n 0.00123617f $X=9.245
+ $Y=1.705 $X2=0 $Y2=0
cc_872 N_A_759_119#_M1040_g N_A_1770_412#_c_1468_n 0.016651f $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_873 N_A_759_119#_M1040_g N_A_1770_412#_c_1470_n 0.0087442f $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_874 N_A_759_119#_M1010_g N_A_1770_412#_c_1481_n 0.00569159f $X=8.775 $Y=2.48
+ $X2=0 $Y2=0
cc_875 N_A_759_119#_M1040_g N_A_1770_412#_c_1472_n 0.0102305f $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_876 N_A_759_119#_c_1183_n N_A_1770_412#_c_1473_n 2.1968e-19 $X=9.245 $Y=1.705
+ $X2=0 $Y2=0
cc_877 N_A_759_119#_M1040_g N_A_1770_412#_c_1473_n 0.00398124f $X=9.32 $Y=0.55
+ $X2=0 $Y2=0
cc_878 N_A_759_119#_c_1209_n N_VPWR_M1042_d 0.00376426f $X=4.345 $Y=2.015 $X2=0
+ $Y2=0
cc_879 N_A_759_119#_c_1188_n N_VPWR_M1042_d 0.00128318f $X=4.43 $Y=1.93 $X2=0
+ $Y2=0
cc_880 N_A_759_119#_M1017_g N_VPWR_c_1704_n 0.0102678f $X=4.595 $Y=2.465 $X2=0
+ $Y2=0
cc_881 N_A_759_119#_c_1178_n N_VPWR_c_1704_n 0.00237213f $X=5.085 $Y=3.075 $X2=0
+ $Y2=0
cc_882 N_A_759_119#_M1023_g N_VPWR_c_1705_n 0.00604888f $X=6.165 $Y=2.525 $X2=0
+ $Y2=0
cc_883 N_A_759_119#_c_1196_n N_VPWR_c_1705_n 0.0253068f $X=8.7 $Y=3.15 $X2=0
+ $Y2=0
cc_884 N_A_759_119#_c_1196_n N_VPWR_c_1706_n 0.0216291f $X=8.7 $Y=3.15 $X2=0
+ $Y2=0
cc_885 N_A_759_119#_M1010_g N_VPWR_c_1706_n 0.00357722f $X=8.775 $Y=2.48 $X2=0
+ $Y2=0
cc_886 N_A_759_119#_M1017_g N_VPWR_c_1716_n 0.00358332f $X=4.595 $Y=2.465 $X2=0
+ $Y2=0
cc_887 N_A_759_119#_c_1194_n N_VPWR_c_1716_n 0.0472789f $X=5.16 $Y=3.15 $X2=0
+ $Y2=0
cc_888 N_A_759_119#_c_1196_n N_VPWR_c_1719_n 0.0226041f $X=8.7 $Y=3.15 $X2=0
+ $Y2=0
cc_889 N_A_759_119#_c_1196_n N_VPWR_c_1720_n 0.0255173f $X=8.7 $Y=3.15 $X2=0
+ $Y2=0
cc_890 N_A_759_119#_M1042_s N_VPWR_c_1701_n 0.00326452f $X=3.825 $Y=1.835 $X2=0
+ $Y2=0
cc_891 N_A_759_119#_M1017_g N_VPWR_c_1701_n 0.00443322f $X=4.595 $Y=2.465 $X2=0
+ $Y2=0
cc_892 N_A_759_119#_c_1193_n N_VPWR_c_1701_n 0.0272026f $X=6.09 $Y=3.15 $X2=0
+ $Y2=0
cc_893 N_A_759_119#_c_1194_n N_VPWR_c_1701_n 0.00542487f $X=5.16 $Y=3.15 $X2=0
+ $Y2=0
cc_894 N_A_759_119#_c_1196_n N_VPWR_c_1701_n 0.07319f $X=8.7 $Y=3.15 $X2=0 $Y2=0
cc_895 N_A_759_119#_c_1200_n N_VPWR_c_1701_n 0.00431118f $X=6.165 $Y=3.15 $X2=0
+ $Y2=0
cc_896 N_A_759_119#_c_1189_n N_A_359_489#_c_1903_n 0.00143236f $X=3.935 $Y=0.82
+ $X2=0 $Y2=0
cc_897 N_A_759_119#_M1042_s N_A_359_489#_c_1907_n 0.00694903f $X=3.825 $Y=1.835
+ $X2=0 $Y2=0
cc_898 N_A_759_119#_M1017_g N_A_359_489#_c_1907_n 0.0128823f $X=4.595 $Y=2.465
+ $X2=0 $Y2=0
cc_899 N_A_759_119#_c_1178_n N_A_359_489#_c_1907_n 0.0129087f $X=5.085 $Y=3.075
+ $X2=0 $Y2=0
cc_900 N_A_759_119#_c_1193_n N_A_359_489#_c_1907_n 0.00179868f $X=6.09 $Y=3.15
+ $X2=0 $Y2=0
cc_901 N_A_759_119#_c_1209_n N_A_359_489#_c_1907_n 0.00819849f $X=4.345 $Y=2.015
+ $X2=0 $Y2=0
cc_902 N_A_759_119#_c_1219_n N_A_359_489#_c_1907_n 0.0139554f $X=3.99 $Y=2.015
+ $X2=0 $Y2=0
cc_903 N_A_759_119#_M1023_g N_A_359_489#_c_1909_n 2.89603e-19 $X=6.165 $Y=2.525
+ $X2=0 $Y2=0
cc_904 N_A_759_119#_c_1178_n N_A_359_489#_c_1910_n 0.0011732f $X=5.085 $Y=3.075
+ $X2=0 $Y2=0
cc_905 N_A_759_119#_c_1180_n N_A_359_489#_c_1904_n 0.0108241f $X=6.165 $Y=1.165
+ $X2=0 $Y2=0
cc_906 N_A_759_119#_c_1182_n N_A_359_489#_c_1904_n 0.00171886f $X=6.24 $Y=1.09
+ $X2=0 $Y2=0
cc_907 N_A_759_119#_c_1178_n N_A_359_489#_c_1914_n 0.00411454f $X=5.085 $Y=3.075
+ $X2=0 $Y2=0
cc_908 N_A_759_119#_c_1193_n N_A_359_489#_c_1914_n 0.00487376f $X=6.09 $Y=3.15
+ $X2=0 $Y2=0
cc_909 N_A_759_119#_c_1178_n N_A_359_489#_c_1915_n 0.00184742f $X=5.085 $Y=3.075
+ $X2=0 $Y2=0
cc_910 N_A_759_119#_c_1186_n N_VGND_M1022_s 0.00472939f $X=4.345 $Y=0.95 $X2=0
+ $Y2=0
cc_911 N_A_759_119#_c_1177_n N_VGND_c_2085_n 0.0027164f $X=4.7 $Y=1.09 $X2=0
+ $Y2=0
cc_912 N_A_759_119#_c_1181_n N_VGND_c_2085_n 0.00128968f $X=5.205 $Y=1.165 $X2=0
+ $Y2=0
cc_913 N_A_759_119#_c_1186_n N_VGND_c_2085_n 0.0194919f $X=4.345 $Y=0.95 $X2=0
+ $Y2=0
cc_914 N_A_759_119#_c_1190_n N_VGND_c_2085_n 0.00198709f $X=4.685 $Y=1.445 $X2=0
+ $Y2=0
cc_915 N_A_759_119#_c_1179_n N_VGND_c_2086_n 0.00362786f $X=5.13 $Y=1.09 $X2=0
+ $Y2=0
cc_916 N_A_759_119#_c_1180_n N_VGND_c_2086_n 0.0010291f $X=6.165 $Y=1.165 $X2=0
+ $Y2=0
cc_917 N_A_759_119#_M1040_g N_VGND_c_2088_n 7.08958e-19 $X=9.32 $Y=0.55 $X2=0
+ $Y2=0
cc_918 N_A_759_119#_c_1189_n N_VGND_c_2096_n 0.00439599f $X=3.935 $Y=0.82 $X2=0
+ $Y2=0
cc_919 N_A_759_119#_M1040_g N_VGND_c_2100_n 0.00294187f $X=9.32 $Y=0.55 $X2=0
+ $Y2=0
cc_920 N_A_759_119#_c_1177_n N_VGND_c_2113_n 9.39239e-19 $X=4.7 $Y=1.09 $X2=0
+ $Y2=0
cc_921 N_A_759_119#_c_1179_n N_VGND_c_2113_n 9.39239e-19 $X=5.13 $Y=1.09 $X2=0
+ $Y2=0
cc_922 N_A_759_119#_M1040_g N_VGND_c_2113_n 0.00418184f $X=9.32 $Y=0.55 $X2=0
+ $Y2=0
cc_923 N_A_759_119#_c_1186_n N_VGND_c_2113_n 0.00638806f $X=4.345 $Y=0.95 $X2=0
+ $Y2=0
cc_924 N_A_759_119#_c_1189_n N_VGND_c_2113_n 0.00689175f $X=3.935 $Y=0.82 $X2=0
+ $Y2=0
cc_925 N_A_1923_174#_c_1362_n N_A_1770_412#_M1020_g 0.0131965f $X=10.67 $Y=1.06
+ $X2=0 $Y2=0
cc_926 N_A_1923_174#_c_1364_n N_A_1770_412#_M1020_g 0.0117304f $X=10.835 $Y=0.55
+ $X2=0 $Y2=0
cc_927 N_A_1923_174#_c_1365_n N_A_1770_412#_M1020_g 0.00329477f $X=11.15 $Y=1.94
+ $X2=0 $Y2=0
cc_928 N_A_1923_174#_c_1367_n N_A_1770_412#_M1020_g 0.00988847f $X=10.835
+ $Y=1.06 $X2=0 $Y2=0
cc_929 N_A_1923_174#_c_1371_n N_A_1770_412#_M1045_g 0.00534418f $X=10.73 $Y=2.69
+ $X2=0 $Y2=0
cc_930 N_A_1923_174#_c_1372_n N_A_1770_412#_M1045_g 0.00888572f $X=10.76 $Y=2.47
+ $X2=0 $Y2=0
cc_931 N_A_1923_174#_c_1373_n N_A_1770_412#_M1045_g 0.0179254f $X=11.15 $Y=2.025
+ $X2=0 $Y2=0
cc_932 N_A_1923_174#_c_1365_n N_A_1770_412#_c_1456_n 0.0153803f $X=11.15 $Y=1.94
+ $X2=0 $Y2=0
cc_933 N_A_1923_174#_c_1373_n N_A_1770_412#_c_1456_n 3.41143e-19 $X=11.15
+ $Y=2.025 $X2=0 $Y2=0
cc_934 N_A_1923_174#_c_1365_n N_A_1770_412#_M1007_g 0.00356751f $X=11.15 $Y=1.94
+ $X2=0 $Y2=0
cc_935 N_A_1923_174#_c_1372_n N_A_1770_412#_M1007_g 7.35209e-19 $X=10.76 $Y=2.47
+ $X2=0 $Y2=0
cc_936 N_A_1923_174#_c_1373_n N_A_1770_412#_M1007_g 0.00169057f $X=11.15
+ $Y=2.025 $X2=0 $Y2=0
cc_937 N_A_1923_174#_c_1365_n N_A_1770_412#_M1003_g 0.0023134f $X=11.15 $Y=1.94
+ $X2=0 $Y2=0
cc_938 N_A_1923_174#_c_1367_n N_A_1770_412#_M1003_g 0.00670329f $X=10.835
+ $Y=1.06 $X2=0 $Y2=0
cc_939 N_A_1923_174#_M1001_g N_A_1770_412#_c_1490_n 0.00791286f $X=9.89 $Y=2.69
+ $X2=0 $Y2=0
cc_940 N_A_1923_174#_M1001_g N_A_1770_412#_c_1468_n 0.00285248f $X=9.89 $Y=2.69
+ $X2=0 $Y2=0
cc_941 N_A_1923_174#_c_1361_n N_A_1770_412#_c_1468_n 0.00120807f $X=9.78
+ $Y=1.035 $X2=0 $Y2=0
cc_942 N_A_1923_174#_c_1366_n N_A_1770_412#_c_1468_n 0.0266109f $X=10.125
+ $Y=1.06 $X2=0 $Y2=0
cc_943 N_A_1923_174#_c_1368_n N_A_1770_412#_c_1468_n 0.00225767f $X=9.79 $Y=0.87
+ $X2=0 $Y2=0
cc_944 N_A_1923_174#_c_1361_n N_A_1770_412#_c_1469_n 0.0034403f $X=9.78 $Y=1.035
+ $X2=0 $Y2=0
cc_945 N_A_1923_174#_c_1366_n N_A_1770_412#_c_1469_n 0.0112357f $X=10.125
+ $Y=1.06 $X2=0 $Y2=0
cc_946 N_A_1923_174#_M1001_g N_A_1770_412#_c_1479_n 0.0200045f $X=9.89 $Y=2.69
+ $X2=0 $Y2=0
cc_947 N_A_1923_174#_M1001_g N_A_1770_412#_c_1471_n 0.00366258f $X=9.89 $Y=2.69
+ $X2=0 $Y2=0
cc_948 N_A_1923_174#_c_1363_n N_A_1770_412#_c_1471_n 0.0436829f $X=10.325
+ $Y=1.06 $X2=0 $Y2=0
cc_949 N_A_1923_174#_c_1365_n N_A_1770_412#_c_1471_n 0.0237099f $X=11.15 $Y=1.94
+ $X2=0 $Y2=0
cc_950 N_A_1923_174#_c_1366_n N_A_1770_412#_c_1471_n 0.0109833f $X=10.125
+ $Y=1.06 $X2=0 $Y2=0
cc_951 N_A_1923_174#_c_1367_n N_A_1770_412#_c_1471_n 0.0171769f $X=10.835
+ $Y=1.06 $X2=0 $Y2=0
cc_952 N_A_1923_174#_c_1373_n N_A_1770_412#_c_1471_n 0.0143784f $X=11.15
+ $Y=2.025 $X2=0 $Y2=0
cc_953 N_A_1923_174#_c_1368_n N_A_1770_412#_c_1472_n 0.00166262f $X=9.79 $Y=0.87
+ $X2=0 $Y2=0
cc_954 N_A_1923_174#_M1001_g N_A_1770_412#_c_1473_n 0.0130659f $X=9.89 $Y=2.69
+ $X2=0 $Y2=0
cc_955 N_A_1923_174#_c_1361_n N_A_1770_412#_c_1473_n 0.00137822f $X=9.78
+ $Y=1.035 $X2=0 $Y2=0
cc_956 N_A_1923_174#_c_1366_n N_A_1770_412#_c_1473_n 0.0153267f $X=10.125
+ $Y=1.06 $X2=0 $Y2=0
cc_957 N_A_1923_174#_c_1365_n N_A_1770_412#_c_1474_n 0.00745248f $X=11.15
+ $Y=1.94 $X2=0 $Y2=0
cc_958 N_A_1923_174#_c_1371_n N_A_1770_412#_c_1474_n 0.00129642f $X=10.73
+ $Y=2.69 $X2=0 $Y2=0
cc_959 N_A_1923_174#_c_1367_n N_A_1770_412#_c_1474_n 0.0115749f $X=10.835
+ $Y=1.06 $X2=0 $Y2=0
cc_960 N_A_1923_174#_c_1373_n N_A_1770_412#_c_1474_n 0.00496318f $X=11.15
+ $Y=2.025 $X2=0 $Y2=0
cc_961 N_A_1923_174#_c_1365_n N_VPWR_M1045_d 0.00169848f $X=11.15 $Y=1.94 $X2=0
+ $Y2=0
cc_962 N_A_1923_174#_c_1373_n N_VPWR_M1045_d 0.00335436f $X=11.15 $Y=2.025 $X2=0
+ $Y2=0
cc_963 N_A_1923_174#_c_1372_n N_VPWR_c_1707_n 0.0323753f $X=10.76 $Y=2.47 $X2=0
+ $Y2=0
cc_964 N_A_1923_174#_c_1373_n N_VPWR_c_1707_n 0.00685658f $X=11.15 $Y=2.025
+ $X2=0 $Y2=0
cc_965 N_A_1923_174#_c_1371_n N_VPWR_c_1721_n 0.00653045f $X=10.73 $Y=2.69 $X2=0
+ $Y2=0
cc_966 N_A_1923_174#_M1001_g N_VPWR_c_1727_n 0.0196714f $X=9.89 $Y=2.69 $X2=0
+ $Y2=0
cc_967 N_A_1923_174#_c_1371_n N_VPWR_c_1701_n 0.00904861f $X=10.73 $Y=2.69 $X2=0
+ $Y2=0
cc_968 N_A_1923_174#_c_1365_n N_Q_N_c_2043_n 0.0248454f $X=11.15 $Y=1.94 $X2=0
+ $Y2=0
cc_969 N_A_1923_174#_c_1367_n N_Q_N_c_2043_n 0.00861348f $X=10.835 $Y=1.06 $X2=0
+ $Y2=0
cc_970 N_A_1923_174#_c_1361_n N_VGND_c_2088_n 2.70305e-19 $X=9.78 $Y=1.035 $X2=0
+ $Y2=0
cc_971 N_A_1923_174#_c_1364_n N_VGND_c_2088_n 0.0113755f $X=10.835 $Y=0.55 $X2=0
+ $Y2=0
cc_972 N_A_1923_174#_c_1366_n N_VGND_c_2088_n 0.0203737f $X=10.125 $Y=1.06 $X2=0
+ $Y2=0
cc_973 N_A_1923_174#_c_1368_n N_VGND_c_2088_n 0.00995483f $X=9.79 $Y=0.87 $X2=0
+ $Y2=0
cc_974 N_A_1923_174#_c_1364_n N_VGND_c_2089_n 0.0403776f $X=10.835 $Y=0.55 $X2=0
+ $Y2=0
cc_975 N_A_1923_174#_c_1367_n N_VGND_c_2089_n 0.00734563f $X=10.835 $Y=1.06
+ $X2=0 $Y2=0
cc_976 N_A_1923_174#_c_1368_n N_VGND_c_2100_n 0.0040395f $X=9.79 $Y=0.87 $X2=0
+ $Y2=0
cc_977 N_A_1923_174#_c_1364_n N_VGND_c_2104_n 0.0158357f $X=10.835 $Y=0.55 $X2=0
+ $Y2=0
cc_978 N_A_1923_174#_c_1363_n N_VGND_c_2113_n 0.0150349f $X=10.325 $Y=1.06 $X2=0
+ $Y2=0
cc_979 N_A_1923_174#_c_1364_n N_VGND_c_2113_n 0.0121432f $X=10.835 $Y=0.55 $X2=0
+ $Y2=0
cc_980 N_A_1923_174#_c_1366_n N_VGND_c_2113_n 0.00979114f $X=10.125 $Y=1.06
+ $X2=0 $Y2=0
cc_981 N_A_1923_174#_c_1368_n N_VGND_c_2113_n 0.00413919f $X=9.79 $Y=0.87 $X2=0
+ $Y2=0
cc_982 N_A_1770_412#_M1037_g N_A_2516_367#_c_1647_n 6.01505e-19 $X=12 $Y=0.66
+ $X2=0 $Y2=0
cc_983 N_A_1770_412#_M1011_g N_A_2516_367#_c_1647_n 0.0230531f $X=12.525 $Y=0.45
+ $X2=0 $Y2=0
cc_984 N_A_1770_412#_M1039_g N_A_2516_367#_c_1648_n 8.57075e-19 $X=11.98
+ $Y=2.465 $X2=0 $Y2=0
cc_985 N_A_1770_412#_M1029_g N_A_2516_367#_c_1648_n 0.0164902f $X=12.505
+ $Y=2.155 $X2=0 $Y2=0
cc_986 N_A_1770_412#_M1037_g N_A_2516_367#_c_1650_n 4.65144e-19 $X=12 $Y=0.66
+ $X2=0 $Y2=0
cc_987 N_A_1770_412#_M1029_g N_A_2516_367#_c_1650_n 0.00107906f $X=12.505
+ $Y=2.155 $X2=0 $Y2=0
cc_988 N_A_1770_412#_M1011_g N_A_2516_367#_c_1650_n 0.00576739f $X=12.525
+ $Y=0.45 $X2=0 $Y2=0
cc_989 N_A_1770_412#_c_1467_n N_A_2516_367#_c_1650_n 0.00830008f $X=12.515
+ $Y=1.455 $X2=0 $Y2=0
cc_990 N_A_1770_412#_M1029_g N_A_2516_367#_c_1651_n 4.48633e-19 $X=12.505
+ $Y=2.155 $X2=0 $Y2=0
cc_991 N_A_1770_412#_M1011_g N_A_2516_367#_c_1651_n 0.00481104f $X=12.525
+ $Y=0.45 $X2=0 $Y2=0
cc_992 N_A_1770_412#_M1045_g N_VPWR_c_1707_n 0.0101072f $X=10.945 $Y=2.69 $X2=0
+ $Y2=0
cc_993 N_A_1770_412#_M1007_g N_VPWR_c_1707_n 0.0143263f $X=11.55 $Y=2.465 $X2=0
+ $Y2=0
cc_994 N_A_1770_412#_M1039_g N_VPWR_c_1707_n 7.19673e-19 $X=11.98 $Y=2.465 $X2=0
+ $Y2=0
cc_995 N_A_1770_412#_M1039_g N_VPWR_c_1708_n 0.00627385f $X=11.98 $Y=2.465 $X2=0
+ $Y2=0
cc_996 N_A_1770_412#_c_1462_n N_VPWR_c_1708_n 0.00737142f $X=12.43 $Y=1.455
+ $X2=0 $Y2=0
cc_997 N_A_1770_412#_M1029_g N_VPWR_c_1708_n 0.00560522f $X=12.505 $Y=2.155
+ $X2=0 $Y2=0
cc_998 N_A_1770_412#_M1029_g N_VPWR_c_1709_n 0.00401801f $X=12.505 $Y=2.155
+ $X2=0 $Y2=0
cc_999 N_A_1770_412#_c_1490_n N_VPWR_c_1720_n 0.00818831f $X=9.765 $Y=2.58 $X2=0
+ $Y2=0
cc_1000 N_A_1770_412#_c_1481_n N_VPWR_c_1720_n 0.0112865f $X=8.99 $Y=2.58 $X2=0
+ $Y2=0
cc_1001 N_A_1770_412#_M1045_g N_VPWR_c_1721_n 0.00511894f $X=10.945 $Y=2.69
+ $X2=0 $Y2=0
cc_1002 N_A_1770_412#_M1007_g N_VPWR_c_1722_n 0.00564095f $X=11.55 $Y=2.465
+ $X2=0 $Y2=0
cc_1003 N_A_1770_412#_M1039_g N_VPWR_c_1722_n 0.00571722f $X=11.98 $Y=2.465
+ $X2=0 $Y2=0
cc_1004 N_A_1770_412#_M1029_g N_VPWR_c_1723_n 0.00312414f $X=12.505 $Y=2.155
+ $X2=0 $Y2=0
cc_1005 N_A_1770_412#_M1045_g N_VPWR_c_1727_n 7.66279e-19 $X=10.945 $Y=2.69
+ $X2=0 $Y2=0
cc_1006 N_A_1770_412#_c_1490_n N_VPWR_c_1727_n 0.0246271f $X=9.765 $Y=2.58 $X2=0
+ $Y2=0
cc_1007 N_A_1770_412#_c_1481_n N_VPWR_c_1727_n 0.00213775f $X=8.99 $Y=2.58 $X2=0
+ $Y2=0
cc_1008 N_A_1770_412#_M1045_g N_VPWR_c_1701_n 0.00526787f $X=10.945 $Y=2.69
+ $X2=0 $Y2=0
cc_1009 N_A_1770_412#_M1007_g N_VPWR_c_1701_n 0.00948291f $X=11.55 $Y=2.465
+ $X2=0 $Y2=0
cc_1010 N_A_1770_412#_M1039_g N_VPWR_c_1701_n 0.0115803f $X=11.98 $Y=2.465 $X2=0
+ $Y2=0
cc_1011 N_A_1770_412#_M1029_g N_VPWR_c_1701_n 0.00410284f $X=12.505 $Y=2.155
+ $X2=0 $Y2=0
cc_1012 N_A_1770_412#_c_1490_n N_VPWR_c_1701_n 0.0164594f $X=9.765 $Y=2.58 $X2=0
+ $Y2=0
cc_1013 N_A_1770_412#_c_1481_n N_VPWR_c_1701_n 0.0114402f $X=8.99 $Y=2.58 $X2=0
+ $Y2=0
cc_1014 N_A_1770_412#_c_1490_n A_1885_496# 0.00836024f $X=9.765 $Y=2.58
+ $X2=-0.19 $Y2=-0.245
cc_1015 N_A_1770_412#_M1007_g N_Q_N_c_2043_n 0.00429654f $X=11.55 $Y=2.465 $X2=0
+ $Y2=0
cc_1016 N_A_1770_412#_M1003_g N_Q_N_c_2043_n 0.00420574f $X=11.57 $Y=0.66 $X2=0
+ $Y2=0
cc_1017 N_A_1770_412#_c_1459_n N_Q_N_c_2043_n 0.0118528f $X=11.905 $Y=1.455
+ $X2=0 $Y2=0
cc_1018 N_A_1770_412#_M1039_g N_Q_N_c_2043_n 0.0216568f $X=11.98 $Y=2.465 $X2=0
+ $Y2=0
cc_1019 N_A_1770_412#_M1037_g N_Q_N_c_2043_n 0.00500988f $X=12 $Y=0.66 $X2=0
+ $Y2=0
cc_1020 N_A_1770_412#_M1029_g N_Q_N_c_2043_n 9.79397e-19 $X=12.505 $Y=2.155
+ $X2=0 $Y2=0
cc_1021 N_A_1770_412#_c_1466_n N_Q_N_c_2043_n 0.00451321f $X=11.99 $Y=1.455
+ $X2=0 $Y2=0
cc_1022 N_A_1770_412#_M1020_g N_VGND_c_2088_n 0.00164717f $X=10.62 $Y=0.55 $X2=0
+ $Y2=0
cc_1023 N_A_1770_412#_c_1472_n N_VGND_c_2088_n 0.00878624f $X=9.342 $Y=0.452
+ $X2=0 $Y2=0
cc_1024 N_A_1770_412#_M1020_g N_VGND_c_2089_n 0.00405198f $X=10.62 $Y=0.55 $X2=0
+ $Y2=0
cc_1025 N_A_1770_412#_c_1456_n N_VGND_c_2089_n 0.00534154f $X=11.475 $Y=1.455
+ $X2=0 $Y2=0
cc_1026 N_A_1770_412#_M1003_g N_VGND_c_2089_n 0.00338669f $X=11.57 $Y=0.66 $X2=0
+ $Y2=0
cc_1027 N_A_1770_412#_M1037_g N_VGND_c_2090_n 0.00487522f $X=12 $Y=0.66 $X2=0
+ $Y2=0
cc_1028 N_A_1770_412#_c_1462_n N_VGND_c_2090_n 0.00721663f $X=12.43 $Y=1.455
+ $X2=0 $Y2=0
cc_1029 N_A_1770_412#_M1011_g N_VGND_c_2090_n 0.00732113f $X=12.525 $Y=0.45
+ $X2=0 $Y2=0
cc_1030 N_A_1770_412#_M1011_g N_VGND_c_2091_n 0.00499168f $X=12.525 $Y=0.45
+ $X2=0 $Y2=0
cc_1031 N_A_1770_412#_c_1472_n N_VGND_c_2100_n 0.0285769f $X=9.342 $Y=0.452
+ $X2=0 $Y2=0
cc_1032 N_A_1770_412#_M1020_g N_VGND_c_2104_n 0.00457558f $X=10.62 $Y=0.55 $X2=0
+ $Y2=0
cc_1033 N_A_1770_412#_M1003_g N_VGND_c_2105_n 0.0058025f $X=11.57 $Y=0.66 $X2=0
+ $Y2=0
cc_1034 N_A_1770_412#_M1037_g N_VGND_c_2105_n 0.0058025f $X=12 $Y=0.66 $X2=0
+ $Y2=0
cc_1035 N_A_1770_412#_M1011_g N_VGND_c_2106_n 0.00545083f $X=12.525 $Y=0.45
+ $X2=0 $Y2=0
cc_1036 N_A_1770_412#_M1020_g N_VGND_c_2113_n 0.00534903f $X=10.62 $Y=0.55 $X2=0
+ $Y2=0
cc_1037 N_A_1770_412#_M1003_g N_VGND_c_2113_n 0.0118423f $X=11.57 $Y=0.66 $X2=0
+ $Y2=0
cc_1038 N_A_1770_412#_M1037_g N_VGND_c_2113_n 0.0108413f $X=12 $Y=0.66 $X2=0
+ $Y2=0
cc_1039 N_A_1770_412#_M1011_g N_VGND_c_2113_n 0.0113899f $X=12.525 $Y=0.45 $X2=0
+ $Y2=0
cc_1040 N_A_1770_412#_c_1472_n N_VGND_c_2113_n 0.0156018f $X=9.342 $Y=0.452
+ $X2=0 $Y2=0
cc_1041 N_A_2516_367#_c_1648_n N_VPWR_c_1708_n 0.0284172f $X=12.72 $Y=1.98 $X2=0
+ $Y2=0
cc_1042 N_A_2516_367#_M1008_g N_VPWR_c_1709_n 0.0197302f $X=13.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1043 N_A_2516_367#_M1026_g N_VPWR_c_1709_n 7.82599e-19 $X=13.905 $Y=2.465
+ $X2=0 $Y2=0
cc_1044 N_A_2516_367#_c_1648_n N_VPWR_c_1709_n 0.0483698f $X=12.72 $Y=1.98 $X2=0
+ $Y2=0
cc_1045 N_A_2516_367#_c_1649_n N_VPWR_c_1709_n 0.0194308f $X=13.32 $Y=1.395
+ $X2=0 $Y2=0
cc_1046 N_A_2516_367#_c_1651_n N_VPWR_c_1709_n 0.00544712f $X=13.905 $Y=1.395
+ $X2=0 $Y2=0
cc_1047 N_A_2516_367#_M1026_g N_VPWR_c_1711_n 0.0077624f $X=13.905 $Y=2.465
+ $X2=0 $Y2=0
cc_1048 N_A_2516_367#_M1008_g N_VPWR_c_1724_n 0.00564095f $X=13.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1049 N_A_2516_367#_M1026_g N_VPWR_c_1724_n 0.00583607f $X=13.905 $Y=2.465
+ $X2=0 $Y2=0
cc_1050 N_A_2516_367#_M1008_g N_VPWR_c_1701_n 0.00948291f $X=13.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1051 N_A_2516_367#_M1026_g N_VPWR_c_1701_n 0.0114326f $X=13.905 $Y=2.465
+ $X2=0 $Y2=0
cc_1052 N_A_2516_367#_c_1648_n N_VPWR_c_1701_n 0.0121821f $X=12.72 $Y=1.98 $X2=0
+ $Y2=0
cc_1053 N_A_2516_367#_c_1647_n N_Q_N_c_2043_n 0.00368404f $X=12.74 $Y=0.45 $X2=0
+ $Y2=0
cc_1054 N_A_2516_367#_c_1648_n N_Q_N_c_2043_n 0.00554875f $X=12.72 $Y=1.98 $X2=0
+ $Y2=0
cc_1055 N_A_2516_367#_c_1650_n N_Q_N_c_2043_n 0.0088304f $X=12.74 $Y=1.395 $X2=0
+ $Y2=0
cc_1056 N_A_2516_367#_c_1643_n N_Q_c_2065_n 0.00251344f $X=13.475 $Y=1.23 $X2=0
+ $Y2=0
cc_1057 N_A_2516_367#_M1008_g N_Q_c_2065_n 0.00754289f $X=13.475 $Y=2.465 $X2=0
+ $Y2=0
cc_1058 N_A_2516_367#_c_1645_n N_Q_c_2065_n 0.00347385f $X=13.905 $Y=1.23 $X2=0
+ $Y2=0
cc_1059 N_A_2516_367#_M1026_g N_Q_c_2065_n 0.00759462f $X=13.905 $Y=2.465 $X2=0
+ $Y2=0
cc_1060 N_A_2516_367#_c_1647_n N_Q_c_2065_n 0.00430873f $X=12.74 $Y=0.45 $X2=0
+ $Y2=0
cc_1061 N_A_2516_367#_c_1649_n N_Q_c_2065_n 0.0255555f $X=13.32 $Y=1.395 $X2=0
+ $Y2=0
cc_1062 N_A_2516_367#_c_1651_n N_Q_c_2065_n 0.0299442f $X=13.905 $Y=1.395 $X2=0
+ $Y2=0
cc_1063 N_A_2516_367#_c_1647_n N_VGND_c_2090_n 0.0483659f $X=12.74 $Y=0.45 $X2=0
+ $Y2=0
cc_1064 N_A_2516_367#_c_1643_n N_VGND_c_2091_n 0.0125932f $X=13.475 $Y=1.23
+ $X2=0 $Y2=0
cc_1065 N_A_2516_367#_c_1645_n N_VGND_c_2091_n 5.5046e-19 $X=13.905 $Y=1.23
+ $X2=0 $Y2=0
cc_1066 N_A_2516_367#_c_1647_n N_VGND_c_2091_n 0.0593959f $X=12.74 $Y=0.45 $X2=0
+ $Y2=0
cc_1067 N_A_2516_367#_c_1649_n N_VGND_c_2091_n 0.0231351f $X=13.32 $Y=1.395
+ $X2=0 $Y2=0
cc_1068 N_A_2516_367#_c_1651_n N_VGND_c_2091_n 0.00553375f $X=13.905 $Y=1.395
+ $X2=0 $Y2=0
cc_1069 N_A_2516_367#_c_1645_n N_VGND_c_2093_n 0.00710381f $X=13.905 $Y=1.23
+ $X2=0 $Y2=0
cc_1070 N_A_2516_367#_c_1647_n N_VGND_c_2106_n 0.0176612f $X=12.74 $Y=0.45 $X2=0
+ $Y2=0
cc_1071 N_A_2516_367#_c_1643_n N_VGND_c_2107_n 0.00521096f $X=13.475 $Y=1.23
+ $X2=0 $Y2=0
cc_1072 N_A_2516_367#_c_1645_n N_VGND_c_2107_n 0.00539121f $X=13.905 $Y=1.23
+ $X2=0 $Y2=0
cc_1073 N_A_2516_367#_M1011_d N_VGND_c_2113_n 0.00215771f $X=12.6 $Y=0.24 $X2=0
+ $Y2=0
cc_1074 N_A_2516_367#_c_1643_n N_VGND_c_2113_n 0.00936705f $X=13.475 $Y=1.23
+ $X2=0 $Y2=0
cc_1075 N_A_2516_367#_c_1645_n N_VGND_c_2113_n 0.0109079f $X=13.905 $Y=1.23
+ $X2=0 $Y2=0
cc_1076 N_A_2516_367#_c_1647_n N_VGND_c_2113_n 0.0124419f $X=12.74 $Y=0.45 $X2=0
+ $Y2=0
cc_1077 N_VPWR_c_1701_n A_287_489# 0.00899413f $X=14.16 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1078 N_VPWR_c_1701_n N_A_359_489#_M1009_d 0.00223559f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1079 N_VPWR_c_1701_n N_A_359_489#_M1002_d 0.00212301f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1080 N_VPWR_M1034_d N_A_359_489#_c_1916_n 0.00784053f $X=2.695 $Y=2.445 $X2=0
+ $Y2=0
cc_1081 N_VPWR_c_1703_n N_A_359_489#_c_1916_n 0.0181839f $X=2.835 $Y=2.94 $X2=0
+ $Y2=0
cc_1082 N_VPWR_c_1712_n N_A_359_489#_c_1916_n 0.00811461f $X=2.67 $Y=3.33 $X2=0
+ $Y2=0
cc_1083 N_VPWR_c_1701_n N_A_359_489#_c_1916_n 0.0160069f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1084 N_VPWR_M1042_d N_A_359_489#_c_1907_n 0.00413003f $X=4.24 $Y=1.835 $X2=0
+ $Y2=0
cc_1085 N_VPWR_c_1704_n N_A_359_489#_c_1907_n 0.0161939f $X=4.38 $Y=2.93 $X2=0
+ $Y2=0
cc_1086 N_VPWR_c_1714_n N_A_359_489#_c_1907_n 0.0104637f $X=4.215 $Y=3.33 $X2=0
+ $Y2=0
cc_1087 N_VPWR_c_1716_n N_A_359_489#_c_1907_n 0.0124534f $X=6.69 $Y=3.33 $X2=0
+ $Y2=0
cc_1088 N_VPWR_c_1701_n N_A_359_489#_c_1907_n 0.0397619f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1089 N_VPWR_M1034_d N_A_359_489#_c_1908_n 7.97895e-19 $X=2.695 $Y=2.445 $X2=0
+ $Y2=0
cc_1090 N_VPWR_c_1703_n N_A_359_489#_c_1908_n 0.00194376f $X=2.835 $Y=2.94 $X2=0
+ $Y2=0
cc_1091 N_VPWR_c_1714_n N_A_359_489#_c_1908_n 0.00294609f $X=4.215 $Y=3.33 $X2=0
+ $Y2=0
cc_1092 N_VPWR_c_1701_n N_A_359_489#_c_1908_n 0.00560275f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1093 N_VPWR_c_1702_n N_A_359_489#_c_1912_n 0.0211092f $X=1.145 $Y=2.6 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1703_n N_A_359_489#_c_1912_n 0.0066483f $X=2.835 $Y=2.94 $X2=0
+ $Y2=0
cc_1095 N_VPWR_c_1712_n N_A_359_489#_c_1912_n 0.0188411f $X=2.67 $Y=3.33 $X2=0
+ $Y2=0
cc_1096 N_VPWR_c_1701_n N_A_359_489#_c_1912_n 0.0123607f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1097 N_VPWR_c_1703_n N_A_359_489#_c_1913_n 0.0158355f $X=2.835 $Y=2.94 $X2=0
+ $Y2=0
cc_1098 N_VPWR_c_1704_n N_A_359_489#_c_1913_n 0.0069225f $X=4.38 $Y=2.93 $X2=0
+ $Y2=0
cc_1099 N_VPWR_c_1714_n N_A_359_489#_c_1913_n 0.0208498f $X=4.215 $Y=3.33 $X2=0
+ $Y2=0
cc_1100 N_VPWR_c_1701_n N_A_359_489#_c_1913_n 0.012522f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1101 N_VPWR_c_1716_n N_A_359_489#_c_1914_n 0.00454945f $X=6.69 $Y=3.33 $X2=0
+ $Y2=0
cc_1102 N_VPWR_c_1701_n N_A_359_489#_c_1914_n 0.00682782f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1103 N_VPWR_c_1701_n A_445_489# 0.00390756f $X=14.16 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1104 N_VPWR_c_1727_n A_1885_496# 0.00129994f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1105 N_VPWR_c_1701_n N_Q_N_M1007_d 0.00310528f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1106 N_VPWR_c_1708_n N_Q_N_c_2043_n 0.0480563f $X=12.24 $Y=1.96 $X2=0 $Y2=0
cc_1107 N_VPWR_c_1722_n N_Q_N_c_2043_n 0.0153751f $X=12.085 $Y=3.33 $X2=0 $Y2=0
cc_1108 N_VPWR_c_1701_n N_Q_N_c_2043_n 0.0101105f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1109 N_VPWR_c_1701_n N_Q_M1008_s 0.00380103f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1110 N_VPWR_c_1709_n N_Q_c_2065_n 0.0475786f $X=13.26 $Y=1.98 $X2=0 $Y2=0
cc_1111 N_VPWR_c_1711_n N_Q_c_2065_n 0.0446985f $X=14.12 $Y=1.98 $X2=0 $Y2=0
cc_1112 N_VPWR_c_1724_n N_Q_c_2065_n 0.0140491f $X=13.98 $Y=3.33 $X2=0 $Y2=0
cc_1113 N_VPWR_c_1701_n N_Q_c_2065_n 0.0090585f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1114 N_VPWR_c_1711_n N_VGND_c_2093_n 0.0107653f $X=14.12 $Y=1.98 $X2=0 $Y2=0
cc_1115 N_A_359_489#_c_1916_n A_445_489# 0.00984236f $X=2.975 $Y=2.55 $X2=-0.19
+ $Y2=-0.245
cc_1116 N_A_359_489#_c_1902_n N_VGND_c_2113_n 0.00168329f $X=2.975 $Y=0.88 $X2=0
+ $Y2=0
cc_1117 N_A_359_489#_c_1902_n N_noxref_25_M1047_d 0.00182394f $X=2.975 $Y=0.88
+ $X2=0 $Y2=0
cc_1118 N_A_359_489#_M1035_d N_noxref_25_c_2245_n 0.00199854f $X=1.975 $Y=0.405
+ $X2=0 $Y2=0
cc_1119 N_A_359_489#_c_1902_n N_noxref_25_c_2245_n 0.0146573f $X=2.975 $Y=0.88
+ $X2=0 $Y2=0
cc_1120 N_A_359_489#_c_1905_n N_noxref_25_c_2245_n 0.0154818f $X=2.14 $Y=0.7
+ $X2=0 $Y2=0
cc_1121 N_A_359_489#_c_1905_n N_noxref_25_c_2246_n 0.00290675f $X=2.14 $Y=0.7
+ $X2=0 $Y2=0
cc_1122 N_A_359_489#_c_1902_n N_noxref_25_c_2247_n 0.0151225f $X=2.975 $Y=0.88
+ $X2=0 $Y2=0
cc_1123 N_A_359_489#_c_1905_n N_noxref_25_c_2247_n 5.76861e-19 $X=2.14 $Y=0.7
+ $X2=0 $Y2=0
cc_1124 N_A_359_489#_c_1902_n noxref_27 0.00266636f $X=2.975 $Y=0.88 $X2=-0.19
+ $Y2=-0.245
cc_1125 N_Q_N_c_2043_n N_VGND_c_2090_n 0.00114318f $X=11.785 $Y=0.42 $X2=0 $Y2=0
cc_1126 N_Q_N_c_2043_n N_VGND_c_2105_n 0.0151136f $X=11.785 $Y=0.42 $X2=0 $Y2=0
cc_1127 N_Q_N_M1003_s N_VGND_c_2113_n 0.0027574f $X=11.645 $Y=0.24 $X2=0 $Y2=0
cc_1128 N_Q_N_c_2043_n N_VGND_c_2113_n 0.0102248f $X=11.785 $Y=0.42 $X2=0 $Y2=0
cc_1129 N_Q_c_2065_n N_VGND_c_2091_n 0.0308662f $X=13.69 $Y=0.42 $X2=0 $Y2=0
cc_1130 N_Q_c_2065_n N_VGND_c_2093_n 0.0314226f $X=13.69 $Y=0.42 $X2=0 $Y2=0
cc_1131 N_Q_c_2065_n N_VGND_c_2107_n 0.016703f $X=13.69 $Y=0.42 $X2=0 $Y2=0
cc_1132 N_Q_c_2065_n N_VGND_c_2113_n 0.0090585f $X=13.69 $Y=0.42 $X2=0 $Y2=0
cc_1133 N_VGND_c_2094_n N_noxref_25_c_2245_n 0.0820806f $X=3.35 $Y=0 $X2=0 $Y2=0
cc_1134 N_VGND_c_2113_n N_noxref_25_c_2245_n 0.0502516f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1135 N_VGND_c_2083_n N_noxref_25_c_2246_n 0.029516f $X=0.69 $Y=0.6 $X2=0
+ $Y2=0
cc_1136 N_VGND_c_2094_n N_noxref_25_c_2246_n 0.0233489f $X=3.35 $Y=0 $X2=0 $Y2=0
cc_1137 N_VGND_c_2113_n N_noxref_25_c_2246_n 0.0125854f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1138 N_VGND_c_2084_n N_noxref_25_c_2247_n 0.0190884f $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_1139 N_VGND_c_2094_n N_noxref_25_c_2247_n 0.0210242f $X=3.35 $Y=0 $X2=0 $Y2=0
cc_1140 N_VGND_c_2113_n N_noxref_25_c_2247_n 0.0123731f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1141 N_noxref_25_c_2245_n noxref_26 0.00154828f $X=2.85 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_1142 N_noxref_25_c_2245_n noxref_27 0.00270557f $X=2.85 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
