* File: sky130_fd_sc_lp__dlrtn_4.pxi.spice
* Created: Wed Sep  2 09:47:03 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTN_4%D N_D_c_161_n N_D_M1022_g N_D_M1016_g N_D_c_163_n
+ D D D N_D_c_165_n N_D_c_166_n PM_SKY130_FD_SC_LP__DLRTN_4%D
x_PM_SKY130_FD_SC_LP__DLRTN_4%GATE_N N_GATE_N_M1001_g N_GATE_N_M1005_g GATE_N
+ N_GATE_N_c_204_n N_GATE_N_c_205_n PM_SKY130_FD_SC_LP__DLRTN_4%GATE_N
x_PM_SKY130_FD_SC_LP__DLRTN_4%A_27_468# N_A_27_468#_M1016_s N_A_27_468#_M1022_s
+ N_A_27_468#_M1003_g N_A_27_468#_M1010_g N_A_27_468#_c_236_n
+ N_A_27_468#_c_243_n N_A_27_468#_c_237_n N_A_27_468#_c_245_n
+ N_A_27_468#_c_257_n N_A_27_468#_c_246_n N_A_27_468#_c_247_n
+ N_A_27_468#_c_248_n N_A_27_468#_c_273_p N_A_27_468#_c_249_n
+ N_A_27_468#_c_238_n N_A_27_468#_c_239_n N_A_27_468#_c_240_n
+ N_A_27_468#_c_251_n PM_SKY130_FD_SC_LP__DLRTN_4%A_27_468#
x_PM_SKY130_FD_SC_LP__DLRTN_4%A_357_365# N_A_357_365#_M1017_s
+ N_A_357_365#_M1002_s N_A_357_365#_M1013_g N_A_357_365#_M1000_g
+ N_A_357_365#_c_357_n N_A_357_365#_c_345_n N_A_357_365#_c_346_n
+ N_A_357_365#_c_347_n N_A_357_365#_c_348_n N_A_357_365#_c_349_n
+ N_A_357_365#_c_350_n N_A_357_365#_c_351_n N_A_357_365#_c_352_n
+ N_A_357_365#_c_353_n N_A_357_365#_c_354_n N_A_357_365#_c_360_n
+ N_A_357_365#_c_355_n PM_SKY130_FD_SC_LP__DLRTN_4%A_357_365#
x_PM_SKY130_FD_SC_LP__DLRTN_4%A_250_70# N_A_250_70#_M1001_d N_A_250_70#_M1005_d
+ N_A_250_70#_c_459_n N_A_250_70#_c_460_n N_A_250_70#_c_461_n
+ N_A_250_70#_M1017_g N_A_250_70#_M1002_g N_A_250_70#_M1024_g
+ N_A_250_70#_c_464_n N_A_250_70#_c_465_n N_A_250_70#_c_466_n
+ N_A_250_70#_M1020_g N_A_250_70#_c_467_n N_A_250_70#_c_468_n
+ N_A_250_70#_c_469_n N_A_250_70#_c_470_n N_A_250_70#_c_478_n
+ N_A_250_70#_c_471_n N_A_250_70#_c_472_n PM_SKY130_FD_SC_LP__DLRTN_4%A_250_70#
x_PM_SKY130_FD_SC_LP__DLRTN_4%A_789_99# N_A_789_99#_M1018_s N_A_789_99#_M1019_d
+ N_A_789_99#_c_578_n N_A_789_99#_M1004_g N_A_789_99#_M1008_g
+ N_A_789_99#_M1007_g N_A_789_99#_M1011_g N_A_789_99#_M1012_g
+ N_A_789_99#_M1014_g N_A_789_99#_M1021_g N_A_789_99#_M1015_g
+ N_A_789_99#_M1023_g N_A_789_99#_M1025_g N_A_789_99#_c_584_n
+ N_A_789_99#_c_598_n N_A_789_99#_c_585_n N_A_789_99#_c_613_p
+ N_A_789_99#_c_608_n N_A_789_99#_c_586_n N_A_789_99#_c_633_p
+ N_A_789_99#_c_587_n N_A_789_99#_c_636_p N_A_789_99#_c_588_n
+ N_A_789_99#_c_589_n N_A_789_99#_c_693_p N_A_789_99#_c_649_p
+ N_A_789_99#_c_590_n N_A_789_99#_c_591_n PM_SKY130_FD_SC_LP__DLRTN_4%A_789_99#
x_PM_SKY130_FD_SC_LP__DLRTN_4%A_639_125# N_A_639_125#_M1024_d
+ N_A_639_125#_M1013_d N_A_639_125#_c_750_n N_A_639_125#_M1018_g
+ N_A_639_125#_M1019_g N_A_639_125#_c_752_n N_A_639_125#_c_753_n
+ N_A_639_125#_c_764_n N_A_639_125#_c_768_n N_A_639_125#_c_754_n
+ N_A_639_125#_c_755_n N_A_639_125#_c_759_n N_A_639_125#_c_756_n
+ N_A_639_125#_c_757_n PM_SKY130_FD_SC_LP__DLRTN_4%A_639_125#
x_PM_SKY130_FD_SC_LP__DLRTN_4%RESET_B N_RESET_B_M1009_g N_RESET_B_M1006_g
+ RESET_B RESET_B RESET_B N_RESET_B_c_837_n PM_SKY130_FD_SC_LP__DLRTN_4%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTN_4%VPWR N_VPWR_M1022_d N_VPWR_M1002_d N_VPWR_M1008_d
+ N_VPWR_M1006_d N_VPWR_M1014_d N_VPWR_M1025_d N_VPWR_c_881_n N_VPWR_c_882_n
+ N_VPWR_c_883_n N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n
+ N_VPWR_c_888_n N_VPWR_c_889_n N_VPWR_c_890_n VPWR N_VPWR_c_891_n
+ N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n
+ N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_880_n PM_SKY130_FD_SC_LP__DLRTN_4%VPWR
x_PM_SKY130_FD_SC_LP__DLRTN_4%Q N_Q_M1011_d N_Q_M1021_d N_Q_M1007_s N_Q_M1015_s
+ N_Q_c_997_n N_Q_c_1031_n N_Q_c_986_n N_Q_c_987_n N_Q_c_992_n N_Q_c_993_n
+ N_Q_c_1016_n N_Q_c_1035_n N_Q_c_988_n N_Q_c_994_n N_Q_c_1022_n N_Q_c_989_n
+ N_Q_c_995_n Q N_Q_c_990_n Q PM_SKY130_FD_SC_LP__DLRTN_4%Q
x_PM_SKY130_FD_SC_LP__DLRTN_4%VGND N_VGND_M1016_d N_VGND_M1017_d N_VGND_M1004_d
+ N_VGND_M1009_d N_VGND_M1012_s N_VGND_M1023_s N_VGND_c_1048_n N_VGND_c_1049_n
+ N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n N_VGND_c_1053_n
+ N_VGND_c_1054_n N_VGND_c_1055_n N_VGND_c_1056_n N_VGND_c_1057_n
+ N_VGND_c_1058_n VGND N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n
+ N_VGND_c_1062_n N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n
+ N_VGND_c_1066_n PM_SKY130_FD_SC_LP__DLRTN_4%VGND
cc_1 VNB N_D_c_161_n 0.0201985f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.34
cc_2 VNB N_D_M1022_g 0.0060756f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_3 VNB N_D_c_163_n 0.0243765f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.55
cc_4 VNB D 0.00991979f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_5 VNB N_D_c_165_n 0.0245758f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.045
cc_6 VNB N_D_c_166_n 0.0204468f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.88
cc_7 VNB N_GATE_N_M1001_g 0.0614037f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.55
cc_8 VNB N_A_27_468#_M1003_g 0.0265885f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.56
cc_9 VNB N_A_27_468#_c_236_n 0.00640119f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.045
cc_10 VNB N_A_27_468#_c_237_n 0.0527061f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.88
cc_11 VNB N_A_27_468#_c_238_n 0.00171403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_468#_c_239_n 0.0166544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_468#_c_240_n 0.0231449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_357_365#_c_345_n 6.56039e-19 $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.88
cc_15 VNB N_A_357_365#_c_346_n 0.00166744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_357_365#_c_347_n 0.0138281f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.045
cc_17 VNB N_A_357_365#_c_348_n 0.00548938f $X=-0.19 $Y=-0.245 $X2=0.775
+ $Y2=1.295
cc_18 VNB N_A_357_365#_c_349_n 0.00168179f $X=-0.19 $Y=-0.245 $X2=0.775
+ $Y2=1.665
cc_19 VNB N_A_357_365#_c_350_n 0.00248766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_357_365#_c_351_n 0.00749085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_357_365#_c_352_n 0.0402007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_357_365#_c_353_n 0.011473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_357_365#_c_354_n 0.00324024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_357_365#_c_355_n 0.0144761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_250_70#_c_459_n 0.0600248f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.56
cc_26 VNB N_A_250_70#_c_460_n 0.105586f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.56
cc_27 VNB N_A_250_70#_c_461_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.55
cc_28 VNB N_A_250_70#_M1017_g 0.0252683f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_29 VNB N_A_250_70#_M1024_g 0.0373175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_250_70#_c_464_n 0.0266134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_250_70#_c_465_n 0.00644547f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.045
cc_32 VNB N_A_250_70#_c_466_n 0.0159593f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.295
cc_33 VNB N_A_250_70#_c_467_n 0.0105038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_250_70#_c_468_n 0.0208581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_250_70#_c_469_n 0.0113526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_250_70#_c_470_n 0.0156465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_250_70#_c_471_n 0.0030404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_250_70#_c_472_n 0.0032972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_789_99#_c_578_n 0.0326891f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.88
cc_40 VNB N_A_789_99#_M1004_g 0.0210807f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.56
cc_41 VNB N_A_789_99#_M1011_g 0.0243338f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.925
cc_42 VNB N_A_789_99#_M1012_g 0.0226933f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.295
cc_43 VNB N_A_789_99#_M1021_g 0.0226791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_789_99#_M1023_g 0.0279341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_789_99#_c_584_n 0.00686792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_789_99#_c_585_n 0.00144614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_789_99#_c_586_n 0.00499195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_789_99#_c_587_n 0.00178699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_789_99#_c_588_n 0.00266611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_789_99#_c_589_n 3.61316e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_789_99#_c_590_n 0.00103189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_789_99#_c_591_n 0.0667522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_639_125#_c_750_n 0.0188603f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.88
cc_54 VNB N_A_639_125#_M1019_g 0.0080726f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_55 VNB N_A_639_125#_c_752_n 0.0434183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_639_125#_c_753_n 0.00877605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_639_125#_c_754_n 0.0352219f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.045
cc_58 VNB N_A_639_125#_c_755_n 0.00960535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_639_125#_c_756_n 0.0035867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_639_125#_c_757_n 3.98181e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_M1009_g 0.0185464f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.55
cc_62 VNB N_RESET_B_M1006_g 0.00514095f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.88
cc_63 VNB RESET_B 0.0037508f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.56
cc_64 VNB N_RESET_B_c_837_n 0.0323256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VPWR_c_880_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_986_n 0.0086357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_Q_c_987_n 0.00271466f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.045
cc_68 VNB N_Q_c_988_n 0.00353859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_c_989_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_Q_c_990_n 0.0108368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB Q 0.0202259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1048_n 0.00344978f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.925
cc_73 VNB N_VGND_c_1049_n 0.00958361f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.295
cc_74 VNB N_VGND_c_1050_n 0.0161061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1051_n 0.00501995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1052_n 3.22457e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1053_n 0.0106846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1054_n 0.029201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1055_n 0.02285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1056_n 0.00579822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1057_n 0.0333054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1058_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1059_n 0.036123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1060_n 0.0292388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1061_n 0.0157463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1062_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1063_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1064_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1065_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1066_n 0.399889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VPB N_D_M1022_g 0.0554558f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_92 VPB D 0.00497016f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_93 VPB N_GATE_N_M1001_g 0.0124914f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.55
cc_94 VPB N_GATE_N_M1005_g 0.026022f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.88
cc_95 VPB N_GATE_N_c_204_n 0.00404481f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_96 VPB N_GATE_N_c_205_n 0.0453494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_27_468#_M1010_g 0.0190466f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_98 VPB N_A_27_468#_c_236_n 0.0180673f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.045
cc_99 VPB N_A_27_468#_c_243_n 0.0163685f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.045
cc_100 VPB N_A_27_468#_c_237_n 0.0350558f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.88
cc_101 VPB N_A_27_468#_c_245_n 0.00583544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_27_468#_c_246_n 0.0153862f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.665
cc_103 VPB N_A_27_468#_c_247_n 0.00134151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_27_468#_c_248_n 0.00462687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_27_468#_c_249_n 0.00309813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_27_468#_c_238_n 0.00159938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_27_468#_c_251_n 0.0289766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_357_365#_M1013_g 0.0229729f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.56
cc_109 VPB N_A_357_365#_c_357_n 0.00483794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_357_365#_c_346_n 0.00267243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_357_365#_c_354_n 0.00283169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_357_365#_c_360_n 0.0310256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_250_70#_M1002_g 0.0484935f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.045
cc_114 VPB N_A_250_70#_c_466_n 0.00198313f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.295
cc_115 VPB N_A_250_70#_M1020_g 0.0363201f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.665
cc_116 VPB N_A_250_70#_c_467_n 0.00732811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_250_70#_c_468_n 0.0104948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_250_70#_c_478_n 0.0171929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_250_70#_c_471_n 0.0030404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_789_99#_M1008_g 0.0222644f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_121 VPB N_A_789_99#_M1007_g 0.0189309f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.045
cc_122 VPB N_A_789_99#_M1014_g 0.0180412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_789_99#_M1015_g 0.0179089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_789_99#_M1025_g 0.0212849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_789_99#_c_584_n 0.0207673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_789_99#_c_598_n 0.0185997f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_789_99#_c_585_n 0.00232953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_789_99#_c_589_n 0.00110232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_789_99#_c_591_n 0.0111314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_639_125#_M1019_g 0.0230243f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_131 VPB N_A_639_125#_c_759_n 0.00926756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_639_125#_c_756_n 0.00459988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_RESET_B_M1006_g 0.0191571f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.88
cc_134 VPB RESET_B 0.00117856f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.56
cc_135 VPB N_VPWR_c_881_n 0.00538429f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.925
cc_136 VPB N_VPWR_c_882_n 0.0167255f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.295
cc_137 VPB N_VPWR_c_883_n 0.0164981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_884_n 0.0146078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_885_n 0.00431328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_886_n 3.16879e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_887_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_888_n 0.0412014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_889_n 0.0580188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_890_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_891_n 0.0167011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_892_n 0.0403753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_893_n 0.0154186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_894_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_895_n 0.00445824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_896_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_897_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_898_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_880_n 0.104535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_Q_c_992_n 0.00304538f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.295
cc_155 VPB N_Q_c_993_n 0.00191919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_Q_c_994_n 0.0100496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_Q_c_995_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB Q 0.00555106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 N_D_M1022_g N_GATE_N_M1001_g 0.00556423f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_160 D N_GATE_N_M1001_g 0.00891973f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_161 N_D_c_166_n N_GATE_N_M1001_g 0.041348f $X=0.61 $Y=0.88 $X2=0 $Y2=0
cc_162 N_D_M1022_g N_GATE_N_M1005_g 0.0137512f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_163 N_D_M1022_g N_GATE_N_c_204_n 0.00193835f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_164 N_D_c_163_n N_GATE_N_c_204_n 7.1555e-19 $X=0.61 $Y=1.55 $X2=0 $Y2=0
cc_165 D N_GATE_N_c_204_n 0.0318004f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_166 N_D_M1022_g N_GATE_N_c_205_n 0.0172433f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_167 N_D_c_163_n N_GATE_N_c_205_n 0.00116823f $X=0.61 $Y=1.55 $X2=0 $Y2=0
cc_168 D N_GATE_N_c_205_n 0.00517239f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_169 D N_A_27_468#_c_237_n 0.0729416f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_170 N_D_c_165_n N_A_27_468#_c_237_n 0.043141f $X=0.655 $Y=1.045 $X2=0 $Y2=0
cc_171 N_D_c_166_n N_A_27_468#_c_237_n 0.00524177f $X=0.61 $Y=0.88 $X2=0 $Y2=0
cc_172 N_D_M1022_g N_A_27_468#_c_245_n 0.0155356f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_173 D N_A_27_468#_c_245_n 0.00348399f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_174 N_D_M1022_g N_A_27_468#_c_257_n 0.00130649f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_175 N_D_M1022_g N_A_27_468#_c_247_n 3.48984e-19 $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_176 D N_A_27_468#_c_240_n 0.00706386f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_177 N_D_c_165_n N_A_27_468#_c_240_n 0.00635427f $X=0.655 $Y=1.045 $X2=0 $Y2=0
cc_178 N_D_c_166_n N_A_27_468#_c_240_n 4.34564e-19 $X=0.61 $Y=0.88 $X2=0 $Y2=0
cc_179 N_D_M1022_g N_A_27_468#_c_251_n 4.52926e-19 $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_180 D N_A_250_70#_c_470_n 0.0323383f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_181 D N_A_250_70#_c_478_n 0.00553185f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_182 D N_A_250_70#_c_472_n 0.0165394f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_183 N_D_M1022_g N_VPWR_c_881_n 0.00970612f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_184 N_D_M1022_g N_VPWR_c_891_n 0.00428763f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_185 N_D_M1022_g N_VPWR_c_880_n 0.00446945f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_186 D N_VGND_c_1048_n 0.0167671f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_187 N_D_c_166_n N_VGND_c_1048_n 0.0101922f $X=0.61 $Y=0.88 $X2=0 $Y2=0
cc_188 N_D_c_166_n N_VGND_c_1055_n 0.00396895f $X=0.61 $Y=0.88 $X2=0 $Y2=0
cc_189 D N_VGND_c_1066_n 0.00672098f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_190 N_D_c_166_n N_VGND_c_1066_n 0.0041875f $X=0.61 $Y=0.88 $X2=0 $Y2=0
cc_191 N_GATE_N_c_204_n N_A_27_468#_c_237_n 0.0139939f $X=0.955 $Y=2.015 $X2=0
+ $Y2=0
cc_192 N_GATE_N_M1005_g N_A_27_468#_c_245_n 0.00534158f $X=1.175 $Y=2.66 $X2=0
+ $Y2=0
cc_193 N_GATE_N_c_204_n N_A_27_468#_c_245_n 0.0378536f $X=0.955 $Y=2.015 $X2=0
+ $Y2=0
cc_194 N_GATE_N_c_205_n N_A_27_468#_c_245_n 0.00732602f $X=1.175 $Y=2.015 $X2=0
+ $Y2=0
cc_195 N_GATE_N_M1005_g N_A_27_468#_c_257_n 0.00929464f $X=1.175 $Y=2.66 $X2=0
+ $Y2=0
cc_196 N_GATE_N_M1005_g N_A_27_468#_c_246_n 0.0126617f $X=1.175 $Y=2.66 $X2=0
+ $Y2=0
cc_197 N_GATE_N_M1005_g N_A_27_468#_c_247_n 0.00269018f $X=1.175 $Y=2.66 $X2=0
+ $Y2=0
cc_198 N_GATE_N_M1005_g N_A_27_468#_c_248_n 0.00304436f $X=1.175 $Y=2.66 $X2=0
+ $Y2=0
cc_199 N_GATE_N_M1001_g N_A_250_70#_c_461_n 0.0368417f $X=1.175 $Y=0.56 $X2=0
+ $Y2=0
cc_200 N_GATE_N_M1001_g N_A_250_70#_c_470_n 0.00771884f $X=1.175 $Y=0.56 $X2=0
+ $Y2=0
cc_201 N_GATE_N_M1001_g N_A_250_70#_c_478_n 0.0233958f $X=1.175 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_GATE_N_c_204_n N_A_250_70#_c_478_n 0.0180323f $X=0.955 $Y=2.015 $X2=0
+ $Y2=0
cc_203 N_GATE_N_M1001_g N_A_250_70#_c_472_n 0.00288057f $X=1.175 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_GATE_N_M1005_g N_VPWR_c_881_n 0.00310435f $X=1.175 $Y=2.66 $X2=0 $Y2=0
cc_205 N_GATE_N_M1005_g N_VPWR_c_892_n 0.00299966f $X=1.175 $Y=2.66 $X2=0 $Y2=0
cc_206 N_GATE_N_M1005_g N_VPWR_c_880_n 0.00428799f $X=1.175 $Y=2.66 $X2=0 $Y2=0
cc_207 N_GATE_N_M1001_g N_VGND_c_1048_n 0.00882944f $X=1.175 $Y=0.56 $X2=0 $Y2=0
cc_208 N_GATE_N_M1001_g N_VGND_c_1057_n 0.00396895f $X=1.175 $Y=0.56 $X2=0 $Y2=0
cc_209 N_GATE_N_M1001_g N_VGND_c_1066_n 0.00774381f $X=1.175 $Y=0.56 $X2=0 $Y2=0
cc_210 N_A_27_468#_c_246_n N_A_357_365#_M1002_s 0.0010603f $X=1.675 $Y=2.915
+ $X2=0 $Y2=0
cc_211 N_A_27_468#_c_248_n N_A_357_365#_M1002_s 0.00872491f $X=1.842 $Y=2.83
+ $X2=0 $Y2=0
cc_212 N_A_27_468#_c_273_p N_A_357_365#_M1002_s 0.00369196f $X=2.505 $Y=2.36
+ $X2=0 $Y2=0
cc_213 N_A_27_468#_c_249_n N_A_357_365#_M1002_s 0.00398708f $X=2.01 $Y=2.36
+ $X2=0 $Y2=0
cc_214 N_A_27_468#_c_243_n N_A_357_365#_M1013_g 0.0376618f $X=2.67 $Y=2.075
+ $X2=0 $Y2=0
cc_215 N_A_27_468#_c_273_p N_A_357_365#_M1013_g 5.74605e-19 $X=2.505 $Y=2.36
+ $X2=0 $Y2=0
cc_216 N_A_27_468#_c_236_n N_A_357_365#_c_357_n 8.35496e-19 $X=2.67 $Y=1.91
+ $X2=0 $Y2=0
cc_217 N_A_27_468#_c_273_p N_A_357_365#_c_357_n 0.0179531f $X=2.505 $Y=2.36
+ $X2=0 $Y2=0
cc_218 N_A_27_468#_c_249_n N_A_357_365#_c_357_n 0.0224396f $X=2.01 $Y=2.36 $X2=0
+ $Y2=0
cc_219 N_A_27_468#_c_238_n N_A_357_365#_c_357_n 0.0169812f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_220 N_A_27_468#_M1003_g N_A_357_365#_c_346_n 9.96596e-19 $X=2.76 $Y=0.835
+ $X2=0 $Y2=0
cc_221 N_A_27_468#_c_238_n N_A_357_365#_c_346_n 0.0230739f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_222 N_A_27_468#_c_239_n N_A_357_365#_c_346_n 0.00140979f $X=2.67 $Y=1.57
+ $X2=0 $Y2=0
cc_223 N_A_27_468#_M1003_g N_A_357_365#_c_347_n 0.0121848f $X=2.76 $Y=0.835
+ $X2=0 $Y2=0
cc_224 N_A_27_468#_c_238_n N_A_357_365#_c_347_n 0.0245023f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_225 N_A_27_468#_c_239_n N_A_357_365#_c_347_n 0.00123144f $X=2.67 $Y=1.57
+ $X2=0 $Y2=0
cc_226 N_A_27_468#_M1003_g N_A_357_365#_c_349_n 0.0104246f $X=2.76 $Y=0.835
+ $X2=0 $Y2=0
cc_227 N_A_27_468#_M1003_g N_A_357_365#_c_353_n 0.00198306f $X=2.76 $Y=0.835
+ $X2=0 $Y2=0
cc_228 N_A_27_468#_M1003_g N_A_357_365#_c_354_n 0.00164614f $X=2.76 $Y=0.835
+ $X2=0 $Y2=0
cc_229 N_A_27_468#_c_236_n N_A_357_365#_c_354_n 0.00114651f $X=2.67 $Y=1.91
+ $X2=0 $Y2=0
cc_230 N_A_27_468#_c_238_n N_A_357_365#_c_354_n 0.0432786f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_231 N_A_27_468#_c_239_n N_A_357_365#_c_354_n 0.00465147f $X=2.67 $Y=1.57
+ $X2=0 $Y2=0
cc_232 N_A_27_468#_c_236_n N_A_357_365#_c_360_n 0.0376618f $X=2.67 $Y=1.91 $X2=0
+ $Y2=0
cc_233 N_A_27_468#_c_238_n N_A_357_365#_c_360_n 0.00237622f $X=2.67 $Y=1.57
+ $X2=0 $Y2=0
cc_234 N_A_27_468#_c_246_n N_A_250_70#_M1005_d 0.00321487f $X=1.675 $Y=2.915
+ $X2=0 $Y2=0
cc_235 N_A_27_468#_M1003_g N_A_250_70#_c_460_n 0.0089911f $X=2.76 $Y=0.835 $X2=0
+ $Y2=0
cc_236 N_A_27_468#_M1003_g N_A_250_70#_M1017_g 0.0206778f $X=2.76 $Y=0.835 $X2=0
+ $Y2=0
cc_237 N_A_27_468#_M1010_g N_A_250_70#_M1002_g 0.0158123f $X=2.76 $Y=2.555 $X2=0
+ $Y2=0
cc_238 N_A_27_468#_c_236_n N_A_250_70#_M1002_g 0.0202042f $X=2.67 $Y=1.91 $X2=0
+ $Y2=0
cc_239 N_A_27_468#_c_246_n N_A_250_70#_M1002_g 0.00395685f $X=1.675 $Y=2.915
+ $X2=0 $Y2=0
cc_240 N_A_27_468#_c_248_n N_A_250_70#_M1002_g 0.0113396f $X=1.842 $Y=2.83 $X2=0
+ $Y2=0
cc_241 N_A_27_468#_c_273_p N_A_250_70#_M1002_g 0.0177646f $X=2.505 $Y=2.36 $X2=0
+ $Y2=0
cc_242 N_A_27_468#_c_238_n N_A_250_70#_M1002_g 0.00419199f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_243 N_A_27_468#_M1003_g N_A_250_70#_M1024_g 0.0314158f $X=2.76 $Y=0.835 $X2=0
+ $Y2=0
cc_244 N_A_27_468#_c_238_n N_A_250_70#_c_465_n 5.20602e-19 $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_245 N_A_27_468#_c_239_n N_A_250_70#_c_465_n 0.0314158f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_246 N_A_27_468#_c_249_n N_A_250_70#_c_467_n 0.00171197f $X=2.01 $Y=2.36 $X2=0
+ $Y2=0
cc_247 N_A_27_468#_c_238_n N_A_250_70#_c_469_n 0.00231268f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_248 N_A_27_468#_c_239_n N_A_250_70#_c_469_n 0.0202042f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_249 N_A_27_468#_c_245_n N_A_250_70#_c_478_n 0.00790237f $X=0.955 $Y=2.405
+ $X2=0 $Y2=0
cc_250 N_A_27_468#_c_246_n N_A_250_70#_c_478_n 0.015221f $X=1.675 $Y=2.915 $X2=0
+ $Y2=0
cc_251 N_A_27_468#_c_248_n N_A_250_70#_c_478_n 0.0169892f $X=1.842 $Y=2.83 $X2=0
+ $Y2=0
cc_252 N_A_27_468#_c_249_n N_A_250_70#_c_478_n 0.0144216f $X=2.01 $Y=2.36 $X2=0
+ $Y2=0
cc_253 N_A_27_468#_c_249_n N_A_250_70#_c_471_n 0.00217628f $X=2.01 $Y=2.36 $X2=0
+ $Y2=0
cc_254 N_A_27_468#_M1010_g N_A_639_125#_c_759_n 0.00179067f $X=2.76 $Y=2.555
+ $X2=0 $Y2=0
cc_255 N_A_27_468#_c_273_p N_A_639_125#_c_759_n 0.00776834f $X=2.505 $Y=2.36
+ $X2=0 $Y2=0
cc_256 N_A_27_468#_c_238_n N_A_639_125#_c_759_n 0.0012738f $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_257 N_A_27_468#_c_245_n N_VPWR_M1022_d 0.00684084f $X=0.955 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_258 N_A_27_468#_c_257_n N_VPWR_M1022_d 0.00404186f $X=1.04 $Y=2.83 $X2=-0.19
+ $Y2=-0.245
cc_259 N_A_27_468#_c_247_n N_VPWR_M1022_d 0.00143095f $X=1.125 $Y=2.915
+ $X2=-0.19 $Y2=-0.245
cc_260 N_A_27_468#_c_273_p N_VPWR_M1002_d 0.00903518f $X=2.505 $Y=2.36 $X2=0
+ $Y2=0
cc_261 N_A_27_468#_c_238_n N_VPWR_M1002_d 5.04244e-19 $X=2.67 $Y=1.57 $X2=0
+ $Y2=0
cc_262 N_A_27_468#_c_245_n N_VPWR_c_881_n 0.015086f $X=0.955 $Y=2.405 $X2=0
+ $Y2=0
cc_263 N_A_27_468#_c_257_n N_VPWR_c_881_n 0.0126784f $X=1.04 $Y=2.83 $X2=0 $Y2=0
cc_264 N_A_27_468#_c_247_n N_VPWR_c_881_n 0.0142637f $X=1.125 $Y=2.915 $X2=0
+ $Y2=0
cc_265 N_A_27_468#_c_251_n N_VPWR_c_881_n 0.0129931f $X=0.26 $Y=2.485 $X2=0
+ $Y2=0
cc_266 N_A_27_468#_M1010_g N_VPWR_c_882_n 0.00367204f $X=2.76 $Y=2.555 $X2=0
+ $Y2=0
cc_267 N_A_27_468#_c_243_n N_VPWR_c_882_n 4.97572e-19 $X=2.67 $Y=2.075 $X2=0
+ $Y2=0
cc_268 N_A_27_468#_c_246_n N_VPWR_c_882_n 0.00843167f $X=1.675 $Y=2.915 $X2=0
+ $Y2=0
cc_269 N_A_27_468#_c_273_p N_VPWR_c_882_n 0.0234562f $X=2.505 $Y=2.36 $X2=0
+ $Y2=0
cc_270 N_A_27_468#_M1010_g N_VPWR_c_889_n 0.00517164f $X=2.76 $Y=2.555 $X2=0
+ $Y2=0
cc_271 N_A_27_468#_c_251_n N_VPWR_c_891_n 0.0129995f $X=0.26 $Y=2.485 $X2=0
+ $Y2=0
cc_272 N_A_27_468#_c_246_n N_VPWR_c_892_n 0.0399938f $X=1.675 $Y=2.915 $X2=0
+ $Y2=0
cc_273 N_A_27_468#_c_247_n N_VPWR_c_892_n 0.00814802f $X=1.125 $Y=2.915 $X2=0
+ $Y2=0
cc_274 N_A_27_468#_M1010_g N_VPWR_c_880_n 0.00519032f $X=2.76 $Y=2.555 $X2=0
+ $Y2=0
cc_275 N_A_27_468#_c_245_n N_VPWR_c_880_n 0.0115759f $X=0.955 $Y=2.405 $X2=0
+ $Y2=0
cc_276 N_A_27_468#_c_246_n N_VPWR_c_880_n 0.0316348f $X=1.675 $Y=2.915 $X2=0
+ $Y2=0
cc_277 N_A_27_468#_c_247_n N_VPWR_c_880_n 0.00622816f $X=1.125 $Y=2.915 $X2=0
+ $Y2=0
cc_278 N_A_27_468#_c_251_n N_VPWR_c_880_n 0.0100156f $X=0.26 $Y=2.485 $X2=0
+ $Y2=0
cc_279 N_A_27_468#_c_240_n N_VGND_c_1048_n 0.0135511f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_280 N_A_27_468#_M1003_g N_VGND_c_1049_n 0.00348057f $X=2.76 $Y=0.835 $X2=0
+ $Y2=0
cc_281 N_A_27_468#_c_240_n N_VGND_c_1055_n 0.0243469f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_282 N_A_27_468#_M1003_g N_VGND_c_1066_n 8.54987e-19 $X=2.76 $Y=0.835 $X2=0
+ $Y2=0
cc_283 N_A_27_468#_c_240_n N_VGND_c_1066_n 0.01937f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_284 N_A_357_365#_c_345_n N_A_250_70#_c_459_n 0.00313006f $X=2.005 $Y=0.9
+ $X2=0 $Y2=0
cc_285 N_A_357_365#_c_348_n N_A_250_70#_c_459_n 0.00192424f $X=2.27 $Y=1.14
+ $X2=0 $Y2=0
cc_286 N_A_357_365#_c_345_n N_A_250_70#_c_460_n 0.00342288f $X=2.005 $Y=0.9
+ $X2=0 $Y2=0
cc_287 N_A_357_365#_c_350_n N_A_250_70#_c_460_n 0.00449971f $X=2.99 $Y=0.375
+ $X2=0 $Y2=0
cc_288 N_A_357_365#_c_352_n N_A_250_70#_c_460_n 0.0218994f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_289 N_A_357_365#_c_345_n N_A_250_70#_M1017_g 2.50028e-19 $X=2.005 $Y=0.9
+ $X2=0 $Y2=0
cc_290 N_A_357_365#_c_346_n N_A_250_70#_M1017_g 0.00437748f $X=2.185 $Y=1.825
+ $X2=0 $Y2=0
cc_291 N_A_357_365#_c_347_n N_A_250_70#_M1017_g 0.00463491f $X=2.82 $Y=1.14
+ $X2=0 $Y2=0
cc_292 N_A_357_365#_c_348_n N_A_250_70#_M1017_g 0.00966556f $X=2.27 $Y=1.14
+ $X2=0 $Y2=0
cc_293 N_A_357_365#_c_349_n N_A_250_70#_M1017_g 7.65731e-19 $X=2.905 $Y=1.055
+ $X2=0 $Y2=0
cc_294 N_A_357_365#_c_357_n N_A_250_70#_M1002_g 0.0128592f $X=2.1 $Y=1.965 $X2=0
+ $Y2=0
cc_295 N_A_357_365#_c_346_n N_A_250_70#_M1002_g 0.00554646f $X=2.185 $Y=1.825
+ $X2=0 $Y2=0
cc_296 N_A_357_365#_c_349_n N_A_250_70#_M1024_g 0.00440623f $X=2.905 $Y=1.055
+ $X2=0 $Y2=0
cc_297 N_A_357_365#_c_351_n N_A_250_70#_M1024_g 0.0148264f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_298 N_A_357_365#_c_353_n N_A_250_70#_M1024_g 0.00973137f $X=3.21 $Y=1.225
+ $X2=0 $Y2=0
cc_299 N_A_357_365#_c_354_n N_A_250_70#_M1024_g 0.00763076f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_300 N_A_357_365#_c_355_n N_A_250_70#_M1024_g 0.0131527f $X=3.57 $Y=0.515
+ $X2=0 $Y2=0
cc_301 N_A_357_365#_c_353_n N_A_250_70#_c_464_n 9.17726e-19 $X=3.21 $Y=1.225
+ $X2=0 $Y2=0
cc_302 N_A_357_365#_c_354_n N_A_250_70#_c_464_n 0.00927475f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_303 N_A_357_365#_c_355_n N_A_250_70#_c_464_n 0.0101968f $X=3.57 $Y=0.515
+ $X2=0 $Y2=0
cc_304 N_A_357_365#_c_354_n N_A_250_70#_c_465_n 0.00440067f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_305 N_A_357_365#_c_360_n N_A_250_70#_c_465_n 0.0214353f $X=3.21 $Y=1.91 $X2=0
+ $Y2=0
cc_306 N_A_357_365#_c_354_n N_A_250_70#_c_466_n 0.00100968f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_307 N_A_357_365#_M1013_g N_A_250_70#_M1020_g 0.0112112f $X=3.12 $Y=2.555
+ $X2=0 $Y2=0
cc_308 N_A_357_365#_c_354_n N_A_250_70#_M1020_g 7.76758e-19 $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_309 N_A_357_365#_c_360_n N_A_250_70#_M1020_g 0.0199364f $X=3.21 $Y=1.91 $X2=0
+ $Y2=0
cc_310 N_A_357_365#_c_357_n N_A_250_70#_c_468_n 0.00943647f $X=2.1 $Y=1.965
+ $X2=0 $Y2=0
cc_311 N_A_357_365#_c_346_n N_A_250_70#_c_468_n 0.00764743f $X=2.185 $Y=1.825
+ $X2=0 $Y2=0
cc_312 N_A_357_365#_c_348_n N_A_250_70#_c_468_n 0.00443992f $X=2.27 $Y=1.14
+ $X2=0 $Y2=0
cc_313 N_A_357_365#_c_346_n N_A_250_70#_c_469_n 0.00663031f $X=2.185 $Y=1.825
+ $X2=0 $Y2=0
cc_314 N_A_357_365#_c_345_n N_A_250_70#_c_470_n 0.0130273f $X=2.005 $Y=0.9 $X2=0
+ $Y2=0
cc_315 N_A_357_365#_c_346_n N_A_250_70#_c_470_n 0.00504148f $X=2.185 $Y=1.825
+ $X2=0 $Y2=0
cc_316 N_A_357_365#_c_348_n N_A_250_70#_c_470_n 0.0078194f $X=2.27 $Y=1.14 $X2=0
+ $Y2=0
cc_317 N_A_357_365#_c_357_n N_A_250_70#_c_478_n 0.0183166f $X=2.1 $Y=1.965 $X2=0
+ $Y2=0
cc_318 N_A_357_365#_c_346_n N_A_250_70#_c_478_n 0.00541304f $X=2.185 $Y=1.825
+ $X2=0 $Y2=0
cc_319 N_A_357_365#_c_357_n N_A_250_70#_c_471_n 0.0132375f $X=2.1 $Y=1.965 $X2=0
+ $Y2=0
cc_320 N_A_357_365#_c_346_n N_A_250_70#_c_471_n 0.0186352f $X=2.185 $Y=1.825
+ $X2=0 $Y2=0
cc_321 N_A_357_365#_c_348_n N_A_250_70#_c_471_n 0.00147608f $X=2.27 $Y=1.14
+ $X2=0 $Y2=0
cc_322 N_A_357_365#_c_352_n N_A_789_99#_M1004_g 0.00129738f $X=3.57 $Y=0.35
+ $X2=0 $Y2=0
cc_323 N_A_357_365#_c_353_n N_A_789_99#_M1004_g 2.09531e-19 $X=3.21 $Y=1.225
+ $X2=0 $Y2=0
cc_324 N_A_357_365#_c_355_n N_A_789_99#_M1004_g 0.0237861f $X=3.57 $Y=0.515
+ $X2=0 $Y2=0
cc_325 N_A_357_365#_c_351_n N_A_639_125#_c_764_n 0.0341169f $X=3.57 $Y=0.35
+ $X2=0 $Y2=0
cc_326 N_A_357_365#_c_352_n N_A_639_125#_c_764_n 0.00368391f $X=3.57 $Y=0.35
+ $X2=0 $Y2=0
cc_327 N_A_357_365#_c_353_n N_A_639_125#_c_764_n 0.0131135f $X=3.21 $Y=1.225
+ $X2=0 $Y2=0
cc_328 N_A_357_365#_c_355_n N_A_639_125#_c_764_n 0.00786284f $X=3.57 $Y=0.515
+ $X2=0 $Y2=0
cc_329 N_A_357_365#_c_349_n N_A_639_125#_c_768_n 0.00233108f $X=2.905 $Y=1.055
+ $X2=0 $Y2=0
cc_330 N_A_357_365#_c_353_n N_A_639_125#_c_768_n 6.94436e-19 $X=3.21 $Y=1.225
+ $X2=0 $Y2=0
cc_331 N_A_357_365#_c_355_n N_A_639_125#_c_768_n 0.00501052f $X=3.57 $Y=0.515
+ $X2=0 $Y2=0
cc_332 N_A_357_365#_c_351_n N_A_639_125#_c_754_n 2.78145e-19 $X=3.57 $Y=0.35
+ $X2=0 $Y2=0
cc_333 N_A_357_365#_M1013_g N_A_639_125#_c_759_n 0.0140939f $X=3.12 $Y=2.555
+ $X2=0 $Y2=0
cc_334 N_A_357_365#_c_354_n N_A_639_125#_c_759_n 0.0133637f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_335 N_A_357_365#_c_360_n N_A_639_125#_c_759_n 0.0012342f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_336 N_A_357_365#_M1013_g N_A_639_125#_c_756_n 0.00285432f $X=3.12 $Y=2.555
+ $X2=0 $Y2=0
cc_337 N_A_357_365#_c_354_n N_A_639_125#_c_756_n 0.0642867f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_338 N_A_357_365#_c_360_n N_A_639_125#_c_756_n 0.00177198f $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_339 N_A_357_365#_c_353_n N_A_639_125#_c_757_n 0.014397f $X=3.21 $Y=1.225
+ $X2=0 $Y2=0
cc_340 N_A_357_365#_c_354_n N_A_639_125#_c_757_n 8.84571e-19 $X=3.21 $Y=1.91
+ $X2=0 $Y2=0
cc_341 N_A_357_365#_c_355_n N_A_639_125#_c_757_n 0.00369519f $X=3.57 $Y=0.515
+ $X2=0 $Y2=0
cc_342 N_A_357_365#_M1013_g N_VPWR_c_889_n 0.00513466f $X=3.12 $Y=2.555 $X2=0
+ $Y2=0
cc_343 N_A_357_365#_M1013_g N_VPWR_c_880_n 0.00519032f $X=3.12 $Y=2.555 $X2=0
+ $Y2=0
cc_344 N_A_357_365#_c_347_n N_VGND_c_1049_n 0.0234958f $X=2.82 $Y=1.14 $X2=0
+ $Y2=0
cc_345 N_A_357_365#_c_349_n N_VGND_c_1049_n 0.0249893f $X=2.905 $Y=1.055 $X2=0
+ $Y2=0
cc_346 N_A_357_365#_c_350_n N_VGND_c_1049_n 0.0189285f $X=2.99 $Y=0.375 $X2=0
+ $Y2=0
cc_347 N_A_357_365#_c_351_n N_VGND_c_1050_n 0.0120133f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_348 N_A_357_365#_c_352_n N_VGND_c_1050_n 0.00337756f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_349 N_A_357_365#_c_355_n N_VGND_c_1050_n 9.36255e-19 $X=3.57 $Y=0.515 $X2=0
+ $Y2=0
cc_350 N_A_357_365#_c_345_n N_VGND_c_1057_n 0.00293469f $X=2.005 $Y=0.9 $X2=0
+ $Y2=0
cc_351 N_A_357_365#_c_350_n N_VGND_c_1059_n 0.0115893f $X=2.99 $Y=0.375 $X2=0
+ $Y2=0
cc_352 N_A_357_365#_c_351_n N_VGND_c_1059_n 0.0476644f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_353 N_A_357_365#_c_352_n N_VGND_c_1059_n 0.00647615f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_354 N_A_357_365#_c_345_n N_VGND_c_1066_n 0.00485186f $X=2.005 $Y=0.9 $X2=0
+ $Y2=0
cc_355 N_A_357_365#_c_350_n N_VGND_c_1066_n 0.00583135f $X=2.99 $Y=0.375 $X2=0
+ $Y2=0
cc_356 N_A_357_365#_c_351_n N_VGND_c_1066_n 0.0257792f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_357 N_A_357_365#_c_352_n N_VGND_c_1066_n 0.00941423f $X=3.57 $Y=0.35 $X2=0
+ $Y2=0
cc_358 N_A_250_70#_c_466_n N_A_789_99#_c_578_n 0.0456558f $X=3.665 $Y=1.685
+ $X2=0 $Y2=0
cc_359 N_A_250_70#_M1020_g N_A_789_99#_c_598_n 0.036136f $X=3.665 $Y=2.445 $X2=0
+ $Y2=0
cc_360 N_A_250_70#_c_466_n N_A_789_99#_c_585_n 0.00286462f $X=3.665 $Y=1.685
+ $X2=0 $Y2=0
cc_361 N_A_250_70#_M1020_g N_A_789_99#_c_608_n 5.17944e-19 $X=3.665 $Y=2.445
+ $X2=0 $Y2=0
cc_362 N_A_250_70#_M1024_g N_A_639_125#_c_764_n 0.00289485f $X=3.12 $Y=0.835
+ $X2=0 $Y2=0
cc_363 N_A_250_70#_c_464_n N_A_639_125#_c_764_n 0.00202333f $X=3.585 $Y=1.46
+ $X2=0 $Y2=0
cc_364 N_A_250_70#_M1024_g N_A_639_125#_c_768_n 3.65619e-19 $X=3.12 $Y=0.835
+ $X2=0 $Y2=0
cc_365 N_A_250_70#_c_466_n N_A_639_125#_c_754_n 5.87044e-19 $X=3.665 $Y=1.685
+ $X2=0 $Y2=0
cc_366 N_A_250_70#_M1020_g N_A_639_125#_c_759_n 0.017902f $X=3.665 $Y=2.445
+ $X2=0 $Y2=0
cc_367 N_A_250_70#_M1024_g N_A_639_125#_c_756_n 6.96382e-19 $X=3.12 $Y=0.835
+ $X2=0 $Y2=0
cc_368 N_A_250_70#_c_464_n N_A_639_125#_c_756_n 0.00385089f $X=3.585 $Y=1.46
+ $X2=0 $Y2=0
cc_369 N_A_250_70#_c_466_n N_A_639_125#_c_756_n 0.0110063f $X=3.665 $Y=1.685
+ $X2=0 $Y2=0
cc_370 N_A_250_70#_M1020_g N_A_639_125#_c_756_n 0.0132171f $X=3.665 $Y=2.445
+ $X2=0 $Y2=0
cc_371 N_A_250_70#_M1024_g N_A_639_125#_c_757_n 4.03666e-19 $X=3.12 $Y=0.835
+ $X2=0 $Y2=0
cc_372 N_A_250_70#_M1002_g N_VPWR_c_882_n 0.00161341f $X=2.22 $Y=2.555 $X2=0
+ $Y2=0
cc_373 N_A_250_70#_M1020_g N_VPWR_c_889_n 9.55248e-19 $X=3.665 $Y=2.445 $X2=0
+ $Y2=0
cc_374 N_A_250_70#_M1002_g N_VPWR_c_892_n 0.00517164f $X=2.22 $Y=2.555 $X2=0
+ $Y2=0
cc_375 N_A_250_70#_M1002_g N_VPWR_c_880_n 0.00519032f $X=2.22 $Y=2.555 $X2=0
+ $Y2=0
cc_376 N_A_250_70#_M1020_g N_VPWR_c_880_n 4.8622e-19 $X=3.665 $Y=2.445 $X2=0
+ $Y2=0
cc_377 N_A_250_70#_c_461_n N_VGND_c_1048_n 0.00288221f $X=1.74 $Y=0.18 $X2=0
+ $Y2=0
cc_378 N_A_250_70#_c_470_n N_VGND_c_1048_n 0.0134903f $X=1.39 $Y=0.495 $X2=0
+ $Y2=0
cc_379 N_A_250_70#_c_459_n N_VGND_c_1049_n 0.00483978f $X=1.665 $Y=1.325 $X2=0
+ $Y2=0
cc_380 N_A_250_70#_c_460_n N_VGND_c_1049_n 0.0257163f $X=3.045 $Y=0.18 $X2=0
+ $Y2=0
cc_381 N_A_250_70#_M1017_g N_VGND_c_1049_n 0.00746159f $X=2.22 $Y=0.835 $X2=0
+ $Y2=0
cc_382 N_A_250_70#_M1024_g N_VGND_c_1049_n 0.00108545f $X=3.12 $Y=0.835 $X2=0
+ $Y2=0
cc_383 N_A_250_70#_c_461_n N_VGND_c_1057_n 0.0235357f $X=1.74 $Y=0.18 $X2=0
+ $Y2=0
cc_384 N_A_250_70#_c_470_n N_VGND_c_1057_n 0.00960412f $X=1.39 $Y=0.495 $X2=0
+ $Y2=0
cc_385 N_A_250_70#_c_460_n N_VGND_c_1059_n 0.0154621f $X=3.045 $Y=0.18 $X2=0
+ $Y2=0
cc_386 N_A_250_70#_c_460_n N_VGND_c_1066_n 0.0401241f $X=3.045 $Y=0.18 $X2=0
+ $Y2=0
cc_387 N_A_250_70#_c_461_n N_VGND_c_1066_n 0.0113745f $X=1.74 $Y=0.18 $X2=0
+ $Y2=0
cc_388 N_A_250_70#_M1017_g N_VGND_c_1066_n 9.24653e-19 $X=2.22 $Y=0.835 $X2=0
+ $Y2=0
cc_389 N_A_250_70#_c_470_n N_VGND_c_1066_n 0.00739956f $X=1.39 $Y=0.495 $X2=0
+ $Y2=0
cc_390 N_A_789_99#_c_586_n N_A_639_125#_c_750_n 0.00817817f $X=4.755 $Y=0.42
+ $X2=0 $Y2=0
cc_391 N_A_789_99#_c_587_n N_A_639_125#_c_750_n 0.0189547f $X=5.115 $Y=0.955
+ $X2=0 $Y2=0
cc_392 N_A_789_99#_c_578_n N_A_639_125#_M1019_g 0.00893987f $X=4.02 $Y=1.175
+ $X2=0 $Y2=0
cc_393 N_A_789_99#_c_585_n N_A_639_125#_M1019_g 0.00678987f $X=4.115 $Y=1.57
+ $X2=0 $Y2=0
cc_394 N_A_789_99#_c_613_p N_A_639_125#_M1019_g 0.0133814f $X=5.09 $Y=2.385
+ $X2=0 $Y2=0
cc_395 N_A_789_99#_c_578_n N_A_639_125#_c_752_n 0.0130664f $X=4.02 $Y=1.175
+ $X2=0 $Y2=0
cc_396 N_A_789_99#_c_585_n N_A_639_125#_c_752_n 4.45052e-19 $X=4.115 $Y=1.57
+ $X2=0 $Y2=0
cc_397 N_A_789_99#_c_587_n N_A_639_125#_c_752_n 0.00450116f $X=5.115 $Y=0.955
+ $X2=0 $Y2=0
cc_398 N_A_789_99#_M1004_g N_A_639_125#_c_764_n 0.00184053f $X=4.02 $Y=0.835
+ $X2=0 $Y2=0
cc_399 N_A_789_99#_M1004_g N_A_639_125#_c_768_n 0.00346297f $X=4.02 $Y=0.835
+ $X2=0 $Y2=0
cc_400 N_A_789_99#_M1018_s N_A_639_125#_c_754_n 0.00170668f $X=4.63 $Y=0.235
+ $X2=0 $Y2=0
cc_401 N_A_789_99#_c_578_n N_A_639_125#_c_754_n 0.00736291f $X=4.02 $Y=1.175
+ $X2=0 $Y2=0
cc_402 N_A_789_99#_M1004_g N_A_639_125#_c_754_n 0.0111436f $X=4.02 $Y=0.835
+ $X2=0 $Y2=0
cc_403 N_A_789_99#_c_585_n N_A_639_125#_c_754_n 0.0255615f $X=4.115 $Y=1.57
+ $X2=0 $Y2=0
cc_404 N_A_789_99#_c_587_n N_A_639_125#_c_754_n 0.0162475f $X=5.115 $Y=0.955
+ $X2=0 $Y2=0
cc_405 N_A_789_99#_c_578_n N_A_639_125#_c_755_n 0.00140552f $X=4.02 $Y=1.175
+ $X2=0 $Y2=0
cc_406 N_A_789_99#_c_585_n N_A_639_125#_c_755_n 0.00603611f $X=4.115 $Y=1.57
+ $X2=0 $Y2=0
cc_407 N_A_789_99#_M1008_g N_A_639_125#_c_759_n 0.00221633f $X=4.025 $Y=2.445
+ $X2=0 $Y2=0
cc_408 N_A_789_99#_c_598_n N_A_639_125#_c_759_n 0.00154238f $X=4.115 $Y=2.075
+ $X2=0 $Y2=0
cc_409 N_A_789_99#_c_608_n N_A_639_125#_c_759_n 0.0112256f $X=4.28 $Y=2.385
+ $X2=0 $Y2=0
cc_410 N_A_789_99#_c_578_n N_A_639_125#_c_756_n 0.00650992f $X=4.02 $Y=1.175
+ $X2=0 $Y2=0
cc_411 N_A_789_99#_c_585_n N_A_639_125#_c_756_n 0.0513966f $X=4.115 $Y=1.57
+ $X2=0 $Y2=0
cc_412 N_A_789_99#_M1011_g N_RESET_B_M1009_g 0.0261492f $X=5.905 $Y=0.655 $X2=0
+ $Y2=0
cc_413 N_A_789_99#_c_586_n N_RESET_B_M1009_g 0.00137743f $X=4.755 $Y=0.42 $X2=0
+ $Y2=0
cc_414 N_A_789_99#_c_633_p N_RESET_B_M1009_g 0.0152346f $X=5.685 $Y=0.955 $X2=0
+ $Y2=0
cc_415 N_A_789_99#_c_587_n N_RESET_B_M1009_g 0.00376871f $X=5.115 $Y=0.955 $X2=0
+ $Y2=0
cc_416 N_A_789_99#_c_588_n N_RESET_B_M1009_g 0.00326623f $X=5.77 $Y=1.425 $X2=0
+ $Y2=0
cc_417 N_A_789_99#_c_636_p N_RESET_B_M1006_g 0.0103491f $X=5.685 $Y=2.385 $X2=0
+ $Y2=0
cc_418 N_A_789_99#_c_589_n N_RESET_B_M1006_g 0.00505947f $X=5.77 $Y=2.3 $X2=0
+ $Y2=0
cc_419 N_A_789_99#_c_590_n N_RESET_B_M1006_g 2.0934e-19 $X=5.77 $Y=1.51 $X2=0
+ $Y2=0
cc_420 N_A_789_99#_c_591_n N_RESET_B_M1006_g 0.0432689f $X=7.195 $Y=1.51 $X2=0
+ $Y2=0
cc_421 N_A_789_99#_M1019_d RESET_B 0.001837f $X=5.045 $Y=1.835 $X2=0 $Y2=0
cc_422 N_A_789_99#_c_578_n RESET_B 0.00218717f $X=4.02 $Y=1.175 $X2=0 $Y2=0
cc_423 N_A_789_99#_c_585_n RESET_B 0.0155964f $X=4.115 $Y=1.57 $X2=0 $Y2=0
cc_424 N_A_789_99#_c_613_p RESET_B 0.0075073f $X=5.09 $Y=2.385 $X2=0 $Y2=0
cc_425 N_A_789_99#_c_633_p RESET_B 0.027437f $X=5.685 $Y=0.955 $X2=0 $Y2=0
cc_426 N_A_789_99#_c_587_n RESET_B 0.0117197f $X=5.115 $Y=0.955 $X2=0 $Y2=0
cc_427 N_A_789_99#_c_636_p RESET_B 0.0113922f $X=5.685 $Y=2.385 $X2=0 $Y2=0
cc_428 N_A_789_99#_c_588_n RESET_B 0.0168226f $X=5.77 $Y=1.425 $X2=0 $Y2=0
cc_429 N_A_789_99#_c_589_n RESET_B 0.0305142f $X=5.77 $Y=2.3 $X2=0 $Y2=0
cc_430 N_A_789_99#_c_649_p RESET_B 0.0149669f $X=5.185 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A_789_99#_c_590_n RESET_B 0.0151373f $X=5.77 $Y=1.51 $X2=0 $Y2=0
cc_432 N_A_789_99#_c_591_n RESET_B 0.00125685f $X=7.195 $Y=1.51 $X2=0 $Y2=0
cc_433 N_A_789_99#_M1011_g N_RESET_B_c_837_n 0.00679965f $X=5.905 $Y=0.655 $X2=0
+ $Y2=0
cc_434 N_A_789_99#_c_633_p N_RESET_B_c_837_n 0.00330464f $X=5.685 $Y=0.955 $X2=0
+ $Y2=0
cc_435 N_A_789_99#_c_588_n N_RESET_B_c_837_n 0.0014059f $X=5.77 $Y=1.425 $X2=0
+ $Y2=0
cc_436 N_A_789_99#_c_590_n N_RESET_B_c_837_n 8.56548e-19 $X=5.77 $Y=1.51 $X2=0
+ $Y2=0
cc_437 N_A_789_99#_c_591_n N_RESET_B_c_837_n 0.0104992f $X=7.195 $Y=1.51 $X2=0
+ $Y2=0
cc_438 N_A_789_99#_c_585_n N_VPWR_M1008_d 0.00117668f $X=4.115 $Y=1.57 $X2=0
+ $Y2=0
cc_439 N_A_789_99#_c_613_p N_VPWR_M1008_d 0.0342201f $X=5.09 $Y=2.385 $X2=0
+ $Y2=0
cc_440 N_A_789_99#_c_608_n N_VPWR_M1008_d 0.00294652f $X=4.28 $Y=2.385 $X2=0
+ $Y2=0
cc_441 N_A_789_99#_c_636_p N_VPWR_M1006_d 0.00823753f $X=5.685 $Y=2.385 $X2=0
+ $Y2=0
cc_442 N_A_789_99#_c_589_n N_VPWR_M1006_d 0.00452115f $X=5.77 $Y=2.3 $X2=0 $Y2=0
cc_443 N_A_789_99#_M1008_g N_VPWR_c_883_n 0.00384439f $X=4.025 $Y=2.445 $X2=0
+ $Y2=0
cc_444 N_A_789_99#_c_613_p N_VPWR_c_883_n 0.0214369f $X=5.09 $Y=2.385 $X2=0
+ $Y2=0
cc_445 N_A_789_99#_c_649_p N_VPWR_c_884_n 0.0135169f $X=5.185 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_A_789_99#_M1007_g N_VPWR_c_885_n 0.0024778f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_789_99#_c_636_p N_VPWR_c_885_n 0.0189931f $X=5.685 $Y=2.385 $X2=0
+ $Y2=0
cc_448 N_A_789_99#_M1007_g N_VPWR_c_886_n 7.29879e-19 $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A_789_99#_M1014_g N_VPWR_c_886_n 0.0142382f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_789_99#_M1015_g N_VPWR_c_886_n 0.0141179f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_451 N_A_789_99#_M1025_g N_VPWR_c_886_n 7.24342e-19 $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_452 N_A_789_99#_M1015_g N_VPWR_c_888_n 7.24342e-19 $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_453 N_A_789_99#_M1025_g N_VPWR_c_888_n 0.0151814f $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_454 N_A_789_99#_M1008_g N_VPWR_c_889_n 0.00389919f $X=4.025 $Y=2.445 $X2=0
+ $Y2=0
cc_455 N_A_789_99#_M1007_g N_VPWR_c_893_n 0.00585385f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A_789_99#_M1014_g N_VPWR_c_893_n 0.00486043f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_457 N_A_789_99#_M1015_g N_VPWR_c_894_n 0.00486043f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_458 N_A_789_99#_M1025_g N_VPWR_c_894_n 0.00486043f $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_459 N_A_789_99#_M1019_d N_VPWR_c_880_n 0.00262154f $X=5.045 $Y=1.835 $X2=0
+ $Y2=0
cc_460 N_A_789_99#_M1008_g N_VPWR_c_880_n 0.00455831f $X=4.025 $Y=2.445 $X2=0
+ $Y2=0
cc_461 N_A_789_99#_M1007_g N_VPWR_c_880_n 0.00981659f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_462 N_A_789_99#_M1014_g N_VPWR_c_880_n 0.00827314f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_463 N_A_789_99#_M1015_g N_VPWR_c_880_n 0.00824727f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_464 N_A_789_99#_M1025_g N_VPWR_c_880_n 0.00824727f $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_465 N_A_789_99#_c_613_p N_VPWR_c_880_n 0.0163929f $X=5.09 $Y=2.385 $X2=0
+ $Y2=0
cc_466 N_A_789_99#_c_608_n N_VPWR_c_880_n 0.0121659f $X=4.28 $Y=2.385 $X2=0
+ $Y2=0
cc_467 N_A_789_99#_c_636_p N_VPWR_c_880_n 0.00715468f $X=5.685 $Y=2.385 $X2=0
+ $Y2=0
cc_468 N_A_789_99#_c_649_p N_VPWR_c_880_n 0.00847534f $X=5.185 $Y=2.465 $X2=0
+ $Y2=0
cc_469 N_A_789_99#_M1011_g N_Q_c_997_n 5.81897e-19 $X=5.905 $Y=0.655 $X2=0 $Y2=0
cc_470 N_A_789_99#_M1012_g N_Q_c_997_n 6.32385e-19 $X=6.335 $Y=0.655 $X2=0 $Y2=0
cc_471 N_A_789_99#_c_588_n N_Q_c_997_n 0.00179729f $X=5.77 $Y=1.425 $X2=0 $Y2=0
cc_472 N_A_789_99#_M1012_g N_Q_c_986_n 0.0138902f $X=6.335 $Y=0.655 $X2=0 $Y2=0
cc_473 N_A_789_99#_M1021_g N_Q_c_986_n 0.0142932f $X=6.765 $Y=0.655 $X2=0 $Y2=0
cc_474 N_A_789_99#_c_693_p N_Q_c_986_n 0.0467265f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_475 N_A_789_99#_c_591_n N_Q_c_986_n 0.00246472f $X=7.195 $Y=1.51 $X2=0 $Y2=0
cc_476 N_A_789_99#_M1011_g N_Q_c_987_n 0.0014023f $X=5.905 $Y=0.655 $X2=0 $Y2=0
cc_477 N_A_789_99#_c_588_n N_Q_c_987_n 0.013714f $X=5.77 $Y=1.425 $X2=0 $Y2=0
cc_478 N_A_789_99#_c_693_p N_Q_c_987_n 0.0153308f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_479 N_A_789_99#_c_591_n N_Q_c_987_n 0.00256759f $X=7.195 $Y=1.51 $X2=0 $Y2=0
cc_480 N_A_789_99#_M1014_g N_Q_c_992_n 0.0129257f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_481 N_A_789_99#_M1015_g N_Q_c_992_n 0.0130453f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_482 N_A_789_99#_c_693_p N_Q_c_992_n 0.0467265f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_483 N_A_789_99#_c_591_n N_Q_c_992_n 0.00246472f $X=7.195 $Y=1.51 $X2=0 $Y2=0
cc_484 N_A_789_99#_M1007_g N_Q_c_993_n 5.70797e-19 $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_485 N_A_789_99#_c_589_n N_Q_c_993_n 0.00900549f $X=5.77 $Y=2.3 $X2=0 $Y2=0
cc_486 N_A_789_99#_c_693_p N_Q_c_993_n 0.0153305f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_487 N_A_789_99#_c_591_n N_Q_c_993_n 0.00286738f $X=7.195 $Y=1.51 $X2=0 $Y2=0
cc_488 N_A_789_99#_M1021_g N_Q_c_1016_n 6.32385e-19 $X=6.765 $Y=0.655 $X2=0
+ $Y2=0
cc_489 N_A_789_99#_M1023_g N_Q_c_1016_n 7.21728e-19 $X=7.195 $Y=0.655 $X2=0
+ $Y2=0
cc_490 N_A_789_99#_M1023_g N_Q_c_988_n 0.0167803f $X=7.195 $Y=0.655 $X2=0 $Y2=0
cc_491 N_A_789_99#_c_693_p N_Q_c_988_n 0.0069096f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_492 N_A_789_99#_M1025_g N_Q_c_994_n 0.0155324f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_493 N_A_789_99#_c_693_p N_Q_c_994_n 0.0069096f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_494 N_A_789_99#_M1011_g N_Q_c_1022_n 0.00478077f $X=5.905 $Y=0.655 $X2=0
+ $Y2=0
cc_495 N_A_789_99#_c_693_p N_Q_c_989_n 0.0153308f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_496 N_A_789_99#_c_591_n N_Q_c_989_n 0.00256759f $X=7.195 $Y=1.51 $X2=0 $Y2=0
cc_497 N_A_789_99#_c_693_p N_Q_c_995_n 0.0153308f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_498 N_A_789_99#_c_591_n N_Q_c_995_n 0.00256759f $X=7.195 $Y=1.51 $X2=0 $Y2=0
cc_499 N_A_789_99#_M1023_g Q 0.0198116f $X=7.195 $Y=0.655 $X2=0 $Y2=0
cc_500 N_A_789_99#_c_693_p Q 0.0138072f $X=7.01 $Y=1.51 $X2=0 $Y2=0
cc_501 N_A_789_99#_c_633_p N_VGND_M1009_d 0.0089409f $X=5.685 $Y=0.955 $X2=0
+ $Y2=0
cc_502 N_A_789_99#_c_588_n N_VGND_M1009_d 4.29653e-19 $X=5.77 $Y=1.425 $X2=0
+ $Y2=0
cc_503 N_A_789_99#_M1004_g N_VGND_c_1050_n 0.00992362f $X=4.02 $Y=0.835 $X2=0
+ $Y2=0
cc_504 N_A_789_99#_c_586_n N_VGND_c_1050_n 0.0361528f $X=4.755 $Y=0.42 $X2=0
+ $Y2=0
cc_505 N_A_789_99#_c_587_n N_VGND_c_1050_n 0.0136615f $X=5.115 $Y=0.955 $X2=0
+ $Y2=0
cc_506 N_A_789_99#_M1011_g N_VGND_c_1051_n 0.00448009f $X=5.905 $Y=0.655 $X2=0
+ $Y2=0
cc_507 N_A_789_99#_c_633_p N_VGND_c_1051_n 0.0260407f $X=5.685 $Y=0.955 $X2=0
+ $Y2=0
cc_508 N_A_789_99#_M1011_g N_VGND_c_1052_n 4.81961e-19 $X=5.905 $Y=0.655 $X2=0
+ $Y2=0
cc_509 N_A_789_99#_M1012_g N_VGND_c_1052_n 0.0118875f $X=6.335 $Y=0.655 $X2=0
+ $Y2=0
cc_510 N_A_789_99#_M1021_g N_VGND_c_1052_n 0.0117077f $X=6.765 $Y=0.655 $X2=0
+ $Y2=0
cc_511 N_A_789_99#_M1023_g N_VGND_c_1052_n 6.36641e-19 $X=7.195 $Y=0.655 $X2=0
+ $Y2=0
cc_512 N_A_789_99#_M1021_g N_VGND_c_1054_n 6.36641e-19 $X=6.765 $Y=0.655 $X2=0
+ $Y2=0
cc_513 N_A_789_99#_M1023_g N_VGND_c_1054_n 0.0132658f $X=7.195 $Y=0.655 $X2=0
+ $Y2=0
cc_514 N_A_789_99#_M1004_g N_VGND_c_1059_n 0.00345209f $X=4.02 $Y=0.835 $X2=0
+ $Y2=0
cc_515 N_A_789_99#_c_586_n N_VGND_c_1060_n 0.0209621f $X=4.755 $Y=0.42 $X2=0
+ $Y2=0
cc_516 N_A_789_99#_c_587_n N_VGND_c_1060_n 0.00237032f $X=5.115 $Y=0.955 $X2=0
+ $Y2=0
cc_517 N_A_789_99#_M1011_g N_VGND_c_1061_n 0.0054895f $X=5.905 $Y=0.655 $X2=0
+ $Y2=0
cc_518 N_A_789_99#_M1012_g N_VGND_c_1061_n 0.00486043f $X=6.335 $Y=0.655 $X2=0
+ $Y2=0
cc_519 N_A_789_99#_M1021_g N_VGND_c_1062_n 0.00486043f $X=6.765 $Y=0.655 $X2=0
+ $Y2=0
cc_520 N_A_789_99#_M1023_g N_VGND_c_1062_n 0.00486043f $X=7.195 $Y=0.655 $X2=0
+ $Y2=0
cc_521 N_A_789_99#_M1018_s N_VGND_c_1066_n 0.00215158f $X=4.63 $Y=0.235 $X2=0
+ $Y2=0
cc_522 N_A_789_99#_M1004_g N_VGND_c_1066_n 0.00394323f $X=4.02 $Y=0.835 $X2=0
+ $Y2=0
cc_523 N_A_789_99#_M1011_g N_VGND_c_1066_n 0.0102611f $X=5.905 $Y=0.655 $X2=0
+ $Y2=0
cc_524 N_A_789_99#_M1012_g N_VGND_c_1066_n 0.00824727f $X=6.335 $Y=0.655 $X2=0
+ $Y2=0
cc_525 N_A_789_99#_M1021_g N_VGND_c_1066_n 0.00824727f $X=6.765 $Y=0.655 $X2=0
+ $Y2=0
cc_526 N_A_789_99#_M1023_g N_VGND_c_1066_n 0.00824727f $X=7.195 $Y=0.655 $X2=0
+ $Y2=0
cc_527 N_A_789_99#_c_586_n N_VGND_c_1066_n 0.0125487f $X=4.755 $Y=0.42 $X2=0
+ $Y2=0
cc_528 N_A_789_99#_c_587_n N_VGND_c_1066_n 0.00469036f $X=5.115 $Y=0.955 $X2=0
+ $Y2=0
cc_529 N_A_789_99#_c_633_p A_1009_47# 0.00400043f $X=5.685 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_530 N_A_789_99#_c_587_n A_1009_47# 0.00228619f $X=5.115 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_531 N_A_639_125#_c_750_n N_RESET_B_M1009_g 0.0443375f $X=4.97 $Y=1.185 $X2=0
+ $Y2=0
cc_532 N_A_639_125#_M1019_g N_RESET_B_M1006_g 0.041662f $X=4.97 $Y=2.465 $X2=0
+ $Y2=0
cc_533 N_A_639_125#_M1019_g RESET_B 0.0246926f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_534 N_A_639_125#_c_753_n RESET_B 0.0114184f $X=4.97 $Y=1.35 $X2=0 $Y2=0
cc_535 N_A_639_125#_c_754_n RESET_B 0.00207776f $X=4.525 $Y=1.15 $X2=0 $Y2=0
cc_536 N_A_639_125#_c_755_n RESET_B 0.0214546f $X=4.69 $Y=1.35 $X2=0 $Y2=0
cc_537 N_A_639_125#_c_753_n N_RESET_B_c_837_n 0.0443375f $X=4.97 $Y=1.35 $X2=0
+ $Y2=0
cc_538 N_A_639_125#_c_759_n N_VPWR_c_882_n 0.00442838f $X=3.4 $Y=2.38 $X2=0
+ $Y2=0
cc_539 N_A_639_125#_M1019_g N_VPWR_c_883_n 0.0126028f $X=4.97 $Y=2.465 $X2=0
+ $Y2=0
cc_540 N_A_639_125#_M1019_g N_VPWR_c_884_n 0.00486043f $X=4.97 $Y=2.465 $X2=0
+ $Y2=0
cc_541 N_A_639_125#_c_759_n N_VPWR_c_889_n 0.0171103f $X=3.4 $Y=2.38 $X2=0 $Y2=0
cc_542 N_A_639_125#_M1019_g N_VPWR_c_880_n 0.00460797f $X=4.97 $Y=2.465 $X2=0
+ $Y2=0
cc_543 N_A_639_125#_c_759_n N_VPWR_c_880_n 0.0184879f $X=3.4 $Y=2.38 $X2=0 $Y2=0
cc_544 N_A_639_125#_c_750_n N_VGND_c_1050_n 0.00230008f $X=4.97 $Y=1.185 $X2=0
+ $Y2=0
cc_545 N_A_639_125#_c_764_n N_VGND_c_1050_n 0.0103719f $X=3.545 $Y=0.775 $X2=0
+ $Y2=0
cc_546 N_A_639_125#_c_768_n N_VGND_c_1050_n 4.08582e-19 $X=3.635 $Y=1.065 $X2=0
+ $Y2=0
cc_547 N_A_639_125#_c_754_n N_VGND_c_1050_n 0.0244345f $X=4.525 $Y=1.15 $X2=0
+ $Y2=0
cc_548 N_A_639_125#_c_750_n N_VGND_c_1060_n 0.00425893f $X=4.97 $Y=1.185 $X2=0
+ $Y2=0
cc_549 N_A_639_125#_c_750_n N_VGND_c_1066_n 0.00715856f $X=4.97 $Y=1.185 $X2=0
+ $Y2=0
cc_550 N_A_639_125#_c_764_n A_725_125# 0.00294324f $X=3.545 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_551 N_A_639_125#_c_768_n A_725_125# 0.00191939f $X=3.635 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_552 N_RESET_B_M1006_g N_VPWR_c_883_n 5.85194e-19 $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_553 N_RESET_B_M1006_g N_VPWR_c_884_n 0.00585385f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_554 N_RESET_B_M1006_g N_VPWR_c_885_n 0.00248719f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_555 N_RESET_B_M1006_g N_VPWR_c_880_n 0.00646082f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_556 N_RESET_B_M1009_g N_VGND_c_1051_n 0.00607769f $X=5.33 $Y=0.655 $X2=0
+ $Y2=0
cc_557 N_RESET_B_M1009_g N_VGND_c_1060_n 0.00585385f $X=5.33 $Y=0.655 $X2=0
+ $Y2=0
cc_558 N_RESET_B_M1009_g N_VGND_c_1066_n 0.0110123f $X=5.33 $Y=0.655 $X2=0 $Y2=0
cc_559 N_VPWR_c_880_n N_Q_M1007_s 0.00579476f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_560 N_VPWR_c_880_n N_Q_M1015_s 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_561 N_VPWR_c_893_n N_Q_c_1031_n 0.0128008f $X=6.385 $Y=3.33 $X2=0 $Y2=0
cc_562 N_VPWR_c_880_n N_Q_c_1031_n 0.00730372f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_M1014_d N_Q_c_992_n 0.00176461f $X=6.41 $Y=1.835 $X2=0 $Y2=0
cc_564 N_VPWR_c_886_n N_Q_c_992_n 0.0170777f $X=6.55 $Y=2.19 $X2=0 $Y2=0
cc_565 N_VPWR_c_894_n N_Q_c_1035_n 0.0124525f $X=7.245 $Y=3.33 $X2=0 $Y2=0
cc_566 N_VPWR_c_880_n N_Q_c_1035_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_567 N_VPWR_M1025_d N_Q_c_994_n 0.00275378f $X=7.27 $Y=1.835 $X2=0 $Y2=0
cc_568 N_VPWR_c_888_n N_Q_c_994_n 0.023999f $X=7.41 $Y=2.19 $X2=0 $Y2=0
cc_569 N_Q_c_986_n N_VGND_c_1052_n 0.0216087f $X=6.885 $Y=1.17 $X2=0 $Y2=0
cc_570 N_Q_c_988_n N_VGND_c_1054_n 0.00539173f $X=7.345 $Y=1.17 $X2=0 $Y2=0
cc_571 N_Q_c_990_n N_VGND_c_1054_n 0.0211208f $X=7.47 $Y=1.255 $X2=0 $Y2=0
cc_572 N_Q_c_1022_n N_VGND_c_1061_n 0.0156097f $X=6.12 $Y=0.42 $X2=0 $Y2=0
cc_573 N_Q_c_1016_n N_VGND_c_1062_n 0.0124525f $X=6.98 $Y=0.42 $X2=0 $Y2=0
cc_574 N_Q_M1011_d N_VGND_c_1066_n 0.00380103f $X=5.98 $Y=0.235 $X2=0 $Y2=0
cc_575 N_Q_M1021_d N_VGND_c_1066_n 0.00536646f $X=6.84 $Y=0.235 $X2=0 $Y2=0
cc_576 N_Q_c_1016_n N_VGND_c_1066_n 0.00730901f $X=6.98 $Y=0.42 $X2=0 $Y2=0
cc_577 N_Q_c_1022_n N_VGND_c_1066_n 0.00980127f $X=6.12 $Y=0.42 $X2=0 $Y2=0
cc_578 N_VGND_c_1066_n A_1009_47# 0.00690169f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
