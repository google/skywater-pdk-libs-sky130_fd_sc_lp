* NGSPICE file created from sky130_fd_sc_lp__bufkapwr_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__bufkapwr_1 A KAPWR VGND VNB VPB VPWR X
M1000 a_69_161# A KAPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=3.528e+11p ps=3.08e+06u
M1001 VGND a_69_161# X VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.113e+11p ps=1.37e+06u
M1002 a_69_161# A VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 KAPWR a_69_161# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

