* File: sky130_fd_sc_lp__decap_6.pex.spice
* Created: Fri Aug 28 10:20:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAP_6%VGND 1 7 10 13 15 16 18 20 24 28 29 42
r26 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r27 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 36 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r29 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r30 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r31 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r32 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 30 38 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.25
+ $Y2=0
r34 30 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.72
+ $Y2=0
r35 29 41 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.665
+ $Y2=0
r36 29 35 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.16
+ $Y2=0
r37 24 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r38 24 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r39 20 22 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.615 $Y=0.405
+ $X2=2.615 $Y2=1.085
r40 18 41 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.665 $Y2=0
r41 18 20 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.405
r42 16 28 22.4154 $w=1.774e-06 $l=1.03959e-06 $layer=POLY_cond $X=0.915 $Y=1.77
+ $X2=1.4 $Y2=2.595
r43 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.915
+ $Y=1.77 $X2=0.915 $Y2=1.77
r44 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.5 $Y=1.77
+ $X2=0.915 $Y2=1.77
r45 10 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.335 $Y=0.38
+ $X2=0.335 $Y2=1.06
r46 8 13 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.5 $Y2=1.77
r47 8 12 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.335 $Y2=1.06
r48 7 38 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.25 $Y2=0
r49 7 10 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r50 1 22 121.333 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.615 $Y2=1.085
r51 1 20 121.333 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.615 $Y2=0.405
r52 1 12 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=0.335 $Y2=1.06
r53 1 10 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=0.335 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAP_6%VPWR 1 7 9 13 16 22 24 27 30 32 45
r25 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r26 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r28 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 36 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 35 38 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 33 41 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r33 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 32 44 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.632 $Y2=3.33
r35 32 38 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 27 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 27 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 24 26 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.55 $Y=2.29
+ $X2=2.55 $Y2=2.97
r39 22 44 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=2.55 $Y=3.245
+ $X2=2.632 $Y2=3.33
r40 22 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.55 $Y=3.245
+ $X2=2.55 $Y2=2.97
r41 21 24 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.55 $Y=1.675
+ $X2=2.55 $Y2=2.29
r42 16 30 20.7068 $w=1.804e-06 $l=7.75e-07 $layer=POLY_cond $X=1.48 $Y=1.51
+ $X2=1.48 $Y2=0.735
r43 16 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.51 $X2=2.32 $Y2=1.51
r44 15 19 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=1.64 $Y=1.507
+ $X2=2.32 $Y2=1.507
r45 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.64
+ $Y=1.51 $X2=1.64 $Y2=1.51
r46 13 21 6.81699 $w=3.35e-07 $l=2.36525e-07 $layer=LI1_cond $X=2.385 $Y=1.507
+ $X2=2.55 $Y2=1.675
r47 13 19 2.23608 $w=3.33e-07 $l=6.5e-08 $layer=LI1_cond $X=2.385 $Y=1.507
+ $X2=2.32 $Y2=1.507
r48 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.27 $X2=0.26
+ $Y2=2.95
r49 7 41 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r50 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r51 1 26 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=2.55 $Y2=2.97
r52 1 24 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=2.55 $Y2=2.29
r53 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=0.26 $Y2=2.95
r54 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=0.26 $Y2=2.27
.ends

