* File: sky130_fd_sc_lp__o2111a_lp.pxi.spice
* Created: Wed Sep  2 10:12:37 2020
* 
x_PM_SKY130_FD_SC_LP__O2111A_LP%A1 N_A1_M1011_g N_A1_M1012_g N_A1_c_83_n
+ N_A1_c_88_n A1 N_A1_c_84_n N_A1_c_85_n PM_SKY130_FD_SC_LP__O2111A_LP%A1
x_PM_SKY130_FD_SC_LP__O2111A_LP%A2 N_A2_M1000_g N_A2_M1010_g N_A2_c_114_n
+ N_A2_c_119_n A2 N_A2_c_116_n PM_SKY130_FD_SC_LP__O2111A_LP%A2
x_PM_SKY130_FD_SC_LP__O2111A_LP%B1 N_B1_M1005_g N_B1_M1009_g B1 B1 B1 B1
+ N_B1_c_153_n PM_SKY130_FD_SC_LP__O2111A_LP%B1
x_PM_SKY130_FD_SC_LP__O2111A_LP%C1 N_C1_M1003_g N_C1_c_196_n N_C1_M1007_g
+ N_C1_c_197_n C1 N_C1_c_201_n N_C1_c_198_n PM_SKY130_FD_SC_LP__O2111A_LP%C1
x_PM_SKY130_FD_SC_LP__O2111A_LP%D1 N_D1_c_248_n N_D1_M1004_g N_D1_c_249_n
+ N_D1_c_250_n N_D1_M1008_g D1 D1 N_D1_c_253_n PM_SKY130_FD_SC_LP__O2111A_LP%D1
x_PM_SKY130_FD_SC_LP__O2111A_LP%A_232_419# N_A_232_419#_M1004_d
+ N_A_232_419#_M1000_d N_A_232_419#_M1007_d N_A_232_419#_M1006_g
+ N_A_232_419#_M1002_g N_A_232_419#_M1001_g N_A_232_419#_c_301_n
+ N_A_232_419#_c_309_n N_A_232_419#_c_318_n N_A_232_419#_c_302_n
+ N_A_232_419#_c_331_n N_A_232_419#_c_303_n N_A_232_419#_c_304_n
+ N_A_232_419#_c_322_n N_A_232_419#_c_305_n N_A_232_419#_c_342_n
+ N_A_232_419#_c_311_n N_A_232_419#_c_306_n N_A_232_419#_c_307_n
+ N_A_232_419#_c_313_n N_A_232_419#_c_325_n N_A_232_419#_c_314_n
+ N_A_232_419#_c_348_n PM_SKY130_FD_SC_LP__O2111A_LP%A_232_419#
x_PM_SKY130_FD_SC_LP__O2111A_LP%VPWR N_VPWR_M1011_s N_VPWR_M1009_d
+ N_VPWR_M1008_d N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n
+ N_VPWR_c_424_n N_VPWR_c_425_n VPWR N_VPWR_c_426_n N_VPWR_c_427_n
+ N_VPWR_c_419_n N_VPWR_c_429_n PM_SKY130_FD_SC_LP__O2111A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O2111A_LP%X N_X_M1001_d N_X_M1002_d X X X X X X X X X
+ PM_SKY130_FD_SC_LP__O2111A_LP%X
x_PM_SKY130_FD_SC_LP__O2111A_LP%A_29_51# N_A_29_51#_M1012_s N_A_29_51#_M1010_d
+ N_A_29_51#_c_500_n N_A_29_51#_c_501_n N_A_29_51#_c_502_n N_A_29_51#_c_503_n
+ PM_SKY130_FD_SC_LP__O2111A_LP%A_29_51#
x_PM_SKY130_FD_SC_LP__O2111A_LP%VGND N_VGND_M1012_d N_VGND_M1006_s
+ N_VGND_c_526_n N_VGND_c_527_n VGND N_VGND_c_528_n N_VGND_c_529_n
+ N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n
+ PM_SKY130_FD_SC_LP__O2111A_LP%VGND
cc_1 VNB N_A1_M1012_g 0.0508978f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.465
cc_2 VNB N_A1_c_83_n 0.0198555f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.73
cc_3 VNB N_A1_c_84_n 0.0170919f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_4 VNB N_A1_c_85_n 0.0226492f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_5 VNB N_A2_M1010_g 0.0420751f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.465
cc_6 VNB N_A2_c_114_n 0.0153701f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.895
cc_7 VNB A2 0.00638022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_116_n 0.0143038f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_9 VNB N_B1_M1005_g 0.0556808f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_10 VNB B1 0.00754278f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_11 VNB N_B1_c_153_n 0.012055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C1_M1003_g 0.0369403f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_13 VNB N_C1_c_196_n 0.0299333f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.465
cc_14 VNB N_C1_c_197_n 0.0428962f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_C1_c_198_n 5.01531e-19 $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.56
cc_16 VNB N_D1_c_248_n 0.0198005f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.895
cc_17 VNB N_D1_c_249_n 0.0262257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D1_c_250_n 0.00641428f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.225
cc_19 VNB N_D1_M1008_g 0.0371788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB D1 0.0101453f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.895
cc_21 VNB N_D1_c_253_n 0.034576f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_22 VNB N_A_232_419#_M1006_g 0.0420776f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_A_232_419#_M1001_g 0.0418856f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.56
cc_24 VNB N_A_232_419#_c_301_n 0.0240228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_232_419#_c_302_n 0.00623401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_232_419#_c_303_n 0.00329266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_232_419#_c_304_n 0.00263251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_232_419#_c_305_n 0.00193136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_232_419#_c_306_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_232_419#_c_307_n 0.0235911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_419_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 0.0182758f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.465
cc_33 VNB X 0.0509701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_29_51#_c_500_n 0.0251921f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_35 VNB N_A_29_51#_c_501_n 0.0189359f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.895
cc_36 VNB N_A_29_51#_c_502_n 0.00998804f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_A_29_51#_c_503_n 0.00154554f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_38 VNB N_VGND_c_526_n 0.00634717f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.39
cc_39 VNB N_VGND_c_527_n 0.00727047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_528_n 0.0166014f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.56
cc_41 VNB N_VGND_c_529_n 0.0609979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_530_n 0.0268694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_531_n 0.261969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_532_n 0.00528596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_533_n 0.00510792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_A1_M1011_g 0.03531f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_47 VPB N_A1_c_83_n 0.00556555f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.73
cc_48 VPB N_A1_c_88_n 0.0144588f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.895
cc_49 VPB N_A1_c_85_n 0.0135265f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.39
cc_50 VPB N_A2_M1000_g 0.0285266f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_51 VPB N_A2_c_114_n 0.00430828f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.895
cc_52 VPB N_A2_c_119_n 0.0121324f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_53 VPB A2 0.00386934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B1_M1009_g 0.0314027f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.465
cc_55 VPB B1 0.0013085f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.39
cc_56 VPB N_B1_c_153_n 0.0200178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_C1_c_196_n 0.00176778f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.465
cc_58 VPB N_C1_M1007_g 0.0268409f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.39
cc_59 VPB N_C1_c_201_n 0.0283387f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.39
cc_60 VPB N_C1_c_198_n 0.00395059f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.56
cc_61 VPB N_D1_M1008_g 0.040772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_232_419#_M1002_g 0.0327794f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.39
cc_63 VPB N_A_232_419#_c_309_n 0.0168882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_232_419#_c_305_n 5.20321e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_232_419#_c_311_n 0.0120057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_232_419#_c_307_n 0.00424476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_232_419#_c_313_n 0.00811603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_232_419#_c_314_n 0.00203654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_420_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.73
cc_70 VPB N_VPWR_c_421_n 0.0443377f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_71 VPB N_VPWR_c_422_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_423_n 0.00315487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_424_n 0.0349125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_425_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_426_n 0.0298988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_427_n 0.0240188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_419_n 0.0477987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_429_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.0223616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB X 0.0236679f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.895
cc_81 VPB X 0.0367137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 N_A1_M1011_g N_A2_M1000_g 0.0280015f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_83 N_A1_M1012_g N_A2_M1010_g 0.0288693f $X=0.505 $Y=0.465 $X2=0 $Y2=0
cc_84 N_A1_c_83_n N_A2_c_114_n 0.0280015f $X=0.505 $Y=1.73 $X2=0 $Y2=0
cc_85 N_A1_c_88_n N_A2_c_119_n 0.0280015f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_86 N_A1_c_84_n A2 8.50898e-19 $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_87 N_A1_c_85_n A2 0.0403537f $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_88 N_A1_c_84_n N_A2_c_116_n 0.0280015f $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_89 N_A1_c_85_n N_A2_c_116_n 8.47756e-19 $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_90 N_A1_M1011_g N_VPWR_c_421_n 0.0268566f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_91 N_A1_c_88_n N_VPWR_c_421_n 0.00213543f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_92 N_A1_c_85_n N_VPWR_c_421_n 0.0279579f $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_93 N_A1_M1011_g N_VPWR_c_424_n 0.008763f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_94 N_A1_M1011_g N_VPWR_c_419_n 0.0144563f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_95 N_A1_M1012_g N_A_29_51#_c_500_n 0.00812036f $X=0.505 $Y=0.465 $X2=0 $Y2=0
cc_96 N_A1_M1012_g N_A_29_51#_c_501_n 0.0161798f $X=0.505 $Y=0.465 $X2=0 $Y2=0
cc_97 N_A1_c_84_n N_A_29_51#_c_501_n 0.00377547f $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_98 N_A1_c_85_n N_A_29_51#_c_501_n 0.0218428f $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_99 N_A1_c_84_n N_A_29_51#_c_502_n 9.34252e-19 $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_100 N_A1_c_85_n N_A_29_51#_c_502_n 0.0222093f $X=0.505 $Y=1.39 $X2=0 $Y2=0
cc_101 N_A1_M1012_g N_A_29_51#_c_503_n 9.70813e-19 $X=0.505 $Y=0.465 $X2=0 $Y2=0
cc_102 N_A1_M1012_g N_VGND_c_526_n 0.0111508f $X=0.505 $Y=0.465 $X2=0 $Y2=0
cc_103 N_A1_M1012_g N_VGND_c_528_n 0.00469214f $X=0.505 $Y=0.465 $X2=0 $Y2=0
cc_104 N_A1_M1012_g N_VGND_c_531_n 0.00913919f $X=0.505 $Y=0.465 $X2=0 $Y2=0
cc_105 N_A2_M1010_g N_B1_M1005_g 0.0247267f $X=1.015 $Y=0.465 $X2=0 $Y2=0
cc_106 A2 N_B1_M1005_g 0.00406525f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A2_c_116_n N_B1_M1005_g 0.0171548f $X=1.075 $Y=1.39 $X2=0 $Y2=0
cc_108 N_A2_M1000_g N_B1_M1009_g 0.0244511f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_109 N_A2_M1010_g B1 0.00141833f $X=1.015 $Y=0.465 $X2=0 $Y2=0
cc_110 A2 B1 0.0516819f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A2_c_116_n B1 7.1475e-19 $X=1.075 $Y=1.39 $X2=0 $Y2=0
cc_112 N_A2_c_114_n N_B1_c_153_n 0.0171548f $X=1.075 $Y=1.73 $X2=0 $Y2=0
cc_113 N_A2_M1000_g N_A_232_419#_c_313_n 0.00212895f $X=1.035 $Y=2.595 $X2=0
+ $Y2=0
cc_114 N_A2_c_119_n N_A_232_419#_c_313_n 0.00170835f $X=1.075 $Y=1.895 $X2=0
+ $Y2=0
cc_115 A2 N_A_232_419#_c_313_n 0.0121443f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A2_M1000_g N_VPWR_c_421_n 0.0053152f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_117 N_A2_M1000_g N_VPWR_c_422_n 9.76482e-19 $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_118 N_A2_M1000_g N_VPWR_c_424_n 0.00975641f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_119 N_A2_M1000_g N_VPWR_c_419_n 0.0170985f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_120 N_A2_M1010_g N_A_29_51#_c_501_n 0.0142897f $X=1.015 $Y=0.465 $X2=0 $Y2=0
cc_121 A2 N_A_29_51#_c_501_n 0.0327429f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_122 N_A2_c_116_n N_A_29_51#_c_501_n 0.00481644f $X=1.075 $Y=1.39 $X2=0 $Y2=0
cc_123 N_A2_M1010_g N_A_29_51#_c_503_n 0.0105866f $X=1.015 $Y=0.465 $X2=0 $Y2=0
cc_124 N_A2_M1010_g N_VGND_c_526_n 0.00534205f $X=1.015 $Y=0.465 $X2=0 $Y2=0
cc_125 N_A2_M1010_g N_VGND_c_529_n 0.00530134f $X=1.015 $Y=0.465 $X2=0 $Y2=0
cc_126 N_A2_M1010_g N_VGND_c_531_n 0.0101885f $X=1.015 $Y=0.465 $X2=0 $Y2=0
cc_127 N_B1_M1005_g N_C1_M1003_g 0.0617296f $X=1.555 $Y=0.465 $X2=0 $Y2=0
cc_128 B1 N_C1_M1003_g 0.00761472f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_129 N_B1_M1005_g N_C1_c_196_n 0.00571611f $X=1.555 $Y=0.465 $X2=0 $Y2=0
cc_130 B1 N_C1_c_196_n 0.00497255f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_131 N_B1_c_153_n N_C1_c_196_n 0.0179854f $X=1.66 $Y=1.73 $X2=0 $Y2=0
cc_132 N_B1_M1009_g N_C1_M1007_g 0.0201081f $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_133 N_B1_M1009_g N_C1_c_201_n 0.00135686f $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_134 N_B1_M1009_g N_C1_c_198_n 0.00488135f $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_135 B1 N_C1_c_198_n 0.0183642f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_B1_c_153_n N_C1_c_198_n 0.00172594f $X=1.66 $Y=1.73 $X2=0 $Y2=0
cc_137 N_B1_M1009_g N_A_232_419#_c_318_n 0.0176196f $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_138 B1 N_A_232_419#_c_318_n 0.0105142f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_B1_c_153_n N_A_232_419#_c_318_n 3.56637e-19 $X=1.66 $Y=1.73 $X2=0 $Y2=0
cc_140 B1 N_A_232_419#_c_302_n 0.0298022f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_141 B1 N_A_232_419#_c_322_n 0.00816666f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_142 N_B1_M1009_g N_A_232_419#_c_313_n 0.0125124f $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_143 B1 N_A_232_419#_c_313_n 6.4651e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_144 N_B1_M1009_g N_A_232_419#_c_325_n 0.0172616f $X=1.605 $Y=2.595 $X2=0
+ $Y2=0
cc_145 N_B1_M1009_g N_VPWR_c_422_n 0.0133867f $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_146 N_B1_M1009_g N_VPWR_c_424_n 0.00840199f $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_147 N_B1_M1009_g N_VPWR_c_419_n 0.00765867f $X=1.605 $Y=2.595 $X2=0 $Y2=0
cc_148 N_B1_M1005_g N_A_29_51#_c_501_n 0.00131922f $X=1.555 $Y=0.465 $X2=0 $Y2=0
cc_149 B1 N_A_29_51#_c_501_n 0.0137323f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_150 N_B1_M1005_g N_A_29_51#_c_503_n 0.00719106f $X=1.555 $Y=0.465 $X2=0 $Y2=0
cc_151 B1 N_A_29_51#_c_503_n 0.031883f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_152 N_B1_M1005_g N_VGND_c_529_n 0.00398294f $X=1.555 $Y=0.465 $X2=0 $Y2=0
cc_153 B1 N_VGND_c_529_n 0.009163f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_154 N_B1_M1005_g N_VGND_c_531_n 0.00613513f $X=1.555 $Y=0.465 $X2=0 $Y2=0
cc_155 B1 N_VGND_c_531_n 0.0107685f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_156 B1 A_326_51# 0.00178904f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_157 N_C1_M1003_g N_D1_c_248_n 0.040991f $X=1.945 $Y=0.465 $X2=-0.19
+ $Y2=-0.245
cc_158 N_C1_c_197_n N_D1_c_250_n 0.0167183f $X=2.225 $Y=1.325 $X2=0 $Y2=0
cc_159 N_C1_c_197_n N_D1_M1008_g 0.0549643f $X=2.225 $Y=1.325 $X2=0 $Y2=0
cc_160 N_C1_c_198_n N_D1_M1008_g 2.54593e-19 $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_161 N_C1_c_197_n D1 4.61465e-19 $X=2.225 $Y=1.325 $X2=0 $Y2=0
cc_162 N_C1_M1007_g N_A_232_419#_c_318_n 0.0218149f $X=2.455 $Y=2.595 $X2=0
+ $Y2=0
cc_163 N_C1_c_201_n N_A_232_419#_c_318_n 0.00103266f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_164 N_C1_c_198_n N_A_232_419#_c_318_n 0.0219176f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_165 N_C1_M1003_g N_A_232_419#_c_302_n 0.00797843f $X=1.945 $Y=0.465 $X2=0
+ $Y2=0
cc_166 N_C1_c_197_n N_A_232_419#_c_302_n 0.00740312f $X=2.225 $Y=1.325 $X2=0
+ $Y2=0
cc_167 N_C1_M1003_g N_A_232_419#_c_331_n 0.00450676f $X=1.945 $Y=0.465 $X2=0
+ $Y2=0
cc_168 N_C1_c_197_n N_A_232_419#_c_303_n 2.61099e-19 $X=2.225 $Y=1.325 $X2=0
+ $Y2=0
cc_169 N_C1_c_196_n N_A_232_419#_c_304_n 0.0119042f $X=2.322 $Y=1.678 $X2=0
+ $Y2=0
cc_170 N_C1_c_197_n N_A_232_419#_c_304_n 0.00468757f $X=2.225 $Y=1.325 $X2=0
+ $Y2=0
cc_171 N_C1_c_198_n N_A_232_419#_c_304_n 0.00346123f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_172 N_C1_c_196_n N_A_232_419#_c_322_n 0.00557689f $X=2.322 $Y=1.678 $X2=0
+ $Y2=0
cc_173 N_C1_c_197_n N_A_232_419#_c_322_n 0.00190612f $X=2.225 $Y=1.325 $X2=0
+ $Y2=0
cc_174 N_C1_c_198_n N_A_232_419#_c_322_n 0.0134922f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_175 N_C1_c_196_n N_A_232_419#_c_305_n 0.0104355f $X=2.322 $Y=1.678 $X2=0
+ $Y2=0
cc_176 N_C1_c_201_n N_A_232_419#_c_305_n 8.03294e-19 $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_177 N_C1_c_198_n N_A_232_419#_c_305_n 0.00675284f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_178 N_C1_M1007_g N_A_232_419#_c_342_n 0.0128275f $X=2.455 $Y=2.595 $X2=0
+ $Y2=0
cc_179 N_C1_c_201_n N_A_232_419#_c_342_n 0.00132828f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_180 N_C1_c_198_n N_A_232_419#_c_342_n 0.018974f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_181 N_C1_c_198_n N_A_232_419#_c_313_n 0.00240729f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_182 N_C1_c_201_n N_A_232_419#_c_314_n 0.00476001f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_183 N_C1_c_198_n N_A_232_419#_c_314_n 0.0130141f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_184 N_C1_M1007_g N_A_232_419#_c_348_n 0.0189481f $X=2.455 $Y=2.595 $X2=0
+ $Y2=0
cc_185 N_C1_c_198_n N_VPWR_M1009_d 0.00358002f $X=2.23 $Y=1.77 $X2=0 $Y2=0
cc_186 N_C1_M1007_g N_VPWR_c_422_n 0.00702976f $X=2.455 $Y=2.595 $X2=0 $Y2=0
cc_187 N_C1_M1007_g N_VPWR_c_423_n 0.00125577f $X=2.455 $Y=2.595 $X2=0 $Y2=0
cc_188 N_C1_M1007_g N_VPWR_c_426_n 0.00969624f $X=2.455 $Y=2.595 $X2=0 $Y2=0
cc_189 N_C1_M1007_g N_VPWR_c_419_n 0.0103115f $X=2.455 $Y=2.595 $X2=0 $Y2=0
cc_190 N_C1_M1003_g N_VGND_c_529_n 0.00565115f $X=1.945 $Y=0.465 $X2=0 $Y2=0
cc_191 N_C1_M1003_g N_VGND_c_531_n 0.0106215f $X=1.945 $Y=0.465 $X2=0 $Y2=0
cc_192 N_D1_M1008_g N_A_232_419#_M1006_g 0.0407639f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_193 D1 N_A_232_419#_M1006_g 0.00874822f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_194 N_D1_c_253_n N_A_232_419#_M1006_g 0.0165982f $X=2.985 $Y=0.84 $X2=0 $Y2=0
cc_195 N_D1_M1008_g N_A_232_419#_M1002_g 0.0163172f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_196 N_D1_c_248_n N_A_232_419#_c_302_n 0.00888336f $X=2.335 $Y=0.765 $X2=0
+ $Y2=0
cc_197 N_D1_c_250_n N_A_232_419#_c_302_n 0.00492264f $X=2.41 $Y=0.84 $X2=0 $Y2=0
cc_198 N_D1_M1008_g N_A_232_419#_c_302_n 0.00235206f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_199 D1 N_A_232_419#_c_302_n 0.0246339f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_200 N_D1_c_253_n N_A_232_419#_c_302_n 9.23355e-19 $X=2.985 $Y=0.84 $X2=0
+ $Y2=0
cc_201 N_D1_c_248_n N_A_232_419#_c_331_n 0.00434901f $X=2.335 $Y=0.765 $X2=0
+ $Y2=0
cc_202 N_D1_c_248_n N_A_232_419#_c_303_n 0.00350267f $X=2.335 $Y=0.765 $X2=0
+ $Y2=0
cc_203 N_D1_c_249_n N_A_232_419#_c_303_n 0.00666746f $X=2.82 $Y=0.84 $X2=0 $Y2=0
cc_204 D1 N_A_232_419#_c_303_n 0.0133764f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_205 N_D1_c_249_n N_A_232_419#_c_304_n 9.34463e-19 $X=2.82 $Y=0.84 $X2=0 $Y2=0
cc_206 N_D1_c_250_n N_A_232_419#_c_304_n 0.00101374f $X=2.41 $Y=0.84 $X2=0 $Y2=0
cc_207 N_D1_M1008_g N_A_232_419#_c_304_n 0.00243433f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_208 D1 N_A_232_419#_c_304_n 0.0179606f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_209 N_D1_M1008_g N_A_232_419#_c_305_n 0.00330684f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_210 N_D1_M1008_g N_A_232_419#_c_342_n 0.0106949f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_211 N_D1_M1008_g N_A_232_419#_c_311_n 0.0208594f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_212 D1 N_A_232_419#_c_311_n 0.0086399f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_213 N_D1_c_253_n N_A_232_419#_c_311_n 3.17332e-19 $X=2.985 $Y=0.84 $X2=0
+ $Y2=0
cc_214 N_D1_M1008_g N_A_232_419#_c_306_n 0.0021794f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_215 N_D1_M1008_g N_A_232_419#_c_314_n 0.00326325f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_216 D1 N_A_232_419#_c_314_n 0.00519405f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_217 N_D1_c_253_n N_A_232_419#_c_314_n 0.00102784f $X=2.985 $Y=0.84 $X2=0
+ $Y2=0
cc_218 N_D1_M1008_g N_A_232_419#_c_348_n 0.0159628f $X=3.005 $Y=2.595 $X2=0
+ $Y2=0
cc_219 N_D1_M1008_g N_VPWR_c_423_n 0.022803f $X=3.005 $Y=2.595 $X2=0 $Y2=0
cc_220 N_D1_M1008_g N_VPWR_c_426_n 0.00840199f $X=3.005 $Y=2.595 $X2=0 $Y2=0
cc_221 N_D1_M1008_g N_VPWR_c_419_n 0.0136513f $X=3.005 $Y=2.595 $X2=0 $Y2=0
cc_222 N_D1_M1008_g X 2.55579e-19 $X=3.005 $Y=2.595 $X2=0 $Y2=0
cc_223 N_D1_c_248_n N_VGND_c_527_n 0.00234637f $X=2.335 $Y=0.765 $X2=0 $Y2=0
cc_224 D1 N_VGND_c_527_n 0.0116883f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_225 N_D1_c_253_n N_VGND_c_527_n 0.00165197f $X=2.985 $Y=0.84 $X2=0 $Y2=0
cc_226 N_D1_c_248_n N_VGND_c_529_n 0.00356196f $X=2.335 $Y=0.765 $X2=0 $Y2=0
cc_227 N_D1_c_249_n N_VGND_c_529_n 0.0069324f $X=2.82 $Y=0.84 $X2=0 $Y2=0
cc_228 N_D1_c_248_n N_VGND_c_531_n 0.0063571f $X=2.335 $Y=0.765 $X2=0 $Y2=0
cc_229 N_D1_c_249_n N_VGND_c_531_n 0.00915314f $X=2.82 $Y=0.84 $X2=0 $Y2=0
cc_230 D1 N_VGND_c_531_n 0.0139772f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_231 N_A_232_419#_c_318_n N_VPWR_M1009_d 0.0207751f $X=2.575 $Y=2.415 $X2=0
+ $Y2=0
cc_232 N_A_232_419#_c_318_n N_VPWR_c_422_n 0.0204369f $X=2.575 $Y=2.415 $X2=0
+ $Y2=0
cc_233 N_A_232_419#_c_325_n N_VPWR_c_422_n 0.0253679f $X=1.34 $Y=2.415 $X2=0
+ $Y2=0
cc_234 N_A_232_419#_c_348_n N_VPWR_c_422_n 0.0121271f $X=2.74 $Y=2.415 $X2=0
+ $Y2=0
cc_235 N_A_232_419#_M1002_g N_VPWR_c_423_n 0.0239884f $X=3.535 $Y=2.595 $X2=0
+ $Y2=0
cc_236 N_A_232_419#_c_309_n N_VPWR_c_423_n 5.38456e-19 $X=3.567 $Y=1.885 $X2=0
+ $Y2=0
cc_237 N_A_232_419#_c_342_n N_VPWR_c_423_n 0.0167692f $X=2.74 $Y=2.24 $X2=0
+ $Y2=0
cc_238 N_A_232_419#_c_311_n N_VPWR_c_423_n 0.0252391f $X=3.415 $Y=1.8 $X2=0
+ $Y2=0
cc_239 N_A_232_419#_c_348_n N_VPWR_c_423_n 0.0491014f $X=2.74 $Y=2.415 $X2=0
+ $Y2=0
cc_240 N_A_232_419#_c_325_n N_VPWR_c_424_n 0.0183971f $X=1.34 $Y=2.415 $X2=0
+ $Y2=0
cc_241 N_A_232_419#_c_348_n N_VPWR_c_426_n 0.0178372f $X=2.74 $Y=2.415 $X2=0
+ $Y2=0
cc_242 N_A_232_419#_M1002_g N_VPWR_c_427_n 0.00840199f $X=3.535 $Y=2.595 $X2=0
+ $Y2=0
cc_243 N_A_232_419#_M1000_d N_VPWR_c_419_n 0.00308191f $X=1.16 $Y=2.095 $X2=0
+ $Y2=0
cc_244 N_A_232_419#_M1007_d N_VPWR_c_419_n 0.00239922f $X=2.58 $Y=2.095 $X2=0
+ $Y2=0
cc_245 N_A_232_419#_M1002_g N_VPWR_c_419_n 0.0146764f $X=3.535 $Y=2.595 $X2=0
+ $Y2=0
cc_246 N_A_232_419#_c_318_n N_VPWR_c_419_n 0.0237356f $X=2.575 $Y=2.415 $X2=0
+ $Y2=0
cc_247 N_A_232_419#_c_325_n N_VPWR_c_419_n 0.012508f $X=1.34 $Y=2.415 $X2=0
+ $Y2=0
cc_248 N_A_232_419#_c_348_n N_VPWR_c_419_n 0.0124168f $X=2.74 $Y=2.415 $X2=0
+ $Y2=0
cc_249 N_A_232_419#_M1006_g X 0.00132239f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A_232_419#_M1001_g X 0.00863077f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_251 N_A_232_419#_M1002_g X 0.00617829f $X=3.535 $Y=2.595 $X2=0 $Y2=0
cc_252 N_A_232_419#_M1001_g X 0.0258726f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_253 N_A_232_419#_c_309_n X 0.00116864f $X=3.567 $Y=1.885 $X2=0 $Y2=0
cc_254 N_A_232_419#_c_311_n X 0.0114669f $X=3.415 $Y=1.8 $X2=0 $Y2=0
cc_255 N_A_232_419#_c_306_n X 0.0317254f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_256 N_A_232_419#_c_307_n X 0.0077371f $X=3.58 $Y=1.38 $X2=0 $Y2=0
cc_257 N_A_232_419#_M1002_g X 0.00567693f $X=3.535 $Y=2.595 $X2=0 $Y2=0
cc_258 N_A_232_419#_c_309_n X 6.55705e-19 $X=3.567 $Y=1.885 $X2=0 $Y2=0
cc_259 N_A_232_419#_c_311_n X 0.00881185f $X=3.415 $Y=1.8 $X2=0 $Y2=0
cc_260 N_A_232_419#_M1002_g X 0.0184472f $X=3.535 $Y=2.595 $X2=0 $Y2=0
cc_261 N_A_232_419#_M1006_g N_VGND_c_527_n 0.0126882f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_262 N_A_232_419#_M1001_g N_VGND_c_527_n 0.00215298f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_263 N_A_232_419#_c_303_n N_VGND_c_527_n 0.0135699f $X=2.55 $Y=0.41 $X2=0
+ $Y2=0
cc_264 N_A_232_419#_c_331_n N_VGND_c_529_n 0.00705866f $X=2.345 $Y=0.45 $X2=0
+ $Y2=0
cc_265 N_A_232_419#_c_303_n N_VGND_c_529_n 0.0161587f $X=2.55 $Y=0.41 $X2=0
+ $Y2=0
cc_266 N_A_232_419#_M1006_g N_VGND_c_530_n 0.00486043f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_267 N_A_232_419#_M1001_g N_VGND_c_530_n 0.00549284f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_268 N_A_232_419#_M1006_g N_VGND_c_531_n 0.00814425f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_269 N_A_232_419#_M1001_g N_VGND_c_531_n 0.010905f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_270 N_A_232_419#_c_331_n N_VGND_c_531_n 0.00600452f $X=2.345 $Y=0.45 $X2=0
+ $Y2=0
cc_271 N_A_232_419#_c_303_n N_VGND_c_531_n 0.0132406f $X=2.55 $Y=0.41 $X2=0
+ $Y2=0
cc_272 N_A_232_419#_c_302_n A_404_51# 9.97626e-19 $X=2.26 $Y=1.265 $X2=-0.19
+ $Y2=-0.245
cc_273 N_A_232_419#_c_331_n A_404_51# 0.00362145f $X=2.345 $Y=0.45 $X2=-0.19
+ $Y2=-0.245
cc_274 N_VPWR_c_419_n A_134_419# 0.010279f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_275 N_VPWR_c_419_n N_X_M1002_d 0.0023218f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_276 N_VPWR_c_423_n X 0.0680384f $X=3.27 $Y=2.24 $X2=0 $Y2=0
cc_277 N_VPWR_c_427_n X 0.0359399f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_278 N_VPWR_c_419_n X 0.0217944f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_279 X N_VGND_c_527_n 0.0107064f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_280 X N_VGND_c_530_n 0.0197155f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_281 N_X_M1001_d N_VGND_c_531_n 0.00232985f $X=3.9 $Y=0.235 $X2=0 $Y2=0
cc_282 X N_VGND_c_531_n 0.0125355f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_283 N_A_29_51#_c_500_n N_VGND_c_526_n 0.0161397f $X=0.29 $Y=0.48 $X2=0 $Y2=0
cc_284 N_A_29_51#_c_501_n N_VGND_c_526_n 0.0264018f $X=1.065 $Y=0.96 $X2=0 $Y2=0
cc_285 N_A_29_51#_c_503_n N_VGND_c_526_n 0.015529f $X=1.23 $Y=0.48 $X2=0 $Y2=0
cc_286 N_A_29_51#_c_500_n N_VGND_c_528_n 0.0163773f $X=0.29 $Y=0.48 $X2=0 $Y2=0
cc_287 N_A_29_51#_c_503_n N_VGND_c_529_n 0.0144775f $X=1.23 $Y=0.48 $X2=0 $Y2=0
cc_288 N_A_29_51#_c_500_n N_VGND_c_531_n 0.00959046f $X=0.29 $Y=0.48 $X2=0 $Y2=0
cc_289 N_A_29_51#_c_503_n N_VGND_c_531_n 0.00948536f $X=1.23 $Y=0.48 $X2=0 $Y2=0
cc_290 N_VGND_c_531_n A_708_47# 0.00899413f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
