* File: sky130_fd_sc_lp__nor2_4.pex.spice
* Created: Fri Aug 28 10:53:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31 43
+ 45
r77 44 45 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.565 $Y=1.395
+ $X2=1.995 $Y2=1.395
r78 42 44 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.44 $Y=1.395
+ $X2=1.565 $Y2=1.395
r79 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.44
+ $Y=1.395 $X2=1.44 $Y2=1.395
r80 40 42 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.135 $Y=1.395
+ $X2=1.44 $Y2=1.395
r81 38 40 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.76 $Y=1.395
+ $X2=1.135 $Y2=1.395
r82 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.395 $X2=0.76 $Y2=1.395
r83 35 38 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.705 $Y=1.395
+ $X2=0.76 $Y2=1.395
r84 31 43 7.90247 $w=3.48e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=1.385
+ $X2=1.44 $Y2=1.385
r85 31 39 14.4879 $w=3.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.2 $Y=1.385
+ $X2=0.76 $Y2=1.385
r86 30 39 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.72 $Y=1.385 $X2=0.76
+ $Y2=1.385
r87 29 30 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.385
+ $X2=0.72 $Y2=1.385
r88 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.995 $Y=1.56
+ $X2=1.995 $Y2=1.395
r89 25 27 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.995 $Y=1.56
+ $X2=1.995 $Y2=2.465
r90 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.995 $Y=1.23
+ $X2=1.995 $Y2=1.395
r91 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.995 $Y=1.23
+ $X2=1.995 $Y2=0.7
r92 18 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=1.56
+ $X2=1.565 $Y2=1.395
r93 18 20 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.565 $Y=1.56
+ $X2=1.565 $Y2=2.465
r94 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=1.23
+ $X2=1.565 $Y2=1.395
r95 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.565 $Y=1.23
+ $X2=1.565 $Y2=0.7
r96 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.56
+ $X2=1.135 $Y2=1.395
r97 11 13 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.135 $Y=1.56
+ $X2=1.135 $Y2=2.465
r98 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.23
+ $X2=1.135 $Y2=1.395
r99 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.135 $Y=1.23
+ $X2=1.135 $Y2=0.7
r100 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.56
+ $X2=0.705 $Y2=1.395
r101 4 6 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=0.705 $Y=1.56
+ $X2=0.705 $Y2=2.465
r102 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.23
+ $X2=0.705 $Y2=1.395
r103 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.705 $Y=1.23
+ $X2=0.705 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_4%B 1 3 6 8 10 13 17 21 23 25 29 31 32 33
r75 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.75
+ $Y=1.51 $X2=3.75 $Y2=1.51
r76 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.51 $X2=3.41 $Y2=1.51
r77 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.51 $X2=3.07 $Y2=1.51
r78 38 40 27.9326 $w=3.71e-07 $l=2.15e-07 $layer=POLY_cond $X=2.855 $Y=1.452
+ $X2=3.07 $Y2=1.452
r79 37 38 55.8652 $w=3.71e-07 $l=4.3e-07 $layer=POLY_cond $X=2.425 $Y=1.452
+ $X2=2.855 $Y2=1.452
r80 33 49 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=4.08 $Y=1.592
+ $X2=3.75 $Y2=1.592
r81 32 49 5.16019 $w=3.33e-07 $l=1.5e-07 $layer=LI1_cond $X=3.6 $Y=1.592
+ $X2=3.75 $Y2=1.592
r82 32 45 6.53624 $w=3.33e-07 $l=1.9e-07 $layer=LI1_cond $X=3.6 $Y=1.592
+ $X2=3.41 $Y2=1.592
r83 31 45 9.97637 $w=3.33e-07 $l=2.9e-07 $layer=LI1_cond $X=3.12 $Y=1.592
+ $X2=3.41 $Y2=1.592
r84 31 41 1.72006 $w=3.33e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.592 $X2=3.07
+ $Y2=1.592
r85 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.715 $Y=1.675
+ $X2=3.715 $Y2=2.465
r86 23 48 4.54717 $w=3.71e-07 $l=3.5e-08 $layer=POLY_cond $X=3.715 $Y=1.452
+ $X2=3.75 $Y2=1.452
r87 23 27 24.032 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.715 $Y=1.452
+ $X2=3.715 $Y2=1.675
r88 23 44 39.6253 $w=3.71e-07 $l=3.05e-07 $layer=POLY_cond $X=3.715 $Y=1.452
+ $X2=3.41 $Y2=1.452
r89 23 25 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.715 $Y=1.345
+ $X2=3.715 $Y2=0.7
r90 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.285 $Y=1.675
+ $X2=3.285 $Y2=2.465
r91 15 44 16.2399 $w=3.71e-07 $l=1.25e-07 $layer=POLY_cond $X=3.285 $Y=1.452
+ $X2=3.41 $Y2=1.452
r92 15 19 24.032 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.285 $Y=1.452
+ $X2=3.285 $Y2=1.675
r93 15 40 27.9326 $w=3.71e-07 $l=2.15e-07 $layer=POLY_cond $X=3.285 $Y=1.452
+ $X2=3.07 $Y2=1.452
r94 15 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.285 $Y=1.345
+ $X2=3.285 $Y2=0.7
r95 11 38 24.032 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.855 $Y=1.675
+ $X2=2.855 $Y2=1.452
r96 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.855 $Y=1.675
+ $X2=2.855 $Y2=2.465
r97 8 38 24.032 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.855 $Y=1.23
+ $X2=2.855 $Y2=1.452
r98 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.855 $Y=1.23
+ $X2=2.855 $Y2=0.7
r99 4 37 24.032 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.425 $Y=1.675
+ $X2=2.425 $Y2=1.452
r100 4 6 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.425 $Y=1.675
+ $X2=2.425 $Y2=2.465
r101 1 37 24.032 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.425 $Y=1.23
+ $X2=2.425 $Y2=1.452
r102 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.425 $Y=1.23
+ $X2=2.425 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_4%A_73_367# 1 2 3 4 5 18 22 23 26 30 33 36 40
+ 42 44 46 48 51
r57 44 53 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=2.905
+ $X2=3.95 $Y2=2.99
r58 44 46 32.1889 $w=2.88e-07 $l=8.1e-07 $layer=LI1_cond $X=3.95 $Y=2.905
+ $X2=3.95 $Y2=2.095
r59 43 51 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=3.205 $Y=2.99
+ $X2=3.077 $Y2=2.99
r60 42 53 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.805 $Y=2.99
+ $X2=3.95 $Y2=2.99
r61 42 43 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.805 $Y=2.99
+ $X2=3.205 $Y2=2.99
r62 38 51 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.077 $Y=2.905
+ $X2=3.077 $Y2=2.99
r63 38 40 19.8853 $w=2.53e-07 $l=4.4e-07 $layer=LI1_cond $X=3.077 $Y=2.905
+ $X2=3.077 $Y2=2.465
r64 37 50 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.335 $Y=2.99
+ $X2=2.225 $Y2=2.99
r65 36 51 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.95 $Y=2.99
+ $X2=3.077 $Y2=2.99
r66 36 37 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.95 $Y=2.99
+ $X2=2.335 $Y2=2.99
r67 33 50 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.905
+ $X2=2.225 $Y2=2.99
r68 33 35 48.455 $w=2.18e-07 $l=9.25e-07 $layer=LI1_cond $X=2.225 $Y=2.905
+ $X2=2.225 $Y2=1.98
r69 32 35 2.88111 $w=2.18e-07 $l=5.5e-08 $layer=LI1_cond $X=2.225 $Y=1.925
+ $X2=2.225 $Y2=1.98
r70 31 48 5.05528 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=1.445 $Y=1.827
+ $X2=1.35 $Y2=1.827
r71 30 32 6.84872 $w=1.95e-07 $l=1.51261e-07 $layer=LI1_cond $X=2.115 $Y=1.827
+ $X2=2.225 $Y2=1.925
r72 30 31 38.1072 $w=1.93e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=1.827
+ $X2=1.445 $Y2=1.827
r73 26 28 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.35 $Y=1.98
+ $X2=1.35 $Y2=2.91
r74 24 48 1.43626 $w=1.9e-07 $l=9.8e-08 $layer=LI1_cond $X=1.35 $Y=1.925
+ $X2=1.35 $Y2=1.827
r75 24 26 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.35 $Y=1.925
+ $X2=1.35 $Y2=1.98
r76 22 48 5.05528 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=1.255 $Y=1.827
+ $X2=1.35 $Y2=1.827
r77 22 23 38.1072 $w=1.93e-07 $l=6.7e-07 $layer=LI1_cond $X=1.255 $Y=1.827
+ $X2=0.585 $Y2=1.827
r78 18 20 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.455 $Y=1.98
+ $X2=0.455 $Y2=2.91
r79 16 23 6.999 $w=1.95e-07 $l=1.72163e-07 $layer=LI1_cond $X=0.455 $Y=1.925
+ $X2=0.585 $Y2=1.827
r80 16 18 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=0.455 $Y=1.925
+ $X2=0.455 $Y2=1.98
r81 5 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.79
+ $Y=1.835 $X2=3.93 $Y2=2.91
r82 5 46 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.79
+ $Y=1.835 $X2=3.93 $Y2=2.095
r83 4 40 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=2.93
+ $Y=1.835 $X2=3.07 $Y2=2.465
r84 3 50 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.07
+ $Y=1.835 $X2=2.21 $Y2=2.91
r85 3 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.07
+ $Y=1.835 $X2=2.21 $Y2=1.98
r86 2 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.21
+ $Y=1.835 $X2=1.35 $Y2=2.91
r87 2 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.21
+ $Y=1.835 $X2=1.35 $Y2=1.98
r88 1 20 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.835 $X2=0.49 $Y2=2.91
r89 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.835 $X2=0.49 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_4%VPWR 1 2 9 13 17 21 22 23 34 35 38
r57 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 31 34 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.78 $Y2=3.33
r61 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 27 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 23 35 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 23 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 23 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r67 21 26 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.92 $Y2=3.33
r69 17 20 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.78 $Y=2.18
+ $X2=1.78 $Y2=2.95
r70 15 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=3.245
+ $X2=1.78 $Y2=3.33
r71 15 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.78 $Y=3.245
+ $X2=1.78 $Y2=2.95
r72 14 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.92 $Y2=3.33
r73 13 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.78 $Y2=3.33
r74 13 14 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.085 $Y2=3.33
r75 9 12 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.92 $Y=2.18 $X2=0.92
+ $Y2=2.95
r76 7 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=3.245 $X2=0.92
+ $Y2=3.33
r77 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=2.95
r78 2 20 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.64
+ $Y=1.835 $X2=1.78 $Y2=2.95
r79 2 17 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.64
+ $Y=1.835 $X2=1.78 $Y2=2.18
r80 1 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.78
+ $Y=1.835 $X2=0.92 $Y2=2.95
r81 1 9 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=0.78
+ $Y=1.835 $X2=0.92 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_4%Y 1 2 3 4 5 6 21 23 24 27 30 31 32 33 35 41
+ 46 47 48 49 50 51 61 67 75
r92 67 80 6.25913 $w=2.3e-07 $l=1.18e-07 $layer=LI1_cond $X=2.62 $Y=1.56
+ $X2=2.62 $Y2=1.442
r93 59 77 4.56828 $w=2.27e-07 $l=8.59942e-08 $layer=LI1_cond $X=2.622 $Y=1.085
+ $X2=2.62 $Y2=1.17
r94 51 75 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=2.642 $Y=2.035
+ $X2=2.642 $Y2=2.12
r95 51 75 0.0388969 $w=6.13e-07 $l=2e-09 $layer=LI1_cond $X=2.64 $Y=2.427
+ $X2=2.642 $Y2=2.427
r96 50 51 10.2753 $w=3.98e-07 $l=2.85e-07 $layer=LI1_cond $X=2.62 $Y=1.665
+ $X2=2.62 $Y2=1.95
r97 50 67 5.26115 $w=2.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.62 $Y=1.665
+ $X2=2.62 $Y2=1.56
r98 49 80 7.90044 $w=2.27e-07 $l=1.47e-07 $layer=LI1_cond $X=2.62 $Y=1.295
+ $X2=2.62 $Y2=1.442
r99 49 77 6.71806 $w=2.27e-07 $l=1.25e-07 $layer=LI1_cond $X=2.62 $Y=1.295
+ $X2=2.62 $Y2=1.17
r100 48 59 8.19515 $w=2.23e-07 $l=1.6e-07 $layer=LI1_cond $X=2.622 $Y=0.925
+ $X2=2.622 $Y2=1.085
r101 47 48 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.622 $Y=0.555
+ $X2=2.622 $Y2=0.925
r102 47 61 6.40246 $w=2.23e-07 $l=1.25e-07 $layer=LI1_cond $X=2.622 $Y=0.555
+ $X2=2.622 $Y2=0.43
r103 39 41 34.3114 $w=2.18e-07 $l=6.55e-07 $layer=LI1_cond $X=3.515 $Y=1.085
+ $X2=3.515 $Y2=0.43
r104 36 51 2.79892 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2.78 $Y=2.035
+ $X2=2.642 $Y2=2.035
r105 35 46 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=3.505 $Y2=2.035
r106 35 36 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=2.78 $Y2=2.035
r107 34 77 2.43258 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.735 $Y=1.17
+ $X2=2.62 $Y2=1.17
r108 33 39 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.405 $Y=1.17
+ $X2=3.515 $Y2=1.085
r109 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.405 $Y=1.17
+ $X2=2.735 $Y2=1.17
r110 31 80 0.531045 $w=2.35e-07 $l=1.15e-07 $layer=LI1_cond $X=2.505 $Y=1.442
+ $X2=2.62 $Y2=1.442
r111 31 32 29.1789 $w=2.33e-07 $l=5.95e-07 $layer=LI1_cond $X=2.505 $Y=1.442
+ $X2=1.91 $Y2=1.442
r112 30 32 6.83402 $w=2.35e-07 $l=1.6225e-07 $layer=LI1_cond $X=1.802 $Y=1.325
+ $X2=1.91 $Y2=1.442
r113 29 44 4.14756 $w=2.2e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.802 $Y=1.04
+ $X2=1.797 $Y2=0.955
r114 29 30 15.2766 $w=2.13e-07 $l=2.85e-07 $layer=LI1_cond $X=1.802 $Y=1.04
+ $X2=1.802 $Y2=1.325
r115 25 44 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.797 $Y=0.87
+ $X2=1.797 $Y2=0.955
r116 25 27 22.5367 $w=2.23e-07 $l=4.4e-07 $layer=LI1_cond $X=1.797 $Y=0.87
+ $X2=1.797 $Y2=0.43
r117 23 44 2.28545 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.685 $Y=0.955
+ $X2=1.797 $Y2=0.955
r118 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.685 $Y=0.955
+ $X2=1.015 $Y2=0.955
r119 19 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.92 $Y=0.87
+ $X2=1.015 $Y2=0.955
r120 19 21 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=0.92 $Y=0.87
+ $X2=0.92 $Y2=0.43
r121 6 46 300 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=2 $X=3.36
+ $Y=1.835 $X2=3.5 $Y2=2.115
r122 5 51 300 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=2 $X=2.5
+ $Y=1.835 $X2=2.64 $Y2=2.115
r123 4 41 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=3.36
+ $Y=0.28 $X2=3.5 $Y2=0.43
r124 3 61 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=2.5
+ $Y=0.28 $X2=2.64 $Y2=0.43
r125 2 44 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.28 $X2=1.78 $Y2=0.975
r126 2 27 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.28 $X2=1.78 $Y2=0.43
r127 1 21 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=0.78
+ $Y=0.28 $X2=0.92 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_4%VGND 1 2 3 4 5 18 20 24 26 30 34 36 38 40 41
+ 42 48 53 59 62 65 69
r72 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r73 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r74 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r75 57 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r76 57 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r77 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r78 54 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.07
+ $Y2=0
r79 54 56 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.6
+ $Y2=0
r80 53 68 4.29113 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=4.057
+ $Y2=0
r81 53 56 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.6
+ $Y2=0
r82 52 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r83 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r84 49 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.21
+ $Y2=0
r85 49 51 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.64
+ $Y2=0
r86 48 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.07
+ $Y2=0
r87 48 51 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r88 46 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r89 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r90 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r91 42 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r92 42 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r93 40 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.325 $Y=0 $X2=0.24
+ $Y2=0
r94 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.325 $Y=0 $X2=0.49
+ $Y2=0
r95 36 68 3.22654 $w=3e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=4.057 $Y2=0
r96 36 38 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=3.945 $Y2=0.425
r97 32 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0
r98 32 34 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.425
r99 28 62 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r100 28 30 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.425
r101 27 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.35
+ $Y2=0
r102 26 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.08 $Y=0 $X2=2.21
+ $Y2=0
r103 26 27 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.08 $Y=0 $X2=1.515
+ $Y2=0
r104 22 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0
r105 22 24 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0.605
r106 21 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.655 $Y=0 $X2=0.49
+ $Y2=0
r107 20 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.35
+ $Y2=0
r108 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=0.655 $Y2=0
r109 16 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.49 $Y=0.085
+ $X2=0.49 $Y2=0
r110 16 18 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.49 $Y=0.085
+ $X2=0.49 $Y2=0.425
r111 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.79
+ $Y=0.28 $X2=3.93 $Y2=0.425
r112 4 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.93
+ $Y=0.28 $X2=3.07 $Y2=0.425
r113 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.07
+ $Y=0.28 $X2=2.21 $Y2=0.425
r114 2 24 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.21
+ $Y=0.28 $X2=1.35 $Y2=0.605
r115 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.365
+ $Y=0.28 $X2=0.49 $Y2=0.425
.ends

