* File: sky130_fd_sc_lp__ha_0.pxi.spice
* Created: Fri Aug 28 10:36:06 2020
* 
x_PM_SKY130_FD_SC_LP__HA_0%A_80_60# N_A_80_60#_M1013_s N_A_80_60#_M1008_d
+ N_A_80_60#_M1003_g N_A_80_60#_c_96_n N_A_80_60#_M1000_g N_A_80_60#_c_98_n
+ N_A_80_60#_c_92_n N_A_80_60#_c_99_n N_A_80_60#_c_143_p N_A_80_60#_c_121_p
+ N_A_80_60#_c_93_n N_A_80_60#_c_94_n N_A_80_60#_c_95_n
+ PM_SKY130_FD_SC_LP__HA_0%A_80_60#
x_PM_SKY130_FD_SC_LP__HA_0%A_204_315# N_A_204_315#_M1002_s N_A_204_315#_M1010_d
+ N_A_204_315#_M1008_g N_A_204_315#_M1013_g N_A_204_315#_c_169_n
+ N_A_204_315#_M1009_g N_A_204_315#_M1007_g N_A_204_315#_c_161_n
+ N_A_204_315#_c_172_n N_A_204_315#_c_162_n N_A_204_315#_c_163_n
+ N_A_204_315#_c_164_n N_A_204_315#_c_174_n N_A_204_315#_c_165_n
+ N_A_204_315#_c_166_n N_A_204_315#_c_167_n N_A_204_315#_c_223_p
+ N_A_204_315#_c_177_n PM_SKY130_FD_SC_LP__HA_0%A_204_315#
x_PM_SKY130_FD_SC_LP__HA_0%B N_B_M1004_g N_B_M1001_g N_B_c_269_n N_B_M1010_g
+ N_B_c_270_n N_B_M1002_g N_B_c_276_n N_B_c_277_n N_B_c_271_n B B B B
+ N_B_c_279_n PM_SKY130_FD_SC_LP__HA_0%B
x_PM_SKY130_FD_SC_LP__HA_0%A N_A_M1005_g N_A_M1012_g N_A_c_341_n N_A_c_342_n
+ N_A_c_343_n N_A_M1006_g N_A_M1011_g N_A_c_345_n N_A_c_346_n N_A_c_347_n A A
+ PM_SKY130_FD_SC_LP__HA_0%A
x_PM_SKY130_FD_SC_LP__HA_0%SUM N_SUM_M1003_s N_SUM_M1000_s SUM SUM SUM SUM SUM
+ SUM SUM SUM N_SUM_c_412_n PM_SKY130_FD_SC_LP__HA_0%SUM
x_PM_SKY130_FD_SC_LP__HA_0%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_M1006_d
+ N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n VPWR
+ N_VPWR_c_434_n N_VPWR_c_429_n N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n
+ PM_SKY130_FD_SC_LP__HA_0%VPWR
x_PM_SKY130_FD_SC_LP__HA_0%COUT N_COUT_M1007_d N_COUT_M1009_d N_COUT_c_487_n
+ COUT COUT COUT COUT COUT COUT PM_SKY130_FD_SC_LP__HA_0%COUT
x_PM_SKY130_FD_SC_LP__HA_0%VGND N_VGND_M1003_d N_VGND_M1004_d N_VGND_M1011_d
+ N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n VGND N_VGND_c_508_n
+ N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n
+ N_VGND_c_514_n N_VGND_c_515_n PM_SKY130_FD_SC_LP__HA_0%VGND
x_PM_SKY130_FD_SC_LP__HA_0%A_307_47# N_A_307_47#_M1013_d N_A_307_47#_M1012_d
+ N_A_307_47#_c_563_n N_A_307_47#_c_564_n N_A_307_47#_c_565_n
+ N_A_307_47#_c_566_n PM_SKY130_FD_SC_LP__HA_0%A_307_47#
cc_1 VNB N_A_80_60#_M1003_g 0.0679065f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_2 VNB N_A_80_60#_c_92_n 0.0215639f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.595
cc_3 VNB N_A_80_60#_c_93_n 0.0102745f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.76
cc_4 VNB N_A_80_60#_c_94_n 0.017278f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.93
cc_5 VNB N_A_80_60#_c_95_n 0.00514634f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.445
cc_6 VNB N_A_204_315#_M1013_g 0.0365827f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.265
cc_7 VNB N_A_204_315#_M1007_g 0.0470146f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.665
cc_8 VNB N_A_204_315#_c_161_n 0.0445585f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.76
cc_9 VNB N_A_204_315#_c_162_n 0.00212069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_204_315#_c_163_n 0.0190193f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.76
cc_11 VNB N_A_204_315#_c_164_n 0.0203447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_204_315#_c_165_n 0.00985709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_204_315#_c_166_n 0.0102696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_204_315#_c_167_n 0.0115222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1004_g 0.059621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_269_n 0.0172823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_270_n 0.0145099f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.775
cc_18 VNB N_B_c_271_n 0.0153426f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.665
cc_19 VNB N_A_M1005_g 0.0166018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_M1012_g 0.0323141f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.595
cc_21 VNB N_A_c_341_n 0.0469747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_342_n 0.0638621f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.772
cc_23 VNB N_A_c_343_n 0.0101948f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=2.088
cc_24 VNB N_A_M1011_g 0.0527461f $X=-0.19 $Y=-0.245 $X2=1.292 $Y2=2.265
cc_25 VNB N_A_c_345_n 0.0125506f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=2.665
cc_26 VNB N_A_c_346_n 0.0405241f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.665
cc_27 VNB N_A_c_347_n 0.00722665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB A 0.0071027f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.76
cc_29 VNB SUM 0.0380275f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.595
cc_30 VNB SUM 0.01137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB SUM 0.00996062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_429_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB COUT 0.040193f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=2.088
cc_34 VNB COUT 0.0117227f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.775
cc_35 VNB COUT 0.00909777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_505_n 0.0112618f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=2.088
cc_37 VNB N_VGND_c_506_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_507_n 0.0225765f $X=-0.19 $Y=-0.245 $X2=1.292 $Y2=2.265
cc_39 VNB N_VGND_c_508_n 0.0186851f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.665
cc_40 VNB N_VGND_c_509_n 0.0287764f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.93
cc_41 VNB N_VGND_c_510_n 0.0441158f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.445
cc_42 VNB N_VGND_c_511_n 0.019051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_512_n 0.273981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_513_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_514_n 0.00436611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_515_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_307_47#_c_563_n 0.00109763f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_48 VNB N_A_307_47#_c_564_n 0.0124893f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.772
cc_49 VNB N_A_307_47#_c_565_n 0.00970103f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=2.088
cc_50 VNB N_A_307_47#_c_566_n 0.00574098f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.775
cc_51 VPB N_A_80_60#_c_96_n 0.0231499f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=2.088
cc_52 VPB N_A_80_60#_M1000_g 0.0274229f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.775
cc_53 VPB N_A_80_60#_c_98_n 0.0187694f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=2.265
cc_54 VPB N_A_80_60#_c_99_n 0.00427276f $X=-0.19 $Y=1.655 $X2=1.292 $Y2=2.5
cc_55 VPB N_A_80_60#_c_93_n 0.00862593f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.76
cc_56 VPB N_A_80_60#_c_94_n 0.00917866f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.93
cc_57 VPB N_A_204_315#_M1008_g 0.0527055f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.64
cc_58 VPB N_A_204_315#_c_169_n 0.0214355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_204_315#_M1009_g 0.0276095f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.595
cc_60 VPB N_A_204_315#_c_161_n 0.015136f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.76
cc_61 VPB N_A_204_315#_c_172_n 0.0221184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_204_315#_c_164_n 0.010739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_204_315#_c_174_n 0.00421774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_204_315#_c_166_n 0.0170817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_204_315#_c_167_n 0.0105534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_204_315#_c_177_n 0.0016774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_B_M1004_g 0.0172004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_B_M1001_g 0.0224222f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.595
cc_69 VPB N_B_c_269_n 0.0127395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_B_M1010_g 0.0336825f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.265
cc_71 VPB N_B_c_276_n 0.0372221f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.61
cc_72 VPB N_B_c_277_n 0.00906445f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.595
cc_73 VPB B 0.0281489f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.76
cc_74 VPB N_B_c_279_n 0.0434388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_M1005_g 0.0618998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_M1006_g 0.0447073f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.775
cc_77 VPB N_A_c_347_n 0.00446172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB SUM 0.0422501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_SUM_c_412_n 0.0254399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_430_n 0.0138517f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.775
cc_81 VPB N_VPWR_c_431_n 0.0104911f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.61
cc_82 VPB N_VPWR_c_432_n 0.0175289f $X=-0.19 $Y=1.655 $X2=1.292 $Y2=2.5
cc_83 VPB N_VPWR_c_433_n 0.00583738f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=2.665
cc_84 VPB N_VPWR_c_434_n 0.0204631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_429_n 0.0808883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_436_n 0.0258599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_437_n 0.0383675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_438_n 0.0311109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_COUT_c_487_n 0.0329043f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.64
cc_90 VPB COUT 0.0413575f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.775
cc_91 N_A_80_60#_c_96_n N_A_204_315#_M1008_g 0.0162189f $X=0.577 $Y=2.088 $X2=0
+ $Y2=0
cc_92 N_A_80_60#_M1000_g N_A_204_315#_M1008_g 0.0113296f $X=0.57 $Y=2.775 $X2=0
+ $Y2=0
cc_93 N_A_80_60#_c_99_n N_A_204_315#_M1008_g 0.0056701f $X=1.292 $Y=2.5 $X2=0
+ $Y2=0
cc_94 N_A_80_60#_c_94_n N_A_204_315#_M1008_g 0.0288148f $X=1.06 $Y=1.93 $X2=0
+ $Y2=0
cc_95 N_A_80_60#_c_92_n N_A_204_315#_M1013_g 0.0103906f $X=1.06 $Y=1.595 $X2=0
+ $Y2=0
cc_96 N_A_80_60#_c_95_n N_A_204_315#_M1013_g 0.00287677f $X=1.225 $Y=0.445 $X2=0
+ $Y2=0
cc_97 N_A_80_60#_M1003_g N_A_204_315#_c_161_n 4.07045e-19 $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_98 N_A_80_60#_c_92_n N_A_204_315#_c_161_n 0.00374515f $X=1.06 $Y=1.595 $X2=0
+ $Y2=0
cc_99 N_A_80_60#_c_93_n N_A_204_315#_c_161_n 0.0162189f $X=0.59 $Y=1.76 $X2=0
+ $Y2=0
cc_100 N_A_80_60#_c_94_n N_A_204_315#_c_161_n 0.0107433f $X=1.06 $Y=1.93 $X2=0
+ $Y2=0
cc_101 N_A_80_60#_c_92_n N_A_204_315#_c_162_n 0.0375676f $X=1.06 $Y=1.595 $X2=0
+ $Y2=0
cc_102 N_A_80_60#_c_95_n N_A_204_315#_c_162_n 0.00173206f $X=1.225 $Y=0.445
+ $X2=0 $Y2=0
cc_103 N_A_80_60#_M1003_g N_A_204_315#_c_163_n 0.0051525f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_104 N_A_80_60#_c_92_n N_A_204_315#_c_163_n 0.00633295f $X=1.06 $Y=1.595 $X2=0
+ $Y2=0
cc_105 N_A_80_60#_c_95_n N_A_204_315#_c_163_n 0.0025507f $X=1.225 $Y=0.445 $X2=0
+ $Y2=0
cc_106 N_A_80_60#_c_92_n N_A_204_315#_c_174_n 0.00224642f $X=1.06 $Y=1.595 $X2=0
+ $Y2=0
cc_107 N_A_80_60#_c_94_n N_A_204_315#_c_174_n 0.0173502f $X=1.06 $Y=1.93 $X2=0
+ $Y2=0
cc_108 N_A_80_60#_c_94_n N_B_M1004_g 9.33427e-19 $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_109 N_A_80_60#_c_99_n N_B_M1001_g 0.00379795f $X=1.292 $Y=2.5 $X2=0 $Y2=0
cc_110 N_A_80_60#_c_121_p N_B_M1001_g 0.00618116f $X=1.675 $Y=2.665 $X2=0 $Y2=0
cc_111 N_A_80_60#_c_99_n N_B_c_276_n 2.84109e-19 $X=1.292 $Y=2.5 $X2=0 $Y2=0
cc_112 N_A_80_60#_c_121_p N_B_c_276_n 0.0102061f $X=1.675 $Y=2.665 $X2=0 $Y2=0
cc_113 N_A_80_60#_c_94_n N_B_c_276_n 0.00223102f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_114 N_A_80_60#_c_99_n B 0.00233983f $X=1.292 $Y=2.5 $X2=0 $Y2=0
cc_115 N_A_80_60#_c_121_p B 0.0151987f $X=1.675 $Y=2.665 $X2=0 $Y2=0
cc_116 N_A_80_60#_c_94_n B 0.0223274f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_117 N_A_80_60#_c_121_p N_A_M1005_g 9.24678e-19 $X=1.675 $Y=2.665 $X2=0 $Y2=0
cc_118 N_A_80_60#_M1003_g SUM 0.0235637f $X=0.475 $Y=0.64 $X2=0 $Y2=0
cc_119 N_A_80_60#_c_92_n SUM 0.0191761f $X=1.06 $Y=1.595 $X2=0 $Y2=0
cc_120 N_A_80_60#_M1003_g SUM 0.0219131f $X=0.475 $Y=0.64 $X2=0 $Y2=0
cc_121 N_A_80_60#_M1000_g SUM 0.00661592f $X=0.57 $Y=2.775 $X2=0 $Y2=0
cc_122 N_A_80_60#_c_92_n SUM 0.00504938f $X=1.06 $Y=1.595 $X2=0 $Y2=0
cc_123 N_A_80_60#_c_94_n SUM 0.0521358f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_124 N_A_80_60#_M1003_g SUM 0.00787801f $X=0.475 $Y=0.64 $X2=0 $Y2=0
cc_125 N_A_80_60#_M1000_g N_SUM_c_412_n 0.00517516f $X=0.57 $Y=2.775 $X2=0 $Y2=0
cc_126 N_A_80_60#_c_98_n N_SUM_c_412_n 0.00297513f $X=0.577 $Y=2.265 $X2=0 $Y2=0
cc_127 N_A_80_60#_M1000_g N_VPWR_c_430_n 0.0067959f $X=0.57 $Y=2.775 $X2=0 $Y2=0
cc_128 N_A_80_60#_c_98_n N_VPWR_c_430_n 6.57628e-19 $X=0.577 $Y=2.265 $X2=0
+ $Y2=0
cc_129 N_A_80_60#_c_99_n N_VPWR_c_430_n 0.00269941f $X=1.292 $Y=2.5 $X2=0 $Y2=0
cc_130 N_A_80_60#_c_94_n N_VPWR_c_430_n 0.0303203f $X=1.06 $Y=1.93 $X2=0 $Y2=0
cc_131 N_A_80_60#_M1000_g N_VPWR_c_429_n 0.0127355f $X=0.57 $Y=2.775 $X2=0 $Y2=0
cc_132 N_A_80_60#_c_143_p N_VPWR_c_429_n 0.00818208f $X=1.415 $Y=2.665 $X2=0
+ $Y2=0
cc_133 N_A_80_60#_c_121_p N_VPWR_c_429_n 0.0137563f $X=1.675 $Y=2.665 $X2=0
+ $Y2=0
cc_134 N_A_80_60#_M1000_g N_VPWR_c_436_n 0.00579312f $X=0.57 $Y=2.775 $X2=0
+ $Y2=0
cc_135 N_A_80_60#_c_143_p N_VPWR_c_437_n 0.00580142f $X=1.415 $Y=2.665 $X2=0
+ $Y2=0
cc_136 N_A_80_60#_c_121_p N_VPWR_c_437_n 0.0100549f $X=1.675 $Y=2.665 $X2=0
+ $Y2=0
cc_137 N_A_80_60#_c_121_p N_VPWR_c_438_n 0.0116388f $X=1.675 $Y=2.665 $X2=0
+ $Y2=0
cc_138 N_A_80_60#_M1003_g N_VGND_c_505_n 0.00471303f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_139 N_A_80_60#_c_92_n N_VGND_c_505_n 0.0146512f $X=1.06 $Y=1.595 $X2=0 $Y2=0
cc_140 N_A_80_60#_c_95_n N_VGND_c_505_n 0.0267632f $X=1.225 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_80_60#_M1003_g N_VGND_c_508_n 0.00510314f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_142 N_A_80_60#_c_95_n N_VGND_c_509_n 0.0223433f $X=1.225 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_80_60#_M1013_s N_VGND_c_512_n 0.00233781f $X=1.1 $Y=0.235 $X2=0 $Y2=0
cc_144 N_A_80_60#_M1003_g N_VGND_c_512_n 0.00526787f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_145 N_A_80_60#_c_95_n N_VGND_c_512_n 0.0155853f $X=1.225 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_80_60#_c_92_n N_A_307_47#_c_563_n 0.00327095f $X=1.06 $Y=1.595 $X2=0
+ $Y2=0
cc_147 N_A_80_60#_c_92_n N_A_307_47#_c_565_n 0.00769282f $X=1.06 $Y=1.595 $X2=0
+ $Y2=0
cc_148 N_A_204_315#_M1008_g N_B_M1004_g 0.00408518f $X=1.095 $Y=2.665 $X2=0
+ $Y2=0
cc_149 N_A_204_315#_M1013_g N_B_M1004_g 0.0247782f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_204_315#_c_162_n N_B_M1004_g 0.0023542f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A_204_315#_c_163_n N_B_M1004_g 0.0355704f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_152 N_A_204_315#_c_164_n N_B_M1004_g 0.0146193f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_153 N_A_204_315#_M1008_g N_B_M1001_g 0.00523505f $X=1.095 $Y=2.665 $X2=0
+ $Y2=0
cc_154 N_A_204_315#_c_165_n N_B_c_269_n 0.00867384f $X=3.115 $Y=0.885 $X2=0
+ $Y2=0
cc_155 N_A_204_315#_c_166_n N_B_c_269_n 0.0199115f $X=3.525 $Y=1.915 $X2=0 $Y2=0
cc_156 N_A_204_315#_c_177_n N_B_M1010_g 0.00449112f $X=3.48 $Y=2.5 $X2=0 $Y2=0
cc_157 N_A_204_315#_c_165_n N_B_c_270_n 0.0138973f $X=3.115 $Y=0.885 $X2=0 $Y2=0
cc_158 N_A_204_315#_M1008_g N_B_c_276_n 0.0142019f $X=1.095 $Y=2.665 $X2=0 $Y2=0
cc_159 N_A_204_315#_c_161_n N_B_c_276_n 0.00668537f $X=1.41 $Y=1.575 $X2=0 $Y2=0
cc_160 N_A_204_315#_c_164_n N_B_c_276_n 0.00173621f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_161 N_A_204_315#_c_174_n N_B_c_276_n 0.00318658f $X=1.575 $Y=1.65 $X2=0 $Y2=0
cc_162 N_A_204_315#_c_165_n N_B_c_271_n 0.0116157f $X=3.115 $Y=0.885 $X2=0 $Y2=0
cc_163 N_A_204_315#_M1008_g B 9.18308e-19 $X=1.095 $Y=2.665 $X2=0 $Y2=0
cc_164 N_A_204_315#_c_164_n B 0.106729f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_165 N_A_204_315#_c_166_n B 0.0517532f $X=3.525 $Y=1.915 $X2=0 $Y2=0
cc_166 N_A_204_315#_c_177_n B 0.00227967f $X=3.48 $Y=2.5 $X2=0 $Y2=0
cc_167 N_A_204_315#_c_164_n N_B_c_279_n 0.00315425f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_168 N_A_204_315#_c_166_n N_B_c_279_n 0.00370505f $X=3.525 $Y=1.915 $X2=0
+ $Y2=0
cc_169 N_A_204_315#_c_164_n N_A_M1005_g 0.0123593f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_170 N_A_204_315#_c_165_n N_A_M1005_g 0.00434699f $X=3.115 $Y=0.885 $X2=0
+ $Y2=0
cc_171 N_A_204_315#_c_165_n N_A_c_341_n 0.00997386f $X=3.115 $Y=0.885 $X2=0
+ $Y2=0
cc_172 N_A_204_315#_c_165_n N_A_c_342_n 0.00753117f $X=3.115 $Y=0.885 $X2=0
+ $Y2=0
cc_173 N_A_204_315#_M1009_g N_A_M1006_g 0.0111781f $X=4.205 $Y=2.775 $X2=0 $Y2=0
cc_174 N_A_204_315#_c_166_n N_A_M1006_g 0.0245314f $X=3.525 $Y=1.915 $X2=0 $Y2=0
cc_175 N_A_204_315#_c_167_n N_A_M1006_g 0.0259794f $X=4.17 $Y=1.76 $X2=0 $Y2=0
cc_176 N_A_204_315#_c_223_p N_A_M1006_g 0.00373622f $X=3.445 $Y=2.665 $X2=0
+ $Y2=0
cc_177 N_A_204_315#_c_177_n N_A_M1006_g 0.00531275f $X=3.48 $Y=2.5 $X2=0 $Y2=0
cc_178 N_A_204_315#_M1007_g N_A_M1011_g 0.0211017f $X=4.325 $Y=0.885 $X2=0 $Y2=0
cc_179 N_A_204_315#_c_165_n N_A_M1011_g 0.015803f $X=3.115 $Y=0.885 $X2=0 $Y2=0
cc_180 N_A_204_315#_c_164_n N_A_c_345_n 0.0142978f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_181 N_A_204_315#_c_166_n N_A_c_347_n 0.0172302f $X=3.525 $Y=1.915 $X2=0 $Y2=0
cc_182 N_A_204_315#_c_167_n N_A_c_347_n 0.00777551f $X=4.17 $Y=1.76 $X2=0 $Y2=0
cc_183 N_A_204_315#_c_162_n A 0.0139522f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_184 N_A_204_315#_c_164_n A 0.0585685f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_185 N_A_204_315#_c_165_n A 0.0245091f $X=3.115 $Y=0.885 $X2=0 $Y2=0
cc_186 N_A_204_315#_M1008_g N_VPWR_c_430_n 0.00447441f $X=1.095 $Y=2.665 $X2=0
+ $Y2=0
cc_187 N_A_204_315#_M1009_g N_VPWR_c_431_n 0.00654842f $X=4.205 $Y=2.775 $X2=0
+ $Y2=0
cc_188 N_A_204_315#_c_172_n N_VPWR_c_431_n 6.18483e-19 $X=4.202 $Y=2.265 $X2=0
+ $Y2=0
cc_189 N_A_204_315#_c_166_n N_VPWR_c_431_n 0.0280006f $X=3.525 $Y=1.915 $X2=0
+ $Y2=0
cc_190 N_A_204_315#_c_177_n N_VPWR_c_431_n 0.0148883f $X=3.48 $Y=2.5 $X2=0 $Y2=0
cc_191 N_A_204_315#_c_223_p N_VPWR_c_432_n 0.00587801f $X=3.445 $Y=2.665 $X2=0
+ $Y2=0
cc_192 N_A_204_315#_M1009_g N_VPWR_c_434_n 0.0054895f $X=4.205 $Y=2.775 $X2=0
+ $Y2=0
cc_193 N_A_204_315#_M1008_g N_VPWR_c_429_n 0.00519032f $X=1.095 $Y=2.665 $X2=0
+ $Y2=0
cc_194 N_A_204_315#_M1009_g N_VPWR_c_429_n 0.0120934f $X=4.205 $Y=2.775 $X2=0
+ $Y2=0
cc_195 N_A_204_315#_c_223_p N_VPWR_c_429_n 0.00850755f $X=3.445 $Y=2.665 $X2=0
+ $Y2=0
cc_196 N_A_204_315#_M1008_g N_VPWR_c_437_n 0.00517164f $X=1.095 $Y=2.665 $X2=0
+ $Y2=0
cc_197 N_A_204_315#_M1009_g N_COUT_c_487_n 0.00812388f $X=4.205 $Y=2.775 $X2=0
+ $Y2=0
cc_198 N_A_204_315#_c_172_n N_COUT_c_487_n 0.00572929f $X=4.202 $Y=2.265 $X2=0
+ $Y2=0
cc_199 N_A_204_315#_c_166_n N_COUT_c_487_n 7.57502e-19 $X=3.525 $Y=1.915 $X2=0
+ $Y2=0
cc_200 N_A_204_315#_M1007_g COUT 0.0183843f $X=4.325 $Y=0.885 $X2=0 $Y2=0
cc_201 N_A_204_315#_M1009_g COUT 0.00624328f $X=4.205 $Y=2.775 $X2=0 $Y2=0
cc_202 N_A_204_315#_M1007_g COUT 0.0256004f $X=4.325 $Y=0.885 $X2=0 $Y2=0
cc_203 N_A_204_315#_c_166_n COUT 0.0554433f $X=3.525 $Y=1.915 $X2=0 $Y2=0
cc_204 N_A_204_315#_M1007_g COUT 0.010019f $X=4.325 $Y=0.885 $X2=0 $Y2=0
cc_205 N_A_204_315#_M1013_g N_VGND_c_505_n 0.00235001f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_204_315#_M1013_g N_VGND_c_506_n 0.00126049f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_204_315#_M1007_g N_VGND_c_507_n 0.00474665f $X=4.325 $Y=0.885 $X2=0
+ $Y2=0
cc_208 N_A_204_315#_c_166_n N_VGND_c_507_n 0.0121579f $X=3.525 $Y=1.915 $X2=0
+ $Y2=0
cc_209 N_A_204_315#_c_167_n N_VGND_c_507_n 0.00116016f $X=4.17 $Y=1.76 $X2=0
+ $Y2=0
cc_210 N_A_204_315#_M1013_g N_VGND_c_509_n 0.00577974f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_204_315#_c_165_n N_VGND_c_510_n 0.00834492f $X=3.115 $Y=0.885 $X2=0
+ $Y2=0
cc_212 N_A_204_315#_M1007_g N_VGND_c_511_n 0.00291987f $X=4.325 $Y=0.885 $X2=0
+ $Y2=0
cc_213 N_A_204_315#_M1013_g N_VGND_c_512_n 0.0122227f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_214 N_A_204_315#_M1007_g N_VGND_c_512_n 0.0032212f $X=4.325 $Y=0.885 $X2=0
+ $Y2=0
cc_215 N_A_204_315#_c_165_n N_VGND_c_512_n 0.0145154f $X=3.115 $Y=0.885 $X2=0
+ $Y2=0
cc_216 N_A_204_315#_M1013_g N_A_307_47#_c_563_n 7.28977e-19 $X=1.46 $Y=0.445
+ $X2=0 $Y2=0
cc_217 N_A_204_315#_c_165_n N_A_307_47#_c_564_n 0.00971087f $X=3.115 $Y=0.885
+ $X2=0 $Y2=0
cc_218 N_A_204_315#_M1013_g N_A_307_47#_c_565_n 0.00229223f $X=1.46 $Y=0.445
+ $X2=0 $Y2=0
cc_219 N_A_204_315#_c_162_n N_A_307_47#_c_565_n 0.00123756f $X=1.41 $Y=1.22
+ $X2=0 $Y2=0
cc_220 N_A_204_315#_c_165_n A_687_135# 0.00164791f $X=3.115 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_221 N_B_c_277_n N_A_M1005_g 0.0521216f $X=1.89 $Y=2.13 $X2=0 $Y2=0
cc_222 B N_A_M1005_g 0.0254137f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_223 N_B_c_279_n N_A_M1005_g 0.00702332f $X=3.23 $Y=2 $X2=0 $Y2=0
cc_224 N_B_M1004_g N_A_M1012_g 0.0259333f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B_c_270_n N_A_c_341_n 0.0123912f $X=3.36 $Y=1.205 $X2=0 $Y2=0
cc_226 N_B_c_270_n N_A_c_342_n 0.00993587f $X=3.36 $Y=1.205 $X2=0 $Y2=0
cc_227 B N_A_M1006_g 3.58746e-19 $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_228 N_B_c_279_n N_A_M1006_g 0.022113f $X=3.23 $Y=2 $X2=0 $Y2=0
cc_229 N_B_c_269_n N_A_M1011_g 0.00639082f $X=3.23 $Y=1.835 $X2=0 $Y2=0
cc_230 N_B_c_270_n N_A_M1011_g 0.0477831f $X=3.36 $Y=1.205 $X2=0 $Y2=0
cc_231 N_B_M1004_g N_A_c_345_n 0.0521216f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_232 N_B_c_271_n N_A_c_346_n 0.00847467f $X=3.36 $Y=1.28 $X2=0 $Y2=0
cc_233 N_B_c_279_n N_A_c_346_n 2.10435e-19 $X=3.23 $Y=2 $X2=0 $Y2=0
cc_234 N_B_c_269_n N_A_c_347_n 0.022113f $X=3.23 $Y=1.835 $X2=0 $Y2=0
cc_235 N_B_M1004_g A 0.00423471f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_236 N_B_M1010_g N_VPWR_c_432_n 0.00429764f $X=3.23 $Y=2.665 $X2=0 $Y2=0
cc_237 N_B_M1001_g N_VPWR_c_429_n 0.00519032f $X=1.89 $Y=2.665 $X2=0 $Y2=0
cc_238 N_B_M1010_g N_VPWR_c_429_n 0.00432527f $X=3.23 $Y=2.665 $X2=0 $Y2=0
cc_239 N_B_M1001_g N_VPWR_c_437_n 0.00494981f $X=1.89 $Y=2.665 $X2=0 $Y2=0
cc_240 N_B_M1001_g N_VPWR_c_438_n 0.00178822f $X=1.89 $Y=2.665 $X2=0 $Y2=0
cc_241 N_B_M1010_g N_VPWR_c_438_n 0.0110263f $X=3.23 $Y=2.665 $X2=0 $Y2=0
cc_242 B N_VPWR_c_438_n 0.0599081f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_243 N_B_c_279_n N_VPWR_c_438_n 0.00146944f $X=3.23 $Y=2 $X2=0 $Y2=0
cc_244 N_B_M1004_g N_VGND_c_506_n 0.00878665f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_245 N_B_M1004_g N_VGND_c_509_n 0.00362954f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_246 N_B_M1004_g N_VGND_c_512_n 0.00438424f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_247 N_B_c_270_n N_VGND_c_512_n 8.49626e-19 $X=3.36 $Y=1.205 $X2=0 $Y2=0
cc_248 N_B_M1004_g N_A_307_47#_c_563_n 8.69692e-19 $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_249 N_B_M1004_g N_A_307_47#_c_564_n 0.0160455f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A_M1006_g N_VPWR_c_431_n 0.00261047f $X=3.66 $Y=2.665 $X2=0 $Y2=0
cc_251 N_A_M1006_g N_VPWR_c_432_n 0.00495853f $X=3.66 $Y=2.665 $X2=0 $Y2=0
cc_252 N_A_M1005_g N_VPWR_c_429_n 0.00432527f $X=2.28 $Y=2.665 $X2=0 $Y2=0
cc_253 N_A_M1006_g N_VPWR_c_429_n 0.00519032f $X=3.66 $Y=2.665 $X2=0 $Y2=0
cc_254 N_A_M1005_g N_VPWR_c_437_n 0.00429764f $X=2.28 $Y=2.665 $X2=0 $Y2=0
cc_255 N_A_M1005_g N_VPWR_c_438_n 0.0132516f $X=2.28 $Y=2.665 $X2=0 $Y2=0
cc_256 N_A_M1006_g N_VPWR_c_438_n 4.62937e-19 $X=3.66 $Y=2.665 $X2=0 $Y2=0
cc_257 N_A_M1011_g COUT 0.00182801f $X=3.72 $Y=0.885 $X2=0 $Y2=0
cc_258 N_A_M1012_g N_VGND_c_506_n 0.00885153f $X=2.32 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_c_343_n N_VGND_c_506_n 7.11401e-19 $X=2.885 $Y=0.26 $X2=0 $Y2=0
cc_260 N_A_c_342_n N_VGND_c_507_n 0.0241653f $X=3.645 $Y=0.26 $X2=0 $Y2=0
cc_261 N_A_M1012_g N_VGND_c_510_n 0.00362954f $X=2.32 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_c_343_n N_VGND_c_510_n 0.0286185f $X=2.885 $Y=0.26 $X2=0 $Y2=0
cc_263 N_A_M1012_g N_VGND_c_512_n 0.0052251f $X=2.32 $Y=0.445 $X2=0 $Y2=0
cc_264 N_A_c_342_n N_VGND_c_512_n 0.0371589f $X=3.645 $Y=0.26 $X2=0 $Y2=0
cc_265 N_A_c_343_n N_VGND_c_512_n 0.00978654f $X=2.885 $Y=0.26 $X2=0 $Y2=0
cc_266 N_A_M1012_g N_A_307_47#_c_564_n 0.0117824f $X=2.32 $Y=0.445 $X2=0 $Y2=0
cc_267 N_A_c_341_n N_A_307_47#_c_564_n 0.00216164f $X=2.81 $Y=1.055 $X2=0 $Y2=0
cc_268 N_A_c_345_n N_A_307_47#_c_564_n 0.00105442f $X=2.3 $Y=1.22 $X2=0 $Y2=0
cc_269 N_A_c_346_n N_A_307_47#_c_564_n 0.00370833f $X=2.735 $Y=1.22 $X2=0 $Y2=0
cc_270 A N_A_307_47#_c_564_n 0.0557912f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_271 N_A_M1012_g N_A_307_47#_c_566_n 9.56419e-19 $X=2.32 $Y=0.445 $X2=0 $Y2=0
cc_272 N_A_c_343_n N_A_307_47#_c_566_n 0.0119937f $X=2.885 $Y=0.26 $X2=0 $Y2=0
cc_273 SUM N_VPWR_c_430_n 0.00184505f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_274 N_SUM_M1000_s N_VPWR_c_429_n 0.00231914f $X=0.21 $Y=2.455 $X2=0 $Y2=0
cc_275 N_SUM_c_412_n N_VPWR_c_429_n 0.0155486f $X=0.335 $Y=2.6 $X2=0 $Y2=0
cc_276 N_SUM_c_412_n N_VPWR_c_436_n 0.0263719f $X=0.335 $Y=2.6 $X2=0 $Y2=0
cc_277 SUM N_VGND_c_505_n 0.0174689f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_278 SUM N_VGND_c_508_n 0.0127604f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_279 SUM N_VGND_c_512_n 0.011834f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_280 N_VPWR_c_429_n N_COUT_M1009_d 0.00215158f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_281 N_VPWR_c_431_n N_COUT_c_487_n 0.026047f $X=3.875 $Y=2.6 $X2=0 $Y2=0
cc_282 N_VPWR_c_434_n N_COUT_c_487_n 0.0303285f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_429_n N_COUT_c_487_n 0.017612f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_284 COUT N_VGND_c_507_n 0.0538996f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_285 COUT N_VGND_c_511_n 0.0145152f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_286 COUT N_VGND_c_512_n 0.0130211f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_287 N_VGND_c_512_n N_A_307_47#_M1013_d 0.00336966f $X=4.56 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_288 N_VGND_c_512_n N_A_307_47#_M1012_d 0.00234495f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_509_n N_A_307_47#_c_563_n 0.0112671f $X=1.94 $Y=0 $X2=0 $Y2=0
cc_290 N_VGND_c_512_n N_A_307_47#_c_563_n 0.0079618f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_291 N_VGND_c_506_n N_A_307_47#_c_564_n 0.0205535f $X=2.105 $Y=0.445 $X2=0
+ $Y2=0
cc_292 N_VGND_c_509_n N_A_307_47#_c_564_n 0.00238864f $X=1.94 $Y=0 $X2=0 $Y2=0
cc_293 N_VGND_c_510_n N_A_307_47#_c_564_n 0.00238864f $X=3.855 $Y=0 $X2=0 $Y2=0
cc_294 N_VGND_c_512_n N_A_307_47#_c_564_n 0.00919325f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_295 N_VGND_c_510_n N_A_307_47#_c_566_n 0.015222f $X=3.855 $Y=0 $X2=0 $Y2=0
cc_296 N_VGND_c_512_n N_A_307_47#_c_566_n 0.00987569f $X=4.56 $Y=0 $X2=0 $Y2=0
