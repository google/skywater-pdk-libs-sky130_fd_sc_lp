* File: sky130_fd_sc_lp__a22oi_lp.pex.spice
* Created: Wed Sep  2 09:23:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22OI_LP%B2 3 7 11 12 13 16
c37 3 0 8.40218e-20 $X=0.73 $Y=2.545
r38 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.24 $X2=0.69 $Y2=1.24
r39 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.69 $Y=1.58
+ $X2=0.69 $Y2=1.24
r40 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.69 $Y=1.58
+ $X2=0.69 $Y2=1.745
r41 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.69 $Y=1.075
+ $X2=0.69 $Y2=1.24
r42 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.78 $Y=0.445
+ $X2=0.78 $Y2=1.075
r43 3 12 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=0.73 $Y=2.545 $X2=0.73
+ $Y2=1.745
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_LP%B1 3 7 11 12 13 16
c44 12 0 6.99559e-20 $X=1.23 $Y=1.745
r45 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=1.24 $X2=1.23 $Y2=1.24
r46 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.23 $Y=1.58
+ $X2=1.23 $Y2=1.24
r47 11 12 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.58
+ $X2=1.23 $Y2=1.745
r48 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.075
+ $X2=1.23 $Y2=1.24
r49 7 12 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=1.26 $Y=2.545 $X2=1.26
+ $Y2=1.745
r50 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.17 $Y=0.445
+ $X2=1.17 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_LP%A1 3 7 11 12 13 16 17
c41 7 0 8.40218e-20 $X=1.79 $Y=2.545
r42 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.8 $Y=1.24
+ $X2=1.8 $Y2=1.24
r43 13 17 2.14223 $w=6.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.68 $Y=1.41 $X2=1.8
+ $Y2=1.41
r44 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.8 $Y=1.58 $X2=1.8
+ $Y2=1.24
r45 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.58 $X2=1.8
+ $Y2=1.745
r46 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.075
+ $X2=1.8 $Y2=1.24
r47 7 12 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=1.79 $Y=2.545 $X2=1.79
+ $Y2=1.745
r48 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.71 $Y=0.445
+ $X2=1.71 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_LP%A2 3 7 9 12
c27 12 0 2.50695e-20 $X=2.495 $Y=1.02
c28 7 0 4.84015e-20 $X=2.33 $Y=2.545
r29 12 15 72.9334 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=2.432 $Y=1.02
+ $X2=2.432 $Y2=1.525
r30 12 14 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=2.432 $Y=1.02
+ $X2=2.432 $Y2=0.855
r31 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.495
+ $Y=1.02 $X2=2.495 $Y2=1.02
r32 9 13 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.19
+ $X2=2.495 $Y2=1.19
r33 7 15 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.33 $Y=2.545
+ $X2=2.33 $Y2=1.525
r34 3 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.28 $Y=0.445
+ $X2=2.28 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_LP%A_64_409# 1 2 3 12 14 15 17 19 20 21 24
c53 21 0 1.53978e-19 $X=1.69 $Y=2.01
c54 17 0 4.84015e-20 $X=1.525 $Y=2.895
r55 24 26 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.595 $Y=2.19
+ $X2=2.595 $Y2=2.9
r56 22 24 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.595 $Y=2.095
+ $X2=2.595 $Y2=2.19
r57 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.43 $Y=2.01
+ $X2=2.595 $Y2=2.095
r58 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.43 $Y=2.01
+ $X2=1.69 $Y2=2.01
r59 17 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=2.895
+ $X2=1.525 $Y2=2.98
r60 17 19 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.525 $Y=2.895
+ $X2=1.525 $Y2=2.19
r61 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.525 $Y=2.095
+ $X2=1.69 $Y2=2.01
r62 16 19 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.525 $Y=2.095
+ $X2=1.525 $Y2=2.19
r63 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=2.98
+ $X2=1.525 $Y2=2.98
r64 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.36 $Y=2.98
+ $X2=0.63 $Y2=2.98
r65 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.465 $Y=2.895
+ $X2=0.63 $Y2=2.98
r66 10 12 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.465 $Y=2.895
+ $X2=0.465 $Y2=2.44
r67 3 26 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=2.045 $X2=2.595 $Y2=2.9
r68 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=2.045 $X2=2.595 $Y2=2.19
r69 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=2.045 $X2=1.525 $Y2=2.9
r70 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=2.045 $X2=1.525 $Y2=2.19
r71 1 12 300 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=2 $X=0.32
+ $Y=2.045 $X2=0.465 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_LP%Y 1 2 7 9 10 13 17 20 21 22 27 29
c48 9 0 8.40218e-20 $X=0.83 $Y=2.01
r49 27 29 1.57151 $w=2.18e-07 $l=3e-08 $layer=LI1_cond $X=0.235 $Y=0.895
+ $X2=0.235 $Y2=0.925
r50 21 22 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r51 20 27 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=0.81
+ $X2=0.235 $Y2=0.895
r52 20 21 17.9676 $w=2.18e-07 $l=3.43e-07 $layer=LI1_cond $X=0.235 $Y=0.952
+ $X2=0.235 $Y2=1.295
r53 20 29 1.41436 $w=2.18e-07 $l=2.7e-08 $layer=LI1_cond $X=0.235 $Y=0.952
+ $X2=0.235 $Y2=0.925
r54 19 22 13.6198 $w=2.18e-07 $l=2.6e-07 $layer=LI1_cond $X=0.235 $Y=1.925
+ $X2=0.235 $Y2=1.665
r55 15 17 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.385 $Y=0.725
+ $X2=1.385 $Y2=0.47
r56 11 13 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.995 $Y=2.095
+ $X2=0.995 $Y2=2.19
r57 10 19 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.345 $Y=2.01
+ $X2=0.235 $Y2=1.925
r58 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.83 $Y=2.01
+ $X2=0.995 $Y2=2.095
r59 9 10 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.83 $Y=2.01
+ $X2=0.345 $Y2=2.01
r60 8 20 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.345 $Y=0.81
+ $X2=0.235 $Y2=0.81
r61 7 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.22 $Y=0.81
+ $X2=1.385 $Y2=0.725
r62 7 8 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.22 $Y=0.81
+ $X2=0.345 $Y2=0.81
r63 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.855
+ $Y=2.045 $X2=0.995 $Y2=2.19
r64 1 17 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.245
+ $Y=0.235 $X2=1.385 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_LP%VPWR 1 6 9 10 11 21 22
r30 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r33 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 11 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 9 18 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=3.33 $X2=1.68
+ $Y2=3.33
r38 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=2.055 $Y2=3.33
r39 8 21 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.22 $Y=3.33 $X2=2.64
+ $Y2=3.33
r40 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.055 $Y2=3.33
r41 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=3.33
r42 4 6 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=2.44
r43 1 6 300 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=2 $X=1.915
+ $Y=2.045 $X2=2.055 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_LP%VGND 1 2 9 11 13 15 17 22 28 32
c34 32 0 2.50695e-20 $X=2.64 $Y=0
r35 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r36 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r38 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0 $X2=0.565
+ $Y2=0
r40 23 25 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=0.73 $Y=0 $X2=2.16
+ $Y2=0
r41 22 31 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.605
+ $Y2=0
r42 22 25 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.16
+ $Y2=0
r43 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r44 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.565
+ $Y2=0
r46 17 19 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.24
+ $Y2=0
r47 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r48 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r49 11 31 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.495 $Y=0.085
+ $X2=2.605 $Y2=0
r50 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.495 $Y=0.085
+ $X2=2.495 $Y2=0.445
r51 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.565 $Y=0.085
+ $X2=0.565 $Y2=0
r52 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.565 $Y=0.085
+ $X2=0.565 $Y2=0.38
r53 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.495 $Y2=0.445
r54 1 9 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.42
+ $Y=0.235 $X2=0.565 $Y2=0.38
.ends

