# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2bb2o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a2bb2o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245000 1.065000 5.040000 1.235000 ;
        RECT 3.245000 1.235000 3.575000 1.435000 ;
        RECT 4.475000 1.235000 5.040000 1.515000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.415000 4.295000 1.750000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.240000 1.345000 0.715000 1.645000 ;
        RECT 0.545000 1.645000 0.715000 1.950000 ;
        RECT 0.545000 1.950000 1.635000 2.120000 ;
        RECT 1.465000 1.405000 1.970000 1.645000 ;
        RECT 1.465000 1.645000 1.635000 1.950000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895000 1.405000 1.295000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.188600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.475000 0.255000 5.705000 1.065000 ;
        RECT 5.475000 1.065000 7.045000 1.235000 ;
        RECT 5.550000 1.755000 7.045000 1.925000 ;
        RECT 5.550000 1.925000 5.740000 3.075000 ;
        RECT 6.375000 0.255000 6.565000 1.065000 ;
        RECT 6.410000 1.925000 6.630000 3.075000 ;
        RECT 6.875000 1.235000 7.045000 1.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.095000  1.815000 0.375000 2.290000 ;
      RECT 0.095000  2.290000 2.175000 2.460000 ;
      RECT 0.095000  2.460000 0.375000 3.075000 ;
      RECT 0.115000  0.085000 0.400000 1.095000 ;
      RECT 0.545000  2.630000 0.875000 3.245000 ;
      RECT 0.570000  0.255000 1.735000 0.425000 ;
      RECT 0.570000  0.425000 0.850000 1.095000 ;
      RECT 1.020000  0.595000 1.235000 1.065000 ;
      RECT 1.020000  1.065000 2.565000 1.235000 ;
      RECT 1.045000  2.460000 1.255000 3.075000 ;
      RECT 1.405000  0.425000 1.735000 0.895000 ;
      RECT 1.425000  2.630000 1.755000 3.245000 ;
      RECT 1.905000  0.085000 2.185000 0.895000 ;
      RECT 1.935000  1.815000 2.175000 2.290000 ;
      RECT 1.935000  2.460000 2.175000 2.905000 ;
      RECT 1.935000  2.905000 3.065000 3.075000 ;
      RECT 2.345000  1.235000 2.565000 2.100000 ;
      RECT 2.345000  2.100000 3.405000 2.270000 ;
      RECT 2.345000  2.270000 2.565000 2.735000 ;
      RECT 2.365000  0.255000 2.565000 1.065000 ;
      RECT 2.735000  0.085000 3.405000 0.555000 ;
      RECT 2.735000  2.440000 3.065000 2.905000 ;
      RECT 2.755000  0.725000 4.855000 0.895000 ;
      RECT 2.755000  0.895000 2.925000 1.760000 ;
      RECT 2.755000  1.760000 3.745000 1.930000 ;
      RECT 3.235000  2.270000 3.405000 2.310000 ;
      RECT 3.235000  2.310000 5.380000 2.480000 ;
      RECT 3.255000  2.650000 3.585000 3.245000 ;
      RECT 3.575000  0.255000 3.835000 0.725000 ;
      RECT 3.575000  1.930000 4.445000 2.140000 ;
      RECT 3.755000  2.670000 4.850000 3.000000 ;
      RECT 4.015000  0.085000 4.345000 0.555000 ;
      RECT 4.525000  0.255000 4.855000 0.725000 ;
      RECT 5.020000  2.650000 5.350000 3.245000 ;
      RECT 5.025000  0.085000 5.305000 0.885000 ;
      RECT 5.210000  1.405000 6.695000 1.585000 ;
      RECT 5.210000  1.585000 5.380000 2.310000 ;
      RECT 5.875000  0.085000 6.205000 0.865000 ;
      RECT 5.910000  2.095000 6.240000 3.245000 ;
      RECT 6.735000  0.085000 7.065000 0.895000 ;
      RECT 6.800000  2.095000 7.100000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__a2bb2o_4
END LIBRARY
