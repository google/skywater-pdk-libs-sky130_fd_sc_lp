* File: sky130_fd_sc_lp__fa_1.pex.spice
* Created: Wed Sep  2 09:53:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FA_1%A_80_27# 1 2 9 12 16 20 23 24 25 28 34 35 38 39
+ 42 43 47 49
c142 47 0 1.62762e-19 $X=1.842 $Y=1.61
c143 20 0 9.76611e-20 $X=5.555 $Y=0.835
c144 16 0 5.8378e-20 $X=5.515 $Y=2.265
r145 42 45 4.17264 $w=2.88e-07 $l=1.05e-07 $layer=LI1_cond $X=1.775 $Y=2.385
+ $X2=1.775 $Y2=2.49
r146 42 43 4.07689 $w=2.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=2.385
+ $X2=1.775 $Y2=2.3
r147 39 50 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.38
+ $X2=0.597 $Y2=1.545
r148 39 49 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.38
+ $X2=0.597 $Y2=1.215
r149 38 41 7.40102 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.665 $Y=1.38
+ $X2=0.665 $Y2=1.545
r150 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.38 $X2=0.63 $Y2=1.38
r151 35 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.61
+ $X2=5.535 $Y2=1.775
r152 35 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.61
+ $X2=5.535 $Y2=1.445
r153 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.535
+ $Y=1.61 $X2=5.535 $Y2=1.61
r154 32 47 2.79892 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.985 $Y=1.61
+ $X2=1.842 $Y2=1.61
r155 32 34 231.604 $w=1.68e-07 $l=3.55e-06 $layer=LI1_cond $X=1.985 $Y=1.61
+ $X2=5.535 $Y2=1.61
r156 30 47 3.67481 $w=2.52e-07 $l=9.97246e-08 $layer=LI1_cond $X=1.81 $Y=1.695
+ $X2=1.842 $Y2=1.61
r157 30 43 31.6922 $w=2.18e-07 $l=6.05e-07 $layer=LI1_cond $X=1.81 $Y=1.695
+ $X2=1.81 $Y2=2.3
r158 26 47 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=1.842 $Y=1.525
+ $X2=1.842 $Y2=1.61
r159 26 28 25.4751 $w=2.83e-07 $l=6.3e-07 $layer=LI1_cond $X=1.842 $Y=1.525
+ $X2=1.842 $Y2=0.895
r160 24 42 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.63 $Y=2.385
+ $X2=1.775 $Y2=2.385
r161 24 25 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.63 $Y=2.385
+ $X2=0.795 $Y2=2.385
r162 23 25 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.675 $Y=2.3
+ $X2=0.795 $Y2=2.385
r163 23 41 36.2539 $w=2.38e-07 $l=7.55e-07 $layer=LI1_cond $X=0.675 $Y=2.3
+ $X2=0.675 $Y2=1.545
r164 20 52 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.555 $Y=0.835
+ $X2=5.555 $Y2=1.445
r165 16 53 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.515 $Y=2.265
+ $X2=5.515 $Y2=1.775
r166 12 50 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.485 $Y=2.465
+ $X2=0.485 $Y2=1.545
r167 9 49 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.685
+ $X2=0.475 $Y2=1.215
r168 2 45 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=2.285 $X2=1.795 $Y2=2.49
r169 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.685 $X2=1.865 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%A 3 7 11 15 20 21 22 25 30 33 37 41 42 43 44 45
+ 46 51 54 57 58 60 61 65 66
c211 60 0 1.03908e-19 $X=1.17 $Y=1.46
c212 58 0 3.79636e-21 $X=7.035 $Y=1.35
c213 46 0 9.79433e-20 $X=2.785 $Y=2.035
c214 3 0 5.88543e-20 $X=1.08 $Y=2.495
r215 65 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.53 $Y=1.96
+ $X2=2.53 $Y2=2.125
r216 65 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.53 $Y=1.96
+ $X2=2.53 $Y2=1.795
r217 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.96 $X2=2.53 $Y2=1.96
r218 61 72 19.4898 $w=3.38e-07 $l=5.75e-07 $layer=LI1_cond $X=1.175 $Y=1.46
+ $X2=1.175 $Y2=2.035
r219 60 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.46
+ $X2=1.17 $Y2=1.625
r220 60 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.46
+ $X2=1.17 $Y2=1.295
r221 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.46 $X2=1.17 $Y2=1.46
r222 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.035
+ $Y=1.35 $X2=7.035 $Y2=1.35
r223 54 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r224 52 58 26.3141 $w=2.98e-07 $l=6.85e-07 $layer=LI1_cond $X=6.97 $Y=2.035
+ $X2=6.97 $Y2=1.35
r225 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=2.035
r226 48 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=2.035
+ $X2=2.64 $Y2=2.035
r227 46 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=2.035
+ $X2=2.64 $Y2=2.035
r228 45 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=6.96 $Y2=2.035
r229 45 46 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=2.785 $Y2=2.035
r230 44 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r231 43 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=2.035
+ $X2=2.64 $Y2=2.035
r232 43 44 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=2.495 $Y=2.035
+ $X2=1.345 $Y2=2.035
r233 41 57 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.035 $Y=1.69
+ $X2=7.035 $Y2=1.35
r234 41 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.035 $Y=1.69
+ $X2=7.035 $Y2=1.855
r235 40 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.035 $Y=1.185
+ $X2=7.035 $Y2=1.35
r236 35 37 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.895 $Y=1.195
+ $X2=5.085 $Y2=1.195
r237 33 42 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=6.945 $Y=2.265
+ $X2=6.945 $Y2=1.855
r238 30 40 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.945 $Y=0.835
+ $X2=6.945 $Y2=1.185
r239 27 30 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.945 $Y=0.255
+ $X2=6.945 $Y2=0.835
r240 23 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.085 $Y=1.27
+ $X2=5.085 $Y2=1.195
r241 23 25 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=5.085 $Y=1.27
+ $X2=5.085 $Y2=2.265
r242 21 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.87 $Y=0.18
+ $X2=6.945 $Y2=0.255
r243 21 22 974.255 $w=1.5e-07 $l=1.9e-06 $layer=POLY_cond $X=6.87 $Y=0.18
+ $X2=4.97 $Y2=0.18
r244 18 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.895 $Y=1.12
+ $X2=4.895 $Y2=1.195
r245 18 20 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.895 $Y=1.12
+ $X2=4.895 $Y2=0.625
r246 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.895 $Y=0.255
+ $X2=4.97 $Y2=0.18
r247 17 20 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.895 $Y=0.255
+ $X2=4.895 $Y2=0.625
r248 15 67 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.51 $Y=0.895
+ $X2=2.51 $Y2=1.795
r249 11 68 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.44 $Y=2.495
+ $X2=2.44 $Y2=2.125
r250 7 62 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.26 $Y=0.895 $X2=1.26
+ $Y2=1.295
r251 3 63 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.08 $Y=2.495
+ $X2=1.08 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%B 3 7 8 9 13 16 18 20 23 26 29 30 32 35 38 41
+ 42 43 46 49 50 51 52 57 61 63 71 76
c167 57 0 9.48662e-20 $X=5.495 $Y=1.27
c168 50 0 1.4009e-19 $X=6.465 $Y=1.66
c169 30 0 1.12751e-19 $X=4.195 $Y=1.98
c170 7 0 1.16441e-19 $X=1.65 $Y=0.895
r171 76 77 9.43864 $w=3.83e-07 $l=7.5e-08 $layer=POLY_cond $X=4.015 $Y=1.23
+ $X2=4.09 $Y2=1.23
r172 63 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.465
+ $Y=1.32 $X2=6.465 $Y2=1.32
r173 61 63 8.69026 $w=6.38e-07 $l=4.65e-07 $layer=LI1_cond $X=6 $Y=1.505
+ $X2=6.465 $Y2=1.505
r174 60 76 1.88773 $w=3.83e-07 $l=1.5e-08 $layer=POLY_cond $X=4 $Y=1.23
+ $X2=4.015 $Y2=1.23
r175 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4 $Y=1.26
+ $X2=4 $Y2=1.26
r176 57 61 16.6933 $w=3.13e-07 $l=4.2e-07 $layer=LI1_cond $X=5.495 $Y=1.27
+ $X2=5.915 $Y2=1.27
r177 57 59 93.7662 $w=1.95e-07 $l=1.51733e-06 $layer=LI1_cond $X=5.495 $Y=1.27
+ $X2=4 $Y2=1.225
r178 55 60 48.4517 $w=3.83e-07 $l=3.85e-07 $layer=POLY_cond $X=3.615 $Y=1.23
+ $X2=4 $Y2=1.23
r179 55 73 11.3264 $w=3.83e-07 $l=9e-08 $layer=POLY_cond $X=3.615 $Y=1.23
+ $X2=3.525 $Y2=1.23
r180 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.26 $X2=3.615 $Y2=1.26
r181 52 59 9.93987 $w=2.6e-07 $l=1.95e-07 $layer=LI1_cond $X=3.805 $Y=1.225
+ $X2=4 $Y2=1.225
r182 52 54 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=1.225
+ $X2=3.615 $Y2=1.225
r183 50 71 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.465 $Y=1.66
+ $X2=6.465 $Y2=1.32
r184 50 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=1.66
+ $X2=6.465 $Y2=1.825
r185 49 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=1.155
+ $X2=6.465 $Y2=1.32
r186 44 46 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=4.09 $Y=1.905
+ $X2=4.195 $Y2=1.905
r187 40 41 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.615 $Y=2.06
+ $X2=1.615 $Y2=2.21
r188 38 51 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.375 $Y=2.265
+ $X2=6.375 $Y2=1.825
r189 35 49 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.375 $Y=0.835
+ $X2=6.375 $Y2=1.155
r190 30 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=1.98
+ $X2=4.195 $Y2=1.905
r191 30 32 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.195 $Y=1.98
+ $X2=4.195 $Y2=2.265
r192 29 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.09 $Y=1.83
+ $X2=4.09 $Y2=1.905
r193 28 77 24.8035 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.09 $Y=1.425
+ $X2=4.09 $Y2=1.23
r194 28 29 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.09 $Y=1.425
+ $X2=4.09 $Y2=1.83
r195 24 76 24.8035 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.015 $Y=1.035
+ $X2=4.015 $Y2=1.23
r196 24 26 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.015 $Y=1.035
+ $X2=4.015 $Y2=0.625
r197 23 73 24.8035 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.525 $Y=1.035
+ $X2=3.525 $Y2=1.23
r198 22 23 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=3.525 $Y=0.315
+ $X2=3.525 $Y2=1.035
r199 21 43 5.30422 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.105 $Y=1.35
+ $X2=2.985 $Y2=1.35
r200 20 73 27.9434 $w=3.83e-07 $l=1.52971e-07 $layer=POLY_cond $X=3.45 $Y=1.35
+ $X2=3.525 $Y2=1.23
r201 20 21 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=3.45 $Y=1.35
+ $X2=3.105 $Y2=1.35
r202 19 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=0.24
+ $X2=2.94 $Y2=0.24
r203 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.45 $Y=0.24
+ $X2=3.525 $Y2=0.315
r204 18 19 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.45 $Y=0.24
+ $X2=3.015 $Y2=0.24
r205 14 43 20.4101 $w=1.5e-07 $l=9.48683e-08 $layer=POLY_cond $X=3.03 $Y=1.425
+ $X2=2.985 $Y2=1.35
r206 14 16 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=3.03 $Y=1.425
+ $X2=3.03 $Y2=2.495
r207 11 43 20.4101 $w=1.5e-07 $l=9.48683e-08 $layer=POLY_cond $X=2.94 $Y=1.275
+ $X2=2.985 $Y2=1.35
r208 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.94 $Y=1.275
+ $X2=2.94 $Y2=0.895
r209 10 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=0.315
+ $X2=2.94 $Y2=0.24
r210 10 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.94 $Y=0.315
+ $X2=2.94 $Y2=0.895
r211 8 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=0.24
+ $X2=2.94 $Y2=0.24
r212 8 9 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.865 $Y=0.24
+ $X2=1.725 $Y2=0.24
r213 7 40 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=1.65 $Y=0.895
+ $X2=1.65 $Y2=2.06
r214 4 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.65 $Y=0.315
+ $X2=1.725 $Y2=0.24
r215 4 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.65 $Y=0.315
+ $X2=1.65 $Y2=0.895
r216 3 41 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.58 $Y=2.495
+ $X2=1.58 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%CIN 4 7 9 10 12 13 17 22 23 27 30 32 33 38 40
+ 43 45 48 49
c132 32 0 9.79433e-20 $X=2.045 $Y=2.21
c133 27 0 9.48662e-20 $X=5.985 $Y=0.835
r134 48 49 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.61 $Y=2.405
+ $X2=3.61 $Y2=2.775
r135 46 48 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=3.61 $Y=2.12
+ $X2=3.61 $Y2=2.405
r136 45 46 1.87632 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=3.61 $Y=1.992
+ $X2=3.61 $Y2=2.12
r137 43 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.96
+ $X2=3.53 $Y2=2.125
r138 42 45 3.61551 $w=2.53e-07 $l=8e-08 $layer=LI1_cond $X=3.53 $Y=1.992
+ $X2=3.61 $Y2=1.992
r139 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.53
+ $Y=1.96 $X2=3.53 $Y2=1.96
r140 36 38 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=4.45 $Y=1.555
+ $X2=4.655 $Y2=1.555
r141 33 34 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.62 $Y=2.89
+ $X2=3.62 $Y2=3.12
r142 31 32 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.045 $Y=2.06
+ $X2=2.045 $Y2=2.21
r143 27 30 733.255 $w=1.5e-07 $l=1.43e-06 $layer=POLY_cond $X=5.985 $Y=0.835
+ $X2=5.985 $Y2=2.265
r144 25 30 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.985 $Y=2.815
+ $X2=5.985 $Y2=2.265
r145 24 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.73 $Y=2.89
+ $X2=4.655 $Y2=2.89
r146 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.91 $Y=2.89
+ $X2=5.985 $Y2=2.815
r147 23 24 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=5.91 $Y=2.89
+ $X2=4.73 $Y2=2.89
r148 20 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.655 $Y=2.815
+ $X2=4.655 $Y2=2.89
r149 20 22 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.655 $Y=2.815
+ $X2=4.655 $Y2=2.265
r150 19 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.655 $Y=1.63
+ $X2=4.655 $Y2=1.555
r151 19 22 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.655 $Y=1.63
+ $X2=4.655 $Y2=2.265
r152 15 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.45 $Y=1.48
+ $X2=4.45 $Y2=1.555
r153 15 17 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=4.45 $Y=1.48
+ $X2=4.45 $Y2=0.625
r154 14 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.695 $Y=2.89
+ $X2=3.62 $Y2=2.89
r155 13 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.58 $Y=2.89
+ $X2=4.655 $Y2=2.89
r156 13 14 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=4.58 $Y=2.89
+ $X2=3.695 $Y2=2.89
r157 12 33 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.62 $Y=2.815
+ $X2=3.62 $Y2=2.89
r158 12 54 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.62 $Y=2.815
+ $X2=3.62 $Y2=2.125
r159 9 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.545 $Y=3.12
+ $X2=3.62 $Y2=3.12
r160 9 10 748.638 $w=1.5e-07 $l=1.46e-06 $layer=POLY_cond $X=3.545 $Y=3.12
+ $X2=2.085 $Y2=3.12
r161 7 31 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=2.08 $Y=0.895
+ $X2=2.08 $Y2=2.06
r162 4 32 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.01 $Y=2.495
+ $X2=2.01 $Y2=2.21
r163 2 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.01 $Y=3.045
+ $X2=2.085 $Y2=3.12
r164 2 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.01 $Y=3.045
+ $X2=2.01 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%A_1118_411# 1 2 9 12 14 18 20 25 27 31 33 34 35
+ 38
c77 38 0 3.79636e-21 $X=7.585 $Y=1.19
c78 27 0 2.36875e-19 $X=5.77 $Y=2.265
r79 34 39 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.585 $Y=1.355
+ $X2=7.585 $Y2=1.52
r80 34 38 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.585 $Y=1.355
+ $X2=7.585 $Y2=1.19
r81 33 36 5.26624 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=1.355
+ $X2=7.475 $Y2=1.52
r82 33 35 8.18509 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=1.355
+ $X2=7.475 $Y2=1.19
r83 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.575
+ $Y=1.355 $X2=7.575 $Y2=1.355
r84 27 29 5.12197 $w=2.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.74 $Y=2.265
+ $X2=5.74 $Y2=2.385
r85 25 36 26.833 $w=3.33e-07 $l=7.8e-07 $layer=LI1_cond $X=7.457 $Y=2.3
+ $X2=7.457 $Y2=1.52
r86 22 35 10.7828 $w=1.78e-07 $l=1.75e-07 $layer=LI1_cond $X=7.38 $Y=1.015
+ $X2=7.38 $Y2=1.19
r87 20 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.29 $Y=0.93
+ $X2=7.38 $Y2=1.015
r88 20 31 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.29 $Y=0.93 $X2=6.97
+ $Y2=0.93
r89 19 29 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.875 $Y=2.385
+ $X2=5.74 $Y2=2.385
r90 18 25 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=7.29 $Y=2.385
+ $X2=7.457 $Y2=2.3
r91 18 19 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=7.29 $Y=2.385
+ $X2=5.875 $Y2=2.385
r92 14 31 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=6.795 $Y=0.84
+ $X2=6.97 $Y2=0.84
r93 14 16 33.7501 $w=3.48e-07 $l=1.025e-06 $layer=LI1_cond $X=6.795 $Y=0.84
+ $X2=5.77 $Y2=0.84
r94 12 39 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=7.685 $Y=2.465
+ $X2=7.685 $Y2=1.52
r95 9 38 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=7.52 $Y=0.655
+ $X2=7.52 $Y2=1.19
r96 2 27 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=5.59
+ $Y=2.055 $X2=5.77 $Y2=2.265
r97 1 16 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.63
+ $Y=0.625 $X2=5.77 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%COUT 1 2 7 8 9 10 11 12 22 35
r16 32 35 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=0.23 $Y=1.96 $X2=0.23
+ $Y2=1.98
r17 12 40 20.0684 $w=2.88e-07 $l=5.05e-07 $layer=LI1_cond $X=0.23 $Y=2.405
+ $X2=0.23 $Y2=2.91
r18 11 32 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=0.23 $Y=1.955
+ $X2=0.23 $Y2=1.96
r19 11 43 5.56352 $w=2.88e-07 $l=1.4e-07 $layer=LI1_cond $X=0.23 $Y=1.955
+ $X2=0.23 $Y2=1.815
r20 11 12 14.5049 $w=2.88e-07 $l=3.65e-07 $layer=LI1_cond $X=0.23 $Y=2.04
+ $X2=0.23 $Y2=2.405
r21 11 35 2.38436 $w=2.88e-07 $l=6e-08 $layer=LI1_cond $X=0.23 $Y=2.04 $X2=0.23
+ $Y2=1.98
r22 10 43 6.1738 $w=2.78e-07 $l=1.5e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=1.815
r23 9 10 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r24 8 9 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r25 7 8 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.925
r26 7 22 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.42
r27 2 40 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.91
r28 2 35 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=1.98
r29 1 22 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%VPWR 1 2 3 4 5 18 22 26 29 32 35 36 38 42 43 44
+ 46 51 63 72 73 76 79 82
c103 38 0 1.12751e-19 $X=4.87 $Y=2.305
r104 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r105 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 73 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r108 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r109 70 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.45 $Y2=3.33
r110 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 69 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r113 66 69 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 65 68 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 63 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=3.33
+ $X2=7.45 $Y2=3.33
r117 63 68 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.285 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 59 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r121 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r122 56 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=2.735 $Y2=3.33
r123 56 58 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=3.6
+ $Y2=3.33
r124 55 80 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r125 55 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 52 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=2.735 $Y2=3.33
r130 51 54 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 49 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 46 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 46 48 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 44 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 44 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 42 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.845 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 42 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.845 $Y=3.33
+ $X2=4.94 $Y2=3.33
r139 41 65 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r140 41 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.94 $Y2=3.33
r141 38 40 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.87 $Y=2.305
+ $X2=4.87 $Y2=2.47
r142 35 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 35 36 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=4.002 $Y2=3.33
r144 34 61 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r145 34 36 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.12 $Y=3.33
+ $X2=4.002 $Y2=3.33
r146 30 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.45 $Y=3.245
+ $X2=7.45 $Y2=3.33
r147 30 32 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=7.45 $Y=3.245
+ $X2=7.45 $Y2=2.77
r148 29 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.94 $Y=3.245
+ $X2=4.94 $Y2=3.33
r149 29 40 45.2392 $w=1.88e-07 $l=7.75e-07 $layer=LI1_cond $X=4.94 $Y=3.245
+ $X2=4.94 $Y2=2.47
r150 24 36 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.002 $Y=3.245
+ $X2=4.002 $Y2=3.33
r151 24 26 48.0593 $w=2.33e-07 $l=9.8e-07 $layer=LI1_cond $X=4.002 $Y=3.245
+ $X2=4.002 $Y2=2.265
r152 20 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=3.245
+ $X2=2.735 $Y2=3.33
r153 20 22 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.735 $Y=3.245
+ $X2=2.735 $Y2=2.755
r154 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r155 16 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.765
r156 5 32 600 $w=1.7e-07 $l=9.04807e-07 $layer=licon1_PDIFF $count=1 $X=7.02
+ $Y=2.055 $X2=7.45 $Y2=2.77
r157 4 38 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=4.73
+ $Y=2.055 $X2=4.87 $Y2=2.305
r158 3 26 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=2.055 $X2=3.98 $Y2=2.265
r159 2 22 600 $w=1.7e-07 $l=5.69473e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=2.285 $X2=2.735 $Y2=2.755
r160 1 18 600 $w=1.7e-07 $l=1.00683e-06 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.72 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%A_417_457# 1 2 7 9
r24 9 12 4.03355 $w=2.98e-07 $l=1.05e-07 $layer=LI1_cond $X=2.24 $Y=2.385
+ $X2=2.24 $Y2=2.49
r25 8 9 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.39 $Y=2.385 $X2=2.24
+ $Y2=2.385
r26 7 17 4.97132 $w=2.53e-07 $l=1.1e-07 $layer=LI1_cond $X=3.207 $Y=2.385
+ $X2=3.207 $Y2=2.495
r27 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.08 $Y=2.385 $X2=2.39
+ $Y2=2.385
r28 2 17 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=2.285 $X2=3.245 $Y2=2.495
r29 1 12 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=2.285 $X2=2.225 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%A_854_411# 1 2 9 11 12 15
c29 15 0 1.78497e-19 $X=5.3 $Y=2.265
r30 13 15 11.5244 $w=2.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.32 $Y=2.035
+ $X2=5.32 $Y2=2.265
r31 11 13 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.205 $Y=1.95
+ $X2=5.32 $Y2=2.035
r32 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.205 $Y=1.95
+ $X2=4.535 $Y2=1.95
r33 7 12 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=4.412 $Y=2.035
+ $X2=4.535 $Y2=1.95
r34 7 9 10.8189 $w=2.43e-07 $l=2.3e-07 $layer=LI1_cond $X=4.412 $Y=2.035
+ $X2=4.412 $Y2=2.265
r35 2 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.16
+ $Y=2.055 $X2=5.3 $Y2=2.265
r36 1 9 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=2.055 $X2=4.44 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%SUM 1 2 7 9 15 16 17 22
r21 17 28 4.9369 $w=4.33e-07 $l=9.5e-08 $layer=LI1_cond $X=7.857 $Y=0.925
+ $X2=7.857 $Y2=1.02
r22 17 20 3.23214 $w=4.33e-07 $l=1.22e-07 $layer=LI1_cond $X=7.857 $Y=0.925
+ $X2=7.857 $Y2=0.803
r23 16 20 6.57025 $w=4.33e-07 $l=2.48e-07 $layer=LI1_cond $X=7.857 $Y=0.555
+ $X2=7.857 $Y2=0.803
r24 16 22 3.57655 $w=4.33e-07 $l=1.35e-07 $layer=LI1_cond $X=7.857 $Y=0.555
+ $X2=7.857 $Y2=0.42
r25 15 28 38.9869 $w=2.33e-07 $l=7.95e-07 $layer=LI1_cond $X=7.957 $Y=1.815
+ $X2=7.957 $Y2=1.02
r26 9 11 38.2776 $w=2.78e-07 $l=9.3e-07 $layer=LI1_cond $X=7.935 $Y=1.98
+ $X2=7.935 $Y2=2.91
r27 7 15 6.09362 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=7.935 $Y=1.955
+ $X2=7.935 $Y2=1.815
r28 7 9 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=7.935 $Y=1.955
+ $X2=7.935 $Y2=1.98
r29 2 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.835 $X2=7.9 $Y2=2.91
r30 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.835 $X2=7.9 $Y2=1.98
r31 1 22 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=7.595
+ $Y=0.235 $X2=7.755 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%VGND 1 2 3 4 5 18 24 28 30 34 38 40 41 43 44 45
+ 47 52 69 70 73 76 79
c96 34 0 9.76611e-20 $X=4.68 $Y=0.54
r97 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r98 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r99 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r100 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r101 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r102 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r103 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r104 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r105 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r106 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r107 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=0 $X2=4.68
+ $Y2=0
r108 61 63 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.845 $Y=0
+ $X2=5.04 $Y2=0
r109 60 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r110 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r111 57 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.725
+ $Y2=0
r112 57 59 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.6
+ $Y2=0
r113 56 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r114 56 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r115 55 73 13.2917 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=0.867
+ $Y2=0
r116 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.725
+ $Y2=0
r118 52 55 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=0 $X2=1.2
+ $Y2=0
r119 50 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r120 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r121 47 73 13.2917 $w=1.7e-07 $l=3.32e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.867 $Y2=0
r122 47 49 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r123 45 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r124 45 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r125 43 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=6.96
+ $Y2=0
r126 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=7.305
+ $Y2=0
r127 42 69 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=7.92
+ $Y2=0
r128 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=7.305
+ $Y2=0
r129 40 59 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.6
+ $Y2=0
r130 40 41 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.785
+ $Y2=0
r131 36 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0
r132 36 38 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0.55
r133 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.68 $Y=0.085
+ $X2=4.68 $Y2=0
r134 32 34 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=4.68 $Y=0.085
+ $X2=4.68 $Y2=0.54
r135 31 41 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.935 $Y=0 $X2=3.785
+ $Y2=0
r136 30 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.515 $Y=0 $X2=4.68
+ $Y2=0
r137 30 31 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.515 $Y=0
+ $X2=3.935 $Y2=0
r138 26 41 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0
r139 26 28 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0.63
r140 22 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0
r141 22 24 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0.895
r142 18 20 8.45349 $w=6.63e-07 $l=4.7e-07 $layer=LI1_cond $X=0.867 $Y=0.41
+ $X2=0.867 $Y2=0.88
r143 16 73 2.7522 $w=6.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.867 $Y=0.085
+ $X2=0.867 $Y2=0
r144 16 18 5.8455 $w=6.63e-07 $l=3.25e-07 $layer=LI1_cond $X=0.867 $Y=0.085
+ $X2=0.867 $Y2=0.41
r145 5 38 182 $w=1.7e-07 $l=3.20312e-07 $layer=licon1_NDIFF $count=1 $X=7.02
+ $Y=0.625 $X2=7.305 $Y2=0.55
r146 4 34 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.415 $X2=4.68 $Y2=0.54
r147 3 28 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=3.675
+ $Y=0.415 $X2=3.8 $Y2=0.63
r148 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.685 $X2=2.725 $Y2=0.895
r149 1 20 91 $w=1.7e-07 $l=8.26226e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.265 $X2=1.045 $Y2=0.88
r150 1 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.265 $X2=0.69 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%A_431_137# 1 2 9 11 12 15
c28 12 0 1.16441e-19 $X=2.39 $Y=1.27
r29 13 15 15.1913 $w=2.18e-07 $l=2.9e-07 $layer=LI1_cond $X=3.17 $Y=1.185
+ $X2=3.17 $Y2=0.895
r30 11 13 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.06 $Y=1.27
+ $X2=3.17 $Y2=1.185
r31 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.06 $Y=1.27
+ $X2=2.39 $Y2=1.27
r32 7 12 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=2.272 $Y=1.185
+ $X2=2.39 $Y2=1.27
r33 7 9 14.2216 $w=2.33e-07 $l=2.9e-07 $layer=LI1_cond $X=2.272 $Y=1.185
+ $X2=2.272 $Y2=0.895
r34 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.685 $X2=3.155 $Y2=0.895
r35 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.685 $X2=2.295 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__FA_1%A_818_83# 1 2 9 11 12 14
r24 14 16 8.97059 $w=4.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.255 $Y=0.55
+ $X2=5.255 $Y2=0.91
r25 11 16 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.015 $Y=0.91
+ $X2=5.255 $Y2=0.91
r26 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.015 $Y=0.91
+ $X2=4.345 $Y2=0.91
r27 7 12 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=4.225 $Y=0.825
+ $X2=4.345 $Y2=0.91
r28 7 9 9.3636 $w=2.38e-07 $l=1.95e-07 $layer=LI1_cond $X=4.225 $Y=0.825
+ $X2=4.225 $Y2=0.63
r29 2 14 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.97
+ $Y=0.415 $X2=5.11 $Y2=0.55
r30 1 9 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.415 $X2=4.23 $Y2=0.63
.ends

