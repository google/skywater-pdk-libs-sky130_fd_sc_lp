* File: sky130_fd_sc_lp__invlp_2.pex.spice
* Created: Fri Aug 28 10:39:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVLP_2%A 1 3 6 8 12 16 18 22 26 28 32 36 38 39 40
+ 41 48
c76 1 0 1.6164e-19 $X=0.505 $Y=1.225
r77 47 48 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=1.39
+ $X2=0.58 $Y2=1.39
r78 44 47 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.29 $Y=1.39
+ $X2=0.505 $Y2=1.39
r79 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.39 $X2=0.29 $Y2=1.39
r80 41 45 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.39
r81 34 40 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.865 $Y=1.405
+ $X2=1.83 $Y2=1.48
r82 34 36 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.865 $Y=1.405
+ $X2=1.865 $Y2=0.695
r83 30 40 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.795 $Y=1.555
+ $X2=1.83 $Y2=1.48
r84 30 32 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.795 $Y=1.555
+ $X2=1.795 $Y2=2.465
r85 29 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.44 $Y=1.48 $X2=1.365
+ $Y2=1.48
r86 28 40 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.72 $Y=1.48
+ $X2=1.83 $Y2=1.48
r87 28 29 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.72 $Y=1.48
+ $X2=1.44 $Y2=1.48
r88 24 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.365 $Y=1.555
+ $X2=1.365 $Y2=1.48
r89 24 26 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.365 $Y=1.555
+ $X2=1.365 $Y2=2.465
r90 20 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.365 $Y=1.405
+ $X2=1.365 $Y2=1.48
r91 20 22 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.365 $Y=1.405
+ $X2=1.365 $Y2=0.695
r92 19 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.01 $Y=1.48 $X2=0.935
+ $Y2=1.48
r93 18 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.48 $X2=1.365
+ $Y2=1.48
r94 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.29 $Y=1.48
+ $X2=1.01 $Y2=1.48
r95 14 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.935 $Y=1.555
+ $X2=0.935 $Y2=1.48
r96 14 16 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=0.935 $Y=1.555
+ $X2=0.935 $Y2=2.465
r97 10 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.935 $Y=1.405
+ $X2=0.935 $Y2=1.48
r98 10 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.935 $Y=1.405
+ $X2=0.935 $Y2=0.695
r99 8 38 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.86 $Y=1.48 $X2=0.935
+ $Y2=1.48
r100 8 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.86 $Y=1.48
+ $X2=0.58 $Y2=1.48
r101 4 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.555
+ $X2=0.505 $Y2=1.39
r102 4 6 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=0.505 $Y=1.555
+ $X2=0.505 $Y2=2.465
r103 1 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.225
+ $X2=0.505 $Y2=1.39
r104 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.505 $Y=1.225
+ $X2=0.505 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_2%VPWR 1 2 7 9 13 15 19 21 34
r33 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r39 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 22 30 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r41 22 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 21 33 4.65202 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.157 $Y2=3.33
r43 21 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 19 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 19 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 15 18 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=2.08 $Y=1.98
+ $X2=2.08 $Y2=2.95
r47 13 33 3.11416 $w=3.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.157 $Y2=3.33
r48 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.95
r49 9 12 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=0.29 $Y=1.98 $X2=0.29
+ $Y2=2.95
r50 7 30 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.227 $Y2=3.33
r51 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.95
r52 2 18 400 $w=1.7e-07 $l=1.21547e-06 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.835 $X2=2.08 $Y2=2.95
r53 2 15 400 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.835 $X2=2.08 $Y2=1.98
r54 1 12 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.29 $Y2=2.95
r55 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.29 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_2%A_116_367# 1 2 7 9 11 13 15
r27 13 20 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.905
+ $X2=1.62 $Y2=2.99
r28 13 15 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=1.62 $Y=2.905
+ $X2=1.62 $Y2=1.98
r29 12 18 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=2.99
+ $X2=0.72 $Y2=2.99
r30 11 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.495 $Y=2.99
+ $X2=1.62 $Y2=2.99
r31 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.495 $Y=2.99
+ $X2=0.805 $Y2=2.99
r32 7 18 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.905 $X2=0.72
+ $Y2=2.99
r33 7 9 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=0.72 $Y=2.905
+ $X2=0.72 $Y2=1.98
r34 2 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.835 $X2=1.58 $Y2=2.91
r35 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.835 $X2=1.58 $Y2=1.98
r36 1 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.91
r37 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_2%Y 1 2 7 8 9 10 11
r21 10 11 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.15 $Y=1.98
+ $X2=1.15 $Y2=2.405
r22 9 10 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.98
r23 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=1.295 $X2=1.15
+ $Y2=1.665
r24 7 8 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.15 $Y=0.865 $X2=1.15
+ $Y2=1.295
r25 2 10 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=1.98
r26 1 7 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.275 $X2=1.15 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_2%VGND 1 2 7 9 11 13 15 17 30
r28 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r29 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r30 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r31 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r33 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r34 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 18 26 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r36 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r37 17 29 3.96406 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.197
+ $Y2=0
r38 17 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=1.68
+ $Y2=0
r39 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r40 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r41 11 29 3.1791 $w=2.5e-07 $l=1.17346e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.197 $Y2=0
r42 11 13 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0.42
r43 7 26 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r44 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.29 $Y=0.085 $X2=0.29
+ $Y2=0.42
r45 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.94
+ $Y=0.275 $X2=2.08 $Y2=0.42
r46 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.275 $X2=0.29 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_2%A_116_55# 1 2 9 14 16
c25 14 0 1.6164e-19 $X=0.72 $Y=0.42
r26 10 14 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.34
+ $X2=0.72 $Y2=0.34
r27 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=0.34
+ $X2=1.65 $Y2=0.34
r28 9 10 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.485 $Y=0.34
+ $X2=0.805 $Y2=0.34
r29 2 16 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.44
+ $Y=0.275 $X2=1.65 $Y2=0.42
r30 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.275 $X2=0.72 $Y2=0.42
.ends

