# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o21ai_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o21ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.375000 0.455000 1.695000 ;
        RECT 0.125000 1.695000 2.355000 1.750000 ;
        RECT 0.125000 1.750000 1.415000 1.865000 ;
        RECT 1.245000 1.345000 2.355000 1.695000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.185000 1.025000 1.515000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.210000 3.265000 1.750000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.940800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 2.035000 2.735000 2.205000 ;
        RECT 1.000000 2.205000 1.300000 2.735000 ;
        RECT 1.595000 1.920000 2.735000 2.035000 ;
        RECT 2.500000 2.205000 2.735000 3.075000 ;
        RECT 2.525000 0.595000 2.735000 1.920000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.110000  0.255000 0.370000 0.845000 ;
      RECT 0.110000  0.845000 1.365000 1.005000 ;
      RECT 0.110000  1.005000 2.355000 1.015000 ;
      RECT 0.110000  2.035000 0.440000 3.245000 ;
      RECT 0.540000  0.085000 0.870000 0.675000 ;
      RECT 0.610000  2.035000 0.830000 2.905000 ;
      RECT 0.610000  2.905000 1.805000 3.075000 ;
      RECT 1.040000  0.255000 1.365000 0.845000 ;
      RECT 1.195000  1.015000 2.355000 1.175000 ;
      RECT 1.475000  2.375000 1.805000 2.905000 ;
      RECT 1.535000  0.085000 1.865000 0.825000 ;
      RECT 2.000000  2.375000 2.330000 3.245000 ;
      RECT 2.035000  0.255000 3.215000 0.425000 ;
      RECT 2.035000  0.425000 2.355000 1.005000 ;
      RECT 2.905000  0.425000 3.215000 1.040000 ;
      RECT 2.905000  1.920000 3.215000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__o21ai_2
