* NGSPICE file created from sky130_fd_sc_lp__a21boi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21boi_lp A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 Y a_298_318# a_29_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=5.65e+11p ps=5.13e+06u
M1001 a_298_318# B1_N VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=5.65e+11p ps=5.13e+06u
M1002 VPWR A2 a_29_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_172_47# A2 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.772e+11p ps=3e+06u
M1004 Y A1 a_172_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1005 a_29_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_298_318# a_336_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_513_47# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_298_318# B1_N a_513_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1009 a_336_47# a_298_318# Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

