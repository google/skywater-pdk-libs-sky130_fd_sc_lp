* File: sky130_fd_sc_lp__a22oi_2.pxi.spice
* Created: Wed Sep  2 09:23:11 2020
* 
x_PM_SKY130_FD_SC_LP__A22OI_2%A1 N_A1_M1004_g N_A1_M1002_g N_A1_M1003_g
+ N_A1_M1014_g A1 A1 A1 A1 N_A1_c_75_n N_A1_c_76_n N_A1_c_77_n N_A1_c_78_n
+ N_A1_c_87_p PM_SKY130_FD_SC_LP__A22OI_2%A1
x_PM_SKY130_FD_SC_LP__A22OI_2%A2 N_A2_M1001_g N_A2_M1007_g N_A2_c_162_n
+ N_A2_M1013_g N_A2_M1009_g N_A2_c_164_n A2 A2 N_A2_c_165_n N_A2_c_166_n
+ PM_SKY130_FD_SC_LP__A22OI_2%A2
x_PM_SKY130_FD_SC_LP__A22OI_2%B1 N_B1_M1008_g N_B1_M1000_g N_B1_M1011_g
+ N_B1_M1015_g N_B1_c_223_n N_B1_c_224_n N_B1_c_241_p N_B1_c_267_p N_B1_c_231_n
+ B1 N_B1_c_225_n N_B1_c_226_n PM_SKY130_FD_SC_LP__A22OI_2%B1
x_PM_SKY130_FD_SC_LP__A22OI_2%B2 N_B2_M1006_g N_B2_M1005_g N_B2_M1012_g
+ N_B2_M1010_g B2 N_B2_c_298_n N_B2_c_299_n PM_SKY130_FD_SC_LP__A22OI_2%B2
x_PM_SKY130_FD_SC_LP__A22OI_2%A_49_367# N_A_49_367#_M1004_d N_A_49_367#_M1001_d
+ N_A_49_367#_M1014_d N_A_49_367#_M1005_s N_A_49_367#_M1015_d
+ N_A_49_367#_c_346_n N_A_49_367#_c_351_n N_A_49_367#_c_355_n
+ N_A_49_367#_c_356_n N_A_49_367#_c_360_n N_A_49_367#_c_383_p
+ N_A_49_367#_c_376_n N_A_49_367#_c_361_n N_A_49_367#_c_373_n
+ N_A_49_367#_c_347_n N_A_49_367#_c_348_n N_A_49_367#_c_349_n
+ N_A_49_367#_c_363_n N_A_49_367#_c_364_n N_A_49_367#_c_378_n
+ PM_SKY130_FD_SC_LP__A22OI_2%A_49_367#
x_PM_SKY130_FD_SC_LP__A22OI_2%VPWR N_VPWR_M1004_s N_VPWR_M1013_s N_VPWR_c_420_n
+ N_VPWR_c_421_n N_VPWR_c_422_n VPWR N_VPWR_c_423_n N_VPWR_c_424_n
+ N_VPWR_c_419_n N_VPWR_c_426_n PM_SKY130_FD_SC_LP__A22OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A22OI_2%Y N_Y_M1002_d N_Y_M1003_d N_Y_M1011_s N_Y_M1000_s
+ N_Y_M1010_d N_Y_c_484_n N_Y_c_485_n N_Y_c_486_n N_Y_c_500_n N_Y_c_520_n
+ N_Y_c_501_n N_Y_c_487_n N_Y_c_488_n N_Y_c_489_n N_Y_c_531_n Y Y
+ PM_SKY130_FD_SC_LP__A22OI_2%Y
x_PM_SKY130_FD_SC_LP__A22OI_2%A_179_47# N_A_179_47#_M1002_s N_A_179_47#_M1009_s
+ N_A_179_47#_c_581_n N_A_179_47#_c_582_n N_A_179_47#_c_583_n
+ N_A_179_47#_c_584_n PM_SKY130_FD_SC_LP__A22OI_2%A_179_47#
x_PM_SKY130_FD_SC_LP__A22OI_2%VGND N_VGND_M1007_d N_VGND_M1006_s N_VGND_c_609_n
+ N_VGND_c_610_n VGND N_VGND_c_611_n N_VGND_c_612_n N_VGND_c_613_n
+ N_VGND_c_614_n N_VGND_c_615_n N_VGND_c_616_n PM_SKY130_FD_SC_LP__A22OI_2%VGND
x_PM_SKY130_FD_SC_LP__A22OI_2%A_595_47# N_A_595_47#_M1008_d N_A_595_47#_M1012_d
+ N_A_595_47#_c_682_n N_A_595_47#_c_673_n N_A_595_47#_c_678_n
+ N_A_595_47#_c_672_n PM_SKY130_FD_SC_LP__A22OI_2%A_595_47#
cc_1 VNB N_A1_M1002_g 0.033251f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=0.655
cc_2 VNB N_A1_M1003_g 0.0267623f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.655
cc_3 VNB N_A1_c_75_n 0.00113831f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_4 VNB N_A1_c_76_n 0.0409546f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.51
cc_5 VNB N_A1_c_77_n 0.0330809f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.51
cc_6 VNB N_A1_c_78_n 9.38405e-19 $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.51
cc_7 VNB N_A2_M1001_g 0.00663386f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_8 VNB N_A2_M1007_g 0.0262126f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=0.655
cc_9 VNB N_A2_c_162_n 0.0111061f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.345
cc_10 VNB N_A2_M1009_g 0.0261906f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_11 VNB N_A2_c_164_n 0.00508929f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.95
cc_12 VNB N_A2_c_165_n 0.0184927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_166_n 0.00490814f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.51
cc_14 VNB N_B1_M1008_g 0.0281749f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_15 VNB N_B1_M1011_g 0.0330085f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.655
cc_16 VNB N_B1_c_223_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.95
cc_17 VNB N_B1_c_224_n 0.0272338f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.95
cc_18 VNB N_B1_c_225_n 0.028158f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_19 VNB N_B1_c_226_n 0.0169326f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.51
cc_20 VNB N_B2_M1006_g 0.0251564f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_21 VNB N_B2_M1012_g 0.0236222f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.655
cc_22 VNB N_B2_c_298_n 9.30763e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B2_c_299_n 0.0332138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_419_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_25 VNB N_Y_c_484_n 0.0279698f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_26 VNB N_Y_c_485_n 0.0186198f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.95
cc_27 VNB N_Y_c_486_n 0.0120381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_487_n 0.0307623f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_29 VNB N_Y_c_488_n 0.0287221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_489_n 0.0025176f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.51
cc_31 VNB Y 0.00668307f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=2.035
cc_32 VNB N_VGND_c_609_n 0.00561774f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.345
cc_33 VNB N_VGND_c_610_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.675
cc_34 VNB N_VGND_c_611_n 0.0399215f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_35 VNB N_VGND_c_612_n 0.044744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_613_n 0.0275477f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_37 VNB N_VGND_c_614_n 0.263973f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.51
cc_38 VNB N_VGND_c_615_n 0.00631563f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.51
cc_39 VNB N_VGND_c_616_n 0.00436333f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.675
cc_40 VPB N_A1_M1004_g 0.0274649f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_41 VPB N_A1_M1014_g 0.0214139f $X=-0.19 $Y=1.655 $X2=2.54 $Y2=2.465
cc_42 VPB N_A1_c_75_n 0.00127391f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_43 VPB N_A1_c_76_n 0.00890466f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.51
cc_44 VPB N_A1_c_77_n 0.0131977f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.51
cc_45 VPB N_A1_c_78_n 0.00238448f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.51
cc_46 VPB N_A2_M1001_g 0.020899f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_47 VPB N_A2_M1013_g 0.0217587f $X=-0.19 $Y=1.655 $X2=2.54 $Y2=1.675
cc_48 VPB N_A2_c_165_n 0.00630671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A2_c_166_n 0.00704089f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.51
cc_50 VPB N_B1_M1000_g 0.0188459f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=0.655
cc_51 VPB N_B1_M1015_g 0.0246094f $X=-0.19 $Y=1.655 $X2=2.54 $Y2=2.465
cc_52 VPB N_B1_c_223_n 0.00137458f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.95
cc_53 VPB N_B1_c_224_n 0.00694395f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.95
cc_54 VPB N_B1_c_231_n 0.00205237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B1_c_225_n 0.00668482f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_56 VPB N_B1_c_226_n 0.00879023f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.51
cc_57 VPB N_B2_M1005_g 0.0191338f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=0.655
cc_58 VPB N_B2_M1010_g 0.0186863f $X=-0.19 $Y=1.655 $X2=2.54 $Y2=2.465
cc_59 VPB N_B2_c_298_n 0.00263177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_B2_c_299_n 0.00481853f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_49_367#_c_346_n 0.0178477f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_62 VPB N_A_49_367#_c_347_n 0.0133753f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.51
cc_63 VPB N_A_49_367#_c_348_n 0.03085f $X=-0.19 $Y=1.655 $X2=2.125 $Y2=2.035
cc_64 VPB N_A_49_367#_c_349_n 0.0312277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_420_n 0.0050648f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.345
cc_66 VPB N_VPWR_c_421_n 0.0227966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_422_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.54 $Y2=1.675
cc_68 VPB N_VPWR_c_423_n 0.0163769f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.95
cc_69 VPB N_VPWR_c_424_n 0.0570031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_419_n 0.0504668f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_71 VPB N_VPWR_c_426_n 0.0160737f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.51
cc_72 VPB Y 0.00107528f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=2.035
cc_73 N_A1_M1004_g N_A2_M1001_g 0.030678f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A1_c_75_n N_A2_M1001_g 0.00401714f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_75 N_A1_c_87_p N_A2_M1001_g 0.0114198f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_76 N_A1_M1002_g N_A2_M1007_g 0.0274722f $X=0.82 $Y=0.655 $X2=0 $Y2=0
cc_77 N_A1_c_87_p N_A2_c_162_n 3.78953e-19 $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_78 N_A1_c_78_n N_A2_M1013_g 0.00533335f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_79 N_A1_c_87_p N_A2_M1013_g 0.0124346f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_80 N_A1_M1003_g N_A2_M1009_g 0.0269021f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_81 N_A1_c_75_n N_A2_c_164_n 3.42925e-19 $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_82 N_A1_c_76_n N_A2_c_164_n 0.0158003f $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_83 N_A1_c_77_n N_A2_c_165_n 0.0211166f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_84 N_A1_c_78_n N_A2_c_165_n 4.15203e-19 $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_85 N_A1_c_87_p N_A2_c_165_n 8.55878e-19 $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_86 N_A1_M1004_g N_A2_c_166_n 2.86795e-19 $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A1_c_75_n N_A2_c_166_n 0.0363451f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_88 N_A1_c_76_n N_A2_c_166_n 0.00232531f $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_89 N_A1_c_77_n N_A2_c_166_n 0.00118738f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_90 N_A1_c_78_n N_A2_c_166_n 0.0294939f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_91 N_A1_c_87_p N_A2_c_166_n 0.0582765f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A1_M1003_g N_B1_M1008_g 0.021819f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_93 N_A1_M1014_g N_B1_M1000_g 0.0505067f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A1_c_77_n N_B1_c_223_n 3.87502e-19 $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_95 N_A1_c_77_n N_B1_c_224_n 0.0142437f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_96 N_A1_c_87_p N_A_49_367#_M1001_d 0.003401f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A1_M1004_g N_A_49_367#_c_351_n 0.0147814f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_98 A1 N_A_49_367#_c_351_n 0.0162474f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_99 N_A1_c_76_n N_A_49_367#_c_351_n 6.05981e-19 $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_100 N_A1_c_87_p N_A_49_367#_c_351_n 0.0238732f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A1_M1004_g N_A_49_367#_c_355_n 8.31902e-19 $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_102 N_A1_M1014_g N_A_49_367#_c_356_n 0.00434033f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_103 A1 N_A_49_367#_c_356_n 0.0213021f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A1_c_77_n N_A_49_367#_c_356_n 8.94051e-19 $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A1_c_87_p N_A_49_367#_c_356_n 0.0342837f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A1_M1014_g N_A_49_367#_c_360_n 0.0054073f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A1_M1014_g N_A_49_367#_c_361_n 0.00702088f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A1_M1004_g N_A_49_367#_c_349_n 0.0118932f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A1_c_87_p N_A_49_367#_c_363_n 0.0153678f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_110 N_A1_M1014_g N_A_49_367#_c_364_n 0.0120235f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_111 A1 N_VPWR_M1004_s 0.00227604f $X=0.635 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_112 N_A1_c_75_n N_VPWR_M1004_s 0.00173249f $X=0.72 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A1_c_87_p N_VPWR_M1004_s 0.00976304f $X=2.125 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_114 A1 N_VPWR_M1013_s 0.00652414f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_115 N_A1_c_78_n N_VPWR_M1013_s 0.00389571f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_116 N_A1_c_87_p N_VPWR_M1013_s 0.0145269f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_117 N_A1_M1004_g N_VPWR_c_420_n 0.00790185f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A1_M1004_g N_VPWR_c_421_n 0.0054895f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A1_M1014_g N_VPWR_c_424_n 0.00403671f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A1_M1004_g N_VPWR_c_419_n 0.0115101f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A1_M1014_g N_VPWR_c_419_n 0.00707251f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A1_M1014_g N_VPWR_c_426_n 0.0112705f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A1_M1002_g N_Y_c_485_n 0.0143432f $X=0.82 $Y=0.655 $X2=0 $Y2=0
cc_124 N_A1_M1003_g N_Y_c_485_n 0.0151801f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_125 N_A1_c_75_n N_Y_c_485_n 0.0142833f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_126 N_A1_c_76_n N_Y_c_485_n 3.8067e-19 $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_127 N_A1_c_77_n N_Y_c_485_n 0.00200301f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A1_c_78_n N_Y_c_485_n 0.0184099f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A1_c_75_n N_Y_c_486_n 0.00546322f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A1_c_76_n N_Y_c_486_n 0.0060521f $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A1_M1003_g N_Y_c_500_n 0.0108295f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_132 N_A1_M1014_g N_Y_c_501_n 0.00612136f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A1_M1003_g N_Y_c_489_n 2.82828e-19 $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_134 N_A1_c_77_n N_Y_c_489_n 0.00577876f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A1_M1003_g Y 0.00371854f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_136 N_A1_M1014_g Y 0.016252f $X=2.54 $Y=2.465 $X2=0 $Y2=0
cc_137 A1 Y 0.0131944f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_138 N_A1_c_77_n Y 0.00683396f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_139 N_A1_c_78_n Y 0.0430841f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_140 N_A1_M1002_g N_A_179_47#_c_581_n 0.00445191f $X=0.82 $Y=0.655 $X2=0 $Y2=0
cc_141 N_A1_M1003_g N_A_179_47#_c_582_n 0.00218559f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_142 N_A1_M1002_g N_A_179_47#_c_583_n 0.00219277f $X=0.82 $Y=0.655 $X2=0 $Y2=0
cc_143 N_A1_M1003_g N_A_179_47#_c_584_n 0.00443498f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_144 N_A1_M1002_g N_VGND_c_611_n 0.00549284f $X=0.82 $Y=0.655 $X2=0 $Y2=0
cc_145 N_A1_M1003_g N_VGND_c_612_n 0.00549284f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_146 N_A1_M1002_g N_VGND_c_614_n 0.0112381f $X=0.82 $Y=0.655 $X2=0 $Y2=0
cc_147 N_A1_M1003_g N_VGND_c_614_n 0.0105121f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_148 N_A2_M1001_g N_A_49_367#_c_351_n 0.0120783f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A2_M1001_g N_A_49_367#_c_355_n 0.0100464f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A2_M1013_g N_A_49_367#_c_356_n 0.0141754f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A2_M1013_g N_A_49_367#_c_360_n 0.00182811f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A2_M1001_g N_A_49_367#_c_349_n 8.35549e-19 $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A2_M1001_g N_A_49_367#_c_363_n 7.32094e-19 $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A2_M1001_g N_VPWR_c_420_n 0.006481f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A2_M1001_g N_VPWR_c_423_n 0.0054895f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A2_M1013_g N_VPWR_c_423_n 0.00486043f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A2_M1001_g N_VPWR_c_419_n 0.0104478f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A2_M1013_g N_VPWR_c_419_n 0.00819843f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A2_M1001_g N_VPWR_c_426_n 6.75001e-19 $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_M1013_g N_VPWR_c_426_n 0.0140822f $X=1.66 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A2_M1007_g N_Y_c_485_n 0.0113078f $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A2_c_162_n N_Y_c_485_n 0.00620606f $X=1.585 $Y=1.42 $X2=0 $Y2=0
cc_163 N_A2_M1009_g N_Y_c_485_n 0.0113078f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A2_c_164_n N_Y_c_485_n 5.23484e-19 $X=1.24 $Y=1.42 $X2=0 $Y2=0
cc_165 N_A2_c_166_n N_Y_c_485_n 0.0624688f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A2_M1007_g N_A_179_47#_c_581_n 0.0060262f $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_167 N_A2_M1009_g N_A_179_47#_c_581_n 8.09583e-19 $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A2_M1007_g N_A_179_47#_c_582_n 0.00937322f $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A2_M1009_g N_A_179_47#_c_582_n 0.010088f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A2_M1007_g N_A_179_47#_c_583_n 7.14816e-19 $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_171 N_A2_M1007_g N_A_179_47#_c_584_n 8.09583e-19 $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_172 N_A2_M1009_g N_A_179_47#_c_584_n 0.0060262f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_173 N_A2_M1007_g N_VGND_c_609_n 0.00466906f $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A2_M1009_g N_VGND_c_609_n 0.00466906f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_175 N_A2_M1007_g N_VGND_c_611_n 0.00418148f $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_176 N_A2_M1009_g N_VGND_c_612_n 0.00418148f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A2_M1007_g N_VGND_c_614_n 0.00617763f $X=1.25 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A2_M1009_g N_VGND_c_614_n 0.00617763f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_179 N_B1_M1008_g N_B2_M1006_g 0.0265294f $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_180 N_B1_M1000_g N_B2_M1005_g 0.0444632f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B1_c_223_n N_B2_M1005_g 0.00422708f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_182 N_B1_c_241_p N_B2_M1005_g 0.0106216f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_183 N_B1_M1011_g N_B2_M1012_g 0.0344971f $X=4.3 $Y=0.655 $X2=0 $Y2=0
cc_184 N_B1_M1015_g N_B2_M1010_g 0.0344971f $X=4.3 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B1_c_241_p N_B2_M1010_g 0.0139831f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_186 N_B1_c_231_n N_B2_M1010_g 0.00246081f $X=4.075 $Y=1.925 $X2=0 $Y2=0
cc_187 N_B1_c_223_n N_B2_c_298_n 0.0260251f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_188 N_B1_c_224_n N_B2_c_298_n 0.00114773f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_189 N_B1_c_241_p N_B2_c_298_n 0.0297397f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_190 N_B1_c_225_n N_B2_c_298_n 2.87961e-19 $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_191 N_B1_c_226_n N_B2_c_298_n 0.0341877f $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_192 N_B1_c_223_n N_B2_c_299_n 0.00127982f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_193 N_B1_c_224_n N_B2_c_299_n 0.0210055f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_194 N_B1_c_241_p N_B2_c_299_n 5.75497e-19 $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_195 N_B1_c_225_n N_B2_c_299_n 0.0344971f $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_196 N_B1_c_226_n N_B2_c_299_n 0.00378915f $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_197 N_B1_c_241_p N_A_49_367#_M1005_s 0.0033488f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_198 N_B1_M1000_g N_A_49_367#_c_361_n 0.0173446f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_199 N_B1_M1015_g N_A_49_367#_c_373_n 0.0157945f $X=4.3 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B1_c_225_n N_A_49_367#_c_348_n 8.63371e-19 $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_201 N_B1_c_226_n N_A_49_367#_c_348_n 0.00915064f $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_202 N_B1_M1000_g N_VPWR_c_424_n 0.00357877f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B1_M1015_g N_VPWR_c_424_n 0.00357877f $X=4.3 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B1_M1000_g N_VPWR_c_419_n 0.00557742f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B1_M1015_g N_VPWR_c_419_n 0.00633391f $X=4.3 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B1_c_223_n N_Y_M1000_s 0.00111282f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_207 N_B1_c_241_p N_Y_M1000_s 0.00741937f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_208 N_B1_c_267_p N_Y_M1000_s 5.76861e-19 $X=3.155 $Y=2.01 $X2=0 $Y2=0
cc_209 N_B1_c_241_p N_Y_M1010_d 0.00397593f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_210 N_B1_c_231_n N_Y_M1010_d 9.85787e-19 $X=4.075 $Y=1.925 $X2=0 $Y2=0
cc_211 N_B1_M1008_g N_Y_c_500_n 0.0105576f $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_212 N_B1_M1000_g N_Y_c_520_n 0.00868225f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B1_c_224_n N_Y_c_520_n 0.00150565f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_214 N_B1_c_241_p N_Y_c_520_n 0.0417055f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_215 N_B1_c_267_p N_Y_c_520_n 0.0148555f $X=3.155 $Y=2.01 $X2=0 $Y2=0
cc_216 N_B1_M1008_g N_Y_c_487_n 0.0187393f $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_217 N_B1_M1011_g N_Y_c_487_n 0.0147729f $X=4.3 $Y=0.655 $X2=0 $Y2=0
cc_218 N_B1_c_223_n N_Y_c_487_n 0.019561f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_219 N_B1_c_224_n N_Y_c_487_n 0.00125527f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_220 N_B1_c_225_n N_Y_c_487_n 0.00416915f $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_221 N_B1_c_226_n N_Y_c_487_n 0.0453626f $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_222 N_B1_M1008_g N_Y_c_489_n 3.28046e-19 $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_223 N_B1_M1015_g N_Y_c_531_n 0.00380644f $X=4.3 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B1_c_241_p N_Y_c_531_n 0.01489f $X=3.985 $Y=2.01 $X2=0 $Y2=0
cc_225 N_B1_c_226_n N_Y_c_531_n 0.00170819f $X=4.39 $Y=1.51 $X2=0 $Y2=0
cc_226 N_B1_M1008_g Y 0.00676863f $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_227 N_B1_M1000_g Y 0.00598307f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_228 N_B1_c_223_n Y 0.0427713f $X=2.99 $Y=1.51 $X2=0 $Y2=0
cc_229 N_B1_c_267_p Y 0.013441f $X=3.155 $Y=2.01 $X2=0 $Y2=0
cc_230 N_B1_M1008_g N_VGND_c_610_n 9.88819e-19 $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_231 N_B1_M1011_g N_VGND_c_610_n 0.00180633f $X=4.3 $Y=0.655 $X2=0 $Y2=0
cc_232 N_B1_M1008_g N_VGND_c_612_n 0.00585385f $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_233 N_B1_M1011_g N_VGND_c_613_n 0.00580562f $X=4.3 $Y=0.655 $X2=0 $Y2=0
cc_234 N_B1_M1008_g N_VGND_c_614_n 0.0116064f $X=2.9 $Y=0.655 $X2=0 $Y2=0
cc_235 N_B1_M1011_g N_VGND_c_614_n 0.0116712f $X=4.3 $Y=0.655 $X2=0 $Y2=0
cc_236 N_B1_M1011_g N_A_595_47#_c_672_n 0.00305845f $X=4.3 $Y=0.655 $X2=0 $Y2=0
cc_237 N_B2_M1005_g N_A_49_367#_c_376_n 0.0143707f $X=3.44 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B2_M1010_g N_A_49_367#_c_373_n 0.012036f $X=3.87 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B2_M1005_g N_A_49_367#_c_378_n 0.00245543f $X=3.44 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B2_M1010_g N_A_49_367#_c_378_n 0.00467378f $X=3.87 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B2_M1005_g N_VPWR_c_424_n 0.00357877f $X=3.44 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B2_M1010_g N_VPWR_c_424_n 0.00357877f $X=3.87 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B2_M1005_g N_VPWR_c_419_n 0.00551022f $X=3.44 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B2_M1010_g N_VPWR_c_419_n 0.00540931f $X=3.87 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B2_M1005_g N_Y_c_520_n 0.00844278f $X=3.44 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B2_M1010_g N_Y_c_520_n 0.00864832f $X=3.87 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B2_M1006_g N_Y_c_487_n 0.0109928f $X=3.44 $Y=0.655 $X2=0 $Y2=0
cc_248 N_B2_M1012_g N_Y_c_487_n 0.0144461f $X=3.87 $Y=0.655 $X2=0 $Y2=0
cc_249 N_B2_c_298_n N_Y_c_487_n 0.0337458f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_250 N_B2_c_299_n N_Y_c_487_n 7.04948e-19 $X=3.87 $Y=1.51 $X2=0 $Y2=0
cc_251 N_B2_M1005_g N_Y_c_531_n 8.61997e-19 $X=3.44 $Y=2.465 $X2=0 $Y2=0
cc_252 N_B2_M1010_g N_Y_c_531_n 0.00444958f $X=3.87 $Y=2.465 $X2=0 $Y2=0
cc_253 N_B2_M1006_g N_VGND_c_610_n 0.00798892f $X=3.44 $Y=0.655 $X2=0 $Y2=0
cc_254 N_B2_M1012_g N_VGND_c_610_n 0.00988541f $X=3.87 $Y=0.655 $X2=0 $Y2=0
cc_255 N_B2_M1006_g N_VGND_c_612_n 0.0035715f $X=3.44 $Y=0.655 $X2=0 $Y2=0
cc_256 N_B2_M1012_g N_VGND_c_613_n 0.0035715f $X=3.87 $Y=0.655 $X2=0 $Y2=0
cc_257 N_B2_M1006_g N_VGND_c_614_n 0.00454122f $X=3.44 $Y=0.655 $X2=0 $Y2=0
cc_258 N_B2_M1012_g N_VGND_c_614_n 0.00428043f $X=3.87 $Y=0.655 $X2=0 $Y2=0
cc_259 N_B2_M1006_g N_A_595_47#_c_673_n 0.0120015f $X=3.44 $Y=0.655 $X2=0 $Y2=0
cc_260 N_B2_M1012_g N_A_595_47#_c_673_n 0.00966879f $X=3.87 $Y=0.655 $X2=0 $Y2=0
cc_261 N_A_49_367#_c_351_n N_VPWR_M1004_s 0.0106548f $X=1.28 $Y=2.375 $X2=-0.19
+ $Y2=1.655
cc_262 N_A_49_367#_c_356_n N_VPWR_M1013_s 0.017262f $X=2.21 $Y=2.375 $X2=0 $Y2=0
cc_263 N_A_49_367#_c_360_n N_VPWR_M1013_s 0.00449677f $X=2.295 $Y=2.605 $X2=0
+ $Y2=0
cc_264 N_A_49_367#_c_383_p N_VPWR_M1013_s 0.00428442f $X=2.38 $Y=2.69 $X2=0
+ $Y2=0
cc_265 N_A_49_367#_c_364_n N_VPWR_M1013_s 0.00130124f $X=2.59 $Y=2.84 $X2=0
+ $Y2=0
cc_266 N_A_49_367#_c_351_n N_VPWR_c_420_n 0.0266856f $X=1.28 $Y=2.375 $X2=0
+ $Y2=0
cc_267 N_A_49_367#_c_355_n N_VPWR_c_420_n 0.0299545f $X=1.445 $Y=2.91 $X2=0
+ $Y2=0
cc_268 N_A_49_367#_c_349_n N_VPWR_c_420_n 0.0288374f $X=0.37 $Y=2.455 $X2=0
+ $Y2=0
cc_269 N_A_49_367#_c_349_n N_VPWR_c_421_n 0.0210467f $X=0.37 $Y=2.455 $X2=0
+ $Y2=0
cc_270 N_A_49_367#_c_355_n N_VPWR_c_423_n 0.015688f $X=1.445 $Y=2.91 $X2=0 $Y2=0
cc_271 N_A_49_367#_c_361_n N_VPWR_c_424_n 0.105298f $X=3.06 $Y=2.84 $X2=0 $Y2=0
cc_272 N_A_49_367#_c_347_n N_VPWR_c_424_n 0.0182731f $X=4.545 $Y=2.765 $X2=0
+ $Y2=0
cc_273 N_A_49_367#_c_364_n N_VPWR_c_424_n 0.00312738f $X=2.59 $Y=2.84 $X2=0
+ $Y2=0
cc_274 N_A_49_367#_M1004_d N_VPWR_c_419_n 0.00215158f $X=0.245 $Y=1.835 $X2=0
+ $Y2=0
cc_275 N_A_49_367#_M1001_d N_VPWR_c_419_n 0.00380103f $X=1.305 $Y=1.835 $X2=0
+ $Y2=0
cc_276 N_A_49_367#_M1014_d N_VPWR_c_419_n 0.00225186f $X=2.615 $Y=1.835 $X2=0
+ $Y2=0
cc_277 N_A_49_367#_M1005_s N_VPWR_c_419_n 0.00223577f $X=3.515 $Y=1.835 $X2=0
+ $Y2=0
cc_278 N_A_49_367#_M1015_d N_VPWR_c_419_n 0.0021516f $X=4.375 $Y=1.835 $X2=0
+ $Y2=0
cc_279 N_A_49_367#_c_355_n N_VPWR_c_419_n 0.00984745f $X=1.445 $Y=2.91 $X2=0
+ $Y2=0
cc_280 N_A_49_367#_c_383_p N_VPWR_c_419_n 9.76525e-19 $X=2.38 $Y=2.69 $X2=0
+ $Y2=0
cc_281 N_A_49_367#_c_361_n N_VPWR_c_419_n 0.0666895f $X=3.06 $Y=2.84 $X2=0 $Y2=0
cc_282 N_A_49_367#_c_347_n N_VPWR_c_419_n 0.010497f $X=4.545 $Y=2.765 $X2=0
+ $Y2=0
cc_283 N_A_49_367#_c_349_n N_VPWR_c_419_n 0.0125689f $X=0.37 $Y=2.455 $X2=0
+ $Y2=0
cc_284 N_A_49_367#_c_364_n N_VPWR_c_419_n 0.00497333f $X=2.59 $Y=2.84 $X2=0
+ $Y2=0
cc_285 N_A_49_367#_c_356_n N_VPWR_c_426_n 0.0281865f $X=2.21 $Y=2.375 $X2=0
+ $Y2=0
cc_286 N_A_49_367#_c_383_p N_VPWR_c_426_n 0.0260015f $X=2.38 $Y=2.69 $X2=0 $Y2=0
cc_287 N_A_49_367#_c_361_n N_VPWR_c_426_n 0.00558206f $X=3.06 $Y=2.84 $X2=0
+ $Y2=0
cc_288 N_A_49_367#_c_364_n N_VPWR_c_426_n 0.00204485f $X=2.59 $Y=2.84 $X2=0
+ $Y2=0
cc_289 N_A_49_367#_c_376_n N_Y_M1000_s 0.00424978f $X=3.49 $Y=2.84 $X2=0 $Y2=0
cc_290 N_A_49_367#_c_373_n N_Y_M1010_d 0.00330391f $X=4.41 $Y=2.92 $X2=0 $Y2=0
cc_291 N_A_49_367#_M1014_d N_Y_c_520_n 0.00469895f $X=2.615 $Y=1.835 $X2=0 $Y2=0
cc_292 N_A_49_367#_M1005_s N_Y_c_520_n 0.00349431f $X=3.515 $Y=1.835 $X2=0 $Y2=0
cc_293 N_A_49_367#_c_361_n N_Y_c_520_n 0.0581364f $X=3.06 $Y=2.84 $X2=0 $Y2=0
cc_294 N_A_49_367#_c_373_n N_Y_c_520_n 0.00578221f $X=4.41 $Y=2.92 $X2=0 $Y2=0
cc_295 N_A_49_367#_M1014_d N_Y_c_501_n 6.87795e-19 $X=2.615 $Y=1.835 $X2=0 $Y2=0
cc_296 N_A_49_367#_c_356_n N_Y_c_501_n 0.0126735f $X=2.21 $Y=2.375 $X2=0 $Y2=0
cc_297 N_A_49_367#_c_364_n N_Y_c_501_n 0.0104369f $X=2.59 $Y=2.84 $X2=0 $Y2=0
cc_298 N_A_49_367#_c_373_n N_Y_c_531_n 0.015511f $X=4.41 $Y=2.92 $X2=0 $Y2=0
cc_299 N_A_49_367#_M1014_d Y 0.00412215f $X=2.615 $Y=1.835 $X2=0 $Y2=0
cc_300 N_VPWR_c_419_n N_Y_M1000_s 0.00257355f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_301 N_VPWR_c_419_n N_Y_M1010_d 0.00225186f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_302 N_Y_c_485_n N_A_179_47#_M1002_s 0.00176461f $X=2.41 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_303 N_Y_c_485_n N_A_179_47#_M1009_s 0.00176461f $X=2.41 $Y=1.08 $X2=0 $Y2=0
cc_304 N_Y_c_485_n N_A_179_47#_c_582_n 0.0575179f $X=2.41 $Y=1.08 $X2=0 $Y2=0
cc_305 N_Y_c_500_n N_A_179_47#_c_582_n 0.0128488f $X=2.575 $Y=0.41 $X2=0 $Y2=0
cc_306 N_Y_c_485_n N_A_179_47#_c_583_n 0.0169621f $X=2.41 $Y=1.08 $X2=0 $Y2=0
cc_307 N_Y_c_500_n N_A_179_47#_c_584_n 0.027752f $X=2.575 $Y=0.41 $X2=0 $Y2=0
cc_308 N_Y_c_485_n N_VGND_M1007_d 0.0038237f $X=2.41 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_309 N_Y_c_487_n N_VGND_M1006_s 0.00176891f $X=4.4 $Y=1.09 $X2=0 $Y2=0
cc_310 N_Y_c_484_n N_VGND_c_611_n 0.0174563f $X=0.605 $Y=0.42 $X2=0 $Y2=0
cc_311 N_Y_c_500_n N_VGND_c_612_n 0.0230625f $X=2.575 $Y=0.41 $X2=0 $Y2=0
cc_312 N_Y_c_488_n N_VGND_c_613_n 0.0185207f $X=4.515 $Y=0.42 $X2=0 $Y2=0
cc_313 N_Y_M1002_d N_VGND_c_614_n 0.0040649f $X=0.48 $Y=0.235 $X2=0 $Y2=0
cc_314 N_Y_M1003_d N_VGND_c_614_n 0.00918806f $X=2.345 $Y=0.235 $X2=0 $Y2=0
cc_315 N_Y_M1011_s N_VGND_c_614_n 0.00302127f $X=4.375 $Y=0.235 $X2=0 $Y2=0
cc_316 N_Y_c_484_n N_VGND_c_614_n 0.00963639f $X=0.605 $Y=0.42 $X2=0 $Y2=0
cc_317 N_Y_c_500_n N_VGND_c_614_n 0.0127519f $X=2.575 $Y=0.41 $X2=0 $Y2=0
cc_318 N_Y_c_488_n N_VGND_c_614_n 0.010808f $X=4.515 $Y=0.42 $X2=0 $Y2=0
cc_319 N_Y_c_487_n N_A_595_47#_M1008_d 0.00304851f $X=4.4 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_320 N_Y_c_487_n N_A_595_47#_M1012_d 0.00176461f $X=4.4 $Y=1.09 $X2=0 $Y2=0
cc_321 N_Y_c_487_n N_A_595_47#_c_673_n 0.0323573f $X=4.4 $Y=1.09 $X2=0 $Y2=0
cc_322 N_Y_c_487_n N_A_595_47#_c_678_n 0.0221661f $X=4.4 $Y=1.09 $X2=0 $Y2=0
cc_323 N_Y_c_487_n N_A_595_47#_c_672_n 0.0129974f $X=4.4 $Y=1.09 $X2=0 $Y2=0
cc_324 N_A_179_47#_c_582_n N_VGND_M1007_d 0.0072679f $X=1.89 $Y=0.74 $X2=0.585
+ $Y2=1.675
cc_325 N_A_179_47#_c_582_n N_VGND_c_609_n 0.025007f $X=1.89 $Y=0.74 $X2=2.27
+ $Y2=1.345
cc_326 N_A_179_47#_c_581_n N_VGND_c_611_n 0.0176009f $X=1.035 $Y=0.37 $X2=0.635
+ $Y2=1.95
cc_327 N_A_179_47#_c_582_n N_VGND_c_611_n 0.00244463f $X=1.89 $Y=0.74 $X2=0.635
+ $Y2=1.95
cc_328 N_A_179_47#_c_582_n N_VGND_c_612_n 0.00244463f $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_329 N_A_179_47#_c_584_n N_VGND_c_612_n 0.0176009f $X=2.055 $Y=0.37 $X2=0
+ $Y2=0
cc_330 N_A_179_47#_M1002_s N_VGND_c_614_n 0.00223819f $X=0.895 $Y=0.235 $X2=0.82
+ $Y2=1.51
cc_331 N_A_179_47#_M1009_s N_VGND_c_614_n 0.00223819f $X=1.915 $Y=0.235 $X2=0.82
+ $Y2=1.51
cc_332 N_A_179_47#_c_581_n N_VGND_c_614_n 0.0122594f $X=1.035 $Y=0.37 $X2=0.82
+ $Y2=1.51
cc_333 N_A_179_47#_c_582_n N_VGND_c_614_n 0.0102757f $X=1.89 $Y=0.74 $X2=0.82
+ $Y2=1.51
cc_334 N_A_179_47#_c_584_n N_VGND_c_614_n 0.0122594f $X=2.055 $Y=0.37 $X2=0.82
+ $Y2=1.51
cc_335 N_VGND_c_614_n N_A_595_47#_M1008_d 0.00348522f $X=4.56 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_336 N_VGND_c_614_n N_A_595_47#_M1012_d 0.00285044f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_337 N_VGND_c_612_n N_A_595_47#_c_682_n 0.021382f $X=3.49 $Y=0 $X2=0 $Y2=0
cc_338 N_VGND_c_614_n N_A_595_47#_c_682_n 0.0130863f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_M1006_s N_A_595_47#_c_673_n 0.00335857f $X=3.515 $Y=0.235 $X2=0
+ $Y2=0
cc_340 N_VGND_c_610_n N_A_595_47#_c_673_n 0.0161464f $X=3.655 $Y=0.395 $X2=0
+ $Y2=0
cc_341 N_VGND_c_612_n N_A_595_47#_c_673_n 0.00230386f $X=3.49 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_c_613_n N_A_595_47#_c_673_n 0.00229766f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_614_n N_A_595_47#_c_673_n 0.00965909f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_344 N_VGND_c_613_n N_A_595_47#_c_672_n 0.00518942f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_345 N_VGND_c_614_n N_A_595_47#_c_672_n 0.00767521f $X=4.56 $Y=0 $X2=0 $Y2=0
