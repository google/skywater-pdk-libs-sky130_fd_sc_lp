* File: sky130_fd_sc_lp__o2111a_2.pxi.spice
* Created: Fri Aug 28 11:00:03 2020
* 
x_PM_SKY130_FD_SC_LP__O2111A_2%A_80_21# N_A_80_21#_M1001_s N_A_80_21#_M1003_d
+ N_A_80_21#_M1004_d N_A_80_21#_c_70_n N_A_80_21#_M1005_g N_A_80_21#_c_76_n
+ N_A_80_21#_M1007_g N_A_80_21#_c_71_n N_A_80_21#_M1008_g N_A_80_21#_c_77_n
+ N_A_80_21#_M1012_g N_A_80_21#_c_72_n N_A_80_21#_c_81_p N_A_80_21#_c_111_p
+ N_A_80_21#_c_73_n N_A_80_21#_c_95_p N_A_80_21#_c_96_p N_A_80_21#_c_107_p
+ N_A_80_21#_c_123_p N_A_80_21#_c_74_n N_A_80_21#_c_75_n N_A_80_21#_c_94_p
+ PM_SKY130_FD_SC_LP__O2111A_2%A_80_21#
x_PM_SKY130_FD_SC_LP__O2111A_2%D1 N_D1_M1003_g N_D1_M1001_g D1 N_D1_c_153_n
+ N_D1_c_151_n PM_SKY130_FD_SC_LP__O2111A_2%D1
x_PM_SKY130_FD_SC_LP__O2111A_2%C1 N_C1_M1002_g N_C1_M1013_g C1 C1 C1 C1
+ N_C1_c_187_n N_C1_c_188_n C1 PM_SKY130_FD_SC_LP__O2111A_2%C1
x_PM_SKY130_FD_SC_LP__O2111A_2%B1 N_B1_M1006_g N_B1_M1004_g B1 N_B1_c_229_n
+ PM_SKY130_FD_SC_LP__O2111A_2%B1
x_PM_SKY130_FD_SC_LP__O2111A_2%A2 N_A2_M1009_g N_A2_M1010_g A2 A2 A2 A2
+ N_A2_c_263_n PM_SKY130_FD_SC_LP__O2111A_2%A2
x_PM_SKY130_FD_SC_LP__O2111A_2%A1 N_A1_M1011_g N_A1_M1000_g A1 N_A1_c_296_n
+ N_A1_c_297_n PM_SKY130_FD_SC_LP__O2111A_2%A1
x_PM_SKY130_FD_SC_LP__O2111A_2%VPWR N_VPWR_M1007_d N_VPWR_M1012_d N_VPWR_M1013_d
+ N_VPWR_M1000_d N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n
+ N_VPWR_c_324_n N_VPWR_c_325_n VPWR N_VPWR_c_326_n N_VPWR_c_327_n
+ N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_319_n VPWR
+ PM_SKY130_FD_SC_LP__O2111A_2%VPWR
x_PM_SKY130_FD_SC_LP__O2111A_2%X N_X_M1005_d N_X_M1007_s X X X X X X X
+ N_X_c_378_n PM_SKY130_FD_SC_LP__O2111A_2%X
x_PM_SKY130_FD_SC_LP__O2111A_2%VGND N_VGND_M1005_s N_VGND_M1008_s N_VGND_M1009_d
+ N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n VGND
+ N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n
+ N_VGND_c_406_n VGND PM_SKY130_FD_SC_LP__O2111A_2%VGND
x_PM_SKY130_FD_SC_LP__O2111A_2%A_566_51# N_A_566_51#_M1006_d N_A_566_51#_M1011_d
+ N_A_566_51#_c_447_n N_A_566_51#_c_448_n N_A_566_51#_c_449_n
+ N_A_566_51#_c_450_n PM_SKY130_FD_SC_LP__O2111A_2%A_566_51#
cc_1 VNB N_A_80_21#_c_70_n 0.0215271f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A_80_21#_c_71_n 0.0191373f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_3 VNB N_A_80_21#_c_72_n 8.41245e-19 $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.955
cc_4 VNB N_A_80_21#_c_73_n 0.0097287f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=0.42
cc_5 VNB N_A_80_21#_c_74_n 0.0841095f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.35
cc_6 VNB N_A_80_21#_c_75_n 0.0196761f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.225
cc_7 VNB N_D1_M1001_g 0.0276752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D1_c_151_n 0.0333387f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_9 VNB N_C1_M1013_g 0.00516517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB C1 0.00318808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB C1 0.00406953f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_12 VNB N_C1_c_187_n 0.0325457f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_13 VNB N_C1_c_188_n 0.0156887f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_14 VNB N_B1_M1006_g 0.0263054f $X=-0.19 $Y=-0.245 $X2=2.83 $Y2=1.835
cc_15 VNB B1 0.00765812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_229_n 0.0242799f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_17 VNB N_A2_M1009_g 0.0260416f $X=-0.19 $Y=-0.245 $X2=2.83 $Y2=1.835
cc_18 VNB A2 0.00452943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_263_n 0.0225053f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.725
cc_20 VNB N_A1_M1011_g 0.0284153f $X=-0.19 $Y=-0.245 $X2=2.83 $Y2=1.835
cc_21 VNB N_A1_M1000_g 0.00176079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_296_n 0.0489658f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_23 VNB N_A1_c_297_n 0.0112304f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_24 VNB N_VPWR_c_319_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_378_n 0.00159056f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.515
cc_26 VNB N_VGND_c_397_n 0.0109056f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_27 VNB N_VGND_c_398_n 0.0496459f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_28 VNB N_VGND_c_399_n 0.00888396f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_29 VNB N_VGND_c_400_n 0.00626856f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_30 VNB N_VGND_c_401_n 0.0152194f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.04
cc_31 VNB N_VGND_c_402_n 0.0573799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_403_n 0.0181857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_404_n 0.263506f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.225
cc_34 VNB N_VGND_c_405_n 0.00486797f $X=-0.19 $Y=-0.245 $X2=2 $Y2=2.04
cc_35 VNB N_VGND_c_406_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.455
cc_36 VNB N_A_566_51#_c_447_n 0.00200919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_566_51#_c_448_n 0.0145907f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_38 VNB N_A_566_51#_c_449_n 0.0101299f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_39 VNB N_A_566_51#_c_450_n 0.031954f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_40 VPB N_A_80_21#_c_76_n 0.0216568f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.725
cc_41 VPB N_A_80_21#_c_77_n 0.0183692f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.725
cc_42 VPB N_A_80_21#_c_72_n 0.00221342f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=1.955
cc_43 VPB N_A_80_21#_c_74_n 0.021422f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.35
cc_44 VPB N_D1_M1003_g 0.022054f $X=-0.19 $Y=1.655 $X2=2.83 $Y2=1.835
cc_45 VPB N_D1_c_153_n 0.00292505f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.725
cc_46 VPB N_D1_c_151_n 0.0103268f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.185
cc_47 VPB N_C1_M1013_g 0.020181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB C1 0.00324567f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_49 VPB N_B1_M1004_g 0.0204014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB B1 0.00481711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B1_c_229_n 0.00638481f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_52 VPB N_A2_M1010_g 0.0215137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB A2 0.00379237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A2_c_263_n 0.00771465f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.725
cc_55 VPB N_A1_M1000_g 0.0264921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A1_c_297_n 0.00714397f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_57 VPB N_VPWR_c_320_n 0.0108797f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.725
cc_58 VPB N_VPWR_c_321_n 0.0654254f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_59 VPB N_VPWR_c_322_n 0.00236779f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_60 VPB N_VPWR_c_323_n 0.00495041f $X=-0.19 $Y=1.655 $X2=1.305 $Y2=2.04
cc_61 VPB N_VPWR_c_324_n 0.0106587f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=0.42
cc_62 VPB N_VPWR_c_325_n 0.0483425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_326_n 0.0152194f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=2.04
cc_64 VPB N_VPWR_c_327_n 0.0151082f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.225
cc_65 VPB N_VPWR_c_328_n 0.0327604f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=2.04
cc_66 VPB N_VPWR_c_329_n 0.0122846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_330_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_319_n 0.0440739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_X_c_378_n 0.0016834f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=1.515
cc_70 N_A_80_21#_c_72_n N_D1_M1003_g 0.00513349f $X=1.175 $Y=1.955 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_81_p N_D1_M1003_g 0.0148287f $X=1.905 $Y=2.04 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_74_n N_D1_M1003_g 0.00101167f $X=1.06 $Y=1.35 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_73_n N_D1_M1001_g 0.0119855f $X=1.64 $Y=0.42 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_74_n N_D1_M1001_g 0.00248384f $X=1.06 $Y=1.35 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_75_n N_D1_M1001_g 0.00668617f $X=1.175 $Y=1.225 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_72_n N_D1_c_153_n 0.0215464f $X=1.175 $Y=1.955 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_81_p N_D1_c_153_n 0.0257028f $X=1.905 $Y=2.04 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_74_n N_D1_c_153_n 4.40467e-19 $X=1.06 $Y=1.35 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_75_n N_D1_c_153_n 0.0284192f $X=1.175 $Y=1.225 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_72_n N_D1_c_151_n 0.00100627f $X=1.175 $Y=1.955 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_81_p N_D1_c_151_n 0.0011446f $X=1.905 $Y=2.04 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_74_n N_D1_c_151_n 0.0169524f $X=1.06 $Y=1.35 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_75_n N_D1_c_151_n 0.0103061f $X=1.175 $Y=1.225 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_94_p N_D1_c_151_n 8.17198e-19 $X=2 $Y=2.04 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_95_p N_C1_M1013_g 0.0115737f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_96_p N_C1_M1013_g 0.0124019f $X=2.865 $Y=2.04 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_94_p N_C1_M1013_g 4.2644e-19 $X=2 $Y=2.04 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_73_n C1 0.0450092f $X=1.64 $Y=0.42 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_75_n C1 0.0129191f $X=1.175 $Y=1.225 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_96_p C1 0.0138692f $X=2.865 $Y=2.04 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_94_p C1 0.0106087f $X=2 $Y=2.04 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_96_p N_C1_c_187_n 0.00262599f $X=2.865 $Y=2.04 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_73_n N_C1_c_188_n 0.00107601f $X=1.64 $Y=0.42 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_95_p N_B1_M1004_g 7.25236e-19 $X=2 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_96_p N_B1_M1004_g 0.0158773f $X=2.865 $Y=2.04 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_96_p B1 0.0196773f $X=2.865 $Y=2.04 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_107_p B1 0.0117185f $X=3.03 $Y=2.125 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_107_p N_B1_c_229_n 8.1826e-19 $X=3.03 $Y=2.125 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_72_n N_VPWR_M1012_d 0.00359679f $X=1.175 $Y=1.955 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_81_p N_VPWR_M1012_d 0.013799f $X=1.905 $Y=2.04 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_111_p N_VPWR_M1012_d 0.00689218f $X=1.305 $Y=2.04 $X2=0
+ $Y2=0
cc_102 N_A_80_21#_c_96_p N_VPWR_M1013_d 0.00891112f $X=2.865 $Y=2.04 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_76_n N_VPWR_c_321_n 0.00749164f $X=0.475 $Y=1.725 $X2=0
+ $Y2=0
cc_104 N_A_80_21#_c_76_n N_VPWR_c_322_n 6.74001e-19 $X=0.475 $Y=1.725 $X2=0
+ $Y2=0
cc_105 N_A_80_21#_c_77_n N_VPWR_c_322_n 0.0161815f $X=0.905 $Y=1.725 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_81_p N_VPWR_c_322_n 0.0300624f $X=1.905 $Y=2.04 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_111_p N_VPWR_c_322_n 0.0233519f $X=1.305 $Y=2.04 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_74_n N_VPWR_c_322_n 0.00173523f $X=1.06 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_96_p N_VPWR_c_323_n 0.022455f $X=2.865 $Y=2.04 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_76_n N_VPWR_c_326_n 0.00585385f $X=0.475 $Y=1.725 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_c_77_n N_VPWR_c_326_n 0.00564095f $X=0.905 $Y=1.725 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_c_95_p N_VPWR_c_327_n 0.0150063f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_123_p N_VPWR_c_328_n 0.0212513f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_114 N_A_80_21#_M1003_d N_VPWR_c_319_n 0.00380103f $X=1.86 $Y=1.835 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_M1004_d N_VPWR_c_319_n 0.00526034f $X=2.83 $Y=1.835 $X2=0
+ $Y2=0
cc_116 N_A_80_21#_c_76_n N_VPWR_c_319_n 0.011455f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_77_n N_VPWR_c_319_n 0.00948291f $X=0.905 $Y=1.725 $X2=0
+ $Y2=0
cc_118 N_A_80_21#_c_95_p N_VPWR_c_319_n 0.00950443f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_123_p N_VPWR_c_319_n 0.0127519f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_70_n N_X_c_378_n 0.00314492f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_76_n N_X_c_378_n 0.00337938f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_71_n N_X_c_378_n 0.00137547f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_77_n N_X_c_378_n 0.00163963f $X=0.905 $Y=1.725 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_72_n N_X_c_378_n 0.0218981f $X=1.175 $Y=1.955 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_74_n N_X_c_378_n 0.0469991f $X=1.06 $Y=1.35 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_75_n N_X_c_378_n 0.0342465f $X=1.175 $Y=1.225 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_75_n N_VGND_M1008_s 0.00230073f $X=1.175 $Y=1.225 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_c_70_n N_VGND_c_398_n 0.0071064f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_70_n N_VGND_c_399_n 6.17162e-19 $X=0.475 $Y=1.185 $X2=0
+ $Y2=0
cc_130 N_A_80_21#_c_71_n N_VGND_c_399_n 0.0100163f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A_80_21#_c_73_n N_VGND_c_399_n 0.0524466f $X=1.64 $Y=0.42 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_74_n N_VGND_c_399_n 0.00126616f $X=1.06 $Y=1.35 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_75_n N_VGND_c_399_n 0.022674f $X=1.175 $Y=1.225 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_70_n N_VGND_c_401_n 0.00585385f $X=0.475 $Y=1.185 $X2=0
+ $Y2=0
cc_135 N_A_80_21#_c_71_n N_VGND_c_401_n 0.00564095f $X=0.905 $Y=1.185 $X2=0
+ $Y2=0
cc_136 N_A_80_21#_c_73_n N_VGND_c_402_n 0.0224804f $X=1.64 $Y=0.42 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_70_n N_VGND_c_404_n 0.011455f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_71_n N_VGND_c_404_n 0.00948291f $X=0.905 $Y=1.185 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_c_73_n N_VGND_c_404_n 0.0134096f $X=1.64 $Y=0.42 $X2=0 $Y2=0
cc_140 N_D1_M1003_g N_C1_M1013_g 0.0176163f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_141 N_D1_M1001_g C1 0.00926873f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_142 N_D1_M1003_g C1 6.67239e-19 $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_143 N_D1_c_153_n C1 0.0288017f $X=1.64 $Y=1.51 $X2=0 $Y2=0
cc_144 N_D1_c_151_n C1 0.00393106f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_145 N_D1_c_153_n N_C1_c_187_n 3.20692e-19 $X=1.64 $Y=1.51 $X2=0 $Y2=0
cc_146 N_D1_c_151_n N_C1_c_187_n 0.0468042f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_147 N_D1_M1001_g N_C1_c_188_n 0.0468042f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_148 N_D1_M1003_g N_VPWR_c_322_n 0.0182543f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_149 N_D1_M1003_g N_VPWR_c_327_n 0.00486043f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_150 N_D1_M1003_g N_VPWR_c_319_n 0.0082726f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_151 N_D1_M1001_g N_VGND_c_399_n 0.00335405f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_152 N_D1_M1001_g N_VGND_c_402_n 0.00529818f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_153 N_D1_M1001_g N_VGND_c_404_n 0.0109271f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_154 C1 N_B1_M1006_g 0.00820107f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_155 N_C1_c_187_n N_B1_M1006_g 0.0214715f $X=2.305 $Y=1.37 $X2=0 $Y2=0
cc_156 N_C1_c_188_n N_B1_M1006_g 0.0301585f $X=2.305 $Y=1.205 $X2=0 $Y2=0
cc_157 N_C1_M1013_g B1 8.72081e-19 $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_158 C1 B1 0.0214993f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_159 N_C1_c_187_n B1 4.07101e-19 $X=2.305 $Y=1.37 $X2=0 $Y2=0
cc_160 N_C1_M1013_g N_B1_c_229_n 0.0367247f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_161 C1 N_B1_c_229_n 0.0014065f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_162 N_C1_M1013_g N_VPWR_c_322_n 7.36032e-19 $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_163 N_C1_M1013_g N_VPWR_c_323_n 0.00636535f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_164 N_C1_M1013_g N_VPWR_c_327_n 0.00564131f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_165 N_C1_M1013_g N_VPWR_c_319_n 0.0105297f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_166 C1 N_VGND_c_402_n 0.0132673f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_167 N_C1_c_188_n N_VGND_c_402_n 0.00364419f $X=2.305 $Y=1.205 $X2=0 $Y2=0
cc_168 C1 N_VGND_c_404_n 0.0131499f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_169 N_C1_c_188_n N_VGND_c_404_n 0.00537159f $X=2.305 $Y=1.205 $X2=0 $Y2=0
cc_170 C1 A_386_51# 0.00748401f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_171 C1 A_458_51# 0.0107478f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_172 C1 N_A_566_51#_c_449_n 0.00591424f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_173 N_B1_M1006_g N_A2_M1009_g 0.0230847f $X=2.755 $Y=0.675 $X2=0 $Y2=0
cc_174 N_B1_M1004_g N_A2_M1010_g 0.0251367f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_175 B1 N_A2_M1010_g 0.00108499f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_176 B1 A2 0.0214156f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_177 N_B1_c_229_n A2 3.12148e-19 $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_178 B1 N_A2_c_263_n 3.13256e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B1_c_229_n N_A2_c_263_n 0.0221755f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_180 N_B1_M1004_g N_VPWR_c_323_n 0.00420302f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B1_M1004_g N_VPWR_c_328_n 0.00585385f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B1_M1004_g N_VPWR_c_319_n 0.0112268f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B1_M1006_g N_VGND_c_402_n 0.00565115f $X=2.755 $Y=0.675 $X2=0 $Y2=0
cc_184 N_B1_M1006_g N_VGND_c_404_n 0.0112546f $X=2.755 $Y=0.675 $X2=0 $Y2=0
cc_185 N_B1_M1006_g N_A_566_51#_c_449_n 0.00206447f $X=2.755 $Y=0.675 $X2=0
+ $Y2=0
cc_186 B1 N_A_566_51#_c_449_n 0.0101785f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_187 N_B1_c_229_n N_A_566_51#_c_449_n 0.00362523f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A2_M1009_g N_A1_M1011_g 0.0243608f $X=3.295 $Y=0.675 $X2=0 $Y2=0
cc_189 N_A2_M1010_g N_A1_M1000_g 0.035618f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_190 A2 N_A1_M1000_g 0.00956472f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_191 A2 N_A1_c_296_n 0.0019107f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A2_c_263_n N_A1_c_296_n 0.0213742f $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_193 A2 N_A1_c_297_n 0.0263023f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A2_c_263_n N_A1_c_297_n 4.6215e-19 $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A2_M1010_g N_VPWR_c_325_n 0.00164342f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A2_M1010_g N_VPWR_c_328_n 0.00585385f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_197 A2 N_VPWR_c_328_n 0.0118455f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A2_M1010_g N_VPWR_c_319_n 0.0114286f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_199 A2 N_VPWR_c_319_n 0.0102675f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_200 A2 A_674_367# 0.0309051f $X=3.515 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_201 N_A2_M1009_g N_VGND_c_400_n 0.00325573f $X=3.295 $Y=0.675 $X2=0 $Y2=0
cc_202 N_A2_M1009_g N_VGND_c_402_n 0.00565115f $X=3.295 $Y=0.675 $X2=0 $Y2=0
cc_203 N_A2_M1009_g N_VGND_c_404_n 0.0110249f $X=3.295 $Y=0.675 $X2=0 $Y2=0
cc_204 N_A2_M1009_g N_A_566_51#_c_448_n 0.015298f $X=3.295 $Y=0.675 $X2=0 $Y2=0
cc_205 A2 N_A_566_51#_c_448_n 0.030133f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_206 N_A2_c_263_n N_A_566_51#_c_448_n 0.00429184f $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_207 N_A2_M1009_g N_A_566_51#_c_450_n 6.50435e-19 $X=3.295 $Y=0.675 $X2=0
+ $Y2=0
cc_208 N_A1_M1000_g N_VPWR_c_325_n 0.0227166f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A1_c_296_n N_VPWR_c_325_n 0.00163377f $X=4.05 $Y=1.46 $X2=0 $Y2=0
cc_210 N_A1_c_297_n N_VPWR_c_325_n 0.0261278f $X=4.05 $Y=1.46 $X2=0 $Y2=0
cc_211 N_A1_M1000_g N_VPWR_c_328_n 0.00486043f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A1_M1000_g N_VPWR_c_319_n 0.00864313f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A1_M1011_g N_VGND_c_400_n 0.00655853f $X=3.835 $Y=0.675 $X2=0 $Y2=0
cc_214 N_A1_M1011_g N_VGND_c_403_n 0.00529818f $X=3.835 $Y=0.675 $X2=0 $Y2=0
cc_215 N_A1_M1011_g N_VGND_c_404_n 0.0108401f $X=3.835 $Y=0.675 $X2=0 $Y2=0
cc_216 N_A1_M1011_g N_A_566_51#_c_448_n 0.0184008f $X=3.835 $Y=0.675 $X2=0 $Y2=0
cc_217 N_A1_c_296_n N_A_566_51#_c_448_n 0.00782521f $X=4.05 $Y=1.46 $X2=0 $Y2=0
cc_218 N_A1_c_297_n N_A_566_51#_c_448_n 0.0280151f $X=4.05 $Y=1.46 $X2=0 $Y2=0
cc_219 N_A1_M1011_g N_A_566_51#_c_450_n 0.0130628f $X=3.835 $Y=0.675 $X2=0 $Y2=0
cc_220 N_VPWR_c_319_n N_X_M1007_s 0.00345315f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_321_n N_X_c_378_n 0.00112943f $X=0.26 $Y=1.985 $X2=0 $Y2=0
cc_222 N_VPWR_c_326_n N_X_c_378_n 0.0144039f $X=0.975 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_319_n N_X_c_378_n 0.00944728f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_c_319_n A_674_367# 0.00713491f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_225 N_X_c_378_n N_VGND_c_398_n 0.0015328f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_226 N_X_c_378_n N_VGND_c_401_n 0.0144039f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_227 N_X_M1005_d N_VGND_c_404_n 0.00345315f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_228 N_X_c_378_n N_VGND_c_404_n 0.00944728f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_229 N_VGND_c_402_n N_A_566_51#_c_447_n 0.0212513f $X=3.385 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_404_n N_A_566_51#_c_447_n 0.0127519f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_M1009_d N_A_566_51#_c_448_n 0.0030319f $X=3.37 $Y=0.255 $X2=0
+ $Y2=0
cc_232 N_VGND_c_400_n N_A_566_51#_c_448_n 0.022455f $X=3.55 $Y=0.4 $X2=0 $Y2=0
cc_233 N_VGND_c_403_n N_A_566_51#_c_450_n 0.0210467f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_404_n N_A_566_51#_c_450_n 0.0126321f $X=4.08 $Y=0 $X2=0 $Y2=0
