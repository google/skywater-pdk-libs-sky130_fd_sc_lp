* NGSPICE file created from sky130_fd_sc_lp__or3b_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or3b_lp A B C_N VGND VNB VPB VPWR X
M1000 X a_350_47# a_804_101# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR C_N a_27_47# VPB phighvt w=1e+06u l=250000u
+  ad=6.75e+11p pd=5.35e+06u as=2.85e+11p ps=2.57e+06u
M1002 a_114_47# C_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1003 a_272_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.549e+11p ps=4.21e+06u
M1004 a_350_47# a_27_47# a_272_47# VNB nshort w=420000u l=150000u
+  ad=3.465e+11p pd=3.81e+06u as=0p ps=0u
M1005 VGND A a_640_101# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_350_47# B a_466_185# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_804_101# a_350_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_628_419# B a_263_373# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=5.7e+11p ps=5.14e+06u
M1009 a_466_185# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_350_47# a_27_47# a_263_373# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1011 X a_350_47# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1012 VPWR A a_628_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_640_101# A a_350_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C_N a_114_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

