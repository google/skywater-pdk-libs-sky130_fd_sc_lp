* File: sky130_fd_sc_lp__a311o_0.spice
* Created: Fri Aug 28 09:57:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311o_0.pex.spice"
.subckt sky130_fd_sc_lp__a311o_0  VNB VPB A3 A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_72_312#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1011 A_246_48# N_A3_M1011_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0819 PD=0.69 PS=0.81 NRD=22.848 NRS=11.424 M=1 R=2.8 SA=75000.7
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1009 A_330_48# N_A2_M1009_g A_246_48# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0567 PD=0.81 PS=0.69 NRD=39.996 NRS=22.848 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1001 N_A_72_312#_M1001_d N_A1_M1001_g A_330_48# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0819 PD=0.99 PS=0.81 NRD=75.708 NRS=39.996 M=1 R=2.8 SA=75001.7
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_B1_M1010_g N_A_72_312#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=0.99 NRD=0 NRS=7.14 M=1 R=2.8 SA=75002.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_72_312#_M1003_d N_C1_M1003_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_72_312#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_224_486#_M1008_d N_A3_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=12.2928 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_224_486#_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1984 AS=0.1024 PD=1.26 PS=0.96 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1007 N_A_224_486#_M1007_d N_A1_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1984 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.9 SB=75001 A=0.096 P=1.58 MULT=1
MM1002 A_558_486# N_B1_M1002_g N_A_224_486#_M1007_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_72_312#_M1000_d N_C1_M1000_g A_558_486# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75002.7
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a311o_0.pxi.spice"
*
.ends
*
*
