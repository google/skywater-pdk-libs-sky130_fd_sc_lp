* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111oi_lp A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VGND C1 a_553_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A1 a_131_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_125_57# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_553_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y D1 a_711_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y A1 a_125_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_131_409# B1 a_539_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_539_409# C1 a_637_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_637_409# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VGND B1 a_289_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_131_409# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_289_57# B1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_711_47# D1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
