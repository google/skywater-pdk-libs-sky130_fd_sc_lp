* File: sky130_fd_sc_lp__a32oi_m.pxi.spice
* Created: Fri Aug 28 10:02:15 2020
* 
x_PM_SKY130_FD_SC_LP__A32OI_M%B2 N_B2_c_71_n N_B2_c_72_n N_B2_c_73_n
+ N_B2_M1000_g N_B2_M1009_g N_B2_c_75_n N_B2_c_80_n B2 B2 B2 B2 B2 N_B2_c_77_n
+ PM_SKY130_FD_SC_LP__A32OI_M%B2
x_PM_SKY130_FD_SC_LP__A32OI_M%B1 N_B1_M1007_g N_B1_M1002_g N_B1_c_111_n
+ N_B1_c_116_n B1 B1 B1 B1 N_B1_c_113_n PM_SKY130_FD_SC_LP__A32OI_M%B1
x_PM_SKY130_FD_SC_LP__A32OI_M%A1 N_A1_M1001_g N_A1_M1003_g N_A1_c_158_n
+ N_A1_c_159_n N_A1_c_160_n A1 A1 A1 A1 A1 N_A1_c_162_n
+ PM_SKY130_FD_SC_LP__A32OI_M%A1
x_PM_SKY130_FD_SC_LP__A32OI_M%A2 N_A2_M1005_g N_A2_c_207_n N_A2_M1004_g
+ N_A2_c_211_n A2 A2 A2 A2 A2 N_A2_c_209_n PM_SKY130_FD_SC_LP__A32OI_M%A2
x_PM_SKY130_FD_SC_LP__A32OI_M%A3 N_A3_c_255_n N_A3_M1006_g N_A3_M1008_g
+ N_A3_c_256_n N_A3_c_261_n N_A3_c_262_n N_A3_c_257_n A3 A3 A3 A3 A3
+ N_A3_c_259_n PM_SKY130_FD_SC_LP__A32OI_M%A3
x_PM_SKY130_FD_SC_LP__A32OI_M%A_40_500# N_A_40_500#_M1000_s N_A_40_500#_M1002_d
+ N_A_40_500#_M1004_d N_A_40_500#_c_294_n N_A_40_500#_c_303_n
+ N_A_40_500#_c_295_n N_A_40_500#_c_296_n N_A_40_500#_c_325_p
+ N_A_40_500#_c_297_n PM_SKY130_FD_SC_LP__A32OI_M%A_40_500#
x_PM_SKY130_FD_SC_LP__A32OI_M%Y N_Y_M1007_d N_Y_M1000_d N_Y_c_330_n N_Y_c_335_n
+ N_Y_c_333_n N_Y_c_331_n Y PM_SKY130_FD_SC_LP__A32OI_M%Y
x_PM_SKY130_FD_SC_LP__A32OI_M%VPWR N_VPWR_M1003_d N_VPWR_M1008_d N_VPWR_c_371_n
+ N_VPWR_c_372_n VPWR N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n
+ N_VPWR_c_370_n N_VPWR_c_377_n N_VPWR_c_378_n PM_SKY130_FD_SC_LP__A32OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A32OI_M%VGND N_VGND_M1009_s N_VGND_M1006_d N_VGND_c_405_n
+ N_VGND_c_406_n N_VGND_c_407_n VGND N_VGND_c_408_n N_VGND_c_409_n
+ N_VGND_c_410_n N_VGND_c_411_n PM_SKY130_FD_SC_LP__A32OI_M%VGND
cc_1 VNB N_B2_c_71_n 0.0100006f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.14
cc_2 VNB N_B2_c_72_n 0.025849f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.915
cc_3 VNB N_B2_c_73_n 0.0232974f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.915
cc_4 VNB N_B2_M1009_g 0.0263686f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.445
cc_5 VNB N_B2_c_75_n 0.0248861f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_6 VNB B2 0.00741547f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_B2_c_77_n 0.0377367f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_8 VNB N_B1_M1007_g 0.0406381f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.915
cc_9 VNB N_B1_c_111_n 0.0186669f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.445
cc_10 VNB B1 0.00700825f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_11 VNB N_B1_c_113_n 0.0171259f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_A1_M1003_g 0.0108882f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.71
cc_13 VNB N_A1_c_158_n 0.0172649f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.84
cc_14 VNB N_A1_c_159_n 0.0243741f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.445
cc_15 VNB N_A1_c_160_n 0.0177567f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.445
cc_16 VNB A1 0.00250438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_162_n 0.0172381f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_18 VNB N_A2_M1005_g 0.0346911f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.915
cc_19 VNB N_A2_c_207_n 0.0242988f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.71
cc_20 VNB A2 0.00415876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_209_n 0.0195505f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_22 VNB N_A3_c_255_n 0.0207382f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.51
cc_23 VNB N_A3_c_256_n 0.0317145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A3_c_257_n 0.0369157f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.215
cc_25 VNB A3 0.0326811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A3_c_259_n 0.0180124f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_27 VNB N_Y_c_330_n 0.00455125f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.71
cc_28 VNB N_Y_c_331_n 0.00333004f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_29 VNB Y 0.014764f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.215
cc_30 VNB N_VPWR_c_370_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_31 VNB N_VGND_c_405_n 0.0125039f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.71
cc_32 VNB N_VGND_c_406_n 0.0155464f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.84
cc_33 VNB N_VGND_c_407_n 0.01277f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_34 VNB N_VGND_c_408_n 0.0558847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_409_n 0.0199636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_410_n 0.207008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_411_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_B2_c_71_n 0.0316504f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.14
cc_39 VPB N_B2_M1000_g 0.0228029f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=2.71
cc_40 VPB N_B2_c_80_n 0.0321856f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=2.215
cc_41 VPB B2 0.0327044f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_42 VPB N_B1_M1002_g 0.043204f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=2.71
cc_43 VPB N_B1_c_111_n 0.00571605f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.445
cc_44 VPB N_B1_c_116_n 0.0172188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB B1 0.00646977f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_46 VPB N_A1_M1003_g 0.0558851f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=2.71
cc_47 VPB A1 0.00482355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_M1004_g 0.0471947f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.84
cc_49 VPB N_A2_c_211_n 0.0187017f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.445
cc_50 VPB A2 0.0033052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A3_M1008_g 0.0304732f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=2.71
cc_52 VPB N_A3_c_261_n 0.0360365f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_53 VPB N_A3_c_262_n 0.0356417f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.215
cc_54 VPB A3 0.0156644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A3_c_259_n 0.00537119f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_56 VPB N_A_40_500#_c_294_n 0.00838459f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.445
cc_57 VPB N_A_40_500#_c_295_n 0.0233645f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.215
cc_58 VPB N_A_40_500#_c_296_n 0.00701731f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_40_500#_c_297_n 0.0190159f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_60 VPB N_Y_c_333_n 0.00474149f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.445
cc_61 VPB Y 0.0102527f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=2.215
cc_62 VPB N_VPWR_c_371_n 0.00763619f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.84
cc_63 VPB N_VPWR_c_372_n 0.0219404f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_64 VPB N_VPWR_c_373_n 0.0421572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_374_n 0.0184085f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_66 VPB N_VPWR_c_375_n 0.0174178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_370_n 0.0854682f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_68 VPB N_VPWR_c_377_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_69 VPB N_VPWR_c_378_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_70 N_B2_M1009_g N_B1_M1007_g 0.0548852f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_71 N_B2_c_77_n N_B1_M1007_g 0.00215545f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_72 N_B2_c_71_n N_B1_M1002_g 0.00199739f $X=0.36 $Y=2.14 $X2=0 $Y2=0
cc_73 N_B2_c_80_n N_B1_M1002_g 0.0256503f $X=0.62 $Y=2.215 $X2=0 $Y2=0
cc_74 N_B2_c_75_n N_B1_c_111_n 0.0039952f $X=0.27 $Y=1.51 $X2=0 $Y2=0
cc_75 N_B2_c_71_n N_B1_c_116_n 0.0039952f $X=0.36 $Y=2.14 $X2=0 $Y2=0
cc_76 N_B2_c_77_n N_B1_c_113_n 0.0039952f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_77 N_B2_M1000_g N_A_40_500#_c_294_n 0.0137004f $X=0.62 $Y=2.71 $X2=0 $Y2=0
cc_78 N_B2_M1000_g N_A_40_500#_c_297_n 0.00142375f $X=0.62 $Y=2.71 $X2=0 $Y2=0
cc_79 N_B2_c_80_n N_A_40_500#_c_297_n 0.00487736f $X=0.62 $Y=2.215 $X2=0 $Y2=0
cc_80 B2 N_A_40_500#_c_297_n 0.0159225f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_81 N_B2_M1009_g N_Y_c_335_n 0.012797f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_82 N_B2_M1000_g N_Y_c_333_n 0.0147553f $X=0.62 $Y=2.71 $X2=0 $Y2=0
cc_83 B2 N_Y_c_333_n 0.00997156f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_B2_c_72_n Y 0.00794884f $X=0.61 $Y=0.915 $X2=0 $Y2=0
cc_85 N_B2_M1009_g Y 0.0090935f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_86 N_B2_c_80_n Y 0.00595609f $X=0.62 $Y=2.215 $X2=0 $Y2=0
cc_87 B2 Y 0.0715848f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_88 N_B2_c_77_n Y 0.0085402f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_89 N_B2_M1000_g N_VPWR_c_373_n 9.21892e-19 $X=0.62 $Y=2.71 $X2=0 $Y2=0
cc_90 B2 N_VPWR_c_370_n 5.71109e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_91 N_B2_c_73_n N_VGND_c_406_n 0.00626709f $X=0.435 $Y=0.915 $X2=0 $Y2=0
cc_92 N_B2_M1009_g N_VGND_c_406_n 0.0131124f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_93 B2 N_VGND_c_406_n 0.00859099f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_94 N_B2_M1009_g N_VGND_c_408_n 0.00432572f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_95 N_B2_c_73_n N_VGND_c_410_n 0.00370238f $X=0.435 $Y=0.915 $X2=0 $Y2=0
cc_96 N_B2_M1009_g N_VGND_c_410_n 0.00757315f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_97 B2 N_VGND_c_410_n 9.40005e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_98 N_B1_M1002_g N_A1_M1003_g 0.0285531f $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_99 N_B1_c_111_n N_A1_M1003_g 0.02206f $X=1.07 $Y=1.735 $X2=0 $Y2=0
cc_100 B1 N_A1_M1003_g 0.00439794f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_101 N_B1_M1007_g N_A1_c_158_n 0.0286199f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_102 N_B1_c_113_n N_A1_c_159_n 0.00636699f $X=1.07 $Y=1.395 $X2=0 $Y2=0
cc_103 N_B1_c_111_n N_A1_c_160_n 0.00636699f $X=1.07 $Y=1.735 $X2=0 $Y2=0
cc_104 N_B1_M1007_g A1 0.00129287f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_105 N_B1_M1002_g A1 2.13949e-19 $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_106 B1 A1 0.0759032f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_107 N_B1_c_113_n A1 7.2391e-19 $X=1.07 $Y=1.395 $X2=0 $Y2=0
cc_108 B1 N_A1_c_162_n 0.00452869f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_109 N_B1_M1002_g N_A_40_500#_c_294_n 0.0139122f $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_110 N_B1_M1002_g N_A_40_500#_c_303_n 3.3835e-19 $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_111 N_B1_M1002_g N_A_40_500#_c_296_n 0.0015792f $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_112 N_B1_c_116_n N_A_40_500#_c_296_n 2.64202e-19 $X=1.07 $Y=1.9 $X2=0 $Y2=0
cc_113 B1 N_A_40_500#_c_296_n 0.00868207f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_114 N_B1_M1007_g N_Y_c_330_n 0.00913052f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_115 B1 N_Y_c_330_n 0.012183f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_116 N_B1_c_113_n N_Y_c_330_n 0.00187052f $X=1.07 $Y=1.395 $X2=0 $Y2=0
cc_117 N_B1_M1002_g N_Y_c_333_n 0.00790374f $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_118 N_B1_c_116_n N_Y_c_333_n 0.00247479f $X=1.07 $Y=1.9 $X2=0 $Y2=0
cc_119 B1 N_Y_c_333_n 0.00108947f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_120 B1 N_Y_c_331_n 0.0105926f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_121 N_B1_c_113_n N_Y_c_331_n 2.59481e-19 $X=1.07 $Y=1.395 $X2=0 $Y2=0
cc_122 N_B1_M1007_g Y 0.00729068f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B1_M1002_g Y 0.00653883f $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_124 B1 Y 0.0913326f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_125 N_B1_c_113_n Y 0.00656052f $X=1.07 $Y=1.395 $X2=0 $Y2=0
cc_126 N_B1_M1002_g N_VPWR_c_373_n 9.21892e-19 $X=1.05 $Y=2.71 $X2=0 $Y2=0
cc_127 N_B1_M1007_g N_VGND_c_408_n 0.00402178f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_128 N_B1_M1007_g N_VGND_c_410_n 0.00567203f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_129 B1 N_VGND_c_410_n 5.66395e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_130 N_A1_c_158_n N_A2_M1005_g 0.0202962f $X=1.61 $Y=0.765 $X2=0 $Y2=0
cc_131 A1 N_A2_M1005_g 0.00456955f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 N_A1_c_162_n N_A2_M1005_g 0.0133861f $X=1.61 $Y=0.93 $X2=0 $Y2=0
cc_133 N_A1_M1003_g N_A2_c_207_n 0.0124291f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_134 N_A1_c_160_n N_A2_c_207_n 0.0133861f $X=1.61 $Y=1.435 $X2=0 $Y2=0
cc_135 A1 N_A2_c_207_n 0.00318015f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_A1_M1003_g N_A2_M1004_g 0.0331113f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_137 A1 N_A2_M1004_g 0.00216718f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_138 N_A1_M1003_g A2 6.6191e-19 $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_139 N_A1_c_158_n A2 2.70084e-19 $X=1.61 $Y=0.765 $X2=0 $Y2=0
cc_140 A1 A2 0.074573f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A1_c_162_n A2 0.00205392f $X=1.61 $Y=0.93 $X2=0 $Y2=0
cc_142 N_A1_c_159_n N_A2_c_209_n 0.0133861f $X=1.61 $Y=1.27 $X2=0 $Y2=0
cc_143 N_A1_M1003_g N_A_40_500#_c_294_n 0.00149267f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_144 N_A1_M1003_g N_A_40_500#_c_303_n 0.00620893f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_145 N_A1_M1003_g N_A_40_500#_c_295_n 0.0134758f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_146 A1 N_A_40_500#_c_295_n 0.0169991f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_147 N_A1_M1003_g N_Y_c_333_n 2.71119e-19 $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_148 N_A1_c_158_n N_Y_c_331_n 0.00322885f $X=1.61 $Y=0.765 $X2=0 $Y2=0
cc_149 A1 N_Y_c_331_n 0.0132161f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_150 N_A1_M1003_g N_VPWR_c_371_n 0.00675938f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_151 N_A1_M1003_g N_VPWR_c_373_n 0.00455951f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_152 N_A1_M1003_g N_VPWR_c_370_n 0.00447788f $X=1.56 $Y=2.71 $X2=0 $Y2=0
cc_153 N_A1_c_158_n N_VGND_c_408_n 0.00499463f $X=1.61 $Y=0.765 $X2=0 $Y2=0
cc_154 A1 N_VGND_c_408_n 0.00601361f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A1_c_162_n N_VGND_c_408_n 6.70397e-19 $X=1.61 $Y=0.93 $X2=0 $Y2=0
cc_156 N_A1_c_158_n N_VGND_c_410_n 0.00896108f $X=1.61 $Y=0.765 $X2=0 $Y2=0
cc_157 A1 N_VGND_c_410_n 0.00778387f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_158 N_A1_c_162_n N_VGND_c_410_n 2.90533e-19 $X=1.61 $Y=0.93 $X2=0 $Y2=0
cc_159 A1 A_319_47# 0.0036712f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_160 N_A2_M1005_g N_A3_c_255_n 0.0500069f $X=2.06 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_161 A2 N_A3_c_255_n 0.00843278f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_162 N_A2_M1004_g N_A3_c_261_n 0.00615982f $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_163 N_A2_c_211_n N_A3_c_261_n 0.0118605f $X=2.155 $Y=1.825 $X2=0 $Y2=0
cc_164 A2 N_A3_c_261_n 8.77149e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_165 N_A2_M1004_g N_A3_c_262_n 0.0277796f $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_166 A2 N_A3_c_262_n 4.37285e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_167 N_A2_M1005_g N_A3_c_257_n 0.00591253f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_168 A2 N_A3_c_257_n 0.00164185f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_169 N_A2_c_209_n N_A3_c_257_n 0.0118605f $X=2.16 $Y=1.32 $X2=0 $Y2=0
cc_170 N_A2_M1005_g A3 8.44411e-19 $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_171 N_A2_M1004_g A3 0.0019424f $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_172 A2 A3 0.0624663f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_173 N_A2_c_209_n A3 0.0045679f $X=2.16 $Y=1.32 $X2=0 $Y2=0
cc_174 N_A2_c_207_n N_A3_c_259_n 0.0118605f $X=2.155 $Y=1.655 $X2=0 $Y2=0
cc_175 N_A2_M1004_g N_A_40_500#_c_295_n 0.0143365f $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_176 N_A2_c_211_n N_A_40_500#_c_295_n 0.0033194f $X=2.155 $Y=1.825 $X2=0 $Y2=0
cc_177 A2 N_A_40_500#_c_295_n 0.0123064f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_178 N_A2_M1004_g N_VPWR_c_371_n 0.00322432f $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_179 N_A2_M1004_g N_VPWR_c_372_n 7.06614e-19 $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_180 N_A2_M1004_g N_VPWR_c_374_n 0.00548708f $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_181 N_A2_M1004_g N_VPWR_c_370_n 0.00533081f $X=2.07 $Y=2.71 $X2=0 $Y2=0
cc_182 N_A2_M1005_g N_VGND_c_407_n 0.00232326f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_183 A2 N_VGND_c_407_n 8.92634e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_184 N_A2_M1005_g N_VGND_c_408_n 0.00511915f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_185 A2 N_VGND_c_408_n 0.00400372f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_186 N_A2_M1005_g N_VGND_c_410_n 0.00900763f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_187 A2 N_VGND_c_410_n 0.00544279f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_188 A2 A_427_47# 0.00279161f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_189 N_A3_M1008_g N_A_40_500#_c_295_n 0.00142609f $X=2.5 $Y=2.71 $X2=0 $Y2=0
cc_190 A3 N_A_40_500#_c_295_n 0.0132356f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_191 N_A3_M1008_g N_VPWR_c_372_n 0.00957179f $X=2.5 $Y=2.71 $X2=0 $Y2=0
cc_192 N_A3_c_262_n N_VPWR_c_372_n 0.003233f $X=2.66 $Y=2.215 $X2=0 $Y2=0
cc_193 A3 N_VPWR_c_372_n 0.0194467f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_194 N_A3_M1008_g N_VPWR_c_374_n 0.00455951f $X=2.5 $Y=2.71 $X2=0 $Y2=0
cc_195 N_A3_M1008_g N_VPWR_c_370_n 0.00447788f $X=2.5 $Y=2.71 $X2=0 $Y2=0
cc_196 A3 N_VPWR_c_370_n 9.58398e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_197 N_A3_c_255_n N_VGND_c_407_n 0.0112017f $X=2.42 $Y=0.765 $X2=0 $Y2=0
cc_198 N_A3_c_256_n N_VGND_c_407_n 0.00508284f $X=2.64 $Y=0.84 $X2=0 $Y2=0
cc_199 A3 N_VGND_c_407_n 0.0108979f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_200 N_A3_c_255_n N_VGND_c_408_n 0.00486043f $X=2.42 $Y=0.765 $X2=0 $Y2=0
cc_201 N_A3_c_255_n N_VGND_c_410_n 0.00818711f $X=2.42 $Y=0.765 $X2=0 $Y2=0
cc_202 A3 N_VGND_c_410_n 0.00180401f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_203 N_A_40_500#_c_294_n N_Y_M1000_d 0.00180746f $X=1.18 $Y=2.975 $X2=0 $Y2=0
cc_204 N_A_40_500#_c_294_n N_Y_c_333_n 0.0160841f $X=1.18 $Y=2.975 $X2=0 $Y2=0
cc_205 N_A_40_500#_c_303_n N_Y_c_333_n 0.00822738f $X=1.285 $Y=2.645 $X2=0 $Y2=0
cc_206 N_A_40_500#_c_296_n N_Y_c_333_n 0.0138775f $X=1.39 $Y=2.405 $X2=0 $Y2=0
cc_207 N_A_40_500#_c_294_n N_VPWR_c_371_n 0.0118055f $X=1.18 $Y=2.975 $X2=0
+ $Y2=0
cc_208 N_A_40_500#_c_303_n N_VPWR_c_371_n 0.0135009f $X=1.285 $Y=2.645 $X2=0
+ $Y2=0
cc_209 N_A_40_500#_c_295_n N_VPWR_c_371_n 0.0226391f $X=2.2 $Y=2.405 $X2=0 $Y2=0
cc_210 N_A_40_500#_c_294_n N_VPWR_c_373_n 0.0543661f $X=1.18 $Y=2.975 $X2=0
+ $Y2=0
cc_211 N_A_40_500#_c_297_n N_VPWR_c_373_n 0.0206108f $X=0.325 $Y=2.775 $X2=0
+ $Y2=0
cc_212 N_A_40_500#_c_325_p N_VPWR_c_374_n 0.00412673f $X=2.285 $Y=2.645 $X2=0
+ $Y2=0
cc_213 N_A_40_500#_c_294_n N_VPWR_c_370_n 0.0338106f $X=1.18 $Y=2.975 $X2=0
+ $Y2=0
cc_214 N_A_40_500#_c_295_n N_VPWR_c_370_n 0.0167623f $X=2.2 $Y=2.405 $X2=0 $Y2=0
cc_215 N_A_40_500#_c_325_p N_VPWR_c_370_n 0.00545208f $X=2.285 $Y=2.645 $X2=0
+ $Y2=0
cc_216 N_A_40_500#_c_297_n N_VPWR_c_370_n 0.0124745f $X=0.325 $Y=2.775 $X2=0
+ $Y2=0
cc_217 N_Y_c_330_n N_VGND_c_408_n 0.00744054f $X=1.155 $Y=0.575 $X2=0 $Y2=0
cc_218 N_Y_c_335_n N_VGND_c_408_n 0.00389f $X=0.805 $Y=0.575 $X2=0 $Y2=0
cc_219 N_Y_c_331_n N_VGND_c_408_n 0.0080317f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_220 N_Y_M1007_d N_VGND_c_410_n 0.00621794f $X=1.12 $Y=0.235 $X2=0 $Y2=0
cc_221 N_Y_c_330_n N_VGND_c_410_n 0.0104212f $X=1.155 $Y=0.575 $X2=0 $Y2=0
cc_222 N_Y_c_335_n N_VGND_c_410_n 0.00509672f $X=0.805 $Y=0.575 $X2=0 $Y2=0
cc_223 N_Y_c_331_n N_VGND_c_410_n 0.00687036f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_224 N_Y_c_330_n A_152_47# 0.00137964f $X=1.155 $Y=0.575 $X2=-0.19 $Y2=-0.245
cc_225 N_VGND_c_410_n A_152_47# 0.00203487f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_226 N_VGND_c_410_n A_319_47# 0.0108187f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_227 N_VGND_c_410_n A_427_47# 0.00535573f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
