* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 a_776_99# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR a_626_125# a_776_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_31_464# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_31_464# a_554_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_776_99# a_626_125# a_996_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_31_464# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_996_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_554_125# a_221_70# a_626_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_776_99# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 Q a_776_99# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND GATE_N a_221_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_726_125# a_776_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_776_99# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_626_125# a_372_397# a_726_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_626_125# a_221_70# a_763_473# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_763_473# a_776_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VPWR a_31_464# a_582_473# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_582_473# a_372_397# a_626_125# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_372_397# a_221_70# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR GATE_N a_221_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_372_397# a_221_70# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 Q a_776_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
