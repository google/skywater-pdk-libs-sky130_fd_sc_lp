* File: sky130_fd_sc_lp__nand3_4.pex.spice
* Created: Fri Aug 28 10:49:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3_4%A 3 7 11 15 19 23 27 31 33 34 35 51
c77 51 0 2.34486e-19 $X=1.795 $Y=1.51
c78 27 0 5.94179e-20 $X=1.795 $Y=0.705
r79 51 52 2.94801 $w=3.27e-07 $l=2e-08 $layer=POLY_cond $X=1.795 $Y=1.51
+ $X2=1.815 $Y2=1.51
r80 50 51 60.4342 $w=3.27e-07 $l=4.1e-07 $layer=POLY_cond $X=1.385 $Y=1.51
+ $X2=1.795 $Y2=1.51
r81 49 50 2.94801 $w=3.27e-07 $l=2e-08 $layer=POLY_cond $X=1.365 $Y=1.51
+ $X2=1.385 $Y2=1.51
r82 47 49 32.4281 $w=3.27e-07 $l=2.2e-07 $layer=POLY_cond $X=1.145 $Y=1.51
+ $X2=1.365 $Y2=1.51
r83 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.145
+ $Y=1.51 $X2=1.145 $Y2=1.51
r84 45 47 28.0061 $w=3.27e-07 $l=1.9e-07 $layer=POLY_cond $X=0.955 $Y=1.51
+ $X2=1.145 $Y2=1.51
r85 44 45 2.94801 $w=3.27e-07 $l=2e-08 $layer=POLY_cond $X=0.935 $Y=1.51
+ $X2=0.955 $Y2=1.51
r86 43 44 60.4342 $w=3.27e-07 $l=4.1e-07 $layer=POLY_cond $X=0.525 $Y=1.51
+ $X2=0.935 $Y2=1.51
r87 42 43 2.94801 $w=3.27e-07 $l=2e-08 $layer=POLY_cond $X=0.505 $Y=1.51
+ $X2=0.525 $Y2=1.51
r88 40 42 5.89602 $w=3.27e-07 $l=4e-08 $layer=POLY_cond $X=0.465 $Y=1.51
+ $X2=0.505 $Y2=1.51
r89 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.465
+ $Y=1.51 $X2=0.465 $Y2=1.51
r90 35 48 1.78548 $w=3.53e-07 $l=5.5e-08 $layer=LI1_cond $X=1.2 $Y=1.572
+ $X2=1.145 $Y2=1.572
r91 34 48 13.7969 $w=3.53e-07 $l=4.25e-07 $layer=LI1_cond $X=0.72 $Y=1.572
+ $X2=1.145 $Y2=1.572
r92 34 41 8.27811 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.72 $Y=1.572
+ $X2=0.465 $Y2=1.572
r93 33 41 7.30422 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=0.24 $Y=1.572
+ $X2=0.465 $Y2=1.572
r94 29 52 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.675
+ $X2=1.815 $Y2=1.51
r95 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.815 $Y=1.675
+ $X2=1.815 $Y2=2.465
r96 25 51 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.345
+ $X2=1.795 $Y2=1.51
r97 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.795 $Y=1.345
+ $X2=1.795 $Y2=0.705
r98 21 50 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.675
+ $X2=1.385 $Y2=1.51
r99 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.385 $Y=1.675
+ $X2=1.385 $Y2=2.465
r100 17 49 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.345
+ $X2=1.365 $Y2=1.51
r101 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.365 $Y=1.345
+ $X2=1.365 $Y2=0.705
r102 13 45 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=1.51
r103 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=2.465
r104 9 44 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.345
+ $X2=0.935 $Y2=1.51
r105 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.935 $Y=1.345
+ $X2=0.935 $Y2=0.705
r106 5 43 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.675
+ $X2=0.525 $Y2=1.51
r107 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.525 $Y=1.675
+ $X2=0.525 $Y2=2.465
r108 1 42 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.345
+ $X2=0.505 $Y2=1.51
r109 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.505 $Y=1.345
+ $X2=0.505 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_4%B 3 7 11 15 19 23 27 31 33 38 39 41 45 47 48
+ 51 52 53 54 55 66
c126 39 0 2.39085e-19 $X=2.987 $Y=1.92
c127 33 0 1.73689e-19 $X=2.795 $Y=1.515
c128 23 0 1.26098e-19 $X=3.105 $Y=2.465
r129 62 63 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=2.245 $Y=1.51
+ $X2=2.655 $Y2=1.51
r130 60 62 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.225 $Y=1.51
+ $X2=2.245 $Y2=1.51
r131 54 55 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=2.02
+ $X2=5.04 $Y2=2.02
r132 53 54 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=2.02
+ $X2=4.56 $Y2=2.02
r133 52 53 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=2.02
+ $X2=4.08 $Y2=2.02
r134 51 55 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=5.2 $Y=2.02
+ $X2=5.04 $Y2=2.02
r135 48 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.375 $Y=1.51
+ $X2=5.375 $Y2=1.675
r136 48 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.375 $Y=1.51
+ $X2=5.375 $Y2=1.345
r137 47 50 7.82185 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=5.37 $Y=1.51
+ $X2=5.37 $Y2=1.705
r138 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.375
+ $Y=1.51 $X2=5.375 $Y2=1.51
r139 45 52 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=3.18 $Y=2.02
+ $X2=3.6 $Y2=2.02
r140 44 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.015 $Y=1.51
+ $X2=3.105 $Y2=1.51
r141 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.015
+ $Y=1.51 $X2=3.015 $Y2=1.51
r142 41 51 6.85974 $w=2e-07 $l=1.57242e-07 $layer=LI1_cond $X=5.315 $Y=1.92
+ $X2=5.2 $Y2=2.02
r143 41 50 10.7728 $w=2.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.315 $Y=1.92
+ $X2=5.315 $Y2=1.705
r144 39 45 7.74296 $w=2e-07 $l=2.378e-07 $layer=LI1_cond $X=2.987 $Y=1.92
+ $X2=3.18 $Y2=2.02
r145 38 43 2.57054 $w=3.85e-07 $l=9e-08 $layer=LI1_cond $X=2.987 $Y=1.605
+ $X2=2.987 $Y2=1.515
r146 38 39 9.42908 $w=3.83e-07 $l=3.15e-07 $layer=LI1_cond $X=2.987 $Y=1.605
+ $X2=2.987 $Y2=1.92
r147 36 44 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.675 $Y=1.51
+ $X2=3.015 $Y2=1.51
r148 36 63 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.675 $Y=1.51
+ $X2=2.655 $Y2=1.51
r149 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.675
+ $Y=1.51 $X2=2.675 $Y2=1.51
r150 33 43 5.48382 $w=1.8e-07 $l=1.92e-07 $layer=LI1_cond $X=2.795 $Y=1.515
+ $X2=2.987 $Y2=1.515
r151 33 35 7.39394 $w=1.78e-07 $l=1.2e-07 $layer=LI1_cond $X=2.795 $Y=1.515
+ $X2=2.675 $Y2=1.515
r152 31 70 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.285 $Y=2.465
+ $X2=5.285 $Y2=1.675
r153 27 69 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.285 $Y=0.705
+ $X2=5.285 $Y2=1.345
r154 21 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.675
+ $X2=3.105 $Y2=1.51
r155 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.105 $Y=1.675
+ $X2=3.105 $Y2=2.465
r156 17 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.345
+ $X2=3.105 $Y2=1.51
r157 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.105 $Y=1.345
+ $X2=3.105 $Y2=0.705
r158 13 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.675
+ $X2=2.675 $Y2=1.51
r159 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.675 $Y=1.675
+ $X2=2.675 $Y2=2.465
r160 9 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.345
+ $X2=2.655 $Y2=1.51
r161 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.655 $Y=1.345
+ $X2=2.655 $Y2=0.705
r162 5 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.245 $Y=1.675
+ $X2=2.245 $Y2=1.51
r163 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.245 $Y=1.675
+ $X2=2.245 $Y2=2.465
r164 1 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.345
+ $X2=2.225 $Y2=1.51
r165 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.225 $Y=1.345
+ $X2=2.225 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_4%C 3 7 11 15 19 23 27 31 33 34 35 52 53
c83 53 0 8.67609e-20 $X=4.855 $Y=1.51
c84 27 0 1.27067e-19 $X=4.855 $Y=0.705
c85 11 0 5.9075e-20 $X=3.995 $Y=0.705
c86 7 0 1.26355e-19 $X=3.565 $Y=0.705
r87 51 53 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=4.575 $Y=1.51
+ $X2=4.855 $Y2=1.51
r88 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=1.51 $X2=4.575 $Y2=1.51
r89 49 51 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.425 $Y=1.51
+ $X2=4.575 $Y2=1.51
r90 47 49 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.235 $Y=1.51
+ $X2=4.425 $Y2=1.51
r91 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.235
+ $Y=1.51 $X2=4.235 $Y2=1.51
r92 45 47 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.995 $Y=1.51
+ $X2=4.235 $Y2=1.51
r93 43 45 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.895 $Y=1.51
+ $X2=3.995 $Y2=1.51
r94 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.895
+ $Y=1.51 $X2=3.895 $Y2=1.51
r95 41 43 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.565 $Y=1.51
+ $X2=3.895 $Y2=1.51
r96 39 41 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.535 $Y=1.51
+ $X2=3.565 $Y2=1.51
r97 35 52 0.531897 $w=3.23e-07 $l=1.5e-08 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.575 $Y2=1.587
r98 35 48 11.5244 $w=3.23e-07 $l=3.25e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.235 $Y2=1.587
r99 34 48 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.235 $Y2=1.587
r100 34 44 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=3.895 $Y2=1.587
r101 33 44 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=3.6 $Y=1.587
+ $X2=3.895 $Y2=1.587
r102 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.675
+ $X2=4.855 $Y2=1.51
r103 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.855 $Y=1.675
+ $X2=4.855 $Y2=2.465
r104 25 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.345
+ $X2=4.855 $Y2=1.51
r105 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.855 $Y=1.345
+ $X2=4.855 $Y2=0.705
r106 21 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.675
+ $X2=4.425 $Y2=1.51
r107 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.425 $Y=1.675
+ $X2=4.425 $Y2=2.465
r108 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.345
+ $X2=4.425 $Y2=1.51
r109 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.425 $Y=1.345
+ $X2=4.425 $Y2=0.705
r110 13 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.675
+ $X2=3.995 $Y2=1.51
r111 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.995 $Y=1.675
+ $X2=3.995 $Y2=2.465
r112 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.345
+ $X2=3.995 $Y2=1.51
r113 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.995 $Y=1.345
+ $X2=3.995 $Y2=0.705
r114 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.345
+ $X2=3.565 $Y2=1.51
r115 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.565 $Y=1.345
+ $X2=3.565 $Y2=0.705
r116 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.675
+ $X2=3.535 $Y2=1.51
r117 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.535 $Y=1.675
+ $X2=3.535 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 40 42 46 50
+ 52 54 57 58 59 60 61 63 75 80 89 92 95 99
c109 4 0 1.52324e-19 $X=2.75 $Y=1.835
r110 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r111 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r114 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r115 84 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r116 84 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 81 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=3.33
+ $X2=4.64 $Y2=3.33
r119 81 83 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.805 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 80 98 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=5.335 $Y=3.33
+ $X2=5.547 $Y2=3.33
r121 80 83 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 79 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r123 79 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 76 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=3.75 $Y2=3.33
r126 76 78 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=4.08 $Y2=3.33
r127 75 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.64 $Y2=3.33
r128 75 78 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r130 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r131 71 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 68 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r134 68 70 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r135 67 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 67 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 64 86 4.66755 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.237 $Y2=3.33
r139 64 66 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 63 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r141 63 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r142 61 93 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 61 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r144 59 73 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.64 $Y2=3.33
r145 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.89 $Y2=3.33
r146 57 70 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.68 $Y2=3.33
r147 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.03 $Y2=3.33
r148 56 73 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.64 $Y2=3.33
r149 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.03 $Y2=3.33
r150 52 98 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=5.5 $Y=3.245
+ $X2=5.547 $Y2=3.33
r151 52 54 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=5.5 $Y=3.245
+ $X2=5.5 $Y2=2.375
r152 48 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=3.245
+ $X2=4.64 $Y2=3.33
r153 48 50 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.64 $Y=3.245
+ $X2=4.64 $Y2=2.755
r154 44 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=3.245
+ $X2=3.75 $Y2=3.33
r155 44 46 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=3.75 $Y=3.245
+ $X2=3.75 $Y2=2.755
r156 43 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=2.89 $Y2=3.33
r157 42 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=3.75 $Y2=3.33
r158 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=3.055 $Y2=3.33
r159 38 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=3.245
+ $X2=2.89 $Y2=3.33
r160 38 40 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.89 $Y=3.245
+ $X2=2.89 $Y2=2.755
r161 34 37 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.03 $Y=2.2
+ $X2=2.03 $Y2=2.97
r162 32 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=3.33
r163 32 37 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=2.97
r164 28 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r165 28 30 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.355
r166 24 27 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.31 $Y=2.005
+ $X2=0.31 $Y2=2.95
r167 22 86 3.09863 $w=3.3e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.237 $Y2=3.33
r168 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.31 $Y2=2.95
r169 7 54 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=2.375
r170 6 50 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=1.835 $X2=4.64 $Y2=2.755
r171 5 46 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=1.835 $X2=3.75 $Y2=2.755
r172 4 40 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=2.75
+ $Y=1.835 $X2=2.89 $Y2=2.755
r173 3 37 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.835 $X2=2.03 $Y2=2.97
r174 3 34 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.835 $X2=2.03 $Y2=2.2
r175 2 30 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.355
r176 1 27 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.95
r177 1 24 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_4%Y 1 2 3 4 5 6 7 8 27 29 31 33 34 35 39 42 43
+ 45 47 52 55 59 63 69 71 73 75 77 78
c101 47 0 1.26098e-19 $X=2.365 $Y=1.86
r102 78 82 5.48157 $w=4.34e-07 $l=1.95e-07 $layer=LI1_cond $X=1.747 $Y=1.665
+ $X2=1.747 $Y2=1.86
r103 64 75 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.305 $Y=2.375
+ $X2=4.205 $Y2=2.375
r104 63 77 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.975 $Y=2.375
+ $X2=5.07 $Y2=2.375
r105 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=2.375
+ $X2=4.305 $Y2=2.375
r106 60 73 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.415 $Y=2.375
+ $X2=3.32 $Y2=2.375
r107 59 75 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.105 $Y=2.375
+ $X2=4.205 $Y2=2.375
r108 59 60 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.105 $Y=2.375
+ $X2=3.415 $Y2=2.375
r109 56 71 2.28545 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.625 $Y=2.375
+ $X2=2.495 $Y2=2.375
r110 55 73 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.225 $Y=2.375
+ $X2=3.32 $Y2=2.375
r111 55 56 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.225 $Y=2.375
+ $X2=2.625 $Y2=2.375
r112 50 71 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=2.29
+ $X2=2.495 $Y2=2.375
r113 50 52 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=2.495 $Y=2.29
+ $X2=2.495 $Y2=1.98
r114 49 52 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=2.495 $Y=1.945
+ $X2=2.495 $Y2=1.98
r115 48 82 6.27713 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=2 $Y=1.86 $X2=1.747
+ $Y2=1.86
r116 47 49 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.365 $Y=1.86
+ $X2=2.495 $Y2=1.945
r117 47 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.365 $Y=1.86
+ $X2=2 $Y2=1.86
r118 43 85 4.34317 $w=4.34e-07 $l=1.5e-08 $layer=LI1_cond $X=1.6 $Y=2.1 $X2=1.6
+ $Y2=2.085
r119 43 45 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=1.6 $Y=2.1 $X2=1.6
+ $Y2=2.91
r120 42 78 9.85388 $w=4.34e-07 $l=3.03974e-07 $layer=LI1_cond $X=1.602 $Y=1.425
+ $X2=1.747 $Y2=1.665
r121 41 69 4.14756 $w=2.2e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.602 $Y=1.225
+ $X2=1.597 $Y2=1.14
r122 41 42 10.7204 $w=2.13e-07 $l=2e-07 $layer=LI1_cond $X=1.602 $Y=1.225
+ $X2=1.602 $Y2=1.425
r123 37 69 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.597 $Y=1.055
+ $X2=1.597 $Y2=1.14
r124 37 39 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.597 $Y=1.055
+ $X2=1.597 $Y2=0.76
r125 36 68 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=0.835 $Y=2.01
+ $X2=0.74 $Y2=2.01
r126 35 85 2.10829 $w=4.34e-07 $l=1.37477e-07 $layer=LI1_cond $X=1.495 $Y=2.01
+ $X2=1.6 $Y2=2.085
r127 35 82 4.21659 $w=4.34e-07 $l=3.18283e-07 $layer=LI1_cond $X=1.495 $Y=2.01
+ $X2=1.747 $Y2=1.86
r128 35 36 40.6667 $w=1.78e-07 $l=6.6e-07 $layer=LI1_cond $X=1.495 $Y=2.01
+ $X2=0.835 $Y2=2.01
r129 33 69 2.28545 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.485 $Y=1.14
+ $X2=1.597 $Y2=1.14
r130 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.485 $Y=1.14
+ $X2=0.815 $Y2=1.14
r131 29 68 3.31928 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=0.74 $Y=2.1 $X2=0.74
+ $Y2=2.01
r132 29 31 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=0.74 $Y=2.1
+ $X2=0.74 $Y2=2.91
r133 25 34 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.705 $Y=1.055
+ $X2=0.815 $Y2=1.14
r134 25 27 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=1.055
+ $X2=0.705 $Y2=0.76
r135 8 77 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=4.93
+ $Y=1.835 $X2=5.07 $Y2=2.455
r136 7 75 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=4.07
+ $Y=1.835 $X2=4.21 $Y2=2.455
r137 6 73 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=3.18
+ $Y=1.835 $X2=3.32 $Y2=2.455
r138 5 71 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.455
r139 5 52 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=1.98
r140 4 85 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.085
r141 4 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.91
r142 3 68 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=2.085
r143 3 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=2.91
r144 2 39 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.285 $X2=1.58 $Y2=0.76
r145 1 27 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.285 $X2=0.72 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_4%A_33_57# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 42 44 45
c84 33 0 6.07968e-20 $X=2.105 $Y=1.17
r85 40 42 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=5.535 $Y=1.085
+ $X2=5.535 $Y2=0.43
r86 39 45 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=1.17
+ $X2=2.89 $Y2=1.17
r87 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.405 $Y=1.17
+ $X2=5.535 $Y2=1.085
r88 38 39 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.405 $Y=1.17
+ $X2=3.005 $Y2=1.17
r89 34 45 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=1.085
+ $X2=2.89 $Y2=1.17
r90 34 36 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.89 $Y=1.085
+ $X2=2.89 $Y2=0.81
r91 32 45 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.775 $Y=1.17
+ $X2=2.89 $Y2=1.17
r92 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.775 $Y=1.17
+ $X2=2.105 $Y2=1.17
r93 29 33 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.992 $Y=1.085
+ $X2=2.105 $Y2=1.17
r94 29 31 33.5489 $w=2.23e-07 $l=6.55e-07 $layer=LI1_cond $X=1.992 $Y=1.085
+ $X2=1.992 $Y2=0.43
r95 28 31 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=1.992 $Y=0.425
+ $X2=1.992 $Y2=0.43
r96 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0.34
+ $X2=1.15 $Y2=0.34
r97 26 28 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.88 $Y=0.34
+ $X2=1.992 $Y2=0.425
r98 26 27 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.88 $Y=0.34
+ $X2=1.315 $Y2=0.34
r99 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.425
+ $X2=1.15 $Y2=0.34
r100 22 24 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=0.425
+ $X2=1.15 $Y2=0.43
r101 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0.34
+ $X2=1.15 $Y2=0.34
r102 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.34
+ $X2=0.425 $Y2=0.34
r103 16 21 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.275 $Y=0.425
+ $X2=0.425 $Y2=0.34
r104 16 18 0.192074 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=0.275 $Y=0.425
+ $X2=0.275 $Y2=0.43
r105 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.285 $X2=5.5 $Y2=0.43
r106 4 36 182 $w=1.7e-07 $l=5.99687e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.285 $X2=2.89 $Y2=0.81
r107 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.285 $X2=2.01 $Y2=0.43
r108 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.285 $X2=1.15 $Y2=0.43
r109 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.285 $X2=0.29 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_4%A_460_57# 1 2 3 4 15 17 18 19 20 22 29 30 32
+ 33
c58 30 0 2.53422e-19 $X=4.355 $Y=0.807
c59 19 0 5.9075e-20 $X=3.34 $Y=0.425
c60 18 0 5.94179e-20 $X=2.605 $Y=0.34
r61 32 33 8.04147 $w=2.13e-07 $l=1.4e-07 $layer=LI1_cond $X=5.07 $Y=0.807
+ $X2=4.93 $Y2=0.807
r62 30 33 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.355 $Y=0.83
+ $X2=4.93 $Y2=0.83
r63 28 30 8.30948 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=4.21 $Y=0.807
+ $X2=4.355 $Y2=0.807
r64 28 29 8.30948 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=4.21 $Y=0.807
+ $X2=4.065 $Y2=0.807
r65 22 29 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.505 $Y=0.83
+ $X2=4.065 $Y2=0.83
r66 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.34 $Y=0.745
+ $X2=3.505 $Y2=0.83
r67 19 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.34 $Y=0.425 $X2=3.34
+ $Y2=0.34
r68 19 20 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.34 $Y=0.425
+ $X2=3.34 $Y2=0.745
r69 17 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=0.34
+ $X2=3.34 $Y2=0.34
r70 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.175 $Y=0.34
+ $X2=2.605 $Y2=0.34
r71 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.44 $Y=0.425
+ $X2=2.605 $Y2=0.34
r72 13 15 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.44 $Y=0.425
+ $X2=2.44 $Y2=0.43
r73 4 32 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.285 $X2=5.07 $Y2=0.83
r74 3 28 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=4.07
+ $Y=0.285 $X2=4.21 $Y2=0.83
r75 2 26 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=3.18
+ $Y=0.285 $X2=3.34 $Y2=0.42
r76 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.285 $X2=2.44 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_4%VGND 1 2 9 13 16 17 18 27 33 34 37
r73 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r74 34 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r75 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r76 31 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.64
+ $Y2=0
r77 31 33 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=5.52
+ $Y2=0
r78 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r79 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r80 27 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.64
+ $Y2=0
r81 27 29 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.08
+ $Y2=0
r82 26 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r83 25 26 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r84 21 25 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r85 21 22 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r86 18 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r87 18 22 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.24
+ $Y2=0
r88 16 25 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.6
+ $Y2=0
r89 16 17 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.81
+ $Y2=0
r90 15 29 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=4.08
+ $Y2=0
r91 15 17 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=3.81
+ $Y2=0
r92 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r93 11 13 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.47
r94 7 17 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=0.085
+ $X2=3.81 $Y2=0
r95 7 9 13.872 $w=2.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.81 $Y=0.085 $X2=3.81
+ $Y2=0.41
r96 2 13 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.5
+ $Y=0.285 $X2=4.64 $Y2=0.47
r97 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.285 $X2=3.78 $Y2=0.41
.ends

