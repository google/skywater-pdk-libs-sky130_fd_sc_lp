* File: sky130_fd_sc_lp__o211ai_m.pex.spice
* Created: Fri Aug 28 11:03:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211AI_M%A1 3 7 11 15 17 18 19 20 26
c32 26 0 1.81115e-19 $X=0.385 $Y=1.49
c33 11 0 1.64738e-19 $X=0.39 $Y=1.475
r34 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.49 $X2=0.385 $Y2=1.49
r35 19 20 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=2.035
+ $X2=0.312 $Y2=2.405
r36 18 19 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=2.035
r37 18 27 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=1.49
r38 17 27 7.13417 $w=3.13e-07 $l=1.95e-07 $layer=LI1_cond $X=0.312 $Y=1.295
+ $X2=0.312 $Y2=1.49
r39 13 26 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.385 $Y=1.845
+ $X2=0.385 $Y2=1.49
r40 13 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.385 $Y=1.92
+ $X2=0.665 $Y2=1.92
r41 11 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.385 $Y=1.475
+ $X2=0.385 $Y2=1.49
r42 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.39 $Y=1.325
+ $X2=0.39 $Y2=1.475
r43 5 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=1.995
+ $X2=0.665 $Y2=1.92
r44 5 7 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.665 $Y=1.995
+ $X2=0.665 $Y2=2.885
r45 3 10 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.485 $Y=0.445
+ $X2=0.485 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_M%A2 3 7 11 12 13 16
c42 13 0 1.81115e-19 $X=1.2 $Y=1.295
r43 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.935
+ $Y=1.1 $X2=0.935 $Y2=1.1
r44 13 17 6.21492 $w=5.08e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=1.27
+ $X2=0.935 $Y2=1.27
r45 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.935 $Y=1.44
+ $X2=0.935 $Y2=1.1
r46 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.44
+ $X2=0.935 $Y2=1.605
r47 10 16 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=0.935
+ $X2=0.935 $Y2=1.1
r48 7 12 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=1.025 $Y=2.885
+ $X2=1.025 $Y2=1.605
r49 3 10 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.955 $Y=0.445
+ $X2=0.955 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_M%B1 3 7 11 12 13 16
c45 3 0 9.23808e-20 $X=1.385 $Y=0.445
r46 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.475
+ $Y=1.79 $X2=1.475 $Y2=1.79
r47 13 17 4.80777 $w=5.08e-07 $l=2.05e-07 $layer=LI1_cond $X=1.68 $Y=1.96
+ $X2=1.475 $Y2=1.96
r48 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.475 $Y=2.13
+ $X2=1.475 $Y2=1.79
r49 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=2.13
+ $X2=1.475 $Y2=2.295
r50 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.625
+ $X2=1.475 $Y2=1.79
r51 7 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.455 $Y=2.885
+ $X2=1.455 $Y2=2.295
r52 3 10 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.385 $Y=0.445
+ $X2=1.385 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_M%C1 1 3 6 8 11
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=0.93 $X2=2.015 $Y2=0.93
r34 11 13 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=1.925 $Y=0.93
+ $X2=2.015 $Y2=0.93
r35 8 14 9.18961 $w=1.73e-07 $l=1.45e-07 $layer=LI1_cond $X=2.16 $Y=0.927
+ $X2=2.015 $Y2=0.927
r36 4 11 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.095
+ $X2=1.925 $Y2=0.93
r37 4 6 917.851 $w=1.5e-07 $l=1.79e-06 $layer=POLY_cond $X=1.925 $Y=1.095
+ $X2=1.925 $Y2=2.885
r38 1 11 32.6165 $w=2.66e-07 $l=2.49199e-07 $layer=POLY_cond $X=1.745 $Y=0.765
+ $X2=1.925 $Y2=0.93
r39 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.745 $Y=0.765
+ $X2=1.745 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_M%VPWR 1 2 9 13 16 17 18 23 29 30 33
r37 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 30 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 27 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=1.69 $Y2=3.33
r41 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.69 $Y2=3.33
r43 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 18 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 18 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 16 21 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=0.285 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=3.33
+ $X2=0.45 $Y2=3.33
r50 15 25 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.45 $Y2=3.33
r52 11 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=3.245
+ $X2=1.69 $Y2=3.33
r53 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.69 $Y=3.245
+ $X2=1.69 $Y2=2.95
r54 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.45 $Y=3.245 $X2=0.45
+ $Y2=3.33
r55 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.45 $Y=3.245
+ $X2=0.45 $Y2=2.95
r56 2 13 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=2.675 $X2=1.69 $Y2=2.95
r57 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=2.675 $X2=0.45 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_M%Y 1 2 3 12 14 15 17 18 19 23 28 29 30 31 32
+ 54
c67 12 0 1.69038e-19 $X=1.24 $Y=2.82
r68 39 54 2.49696 $w=2.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.095 $Y=1.73
+ $X2=2.095 $Y2=1.665
r69 30 31 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.095 $Y=2.035
+ $X2=2.095 $Y2=2.405
r70 29 54 0.384148 $w=2.98e-07 $l=1e-08 $layer=LI1_cond $X=2.095 $Y=1.655
+ $X2=2.095 $Y2=1.665
r71 29 30 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.095 $Y=1.74
+ $X2=2.095 $Y2=2.035
r72 29 39 0.384148 $w=2.98e-07 $l=1e-08 $layer=LI1_cond $X=2.095 $Y=1.74
+ $X2=2.095 $Y2=1.73
r73 27 32 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=2.14 $Y=2.665
+ $X2=2.14 $Y2=2.775
r74 27 28 3.64284 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=2.14 $Y=2.665
+ $X2=2.095 $Y2=2.58
r75 26 31 3.45733 $w=2.98e-07 $l=9e-08 $layer=LI1_cond $X=2.095 $Y=2.495
+ $X2=2.095 $Y2=2.405
r76 26 28 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=2.495
+ $X2=2.095 $Y2=2.58
r77 25 29 11.7899 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.03 $Y=1.365
+ $X2=2.03 $Y2=1.58
r78 20 23 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.585 $Y=0.495
+ $X2=1.96 $Y2=0.495
r79 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.945 $Y=1.28
+ $X2=2.03 $Y2=1.365
r80 18 19 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.945 $Y=1.28
+ $X2=1.67 $Y2=1.28
r81 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.585 $Y=1.195
+ $X2=1.67 $Y2=1.28
r82 16 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0.66
+ $X2=1.585 $Y2=0.495
r83 16 17 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.585 $Y=0.66
+ $X2=1.585 $Y2=1.195
r84 14 28 2.83584 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.945 $Y=2.58
+ $X2=2.095 $Y2=2.58
r85 14 15 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.945 $Y=2.58
+ $X2=1.345 $Y2=2.58
r86 10 15 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.24 $Y=2.665
+ $X2=1.345 $Y2=2.58
r87 10 12 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.24 $Y=2.665
+ $X2=1.24 $Y2=2.82
r88 3 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.675 $X2=2.14 $Y2=2.82
r89 2 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=2.675 $X2=1.24 $Y2=2.82
r90 1 23 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.235 $X2=1.96 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_M%A_29_47# 1 2 9 11 12 15
c26 15 0 1.87164e-19 $X=1.17 $Y=0.51
c27 11 0 1.64738e-19 $X=1.065 $Y=0.75
r28 13 15 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.17 $Y=0.665
+ $X2=1.17 $Y2=0.51
r29 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.065 $Y=0.75
+ $X2=1.17 $Y2=0.665
r30 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.065 $Y=0.75
+ $X2=0.375 $Y2=0.75
r31 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.27 $Y=0.665
+ $X2=0.375 $Y2=0.75
r32 7 9 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.27 $Y=0.665
+ $X2=0.27 $Y2=0.51
r33 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.17 $Y2=0.51
r34 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_M%VGND 1 6 8 10 20 21 24
r33 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r36 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.72
+ $Y2=0
r37 15 17 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.2
+ $Y2=0
r38 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r39 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.72
+ $Y2=0
r41 10 12 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r42 8 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r43 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r44 8 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085 $X2=0.72
+ $Y2=0
r46 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.38
r47 1 6 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.72 $Y2=0.38
.ends

