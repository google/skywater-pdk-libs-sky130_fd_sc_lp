* File: sky130_fd_sc_lp__o41ai_1.spice
* Created: Wed Sep  2 10:28:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o41ai_1  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_A_156_49#_M1004_d N_B1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.2226 PD=1.22 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A4_M1003_g N_A_156_49#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.1596 PD=1.14 PS=1.22 NRD=2.856 NRS=7.14 M=1 R=5.6 SA=75000.7
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1006 N_A_156_49#_M1006_d N_A3_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1302 AS=0.126 PD=1.15 PS=1.14 NRD=0 NRS=0 M=1 R=5.6 SA=75001.2 SB=75001.2
+ A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_156_49#_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1722 AS=0.1302 PD=1.25 PS=1.15 NRD=8.568 NRS=4.284 M=1 R=5.6 SA=75001.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1001 N_A_156_49#_M1001_d N_A1_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1722 PD=2.21 PS=1.25 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.3528 PD=1.65 PS=3.08 NRD=12.4898 NRS=0.7683 M=1 R=8.4
+ SA=75000.2 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1008 A_264_367# N_A4_M1008_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.2457 PD=1.47 PS=1.65 NRD=7.8012 NRS=4.6886 M=1 R=8.4 SA=75000.7
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1009 A_336_367# N_A3_M1009_g A_264_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75001.1
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1002 A_444_367# N_A2_M1002_g A_336_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=21.8867 M=1 R=8.4 SA=75001.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g A_444_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75002.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o41ai_1.pxi.spice"
*
.ends
*
*
