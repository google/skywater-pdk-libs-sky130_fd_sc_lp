* NGSPICE file created from sky130_fd_sc_lp__ha_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__ha_lp A B VGND VNB VPB VPWR COUT SUM
M1000 a_296_286# B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=9.85e+11p ps=7.97e+06u
M1001 VGND A a_743_125# VNB nshort w=420000u l=150000u
+  ad=3.5385e+11p pd=4.21e+06u as=8.82e+10p ps=1.26e+06u
M1002 a_901_125# a_296_286# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 a_743_125# B a_296_286# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1004 VPWR a_83_153# SUM VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1005 a_369_47# a_296_286# a_83_153# VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=1.1865e+11p ps=1.41e+06u
M1006 VGND a_83_153# a_113_179# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 VPWR A a_493_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1008 a_113_179# a_83_153# SUM VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1009 VGND B a_369_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_493_419# B a_83_153# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=4.85e+11p ps=2.97e+06u
M1011 VPWR A a_296_286# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1012 COUT a_296_286# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1013 a_83_153# a_296_286# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1014 COUT a_296_286# a_901_125# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1015 a_369_47# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

