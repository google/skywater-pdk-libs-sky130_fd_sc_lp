* File: sky130_fd_sc_lp__einvp_2.pxi.spice
* Created: Fri Aug 28 10:33:51 2020
* 
x_PM_SKY130_FD_SC_LP__EINVP_2%TE N_TE_M1000_g N_TE_M1006_g N_TE_c_65_n
+ N_TE_c_73_n N_TE_c_66_n N_TE_M1004_g N_TE_c_67_n N_TE_c_68_n N_TE_c_69_n
+ N_TE_M1008_g N_TE_c_70_n N_TE_c_71_n TE N_TE_c_75_n N_TE_c_76_n
+ PM_SKY130_FD_SC_LP__EINVP_2%TE
x_PM_SKY130_FD_SC_LP__EINVP_2%A_30_131# N_A_30_131#_M1000_s N_A_30_131#_M1006_s
+ N_A_30_131#_c_131_n N_A_30_131#_M1003_g N_A_30_131#_c_132_n
+ N_A_30_131#_M1005_g N_A_30_131#_c_126_n N_A_30_131#_c_127_n
+ N_A_30_131#_c_128_n N_A_30_131#_c_129_n N_A_30_131#_c_130_n
+ PM_SKY130_FD_SC_LP__EINVP_2%A_30_131#
x_PM_SKY130_FD_SC_LP__EINVP_2%A N_A_c_174_n N_A_M1002_g N_A_M1001_g N_A_c_176_n
+ N_A_M1009_g N_A_M1007_g N_A_c_178_n A A N_A_c_180_n N_A_c_181_n
+ PM_SKY130_FD_SC_LP__EINVP_2%A
x_PM_SKY130_FD_SC_LP__EINVP_2%VPWR N_VPWR_M1006_d N_VPWR_M1003_d N_VPWR_c_217_n
+ N_VPWR_c_218_n N_VPWR_c_219_n N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n
+ VPWR N_VPWR_c_223_n N_VPWR_c_216_n N_VPWR_c_225_n
+ PM_SKY130_FD_SC_LP__EINVP_2%VPWR
x_PM_SKY130_FD_SC_LP__EINVP_2%A_249_367# N_A_249_367#_M1003_s
+ N_A_249_367#_M1005_s N_A_249_367#_M1007_s N_A_249_367#_c_277_n
+ N_A_249_367#_c_273_n N_A_249_367#_c_274_n N_A_249_367#_c_298_n
+ N_A_249_367#_c_285_n N_A_249_367#_c_275_n N_A_249_367#_c_276_n
+ PM_SKY130_FD_SC_LP__EINVP_2%A_249_367#
x_PM_SKY130_FD_SC_LP__EINVP_2%Z N_Z_M1002_s N_Z_M1001_d Z Z Z Z Z N_Z_c_308_n
+ PM_SKY130_FD_SC_LP__EINVP_2%Z
x_PM_SKY130_FD_SC_LP__EINVP_2%VGND N_VGND_M1000_d N_VGND_M1008_s N_VGND_c_325_n
+ N_VGND_c_326_n VGND N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n PM_SKY130_FD_SC_LP__EINVP_2%VGND
x_PM_SKY130_FD_SC_LP__EINVP_2%A_218_47# N_A_218_47#_M1004_d N_A_218_47#_M1002_d
+ N_A_218_47#_M1009_d N_A_218_47#_c_390_n N_A_218_47#_c_365_n
+ N_A_218_47#_c_366_n N_A_218_47#_c_367_n N_A_218_47#_c_368_n
+ N_A_218_47#_c_369_n N_A_218_47#_c_370_n PM_SKY130_FD_SC_LP__EINVP_2%A_218_47#
cc_1 VNB N_TE_M1000_g 0.0299077f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.865
cc_2 VNB N_TE_M1006_g 0.00865411f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.155
cc_3 VNB N_TE_c_65_n 0.0160043f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.41
cc_4 VNB N_TE_c_66_n 0.0191923f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.185
cc_5 VNB N_TE_c_67_n 0.00816314f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.78
cc_6 VNB N_TE_c_68_n 0.0268866f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.26
cc_7 VNB N_TE_c_69_n 0.0186908f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.185
cc_8 VNB N_TE_c_70_n 0.00630028f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.41
cc_9 VNB N_TE_c_71_n 0.0124883f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.26
cc_10 VNB N_A_30_131#_c_126_n 0.0321391f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_11 VNB N_A_30_131#_c_127_n 0.0030033f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=1.26
cc_12 VNB N_A_30_131#_c_128_n 0.0198688f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.41
cc_13 VNB N_A_30_131#_c_129_n 0.0411308f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.26
cc_14 VNB N_A_30_131#_c_130_n 0.00893146f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.69
cc_15 VNB N_A_c_174_n 0.0197818f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.335
cc_16 VNB N_A_M1001_g 0.0100859f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.78
cc_17 VNB N_A_c_176_n 0.0191005f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.41
cc_18 VNB N_A_M1007_g 0.00146273f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_19 VNB N_A_c_178_n 0.00715336f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.78
cc_20 VNB A 0.00724039f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.26
cc_21 VNB N_A_c_180_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.41
cc_22 VNB N_A_c_181_n 0.0555581f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.41
cc_23 VNB N_VPWR_c_216_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_325_n 0.0205283f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.41
cc_25 VNB N_VGND_c_326_n 0.00956531f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_26 VNB N_VGND_c_327_n 0.0183576f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=1.26
cc_27 VNB N_VGND_c_328_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.26
cc_28 VNB N_VGND_c_329_n 0.0395291f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.865
cc_29 VNB N_VGND_c_330_n 0.212345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_331_n 0.00740538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_332_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_218_47#_c_365_n 0.0190442f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_33 VNB N_A_218_47#_c_366_n 9.77998e-19 $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_34 VNB N_A_218_47#_c_367_n 0.0071775f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=1.26
cc_35 VNB N_A_218_47#_c_368_n 0.011971f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.185
cc_36 VNB N_A_218_47#_c_369_n 0.00385541f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=0.655
cc_37 VNB N_A_218_47#_c_370_n 0.023359f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.26
cc_38 VPB N_TE_M1006_g 0.0316725f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.155
cc_39 VPB N_TE_c_73_n 0.0203752f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=2.855
cc_40 VPB N_TE_c_67_n 0.0573676f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.78
cc_41 VPB N_TE_c_75_n 0.0277816f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.945
cc_42 VPB N_TE_c_76_n 0.0405639f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.945
cc_43 VPB N_A_30_131#_c_131_n 0.0187313f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.155
cc_44 VPB N_A_30_131#_c_132_n 0.0156087f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.41
cc_45 VPB N_A_30_131#_c_127_n 0.0370334f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=1.26
cc_46 VPB N_A_30_131#_c_129_n 0.00976757f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.26
cc_47 VPB N_A_M1001_g 0.0193857f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.78
cc_48 VPB N_A_M1007_g 0.0245703f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.655
cc_49 VPB A 0.00640005f $X=-0.19 $Y=1.655 $X2=1.37 $Y2=1.26
cc_50 VPB N_VPWR_c_217_n 0.0121789f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.155
cc_51 VPB N_VPWR_c_218_n 0.0142107f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.41
cc_52 VPB N_VPWR_c_219_n 4.00916e-19 $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.185
cc_53 VPB N_VPWR_c_220_n 0.011478f $X=-0.19 $Y=1.655 $X2=1.37 $Y2=1.26
cc_54 VPB N_VPWR_c_221_n 0.0252544f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=0.655
cc_55 VPB N_VPWR_c_222_n 0.00353254f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=0.655
cc_56 VPB N_VPWR_c_223_n 0.0346796f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.865
cc_57 VPB N_VPWR_c_216_n 0.0557295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_225_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_249_367#_c_273_n 0.00664288f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.485
cc_60 VPB N_A_249_367#_c_274_n 0.00221093f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.78
cc_61 VPB N_A_249_367#_c_275_n 0.00745909f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.26
cc_62 VPB N_A_249_367#_c_276_n 0.0372906f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.69
cc_63 N_TE_c_73_n N_A_30_131#_c_131_n 0.0121356f $X=0.94 $Y=2.855 $X2=0 $Y2=0
cc_64 N_TE_M1000_g N_A_30_131#_c_126_n 0.0143673f $X=0.49 $Y=0.865 $X2=0 $Y2=0
cc_65 N_TE_M1006_g N_A_30_131#_c_127_n 0.0103867f $X=0.49 $Y=2.155 $X2=0 $Y2=0
cc_66 N_TE_c_75_n N_A_30_131#_c_127_n 0.0240718f $X=0.575 $Y=2.945 $X2=0 $Y2=0
cc_67 N_TE_M1006_g N_A_30_131#_c_128_n 0.0106272f $X=0.49 $Y=2.155 $X2=0 $Y2=0
cc_68 N_TE_c_65_n N_A_30_131#_c_128_n 0.0112071f $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_69 N_TE_c_67_n N_A_30_131#_c_128_n 0.00636695f $X=1.015 $Y=2.78 $X2=0 $Y2=0
cc_70 N_TE_c_68_n N_A_30_131#_c_128_n 0.0115819f $X=1.37 $Y=1.26 $X2=0 $Y2=0
cc_71 N_TE_c_70_n N_A_30_131#_c_128_n 0.00805256f $X=0.49 $Y=1.41 $X2=0 $Y2=0
cc_72 N_TE_c_71_n N_A_30_131#_c_128_n 0.00869539f $X=1.015 $Y=1.26 $X2=0 $Y2=0
cc_73 N_TE_c_67_n N_A_30_131#_c_129_n 0.0121356f $X=1.015 $Y=2.78 $X2=0 $Y2=0
cc_74 N_TE_c_68_n N_A_30_131#_c_129_n 5.54078e-19 $X=1.37 $Y=1.26 $X2=0 $Y2=0
cc_75 N_TE_c_71_n N_A_30_131#_c_129_n 0.00378801f $X=1.015 $Y=1.26 $X2=0 $Y2=0
cc_76 N_TE_M1006_g N_VPWR_c_217_n 0.00308406f $X=0.49 $Y=2.155 $X2=0 $Y2=0
cc_77 N_TE_c_73_n N_VPWR_c_217_n 0.00942558f $X=0.94 $Y=2.855 $X2=0 $Y2=0
cc_78 N_TE_c_67_n N_VPWR_c_217_n 0.0067834f $X=1.015 $Y=2.78 $X2=0 $Y2=0
cc_79 N_TE_c_75_n N_VPWR_c_217_n 0.0317728f $X=0.575 $Y=2.945 $X2=0 $Y2=0
cc_80 N_TE_c_76_n N_VPWR_c_217_n 0.00246181f $X=0.74 $Y=2.945 $X2=0 $Y2=0
cc_81 N_TE_M1006_g N_VPWR_c_220_n 5.21352e-19 $X=0.49 $Y=2.155 $X2=0 $Y2=0
cc_82 N_TE_c_65_n N_VPWR_c_220_n 0.00117741f $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_83 N_TE_c_73_n N_VPWR_c_220_n 0.00394505f $X=0.94 $Y=2.855 $X2=0 $Y2=0
cc_84 N_TE_c_67_n N_VPWR_c_220_n 0.0249162f $X=1.015 $Y=2.78 $X2=0 $Y2=0
cc_85 N_TE_c_75_n N_VPWR_c_220_n 0.014747f $X=0.575 $Y=2.945 $X2=0 $Y2=0
cc_86 N_TE_c_76_n N_VPWR_c_220_n 5.03395e-19 $X=0.74 $Y=2.945 $X2=0 $Y2=0
cc_87 N_TE_c_73_n N_VPWR_c_221_n 0.00460599f $X=0.94 $Y=2.855 $X2=0 $Y2=0
cc_88 N_TE_c_75_n N_VPWR_c_221_n 0.0398431f $X=0.575 $Y=2.945 $X2=0 $Y2=0
cc_89 N_TE_c_76_n N_VPWR_c_221_n 0.00624407f $X=0.74 $Y=2.945 $X2=0 $Y2=0
cc_90 N_TE_c_73_n N_VPWR_c_216_n 0.00490874f $X=0.94 $Y=2.855 $X2=0 $Y2=0
cc_91 N_TE_c_75_n N_VPWR_c_216_n 0.0226965f $X=0.575 $Y=2.945 $X2=0 $Y2=0
cc_92 N_TE_c_76_n N_VPWR_c_216_n 0.00854368f $X=0.74 $Y=2.945 $X2=0 $Y2=0
cc_93 N_TE_c_67_n N_A_249_367#_c_277_n 0.0035558f $X=1.015 $Y=2.78 $X2=0 $Y2=0
cc_94 N_TE_c_67_n N_A_249_367#_c_274_n 0.00196579f $X=1.015 $Y=2.78 $X2=0 $Y2=0
cc_95 N_TE_M1000_g N_VGND_c_325_n 0.0171844f $X=0.49 $Y=0.865 $X2=0 $Y2=0
cc_96 N_TE_c_65_n N_VGND_c_325_n 0.00405635f $X=0.94 $Y=1.41 $X2=0 $Y2=0
cc_97 N_TE_c_66_n N_VGND_c_325_n 0.00671248f $X=1.015 $Y=1.185 $X2=0 $Y2=0
cc_98 N_TE_c_66_n N_VGND_c_326_n 6.47207e-19 $X=1.015 $Y=1.185 $X2=0 $Y2=0
cc_99 N_TE_c_69_n N_VGND_c_326_n 0.0127468f $X=1.445 $Y=1.185 $X2=0 $Y2=0
cc_100 N_TE_M1000_g N_VGND_c_327_n 0.00332367f $X=0.49 $Y=0.865 $X2=0 $Y2=0
cc_101 N_TE_c_66_n N_VGND_c_328_n 0.00585385f $X=1.015 $Y=1.185 $X2=0 $Y2=0
cc_102 N_TE_c_69_n N_VGND_c_328_n 0.00486043f $X=1.445 $Y=1.185 $X2=0 $Y2=0
cc_103 N_TE_M1000_g N_VGND_c_330_n 0.00387424f $X=0.49 $Y=0.865 $X2=0 $Y2=0
cc_104 N_TE_c_66_n N_VGND_c_330_n 0.0118358f $X=1.015 $Y=1.185 $X2=0 $Y2=0
cc_105 N_TE_c_69_n N_VGND_c_330_n 0.00824727f $X=1.445 $Y=1.185 $X2=0 $Y2=0
cc_106 N_TE_c_68_n N_A_218_47#_c_365_n 0.00371913f $X=1.37 $Y=1.26 $X2=0 $Y2=0
cc_107 N_TE_c_69_n N_A_218_47#_c_365_n 0.0114435f $X=1.445 $Y=1.185 $X2=0 $Y2=0
cc_108 N_TE_M1000_g N_A_218_47#_c_366_n 2.2014e-19 $X=0.49 $Y=0.865 $X2=0 $Y2=0
cc_109 N_TE_c_66_n N_A_218_47#_c_366_n 0.0027071f $X=1.015 $Y=1.185 $X2=0 $Y2=0
cc_110 N_TE_c_68_n N_A_218_47#_c_366_n 0.00638501f $X=1.37 $Y=1.26 $X2=0 $Y2=0
cc_111 N_TE_c_69_n N_A_218_47#_c_367_n 0.00374471f $X=1.445 $Y=1.185 $X2=0 $Y2=0
cc_112 N_A_30_131#_c_132_n N_A_M1001_g 0.0176224f $X=2.015 $Y=1.725 $X2=0 $Y2=0
cc_113 N_A_30_131#_c_128_n N_A_c_178_n 6.22636e-19 $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_114 N_A_30_131#_c_129_n N_A_c_178_n 0.0176224f $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_115 N_A_30_131#_c_131_n N_VPWR_c_218_n 0.00486043f $X=1.585 $Y=1.725 $X2=0
+ $Y2=0
cc_116 N_A_30_131#_c_131_n N_VPWR_c_219_n 0.0144311f $X=1.585 $Y=1.725 $X2=0
+ $Y2=0
cc_117 N_A_30_131#_c_132_n N_VPWR_c_219_n 0.0153101f $X=2.015 $Y=1.725 $X2=0
+ $Y2=0
cc_118 N_A_30_131#_c_131_n N_VPWR_c_220_n 0.003564f $X=1.585 $Y=1.725 $X2=0
+ $Y2=0
cc_119 N_A_30_131#_c_127_n N_VPWR_c_220_n 0.00153767f $X=0.275 $Y=1.98 $X2=0
+ $Y2=0
cc_120 N_A_30_131#_c_128_n N_VPWR_c_220_n 0.0344103f $X=1.925 $Y=1.51 $X2=0
+ $Y2=0
cc_121 N_A_30_131#_c_132_n N_VPWR_c_223_n 0.00486043f $X=2.015 $Y=1.725 $X2=0
+ $Y2=0
cc_122 N_A_30_131#_c_131_n N_VPWR_c_216_n 0.00954696f $X=1.585 $Y=1.725 $X2=0
+ $Y2=0
cc_123 N_A_30_131#_c_132_n N_VPWR_c_216_n 0.0082726f $X=2.015 $Y=1.725 $X2=0
+ $Y2=0
cc_124 N_A_30_131#_c_131_n N_A_249_367#_c_273_n 0.0129987f $X=1.585 $Y=1.725
+ $X2=0 $Y2=0
cc_125 N_A_30_131#_c_132_n N_A_249_367#_c_273_n 0.012831f $X=2.015 $Y=1.725
+ $X2=0 $Y2=0
cc_126 N_A_30_131#_c_128_n N_A_249_367#_c_273_n 0.0418287f $X=1.925 $Y=1.51
+ $X2=0 $Y2=0
cc_127 N_A_30_131#_c_129_n N_A_249_367#_c_273_n 0.00263139f $X=1.925 $Y=1.51
+ $X2=0 $Y2=0
cc_128 N_A_30_131#_c_128_n N_A_249_367#_c_274_n 0.0162207f $X=1.925 $Y=1.51
+ $X2=0 $Y2=0
cc_129 N_A_30_131#_c_128_n N_Z_c_308_n 0.00662334f $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A_30_131#_c_129_n N_Z_c_308_n 0.00159303f $X=1.925 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A_30_131#_c_126_n N_VGND_c_325_n 0.0167402f $X=0.275 $Y=0.885 $X2=0
+ $Y2=0
cc_132 N_A_30_131#_c_128_n N_VGND_c_325_n 0.0196654f $X=1.925 $Y=1.51 $X2=0
+ $Y2=0
cc_133 N_A_30_131#_c_126_n N_VGND_c_327_n 0.00412028f $X=0.275 $Y=0.885 $X2=0
+ $Y2=0
cc_134 N_A_30_131#_c_126_n N_VGND_c_330_n 0.00735187f $X=0.275 $Y=0.885 $X2=0
+ $Y2=0
cc_135 N_A_30_131#_c_128_n N_A_218_47#_c_365_n 0.0513656f $X=1.925 $Y=1.51 $X2=0
+ $Y2=0
cc_136 N_A_30_131#_c_129_n N_A_218_47#_c_365_n 0.0102883f $X=1.925 $Y=1.51 $X2=0
+ $Y2=0
cc_137 N_A_30_131#_c_128_n N_A_218_47#_c_366_n 0.0168892f $X=1.925 $Y=1.51 $X2=0
+ $Y2=0
cc_138 N_A_M1001_g N_VPWR_c_219_n 0.00109252f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_M1001_g N_VPWR_c_223_n 0.00357877f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_M1007_g N_VPWR_c_223_n 0.00357877f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_VPWR_c_216_n 0.00537654f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_M1007_g N_VPWR_c_216_n 0.00629314f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_M1001_g N_A_249_367#_c_273_n 4.90985e-19 $X=2.445 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_M1001_g N_A_249_367#_c_285_n 0.0115031f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1007_g N_A_249_367#_c_285_n 0.0114565f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_146 A N_A_249_367#_c_276_n 0.0228788f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A_c_181_n N_A_249_367#_c_276_n 0.00147549f $X=3.09 $Y=1.46 $X2=0 $Y2=0
cc_148 N_A_c_174_n N_Z_c_308_n 0.0109989f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_149 N_A_M1001_g N_Z_c_308_n 0.0228827f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_c_176_n N_Z_c_308_n 0.0146316f $X=2.875 $Y=1.295 $X2=0 $Y2=0
cc_151 N_A_M1007_g N_Z_c_308_n 0.0228514f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_c_178_n N_Z_c_308_n 0.00394947f $X=2.445 $Y=1.37 $X2=0 $Y2=0
cc_153 A N_Z_c_308_n 0.0405526f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A_c_180_n N_Z_c_308_n 0.00871516f $X=2.8 $Y=1.46 $X2=0 $Y2=0
cc_155 N_A_c_181_n N_Z_c_308_n 0.00754517f $X=3.09 $Y=1.46 $X2=0 $Y2=0
cc_156 N_A_c_174_n N_VGND_c_326_n 0.00119067f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_157 N_A_c_174_n N_VGND_c_329_n 0.0029147f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_158 N_A_c_176_n N_VGND_c_329_n 0.0029147f $X=2.875 $Y=1.295 $X2=0 $Y2=0
cc_159 N_A_c_174_n N_VGND_c_330_n 0.00428625f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_160 N_A_c_176_n N_VGND_c_330_n 0.00420369f $X=2.875 $Y=1.295 $X2=0 $Y2=0
cc_161 N_A_c_174_n N_A_218_47#_c_365_n 0.00116263f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_162 N_A_c_174_n N_A_218_47#_c_368_n 0.0128685f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_163 N_A_c_176_n N_A_218_47#_c_368_n 0.0128685f $X=2.875 $Y=1.295 $X2=0 $Y2=0
cc_164 A N_A_218_47#_c_370_n 0.0228786f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A_c_181_n N_A_218_47#_c_370_n 0.00161388f $X=3.09 $Y=1.46 $X2=0 $Y2=0
cc_166 N_VPWR_c_216_n N_A_249_367#_M1003_s 0.00444756f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_167 N_VPWR_c_216_n N_A_249_367#_M1005_s 0.00376627f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_216_n N_A_249_367#_M1007_s 0.00215161f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_218_n N_A_249_367#_c_277_n 0.0135387f $X=1.635 $Y=3.33 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_220_n N_A_249_367#_c_277_n 0.0886544f $X=0.705 $Y=1.99 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_216_n N_A_249_367#_c_277_n 0.00769778f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_172 N_VPWR_M1003_d N_A_249_367#_c_273_n 0.00176461f $X=1.66 $Y=1.835 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_219_n N_A_249_367#_c_273_n 0.0170777f $X=1.8 $Y=2.2 $X2=0 $Y2=0
cc_174 N_VPWR_c_220_n N_A_249_367#_c_274_n 0.0107846f $X=0.705 $Y=1.99 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_223_n N_A_249_367#_c_298_n 0.0125234f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_216_n N_A_249_367#_c_298_n 0.00738676f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_223_n N_A_249_367#_c_285_n 0.0361172f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_216_n N_A_249_367#_c_285_n 0.023676f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_223_n N_A_249_367#_c_275_n 0.017882f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_180 N_VPWR_c_216_n N_A_249_367#_c_275_n 0.0101029f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_216_n N_Z_M1001_d 0.00225186f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_182 N_A_249_367#_c_285_n N_Z_M1001_d 0.00332344f $X=2.995 $Y=2.99 $X2=0 $Y2=0
cc_183 N_A_249_367#_c_273_n N_Z_c_308_n 0.00915965f $X=2.135 $Y=1.86 $X2=0 $Y2=0
cc_184 N_A_249_367#_c_285_n N_Z_c_308_n 0.0159805f $X=2.995 $Y=2.99 $X2=0 $Y2=0
cc_185 N_A_249_367#_c_273_n N_A_218_47#_c_365_n 0.00963073f $X=2.135 $Y=1.86
+ $X2=0 $Y2=0
cc_186 N_Z_c_308_n N_A_218_47#_c_365_n 0.00869346f $X=2.66 $Y=0.68 $X2=0.24
+ $Y2=0.885
cc_187 N_Z_M1002_s N_A_218_47#_c_368_n 0.00176461f $X=2.52 $Y=0.345 $X2=0 $Y2=0
cc_188 N_Z_c_308_n N_A_218_47#_c_368_n 0.0159805f $X=2.66 $Y=0.68 $X2=0 $Y2=0
cc_189 N_VGND_c_330_n N_A_218_47#_M1004_d 0.00397496f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_190 N_VGND_c_328_n N_A_218_47#_c_390_n 0.0138717f $X=1.495 $Y=0 $X2=0 $Y2=0
cc_191 N_VGND_c_330_n N_A_218_47#_c_390_n 0.00886411f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_M1008_s N_A_218_47#_c_365_n 0.00225342f $X=1.52 $Y=0.235 $X2=0
+ $Y2=0
cc_193 N_VGND_c_326_n N_A_218_47#_c_365_n 0.0220026f $X=1.66 $Y=0.38 $X2=0 $Y2=0
cc_194 N_VGND_c_325_n N_A_218_47#_c_366_n 0.0034859f $X=0.8 $Y=0.38 $X2=0 $Y2=0
cc_195 N_VGND_c_326_n N_A_218_47#_c_367_n 0.0301918f $X=1.66 $Y=0.38 $X2=0 $Y2=0
cc_196 N_VGND_c_329_n N_A_218_47#_c_368_n 0.0608672f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_197 N_VGND_c_330_n N_A_218_47#_c_368_n 0.0339255f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_326_n N_A_218_47#_c_369_n 0.0118078f $X=1.66 $Y=0.38 $X2=0 $Y2=0
cc_199 N_VGND_c_329_n N_A_218_47#_c_369_n 0.0186386f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_c_330_n N_A_218_47#_c_369_n 0.0101082f $X=3.12 $Y=0 $X2=0 $Y2=0
