* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 X a_180_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND a_180_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR A1 a_878_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_37_49# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 X a_180_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR a_180_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 X a_180_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VGND a_180_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_575_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_180_23# a_37_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_878_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_180_23# A2 a_878_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_878_367# A2 a_180_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_575_65# a_37_49# a_180_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_180_23# a_37_49# a_575_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 X a_180_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_575_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VGND A1 a_575_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VPWR a_37_49# a_180_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_37_49# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR a_180_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND A2 a_575_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
