* File: sky130_fd_sc_lp__nand2b_4.pxi.spice
* Created: Wed Sep  2 10:03:40 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2B_4%A_N N_A_N_M1011_g N_A_N_M1016_g A_N N_A_N_c_90_n
+ N_A_N_c_91_n PM_SKY130_FD_SC_LP__NAND2B_4%A_N
x_PM_SKY130_FD_SC_LP__NAND2B_4%A_27_51# N_A_27_51#_M1011_s N_A_27_51#_M1016_s
+ N_A_27_51#_M1002_g N_A_27_51#_M1000_g N_A_27_51#_M1006_g N_A_27_51#_M1001_g
+ N_A_27_51#_M1007_g N_A_27_51#_M1008_g N_A_27_51#_M1012_g N_A_27_51#_M1015_g
+ N_A_27_51#_c_125_n N_A_27_51#_c_137_n N_A_27_51#_c_138_n N_A_27_51#_c_126_n
+ N_A_27_51#_c_127_n N_A_27_51#_c_150_n N_A_27_51#_c_128_n N_A_27_51#_c_129_n
+ N_A_27_51#_c_169_p N_A_27_51#_c_130_n N_A_27_51#_c_131_n N_A_27_51#_c_132_n
+ PM_SKY130_FD_SC_LP__NAND2B_4%A_27_51#
x_PM_SKY130_FD_SC_LP__NAND2B_4%B N_B_M1003_g N_B_M1004_g N_B_M1005_g N_B_M1009_g
+ N_B_M1010_g N_B_M1013_g N_B_M1014_g N_B_M1017_g B B B N_B_c_255_n
+ PM_SKY130_FD_SC_LP__NAND2B_4%B
x_PM_SKY130_FD_SC_LP__NAND2B_4%VPWR N_VPWR_M1016_d N_VPWR_M1006_d N_VPWR_M1012_d
+ N_VPWR_M1009_d N_VPWR_M1017_d N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n
+ N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_344_n
+ N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n
+ N_VPWR_c_337_n VPWR N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n
+ N_VPWR_c_324_n PM_SKY130_FD_SC_LP__NAND2B_4%VPWR
x_PM_SKY130_FD_SC_LP__NAND2B_4%Y N_Y_M1000_d N_Y_M1008_d N_Y_M1002_s N_Y_M1007_s
+ N_Y_M1004_s N_Y_M1013_s N_Y_c_468_n N_Y_c_416_n N_Y_c_413_n N_Y_c_414_n
+ N_Y_c_408_n N_Y_c_409_n N_Y_c_437_n N_Y_c_410_n N_Y_c_451_n N_Y_c_455_n
+ N_Y_c_475_n N_Y_c_411_n Y Y Y N_Y_c_459_n N_Y_c_412_n Y N_Y_c_448_n
+ N_Y_c_483_n PM_SKY130_FD_SC_LP__NAND2B_4%Y
x_PM_SKY130_FD_SC_LP__NAND2B_4%VGND N_VGND_M1011_d N_VGND_M1003_d N_VGND_M1010_d
+ N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ N_VGND_c_503_n N_VGND_c_504_n VGND N_VGND_c_505_n N_VGND_c_506_n
+ N_VGND_c_507_n N_VGND_c_508_n PM_SKY130_FD_SC_LP__NAND2B_4%VGND
x_PM_SKY130_FD_SC_LP__NAND2B_4%A_217_65# N_A_217_65#_M1000_s N_A_217_65#_M1001_s
+ N_A_217_65#_M1015_s N_A_217_65#_M1005_s N_A_217_65#_M1014_s
+ N_A_217_65#_c_564_n N_A_217_65#_c_565_n N_A_217_65#_c_566_n
+ N_A_217_65#_c_582_n N_A_217_65#_c_567_n N_A_217_65#_c_568_n
+ N_A_217_65#_c_569_n N_A_217_65#_c_570_n N_A_217_65#_c_571_n
+ N_A_217_65#_c_572_n N_A_217_65#_c_573_n N_A_217_65#_c_574_n
+ PM_SKY130_FD_SC_LP__NAND2B_4%A_217_65#
cc_1 VNB N_A_N_M1011_g 0.0308454f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.675
cc_2 VNB N_A_N_M1016_g 0.00176153f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A_N_c_90_n 0.0425999f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_4 VNB N_A_N_c_91_n 0.010931f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_5 VNB N_A_27_51#_M1000_g 0.0234147f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_6 VNB N_A_27_51#_M1001_g 0.0198126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_51#_M1008_g 0.0206139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_51#_M1015_g 0.0201527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_51#_c_125_n 0.0306079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_51#_c_126_n 0.00613023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_51#_c_127_n 0.0110866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_51#_c_128_n 0.00379243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_51#_c_129_n 3.46832e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_51#_c_130_n 0.00102142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_51#_c_131_n 0.0377509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_51#_c_132_n 0.0738125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_M1003_g 0.0193682f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.675
cc_18 VNB N_B_M1005_g 0.0190876f $X=-0.19 $Y=-0.245 $X2=0.357 $Y2=1.46
cc_19 VNB N_B_M1010_g 0.0190876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_M1014_g 0.0259905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB B 0.0183748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_255_n 0.0881543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_324_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_408_n 0.00313495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_409_n 0.00228483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_410_n 8.75342e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_411_n 0.00131115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_412_n 0.00413361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_498_n 0.00916177f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_30 VNB N_VGND_c_499_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.46
cc_31 VNB N_VGND_c_500_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_501_n 0.0578927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_502_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_503_n 0.0142255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_504_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_505_n 0.0156016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_506_n 0.0235135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_507_n 0.310496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_508_n 0.00528596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_217_65#_c_564_n 0.00983413f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.665
cc_41 VNB N_A_217_65#_c_565_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_217_65#_c_566_n 0.0036506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_217_65#_c_567_n 0.00471508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_217_65#_c_568_n 0.003383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_217_65#_c_569_n 0.00316221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_217_65#_c_570_n 0.00214825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_217_65#_c_571_n 0.0123411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_217_65#_c_572_n 0.0312591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_217_65#_c_573_n 0.00221189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_217_65#_c_574_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_A_N_M1016_g 0.0289984f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_52 VPB N_A_N_c_91_n 0.00619398f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.46
cc_53 VPB N_A_27_51#_M1002_g 0.0224353f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_54 VPB N_A_27_51#_M1006_g 0.0190161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_27_51#_M1007_g 0.0189837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_27_51#_M1012_g 0.0188369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_27_51#_c_137_n 0.00880428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_27_51#_c_138_n 0.0369431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_27_51#_c_129_n 0.00303354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_27_51#_c_131_n 0.0153175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_27_51#_c_132_n 0.0170768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_B_M1004_g 0.0207094f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_63 VPB N_B_M1009_g 0.0187318f $X=-0.19 $Y=1.655 $X2=0.357 $Y2=1.625
cc_64 VPB N_B_M1013_g 0.0180542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B_M1017_g 0.0233606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB B 0.0231017f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_B_c_255_n 0.021496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_325_n 0.00448275f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_326_n 0.00241491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_327_n 0.00444312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_328_n 0.00501089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_329_n 0.00459242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_330_n 0.0157625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_331_n 0.0479818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_332_n 0.0165512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_333_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_334_n 0.0173748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_335_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_336_n 0.0189541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_337_n 0.00507132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_338_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_339_n 0.0146078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_340_n 0.0129947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_324_n 0.0513786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_Y_c_413_n 0.00270367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_Y_c_414_n 0.00281685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_Y_c_412_n 0.00494997f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 N_A_N_M1016_g N_A_27_51#_M1002_g 0.00604141f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_N_c_90_n N_A_27_51#_c_137_n 0.00105438f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_90 N_A_N_c_91_n N_A_27_51#_c_137_n 0.0170218f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_91 N_A_N_M1011_g N_A_27_51#_c_126_n 0.0173038f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_92 N_A_N_c_90_n N_A_27_51#_c_126_n 0.00133621f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_93 N_A_N_c_91_n N_A_27_51#_c_126_n 0.0110197f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_94 N_A_N_c_90_n N_A_27_51#_c_127_n 0.00456171f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_95 N_A_N_c_91_n N_A_27_51#_c_127_n 0.0162521f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_96 N_A_N_M1016_g N_A_27_51#_c_150_n 0.0147913f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_N_c_91_n N_A_27_51#_c_150_n 0.00874699f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_98 N_A_N_M1011_g N_A_27_51#_c_128_n 0.00642795f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_99 N_A_N_c_91_n N_A_27_51#_c_128_n 0.00448175f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_100 N_A_N_c_90_n N_A_27_51#_c_129_n 0.00582009f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_101 N_A_N_c_91_n N_A_27_51#_c_129_n 0.012353f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_102 N_A_N_c_90_n N_A_27_51#_c_130_n 0.00118572f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_103 N_A_N_c_91_n N_A_27_51#_c_130_n 0.0143649f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_104 N_A_N_c_90_n N_A_27_51#_c_131_n 0.0205717f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_105 N_A_N_c_91_n N_A_27_51#_c_131_n 2.94943e-19 $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_106 N_A_N_M1016_g N_VPWR_c_325_n 0.0136363f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_N_M1016_g N_VPWR_c_326_n 0.00164531f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_N_M1016_g N_VPWR_c_344_n 0.00616409f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_N_M1016_g N_VPWR_c_338_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_N_M1016_g N_VPWR_c_324_n 0.00917987f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_N_M1011_g N_VGND_c_498_n 0.01295f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_112 N_A_N_M1011_g N_VGND_c_505_n 0.00469214f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_113 N_A_N_M1011_g N_VGND_c_507_n 0.0091141f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_114 N_A_N_M1011_g N_A_217_65#_c_564_n 0.00367486f $X=0.475 $Y=0.675 $X2=0
+ $Y2=0
cc_115 N_A_27_51#_M1015_g N_B_M1003_g 0.0182358f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_116 N_A_27_51#_M1012_g N_B_M1004_g 0.0343938f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_27_51#_c_132_n B 2.75645e-19 $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A_27_51#_c_132_n N_B_c_255_n 0.0182358f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_119 N_A_27_51#_c_150_n N_VPWR_M1016_d 0.00726746f $X=0.665 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_27_51#_c_129_n N_VPWR_M1016_d 0.00235298f $X=0.75 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_27_51#_M1002_g N_VPWR_c_326_n 0.00491485f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_27_51#_c_150_n N_VPWR_c_326_n 0.0142383f $X=0.665 $Y=2.015 $X2=0
+ $Y2=0
cc_123 N_A_27_51#_c_129_n N_VPWR_c_326_n 0.00981374f $X=0.75 $Y=1.93 $X2=0 $Y2=0
cc_124 N_A_27_51#_c_169_p N_VPWR_c_326_n 0.0180951f $X=2.285 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A_27_51#_c_131_n N_VPWR_c_326_n 0.00650808f $X=1.27 $Y=1.51 $X2=0 $Y2=0
cc_126 N_A_27_51#_M1006_g N_VPWR_c_327_n 0.00177178f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_A_27_51#_M1007_g N_VPWR_c_327_n 0.00182632f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_A_27_51#_M1012_g N_VPWR_c_328_n 0.00665091f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_27_51#_c_132_n N_VPWR_c_328_n 2.86496e-19 $X=2.855 $Y=1.51 $X2=0
+ $Y2=0
cc_130 N_A_27_51#_c_150_n N_VPWR_c_344_n 0.0217057f $X=0.665 $Y=2.015 $X2=0
+ $Y2=0
cc_131 N_A_27_51#_c_169_p N_VPWR_c_344_n 0.00449833f $X=2.285 $Y=1.51 $X2=0
+ $Y2=0
cc_132 N_A_27_51#_c_131_n N_VPWR_c_344_n 0.0033047f $X=1.27 $Y=1.51 $X2=0 $Y2=0
cc_133 N_A_27_51#_M1002_g N_VPWR_c_332_n 0.00585385f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_27_51#_M1006_g N_VPWR_c_332_n 0.00585385f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_27_51#_M1007_g N_VPWR_c_334_n 0.00585385f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_27_51#_M1012_g N_VPWR_c_334_n 0.0054895f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_27_51#_c_138_n N_VPWR_c_338_n 0.0178111f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_138 N_A_27_51#_M1016_s N_VPWR_c_324_n 0.00371702f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_139 N_A_27_51#_M1002_g N_VPWR_c_324_n 0.0112694f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_27_51#_M1006_g N_VPWR_c_324_n 0.0107298f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A_27_51#_M1007_g N_VPWR_c_324_n 0.0107298f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_27_51#_M1012_g N_VPWR_c_324_n 0.0102236f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_27_51#_c_138_n N_VPWR_c_324_n 0.0100304f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_144 N_A_27_51#_M1000_g N_Y_c_416_n 0.00544024f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_145 N_A_27_51#_M1001_g N_Y_c_416_n 0.00688101f $X=1.855 $Y=0.745 $X2=0 $Y2=0
cc_146 N_A_27_51#_M1008_g N_Y_c_416_n 2.75259e-19 $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_147 N_A_27_51#_M1006_g N_Y_c_413_n 0.0141248f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_27_51#_M1007_g N_Y_c_413_n 0.0142694f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_27_51#_c_169_p N_Y_c_413_n 0.0467246f $X=2.285 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A_27_51#_c_132_n N_Y_c_413_n 0.00478035f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A_27_51#_M1002_g N_Y_c_414_n 8.92873e-19 $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_27_51#_c_129_n N_Y_c_414_n 0.00121342f $X=0.75 $Y=1.93 $X2=0 $Y2=0
cc_153 N_A_27_51#_c_169_p N_Y_c_414_n 0.02098f $X=2.285 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A_27_51#_c_132_n N_Y_c_414_n 0.00291181f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A_27_51#_M1001_g N_Y_c_408_n 0.00961273f $X=1.855 $Y=0.745 $X2=0 $Y2=0
cc_156 N_A_27_51#_M1008_g N_Y_c_408_n 0.013136f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_157 N_A_27_51#_c_169_p N_Y_c_408_n 0.0450717f $X=2.285 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A_27_51#_c_132_n N_Y_c_408_n 0.00449089f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A_27_51#_M1000_g N_Y_c_409_n 0.00401488f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_160 N_A_27_51#_M1001_g N_Y_c_409_n 0.00180291f $X=1.855 $Y=0.745 $X2=0 $Y2=0
cc_161 N_A_27_51#_c_126_n N_Y_c_409_n 3.23963e-19 $X=0.665 $Y=1.11 $X2=0 $Y2=0
cc_162 N_A_27_51#_c_128_n N_Y_c_409_n 0.0017168f $X=0.75 $Y=1.425 $X2=0 $Y2=0
cc_163 N_A_27_51#_c_169_p N_Y_c_409_n 0.0263008f $X=2.285 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A_27_51#_c_132_n N_Y_c_409_n 0.00290354f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A_27_51#_M1015_g N_Y_c_437_n 0.00517847f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_166 N_A_27_51#_M1008_g N_Y_c_410_n 0.00188828f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_167 N_A_27_51#_M1015_g N_Y_c_410_n 0.00232961f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_168 N_A_27_51#_c_169_p N_Y_c_410_n 0.0010382f $X=2.285 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A_27_51#_c_132_n N_Y_c_410_n 0.00854843f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A_27_51#_M1015_g N_Y_c_411_n 0.00298575f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_171 N_A_27_51#_c_132_n N_Y_c_411_n 0.00342061f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A_27_51#_M1007_g N_Y_c_412_n 0.00203563f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A_27_51#_M1012_g N_Y_c_412_n 0.0202016f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_27_51#_c_169_p N_Y_c_412_n 0.0195197f $X=2.285 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A_27_51#_c_132_n N_Y_c_412_n 0.0278243f $X=2.855 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A_27_51#_M1012_g N_Y_c_448_n 0.0133604f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A_27_51#_c_126_n N_VGND_M1011_d 0.00259519f $X=0.665 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_27_51#_M1000_g N_VGND_c_498_n 0.00149641f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_179 N_A_27_51#_c_126_n N_VGND_c_498_n 0.0218666f $X=0.665 $Y=1.11 $X2=0 $Y2=0
cc_180 N_A_27_51#_c_169_p N_VGND_c_498_n 6.06678e-19 $X=2.285 $Y=1.51 $X2=0
+ $Y2=0
cc_181 N_A_27_51#_c_131_n N_VGND_c_498_n 6.82252e-19 $X=1.27 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_27_51#_M1015_g N_VGND_c_499_n 5.15399e-19 $X=2.855 $Y=0.745 $X2=0
+ $Y2=0
cc_183 N_A_27_51#_M1000_g N_VGND_c_501_n 0.00302501f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_184 N_A_27_51#_M1001_g N_VGND_c_501_n 0.00302501f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_185 N_A_27_51#_M1008_g N_VGND_c_501_n 0.00302473f $X=2.355 $Y=0.745 $X2=0
+ $Y2=0
cc_186 N_A_27_51#_M1015_g N_VGND_c_501_n 0.00302501f $X=2.855 $Y=0.745 $X2=0
+ $Y2=0
cc_187 N_A_27_51#_c_125_n N_VGND_c_505_n 0.0174563f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_188 N_A_27_51#_M1000_g N_VGND_c_507_n 0.0048466f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_189 N_A_27_51#_M1001_g N_VGND_c_507_n 0.00441253f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_190 N_A_27_51#_M1008_g N_VGND_c_507_n 0.00447833f $X=2.355 $Y=0.745 $X2=0
+ $Y2=0
cc_191 N_A_27_51#_M1015_g N_VGND_c_507_n 0.00442227f $X=2.855 $Y=0.745 $X2=0
+ $Y2=0
cc_192 N_A_27_51#_c_125_n N_VGND_c_507_n 0.00963638f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_193 N_A_27_51#_M1000_g N_A_217_65#_c_564_n 0.00354524f $X=1.425 $Y=0.745
+ $X2=0 $Y2=0
cc_194 N_A_27_51#_c_126_n N_A_217_65#_c_564_n 0.0119909f $X=0.665 $Y=1.11 $X2=0
+ $Y2=0
cc_195 N_A_27_51#_c_169_p N_A_217_65#_c_564_n 0.0160751f $X=2.285 $Y=1.51 $X2=0
+ $Y2=0
cc_196 N_A_27_51#_c_131_n N_A_217_65#_c_564_n 0.00649619f $X=1.27 $Y=1.51 $X2=0
+ $Y2=0
cc_197 N_A_27_51#_M1000_g N_A_217_65#_c_565_n 0.012559f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_198 N_A_27_51#_M1001_g N_A_217_65#_c_565_n 0.0116483f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_199 N_A_27_51#_M1008_g N_A_217_65#_c_582_n 0.00707611f $X=2.355 $Y=0.745
+ $X2=0 $Y2=0
cc_200 N_A_27_51#_M1015_g N_A_217_65#_c_582_n 3.06659e-19 $X=2.855 $Y=0.745
+ $X2=0 $Y2=0
cc_201 N_A_27_51#_M1008_g N_A_217_65#_c_567_n 0.00869988f $X=2.355 $Y=0.745
+ $X2=0 $Y2=0
cc_202 N_A_27_51#_M1015_g N_A_217_65#_c_567_n 0.0122087f $X=2.855 $Y=0.745 $X2=0
+ $Y2=0
cc_203 N_A_27_51#_M1015_g N_A_217_65#_c_569_n 7.3655e-19 $X=2.855 $Y=0.745 $X2=0
+ $Y2=0
cc_204 N_A_27_51#_M1008_g N_A_217_65#_c_573_n 0.00152703f $X=2.355 $Y=0.745
+ $X2=0 $Y2=0
cc_205 N_B_M1004_g N_VPWR_c_328_n 0.0080481f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B_M1009_g N_VPWR_c_329_n 0.00368151f $X=3.775 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B_M1013_g N_VPWR_c_329_n 0.00218677f $X=4.205 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B_M1013_g N_VPWR_c_331_n 7.38245e-19 $X=4.205 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B_M1017_g N_VPWR_c_331_n 0.020143f $X=4.635 $Y=2.465 $X2=0 $Y2=0
cc_210 B N_VPWR_c_331_n 0.0257694f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_211 N_B_c_255_n N_VPWR_c_331_n 0.00132005f $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_212 N_B_M1004_g N_VPWR_c_336_n 0.00585385f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B_M1009_g N_VPWR_c_336_n 0.00585385f $X=3.775 $Y=2.465 $X2=0 $Y2=0
cc_214 N_B_M1013_g N_VPWR_c_339_n 0.00585385f $X=4.205 $Y=2.465 $X2=0 $Y2=0
cc_215 N_B_M1017_g N_VPWR_c_339_n 0.00486043f $X=4.635 $Y=2.465 $X2=0 $Y2=0
cc_216 N_B_M1004_g N_VPWR_c_324_n 0.0112241f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_217 N_B_M1009_g N_VPWR_c_324_n 0.0106705f $X=3.775 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B_M1013_g N_VPWR_c_324_n 0.0105087f $X=4.205 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B_M1017_g N_VPWR_c_324_n 0.00824727f $X=4.635 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B_M1003_g N_Y_c_410_n 9.60448e-19 $X=3.285 $Y=0.745 $X2=0 $Y2=0
cc_221 B N_Y_c_410_n 4.74855e-19 $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B_M1009_g N_Y_c_451_n 0.0129469f $X=3.775 $Y=2.465 $X2=0 $Y2=0
cc_223 N_B_M1013_g N_Y_c_451_n 0.0129934f $X=4.205 $Y=2.465 $X2=0 $Y2=0
cc_224 B N_Y_c_451_n 0.040138f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B_c_255_n N_Y_c_451_n 5.60268e-19 $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_226 B N_Y_c_455_n 0.0166692f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B_c_255_n N_Y_c_455_n 6.3349e-19 $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_228 B Y 0.0239715f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_229 N_B_c_255_n Y 0.00101623f $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_230 N_B_M1004_g N_Y_c_459_n 0.0149492f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_231 B N_Y_c_459_n 0.00789478f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_232 B N_Y_c_412_n 0.0275439f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B_c_255_n N_Y_c_412_n 0.00777515f $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_234 N_B_M1004_g N_Y_c_448_n 9.3101e-19 $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_235 N_B_M1003_g N_VGND_c_499_n 0.0102666f $X=3.285 $Y=0.745 $X2=0 $Y2=0
cc_236 N_B_M1005_g N_VGND_c_499_n 0.0100754f $X=3.715 $Y=0.745 $X2=0 $Y2=0
cc_237 N_B_M1010_g N_VGND_c_499_n 4.59082e-19 $X=4.145 $Y=0.745 $X2=0 $Y2=0
cc_238 N_B_M1005_g N_VGND_c_500_n 4.56253e-19 $X=3.715 $Y=0.745 $X2=0 $Y2=0
cc_239 N_B_M1010_g N_VGND_c_500_n 0.00997431f $X=4.145 $Y=0.745 $X2=0 $Y2=0
cc_240 N_B_M1014_g N_VGND_c_500_n 0.0124264f $X=4.575 $Y=0.745 $X2=0 $Y2=0
cc_241 N_B_M1003_g N_VGND_c_501_n 0.00414769f $X=3.285 $Y=0.745 $X2=0 $Y2=0
cc_242 N_B_M1005_g N_VGND_c_503_n 0.00414769f $X=3.715 $Y=0.745 $X2=0 $Y2=0
cc_243 N_B_M1010_g N_VGND_c_503_n 0.00414769f $X=4.145 $Y=0.745 $X2=0 $Y2=0
cc_244 N_B_M1014_g N_VGND_c_506_n 0.00414769f $X=4.575 $Y=0.745 $X2=0 $Y2=0
cc_245 N_B_M1003_g N_VGND_c_507_n 0.0078848f $X=3.285 $Y=0.745 $X2=0 $Y2=0
cc_246 N_B_M1005_g N_VGND_c_507_n 0.00787505f $X=3.715 $Y=0.745 $X2=0 $Y2=0
cc_247 N_B_M1010_g N_VGND_c_507_n 0.00787505f $X=4.145 $Y=0.745 $X2=0 $Y2=0
cc_248 N_B_M1014_g N_VGND_c_507_n 0.00829411f $X=4.575 $Y=0.745 $X2=0 $Y2=0
cc_249 N_B_M1003_g N_A_217_65#_c_567_n 5.73473e-19 $X=3.285 $Y=0.745 $X2=0 $Y2=0
cc_250 N_B_M1003_g N_A_217_65#_c_568_n 0.013709f $X=3.285 $Y=0.745 $X2=0 $Y2=0
cc_251 N_B_M1005_g N_A_217_65#_c_568_n 0.013286f $X=3.715 $Y=0.745 $X2=0 $Y2=0
cc_252 B N_A_217_65#_c_568_n 0.043009f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_253 N_B_c_255_n N_A_217_65#_c_568_n 0.00246472f $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_254 N_B_M1005_g N_A_217_65#_c_570_n 0.00105889f $X=3.715 $Y=0.745 $X2=0 $Y2=0
cc_255 N_B_M1010_g N_A_217_65#_c_570_n 0.00105889f $X=4.145 $Y=0.745 $X2=0 $Y2=0
cc_256 N_B_M1010_g N_A_217_65#_c_571_n 0.0136351f $X=4.145 $Y=0.745 $X2=0 $Y2=0
cc_257 N_B_M1014_g N_A_217_65#_c_571_n 0.0143594f $X=4.575 $Y=0.745 $X2=0 $Y2=0
cc_258 B N_A_217_65#_c_571_n 0.0714367f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_259 N_B_c_255_n N_A_217_65#_c_571_n 0.0103826f $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_260 N_B_M1014_g N_A_217_65#_c_572_n 0.00354556f $X=4.575 $Y=0.745 $X2=0 $Y2=0
cc_261 B N_A_217_65#_c_574_n 0.0160407f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_262 N_B_c_255_n N_A_217_65#_c_574_n 0.00282576f $X=4.775 $Y=1.51 $X2=0 $Y2=0
cc_263 N_VPWR_c_324_n N_Y_M1002_s 0.00293134f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_264 N_VPWR_c_324_n N_Y_M1007_s 0.00240953f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_c_324_n N_Y_M1004_s 0.00306597f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_266 N_VPWR_c_324_n N_Y_M1013_s 0.00432284f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_332_n N_Y_c_468_n 0.0149362f $X=1.865 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_c_324_n N_Y_c_468_n 0.0100304f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_M1006_d N_Y_c_413_n 0.00261503f $X=1.85 $Y=1.835 $X2=0 $Y2=0
cc_270 N_VPWR_c_327_n N_Y_c_413_n 0.0200142f $X=2.03 $Y=2.19 $X2=0 $Y2=0
cc_271 N_VPWR_c_326_n N_Y_c_414_n 0.00295513f $X=1.13 $Y=1.965 $X2=0 $Y2=0
cc_272 N_VPWR_M1009_d N_Y_c_451_n 0.00333177f $X=3.85 $Y=1.835 $X2=0 $Y2=0
cc_273 N_VPWR_c_329_n N_Y_c_451_n 0.0135055f $X=3.99 $Y=2.435 $X2=0 $Y2=0
cc_274 N_VPWR_c_339_n N_Y_c_475_n 0.0135169f $X=4.685 $Y=3.33 $X2=0 $Y2=0
cc_275 N_VPWR_c_324_n N_Y_c_475_n 0.00847534f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_276 N_VPWR_M1012_d N_Y_c_459_n 0.00229844f $X=2.79 $Y=1.835 $X2=0 $Y2=0
cc_277 N_VPWR_c_328_n N_Y_c_459_n 0.00594688f $X=3 $Y=2.375 $X2=0 $Y2=0
cc_278 N_VPWR_M1012_d N_Y_c_412_n 0.0047294f $X=2.79 $Y=1.835 $X2=0 $Y2=0
cc_279 N_VPWR_c_328_n N_Y_c_412_n 0.0210077f $X=3 $Y=2.375 $X2=0 $Y2=0
cc_280 N_VPWR_c_334_n N_Y_c_448_n 0.0171073f $X=2.835 $Y=3.33 $X2=0 $Y2=0
cc_281 N_VPWR_c_324_n N_Y_c_448_n 0.0114026f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_282 N_VPWR_c_336_n N_Y_c_483_n 0.0195097f $X=3.86 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_324_n N_Y_c_483_n 0.0127519f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_284 N_Y_c_408_n N_A_217_65#_M1001_s 0.00250873f $X=2.475 $Y=1.17 $X2=0 $Y2=0
cc_285 N_Y_c_409_n N_A_217_65#_c_564_n 0.00497809f $X=1.805 $Y=1.17 $X2=0 $Y2=0
cc_286 N_Y_M1000_d N_A_217_65#_c_565_n 0.00180746f $X=1.5 $Y=0.325 $X2=0 $Y2=0
cc_287 N_Y_c_416_n N_A_217_65#_c_565_n 0.015151f $X=1.64 $Y=0.69 $X2=0 $Y2=0
cc_288 N_Y_c_408_n N_A_217_65#_c_565_n 0.00272017f $X=2.475 $Y=1.17 $X2=0 $Y2=0
cc_289 N_Y_c_408_n N_A_217_65#_c_582_n 0.0209355f $X=2.475 $Y=1.17 $X2=0 $Y2=0
cc_290 N_Y_M1008_d N_A_217_65#_c_567_n 0.00256964f $X=2.43 $Y=0.325 $X2=0 $Y2=0
cc_291 N_Y_c_408_n N_A_217_65#_c_567_n 0.00272017f $X=2.475 $Y=1.17 $X2=0 $Y2=0
cc_292 N_Y_c_437_n N_A_217_65#_c_567_n 0.0186552f $X=2.64 $Y=0.69 $X2=0 $Y2=0
cc_293 N_Y_c_459_n N_A_217_65#_c_568_n 0.00149485f $X=3.36 $Y=2.025 $X2=0 $Y2=0
cc_294 N_Y_c_411_n N_A_217_65#_c_569_n 0.011362f $X=2.64 $Y=1.17 $X2=0 $Y2=0
cc_295 N_Y_c_459_n N_A_217_65#_c_569_n 0.00244995f $X=3.36 $Y=2.025 $X2=0 $Y2=0
cc_296 N_Y_c_412_n N_A_217_65#_c_569_n 0.00926285f $X=3.08 $Y=2.025 $X2=0 $Y2=0
cc_297 N_VGND_c_498_n N_A_217_65#_c_564_n 0.032487f $X=0.69 $Y=0.4 $X2=0 $Y2=0
cc_298 N_VGND_c_501_n N_A_217_65#_c_565_n 0.0422287f $X=3.335 $Y=0 $X2=0 $Y2=0
cc_299 N_VGND_c_507_n N_A_217_65#_c_565_n 0.0238173f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_300 N_VGND_c_498_n N_A_217_65#_c_566_n 0.0139f $X=0.69 $Y=0.4 $X2=0 $Y2=0
cc_301 N_VGND_c_501_n N_A_217_65#_c_566_n 0.0186386f $X=3.335 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_507_n N_A_217_65#_c_566_n 0.0101082f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_303 N_VGND_c_499_n N_A_217_65#_c_567_n 0.00962585f $X=3.5 $Y=0.45 $X2=0 $Y2=0
cc_304 N_VGND_c_501_n N_A_217_65#_c_567_n 0.0559248f $X=3.335 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_507_n N_A_217_65#_c_567_n 0.0313184f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_M1003_d N_A_217_65#_c_568_n 0.00176461f $X=3.36 $Y=0.325 $X2=0
+ $Y2=0
cc_307 N_VGND_c_499_n N_A_217_65#_c_568_n 0.0170777f $X=3.5 $Y=0.45 $X2=0 $Y2=0
cc_308 N_VGND_c_499_n N_A_217_65#_c_570_n 0.0251314f $X=3.5 $Y=0.45 $X2=0 $Y2=0
cc_309 N_VGND_c_500_n N_A_217_65#_c_570_n 0.0247562f $X=4.36 $Y=0.45 $X2=0 $Y2=0
cc_310 N_VGND_c_503_n N_A_217_65#_c_570_n 0.0113237f $X=4.195 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_507_n N_A_217_65#_c_570_n 0.00720172f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_M1010_d N_A_217_65#_c_571_n 0.00176773f $X=4.22 $Y=0.325 $X2=0
+ $Y2=0
cc_313 N_VGND_c_500_n N_A_217_65#_c_571_n 0.0171443f $X=4.36 $Y=0.45 $X2=0 $Y2=0
cc_314 N_VGND_c_500_n N_A_217_65#_c_572_n 0.0232759f $X=4.36 $Y=0.45 $X2=0 $Y2=0
cc_315 N_VGND_c_506_n N_A_217_65#_c_572_n 0.0140356f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_507_n N_A_217_65#_c_572_n 0.00977851f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_501_n N_A_217_65#_c_573_n 0.0235159f $X=3.335 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_c_507_n N_A_217_65#_c_573_n 0.0127052f $X=5.04 $Y=0 $X2=0 $Y2=0
