* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o41a_m A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_300_51# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_444_535# A2 a_516_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_516_535# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND A3 a_300_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_300_51# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND A1 a_300_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_80_21# A4 a_329_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_329_535# A3 a_444_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_80_21# B1 a_300_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
