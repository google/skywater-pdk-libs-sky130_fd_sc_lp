* File: sky130_fd_sc_lp__mux4_m.pex.spice
* Created: Fri Aug 28 10:46:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX4_M%A2 3 7 11 12 13 14 15 16 22
c40 11 0 1.4009e-19 $X=1.2 $Y=1.99
r41 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=2.405 $X2=1.2
+ $Y2=2.775
r42 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=2.035 $X2=1.2
+ $Y2=2.405
r43 13 14 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.2 $Y=1.65 $X2=1.2
+ $Y2=2.035
r44 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=1.65
+ $X2=1.2 $Y2=1.65
r45 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.2 $Y=1.99 $X2=1.2
+ $Y2=1.65
r46 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.99 $X2=1.2
+ $Y2=2.155
r47 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.485
+ $X2=1.2 $Y2=1.65
r48 7 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.29 $Y=2.525
+ $X2=1.29 $Y2=2.155
r49 3 10 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=1.29 $Y=0.84
+ $X2=1.29 $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A_59_463# 1 2 9 12 16 20 23 25 27 31 33 36 39
+ 40 42 43 45 46 47 50 54 58 63
c144 58 0 1.02967e-19 $X=1.672 $Y=1.22
c145 50 0 1.36796e-19 $X=3.61 $Y=1.715
c146 16 0 1.94979e-19 $X=3.52 $Y=2.525
r147 56 57 4.90862 $w=3.83e-07 $l=8.5e-08 $layer=LI1_cond $X=0.507 $Y=1.22
+ $X2=0.507 $Y2=1.305
r148 54 56 9.42908 $w=3.83e-07 $l=3.15e-07 $layer=LI1_cond $X=0.507 $Y=0.905
+ $X2=0.507 $Y2=1.22
r149 51 63 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.61 $Y=1.715
+ $X2=3.795 $Y2=1.715
r150 51 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.61 $Y=1.715
+ $X2=3.52 $Y2=1.715
r151 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.61
+ $Y=1.715 $X2=3.61 $Y2=1.715
r152 48 50 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.61 $Y=1.27
+ $X2=3.61 $Y2=1.715
r153 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.525 $Y=1.185
+ $X2=3.61 $Y2=1.27
r154 46 47 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.525 $Y=1.185
+ $X2=2.525 $Y2=1.185
r155 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.44 $Y=1.1
+ $X2=2.525 $Y2=1.185
r156 44 45 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.44 $Y=0.445
+ $X2=2.44 $Y2=1.1
r157 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.355 $Y=0.36
+ $X2=2.44 $Y2=0.445
r158 42 43 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.355 $Y=0.36
+ $X2=1.69 $Y2=0.36
r159 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.74
+ $Y=1.325 $X2=1.74 $Y2=1.325
r160 37 58 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=1.672 $Y=1.305
+ $X2=1.672 $Y2=1.22
r161 37 39 0.7557 $w=3.03e-07 $l=2e-08 $layer=LI1_cond $X=1.672 $Y=1.305
+ $X2=1.672 $Y2=1.325
r162 36 58 3.87901 $w=2.37e-07 $l=1.13666e-07 $layer=LI1_cond $X=1.605 $Y=1.135
+ $X2=1.672 $Y2=1.22
r163 35 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.605 $Y=0.445
+ $X2=1.69 $Y2=0.36
r164 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.605 $Y=0.445
+ $X2=1.605 $Y2=1.135
r165 34 56 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.7 $Y=1.22
+ $X2=0.507 $Y2=1.22
r166 33 58 2.57001 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.52 $Y=1.22
+ $X2=1.672 $Y2=1.22
r167 33 34 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.52 $Y=1.22
+ $X2=0.7 $Y2=1.22
r168 31 57 61 $w=2.08e-07 $l=1.155e-06 $layer=LI1_cond $X=0.42 $Y=2.46 $X2=0.42
+ $Y2=1.305
r169 25 40 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.74 $Y=1.68
+ $X2=1.74 $Y2=1.325
r170 25 27 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.74 $Y=1.755
+ $X2=2.08 $Y2=1.755
r171 23 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.16
+ $X2=1.74 $Y2=1.325
r172 18 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.55
+ $X2=3.795 $Y2=1.715
r173 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.795 $Y=1.55
+ $X2=3.795 $Y2=0.84
r174 14 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.88
+ $X2=3.52 $Y2=1.715
r175 14 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.52 $Y=1.88
+ $X2=3.52 $Y2=2.525
r176 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.08 $Y=1.83
+ $X2=2.08 $Y2=1.755
r177 10 12 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.08 $Y=1.83
+ $X2=2.08 $Y2=2.525
r178 9 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.65 $Y=0.84
+ $X2=1.65 $Y2=1.16
r179 2 31 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.295
+ $Y=2.315 $X2=0.42 $Y2=2.46
r180 1 54 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.41
+ $Y=0.63 $X2=0.535 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A3 3 7 11 12 13 16
r45 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.53
+ $Y=1.555 $X2=2.53 $Y2=1.555
r46 13 17 2.57978 $w=5.08e-07 $l=1.1e-07 $layer=LI1_cond $X=2.64 $Y=1.725
+ $X2=2.53 $Y2=1.725
r47 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.53 $Y=1.895
+ $X2=2.53 $Y2=1.555
r48 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.53 $Y=1.895
+ $X2=2.53 $Y2=2.06
r49 10 16 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.53 $Y=1.39
+ $X2=2.53 $Y2=1.555
r50 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.55 $Y=0.84 $X2=2.55
+ $Y2=1.39
r51 3 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.44 $Y=2.525
+ $X2=2.44 $Y2=2.06
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A1 3 7 11 12 13 16 17
r42 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.07
+ $Y=1.555 $X2=3.07 $Y2=1.555
r43 13 17 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.07 $Y=1.665
+ $X2=3.07 $Y2=1.555
r44 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.07 $Y=1.895
+ $X2=3.07 $Y2=1.555
r45 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.895
+ $X2=3.07 $Y2=2.06
r46 10 16 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.39
+ $X2=3.07 $Y2=1.555
r47 7 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.16 $Y=2.525
+ $X2=3.16 $Y2=2.06
r48 3 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.005 $Y=0.84
+ $X2=3.005 $Y2=1.39
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%S0 3 8 9 13 15 16 19 21 25 27 31 33 36 39 41
+ 42 43 46 49 51 55
c135 19 0 1.02967e-19 $X=2.19 $Y=0.84
r136 49 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.24 $Y=0.555
+ $X2=0.24 $Y2=0.35
r137 47 54 45.9721 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=0.35
+ $X2=0.585 $Y2=0.515
r138 47 51 18.3916 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=0.35
+ $X2=0.585 $Y2=0.185
r139 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=0.35 $X2=0.51 $Y2=0.35
r140 44 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.325 $Y=0.35
+ $X2=0.24 $Y2=0.35
r141 44 46 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.325 $Y=0.35
+ $X2=0.51 $Y2=0.35
r142 37 39 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=0.635 $Y=1.235
+ $X2=0.75 $Y2=1.235
r143 35 36 1443.44 $w=1.5e-07 $l=2.815e-06 $layer=POLY_cond $X=4.935 $Y=0.26
+ $X2=4.935 $Y2=3.075
r144 34 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.025 $Y=3.15
+ $X2=3.95 $Y2=3.15
r145 33 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.86 $Y=3.15
+ $X2=4.935 $Y2=3.075
r146 33 34 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=4.86 $Y=3.15
+ $X2=4.025 $Y2=3.15
r147 29 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.95 $Y=3.075
+ $X2=3.95 $Y2=3.15
r148 29 31 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.95 $Y=3.075
+ $X2=3.95 $Y2=2.525
r149 28 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.44 $Y=0.185
+ $X2=3.365 $Y2=0.185
r150 27 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.86 $Y=0.185
+ $X2=4.935 $Y2=0.26
r151 27 28 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=4.86 $Y=0.185
+ $X2=3.44 $Y2=0.185
r152 23 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=0.26
+ $X2=3.365 $Y2=0.185
r153 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.365 $Y=0.26
+ $X2=3.365 $Y2=0.84
r154 22 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.265 $Y=0.185
+ $X2=2.19 $Y2=0.185
r155 21 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.29 $Y=0.185
+ $X2=3.365 $Y2=0.185
r156 21 22 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=3.29 $Y=0.185
+ $X2=2.265 $Y2=0.185
r157 17 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.19 $Y=0.26
+ $X2=2.19 $Y2=0.185
r158 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.19 $Y=0.26
+ $X2=2.19 $Y2=0.84
r159 15 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.875 $Y=3.15
+ $X2=3.95 $Y2=3.15
r160 15 16 1102.45 $w=1.5e-07 $l=2.15e-06 $layer=POLY_cond $X=3.875 $Y=3.15
+ $X2=1.725 $Y2=3.15
r161 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.65 $Y=3.075
+ $X2=1.725 $Y2=3.15
r162 11 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.65 $Y=3.075
+ $X2=1.65 $Y2=2.525
r163 10 51 30.3798 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.825 $Y=0.185
+ $X2=0.585 $Y2=0.185
r164 9 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.115 $Y=0.185
+ $X2=2.19 $Y2=0.185
r165 9 10 661.468 $w=1.5e-07 $l=1.29e-06 $layer=POLY_cond $X=2.115 $Y=0.185
+ $X2=0.825 $Y2=0.185
r166 8 54 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.75 $Y=0.84
+ $X2=0.75 $Y2=0.515
r167 6 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.75 $Y=1.16
+ $X2=0.75 $Y2=1.235
r168 6 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.75 $Y=1.16 $X2=0.75
+ $Y2=0.84
r169 1 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.635 $Y=1.31
+ $X2=0.635 $Y2=1.235
r170 1 3 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=0.635 $Y=1.31
+ $X2=0.635 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A0 1 3 6 8 11
c33 6 0 1.36796e-19 $X=4.31 $Y=2.525
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.4
+ $Y=1.325 $X2=4.4 $Y2=1.325
r35 11 13 15.9485 $w=2.72e-07 $l=9e-08 $layer=POLY_cond $X=4.31 $Y=1.325 $X2=4.4
+ $Y2=1.325
r36 8 14 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.56 $Y=1.325 $X2=4.4
+ $Y2=1.325
r37 4 11 16.6763 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.31 $Y=1.49
+ $X2=4.31 $Y2=1.325
r38 4 6 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=4.31 $Y=1.49
+ $X2=4.31 $Y2=2.525
r39 1 11 27.4669 $w=2.72e-07 $l=2.29783e-07 $layer=POLY_cond $X=4.155 $Y=1.16
+ $X2=4.31 $Y2=1.325
r40 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.155 $Y=1.16
+ $X2=4.155 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A_1118_37# 1 2 10 12 15 17 20 22 25 29 31 40
r70 39 40 31.0318 $w=3.4e-07 $l=7.5e-08 $layer=POLY_cond $X=6.275 $Y=1.965
+ $X2=6.2 $Y2=1.965
r71 31 34 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=7.04 $Y=0.35 $X2=7.04
+ $Y2=0.43
r72 27 29 38.29 $w=2.08e-07 $l=7.25e-07 $layer=LI1_cond $X=7.04 $Y=2.055
+ $X2=7.04 $Y2=2.78
r73 25 39 39.8838 $w=3.4e-07 $l=2.35e-07 $layer=POLY_cond $X=6.51 $Y=1.965
+ $X2=6.275 $Y2=1.965
r74 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.51
+ $Y=1.97 $X2=6.51 $Y2=1.97
r75 22 27 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.935 $Y=1.97
+ $X2=7.04 $Y2=2.055
r76 22 24 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.935 $Y=1.97
+ $X2=6.51 $Y2=1.97
r77 20 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.755 $Y=0.35
+ $X2=5.755 $Y2=0.515
r78 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.755
+ $Y=0.35 $X2=5.755 $Y2=0.35
r79 17 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.935 $Y=0.35
+ $X2=7.04 $Y2=0.35
r80 17 19 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=6.935 $Y=0.35
+ $X2=5.755 $Y2=0.35
r81 13 39 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.275 $Y=2.135
+ $X2=6.275 $Y2=1.965
r82 13 15 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.275 $Y=2.135
+ $X2=6.275 $Y2=2.525
r83 12 40 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.92 $Y=1.87 $X2=6.2
+ $Y2=1.87
r84 10 38 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.845 $Y=1.065
+ $X2=5.845 $Y2=0.515
r85 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.845 $Y=1.795
+ $X2=5.92 $Y2=1.87
r86 8 10 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.845 $Y=1.795
+ $X2=5.845 $Y2=1.065
r87 2 29 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.915
+ $Y=2.635 $X2=7.04 $Y2=2.78
r88 1 34 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=6.915
+ $Y=0.235 $X2=7.04 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%S1 3 5 6 7 9 10 11 13 15 16 18 19 21 25 30 33
+ 34 37
c84 25 0 1.248e-19 $X=7.255 $Y=2.45
r85 34 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.96
+ $Y=0.93 $X2=6.96 $Y2=0.93
r86 32 37 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=6.96 $Y=1.385
+ $X2=6.96 $Y2=0.93
r87 32 33 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=6.96 $Y=1.385
+ $X2=6.96 $Y2=1.46
r88 28 37 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.96 $Y=0.915
+ $X2=6.96 $Y2=0.93
r89 28 30 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=6.96 $Y=0.84
+ $X2=7.255 $Y2=0.84
r90 24 25 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=7.05 $Y=2.45
+ $X2=7.255 $Y2=2.45
r91 22 24 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.765 $Y=2.45
+ $X2=7.05 $Y2=2.45
r92 19 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.255 $Y=2.525
+ $X2=7.255 $Y2=2.45
r93 19 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.255 $Y=2.525
+ $X2=7.255 $Y2=2.845
r94 16 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.255 $Y=0.765
+ $X2=7.255 $Y2=0.84
r95 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.255 $Y=0.765
+ $X2=7.255 $Y2=0.445
r96 15 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.05 $Y=2.375
+ $X2=7.05 $Y2=2.45
r97 14 33 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.05 $Y=1.535
+ $X2=6.96 $Y2=1.46
r98 14 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.05 $Y=1.535
+ $X2=7.05 $Y2=2.375
r99 12 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.765 $Y=2.525
+ $X2=6.765 $Y2=2.45
r100 12 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.765 $Y=2.525
+ $X2=6.765 $Y2=3.075
r101 10 33 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.46
+ $X2=6.96 $Y2=1.46
r102 10 11 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.795 $Y=1.46
+ $X2=6.35 $Y2=1.46
r103 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.275 $Y=1.385
+ $X2=6.35 $Y2=1.46
r104 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.275 $Y=1.385
+ $X2=6.275 $Y2=1.065
r105 5 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.69 $Y=3.15
+ $X2=6.765 $Y2=3.075
r106 5 6 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.69 $Y=3.15 $X2=5.92
+ $Y2=3.15
r107 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.845 $Y=3.075
+ $X2=5.92 $Y2=3.15
r108 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.845 $Y=3.075
+ $X2=5.845 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A_1184_171# 1 2 8 11 15 19 23 25 27 29 30 32
+ 35
r61 35 39 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=7.562 $Y=1.695
+ $X2=7.562 $Y2=1.86
r62 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.53
+ $Y=1.695 $X2=7.53 $Y2=1.695
r63 30 37 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=7.562 $Y=1.355
+ $X2=7.562 $Y2=1.19
r64 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.53
+ $Y=1.355 $X2=7.53 $Y2=1.355
r65 27 34 3.40825 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=7.53 $Y=1.535
+ $X2=7.53 $Y2=1.697
r66 27 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.53 $Y=1.535
+ $X2=7.53 $Y2=1.355
r67 26 32 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.165 $Y=1.62
+ $X2=6.07 $Y2=1.62
r68 25 34 3.40825 $w=1.7e-07 $l=1.17346e-07 $layer=LI1_cond $X=7.445 $Y=1.62
+ $X2=7.53 $Y2=1.697
r69 25 26 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=7.445 $Y=1.62
+ $X2=6.165 $Y2=1.62
r70 21 32 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=1.705
+ $X2=6.07 $Y2=1.62
r71 21 23 44.0718 $w=1.88e-07 $l=7.55e-07 $layer=LI1_cond $X=6.07 $Y=1.705
+ $X2=6.07 $Y2=2.46
r72 17 32 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=1.535
+ $X2=6.07 $Y2=1.62
r73 17 19 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=6.07 $Y=1.535
+ $X2=6.07 $Y2=1.13
r74 15 39 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=7.685 $Y=2.845
+ $X2=7.685 $Y2=1.86
r75 11 37 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=7.685 $Y=0.445
+ $X2=7.685 $Y2=1.19
r76 8 35 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=7.562 $Y=1.663
+ $X2=7.562 $Y2=1.695
r77 7 30 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=7.562 $Y=1.387
+ $X2=7.562 $Y2=1.355
r78 7 8 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=7.562 $Y=1.387
+ $X2=7.562 $Y2=1.663
r79 2 23 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=2.315 $X2=6.06 $Y2=2.46
r80 1 19 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.92
+ $Y=0.855 $X2=6.06 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 35 41 55
+ 61 62 65 68
c84 62 0 1.248e-19 $X=7.92 $Y=3.33
r85 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r86 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 62 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r88 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r89 59 68 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.47 $Y2=3.33
r90 59 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.92 $Y2=3.33
r91 58 69 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r92 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r93 55 68 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.365 $Y=3.33
+ $X2=7.47 $Y2=3.33
r94 55 57 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=7.365 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 54 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r96 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 51 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 48 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.66 $Y2=3.33
r101 48 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=3.12 $Y2=3.33
r102 47 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r106 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 41 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=3.33
+ $X2=2.66 $Y2=3.33
r108 41 46 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 39 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 35 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 35 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 33 53 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.66 $Y2=3.33
r115 32 57 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.66 $Y2=3.33
r117 30 38 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 30 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.84 $Y2=3.33
r119 29 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 29 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.84 $Y2=3.33
r121 25 68 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=3.245
+ $X2=7.47 $Y2=3.33
r122 25 27 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=7.47 $Y=3.245
+ $X2=7.47 $Y2=2.91
r123 21 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=3.245
+ $X2=4.66 $Y2=3.33
r124 21 23 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.66 $Y=3.245
+ $X2=4.66 $Y2=2.59
r125 17 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=3.245
+ $X2=2.66 $Y2=3.33
r126 17 19 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.66 $Y=3.245
+ $X2=2.66 $Y2=2.61
r127 13 31 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=3.245
+ $X2=0.84 $Y2=3.33
r128 13 15 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=0.84 $Y=3.245
+ $X2=0.84 $Y2=2.59
r129 4 27 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=7.33
+ $Y=2.635 $X2=7.47 $Y2=2.91
r130 3 23 600 $w=1.7e-07 $l=3.88909e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=2.315 $X2=4.66 $Y2=2.59
r131 2 19 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=2.315 $X2=2.66 $Y2=2.61
r132 1 15 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=2.315 $X2=0.85 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A_345_126# 1 2 3 4 15 18 19 20 22 23 24 26 27
+ 28 30 31 32 34 35 36 37 41 45 53 55
c156 22 0 6.53158e-20 $X=3.09 $Y=2.745
r157 51 53 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.975 $Y=0.79
+ $X2=2.09 $Y2=0.79
r158 43 45 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=6.49 $Y=2.805
+ $X2=6.49 $Y2=2.59
r159 39 41 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=6.49 $Y=0.785
+ $X2=6.49 $Y2=1
r160 38 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.795 $Y=2.89
+ $X2=5.71 $Y2=2.89
r161 37 43 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.385 $Y=2.89
+ $X2=6.49 $Y2=2.805
r162 37 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.385 $Y=2.89
+ $X2=5.795 $Y2=2.89
r163 35 39 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.385 $Y=0.7
+ $X2=6.49 $Y2=0.785
r164 35 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.385 $Y=0.7
+ $X2=5.795 $Y2=0.7
r165 34 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=2.805
+ $X2=5.71 $Y2=2.89
r166 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.71 $Y=0.785
+ $X2=5.795 $Y2=0.7
r167 33 34 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=5.71 $Y=0.785
+ $X2=5.71 $Y2=2.805
r168 31 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=2.89
+ $X2=5.71 $Y2=2.89
r169 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.625 $Y=2.89
+ $X2=5.095 $Y2=2.89
r170 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.01 $Y=2.805
+ $X2=5.095 $Y2=2.89
r171 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.01 $Y=2.245
+ $X2=5.01 $Y2=2.805
r172 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.925 $Y=2.16
+ $X2=5.01 $Y2=2.245
r173 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.925 $Y=2.16
+ $X2=4.395 $Y2=2.16
r174 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.31 $Y=2.245
+ $X2=4.395 $Y2=2.16
r175 25 26 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.31 $Y=2.245
+ $X2=4.31 $Y2=2.745
r176 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.225 $Y=2.83
+ $X2=4.31 $Y2=2.745
r177 23 24 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=4.225 $Y=2.83
+ $X2=3.175 $Y2=2.83
r178 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.09 $Y=2.745
+ $X2=3.175 $Y2=2.83
r179 21 22 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.09 $Y=2.345
+ $X2=3.09 $Y2=2.745
r180 20 49 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=2.26
+ $X2=2.09 $Y2=2.26
r181 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.005 $Y=2.26
+ $X2=3.09 $Y2=2.345
r182 19 20 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.005 $Y=2.26
+ $X2=2.175 $Y2=2.26
r183 18 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=2.175
+ $X2=2.09 $Y2=2.26
r184 17 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=0.955
+ $X2=2.09 $Y2=0.79
r185 17 18 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=2.09 $Y=0.955
+ $X2=2.09 $Y2=2.175
r186 13 49 13.5701 $w=1.68e-07 $l=2.08e-07 $layer=LI1_cond $X=1.882 $Y=2.26
+ $X2=2.09 $Y2=2.26
r187 13 15 5.40943 $w=2.43e-07 $l=1.15e-07 $layer=LI1_cond $X=1.882 $Y=2.345
+ $X2=1.882 $Y2=2.46
r188 4 45 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=2.315 $X2=6.49 $Y2=2.59
r189 3 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=2.315 $X2=1.865 $Y2=2.46
r190 2 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.35
+ $Y=0.855 $X2=6.49 $Y2=1
r191 1 51 182 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.63 $X2=1.975 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%A_688_126# 1 2 3 4 13 17 22 24 25 29 33 35 36
c61 35 0 1.94979e-19 $X=3.96 $Y=1.81
r62 31 36 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=5.36 $Y=1.895
+ $X2=5.35 $Y2=1.81
r63 31 33 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.36 $Y=1.895
+ $X2=5.36 $Y2=2.46
r64 27 36 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=1.725
+ $X2=5.35 $Y2=1.81
r65 27 29 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=5.35 $Y=1.725
+ $X2=5.35 $Y2=1.13
r66 26 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=1.81
+ $X2=3.96 $Y2=1.81
r67 25 36 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.255 $Y=1.81
+ $X2=5.35 $Y2=1.81
r68 25 26 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=5.255 $Y=1.81
+ $X2=4.045 $Y2=1.81
r69 23 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=1.895
+ $X2=3.96 $Y2=1.81
r70 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.96 $Y=1.895
+ $X2=3.96 $Y2=2.355
r71 22 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=1.725
+ $X2=3.96 $Y2=1.81
r72 21 22 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=3.96 $Y=0.92
+ $X2=3.96 $Y2=1.725
r73 17 24 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.875 $Y=2.46
+ $X2=3.96 $Y2=2.355
r74 17 19 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=3.875 $Y=2.46
+ $X2=3.735 $Y2=2.46
r75 13 21 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.875 $Y=0.815
+ $X2=3.96 $Y2=0.92
r76 13 15 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.875 $Y=0.815
+ $X2=3.58 $Y2=0.815
r77 4 33 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=2.315 $X2=5.36 $Y2=2.46
r78 3 19 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.595
+ $Y=2.315 $X2=3.735 $Y2=2.46
r79 2 29 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=5.235
+ $Y=0.855 $X2=5.36 $Y2=1.13
r80 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.63 $X2=3.58 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%X 1 2 7 8 9 10 11 12 20
r13 11 12 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=7.9 $Y=2.405 $X2=7.9
+ $Y2=2.775
r14 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=7.9 $Y=2.035 $X2=7.9
+ $Y2=2.405
r15 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=7.9 $Y=1.665 $X2=7.9
+ $Y2=2.035
r16 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=7.9 $Y=1.295 $X2=7.9
+ $Y2=1.665
r17 7 8 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=7.9 $Y=0.925 $X2=7.9
+ $Y2=1.295
r18 7 20 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=7.9 $Y=0.925 $X2=7.9
+ $Y2=0.51
r19 2 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.635 $X2=7.9 $Y2=2.78
r20 1 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.235 $X2=7.9 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_M%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 37 52
+ 58 59 62 65
r82 65 66 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r83 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r84 59 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r85 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r86 56 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.575 $Y=0 $X2=7.48
+ $Y2=0
r87 56 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.575 $Y=0 $X2=7.92
+ $Y2=0
r88 55 66 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=7.44
+ $Y2=0
r89 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r90 52 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.385 $Y=0 $X2=7.48
+ $Y2=0
r91 52 54 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=7.385 $Y=0
+ $X2=4.56 $Y2=0
r92 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r93 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r94 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r95 45 63 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.2
+ $Y2=0
r96 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r97 42 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=0 $X2=1.045
+ $Y2=0
r98 42 44 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.21 $Y=0 $X2=2.64
+ $Y2=0
r99 40 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r100 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 37 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.045
+ $Y2=0
r102 37 39 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.72
+ $Y2=0
r103 35 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r104 35 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r105 35 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r106 33 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.265 $Y=0
+ $X2=4.08 $Y2=0
r107 33 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.37
+ $Y2=0
r108 32 54 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.56
+ $Y2=0
r109 32 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.37
+ $Y2=0
r110 30 44 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.64
+ $Y2=0
r111 30 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.8
+ $Y2=0
r112 29 47 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.895 $Y=0
+ $X2=3.12 $Y2=0
r113 29 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.895 $Y=0 $X2=2.8
+ $Y2=0
r114 25 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.48 $Y=0.085
+ $X2=7.48 $Y2=0
r115 25 27 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=7.48 $Y=0.085
+ $X2=7.48 $Y2=0.38
r116 21 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0
r117 21 23 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0.775
r118 17 31 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0
r119 17 19 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0.755
r120 13 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=0.085
+ $X2=1.045 $Y2=0
r121 13 15 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=1.045 $Y=0.085
+ $X2=1.045 $Y2=0.775
r122 4 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.235 $X2=7.47 $Y2=0.38
r123 3 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.23
+ $Y=0.63 $X2=4.37 $Y2=0.775
r124 2 19 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.63 $X2=2.79 $Y2=0.755
r125 1 15 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=0.825
+ $Y=0.63 $X2=1.045 $Y2=0.775
.ends

