* File: sky130_fd_sc_lp__dlrbp_lp.pex.spice
* Created: Wed Sep  2 09:46:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%D 3 7 11 15 17 18 19 23
r40 18 19 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.667 $Y=1.295
+ $X2=0.667 $Y2=1.665
r41 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.665
+ $Y=1.345 $X2=0.665 $Y2=1.345
r42 16 23 40.6942 $w=4.1e-07 $l=3e-07 $layer=POLY_cond $X=0.625 $Y=1.645
+ $X2=0.625 $Y2=1.345
r43 16 17 36.2176 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.625 $Y=1.645
+ $X2=0.625 $Y2=1.85
r44 15 23 2.03471 $w=4.1e-07 $l=1.5e-08 $layer=POLY_cond $X=0.625 $Y=1.33
+ $X2=0.625 $Y2=1.345
r45 7 17 185.098 $w=2.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.705 $Y=2.595
+ $X2=0.705 $Y2=1.85
r46 1 15 24.4548 $w=4.1e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=1.18
+ $X2=0.675 $Y2=1.33
r47 1 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.855 $Y=1.18
+ $X2=0.855 $Y2=0.77
r48 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%GATE 3 7 13 15 16 17 18 22
c47 13 0 1.42163e-19 $X=1.645 $Y=0.77
r48 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.51
+ $Y=1.345 $X2=1.51 $Y2=1.345
r49 18 23 6.48721 $w=5.88e-07 $l=3.2e-07 $layer=LI1_cond $X=1.38 $Y=1.665
+ $X2=1.38 $Y2=1.345
r50 17 23 1.01363 $w=5.88e-07 $l=5e-08 $layer=LI1_cond $X=1.38 $Y=1.295 $X2=1.38
+ $Y2=1.345
r51 15 16 29.6612 $w=5.1e-07 $l=1.5e-07 $layer=POLY_cond $X=1.415 $Y=1.7
+ $X2=1.415 $Y2=1.85
r52 11 22 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=1.645 $Y=1.18
+ $X2=1.465 $Y2=1.345
r53 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.645 $Y=1.18
+ $X2=1.645 $Y2=0.77
r54 9 22 9.4417 $w=5.1e-07 $l=9e-08 $layer=POLY_cond $X=1.465 $Y=1.435 $X2=1.465
+ $Y2=1.345
r55 9 15 27.8006 $w=5.1e-07 $l=2.65e-07 $layer=POLY_cond $X=1.465 $Y=1.435
+ $X2=1.465 $Y2=1.7
r56 5 22 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=1.285 $Y=1.18
+ $X2=1.465 $Y2=1.345
r57 5 7 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.285 $Y=1.18
+ $X2=1.285 $Y2=0.77
r58 3 16 185.098 $w=2.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.235 $Y=2.595
+ $X2=1.235 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%A_272_419# 1 2 9 13 17 21 25 27 30 31 33 34
+ 35 37 38 39 40 42 46 48 51 58 60 61 68
c161 27 0 1.20621e-19 $X=1.855 $Y=2.25
r162 64 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.635 $Y=1.3
+ $X2=2.725 $Y2=1.3
r163 61 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.03
+ $X2=4.735 $Y2=0.865
r164 60 63 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=1.03
+ $X2=4.735 $Y2=1.195
r165 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.735
+ $Y=1.03 $X2=4.735 $Y2=1.03
r166 58 72 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.51
+ $X2=3.835 $Y2=1.675
r167 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.835
+ $Y=1.51 $X2=3.835 $Y2=1.51
r168 54 68 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.81 $Y=1.3
+ $X2=2.995 $Y2=1.3
r169 54 66 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=2.81 $Y=1.3
+ $X2=2.725 $Y2=1.3
r170 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=1.3 $X2=2.81 $Y2=1.3
r171 48 50 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.86 $Y=0.77
+ $X2=1.86 $Y2=1
r172 44 46 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.5 $Y=2.205
+ $X2=1.665 $Y2=2.205
r173 42 63 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=4.815 $Y=2.895
+ $X2=4.815 $Y2=1.195
r174 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.73 $Y=2.98
+ $X2=4.815 $Y2=2.895
r175 39 40 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.73 $Y=2.98 $X2=4
+ $Y2=2.98
r176 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.835 $Y=2.895
+ $X2=4 $Y2=2.98
r177 37 57 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=1.675
+ $X2=3.835 $Y2=1.51
r178 37 38 42.6055 $w=3.28e-07 $l=1.22e-06 $layer=LI1_cond $X=3.835 $Y=1.675
+ $X2=3.835 $Y2=2.895
r179 36 53 9.59551 $w=2.67e-07 $l=2.1e-07 $layer=LI1_cond $X=2.81 $Y=1.51
+ $X2=2.81 $Y2=1.3
r180 35 57 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.67 $Y=1.51
+ $X2=3.835 $Y2=1.51
r181 35 36 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.67 $Y=1.51
+ $X2=2.975 $Y2=1.51
r182 33 36 9.14344 $w=2.67e-07 $l=2.0106e-07 $layer=LI1_cond $X=2.89 $Y=1.675
+ $X2=2.81 $Y2=1.51
r183 33 34 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.89 $Y=1.675
+ $X2=2.89 $Y2=2.165
r184 32 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.25
+ $X2=1.94 $Y2=2.25
r185 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.805 $Y=2.25
+ $X2=2.89 $Y2=2.165
r186 31 32 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.805 $Y=2.25
+ $X2=2.025 $Y2=2.25
r187 30 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.165
+ $X2=1.94 $Y2=2.25
r188 30 50 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=1.94 $Y=2.165
+ $X2=1.94 $Y2=1
r189 27 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.25
+ $X2=1.94 $Y2=2.25
r190 27 46 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=2.25
+ $X2=1.665 $Y2=2.25
r191 25 74 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.645 $Y=0.455
+ $X2=4.645 $Y2=0.865
r192 21 72 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.825 $Y=2.335
+ $X2=3.825 $Y2=1.675
r193 15 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.995 $Y=1.135
+ $X2=2.995 $Y2=1.3
r194 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.995 $Y=1.135
+ $X2=2.995 $Y2=0.455
r195 11 66 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.465
+ $X2=2.725 $Y2=1.3
r196 11 13 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.725 $Y=1.465
+ $X2=2.725 $Y2=2.175
r197 7 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.135
+ $X2=2.635 $Y2=1.3
r198 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.635 $Y=1.135
+ $X2=2.635 $Y2=0.455
r199 2 44 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=2.095 $X2=1.5 $Y2=2.245
r200 1 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.56 $X2=1.86 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%A_27_112# 1 2 7 9 12 17 19 21 24 28 29 32
+ 36 37
c85 29 0 1.20621e-19 $X=1.99 $Y=2.9
c86 19 0 1.62324e-20 $X=3.335 $Y=1.705
c87 17 0 6.01512e-20 $X=3.425 $Y=0.455
r88 36 38 8.78751 $w=4.88e-07 $l=3.6e-07 $layer=LI1_cond $X=0.36 $Y=2.24
+ $X2=0.36 $Y2=2.6
r89 36 37 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.36 $Y=2.24
+ $X2=0.36 $Y2=2.075
r90 34 37 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=0.2 $Y=1 $X2=0.2
+ $Y2=2.075
r91 32 34 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.28 $Y=0.77
+ $X2=0.28 $Y2=1
r92 29 42 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.99 $Y=2.9 $X2=1.99
+ $Y2=3.12
r93 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=2.9 $X2=1.99 $Y2=2.9
r94 26 28 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.99 $Y=2.685
+ $X2=1.99 $Y2=2.9
r95 25 38 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.605 $Y=2.6
+ $X2=0.36 $Y2=2.6
r96 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.825 $Y=2.6
+ $X2=1.99 $Y2=2.685
r97 24 25 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=1.825 $Y=2.6
+ $X2=0.605 $Y2=2.6
r98 20 21 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=3.405 $Y=0.955
+ $X2=3.405 $Y2=1.105
r99 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.385 $Y=1.705
+ $X2=3.385 $Y2=1.105
r100 17 20 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.425 $Y=0.455
+ $X2=3.425 $Y2=0.955
r101 10 12 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.335 $Y=3.045
+ $X2=3.335 $Y2=2.335
r102 9 19 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.335 $Y=1.83
+ $X2=3.335 $Y2=1.705
r103 9 12 125.469 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.335 $Y=1.83
+ $X2=3.335 $Y2=2.335
r104 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=3.12
+ $X2=1.99 $Y2=3.12
r105 7 10 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.21 $Y=3.12
+ $X2=3.335 $Y2=3.045
r106 7 8 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=3.21 $Y=3.12
+ $X2=2.155 $Y2=3.12
r107 2 36 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.295
+ $Y=2.095 $X2=0.44 $Y2=2.24
r108 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%A_455_49# 1 2 9 10 13 14 15 18 22 25 28 32
+ 35 36 37 40
c94 35 0 6.01512e-20 $X=3.875 $Y=0.94
c95 32 0 1.62324e-20 $X=2.46 $Y=1.82
c96 25 0 1.42163e-19 $X=2.34 $Y=1.655
c97 18 0 1.80631e-19 $X=4.65 $Y=2.335
r98 36 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.875 $Y=0.94
+ $X2=3.875 $Y2=1.03
r99 36 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=0.94
+ $X2=3.875 $Y2=0.775
r100 35 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=0.94
+ $X2=3.71 $Y2=0.94
r101 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.875
+ $Y=0.94 $X2=3.875 $Y2=0.94
r102 29 32 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.34 $Y=1.82
+ $X2=2.46 $Y2=1.82
r103 27 28 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=0.87
+ $X2=2.42 $Y2=0.87
r104 27 37 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=2.585 $Y=0.87
+ $X2=3.71 $Y2=0.87
r105 25 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=1.655
+ $X2=2.34 $Y2=1.82
r106 24 28 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.34 $Y=0.955
+ $X2=2.42 $Y2=0.87
r107 24 25 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.34 $Y=0.955
+ $X2=2.34 $Y2=1.655
r108 20 28 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=0.785
+ $X2=2.42 $Y2=0.87
r109 20 22 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.42 $Y=0.785
+ $X2=2.42 $Y2=0.475
r110 16 18 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=4.65 $Y=1.585
+ $X2=4.65 $Y2=2.335
r111 14 16 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=4.525 $Y=1.51
+ $X2=4.65 $Y2=1.585
r112 14 15 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.525 $Y=1.51
+ $X2=4.36 $Y2=1.51
r113 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.285 $Y=1.435
+ $X2=4.36 $Y2=1.51
r114 12 13 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.285 $Y=1.105
+ $X2=4.285 $Y2=1.435
r115 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.04 $Y=1.03
+ $X2=3.875 $Y2=1.03
r116 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.21 $Y=1.03
+ $X2=4.285 $Y2=1.105
r117 10 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.21 $Y=1.03
+ $X2=4.04 $Y2=1.03
r118 9 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.815 $Y=0.455
+ $X2=3.815 $Y2=0.775
r119 2 32 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.675 $X2=2.46 $Y2=1.82
r120 1 22 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.245 $X2=2.42 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%A_1028_23# 1 2 9 13 17 21 25 27 28 29 31 34
+ 36 38 45 48 52 53 55 56 59 62 64 65 69 70 75 78 79
c169 78 0 1.86549e-19 $X=6.18 $Y=1.88
c170 56 0 1.80631e-19 $X=5.47 $Y=1.8
c171 34 0 1.76362e-19 $X=8.74 $Y=2.37
c172 17 0 1.87193e-19 $X=7.06 $Y=2.235
r173 73 75 6.97531 $w=3.78e-07 $l=2.3e-07 $layer=LI1_cond $X=6.075 $Y=0.495
+ $X2=6.305 $Y2=0.495
r174 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.1
+ $Y=1.03 $X2=7.1 $Y2=1.03
r175 67 69 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.1 $Y=1.365
+ $X2=7.1 $Y2=1.03
r176 66 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.45
+ $X2=6.305 $Y2=1.45
r177 65 67 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.935 $Y=1.45
+ $X2=7.1 $Y2=1.365
r178 65 66 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.935 $Y=1.45
+ $X2=6.39 $Y2=1.45
r179 64 78 3.43356 $w=2.72e-07 $l=1.39155e-07 $layer=LI1_cond $X=6.305 $Y=1.715
+ $X2=6.202 $Y2=1.8
r180 63 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=1.535
+ $X2=6.305 $Y2=1.45
r181 63 64 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.305 $Y=1.535
+ $X2=6.305 $Y2=1.715
r182 62 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=1.365
+ $X2=6.305 $Y2=1.45
r183 61 75 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.305 $Y=0.685
+ $X2=6.305 $Y2=0.495
r184 61 62 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.305 $Y=0.685
+ $X2=6.305 $Y2=1.365
r185 57 78 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=6.202 $Y=1.885
+ $X2=6.202 $Y2=1.8
r186 57 59 24.7391 $w=3.73e-07 $l=8.05e-07 $layer=LI1_cond $X=6.202 $Y=1.885
+ $X2=6.202 $Y2=2.69
r187 55 78 3.08518 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=6.015 $Y=1.8
+ $X2=6.202 $Y2=1.8
r188 55 56 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.015 $Y=1.8
+ $X2=5.47 $Y2=1.8
r189 53 83 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.51
+ $X2=5.305 $Y2=1.675
r190 53 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.51
+ $X2=5.305 $Y2=1.345
r191 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.305
+ $Y=1.51 $X2=5.305 $Y2=1.51
r192 50 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.305 $Y=1.715
+ $X2=5.47 $Y2=1.8
r193 50 52 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.305 $Y=1.715
+ $X2=5.305 $Y2=1.51
r194 44 70 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.1 $Y=1.37 $X2=7.1
+ $Y2=1.03
r195 44 45 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.1 $Y=1.37
+ $X2=7.1 $Y2=1.535
r196 42 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.1 $Y=1.015
+ $X2=7.1 $Y2=1.03
r197 42 43 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.1 $Y=0.94 $X2=7.44
+ $Y2=0.94
r198 39 42 10.2553 $w=1.5e-07 $l=2e-08 $layer=POLY_cond $X=7.08 $Y=0.94 $X2=7.1
+ $Y2=0.94
r199 36 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.79 $Y=0.865
+ $X2=8.79 $Y2=0.94
r200 36 38 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.79 $Y=0.865
+ $X2=8.79 $Y2=0.58
r201 32 48 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=8.74 $Y=0.94 $X2=8.79
+ $Y2=0.94
r202 32 46 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=8.74 $Y=0.94
+ $X2=8.43 $Y2=0.94
r203 32 34 336.655 $w=2.5e-07 $l=1.355e-06 $layer=POLY_cond $X=8.74 $Y=1.015
+ $X2=8.74 $Y2=2.37
r204 29 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.43 $Y=0.865
+ $X2=8.43 $Y2=0.94
r205 29 31 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.43 $Y=0.865
+ $X2=8.43 $Y2=0.58
r206 28 43 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.515 $Y=0.94
+ $X2=7.44 $Y2=0.94
r207 27 46 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.355 $Y=0.94
+ $X2=8.43 $Y2=0.94
r208 27 28 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.355 $Y=0.94
+ $X2=7.515 $Y2=0.94
r209 23 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.44 $Y=0.865
+ $X2=7.44 $Y2=0.94
r210 23 25 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.44 $Y=0.865
+ $X2=7.44 $Y2=0.455
r211 19 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.08 $Y=0.865
+ $X2=7.08 $Y2=0.94
r212 19 21 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.08 $Y=0.865
+ $X2=7.08 $Y2=0.455
r213 17 45 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=7.06 $Y=2.235
+ $X2=7.06 $Y2=1.535
r214 13 83 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.265 $Y=2.335
+ $X2=5.265 $Y2=1.675
r215 9 82 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.215 $Y=0.455
+ $X2=5.215 $Y2=1.345
r216 2 78 300 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_PDIFF $count=2 $X=5.96
+ $Y=1.835 $X2=6.18 $Y2=1.88
r217 2 59 600 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=5.96
+ $Y=1.835 $X2=6.18 $Y2=2.69
r218 1 73 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.93
+ $Y=0.245 $X2=6.075 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%A_778_49# 1 2 9 11 12 15 19 22 26 29 30 31
+ 34 39 41 42
c100 41 0 2.33725e-19 $X=5.875 $Y=1.03
c101 19 0 1.86549e-19 $X=5.875 $Y=1.535
r102 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.875
+ $Y=1.03 $X2=5.875 $Y2=1.03
r103 38 39 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=0.475
+ $X2=4.55 $Y2=0.475
r104 35 38 2.19513 $w=4.18e-07 $l=8e-08 $layer=LI1_cond $X=4.305 $Y=0.475
+ $X2=4.385 $Y2=0.475
r105 30 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=0.95
+ $X2=5.875 $Y2=0.95
r106 30 31 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.71 $Y=0.95
+ $X2=5.25 $Y2=0.95
r107 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.165 $Y=0.865
+ $X2=5.25 $Y2=0.95
r108 28 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.165 $Y=0.685
+ $X2=5.165 $Y2=0.865
r109 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.08 $Y=0.6
+ $X2=5.165 $Y2=0.685
r110 26 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.08 $Y=0.6
+ $X2=4.55 $Y2=0.6
r111 24 35 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=4.305 $Y=0.685
+ $X2=4.305 $Y2=0.475
r112 24 34 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=4.305 $Y=0.685
+ $X2=4.305 $Y2=1.815
r113 22 34 7.56219 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=1.98
+ $X2=4.345 $Y2=1.815
r114 18 42 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.875 $Y=1.37
+ $X2=5.875 $Y2=1.03
r115 18 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.875 $Y=1.37
+ $X2=5.875 $Y2=1.535
r116 17 42 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.875 $Y=1.015
+ $X2=5.875 $Y2=1.03
r117 13 15 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=6.29 $Y=0.865
+ $X2=6.29 $Y2=0.455
r118 12 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.04 $Y=0.94
+ $X2=5.875 $Y2=1.015
r119 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.215 $Y=0.94
+ $X2=6.29 $Y2=0.865
r120 11 12 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.215 $Y=0.94
+ $X2=6.04 $Y2=0.94
r121 9 19 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=5.835 $Y=2.335
+ $X2=5.835 $Y2=1.535
r122 2 22 300 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.835 $X2=4.345 $Y2=1.98
r123 1 38 182 $w=1.7e-07 $l=5.99062e-07 $layer=licon1_NDIFF $count=1 $X=3.89
+ $Y=0.245 $X2=4.385 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%RESET_B 4 7 9 10 12 14 16 17 18 19 24
c51 17 0 3.63555e-19 $X=7.92 $Y=2.035
c52 16 0 3.19502e-20 $X=7.96 $Y=2.89
c53 14 0 1.53358e-19 $X=6.562 $Y=1.525
c54 7 0 8.03672e-20 $X=6.65 $Y=0.455
c55 4 0 1.0017e-19 $X=6.525 $Y=2.235
r56 18 19 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=7.96 $Y=2.385
+ $X2=7.96 $Y2=2.775
r57 18 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.96
+ $Y=2.385 $X2=7.96 $Y2=2.385
r58 17 18 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=7.96 $Y=2.035
+ $X2=7.96 $Y2=2.385
r59 15 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.96 $Y=2.725
+ $X2=7.96 $Y2=2.385
r60 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.96 $Y=2.725
+ $X2=7.96 $Y2=2.89
r61 13 14 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.562 $Y=1.375
+ $X2=6.562 $Y2=1.525
r62 12 16 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=7.87 $Y=3.075
+ $X2=7.87 $Y2=2.89
r63 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.795 $Y=3.15
+ $X2=7.87 $Y2=3.075
r64 9 10 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=7.795 $Y=3.15
+ $X2=6.65 $Y2=3.15
r65 7 13 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=6.65 $Y=0.455
+ $X2=6.65 $Y2=1.375
r66 4 14 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.525 $Y=2.235
+ $X2=6.525 $Y2=1.525
r67 2 10 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=6.525 $Y=3.075
+ $X2=6.65 $Y2=3.15
r68 2 4 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.525 $Y=3.075
+ $X2=6.525 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%A_1614_74# 1 2 9 13 17 23 26 29 33 37 38 45
+ 46
r63 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.31
+ $Y=1.155 $X2=9.31 $Y2=1.155
r64 37 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=1.075
+ $X2=9.31 $Y2=1.075
r65 37 38 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=9.145 $Y=1.075
+ $X2=8.64 $Y2=1.075
r66 33 35 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.475 $Y=2.015
+ $X2=8.475 $Y2=2.725
r67 31 38 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.475 $Y=1.075
+ $X2=8.64 $Y2=1.075
r68 31 33 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=8.475 $Y=1.16
+ $X2=8.475 $Y2=2.015
r69 27 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.215 $Y=1.075
+ $X2=8.475 $Y2=1.075
r70 27 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=8.215 $Y=0.99
+ $X2=8.215 $Y2=0.58
r71 25 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.31 $Y=1.495
+ $X2=9.31 $Y2=1.155
r72 25 26 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.31 $Y=1.495
+ $X2=9.31 $Y2=1.66
r73 22 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.31 $Y=1.14
+ $X2=9.31 $Y2=1.155
r74 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.31 $Y=1.065
+ $X2=9.58 $Y2=1.065
r75 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.22 $Y=1.065 $X2=9.31
+ $Y2=1.065
r76 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.58 $Y=0.99
+ $X2=9.58 $Y2=1.065
r77 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.58 $Y=0.99
+ $X2=9.58 $Y2=0.58
r78 13 26 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=9.27 $Y=2.37
+ $X2=9.27 $Y2=1.66
r79 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.22 $Y=0.99 $X2=9.22
+ $Y2=1.065
r80 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.22 $Y=0.99 $X2=9.22
+ $Y2=0.58
r81 2 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.33
+ $Y=1.87 $X2=8.475 $Y2=2.725
r82 2 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.33
+ $Y=1.87 $X2=8.475 $Y2=2.015
r83 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.07
+ $Y=0.37 $X2=8.215 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%VPWR 1 2 3 4 5 18 22 26 30 36 41 42 44 45
+ 46 52 59 71 77 78 81 84 87
c107 78 0 3.19502e-20 $X=9.84 $Y=3.33
r108 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r109 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r111 78 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r112 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r113 75 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.17 $Y=3.33
+ $X2=9.005 $Y2=3.33
r114 75 77 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.17 $Y=3.33
+ $X2=9.84 $Y2=3.33
r115 74 88 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 71 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.84 $Y=3.33
+ $X2=9.005 $Y2=3.33
r118 71 73 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=8.84 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 70 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r120 70 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 67 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=3.33
+ $X2=5.53 $Y2=3.33
r123 67 69 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=5.695 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r126 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r127 60 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=3.33
+ $X2=3.07 $Y2=3.33
r128 60 62 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.235 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 59 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=3.33
+ $X2=5.53 $Y2=3.33
r130 59 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.365 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 55 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 54 57 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 52 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=3.07 $Y2=3.33
r137 52 57 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 50 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 46 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r141 46 63 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r142 46 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r143 44 69 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.48 $Y2=3.33
r144 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.79 $Y2=3.33
r145 43 73 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.96 $Y2=3.33
r146 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.79 $Y2=3.33
r147 41 49 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.72 $Y2=3.33
r148 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.97 $Y2=3.33
r149 40 54 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=1.2 $Y2=3.33
r150 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.97 $Y2=3.33
r151 36 39 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.005 $Y=2.015
+ $X2=9.005 $Y2=2.725
r152 34 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=3.245
+ $X2=9.005 $Y2=3.33
r153 34 39 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=9.005 $Y=3.245
+ $X2=9.005 $Y2=2.725
r154 30 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.79 $Y=1.88
+ $X2=6.79 $Y2=2.59
r155 28 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.79 $Y=3.245
+ $X2=6.79 $Y2=3.33
r156 28 33 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=6.79 $Y=3.245
+ $X2=6.79 $Y2=2.59
r157 24 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=3.33
r158 24 26 35.4464 $w=3.28e-07 $l=1.015e-06 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=2.23
r159 20 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=3.245
+ $X2=3.07 $Y2=3.33
r160 20 22 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.07 $Y=3.245
+ $X2=3.07 $Y2=2.685
r161 16 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=3.245
+ $X2=0.97 $Y2=3.33
r162 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.97 $Y=3.245
+ $X2=0.97 $Y2=2.95
r163 5 39 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.865
+ $Y=1.87 $X2=9.005 $Y2=2.725
r164 5 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.865
+ $Y=1.87 $X2=9.005 $Y2=2.015
r165 4 33 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.65
+ $Y=1.735 $X2=6.79 $Y2=2.59
r166 4 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.65
+ $Y=1.735 $X2=6.79 $Y2=1.88
r167 3 26 300 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=2 $X=5.39
+ $Y=1.835 $X2=5.53 $Y2=2.23
r168 2 22 600 $w=1.7e-07 $l=1.11459e-06 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.675 $X2=3.07 $Y2=2.685
r169 1 18 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.83
+ $Y=2.095 $X2=0.97 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%Q 1 2 11 12 14 17 18 19
c35 17 0 1.0017e-19 $X=7.44 $Y=2.035
r36 19 28 4.86318 $w=4.53e-07 $l=1.85e-07 $layer=LI1_cond $X=7.387 $Y=2.775
+ $X2=7.387 $Y2=2.59
r37 18 28 4.86318 $w=4.53e-07 $l=1.85e-07 $layer=LI1_cond $X=7.387 $Y=2.405
+ $X2=7.387 $Y2=2.59
r38 17 18 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=7.387 $Y=2.035
+ $X2=7.387 $Y2=2.405
r39 14 16 9.9374 $w=3.73e-07 $l=2.1e-07 $layer=LI1_cond $X=7.632 $Y=0.475
+ $X2=7.632 $Y2=0.685
r40 12 16 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=7.53 $Y=1.715
+ $X2=7.53 $Y2=0.685
r41 11 12 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.387 $Y=1.88
+ $X2=7.387 $Y2=1.715
r42 9 17 2.44473 $w=4.53e-07 $l=9.3e-08 $layer=LI1_cond $X=7.387 $Y=1.942
+ $X2=7.387 $Y2=2.035
r43 9 11 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=7.387 $Y=1.942
+ $X2=7.387 $Y2=1.88
r44 2 28 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.185
+ $Y=1.735 $X2=7.325 $Y2=2.59
r45 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.185
+ $Y=1.735 $X2=7.325 $Y2=1.88
r46 1 14 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=7.515
+ $Y=0.245 $X2=7.655 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%Q_N 1 2 7 8 9 10 11 12 13 43
r22 43 44 7.82231 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=2.015
+ $X2=9.665 $Y2=1.85
r23 13 33 1.01363 $w=5.88e-07 $l=5e-08 $layer=LI1_cond $X=9.665 $Y=2.775
+ $X2=9.665 $Y2=2.725
r24 12 33 6.48721 $w=5.88e-07 $l=3.2e-07 $layer=LI1_cond $X=9.665 $Y=2.405
+ $X2=9.665 $Y2=2.725
r25 12 29 5.27085 $w=5.88e-07 $l=2.6e-07 $layer=LI1_cond $X=9.665 $Y=2.405
+ $X2=9.665 $Y2=2.145
r26 11 29 2.22998 $w=5.88e-07 $l=1.1e-07 $layer=LI1_cond $X=9.665 $Y=2.035
+ $X2=9.665 $Y2=2.145
r27 11 43 0.40545 $w=5.88e-07 $l=2e-08 $layer=LI1_cond $X=9.665 $Y=2.035
+ $X2=9.665 $Y2=2.015
r28 10 44 9.07242 $w=2.33e-07 $l=1.85e-07 $layer=LI1_cond $X=9.842 $Y=1.665
+ $X2=9.842 $Y2=1.85
r29 9 10 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=9.842 $Y=1.295
+ $X2=9.842 $Y2=1.665
r30 8 9 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=9.842 $Y=0.925
+ $X2=9.842 $Y2=1.295
r31 8 41 5.63961 $w=2.33e-07 $l=1.15e-07 $layer=LI1_cond $X=9.842 $Y=0.925
+ $X2=9.842 $Y2=0.81
r32 7 41 9.87681 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.795 $Y=0.555
+ $X2=9.795 $Y2=0.81
r33 2 43 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.395
+ $Y=1.87 $X2=9.535 $Y2=2.015
r34 2 33 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.395
+ $Y=1.87 $X2=9.535 $Y2=2.725
r35 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.655
+ $Y=0.37 $X2=9.795 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_LP%VGND 1 2 3 4 5 18 20 24 28 32 34 38 40 42
+ 47 55 62 63 66 69 72 75 78
r124 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r125 76 79 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r126 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r127 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r128 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r129 67 70 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r130 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r131 63 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=8.88
+ $Y2=0
r132 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r133 60 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.17 $Y=0 $X2=9.005
+ $Y2=0
r134 60 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.17 $Y=0 $X2=9.84
+ $Y2=0
r135 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r136 59 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=5.52
+ $Y2=0
r137 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r138 56 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=5.555
+ $Y2=0
r139 56 58 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=6.48
+ $Y2=0
r140 55 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.7 $Y=0 $X2=6.865
+ $Y2=0
r141 55 58 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.7 $Y=0 $X2=6.48
+ $Y2=0
r142 51 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r143 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r144 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r145 48 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.21
+ $Y2=0
r146 48 50 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.6
+ $Y2=0
r147 47 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.43 $Y=0 $X2=5.555
+ $Y2=0
r148 47 53 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.43 $Y=0 $X2=5.04
+ $Y2=0
r149 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r150 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r151 42 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r152 42 44 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r153 40 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r154 40 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r155 40 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r156 36 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=0.085
+ $X2=9.005 $Y2=0
r157 36 38 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.005 $Y=0.085
+ $X2=9.005 $Y2=0.58
r158 35 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.03 $Y=0 $X2=6.865
+ $Y2=0
r159 34 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=9.005
+ $Y2=0
r160 34 35 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=8.84 $Y=0 $X2=7.03
+ $Y2=0
r161 30 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=0.085
+ $X2=6.865 $Y2=0
r162 30 32 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.865 $Y=0.085
+ $X2=6.865 $Y2=0.455
r163 26 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.555 $Y=0.085
+ $X2=5.555 $Y2=0
r164 26 28 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=5.555 $Y=0.085
+ $X2=5.555 $Y2=0.455
r165 22 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r166 22 24 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.415
r167 21 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r168 20 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.21
+ $Y2=0
r169 20 21 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=3.045 $Y=0
+ $X2=1.235 $Y2=0
r170 16 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r171 16 18 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.77
r172 5 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.865
+ $Y=0.37 $X2=9.005 $Y2=0.58
r173 4 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.725
+ $Y=0.245 $X2=6.865 $Y2=0.455
r174 3 28 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.245 $X2=5.515 $Y2=0.455
r175 2 24 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.245 $X2=3.21 $Y2=0.415
r176 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.56 $X2=1.07 $Y2=0.77
.ends

