* File: sky130_fd_sc_lp__sleep_pargate_plv_7.spice
* Created: Fri Aug 28 11:32:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sleep_pargate_plv_7.pex.spice"
.subckt sky130_fd_sc_lp__sleep_pargate_plv_7  VPB SLEEP VPWR VIRTPWR
* 
* VIRTPWR	VIRTPWR
* VPWR	VPWR
* SLEEP	SLEEP
* VPB	VPB
MM1000 N_VIRTPWR_M1000_d N_SLEEP_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=7
+ AD=1.855 AS=1.855 PD=14.53 PS=14.53 NRD=0 NRS=0 M=1 R=46.6667 SA=75000.2
+ SB=75000.2 A=1.05 P=14.3 MULT=1
DX1_noxref noxref_1 VPB NWDIODE A=17.7175 P=22.73
c_29 VPB 0 8.20372e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sleep_pargate_plv_7.pxi.spice"
*
.ends
*
*
