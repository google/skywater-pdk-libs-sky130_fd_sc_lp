* File: sky130_fd_sc_lp__inv_0.pxi.spice
* Created: Wed Sep  2 09:55:32 2020
* 
x_PM_SKY130_FD_SC_LP__INV_0%A N_A_M1000_g N_A_M1001_g A A A N_A_c_20_n
+ N_A_c_21_n PM_SKY130_FD_SC_LP__INV_0%A
x_PM_SKY130_FD_SC_LP__INV_0%VPWR N_VPWR_M1001_s N_VPWR_c_37_n N_VPWR_c_38_n VPWR
+ N_VPWR_c_39_n N_VPWR_c_36_n PM_SKY130_FD_SC_LP__INV_0%VPWR
x_PM_SKY130_FD_SC_LP__INV_0%Y N_Y_M1000_d N_Y_M1001_d Y Y Y Y Y Y N_Y_c_49_n
+ PM_SKY130_FD_SC_LP__INV_0%Y
x_PM_SKY130_FD_SC_LP__INV_0%VGND N_VGND_M1000_s N_VGND_c_58_n N_VGND_c_59_n VGND
+ N_VGND_c_60_n N_VGND_c_61_n PM_SKY130_FD_SC_LP__INV_0%VGND
cc_1 VNB N_A_M1000_g 0.031511f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.56
cc_2 VNB N_A_M1001_g 0.00168831f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.63
cc_3 VNB N_A_c_20_n 0.0852989f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_4 VNB N_A_c_21_n 0.0299547f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_5 VNB N_VPWR_c_36_n 0.0442671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_Y_c_49_n 0.0631531f $X=-0.19 $Y=-0.245 $X2=0.242 $Y2=1.12
cc_7 VNB N_VGND_c_58_n 0.0112246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_VGND_c_59_n 0.02641f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.63
cc_9 VNB N_VGND_c_60_n 0.0177966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_61_n 0.0909177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VPB N_A_M1001_g 0.0568781f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.63
cc_12 VPB N_A_c_21_n 0.0271461f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_13 VPB N_VPWR_c_37_n 0.0111987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_14 VPB N_VPWR_c_38_n 0.0414032f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.63
cc_15 VPB N_VPWR_c_39_n 0.0176425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_16 VPB N_VPWR_c_36_n 0.0492901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_17 VPB N_Y_c_49_n 0.0644325f $X=-0.19 $Y=1.655 $X2=0.242 $Y2=1.12
cc_18 N_A_M1001_g N_VPWR_c_38_n 0.00573149f $X=0.485 $Y=2.63 $X2=0 $Y2=0
cc_19 N_A_c_20_n N_VPWR_c_38_n 8.68804e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_20 N_A_c_21_n N_VPWR_c_38_n 0.0274534f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_21 N_A_M1001_g N_VPWR_c_39_n 0.00570944f $X=0.485 $Y=2.63 $X2=0 $Y2=0
cc_22 N_A_M1001_g N_VPWR_c_36_n 0.00542671f $X=0.485 $Y=2.63 $X2=0 $Y2=0
cc_23 N_A_M1000_g N_Y_c_49_n 0.0481293f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_24 N_A_c_21_n N_Y_c_49_n 0.0933055f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_25 N_A_M1000_g N_VGND_c_59_n 0.00578496f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_26 N_A_c_20_n N_VGND_c_59_n 0.00204967f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_27 N_A_c_21_n N_VGND_c_59_n 0.0186726f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_28 N_A_M1000_g N_VGND_c_60_n 0.00478016f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_29 N_A_M1000_g N_VGND_c_61_n 0.00971575f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_30 N_VPWR_c_38_n N_Y_c_49_n 0.00311658f $X=0.27 $Y=2.455 $X2=0 $Y2=0
cc_31 N_VPWR_c_39_n N_Y_c_49_n 0.0129982f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_32 N_VPWR_c_36_n N_Y_c_49_n 0.0111232f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_33 N_Y_c_49_n N_VGND_c_60_n 0.0103721f $X=0.7 $Y=0.56 $X2=0 $Y2=0
cc_34 N_Y_c_49_n N_VGND_c_61_n 0.0108819f $X=0.7 $Y=0.56 $X2=0 $Y2=0
