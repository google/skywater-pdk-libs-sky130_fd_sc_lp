* File: sky130_fd_sc_lp__o21bai_4.pex.spice
* Created: Fri Aug 28 11:06:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BAI_4%B1_N 3 5 7 9 13
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.51 $X2=0.385 $Y2=1.51
r31 9 13 4.52224 $w=3.93e-07 $l=1.55e-07 $layer=LI1_cond $X=0.352 $Y=1.665
+ $X2=0.352 $Y2=1.51
r32 5 12 38.9103 $w=3.6e-07 $l=2.1609e-07 $layer=POLY_cond $X=0.53 $Y=1.675
+ $X2=0.412 $Y2=1.51
r33 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.53 $Y=1.675 $X2=0.53
+ $Y2=2.465
r34 1 12 38.9103 $w=3.6e-07 $l=1.93959e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.412 $Y2=1.51
r35 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%A_27_49# 1 2 9 11 13 16 18 20 23 25 27 30
+ 32 34 37 39 41 43 44 45 48 49 54 56 61 67 75
c126 67 0 1.7643e-19 $X=1.355 $Y=1.525
c127 32 0 7.6897e-20 $X=2.72 $Y=1.725
c128 18 0 1.39677e-19 $X=1.86 $Y=1.725
r129 74 75 59.7865 $w=4e-07 $l=4.3e-07 $layer=POLY_cond $X=2.29 $Y=1.525
+ $X2=2.72 $Y2=1.525
r130 71 72 59.7865 $w=4e-07 $l=4.3e-07 $layer=POLY_cond $X=1.43 $Y=1.525
+ $X2=1.86 $Y2=1.525
r131 67 71 10.4279 $w=4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.355 $Y=1.525
+ $X2=1.43 $Y2=1.525
r132 66 67 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=1.32 $Y=1.525
+ $X2=1.355 $Y2=1.525
r133 65 66 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.32
+ $Y=1.49 $X2=1.32 $Y2=1.49
r134 57 74 40.3212 $w=4e-07 $l=2.9e-07 $layer=POLY_cond $X=2 $Y=1.525 $X2=2.29
+ $Y2=1.525
r135 57 72 19.4654 $w=4e-07 $l=1.4e-07 $layer=POLY_cond $X=2 $Y=1.525 $X2=1.86
+ $Y2=1.525
r136 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2
+ $Y=1.49 $X2=2 $Y2=1.49
r137 54 65 3.24197 $w=3.16e-07 $l=6.9282e-08 $layer=LI1_cond $X=1.38 $Y=1.47
+ $X2=1.32 $Y2=1.49
r138 54 56 31.0659 $w=2.28e-07 $l=6.2e-07 $layer=LI1_cond $X=1.38 $Y=1.47 $X2=2
+ $Y2=1.47
r139 53 66 47.2731 $w=4e-07 $l=3.4e-07 $layer=POLY_cond $X=0.98 $Y=1.525
+ $X2=1.32 $Y2=1.525
r140 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.49 $X2=0.98 $Y2=1.49
r141 50 61 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.845 $Y=1.49
+ $X2=0.845 $Y2=1.16
r142 50 52 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.93 $Y=1.49 $X2=0.98
+ $Y2=1.49
r143 49 65 5.36061 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=1.175 $Y=1.49
+ $X2=1.32 $Y2=1.49
r144 49 52 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.175 $Y=1.49
+ $X2=0.98 $Y2=1.49
r145 47 50 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.655
+ $X2=0.845 $Y2=1.49
r146 47 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.845 $Y=1.655
+ $X2=0.845 $Y2=1.93
r147 46 60 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.445 $Y=2.015
+ $X2=0.297 $Y2=2.015
r148 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=2.015
+ $X2=0.845 $Y2=1.93
r149 45 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.76 $Y=2.015
+ $X2=0.445 $Y2=2.015
r150 43 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=1.16
+ $X2=0.845 $Y2=1.16
r151 43 44 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.76 $Y=1.16
+ $X2=0.355 $Y2=1.16
r152 39 60 2.72785 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=2.1
+ $X2=0.297 $Y2=2.015
r153 39 41 31.6434 $w=2.93e-07 $l=8.1e-07 $layer=LI1_cond $X=0.297 $Y=2.1
+ $X2=0.297 $Y2=2.91
r154 35 44 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.355 $Y2=1.16
r155 35 37 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.225 $Y2=0.42
r156 32 75 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.72 $Y=1.725
+ $X2=2.72 $Y2=1.525
r157 32 34 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.72 $Y=1.725
+ $X2=2.72 $Y2=2.465
r158 28 75 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.72 $Y=1.325
+ $X2=2.72 $Y2=1.525
r159 28 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.72 $Y=1.325
+ $X2=2.72 $Y2=0.665
r160 25 74 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.29 $Y=1.725
+ $X2=2.29 $Y2=1.525
r161 25 27 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.29 $Y=1.725
+ $X2=2.29 $Y2=2.465
r162 21 74 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.29 $Y=1.325
+ $X2=2.29 $Y2=1.525
r163 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.29 $Y=1.325
+ $X2=2.29 $Y2=0.665
r164 18 72 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.86 $Y=1.725
+ $X2=1.86 $Y2=1.525
r165 18 20 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.86 $Y=1.725
+ $X2=1.86 $Y2=2.465
r166 14 72 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.86 $Y=1.325
+ $X2=1.86 $Y2=1.525
r167 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.86 $Y=1.325
+ $X2=1.86 $Y2=0.665
r168 11 71 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.43 $Y=1.725
+ $X2=1.43 $Y2=1.525
r169 11 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.43 $Y=1.725
+ $X2=1.43 $Y2=2.465
r170 7 71 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.43 $Y=1.325 $X2=1.43
+ $Y2=1.525
r171 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.43 $Y2=0.665
r172 2 60 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.835 $X2=0.315 $Y2=2.095
r173 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.835 $X2=0.315 $Y2=2.91
r174 1 37 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%A1 3 7 11 15 19 23 27 31 35 36 38 39 41 42
+ 43 44 65
c121 39 0 1.36343e-19 $X=3.335 $Y=2.015
c122 36 0 1.46082e-19 $X=3.17 $Y=1.51
c123 7 0 8.90405e-20 $X=3.205 $Y=0.665
c124 3 0 2.4715e-19 $X=3.19 $Y=2.465
r125 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.46 $X2=6.45 $Y2=1.46
r126 63 65 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=6.215 $Y=1.46
+ $X2=6.45 $Y2=1.46
r127 62 63 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.2 $Y=1.46
+ $X2=6.215 $Y2=1.46
r128 61 66 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=6.11 $Y=1.567
+ $X2=6.45 $Y2=1.567
r129 60 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.11 $Y=1.46 $X2=6.2
+ $Y2=1.46
r130 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.46 $X2=6.11 $Y2=1.46
r131 58 60 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=5.785 $Y=1.46
+ $X2=6.11 $Y2=1.46
r132 56 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.77 $Y=1.46
+ $X2=5.785 $Y2=1.46
r133 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.77
+ $Y=1.46 $X2=5.77 $Y2=1.46
r134 54 56 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=5.355 $Y=1.46
+ $X2=5.77 $Y2=1.46
r135 52 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.34 $Y=1.46
+ $X2=5.355 $Y2=1.46
r136 44 66 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=6.48 $Y=1.567
+ $X2=6.45 $Y2=1.567
r137 43 61 3.29269 $w=3.83e-07 $l=1.1e-07 $layer=LI1_cond $X=6 $Y=1.567 $X2=6.11
+ $Y2=1.567
r138 43 57 6.88472 $w=3.83e-07 $l=2.3e-07 $layer=LI1_cond $X=6 $Y=1.567 $X2=5.77
+ $Y2=1.567
r139 42 57 7.4834 $w=3.83e-07 $l=2.5e-07 $layer=LI1_cond $X=5.52 $Y=1.567
+ $X2=5.77 $Y2=1.567
r140 40 42 9.6854 $w=5.55e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.35 $Y=1.76
+ $X2=5.435 $Y2=1.665
r141 40 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.35 $Y=1.76
+ $X2=5.35 $Y2=1.93
r142 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.265 $Y=2.015
+ $X2=5.35 $Y2=1.93
r143 38 39 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=5.265 $Y=2.015
+ $X2=3.335 $Y2=2.015
r144 36 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.51
+ $X2=3.17 $Y2=1.675
r145 36 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.51
+ $X2=3.17 $Y2=1.345
r146 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.51 $X2=3.17 $Y2=1.51
r147 33 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.17 $Y=1.93
+ $X2=3.335 $Y2=2.015
r148 33 35 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.17 $Y=1.93
+ $X2=3.17 $Y2=1.51
r149 29 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.215 $Y=1.295
+ $X2=6.215 $Y2=1.46
r150 29 31 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=6.215 $Y=1.295
+ $X2=6.215 $Y2=0.665
r151 25 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.2 $Y=1.625
+ $X2=6.2 $Y2=1.46
r152 25 27 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.2 $Y=1.625
+ $X2=6.2 $Y2=2.465
r153 21 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.785 $Y=1.295
+ $X2=5.785 $Y2=1.46
r154 21 23 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=5.785 $Y=1.295
+ $X2=5.785 $Y2=0.665
r155 17 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.77 $Y=1.625
+ $X2=5.77 $Y2=1.46
r156 17 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.77 $Y=1.625
+ $X2=5.77 $Y2=2.465
r157 13 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.355 $Y=1.295
+ $X2=5.355 $Y2=1.46
r158 13 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=5.355 $Y=1.295
+ $X2=5.355 $Y2=0.665
r159 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.34 $Y=1.625
+ $X2=5.34 $Y2=1.46
r160 9 11 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.34 $Y=1.625
+ $X2=5.34 $Y2=2.465
r161 7 50 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.205 $Y=0.665
+ $X2=3.205 $Y2=1.345
r162 3 51 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.19 $Y=2.465
+ $X2=3.19 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%A2 3 7 11 15 19 23 27 31 33 34 35 53 54
c83 54 0 7.96714e-20 $X=4.91 $Y=1.51
r84 54 55 2.21779 $w=3.26e-07 $l=1.5e-08 $layer=POLY_cond $X=4.91 $Y=1.51
+ $X2=4.925 $Y2=1.51
r85 52 54 24.3957 $w=3.26e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.51
+ $X2=4.91 $Y2=1.51
r86 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.745
+ $Y=1.51 $X2=4.745 $Y2=1.51
r87 50 52 36.9632 $w=3.26e-07 $l=2.5e-07 $layer=POLY_cond $X=4.495 $Y=1.51
+ $X2=4.745 $Y2=1.51
r88 49 50 2.21779 $w=3.26e-07 $l=1.5e-08 $layer=POLY_cond $X=4.48 $Y=1.51
+ $X2=4.495 $Y2=1.51
r89 47 49 11.089 $w=3.26e-07 $l=7.5e-08 $layer=POLY_cond $X=4.405 $Y=1.51
+ $X2=4.48 $Y2=1.51
r90 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.405
+ $Y=1.51 $X2=4.405 $Y2=1.51
r91 45 47 50.2699 $w=3.26e-07 $l=3.4e-07 $layer=POLY_cond $X=4.065 $Y=1.51
+ $X2=4.405 $Y2=1.51
r92 44 45 2.21779 $w=3.26e-07 $l=1.5e-08 $layer=POLY_cond $X=4.05 $Y=1.51
+ $X2=4.065 $Y2=1.51
r93 42 44 48.0521 $w=3.26e-07 $l=3.25e-07 $layer=POLY_cond $X=3.725 $Y=1.51
+ $X2=4.05 $Y2=1.51
r94 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.725
+ $Y=1.51 $X2=3.725 $Y2=1.51
r95 40 42 13.3067 $w=3.26e-07 $l=9e-08 $layer=POLY_cond $X=3.635 $Y=1.51
+ $X2=3.725 $Y2=1.51
r96 39 40 2.21779 $w=3.26e-07 $l=1.5e-08 $layer=POLY_cond $X=3.62 $Y=1.51
+ $X2=3.635 $Y2=1.51
r97 35 53 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.745 $Y2=1.587
r98 35 48 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.405 $Y2=1.587
r99 34 48 11.5244 $w=3.23e-07 $l=3.25e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.405 $Y2=1.587
r100 34 43 12.5882 $w=3.23e-07 $l=3.55e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=3.725 $Y2=1.587
r101 33 43 4.43247 $w=3.23e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=1.587
+ $X2=3.725 $Y2=1.587
r102 29 55 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.925 $Y=1.345
+ $X2=4.925 $Y2=1.51
r103 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.925 $Y=1.345
+ $X2=4.925 $Y2=0.665
r104 25 54 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.91 $Y=1.675
+ $X2=4.91 $Y2=1.51
r105 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.91 $Y=1.675
+ $X2=4.91 $Y2=2.465
r106 21 50 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.495 $Y=1.345
+ $X2=4.495 $Y2=1.51
r107 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.495 $Y=1.345
+ $X2=4.495 $Y2=0.665
r108 17 49 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=1.675
+ $X2=4.48 $Y2=1.51
r109 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.48 $Y=1.675
+ $X2=4.48 $Y2=2.465
r110 13 45 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.065 $Y=1.345
+ $X2=4.065 $Y2=1.51
r111 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.065 $Y=1.345
+ $X2=4.065 $Y2=0.665
r112 9 44 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=1.675
+ $X2=4.05 $Y2=1.51
r113 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.05 $Y=1.675
+ $X2=4.05 $Y2=2.465
r114 5 40 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.635 $Y=1.345
+ $X2=3.635 $Y2=1.51
r115 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.635 $Y=1.345
+ $X2=3.635 $Y2=0.665
r116 1 39 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.62 $Y=1.675
+ $X2=3.62 $Y2=1.51
r117 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.62 $Y=1.675
+ $X2=3.62 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%VPWR 1 2 3 4 5 17 20 24 30 34 36 38 43 46
+ 47 49 50 51 53 65 72 78 81 85
r104 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 76 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r108 76 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r109 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r110 73 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.72 $Y=3.33
+ $X2=5.555 $Y2=3.33
r111 73 75 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.72 $Y=3.33 $X2=6
+ $Y2=3.33
r112 72 84 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=6.25 $Y=3.33
+ $X2=6.485 $Y2=3.33
r113 72 75 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=3.33 $X2=6
+ $Y2=3.33
r114 71 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r115 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 67 70 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 65 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.39 $Y=3.33
+ $X2=5.555 $Y2=3.33
r119 65 70 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.39 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 64 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r121 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r123 61 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 58 78 13.9156 $w=1.7e-07 $l=3.63e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=0.977 $Y2=3.33
r126 58 60 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 56 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r129 53 78 13.9156 $w=1.7e-07 $l=3.62e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.977 $Y2=3.33
r130 53 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 51 71 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 51 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r133 49 63 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 49 50 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.92 $Y2=3.33
r135 48 67 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.07 $Y=3.33 $X2=3.12
+ $Y2=3.33
r136 48 50 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=2.92 $Y2=3.33
r137 46 60 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=1.68 $Y2=3.33
r138 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=2.075 $Y2=3.33
r139 45 63 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.24 $Y=3.33 $X2=2.64
+ $Y2=3.33
r140 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=3.33
+ $X2=2.075 $Y2=3.33
r141 43 44 8.89246 $w=7.23e-07 $l=1.9e-07 $layer=LI1_cond $X=0.977 $Y=2.46
+ $X2=0.977 $Y2=2.27
r142 38 41 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=6.415 $Y=2.015
+ $X2=6.415 $Y2=2.95
r143 36 84 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.485 $Y2=3.33
r144 36 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.415 $Y2=2.95
r145 32 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.555 $Y=3.245
+ $X2=5.555 $Y2=3.33
r146 32 34 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.555 $Y=3.245
+ $X2=5.555 $Y2=2.765
r147 28 50 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=3.33
r148 28 30 14.5976 $w=2.98e-07 $l=3.8e-07 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=2.865
r149 24 27 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.075 $Y=2.19
+ $X2=2.075 $Y2=2.95
r150 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=3.33
r151 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=2.95
r152 20 44 13.4452 $w=2.38e-07 $l=2.8e-07 $layer=LI1_cond $X=1.22 $Y=1.99
+ $X2=1.22 $Y2=2.27
r153 17 78 2.93543 $w=7.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.977 $Y=3.245
+ $X2=0.977 $Y2=3.33
r154 16 43 2.83759 $w=7.23e-07 $l=1.72e-07 $layer=LI1_cond $X=0.977 $Y=2.632
+ $X2=0.977 $Y2=2.46
r155 16 17 10.113 $w=7.23e-07 $l=6.13e-07 $layer=LI1_cond $X=0.977 $Y=2.632
+ $X2=0.977 $Y2=3.245
r156 5 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.835 $X2=6.415 $Y2=2.95
r157 5 38 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.835 $X2=6.415 $Y2=2.015
r158 4 34 600 $w=1.7e-07 $l=9.97547e-07 $layer=licon1_PDIFF $count=1 $X=5.415
+ $Y=1.835 $X2=5.555 $Y2=2.765
r159 3 30 600 $w=1.7e-07 $l=1.10711e-06 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.835 $X2=2.955 $Y2=2.865
r160 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.835 $X2=2.075 $Y2=2.95
r161 2 24 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.835 $X2=2.075 $Y2=2.19
r162 1 43 150 $w=1.7e-07 $l=8.78564e-07 $layer=licon1_PDIFF $count=4 $X=0.605
+ $Y=1.835 $X2=1.215 $Y2=2.46
r163 1 20 600 $w=1.7e-07 $l=6.83118e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.835 $X2=1.215 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%Y 1 2 3 4 5 6 21 25 26 27 28 32 35 39 43 45
+ 46 47 48 49 50 54
c80 45 0 1.68735e-19 $X=2.53 $Y=1.84
c81 39 0 1.46082e-19 $X=3.57 $Y=2.445
c82 28 0 2.18092e-19 $X=2.53 $Y=1.755
c83 27 0 8.90405e-20 $X=2.53 $Y=1.185
r84 50 54 3.32574 $w=4.1e-07 $l=1.95e-07 $layer=LI1_cond $X=2.53 $Y=0.98
+ $X2=2.335 $Y2=0.98
r85 49 54 4.91896 $w=4.08e-07 $l=1.75e-07 $layer=LI1_cond $X=2.16 $Y=0.98
+ $X2=2.335 $Y2=0.98
r86 48 49 14.4758 $w=4.08e-07 $l=5.15e-07 $layer=LI1_cond $X=1.645 $Y=0.98
+ $X2=2.16 $Y2=0.98
r87 41 43 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=3.835 $Y=2.445
+ $X2=4.695 $Y2=2.445
r88 39 47 12.2291 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.57 $Y=2.445
+ $X2=3.24 $Y2=2.445
r89 39 41 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.57 $Y=2.445
+ $X2=3.835 $Y2=2.445
r90 38 46 1.37842 $w=2.5e-07 $l=1.58e-07 $layer=LI1_cond $X=2.725 $Y=2.405
+ $X2=2.567 $Y2=2.405
r91 38 47 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=2.725 $Y=2.405
+ $X2=3.24 $Y2=2.405
r92 33 46 5.12339 $w=2.52e-07 $l=1.52889e-07 $layer=LI1_cond $X=2.505 $Y=2.53
+ $X2=2.567 $Y2=2.405
r93 33 35 22.1818 $w=1.88e-07 $l=3.8e-07 $layer=LI1_cond $X=2.505 $Y=2.53
+ $X2=2.505 $Y2=2.91
r94 30 46 5.12339 $w=2.52e-07 $l=1.25e-07 $layer=LI1_cond $X=2.567 $Y=2.28
+ $X2=2.567 $Y2=2.405
r95 30 32 10.9756 $w=3.13e-07 $l=3e-07 $layer=LI1_cond $X=2.567 $Y=2.28
+ $X2=2.567 $Y2=1.98
r96 29 45 2.71818 $w=3.52e-07 $l=1.01833e-07 $layer=LI1_cond $X=2.567 $Y=1.925
+ $X2=2.53 $Y2=1.84
r97 29 32 2.0122 $w=3.13e-07 $l=5.5e-08 $layer=LI1_cond $X=2.567 $Y=1.925
+ $X2=2.567 $Y2=1.98
r98 28 45 2.71818 $w=3.52e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.755
+ $X2=2.53 $Y2=1.84
r99 27 50 3.49629 $w=3.9e-07 $l=2.05e-07 $layer=LI1_cond $X=2.53 $Y=1.185
+ $X2=2.53 $Y2=0.98
r100 27 28 16.8434 $w=3.88e-07 $l=5.7e-07 $layer=LI1_cond $X=2.53 $Y=1.185
+ $X2=2.53 $Y2=1.755
r101 25 45 4.06059 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.335 $Y=1.84
+ $X2=2.53 $Y2=1.84
r102 25 26 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.335 $Y=1.84
+ $X2=1.74 $Y2=1.84
r103 21 23 46.5988 $w=2.28e-07 $l=9.3e-07 $layer=LI1_cond $X=1.625 $Y=1.98
+ $X2=1.625 $Y2=2.91
r104 19 26 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.625 $Y=1.925
+ $X2=1.74 $Y2=1.84
r105 19 21 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.625 $Y=1.925
+ $X2=1.625 $Y2=1.98
r106 6 43 600 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=1 $X=4.555
+ $Y=1.835 $X2=4.695 $Y2=2.445
r107 5 41 600 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=1 $X=3.695
+ $Y=1.835 $X2=3.835 $Y2=2.445
r108 4 35 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=1.835 $X2=2.505 $Y2=2.91
r109 4 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.835 $X2=2.505 $Y2=1.98
r110 3 23 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.835 $X2=1.645 $Y2=2.91
r111 3 21 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.835 $X2=1.645 $Y2=1.98
r112 2 50 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.245 $X2=2.505 $Y2=0.94
r113 1 48 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.245 $X2=1.645 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%A_653_367# 1 2 3 4 13 19 20 21 25 29
c37 13 0 7.6897e-20 $X=4.96 $Y=2.932
c38 1 0 1.36343e-19 $X=3.265 $Y=1.835
r39 27 35 5.05528 $w=1.95e-07 $l=9.74679e-08 $layer=LI1_cond $X=5.985 $Y=2.46
+ $X2=5.98 $Y2=2.365
r40 27 29 1.16746 $w=1.88e-07 $l=2e-08 $layer=LI1_cond $X=5.985 $Y=2.46
+ $X2=5.985 $Y2=2.48
r41 23 35 5.05528 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=5.98 $Y=2.27
+ $X2=5.98 $Y2=2.365
r42 23 25 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=5.98 $Y=2.27
+ $X2=5.98 $Y2=2.095
r43 22 32 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=5.22 $Y=2.365
+ $X2=5.09 $Y2=2.365
r44 21 35 1.43626 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=5.88 $Y=2.365 $X2=5.98
+ $Y2=2.365
r45 21 22 38.5263 $w=1.88e-07 $l=6.6e-07 $layer=LI1_cond $X=5.88 $Y=2.365
+ $X2=5.22 $Y2=2.365
r46 20 34 3.56836 $w=2.6e-07 $l=1.42e-07 $layer=LI1_cond $X=5.09 $Y=2.79
+ $X2=5.09 $Y2=2.932
r47 19 32 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=5.09 $Y=2.46 $X2=5.09
+ $Y2=2.365
r48 19 20 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=5.09 $Y=2.46
+ $X2=5.09 $Y2=2.79
r49 15 18 34.7755 $w=2.83e-07 $l=8.6e-07 $layer=LI1_cond $X=3.405 $Y=2.932
+ $X2=4.265 $Y2=2.932
r50 13 34 3.26681 $w=2.85e-07 $l=1.3e-07 $layer=LI1_cond $X=4.96 $Y=2.932
+ $X2=5.09 $Y2=2.932
r51 13 18 28.1034 $w=2.83e-07 $l=6.95e-07 $layer=LI1_cond $X=4.96 $Y=2.932
+ $X2=4.265 $Y2=2.932
r52 4 29 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=5.845
+ $Y=1.835 $X2=5.985 $Y2=2.48
r53 4 25 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.835 $X2=5.985 $Y2=2.095
r54 3 34 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=1.835 $X2=5.125 $Y2=2.91
r55 3 32 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=1.835 $X2=5.125 $Y2=2.37
r56 2 18 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=1.835 $X2=4.265 $Y2=2.895
r57 1 15 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.835 $X2=3.405 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%VGND 1 2 3 4 5 18 22 26 28 32 36 39 40 41
+ 42 43 45 60 67 68 71 74 77
c99 18 0 1.7643e-19 $X=0.69 $Y=0.39
r100 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r101 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r103 68 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r104 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r105 65 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=0 $X2=6
+ $Y2=0
r106 65 67 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.165 $Y=0
+ $X2=6.48 $Y2=0
r107 64 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r108 64 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r109 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r110 61 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.305 $Y=0 $X2=5.14
+ $Y2=0
r111 61 63 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.305 $Y=0
+ $X2=5.52 $Y2=0
r112 60 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=0 $X2=6
+ $Y2=0
r113 60 63 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=0
+ $X2=5.52 $Y2=0
r114 59 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r115 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r116 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r117 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r118 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r119 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r120 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 50 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r122 50 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r123 48 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r124 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r125 45 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r126 45 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r127 43 59 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r128 43 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r129 41 58 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.08
+ $Y2=0
r130 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.28
+ $Y2=0
r131 39 55 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0
+ $X2=3.12 $Y2=0
r132 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r133 38 58 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.585 $Y=0
+ $X2=4.08 $Y2=0
r134 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r135 34 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6 $Y=0.085 $X2=6
+ $Y2=0
r136 34 36 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6 $Y=0.085 $X2=6
+ $Y2=0.39
r137 30 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.085
+ $X2=5.14 $Y2=0
r138 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.14 $Y=0.085
+ $X2=5.14 $Y2=0.39
r139 29 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.28
+ $Y2=0
r140 28 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=0 $X2=5.14
+ $Y2=0
r141 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=4.445 $Y2=0
r142 24 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0
r143 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0.39
r144 20 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r145 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.37
r146 16 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r147 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.39
r148 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.86
+ $Y=0.245 $X2=6 $Y2=0.39
r149 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5
+ $Y=0.245 $X2=5.14 $Y2=0.39
r150 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.245 $X2=4.28 $Y2=0.39
r151 2 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.28
+ $Y=0.245 $X2=3.42 $Y2=0.37
r152 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.245 $X2=0.69 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_4%A_218_49# 1 2 3 4 5 6 7 24 28 31 32 33 36
+ 38 42 44 48 50 54 57 60 61 62
c88 32 0 7.96714e-20 $X=3.755 $Y=1.14
r89 52 54 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=6.465 $Y=1.035
+ $X2=6.465 $Y2=0.42
r90 51 62 5.40251 $w=1.8e-07 $l=9.98749e-08 $layer=LI1_cond $X=5.665 $Y=1.12
+ $X2=5.57 $Y2=1.11
r91 50 52 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.335 $Y=1.12
+ $X2=6.465 $Y2=1.035
r92 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.335 $Y=1.12
+ $X2=5.665 $Y2=1.12
r93 46 62 1.14861 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=5.57 $Y=1.015
+ $X2=5.57 $Y2=1.11
r94 46 48 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=5.57 $Y=1.015
+ $X2=5.57 $Y2=0.42
r95 45 61 5.40251 $w=1.8e-07 $l=2.32702e-07 $layer=LI1_cond $X=4.805 $Y=1.11
+ $X2=4.615 $Y2=1.015
r96 44 62 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.475 $Y=1.11
+ $X2=5.57 $Y2=1.11
r97 44 45 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=5.475 $Y=1.11
+ $X2=4.805 $Y2=1.11
r98 40 61 1.14861 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=4.71 $Y=1.015
+ $X2=4.615 $Y2=1.015
r99 40 42 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=4.71 $Y=1.015
+ $X2=4.71 $Y2=0.42
r100 39 60 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.945 $Y=1.14
+ $X2=3.85 $Y2=1.14
r101 38 61 5.40251 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.615 $Y=1.14
+ $X2=4.615 $Y2=1.015
r102 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.615 $Y=1.14
+ $X2=3.945 $Y2=1.14
r103 34 60 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=1.055
+ $X2=3.85 $Y2=1.14
r104 34 36 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=3.85 $Y=1.055
+ $X2=3.85 $Y2=0.42
r105 32 60 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.755 $Y=1.14
+ $X2=3.85 $Y2=1.14
r106 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.755 $Y=1.14
+ $X2=3.085 $Y2=1.14
r107 29 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.99 $Y=1.055
+ $X2=3.085 $Y2=1.14
r108 29 31 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=2.99 $Y=1.055
+ $X2=2.99 $Y2=0.94
r109 28 59 4.84456 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=2.99 $Y=0.595
+ $X2=2.99 $Y2=0.425
r110 28 31 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=2.99 $Y=0.595
+ $X2=2.99 $Y2=0.94
r111 25 57 3.35835 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=0.425
+ $X2=1.215 $Y2=0.425
r112 25 27 23.5573 $w=3.38e-07 $l=6.95e-07 $layer=LI1_cond $X=1.38 $Y=0.425
+ $X2=2.075 $Y2=0.425
r113 24 59 2.70725 $w=3.4e-07 $l=9.5e-08 $layer=LI1_cond $X=2.895 $Y=0.425
+ $X2=2.99 $Y2=0.425
r114 24 27 27.7942 $w=3.38e-07 $l=8.2e-07 $layer=LI1_cond $X=2.895 $Y=0.425
+ $X2=2.075 $Y2=0.425
r115 7 54 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=6.29
+ $Y=0.245 $X2=6.43 $Y2=0.42
r116 6 48 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=5.43
+ $Y=0.245 $X2=5.57 $Y2=0.42
r117 5 42 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.57
+ $Y=0.245 $X2=4.71 $Y2=0.42
r118 4 36 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.245 $X2=3.85 $Y2=0.42
r119 3 59 182 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.245 $X2=2.99 $Y2=0.42
r120 3 31 182 $w=1.7e-07 $l=7.86479e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.245 $X2=2.99 $Y2=0.94
r121 2 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.245 $X2=2.075 $Y2=0.43
r122 1 57 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.245 $X2=1.215 $Y2=0.39
.ends

