* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND D_N a_286_512# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Y a_286_512# a_463_355# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND a_45_164# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 Y a_45_164# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_718_355# B a_919_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_45_164# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_45_164# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND a_286_512# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Y a_286_512# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_919_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_718_355# a_45_164# a_463_355# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_919_367# B a_718_355# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VPWR D_N a_286_512# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_463_355# a_45_164# a_718_355# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR A a_919_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_463_355# a_286_512# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
