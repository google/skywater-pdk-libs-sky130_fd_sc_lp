* File: sky130_fd_sc_lp__a32o_m.pxi.spice
* Created: Fri Aug 28 10:01:23 2020
* 
x_PM_SKY130_FD_SC_LP__A32O_M%A_84_153# N_A_84_153#_M1007_d N_A_84_153#_M1002_d
+ N_A_84_153#_M1001_g N_A_84_153#_M1006_g N_A_84_153#_c_71_n N_A_84_153#_c_72_n
+ N_A_84_153#_c_73_n N_A_84_153#_c_100_p N_A_84_153#_c_74_n N_A_84_153#_c_75_n
+ N_A_84_153#_c_76_n N_A_84_153#_c_77_n N_A_84_153#_c_115_p N_A_84_153#_c_78_n
+ N_A_84_153#_c_79_n PM_SKY130_FD_SC_LP__A32O_M%A_84_153#
x_PM_SKY130_FD_SC_LP__A32O_M%A3 N_A3_M1003_g N_A3_M1004_g A3 N_A3_c_161_n
+ N_A3_c_162_n N_A3_c_163_n PM_SKY130_FD_SC_LP__A32O_M%A3
x_PM_SKY130_FD_SC_LP__A32O_M%A2 N_A2_M1000_g N_A2_M1011_g A2 A2 N_A2_c_199_n
+ N_A2_c_200_n PM_SKY130_FD_SC_LP__A32O_M%A2
x_PM_SKY130_FD_SC_LP__A32O_M%A1 N_A1_M1005_g N_A1_M1007_g N_A1_c_232_n
+ N_A1_c_233_n A1 N_A1_c_235_n N_A1_c_236_n PM_SKY130_FD_SC_LP__A32O_M%A1
x_PM_SKY130_FD_SC_LP__A32O_M%B1 N_B1_M1002_g N_B1_M1009_g N_B1_c_277_n B1 B1 B1
+ B1 B1 N_B1_c_280_n PM_SKY130_FD_SC_LP__A32O_M%B1
x_PM_SKY130_FD_SC_LP__A32O_M%B2 N_B2_c_328_n N_B2_M1008_g N_B2_M1010_g
+ N_B2_c_323_n N_B2_c_330_n N_B2_c_324_n N_B2_c_325_n B2 B2 B2 N_B2_c_327_n
+ PM_SKY130_FD_SC_LP__A32O_M%B2
x_PM_SKY130_FD_SC_LP__A32O_M%X N_X_M1001_s N_X_M1006_s N_X_c_360_n N_X_c_362_n X
+ PM_SKY130_FD_SC_LP__A32O_M%X
x_PM_SKY130_FD_SC_LP__A32O_M%VPWR N_VPWR_M1006_d N_VPWR_M1011_d N_VPWR_c_382_n
+ N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_399_p N_VPWR_c_377_n VPWR
+ N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_374_n N_VPWR_c_381_n
+ PM_SKY130_FD_SC_LP__A32O_M%VPWR
x_PM_SKY130_FD_SC_LP__A32O_M%A_228_385# N_A_228_385#_M1004_d
+ N_A_228_385#_M1005_d N_A_228_385#_M1008_d N_A_228_385#_c_402_n
+ N_A_228_385#_c_403_n N_A_228_385#_c_404_n N_A_228_385#_c_405_n
+ N_A_228_385#_c_430_n N_A_228_385#_c_406_n
+ PM_SKY130_FD_SC_LP__A32O_M%A_228_385#
x_PM_SKY130_FD_SC_LP__A32O_M%VGND N_VGND_M1001_d N_VGND_M1010_d N_VGND_c_438_n
+ N_VGND_c_439_n N_VGND_c_440_n VGND N_VGND_c_441_n N_VGND_c_442_n
+ N_VGND_c_443_n N_VGND_c_444_n PM_SKY130_FD_SC_LP__A32O_M%VGND
cc_1 VNB N_A_84_153#_c_71_n 0.0202506f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.765
cc_2 VNB N_A_84_153#_c_72_n 0.0103985f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.915
cc_3 VNB N_A_84_153#_c_73_n 0.0324272f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=1.42
cc_4 VNB N_A_84_153#_c_74_n 0.00510859f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.335
cc_5 VNB N_A_84_153#_c_75_n 0.00245088f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.945
cc_6 VNB N_A_84_153#_c_76_n 0.00215662f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.5
cc_7 VNB N_A_84_153#_c_77_n 0.0282793f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.5
cc_8 VNB N_A_84_153#_c_78_n 0.00122896f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.42
cc_9 VNB N_A_84_153#_c_79_n 0.0245269f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.335
cc_10 VNB N_A3_M1004_g 0.0288869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_c_161_n 0.0304693f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.445
cc_12 VNB N_A3_c_162_n 0.00601811f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.665
cc_13 VNB N_A3_c_163_n 0.0169103f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.135
cc_14 VNB N_A2_M1011_g 0.0286959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A2 0.00374272f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.335
cc_16 VNB N_A2_c_199_n 0.0307423f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.135
cc_17 VNB N_A2_c_200_n 0.0162464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1005_g 0.00893715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_232_n 0.0140224f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.445
cc_20 VNB N_A1_c_233_n 0.0100974f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.445
cc_21 VNB A1 0.00296158f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.665
cc_22 VNB N_A1_c_235_n 0.030147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_236_n 0.0184897f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.915
cc_24 VNB N_B1_M1002_g 0.0114264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_M1009_g 0.0422775f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.915
cc_26 VNB N_B1_c_277_n 0.0215797f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.445
cc_27 VNB N_B2_M1010_g 0.0266578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B2_c_323_n 0.0100904f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.765
cc_29 VNB N_B2_c_324_n 0.0311688f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.765
cc_30 VNB N_B2_c_325_n 0.0245005f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=1.42
cc_31 VNB B2 0.00741547f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.42
cc_32 VNB N_B2_c_327_n 0.0380056f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.505
cc_33 VNB N_X_c_360_n 0.0146279f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.765
cc_34 VNB X 0.0480799f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=1.42
cc_35 VNB N_VPWR_c_374_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=2.05
cc_36 VNB N_VGND_c_438_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.765
cc_37 VNB N_VGND_c_439_n 0.0109718f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.445
cc_38 VNB N_VGND_c_440_n 0.0127868f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.135
cc_39 VNB N_VGND_c_441_n 0.0174606f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.915
cc_40 VNB N_VGND_c_442_n 0.0557596f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=0.48
cc_41 VNB N_VGND_c_443_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.5
cc_42 VNB N_VGND_c_444_n 0.19078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A_84_153#_M1006_g 0.0318405f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.135
cc_44 VPB N_A_84_153#_c_75_n 0.00213533f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=1.945
cc_45 VPB N_A_84_153#_c_76_n 4.92577e-19 $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.5
cc_46 VPB N_A_84_153#_c_77_n 0.00730619f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.5
cc_47 VPB N_A3_M1004_g 0.024097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_M1011_g 0.0220217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A1_M1005_g 0.0236447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B1_M1002_g 0.0444455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB B1 0.0647f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.915
cc_52 VPB N_B1_c_280_n 0.0476351f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=0.585
cc_53 VPB N_B2_c_328_n 0.0200601f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=0.235
cc_54 VPB N_B2_c_323_n 6.30649e-19 $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.765
cc_55 VPB N_B2_c_330_n 0.0272738f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.665
cc_56 VPB B2 0.00714791f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.42
cc_57 VPB N_X_c_362_n 0.0192977f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.765
cc_58 VPB X 0.0129619f $X=-0.19 $Y=1.655 $X2=2.565 $Y2=1.42
cc_59 VPB N_VPWR_c_375_n 0.0468031f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.665
cc_60 VPB N_VPWR_c_376_n 0.0107433f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.135
cc_61 VPB N_VPWR_c_377_n 0.00122182f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.42
cc_62 VPB N_VPWR_c_378_n 0.0213956f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=0.48
cc_63 VPB N_VPWR_c_379_n 0.0634837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_374_n 0.0856674f $X=-0.19 $Y=1.655 $X2=2.57 $Y2=2.05
cc_65 VPB N_VPWR_c_381_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=2.05
cc_66 VPB N_A_228_385#_c_402_n 0.0106212f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.445
cc_67 VPB N_A_228_385#_c_403_n 0.00115793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_228_385#_c_404_n 0.0135623f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.765
cc_69 VPB N_A_228_385#_c_405_n 0.0028715f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.915
cc_70 VPB N_A_228_385#_c_406_n 0.00253089f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=0.48
cc_71 N_A_84_153#_M1006_g N_A3_M1004_g 0.0192266f $X=0.555 $Y=2.135 $X2=0 $Y2=0
cc_72 N_A_84_153#_c_73_n N_A3_M1004_g 0.014816f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_73 N_A_84_153#_c_76_n N_A3_M1004_g 9.69445e-19 $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_74 N_A_84_153#_c_77_n N_A3_M1004_g 0.0188436f $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_75 N_A_84_153#_c_79_n N_A3_M1004_g 0.00739122f $X=0.587 $Y=1.335 $X2=0 $Y2=0
cc_76 N_A_84_153#_c_72_n N_A3_c_161_n 0.009498f $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_77 N_A_84_153#_c_73_n N_A3_c_161_n 0.00398806f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_78 N_A_84_153#_c_79_n N_A3_c_161_n 0.00953438f $X=0.587 $Y=1.335 $X2=0 $Y2=0
cc_79 N_A_84_153#_c_72_n N_A3_c_162_n 7.32603e-19 $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_80 N_A_84_153#_c_73_n N_A3_c_162_n 0.0204651f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_81 N_A_84_153#_c_76_n N_A3_c_162_n 0.00183809f $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_82 N_A_84_153#_c_77_n N_A3_c_162_n 0.00188794f $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_83 N_A_84_153#_c_79_n N_A3_c_162_n 9.44371e-19 $X=0.587 $Y=1.335 $X2=0 $Y2=0
cc_84 N_A_84_153#_c_71_n N_A3_c_163_n 0.0144465f $X=0.51 $Y=0.765 $X2=0 $Y2=0
cc_85 N_A_84_153#_c_73_n N_A2_M1011_g 0.0112831f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_86 N_A_84_153#_c_73_n A2 0.0199689f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_87 N_A_84_153#_c_100_p A2 0.00561741f $X=2.565 $Y=0.48 $X2=0 $Y2=0
cc_88 N_A_84_153#_c_73_n N_A2_c_199_n 0.0042549f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_89 N_A_84_153#_c_73_n N_A1_M1005_g 0.0027888f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_90 N_A_84_153#_c_74_n N_A1_c_232_n 0.00106863f $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_91 N_A_84_153#_c_73_n N_A1_c_233_n 0.0126488f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_92 N_A_84_153#_c_73_n A1 0.0158056f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_93 N_A_84_153#_c_100_p A1 0.00837903f $X=2.565 $Y=0.48 $X2=0 $Y2=0
cc_94 N_A_84_153#_c_74_n A1 0.0152998f $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_95 N_A_84_153#_c_73_n N_A1_c_235_n 0.00384951f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_96 N_A_84_153#_c_100_p N_A1_c_235_n 0.00212703f $X=2.565 $Y=0.48 $X2=0 $Y2=0
cc_97 N_A_84_153#_c_74_n N_A1_c_235_n 3.30974e-19 $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_98 N_A_84_153#_c_100_p N_A1_c_236_n 0.00427658f $X=2.565 $Y=0.48 $X2=0 $Y2=0
cc_99 N_A_84_153#_c_74_n N_A1_c_236_n 8.22248e-19 $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_100 N_A_84_153#_c_73_n N_B1_M1002_g 0.00797418f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_101 N_A_84_153#_c_75_n N_B1_M1002_g 0.00622204f $X=2.65 $Y=1.945 $X2=0 $Y2=0
cc_102 N_A_84_153#_c_115_p N_B1_M1002_g 0.00305983f $X=2.65 $Y=2.05 $X2=0 $Y2=0
cc_103 N_A_84_153#_c_100_p N_B1_M1009_g 0.0121809f $X=2.565 $Y=0.48 $X2=0 $Y2=0
cc_104 N_A_84_153#_c_74_n N_B1_M1009_g 0.0162359f $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_105 N_A_84_153#_c_73_n N_B1_c_277_n 0.0178723f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_106 N_A_84_153#_c_74_n N_B1_c_277_n 8.00161e-19 $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_107 N_A_84_153#_c_115_p N_B1_c_277_n 6.05408e-19 $X=2.65 $Y=2.05 $X2=0 $Y2=0
cc_108 N_A_84_153#_c_78_n N_B1_c_277_n 0.00155932f $X=2.65 $Y=1.42 $X2=0 $Y2=0
cc_109 N_A_84_153#_c_75_n N_B2_c_328_n 0.00606295f $X=2.65 $Y=1.945 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_84_153#_c_115_p N_B2_c_328_n 0.00557035f $X=2.65 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_111 N_A_84_153#_c_74_n N_B2_M1010_g 0.00570585f $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_112 N_A_84_153#_c_75_n N_B2_c_330_n 0.00615314f $X=2.65 $Y=1.945 $X2=0 $Y2=0
cc_113 N_A_84_153#_c_75_n N_B2_c_325_n 0.00134514f $X=2.65 $Y=1.945 $X2=0 $Y2=0
cc_114 N_A_84_153#_c_74_n B2 0.0253256f $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_115 N_A_84_153#_c_75_n B2 0.0121599f $X=2.65 $Y=1.945 $X2=0 $Y2=0
cc_116 N_A_84_153#_c_78_n B2 0.00980344f $X=2.65 $Y=1.42 $X2=0 $Y2=0
cc_117 N_A_84_153#_c_74_n N_B2_c_327_n 0.00269599f $X=2.65 $Y=1.335 $X2=0 $Y2=0
cc_118 N_A_84_153#_c_78_n N_B2_c_327_n 0.00162615f $X=2.65 $Y=1.42 $X2=0 $Y2=0
cc_119 N_A_84_153#_M1006_g N_X_c_362_n 7.59046e-19 $X=0.555 $Y=2.135 $X2=0 $Y2=0
cc_120 N_A_84_153#_c_77_n N_X_c_362_n 2.0576e-19 $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_121 N_A_84_153#_M1006_g X 0.00833406f $X=0.555 $Y=2.135 $X2=0 $Y2=0
cc_122 N_A_84_153#_c_71_n X 0.0037387f $X=0.51 $Y=0.765 $X2=0 $Y2=0
cc_123 N_A_84_153#_c_72_n X 0.0269086f $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_124 N_A_84_153#_c_76_n X 0.0226083f $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_125 N_A_84_153#_M1006_g N_VPWR_c_382_n 0.00901074f $X=0.555 $Y=2.135 $X2=0
+ $Y2=0
cc_126 N_A_84_153#_c_73_n N_VPWR_c_382_n 0.0102168f $X=2.565 $Y=1.42 $X2=0 $Y2=0
cc_127 N_A_84_153#_c_76_n N_VPWR_c_382_n 0.00237481f $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_128 N_A_84_153#_c_77_n N_VPWR_c_382_n 0.00185142f $X=0.59 $Y=1.5 $X2=0 $Y2=0
cc_129 N_A_84_153#_M1006_g N_VPWR_c_377_n 0.00922208f $X=0.555 $Y=2.135 $X2=0
+ $Y2=0
cc_130 N_A_84_153#_M1006_g N_VPWR_c_374_n 0.00318254f $X=0.555 $Y=2.135 $X2=0
+ $Y2=0
cc_131 N_A_84_153#_c_73_n N_A_228_385#_c_402_n 0.0559609f $X=2.565 $Y=1.42 $X2=0
+ $Y2=0
cc_132 N_A_84_153#_c_75_n N_A_228_385#_c_402_n 0.00883968f $X=2.65 $Y=1.945
+ $X2=0 $Y2=0
cc_133 N_A_84_153#_c_75_n N_A_228_385#_c_403_n 0.0036687f $X=2.65 $Y=1.945 $X2=0
+ $Y2=0
cc_134 N_A_84_153#_M1002_d N_A_228_385#_c_404_n 0.00181172f $X=2.43 $Y=1.925
+ $X2=0 $Y2=0
cc_135 N_A_84_153#_c_115_p N_A_228_385#_c_404_n 0.0149318f $X=2.65 $Y=2.05 $X2=0
+ $Y2=0
cc_136 N_A_84_153#_M1006_g N_A_228_385#_c_406_n 0.00117556f $X=0.555 $Y=2.135
+ $X2=0 $Y2=0
cc_137 N_A_84_153#_c_73_n N_A_228_385#_c_406_n 0.0254179f $X=2.565 $Y=1.42 $X2=0
+ $Y2=0
cc_138 N_A_84_153#_c_71_n N_VGND_c_438_n 0.0115631f $X=0.51 $Y=0.765 $X2=0 $Y2=0
cc_139 N_A_84_153#_c_71_n N_VGND_c_441_n 0.00486043f $X=0.51 $Y=0.765 $X2=0
+ $Y2=0
cc_140 N_A_84_153#_c_72_n N_VGND_c_441_n 5.95547e-19 $X=0.51 $Y=0.915 $X2=0
+ $Y2=0
cc_141 N_A_84_153#_c_100_p N_VGND_c_442_n 0.0204358f $X=2.565 $Y=0.48 $X2=0
+ $Y2=0
cc_142 N_A_84_153#_M1007_d N_VGND_c_444_n 0.00377053f $X=2.04 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_A_84_153#_c_71_n N_VGND_c_444_n 0.00940677f $X=0.51 $Y=0.765 $X2=0
+ $Y2=0
cc_144 N_A_84_153#_c_72_n N_VGND_c_444_n 8.01698e-19 $X=0.51 $Y=0.915 $X2=0
+ $Y2=0
cc_145 N_A_84_153#_c_100_p N_VGND_c_444_n 0.0208169f $X=2.565 $Y=0.48 $X2=0
+ $Y2=0
cc_146 N_A_84_153#_c_100_p A_516_47# 0.00119247f $X=2.565 $Y=0.48 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A3_M1004_g N_A2_M1011_g 0.0498357f $X=1.065 $Y=2.135 $X2=0 $Y2=0
cc_148 N_A3_c_161_n A2 2.17885e-19 $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_149 N_A3_c_162_n A2 0.0115753f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_150 N_A3_c_163_n A2 0.00244762f $X=0.975 $Y=0.765 $X2=0 $Y2=0
cc_151 N_A3_c_161_n N_A2_c_199_n 0.0316786f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_152 N_A3_c_162_n N_A2_c_199_n 6.02259e-19 $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_153 N_A3_c_163_n N_A2_c_200_n 0.0316786f $X=0.975 $Y=0.765 $X2=0 $Y2=0
cc_154 N_A3_c_162_n X 0.00935866f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_155 N_A3_M1004_g N_VPWR_c_376_n 0.0136444f $X=1.065 $Y=2.135 $X2=0 $Y2=0
cc_156 N_A3_M1004_g N_A_228_385#_c_406_n 0.0107456f $X=1.065 $Y=2.135 $X2=0
+ $Y2=0
cc_157 N_A3_c_161_n N_VGND_c_438_n 0.00212039f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_158 N_A3_c_162_n N_VGND_c_438_n 0.0106804f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_159 N_A3_c_163_n N_VGND_c_438_n 0.00938678f $X=0.975 $Y=0.765 $X2=0 $Y2=0
cc_160 N_A3_c_161_n N_VGND_c_442_n 0.00148371f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_161 N_A3_c_163_n N_VGND_c_442_n 0.00585385f $X=0.975 $Y=0.765 $X2=0 $Y2=0
cc_162 N_A3_c_161_n N_VGND_c_444_n 0.00203757f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_163 N_A3_c_162_n N_VGND_c_444_n 0.00798778f $X=0.975 $Y=0.93 $X2=0 $Y2=0
cc_164 N_A3_c_163_n N_VGND_c_444_n 0.00661536f $X=0.975 $Y=0.765 $X2=0 $Y2=0
cc_165 N_A2_M1011_g N_A1_c_232_n 0.0107393f $X=1.495 $Y=2.135 $X2=0 $Y2=0
cc_166 N_A2_M1011_g N_A1_c_233_n 0.0357956f $X=1.495 $Y=2.135 $X2=0 $Y2=0
cc_167 A2 A1 0.0172972f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_168 N_A2_c_199_n A1 7.0674e-19 $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_169 N_A2_c_199_n N_A1_c_235_n 0.0210193f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_170 A2 N_A1_c_236_n 0.00786481f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_171 N_A2_c_200_n N_A1_c_236_n 0.0203159f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_172 N_A2_M1011_g B1 9.85313e-19 $X=1.495 $Y=2.135 $X2=0 $Y2=0
cc_173 N_A2_M1011_g N_VPWR_c_376_n 0.0103178f $X=1.495 $Y=2.135 $X2=0 $Y2=0
cc_174 N_A2_M1011_g N_A_228_385#_c_402_n 0.00922477f $X=1.495 $Y=2.135 $X2=0
+ $Y2=0
cc_175 N_A2_M1011_g N_A_228_385#_c_406_n 0.00892878f $X=1.495 $Y=2.135 $X2=0
+ $Y2=0
cc_176 A2 N_VGND_c_438_n 5.62159e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_177 A2 N_VGND_c_442_n 0.0108059f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_178 N_A2_c_199_n N_VGND_c_442_n 4.87387e-19 $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_179 N_A2_c_200_n N_VGND_c_442_n 0.00399843f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_180 A2 N_VGND_c_444_n 0.013237f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_181 N_A2_c_200_n N_VGND_c_444_n 0.00576827f $X=1.515 $Y=0.765 $X2=0 $Y2=0
cc_182 A2 A_300_47# 0.00573959f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_183 N_A1_M1005_g N_B1_M1002_g 0.026574f $X=1.925 $Y=2.135 $X2=0 $Y2=0
cc_184 N_A1_c_233_n N_B1_M1002_g 0.00495856f $X=1.945 $Y=1.485 $X2=0 $Y2=0
cc_185 N_A1_c_232_n N_B1_M1009_g 0.00680555f $X=1.945 $Y=1.335 $X2=0 $Y2=0
cc_186 A1 N_B1_M1009_g 0.00220277f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_187 N_A1_c_235_n N_B1_M1009_g 0.0195734f $X=2.055 $Y=0.93 $X2=0 $Y2=0
cc_188 N_A1_c_236_n N_B1_M1009_g 0.0143851f $X=2.055 $Y=0.765 $X2=0 $Y2=0
cc_189 N_A1_c_232_n N_B1_c_277_n 0.00495856f $X=1.945 $Y=1.335 $X2=0 $Y2=0
cc_190 N_A1_M1005_g B1 0.00622176f $X=1.925 $Y=2.135 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_VPWR_c_376_n 0.00122585f $X=1.925 $Y=2.135 $X2=0 $Y2=0
cc_192 N_A1_M1005_g N_A_228_385#_c_402_n 0.0143605f $X=1.925 $Y=2.135 $X2=0
+ $Y2=0
cc_193 N_A1_c_233_n N_A_228_385#_c_402_n 2.62616e-19 $X=1.945 $Y=1.485 $X2=0
+ $Y2=0
cc_194 N_A1_M1005_g N_A_228_385#_c_403_n 0.00124012f $X=1.925 $Y=2.135 $X2=0
+ $Y2=0
cc_195 N_A1_M1005_g N_A_228_385#_c_405_n 0.00122585f $X=1.925 $Y=2.135 $X2=0
+ $Y2=0
cc_196 N_A1_M1005_g N_A_228_385#_c_406_n 5.95433e-19 $X=1.925 $Y=2.135 $X2=0
+ $Y2=0
cc_197 N_A1_c_235_n N_VGND_c_442_n 0.00156426f $X=2.055 $Y=0.93 $X2=0 $Y2=0
cc_198 N_A1_c_236_n N_VGND_c_442_n 0.00585385f $X=2.055 $Y=0.765 $X2=0 $Y2=0
cc_199 A1 N_VGND_c_444_n 0.00543185f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_200 N_A1_c_235_n N_VGND_c_444_n 0.00201388f $X=2.055 $Y=0.93 $X2=0 $Y2=0
cc_201 N_A1_c_236_n N_VGND_c_444_n 0.00939409f $X=2.055 $Y=0.765 $X2=0 $Y2=0
cc_202 B1 N_B2_c_328_n 9.85313e-19 $X=3.035 $Y=2.69 $X2=-0.19 $Y2=-0.245
cc_203 N_B1_M1009_g N_B2_M1010_g 0.0541402f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_204 N_B1_M1002_g N_B2_c_330_n 0.0205792f $X=2.355 $Y=2.135 $X2=0 $Y2=0
cc_205 N_B1_M1002_g N_B2_c_325_n 0.00333873f $X=2.355 $Y=2.135 $X2=0 $Y2=0
cc_206 N_B1_c_277_n N_B2_c_325_n 0.00749625f $X=2.505 $Y=1.38 $X2=0 $Y2=0
cc_207 N_B1_M1009_g B2 5.47128e-19 $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_208 N_B1_M1009_g N_B2_c_327_n 0.00749625f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_209 B1 N_VPWR_c_375_n 0.0231906f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_210 B1 N_VPWR_c_376_n 0.0509719f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_211 B1 N_VPWR_c_379_n 0.0813186f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_212 N_B1_c_280_n N_VPWR_c_379_n 0.00786248f $X=2.265 $Y=2.88 $X2=0 $Y2=0
cc_213 B1 N_VPWR_c_374_n 0.0739144f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_214 N_B1_c_280_n N_VPWR_c_374_n 0.0109697f $X=2.265 $Y=2.88 $X2=0 $Y2=0
cc_215 N_B1_M1002_g N_A_228_385#_c_402_n 0.00193392f $X=2.355 $Y=2.135 $X2=0
+ $Y2=0
cc_216 N_B1_M1002_g N_A_228_385#_c_403_n 9.8981e-19 $X=2.355 $Y=2.135 $X2=0
+ $Y2=0
cc_217 N_B1_M1002_g N_A_228_385#_c_404_n 0.0144348f $X=2.355 $Y=2.135 $X2=0
+ $Y2=0
cc_218 B1 N_A_228_385#_c_404_n 0.0641676f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_219 N_B1_c_280_n N_A_228_385#_c_404_n 3.54189e-19 $X=2.265 $Y=2.88 $X2=0
+ $Y2=0
cc_220 B1 N_A_228_385#_c_405_n 0.0150744f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_221 N_B1_c_280_n N_A_228_385#_c_405_n 9.1826e-19 $X=2.265 $Y=2.88 $X2=0 $Y2=0
cc_222 N_B1_M1009_g N_VGND_c_440_n 0.00192016f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_223 N_B1_M1009_g N_VGND_c_442_n 0.00381677f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_224 N_B1_M1009_g N_VGND_c_444_n 0.00562796f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B2_c_328_n N_A_228_385#_c_404_n 0.0139375f $X=2.785 $Y=1.815 $X2=0
+ $Y2=0
cc_226 N_B2_c_330_n N_A_228_385#_c_430_n 0.00571065f $X=3 $Y=1.74 $X2=0 $Y2=0
cc_227 N_B2_c_325_n N_A_228_385#_c_430_n 2.19054e-19 $X=3.09 $Y=1.51 $X2=0 $Y2=0
cc_228 B2 N_A_228_385#_c_430_n 0.00695366f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_229 N_B2_M1010_g N_VGND_c_440_n 0.0105667f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_230 N_B2_c_324_n N_VGND_c_440_n 0.00438825f $X=3.022 $Y=0.99 $X2=0 $Y2=0
cc_231 B2 N_VGND_c_440_n 0.00857445f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_232 N_B2_M1010_g N_VGND_c_442_n 0.00486043f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_233 N_B2_M1010_g N_VGND_c_444_n 0.00818711f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_234 N_B2_c_324_n N_VGND_c_444_n 2.78168e-19 $X=3.022 $Y=0.99 $X2=0 $Y2=0
cc_235 B2 N_VGND_c_444_n 9.40005e-19 $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_236 N_X_c_360_n N_VGND_c_441_n 0.0110831f $X=0.29 $Y=0.495 $X2=0 $Y2=0
cc_237 N_X_M1001_s N_VGND_c_444_n 0.00363392f $X=0.165 $Y=0.235 $X2=0 $Y2=0
cc_238 N_X_c_360_n N_VGND_c_444_n 0.00883188f $X=0.29 $Y=0.495 $X2=0 $Y2=0
cc_239 N_VPWR_c_376_n N_A_228_385#_M1004_d 0.00180746f $X=1.625 $Y=2.42
+ $X2=-0.19 $Y2=-0.245
cc_240 N_VPWR_c_376_n N_A_228_385#_c_402_n 0.00463836f $X=1.625 $Y=2.42 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_399_p N_A_228_385#_c_402_n 0.0135835f $X=1.71 $Y=2.2 $X2=0 $Y2=0
cc_242 N_VPWR_c_376_n N_A_228_385#_c_405_n 0.012401f $X=1.625 $Y=2.42 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_376_n N_A_228_385#_c_406_n 0.0158698f $X=1.625 $Y=2.42 $X2=0
+ $Y2=0
cc_244 N_VGND_c_444_n A_228_47# 0.00899413f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_245 N_VGND_c_444_n A_300_47# 0.00790119f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_246 N_VGND_c_444_n A_516_47# 0.00368015f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
