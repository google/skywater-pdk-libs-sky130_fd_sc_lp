* File: sky130_fd_sc_lp__a311o_1.pxi.spice
* Created: Wed Sep  2 09:25:02 2020
* 
x_PM_SKY130_FD_SC_LP__A311O_1%A_80_21# N_A_80_21#_M1002_d N_A_80_21#_M1008_d
+ N_A_80_21#_M1010_d N_A_80_21#_c_58_n N_A_80_21#_M1004_g N_A_80_21#_M1003_g
+ N_A_80_21#_c_60_n N_A_80_21#_c_61_n N_A_80_21#_c_75_p N_A_80_21#_c_145_p
+ N_A_80_21#_c_68_n N_A_80_21#_c_69_n N_A_80_21#_c_93_p N_A_80_21#_c_62_n
+ N_A_80_21#_c_63_n N_A_80_21#_c_70_n N_A_80_21#_c_64_n N_A_80_21#_c_97_p
+ N_A_80_21#_c_65_n PM_SKY130_FD_SC_LP__A311O_1%A_80_21#
x_PM_SKY130_FD_SC_LP__A311O_1%A3 N_A3_M1005_g N_A3_M1009_g A3 N_A3_c_166_n
+ N_A3_c_167_n PM_SKY130_FD_SC_LP__A311O_1%A3
x_PM_SKY130_FD_SC_LP__A311O_1%A2 N_A2_M1000_g N_A2_c_201_n N_A2_M1001_g A2
+ N_A2_c_203_n PM_SKY130_FD_SC_LP__A311O_1%A2
x_PM_SKY130_FD_SC_LP__A311O_1%A1 N_A1_c_232_n N_A1_M1002_g N_A1_M1006_g A1
+ N_A1_c_234_n N_A1_c_235_n PM_SKY130_FD_SC_LP__A311O_1%A1
x_PM_SKY130_FD_SC_LP__A311O_1%B1 N_B1_M1007_g N_B1_M1011_g B1 B1 N_B1_c_266_n
+ N_B1_c_267_n PM_SKY130_FD_SC_LP__A311O_1%B1
x_PM_SKY130_FD_SC_LP__A311O_1%C1 N_C1_c_297_n N_C1_M1008_g N_C1_M1010_g C1
+ N_C1_c_300_n PM_SKY130_FD_SC_LP__A311O_1%C1
x_PM_SKY130_FD_SC_LP__A311O_1%X N_X_M1004_s N_X_M1003_s X X X X X X X
+ N_X_c_321_n X X PM_SKY130_FD_SC_LP__A311O_1%X
x_PM_SKY130_FD_SC_LP__A311O_1%VPWR N_VPWR_M1003_d N_VPWR_M1000_d N_VPWR_c_342_n
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n VPWR N_VPWR_c_346_n
+ N_VPWR_c_347_n N_VPWR_c_341_n N_VPWR_c_349_n PM_SKY130_FD_SC_LP__A311O_1%VPWR
x_PM_SKY130_FD_SC_LP__A311O_1%A_259_367# N_A_259_367#_M1005_d
+ N_A_259_367#_M1006_d N_A_259_367#_c_388_n N_A_259_367#_c_392_n
+ N_A_259_367#_c_389_n N_A_259_367#_c_390_n N_A_259_367#_c_401_n
+ PM_SKY130_FD_SC_LP__A311O_1%A_259_367#
x_PM_SKY130_FD_SC_LP__A311O_1%VGND N_VGND_M1004_d N_VGND_M1007_d N_VGND_c_405_n
+ VGND N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n
+ N_VGND_c_410_n PM_SKY130_FD_SC_LP__A311O_1%VGND
cc_1 VNB N_A_80_21#_c_58_n 0.0209655f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A_80_21#_M1003_g 0.00837681f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.465
cc_3 VNB N_A_80_21#_c_60_n 0.00247457f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.35
cc_4 VNB N_A_80_21#_c_61_n 0.00298409f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.695
cc_5 VNB N_A_80_21#_c_62_n 0.00740554f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=0.94
cc_6 VNB N_A_80_21#_c_63_n 0.0234718f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=0.38
cc_7 VNB N_A_80_21#_c_64_n 0.00216494f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.515
cc_8 VNB N_A_80_21#_c_65_n 0.0400493f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_9 VNB N_A3_M1005_g 0.00729831f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=1.835
cc_10 VNB A3 0.00582694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_c_166_n 0.0310785f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_12 VNB N_A3_c_167_n 0.0196479f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.515
cc_13 VNB N_A2_M1000_g 0.00881389f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=1.835
cc_14 VNB N_A2_c_201_n 0.0170504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A2 0.00643684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_203_n 0.0280639f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_17 VNB N_A1_c_232_n 0.0188291f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.235
cc_18 VNB N_A1_M1006_g 0.00889145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_234_n 0.0027301f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.465
cc_20 VNB N_A1_c_235_n 0.0347587f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.465
cc_21 VNB N_B1_M1011_g 0.00760125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B1 0.0120425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_266_n 0.0282525f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.515
cc_24 VNB N_B1_c_267_n 0.0190096f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.465
cc_25 VNB N_C1_c_297_n 0.0240612f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.235
cc_26 VNB N_C1_M1010_g 0.0102389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB C1 0.0214008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C1_c_300_n 0.0505818f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.515
cc_29 VNB N_X_c_321_n 0.0619051f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.94
cc_30 VNB N_VPWR_c_341_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=0.38
cc_31 VNB N_VGND_c_405_n 0.0055721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_406_n 0.0288393f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.515
cc_33 VNB N_VGND_c_407_n 0.0480179f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.358
cc_34 VNB N_VGND_c_408_n 0.0189813f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.94
cc_35 VNB N_VGND_c_409_n 0.209659f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=1.78
cc_36 VNB N_VGND_c_410_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=1.865
cc_37 VPB N_A_80_21#_M1003_g 0.0244956f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.465
cc_38 VPB N_A_80_21#_c_61_n 8.49974e-19 $X=-0.19 $Y=1.655 $X2=0.722 $Y2=1.695
cc_39 VPB N_A_80_21#_c_68_n 0.0286012f $X=-0.19 $Y=1.655 $X2=3.38 $Y2=1.78
cc_40 VPB N_A_80_21#_c_69_n 0.00150659f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.78
cc_41 VPB N_A_80_21#_c_70_n 0.0470856f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=1.98
cc_42 VPB N_A3_M1005_g 0.0196528f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=1.835
cc_43 VPB N_A2_M1000_g 0.0215834f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=1.835
cc_44 VPB N_A1_M1006_g 0.0227996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B1_M1011_g 0.0191528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_C1_M1010_g 0.0237659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB X 0.0158651f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_48 VPB N_X_c_321_n 0.0209509f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=0.94
cc_49 VPB X 0.0401219f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=1.98
cc_50 VPB N_VPWR_c_342_n 0.00453068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_343_n 0.00190031f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.465
cc_52 VPB N_VPWR_c_344_n 0.0232649f $X=-0.19 $Y=1.655 $X2=0.682 $Y2=1.358
cc_53 VPB N_VPWR_c_345_n 0.00496849f $X=-0.19 $Y=1.655 $X2=0.682 $Y2=1.35
cc_54 VPB N_VPWR_c_346_n 0.0154314f $X=-0.19 $Y=1.655 $X2=3.38 $Y2=1.78
cc_55 VPB N_VPWR_c_347_n 0.0412577f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=0.38
cc_56 VPB N_VPWR_c_341_n 0.0480006f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=0.38
cc_57 VPB N_VPWR_c_349_n 0.0106274f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=1.98
cc_58 N_A_80_21#_M1003_g N_A3_M1005_g 0.0218525f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_80_21#_c_61_n N_A3_M1005_g 0.00326716f $X=0.722 $Y=1.695 $X2=0 $Y2=0
cc_60 N_A_80_21#_c_68_n N_A3_M1005_g 0.014589f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_60_n A3 0.0274271f $X=0.61 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_75_p A3 0.0238548f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_68_n A3 0.0261991f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_65_n A3 0.0010165f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_60_n N_A3_c_166_n 0.001037f $X=0.61 $Y=1.35 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_75_p N_A3_c_166_n 0.00113794f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_68_n N_A3_c_166_n 0.00125536f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_65_n N_A3_c_166_n 0.0181368f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_58_n N_A3_c_167_n 0.0088162f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_60_n N_A3_c_167_n 0.00351468f $X=0.61 $Y=1.35 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_75_p N_A3_c_167_n 0.0132762f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_65_n N_A3_c_167_n 2.31016e-19 $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_68_n N_A2_M1000_g 0.0117585f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_75_p N_A2_c_201_n 0.0122311f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_75_p A2 0.0229808f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_68_n A2 0.0281519f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_75_p N_A2_c_203_n 0.00418655f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_68_n N_A2_c_203_n 0.00122615f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_75_p N_A1_c_232_n 0.0129291f $X=2.325 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_80_21#_c_93_p N_A1_c_232_n 0.0173822f $X=2.49 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_80_21#_c_68_n N_A1_M1006_g 0.0140335f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_75_p N_A1_c_234_n 0.0146286f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_68_n N_A1_c_234_n 0.0219231f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_97_p N_A1_c_234_n 0.00330322f $X=2.49 $Y=0.94 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_68_n N_A1_c_235_n 0.00597192f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_97_p N_A1_c_235_n 0.00574813f $X=2.49 $Y=0.94 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_68_n N_B1_M1011_g 0.0150921f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_70_n N_B1_M1011_g 0.00374372f $X=3.545 $Y=1.98 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_68_n B1 0.0527304f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_62_n B1 0.0370651f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_97_p B1 0.0104029f $X=2.49 $Y=0.94 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_68_n N_B1_c_266_n 0.00122069f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_62_n N_B1_c_266_n 0.00455309f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_93_p N_B1_c_267_n 0.00936545f $X=2.49 $Y=0.42 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_62_n N_B1_c_267_n 0.0133802f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_63_n N_B1_c_267_n 7.08516e-19 $X=3.545 $Y=0.38 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_62_n N_C1_c_297_n 0.0118487f $X=3.38 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_80_21#_c_63_n N_C1_c_297_n 0.011224f $X=3.545 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_80_21#_c_68_n N_C1_M1010_g 0.0161267f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_70_n N_C1_M1010_g 0.0242312f $X=3.545 $Y=1.98 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_68_n C1 0.0273718f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_62_n C1 0.0242962f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_68_n N_C1_c_300_n 0.00241399f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_62_n N_C1_c_300_n 0.00224126f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_105 N_A_80_21#_M1003_g X 0.00331613f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_69_n X 0.0019893f $X=0.84 $Y=1.78 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_64_n X 0.00253833f $X=0.682 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_65_n X 0.00467527f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_58_n N_X_c_321_n 0.013792f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_110 N_A_80_21#_M1003_g N_X_c_321_n 0.00597029f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_60_n N_X_c_321_n 0.0358619f $X=0.61 $Y=1.35 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_61_n N_X_c_321_n 0.0109355f $X=0.722 $Y=1.695 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_69_n N_X_c_321_n 0.0102104f $X=0.84 $Y=1.78 $X2=0 $Y2=0
cc_114 N_A_80_21#_M1003_g X 0.00806094f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_68_n N_VPWR_M1003_d 0.00250873f $X=3.38 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_80_21#_c_68_n N_VPWR_M1000_d 0.00593194f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_117 N_A_80_21#_M1003_g N_VPWR_c_342_n 0.00299807f $X=0.72 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_80_21#_c_68_n N_VPWR_c_342_n 0.0192006f $X=3.38 $Y=1.78 $X2=0 $Y2=0
cc_119 N_A_80_21#_M1003_g N_VPWR_c_344_n 0.0054895f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_70_n N_VPWR_c_347_n 0.0210467f $X=3.545 $Y=1.98 $X2=0 $Y2=0
cc_121 N_A_80_21#_M1010_d N_VPWR_c_341_n 0.00215158f $X=3.405 $Y=1.835 $X2=0
+ $Y2=0
cc_122 N_A_80_21#_M1003_g N_VPWR_c_341_n 0.0110471f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_70_n N_VPWR_c_341_n 0.0125689f $X=3.545 $Y=1.98 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_68_n N_A_259_367#_M1005_d 0.00176461f $X=3.38 $Y=1.78
+ $X2=-0.19 $Y2=-0.245
cc_125 N_A_80_21#_c_68_n N_A_259_367#_M1006_d 0.00298209f $X=3.38 $Y=1.78 $X2=0
+ $Y2=0
cc_126 N_A_80_21#_c_68_n N_A_259_367#_c_388_n 0.0153678f $X=3.38 $Y=1.78 $X2=0
+ $Y2=0
cc_127 N_A_80_21#_c_68_n N_A_259_367#_c_389_n 0.057779f $X=3.38 $Y=1.78 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_c_68_n N_A_259_367#_c_390_n 0.022455f $X=3.38 $Y=1.78 $X2=0
+ $Y2=0
cc_129 N_A_80_21#_c_68_n A_609_367# 0.00366293f $X=3.38 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_80_21#_c_60_n N_VGND_M1004_d 7.26477e-19 $X=0.61 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_80_21#_c_75_p N_VGND_M1004_d 0.00964959f $X=2.325 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_80_21#_c_145_p N_VGND_M1004_d 0.00345945f $X=0.84 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_80_21#_c_62_n N_VGND_M1007_d 0.00581937f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_62_n N_VGND_c_405_n 0.0219905f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_58_n N_VGND_c_406_n 0.0187867f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_75_p N_VGND_c_406_n 0.0270504f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_145_p N_VGND_c_406_n 0.0224686f $X=0.84 $Y=0.94 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_65_n N_VGND_c_406_n 8.62299e-19 $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_93_p N_VGND_c_407_n 0.0230625f $X=2.49 $Y=0.42 $X2=0 $Y2=0
cc_140 N_A_80_21#_c_63_n N_VGND_c_408_n 0.0210467f $X=3.545 $Y=0.38 $X2=0 $Y2=0
cc_141 N_A_80_21#_M1002_d N_VGND_c_409_n 0.00445577f $X=2.265 $Y=0.235 $X2=0
+ $Y2=0
cc_142 N_A_80_21#_M1008_d N_VGND_c_409_n 0.00215158f $X=3.405 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_c_58_n N_VGND_c_409_n 0.00917991f $X=0.475 $Y=1.185 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_c_75_p N_VGND_c_409_n 0.0351962f $X=2.325 $Y=0.94 $X2=0 $Y2=0
cc_145 N_A_80_21#_c_145_p N_VGND_c_409_n 0.00110872f $X=0.84 $Y=0.94 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_93_p N_VGND_c_409_n 0.0127519f $X=2.49 $Y=0.42 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_62_n N_VGND_c_409_n 0.012473f $X=3.38 $Y=0.94 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_63_n N_VGND_c_409_n 0.0125689f $X=3.545 $Y=0.38 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_75_p A_273_47# 0.00675285f $X=2.325 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_80_21#_c_75_p A_363_47# 0.00712813f $X=2.325 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A3_M1005_g N_A2_M1000_g 0.0264649f $X=1.22 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A3_c_166_n N_A2_M1000_g 0.0106398f $X=1.2 $Y=1.36 $X2=0 $Y2=0
cc_153 N_A3_c_167_n N_A2_c_201_n 0.0479754f $X=1.2 $Y=1.195 $X2=0 $Y2=0
cc_154 A3 A2 0.0264628f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_155 N_A3_c_166_n A2 0.00187066f $X=1.2 $Y=1.36 $X2=0 $Y2=0
cc_156 A3 N_A2_c_203_n 3.76596e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A3_c_167_n N_A2_c_203_n 0.0106398f $X=1.2 $Y=1.195 $X2=0 $Y2=0
cc_158 N_A3_M1005_g N_VPWR_c_342_n 0.00159201f $X=1.22 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A3_M1005_g N_VPWR_c_343_n 4.97243e-19 $X=1.22 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A3_M1005_g N_VPWR_c_346_n 0.0054895f $X=1.22 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A3_M1005_g N_VPWR_c_341_n 0.009976f $X=1.22 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A3_M1005_g N_A_259_367#_c_388_n 0.00209265f $X=1.22 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A3_M1005_g N_A_259_367#_c_392_n 0.00921684f $X=1.22 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A3_c_167_n N_VGND_c_406_n 0.0177068f $X=1.2 $Y=1.195 $X2=0 $Y2=0
cc_165 N_A3_c_167_n N_VGND_c_407_n 0.00487821f $X=1.2 $Y=1.195 $X2=0 $Y2=0
cc_166 N_A3_c_167_n N_VGND_c_409_n 0.00472938f $X=1.2 $Y=1.195 $X2=0 $Y2=0
cc_167 N_A2_c_201_n N_A1_c_232_n 0.0475941f $X=1.74 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A2_c_203_n N_A1_c_232_n 0.0214601f $X=1.74 $Y=1.35 $X2=-0.19 $Y2=-0.245
cc_169 N_A2_M1000_g N_A1_M1006_g 0.0168621f $X=1.65 $Y=2.465 $X2=0 $Y2=0
cc_170 A2 N_A1_c_234_n 0.026205f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A2_c_203_n N_A1_c_234_n 0.00102303f $X=1.74 $Y=1.35 $X2=0 $Y2=0
cc_172 N_A2_M1000_g N_A1_c_235_n 2.85986e-19 $X=1.65 $Y=2.465 $X2=0 $Y2=0
cc_173 A2 N_A1_c_235_n 3.97745e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A2_M1000_g N_VPWR_c_343_n 0.0141436f $X=1.65 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A2_M1000_g N_VPWR_c_346_n 0.00486043f $X=1.65 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A2_M1000_g N_VPWR_c_341_n 0.0082726f $X=1.65 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A2_M1000_g N_A_259_367#_c_389_n 0.0135719f $X=1.65 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A2_c_201_n N_VGND_c_406_n 0.00321926f $X=1.74 $Y=1.185 $X2=0 $Y2=0
cc_179 N_A2_c_201_n N_VGND_c_407_n 0.00585385f $X=1.74 $Y=1.185 $X2=0 $Y2=0
cc_180 N_A2_c_201_n N_VGND_c_409_n 0.00672817f $X=1.74 $Y=1.185 $X2=0 $Y2=0
cc_181 N_A1_c_235_n N_B1_M1011_g 0.0329663f $X=2.43 $Y=1.36 $X2=0 $Y2=0
cc_182 N_A1_c_234_n B1 0.0275497f $X=2.28 $Y=1.36 $X2=0 $Y2=0
cc_183 N_A1_c_235_n B1 0.0027403f $X=2.43 $Y=1.36 $X2=0 $Y2=0
cc_184 N_A1_c_234_n N_B1_c_266_n 2.32047e-19 $X=2.28 $Y=1.36 $X2=0 $Y2=0
cc_185 N_A1_c_235_n N_B1_c_266_n 0.0199836f $X=2.43 $Y=1.36 $X2=0 $Y2=0
cc_186 N_A1_c_232_n N_B1_c_267_n 0.0240858f $X=2.19 $Y=1.195 $X2=0 $Y2=0
cc_187 N_A1_M1006_g N_VPWR_c_343_n 0.0153317f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A1_M1006_g N_VPWR_c_347_n 0.00486043f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A1_M1006_g N_VPWR_c_341_n 0.00864313f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A1_M1006_g N_A_259_367#_c_389_n 0.015964f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A1_c_232_n N_VGND_c_407_n 0.00585385f $X=2.19 $Y=1.195 $X2=0 $Y2=0
cc_192 N_A1_c_232_n N_VGND_c_409_n 0.00705933f $X=2.19 $Y=1.195 $X2=0 $Y2=0
cc_193 N_B1_c_266_n N_C1_c_297_n 0.0618839f $X=2.88 $Y=1.35 $X2=-0.19 $Y2=-0.245
cc_194 N_B1_c_267_n N_C1_c_297_n 0.0254916f $X=2.88 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_195 B1 C1 0.0278754f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_196 N_B1_c_266_n C1 2.44563e-19 $X=2.88 $Y=1.35 $X2=0 $Y2=0
cc_197 N_B1_M1011_g N_C1_c_300_n 0.0618839f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_198 B1 N_C1_c_300_n 0.00272892f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_199 N_B1_M1011_g N_VPWR_c_343_n 0.00113392f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B1_M1011_g N_VPWR_c_347_n 0.00585385f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_201 N_B1_M1011_g N_VPWR_c_341_n 0.0109726f $X=2.97 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B1_c_267_n N_VGND_c_405_n 0.00409792f $X=2.88 $Y=1.185 $X2=0 $Y2=0
cc_203 N_B1_c_267_n N_VGND_c_407_n 0.00585385f $X=2.88 $Y=1.185 $X2=0 $Y2=0
cc_204 N_B1_c_267_n N_VGND_c_409_n 0.00703912f $X=2.88 $Y=1.185 $X2=0 $Y2=0
cc_205 N_C1_M1010_g N_VPWR_c_347_n 0.0054895f $X=3.33 $Y=2.465 $X2=0 $Y2=0
cc_206 N_C1_M1010_g N_VPWR_c_341_n 0.0108168f $X=3.33 $Y=2.465 $X2=0 $Y2=0
cc_207 N_C1_c_297_n N_VGND_c_405_n 0.00568878f $X=3.33 $Y=1.195 $X2=0 $Y2=0
cc_208 N_C1_c_297_n N_VGND_c_408_n 0.0054895f $X=3.33 $Y=1.195 $X2=0 $Y2=0
cc_209 N_C1_c_297_n N_VGND_c_409_n 0.00740406f $X=3.33 $Y=1.195 $X2=0 $Y2=0
cc_210 X N_VPWR_c_344_n 0.0393268f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_211 N_X_M1003_s N_VPWR_c_341_n 0.00215158f $X=0.38 $Y=1.835 $X2=0 $Y2=0
cc_212 X N_VPWR_c_341_n 0.0224827f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_213 N_X_c_321_n N_VGND_c_406_n 0.018528f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_214 N_X_M1004_s N_VGND_c_409_n 0.00371702f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_215 N_X_c_321_n N_VGND_c_409_n 0.0104192f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_216 N_VPWR_c_341_n N_A_259_367#_M1005_d 0.00380103f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_217 N_VPWR_c_341_n N_A_259_367#_M1006_d 0.00526034f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_346_n N_A_259_367#_c_392_n 0.015688f $X=1.7 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_c_341_n N_A_259_367#_c_392_n 0.00984745f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_220 N_VPWR_M1000_d N_A_259_367#_c_389_n 0.0131443f $X=1.725 $Y=1.835 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_343_n N_A_259_367#_c_389_n 0.0455532f $X=2.215 $Y=2.48 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_347_n N_A_259_367#_c_401_n 0.0212513f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_341_n N_A_259_367#_c_401_n 0.0127519f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_c_341_n A_609_367# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_225 N_VGND_c_409_n A_273_47# 0.0044696f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_226 N_VGND_c_409_n A_363_47# 0.0044696f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
