* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Y a_27_51# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_27_51# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_644_51# C a_1025_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_1025_65# C a_644_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_27_51# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y a_27_51# a_217_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_644_51# C a_1025_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR a_27_51# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_1025_65# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_217_51# a_27_51# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_644_51# B a_217_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 Y a_27_51# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VGND D a_1025_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 Y a_27_51# a_217_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_1025_65# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_217_51# B a_644_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VGND D a_1025_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_644_51# B a_217_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 a_217_51# B a_644_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_1025_65# C a_644_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 VPWR a_27_51# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_217_51# a_27_51# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
