* File: sky130_fd_sc_lp__a311o_m.pex.spice
* Created: Wed Sep  2 09:25:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311O_M%A3 3 7 9 12 14 15 16 21 23
c47 14 0 1.61905e-19 $X=0.72 $Y=0.925
r48 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=1.325
+ $X2=0.825 $Y2=1.49
r49 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=1.325
+ $X2=0.825 $Y2=1.16
r50 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.825
+ $Y=1.325 $X2=0.825 $Y2=1.325
r51 16 22 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=0.772 $Y=1.665
+ $X2=0.772 $Y2=1.325
r52 15 22 1.25721 $w=2.73e-07 $l=3e-08 $layer=LI1_cond $X=0.772 $Y=1.295
+ $X2=0.772 $Y2=1.325
r53 14 15 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.772 $Y=0.925
+ $X2=0.772 $Y2=1.295
r54 10 12 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=0.915 $Y=0.845
+ $X2=1.025 $Y2=0.845
r55 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.025 $Y=0.77
+ $X2=1.025 $Y2=0.845
r56 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.025 $Y=0.77
+ $X2=1.025 $Y2=0.45
r57 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.915 $Y=0.92
+ $X2=0.915 $Y2=0.845
r58 5 23 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.915 $Y=0.92
+ $X2=0.915 $Y2=1.16
r59 3 24 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=0.905 $Y=2.225
+ $X2=0.905 $Y2=1.49
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%A2 3 7 11 12 13 14 15 16 22
c46 7 0 4.37395e-20 $X=1.385 $Y=0.45
r47 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.365
+ $Y=1.325 $X2=1.365 $Y2=1.325
r48 16 23 9.4417 $w=4.13e-07 $l=3.4e-07 $layer=LI1_cond $X=1.322 $Y=1.665
+ $X2=1.322 $Y2=1.325
r49 15 23 0.833091 $w=4.13e-07 $l=3e-08 $layer=LI1_cond $X=1.322 $Y=1.295
+ $X2=1.322 $Y2=1.325
r50 14 15 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.322 $Y=0.925
+ $X2=1.322 $Y2=1.295
r51 13 14 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.322 $Y=0.555
+ $X2=1.322 $Y2=0.925
r52 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.365 $Y=1.665
+ $X2=1.365 $Y2=1.325
r53 11 12 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.665
+ $X2=1.365 $Y2=1.83
r54 10 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.16
+ $X2=1.365 $Y2=1.325
r55 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.385 $Y=0.45
+ $X2=1.385 $Y2=1.16
r56 3 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.335 $Y=2.225
+ $X2=1.335 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%A_54_154# 1 2 3 11 15 16 18 19 20 23 27 31
+ 33 36 38 39 41 43 46 48 50 55
c96 39 0 4.37395e-20 $X=2.065 $Y=0.735
c97 38 0 1.00858e-19 $X=2.61 $Y=0.735
c98 36 0 7.33235e-20 $X=2.14 $Y=2.94
c99 33 0 1.61348e-19 $X=2.61 $Y=2.94
c100 27 0 1.61905e-19 $X=0.475 $Y=1.805
r101 48 52 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.93 $Y=0.735
+ $X2=2.695 $Y2=0.735
r102 48 50 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2.93 $Y=0.65
+ $X2=2.93 $Y2=0.515
r103 44 55 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.16
+ $X2=2.695 $Y2=2.16
r104 44 46 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=2.78 $Y=2.16
+ $X2=2.93 $Y2=2.16
r105 42 55 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.695 $Y=2.265
+ $X2=2.695 $Y2=2.16
r106 42 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.695 $Y=2.265
+ $X2=2.695 $Y2=2.855
r107 41 55 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.695 $Y=2.055
+ $X2=2.695 $Y2=2.16
r108 40 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.82
+ $X2=2.695 $Y2=0.735
r109 40 41 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.695 $Y=0.82
+ $X2=2.695 $Y2=2.055
r110 38 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.735
+ $X2=2.695 $Y2=0.735
r111 38 39 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.61 $Y=0.735
+ $X2=2.065 $Y2=0.735
r112 36 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.14 $Y=2.94 $X2=2.14
+ $Y2=3.03
r113 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=2.94 $X2=2.14 $Y2=2.94
r114 33 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=2.94
+ $X2=2.695 $Y2=2.855
r115 33 35 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.61 $Y=2.94
+ $X2=2.14 $Y2=2.94
r116 29 39 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.96 $Y=0.65
+ $X2=2.065 $Y2=0.735
r117 29 31 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.96 $Y=0.65
+ $X2=1.96 $Y2=0.515
r118 25 27 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=0.345 $Y=1.805
+ $X2=0.475 $Y2=1.805
r119 21 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.345 $Y=0.845
+ $X2=0.555 $Y2=0.845
r120 19 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=3.03
+ $X2=2.14 $Y2=3.03
r121 19 20 730.691 $w=1.5e-07 $l=1.425e-06 $layer=POLY_cond $X=1.975 $Y=3.03
+ $X2=0.55 $Y2=3.03
r122 16 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.555 $Y=0.77
+ $X2=0.555 $Y2=0.845
r123 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.555 $Y=0.77
+ $X2=0.555 $Y2=0.45
r124 13 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=2.955
+ $X2=0.55 $Y2=3.03
r125 13 15 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.475 $Y=2.955
+ $X2=0.475 $Y2=2.225
r126 12 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.88
+ $X2=0.475 $Y2=1.805
r127 12 15 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.475 $Y=1.88
+ $X2=0.475 $Y2=2.225
r128 11 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.345 $Y=1.73
+ $X2=0.345 $Y2=1.805
r129 10 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.345 $Y=0.92
+ $X2=0.345 $Y2=0.845
r130 10 11 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.345 $Y=0.92
+ $X2=0.345 $Y2=1.73
r131 3 46 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=2.015 $X2=2.93 $Y2=2.16
r132 2 50 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.24 $X2=2.93 $Y2=0.515
r133 1 31 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.24 $X2=1.96 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%A1 3 8 10 11 12 15 17
c47 15 0 1.00858e-19 $X=1.905 $Y=1.665
c48 8 0 1.61348e-19 $X=1.925 $Y=2.225
r49 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.665
+ $X2=1.905 $Y2=1.83
r50 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.665
+ $X2=1.905 $Y2=1.5
r51 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.905
+ $Y=1.665 $X2=1.905 $Y2=1.665
r52 12 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=1.905 $Y2=1.665
r53 11 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.815 $Y=0.92
+ $X2=1.815 $Y2=1.5
r54 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.78 $Y=0.77
+ $X2=1.78 $Y2=0.92
r55 8 18 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.925 $Y=2.225
+ $X2=1.925 $Y2=1.83
r56 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.745 $Y=0.45
+ $X2=1.745 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%B1 3 7 9 12 13
r32 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.095
+ $X2=2.265 $Y2=1.26
r33 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.095
+ $X2=2.265 $Y2=0.93
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=1.095 $X2=2.265 $Y2=1.095
r35 9 13 6.49264 $w=3.53e-07 $l=2e-07 $layer=LI1_cond $X=2.252 $Y=1.295
+ $X2=2.252 $Y2=1.095
r36 7 15 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=2.355 $Y=2.225
+ $X2=2.355 $Y2=1.26
r37 3 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.175 $Y=0.45
+ $X2=2.175 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%C1 1 3 6 9 12 14 15 19
c32 6 0 6.36774e-20 $X=2.715 $Y=2.225
r33 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.425 $X2=3.09 $Y2=1.425
r34 19 21 15.6043 $w=2.78e-07 $l=9e-08 $layer=POLY_cond $X=3 $Y=1.455 $X2=3.09
+ $Y2=1.455
r35 15 22 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=3.105 $Y=1.665
+ $X2=3.105 $Y2=1.425
r36 14 22 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=3.105 $Y=1.295
+ $X2=3.105 $Y2=1.425
r37 10 12 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.715 $Y=0.845
+ $X2=3 $Y2=0.845
r38 9 19 17.1848 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3 $Y=1.26 $X2=3
+ $Y2=1.455
r39 8 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3 $Y=0.92 $X2=3
+ $Y2=0.845
r40 8 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3 $Y=0.92 $X2=3
+ $Y2=1.26
r41 4 19 49.4137 $w=2.78e-07 $l=3.69865e-07 $layer=POLY_cond $X=2.715 $Y=1.65
+ $X2=3 $Y2=1.455
r42 4 6 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.715 $Y=1.65
+ $X2=2.715 $Y2=2.225
r43 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.715 $Y=0.77
+ $X2=2.715 $Y2=0.845
r44 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.715 $Y=0.77
+ $X2=2.715 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%X 1 2 7 8 9 10 11 12 13 22
r19 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=2.405
+ $X2=0.29 $Y2=2.775
r20 12 35 10.4574 $w=2.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.29 $Y=2.405
+ $X2=0.29 $Y2=2.16
r21 11 35 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.29 $Y=2.035
+ $X2=0.29 $Y2=2.16
r22 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=2.035
r23 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r24 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.925 $X2=0.29
+ $Y2=1.295
r25 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.555 $X2=0.29
+ $Y2=0.925
r26 7 22 1.70732 $w=2.68e-07 $l=4e-08 $layer=LI1_cond $X=0.29 $Y=0.555 $X2=0.29
+ $Y2=0.515
r27 2 35 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.015 $X2=0.26 $Y2=2.16
r28 1 22 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.24 $X2=0.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%VPWR 1 2 9 13 16 17 18 24 33 34 37
r37 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r40 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.63 $Y2=3.33
r42 28 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.63 $Y2=3.33
r45 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 18 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 16 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 16 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.605 $Y=3.33 $X2=0.7
+ $Y2=3.33
r53 15 26 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 15 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.795 $Y=3.33 $X2=0.7
+ $Y2=3.33
r55 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r56 11 13 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.365
r57 7 17 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=3.33
r58 7 9 55.7464 $w=1.88e-07 $l=9.55e-07 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=2.29
r59 2 13 600 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.015 $X2=1.63 $Y2=2.365
r60 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.015 $X2=0.69 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%A_196_403# 1 2 7 9 14
c24 7 0 7.33235e-20 $X=2.035 $Y=2.015
r25 14 17 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=2.14 $Y=2.015
+ $X2=2.14 $Y2=2.16
r26 9 12 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=1.12 $Y=2.015
+ $X2=1.12 $Y2=2.16
r27 8 9 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.225 $Y=2.015 $X2=1.12
+ $Y2=2.015
r28 7 14 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.035 $Y=2.015
+ $X2=2.14 $Y2=2.015
r29 7 8 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.035 $Y=2.015
+ $X2=1.225 $Y2=2.015
r30 2 17 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.015 $X2=2.14 $Y2=2.16
r31 1 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.015 $X2=1.12 $Y2=2.16
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_M%VGND 1 2 9 13 16 17 18 20 33 34 37
r55 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r56 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r58 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r59 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r60 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r61 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r62 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.77
+ $Y2=0
r63 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.2
+ $Y2=0
r64 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r65 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r66 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.77
+ $Y2=0
r67 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r68 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r69 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r70 16 30 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r71 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.41
+ $Y2=0
r72 15 33 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=3.12
+ $Y2=0
r73 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.41
+ $Y2=0
r74 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0
r75 11 13 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0.365
r76 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085 $X2=0.77
+ $Y2=0
r77 7 9 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.77 $Y=0.085 $X2=0.77
+ $Y2=0.385
r78 2 13 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.24 $X2=2.41 $Y2=0.365
r79 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.24 $X2=0.77 $Y2=0.385
.ends

