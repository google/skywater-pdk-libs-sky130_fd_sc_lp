* File: sky130_fd_sc_lp__nor2_4.pxi.spice
* Created: Fri Aug 28 10:53:36 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_4%A N_A_c_69_n N_A_M1004_g N_A_M1000_g N_A_c_71_n
+ N_A_M1007_g N_A_M1003_g N_A_c_73_n N_A_M1013_g N_A_M1006_g N_A_c_75_n
+ N_A_M1014_g N_A_M1008_g A A A N_A_c_77_n N_A_c_78_n
+ PM_SKY130_FD_SC_LP__NOR2_4%A
x_PM_SKY130_FD_SC_LP__NOR2_4%B N_B_c_146_n N_B_M1001_g N_B_M1005_g N_B_c_147_n
+ N_B_M1002_g N_B_M1009_g N_B_M1011_g N_B_M1010_g N_B_c_149_n N_B_M1012_g
+ N_B_M1015_g B B B PM_SKY130_FD_SC_LP__NOR2_4%B
x_PM_SKY130_FD_SC_LP__NOR2_4%A_73_367# N_A_73_367#_M1000_d N_A_73_367#_M1003_d
+ N_A_73_367#_M1008_d N_A_73_367#_M1009_d N_A_73_367#_M1015_d
+ N_A_73_367#_c_221_n N_A_73_367#_c_222_n N_A_73_367#_c_223_n
+ N_A_73_367#_c_249_p N_A_73_367#_c_224_n N_A_73_367#_c_252_p
+ N_A_73_367#_c_240_n N_A_73_367#_c_274_p N_A_73_367#_c_242_n
+ N_A_73_367#_c_225_n N_A_73_367#_c_226_n N_A_73_367#_c_227_n
+ N_A_73_367#_c_256_p PM_SKY130_FD_SC_LP__NOR2_4%A_73_367#
x_PM_SKY130_FD_SC_LP__NOR2_4%VPWR N_VPWR_M1000_s N_VPWR_M1006_s N_VPWR_c_279_n
+ N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n VPWR
+ N_VPWR_c_284_n N_VPWR_c_278_n N_VPWR_c_286_n PM_SKY130_FD_SC_LP__NOR2_4%VPWR
x_PM_SKY130_FD_SC_LP__NOR2_4%Y N_Y_M1004_s N_Y_M1013_s N_Y_M1001_d N_Y_M1011_d
+ N_Y_M1005_s N_Y_M1010_s N_Y_c_335_n N_Y_c_347_n N_Y_c_351_n N_Y_c_336_n
+ N_Y_c_337_n N_Y_c_338_n N_Y_c_339_n N_Y_c_340_n N_Y_c_371_n N_Y_c_341_n
+ N_Y_c_377_n Y Y Y Y Y N_Y_c_342_n N_Y_c_343_n N_Y_c_389_n
+ PM_SKY130_FD_SC_LP__NOR2_4%Y
x_PM_SKY130_FD_SC_LP__NOR2_4%VGND N_VGND_M1004_d N_VGND_M1007_d N_VGND_M1014_d
+ N_VGND_M1002_s N_VGND_M1012_s N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n
+ N_VGND_c_430_n N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n
+ N_VGND_c_435_n N_VGND_c_436_n VGND N_VGND_c_437_n N_VGND_c_438_n
+ N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n
+ PM_SKY130_FD_SC_LP__NOR2_4%VGND
cc_1 VNB N_A_c_69_n 0.0209431f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.23
cc_2 VNB N_A_M1000_g 0.00756458f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_3 VNB N_A_c_71_n 0.0159873f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.23
cc_4 VNB N_A_M1003_g 0.0047805f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.465
cc_5 VNB N_A_c_73_n 0.0160323f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.23
cc_6 VNB N_A_M1006_g 0.0047805f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=2.465
cc_7 VNB N_A_c_75_n 0.0167005f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.23
cc_8 VNB N_A_M1008_g 0.0049341f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.465
cc_9 VNB N_A_c_77_n 0.0469624f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.395
cc_10 VNB N_A_c_78_n 0.0841593f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.395
cc_11 VNB N_B_c_146_n 0.0167005f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.23
cc_12 VNB N_B_c_147_n 0.015188f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.23
cc_13 VNB N_B_M1011_g 0.0208058f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.7
cc_14 VNB N_B_c_149_n 0.092589f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.7
cc_15 VNB N_B_M1012_g 0.0304659f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.56
cc_16 VNB B 0.0134068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_278_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.395
cc_18 VNB N_Y_c_335_n 0.00165022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_336_n 0.00193203f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.465
cc_20 VNB N_Y_c_337_n 0.0017546f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_21 VNB N_Y_c_338_n 0.00614561f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_22 VNB N_Y_c_339_n 9.39049e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_340_n 0.00610079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_341_n 0.00189235f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.395
cc_25 VNB N_Y_c_342_n 0.00193203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_343_n 8.0662e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_427_n 0.0345481f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.56
cc_28 VNB N_VGND_c_428_n 0.0135665f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=2.465
cc_29 VNB N_VGND_c_429_n 0.00106177f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.7
cc_30 VNB N_VGND_c_430_n 0.0151079f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.465
cc_31 VNB N_VGND_c_431_n 0.00802119f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_32 VNB N_VGND_c_432_n 0.00107947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_433_n 0.0151486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_434_n 0.0429576f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.395
cc_35 VNB N_VGND_c_435_n 0.0124854f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.395
cc_36 VNB N_VGND_c_436_n 0.00547551f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.395
cc_37 VNB N_VGND_c_437_n 0.0151079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_438_n 0.0149437f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.385
cc_39 VNB N_VGND_c_439_n 0.00494383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_440_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_441_n 0.00494383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_442_n 0.259955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A_M1000_g 0.0251848f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.465
cc_44 VPB N_A_M1003_g 0.018705f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.465
cc_45 VPB N_A_M1006_g 0.018705f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=2.465
cc_46 VPB N_A_M1008_g 0.0188897f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.465
cc_47 VPB N_B_M1005_g 0.0189822f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.465
cc_48 VPB N_B_M1009_g 0.0183504f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.465
cc_49 VPB N_B_M1010_g 0.0180507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B_c_149_n 0.0182847f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=0.7
cc_51 VPB N_B_M1015_g 0.024227f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_52 VPB B 0.0157359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_73_367#_c_221_n 0.0435297f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.56
cc_54 VPB N_A_73_367#_c_222_n 0.00295854f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=1.23
cc_55 VPB N_A_73_367#_c_223_n 0.0109903f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=0.7
cc_56 VPB N_A_73_367#_c_224_n 0.00742928f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_57 VPB N_A_73_367#_c_225_n 0.00746637f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.395
cc_58 VPB N_A_73_367#_c_226_n 0.0375006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_73_367#_c_227_n 0.00145912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_279_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.135 $Y2=0.7
cc_61 VPB N_VPWR_c_280_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.465
cc_62 VPB N_VPWR_c_281_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.565 $Y2=0.7
cc_63 VPB N_VPWR_c_282_n 0.0226949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_283_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=1.23
cc_65 VPB N_VPWR_c_284_n 0.0575369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_278_n 0.0597662f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.395
cc_67 VPB N_VPWR_c_286_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.395
cc_68 VPB Y 0.00230254f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.385
cc_69 N_A_c_75_n N_B_c_146_n 0.0188332f $X=1.995 $Y=1.23 $X2=-0.19 $Y2=-0.245
cc_70 N_A_M1008_g N_B_M1005_g 0.0188332f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_c_78_n N_B_c_149_n 0.0188332f $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_A_73_367#_c_222_n 0.0151162f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_A_73_367#_c_222_n 0.0142654f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A_c_77_n N_A_73_367#_c_222_n 0.049938f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_75 N_A_c_78_n N_A_73_367#_c_222_n 0.0030363f $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_76 N_A_c_77_n N_A_73_367#_c_223_n 0.0230972f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_A_73_367#_c_224_n 0.0177962f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_M1008_g N_A_73_367#_c_224_n 0.0140463f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_c_77_n N_A_73_367#_c_224_n 0.00593195f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_80 N_A_c_78_n N_A_73_367#_c_224_n 7.11963e-19 $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_81 N_A_c_77_n N_A_73_367#_c_227_n 0.0160899f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_82 N_A_c_78_n N_A_73_367#_c_227_n 0.00232957f $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_VPWR_c_279_n 0.0162594f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_84 N_A_M1003_g N_VPWR_c_279_n 0.0142791f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_M1006_g N_VPWR_c_279_n 7.27171e-19 $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_M1003_g N_VPWR_c_280_n 0.00486043f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_M1006_g N_VPWR_c_280_n 0.00486043f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VPWR_c_281_n 7.27171e-19 $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_M1006_g N_VPWR_c_281_n 0.0145199f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_M1008_g N_VPWR_c_281_n 0.0156848f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A_M1000_g N_VPWR_c_282_n 0.00486043f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A_M1008_g N_VPWR_c_284_n 0.00486043f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_93 N_A_M1000_g N_VPWR_c_278_n 0.0093368f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_M1003_g N_VPWR_c_278_n 0.00824727f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_M1006_g N_VPWR_c_278_n 0.00824727f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A_M1008_g N_VPWR_c_278_n 0.0082726f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_c_69_n N_Y_c_335_n 3.41554e-19 $X=0.705 $Y=1.23 $X2=0 $Y2=0
cc_98 N_A_c_71_n N_Y_c_335_n 3.41554e-19 $X=1.135 $Y=1.23 $X2=0 $Y2=0
cc_99 N_A_c_71_n N_Y_c_347_n 0.0122129f $X=1.135 $Y=1.23 $X2=0 $Y2=0
cc_100 N_A_c_73_n N_Y_c_347_n 0.0156946f $X=1.565 $Y=1.23 $X2=0 $Y2=0
cc_101 N_A_c_77_n N_Y_c_347_n 0.032921f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_102 N_A_c_78_n N_Y_c_347_n 6.666e-19 $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_103 N_A_c_77_n N_Y_c_351_n 0.0154649f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_104 N_A_c_78_n N_Y_c_351_n 7.50045e-19 $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_105 N_A_c_73_n N_Y_c_336_n 7.72865e-19 $X=1.565 $Y=1.23 $X2=0 $Y2=0
cc_106 N_A_c_75_n N_Y_c_336_n 8.31937e-19 $X=1.995 $Y=1.23 $X2=0 $Y2=0
cc_107 N_A_c_73_n N_Y_c_337_n 0.00238169f $X=1.565 $Y=1.23 $X2=0 $Y2=0
cc_108 N_A_c_75_n N_Y_c_337_n 0.00131553f $X=1.995 $Y=1.23 $X2=0 $Y2=0
cc_109 N_A_c_77_n N_Y_c_337_n 0.00882247f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_110 N_A_c_78_n N_Y_c_337_n 0.00726591f $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_111 N_A_c_78_n N_Y_c_338_n 0.0157832f $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_112 N_A_c_77_n N_Y_c_339_n 0.0198083f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_113 N_A_c_78_n N_Y_c_339_n 0.00980647f $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_114 N_A_M1008_g Y 5.28685e-19 $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_c_78_n N_Y_c_343_n 3.52244e-19 $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_116 N_A_c_69_n N_VGND_c_427_n 0.015641f $X=0.705 $Y=1.23 $X2=0 $Y2=0
cc_117 N_A_c_71_n N_VGND_c_427_n 5.40202e-19 $X=1.135 $Y=1.23 $X2=0 $Y2=0
cc_118 N_A_c_77_n N_VGND_c_427_n 0.0258603f $X=1.44 $Y=1.395 $X2=0 $Y2=0
cc_119 N_A_c_69_n N_VGND_c_428_n 0.00448994f $X=0.705 $Y=1.23 $X2=0 $Y2=0
cc_120 N_A_c_71_n N_VGND_c_428_n 0.00448994f $X=1.135 $Y=1.23 $X2=0 $Y2=0
cc_121 N_A_c_69_n N_VGND_c_429_n 4.91826e-19 $X=0.705 $Y=1.23 $X2=0 $Y2=0
cc_122 N_A_c_71_n N_VGND_c_429_n 0.009899f $X=1.135 $Y=1.23 $X2=0 $Y2=0
cc_123 N_A_c_73_n N_VGND_c_429_n 0.00996113f $X=1.565 $Y=1.23 $X2=0 $Y2=0
cc_124 N_A_c_75_n N_VGND_c_429_n 5.0204e-19 $X=1.995 $Y=1.23 $X2=0 $Y2=0
cc_125 N_A_c_73_n N_VGND_c_430_n 0.00448994f $X=1.565 $Y=1.23 $X2=0 $Y2=0
cc_126 N_A_c_75_n N_VGND_c_430_n 0.00540763f $X=1.995 $Y=1.23 $X2=0 $Y2=0
cc_127 N_A_c_75_n N_VGND_c_431_n 0.00261519f $X=1.995 $Y=1.23 $X2=0 $Y2=0
cc_128 N_A_c_69_n N_VGND_c_442_n 0.00812427f $X=0.705 $Y=1.23 $X2=0 $Y2=0
cc_129 N_A_c_71_n N_VGND_c_442_n 0.00812427f $X=1.135 $Y=1.23 $X2=0 $Y2=0
cc_130 N_A_c_73_n N_VGND_c_442_n 0.00812427f $X=1.565 $Y=1.23 $X2=0 $Y2=0
cc_131 N_A_c_75_n N_VGND_c_442_n 0.0102588f $X=1.995 $Y=1.23 $X2=0 $Y2=0
cc_132 N_B_M1005_g N_A_73_367#_c_224_n 9.18928e-19 $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_133 N_B_M1005_g N_A_73_367#_c_240_n 0.012237f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B_M1009_g N_A_73_367#_c_240_n 0.0121905f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B_M1010_g N_A_73_367#_c_242_n 0.012237f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B_M1015_g N_A_73_367#_c_242_n 0.012237f $X=3.715 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B_c_149_n N_A_73_367#_c_226_n 9.72225e-19 $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_138 B N_A_73_367#_c_226_n 0.0232232f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_139 N_B_M1005_g N_VPWR_c_281_n 0.00109252f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_140 N_B_M1005_g N_VPWR_c_284_n 0.00357877f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_141 N_B_M1009_g N_VPWR_c_284_n 0.00357877f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_142 N_B_M1010_g N_VPWR_c_284_n 0.00357877f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_143 N_B_M1015_g N_VPWR_c_284_n 0.00357877f $X=3.715 $Y=2.465 $X2=0 $Y2=0
cc_144 N_B_M1005_g N_VPWR_c_278_n 0.00537654f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_145 N_B_M1009_g N_VPWR_c_278_n 0.0053512f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B_M1010_g N_VPWR_c_278_n 0.0053512f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B_M1015_g N_VPWR_c_278_n 0.00638567f $X=3.715 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B_c_149_n N_Y_c_337_n 3.38162e-19 $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_149 N_B_c_149_n N_Y_c_338_n 0.0203073f $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_150 N_B_c_147_n N_Y_c_340_n 0.0106108f $X=2.855 $Y=1.23 $X2=0 $Y2=0
cc_151 N_B_M1011_g N_Y_c_340_n 0.0135515f $X=3.285 $Y=0.7 $X2=0 $Y2=0
cc_152 N_B_c_149_n N_Y_c_340_n 0.0135738f $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_153 N_B_M1012_g N_Y_c_340_n 0.00399542f $X=3.715 $Y=0.7 $X2=0 $Y2=0
cc_154 B N_Y_c_340_n 0.0555055f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_155 N_B_M1009_g N_Y_c_371_n 0.0167543f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B_M1010_g N_Y_c_371_n 0.013068f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_157 N_B_c_149_n N_Y_c_371_n 5.58524e-19 $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_158 B N_Y_c_371_n 0.0283495f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_159 N_B_M1011_g N_Y_c_341_n 7.72646e-19 $X=3.285 $Y=0.7 $X2=0 $Y2=0
cc_160 N_B_M1012_g N_Y_c_341_n 8.22925e-19 $X=3.715 $Y=0.7 $X2=0 $Y2=0
cc_161 N_B_c_149_n N_Y_c_377_n 6.36674e-19 $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_162 B N_Y_c_377_n 0.0169271f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_163 N_B_M1005_g Y 0.00270861f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_164 N_B_M1009_g Y 0.00290081f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B_c_149_n Y 0.00804807f $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_166 B Y 0.0157298f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_167 N_B_c_146_n N_Y_c_342_n 8.31937e-19 $X=2.425 $Y=1.23 $X2=0 $Y2=0
cc_168 N_B_c_147_n N_Y_c_342_n 7.72865e-19 $X=2.855 $Y=1.23 $X2=0 $Y2=0
cc_169 N_B_c_146_n N_Y_c_343_n 0.00157784f $X=2.425 $Y=1.23 $X2=0 $Y2=0
cc_170 N_B_M1011_g N_Y_c_343_n 3.8605e-19 $X=3.285 $Y=0.7 $X2=0 $Y2=0
cc_171 N_B_c_149_n N_Y_c_343_n 0.0191749f $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_172 B N_Y_c_343_n 0.0113432f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B_M1009_g N_Y_c_389_n 5.3453e-19 $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_174 N_B_M1010_g N_Y_c_389_n 3.25901e-19 $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B_c_149_n N_Y_c_389_n 2.50825e-19 $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_176 N_B_c_146_n N_VGND_c_431_n 0.00261457f $X=2.425 $Y=1.23 $X2=0 $Y2=0
cc_177 N_B_c_146_n N_VGND_c_432_n 5.62865e-19 $X=2.425 $Y=1.23 $X2=0 $Y2=0
cc_178 N_B_c_147_n N_VGND_c_432_n 0.0107373f $X=2.855 $Y=1.23 $X2=0 $Y2=0
cc_179 N_B_M1011_g N_VGND_c_432_n 0.0107286f $X=3.285 $Y=0.7 $X2=0 $Y2=0
cc_180 N_B_M1012_g N_VGND_c_432_n 5.6142e-19 $X=3.715 $Y=0.7 $X2=0 $Y2=0
cc_181 N_B_c_149_n N_VGND_c_434_n 0.00430618f $X=3.715 $Y=1.345 $X2=0 $Y2=0
cc_182 N_B_M1012_g N_VGND_c_434_n 0.00713368f $X=3.715 $Y=0.7 $X2=0 $Y2=0
cc_183 B N_VGND_c_434_n 0.0176324f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_184 N_B_c_146_n N_VGND_c_437_n 0.00540763f $X=2.425 $Y=1.23 $X2=0 $Y2=0
cc_185 N_B_c_147_n N_VGND_c_437_n 0.00448994f $X=2.855 $Y=1.23 $X2=0 $Y2=0
cc_186 N_B_M1011_g N_VGND_c_438_n 0.00448994f $X=3.285 $Y=0.7 $X2=0 $Y2=0
cc_187 N_B_M1012_g N_VGND_c_438_n 0.00540763f $X=3.715 $Y=0.7 $X2=0 $Y2=0
cc_188 N_B_c_146_n N_VGND_c_442_n 0.0102588f $X=2.425 $Y=1.23 $X2=0 $Y2=0
cc_189 N_B_c_147_n N_VGND_c_442_n 0.00812427f $X=2.855 $Y=1.23 $X2=0 $Y2=0
cc_190 N_B_M1011_g N_VGND_c_442_n 0.00812427f $X=3.285 $Y=0.7 $X2=0 $Y2=0
cc_191 N_B_M1012_g N_VGND_c_442_n 0.0109826f $X=3.715 $Y=0.7 $X2=0 $Y2=0
cc_192 N_A_73_367#_c_222_n N_VPWR_M1000_s 0.0017721f $X=1.255 $Y=1.827 $X2=-0.19
+ $Y2=1.655
cc_193 N_A_73_367#_c_224_n N_VPWR_M1006_s 0.0017721f $X=2.115 $Y=1.827 $X2=0
+ $Y2=0
cc_194 N_A_73_367#_c_222_n N_VPWR_c_279_n 0.0172384f $X=1.255 $Y=1.827 $X2=0
+ $Y2=0
cc_195 N_A_73_367#_c_249_p N_VPWR_c_280_n 0.0124525f $X=1.35 $Y=1.98 $X2=0 $Y2=0
cc_196 N_A_73_367#_c_224_n N_VPWR_c_281_n 0.0172384f $X=2.115 $Y=1.827 $X2=0
+ $Y2=0
cc_197 N_A_73_367#_c_221_n N_VPWR_c_282_n 0.0178111f $X=0.49 $Y=1.98 $X2=0 $Y2=0
cc_198 N_A_73_367#_c_252_p N_VPWR_c_284_n 0.0135879f $X=2.225 $Y=2.905 $X2=0
+ $Y2=0
cc_199 N_A_73_367#_c_240_n N_VPWR_c_284_n 0.0341772f $X=2.95 $Y=2.99 $X2=0 $Y2=0
cc_200 N_A_73_367#_c_242_n N_VPWR_c_284_n 0.0336481f $X=3.805 $Y=2.99 $X2=0
+ $Y2=0
cc_201 N_A_73_367#_c_225_n N_VPWR_c_284_n 0.0189827f $X=3.95 $Y=2.905 $X2=0
+ $Y2=0
cc_202 N_A_73_367#_c_256_p N_VPWR_c_284_n 0.0148297f $X=3.077 $Y=2.99 $X2=0
+ $Y2=0
cc_203 N_A_73_367#_M1000_d N_VPWR_c_278_n 0.00371702f $X=0.365 $Y=1.835 $X2=0
+ $Y2=0
cc_204 N_A_73_367#_M1003_d N_VPWR_c_278_n 0.00536646f $X=1.21 $Y=1.835 $X2=0
+ $Y2=0
cc_205 N_A_73_367#_M1008_d N_VPWR_c_278_n 0.00376625f $X=2.07 $Y=1.835 $X2=0
+ $Y2=0
cc_206 N_A_73_367#_M1009_d N_VPWR_c_278_n 0.00220343f $X=2.93 $Y=1.835 $X2=0
+ $Y2=0
cc_207 N_A_73_367#_M1015_d N_VPWR_c_278_n 0.00215159f $X=3.79 $Y=1.835 $X2=0
+ $Y2=0
cc_208 N_A_73_367#_c_221_n N_VPWR_c_278_n 0.0100304f $X=0.49 $Y=1.98 $X2=0 $Y2=0
cc_209 N_A_73_367#_c_249_p N_VPWR_c_278_n 0.00730901f $X=1.35 $Y=1.98 $X2=0
+ $Y2=0
cc_210 N_A_73_367#_c_252_p N_VPWR_c_278_n 0.00855309f $X=2.225 $Y=2.905 $X2=0
+ $Y2=0
cc_211 N_A_73_367#_c_240_n N_VPWR_c_278_n 0.0216081f $X=2.95 $Y=2.99 $X2=0 $Y2=0
cc_212 N_A_73_367#_c_242_n N_VPWR_c_278_n 0.0210442f $X=3.805 $Y=2.99 $X2=0
+ $Y2=0
cc_213 N_A_73_367#_c_225_n N_VPWR_c_278_n 0.0112745f $X=3.95 $Y=2.905 $X2=0
+ $Y2=0
cc_214 N_A_73_367#_c_256_p N_VPWR_c_278_n 0.00991381f $X=3.077 $Y=2.99 $X2=0
+ $Y2=0
cc_215 N_A_73_367#_c_240_n N_Y_M1005_s 0.00332774f $X=2.95 $Y=2.99 $X2=0 $Y2=0
cc_216 N_A_73_367#_c_242_n N_Y_M1010_s 0.00332344f $X=3.805 $Y=2.99 $X2=0 $Y2=0
cc_217 N_A_73_367#_c_224_n N_Y_c_338_n 0.0337117f $X=2.115 $Y=1.827 $X2=0 $Y2=0
cc_218 N_A_73_367#_c_224_n N_Y_c_339_n 0.0173551f $X=2.115 $Y=1.827 $X2=0 $Y2=0
cc_219 N_A_73_367#_M1009_d N_Y_c_371_n 0.0034107f $X=2.93 $Y=1.835 $X2=0 $Y2=0
cc_220 N_A_73_367#_c_274_p N_Y_c_371_n 0.0135055f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A_73_367#_c_242_n N_Y_c_377_n 0.0126348f $X=3.805 $Y=2.99 $X2=0 $Y2=0
cc_222 N_A_73_367#_c_224_n Y 0.00896206f $X=2.115 $Y=1.827 $X2=0 $Y2=0
cc_223 N_A_73_367#_c_240_n N_Y_c_389_n 0.0124713f $X=2.95 $Y=2.99 $X2=0 $Y2=0
cc_224 N_VPWR_c_278_n N_Y_M1005_s 0.00225186f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_225 N_VPWR_c_278_n N_Y_M1010_s 0.00225186f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_226 N_Y_c_347_n N_VGND_M1007_d 0.00331065f $X=1.685 $Y=0.955 $X2=0 $Y2=0
cc_227 N_Y_c_340_n N_VGND_M1002_s 0.00176461f $X=3.405 $Y=1.17 $X2=0 $Y2=0
cc_228 N_Y_c_335_n N_VGND_c_427_n 0.0232367f $X=0.92 $Y=0.43 $X2=0 $Y2=0
cc_229 N_Y_c_335_n N_VGND_c_428_n 0.0126758f $X=0.92 $Y=0.43 $X2=0 $Y2=0
cc_230 N_Y_c_335_n N_VGND_c_429_n 0.0168579f $X=0.92 $Y=0.43 $X2=0 $Y2=0
cc_231 N_Y_c_347_n N_VGND_c_429_n 0.0170777f $X=1.685 $Y=0.955 $X2=0 $Y2=0
cc_232 N_Y_c_336_n N_VGND_c_429_n 0.0168719f $X=1.78 $Y=0.43 $X2=0 $Y2=0
cc_233 N_Y_c_336_n N_VGND_c_430_n 0.0150357f $X=1.78 $Y=0.43 $X2=0 $Y2=0
cc_234 N_Y_c_336_n N_VGND_c_431_n 0.00111144f $X=1.78 $Y=0.43 $X2=0 $Y2=0
cc_235 N_Y_c_337_n N_VGND_c_431_n 0.00269003f $X=1.802 $Y=1.325 $X2=0 $Y2=0
cc_236 N_Y_c_338_n N_VGND_c_431_n 0.0222825f $X=2.505 $Y=1.442 $X2=0 $Y2=0
cc_237 N_Y_c_342_n N_VGND_c_431_n 0.00111144f $X=2.64 $Y=0.43 $X2=0 $Y2=0
cc_238 N_Y_c_343_n N_VGND_c_431_n 0.00295513f $X=2.62 $Y=1.56 $X2=0 $Y2=0
cc_239 N_Y_c_340_n N_VGND_c_432_n 0.0170777f $X=3.405 $Y=1.17 $X2=0 $Y2=0
cc_240 N_Y_c_341_n N_VGND_c_432_n 0.0249373f $X=3.5 $Y=0.43 $X2=0 $Y2=0
cc_241 N_Y_c_342_n N_VGND_c_432_n 0.0249392f $X=2.64 $Y=0.43 $X2=0 $Y2=0
cc_242 N_Y_c_340_n N_VGND_c_434_n 0.00166817f $X=3.405 $Y=1.17 $X2=0 $Y2=0
cc_243 N_Y_c_341_n N_VGND_c_434_n 0.00112187f $X=3.5 $Y=0.43 $X2=0 $Y2=0
cc_244 N_Y_c_342_n N_VGND_c_437_n 0.0150357f $X=2.64 $Y=0.43 $X2=0 $Y2=0
cc_245 N_Y_c_341_n N_VGND_c_438_n 0.0146985f $X=3.5 $Y=0.43 $X2=0 $Y2=0
cc_246 N_Y_c_335_n N_VGND_c_442_n 0.00727431f $X=0.92 $Y=0.43 $X2=0 $Y2=0
cc_247 N_Y_c_336_n N_VGND_c_442_n 0.00862857f $X=1.78 $Y=0.43 $X2=0 $Y2=0
cc_248 N_Y_c_341_n N_VGND_c_442_n 0.00843511f $X=3.5 $Y=0.43 $X2=0 $Y2=0
cc_249 N_Y_c_342_n N_VGND_c_442_n 0.00862857f $X=2.64 $Y=0.43 $X2=0 $Y2=0
