* File: sky130_fd_sc_lp__mux2i_0.pxi.spice
* Created: Wed Sep  2 10:00:55 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2I_0%S N_S_M1006_g N_S_M1002_g N_S_c_68_n N_S_M1003_g
+ N_S_M1004_g N_S_c_69_n N_S_c_77_n N_S_c_78_n N_S_c_111_p N_S_c_124_p
+ N_S_c_112_p N_S_c_79_n N_S_c_113_p N_S_c_70_n N_S_c_71_n S S N_S_c_83_n
+ N_S_c_73_n N_S_c_84_n PM_SKY130_FD_SC_LP__MUX2I_0%S
x_PM_SKY130_FD_SC_LP__MUX2I_0%A_47_48# N_A_47_48#_M1006_s N_A_47_48#_M1002_s
+ N_A_47_48#_M1001_g N_A_47_48#_c_181_n N_A_47_48#_M1007_g N_A_47_48#_c_182_n
+ N_A_47_48#_c_183_n N_A_47_48#_c_184_n N_A_47_48#_c_192_n N_A_47_48#_c_185_n
+ N_A_47_48#_c_186_n N_A_47_48#_c_187_n N_A_47_48#_c_188_n N_A_47_48#_c_193_n
+ N_A_47_48#_c_189_n PM_SKY130_FD_SC_LP__MUX2I_0%A_47_48#
x_PM_SKY130_FD_SC_LP__MUX2I_0%A0 N_A0_M1008_g N_A0_M1000_g A0 A0 N_A0_c_252_n
+ N_A0_c_253_n N_A0_c_257_n N_A0_c_254_n N_A0_c_255_n
+ PM_SKY130_FD_SC_LP__MUX2I_0%A0
x_PM_SKY130_FD_SC_LP__MUX2I_0%A1 N_A1_M1009_g N_A1_c_311_n N_A1_M1005_g A1 A1
+ N_A1_c_314_n PM_SKY130_FD_SC_LP__MUX2I_0%A1
x_PM_SKY130_FD_SC_LP__MUX2I_0%VPWR N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_c_363_n
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n VPWR
+ N_VPWR_c_368_n N_VPWR_c_362_n N_VPWR_c_370_n PM_SKY130_FD_SC_LP__MUX2I_0%VPWR
x_PM_SKY130_FD_SC_LP__MUX2I_0%Y N_Y_M1008_d N_Y_M1009_d N_Y_c_410_n N_Y_c_411_n
+ N_Y_c_412_n N_Y_c_409_n N_Y_c_430_n Y PM_SKY130_FD_SC_LP__MUX2I_0%Y
x_PM_SKY130_FD_SC_LP__MUX2I_0%VGND N_VGND_M1006_d N_VGND_M1003_d N_VGND_c_462_n
+ N_VGND_c_463_n N_VGND_c_464_n VGND N_VGND_c_465_n N_VGND_c_466_n
+ N_VGND_c_467_n PM_SKY130_FD_SC_LP__MUX2I_0%VGND
cc_1 VNB N_S_M1006_g 0.0729955f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.45
cc_2 VNB N_S_c_68_n 0.019889f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.77
cc_3 VNB N_S_c_69_n 0.029273f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=0.845
cc_4 VNB N_S_c_70_n 0.010915f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.79
cc_5 VNB N_S_c_71_n 0.0184747f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.79
cc_6 VNB S 0.00310299f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_S_c_73_n 0.0584013f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=1.625
cc_8 VNB N_A_47_48#_c_181_n 0.0110762f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.45
cc_9 VNB N_A_47_48#_c_182_n 0.0174537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_47_48#_c_183_n 0.0226346f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.845
cc_11 VNB N_A_47_48#_c_184_n 0.0179458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_47_48#_c_185_n 0.0243895f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=2.99
cc_13 VNB N_A_47_48#_c_186_n 0.0094722f $X=-0.19 $Y=-0.245 $X2=3.005 $Y2=2.505
cc_14 VNB N_A_47_48#_c_187_n 0.0147956f $X=-0.19 $Y=-0.245 $X2=3.005 $Y2=1.79
cc_15 VNB N_A_47_48#_c_188_n 0.0339143f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.79
cc_16 VNB N_A_47_48#_c_189_n 0.0155868f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_17 VNB N_A0_c_252_n 0.0284302f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.845
cc_18 VNB N_A0_c_253_n 0.0174643f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=0.845
cc_19 VNB N_A0_c_254_n 0.00348478f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=2.245
cc_20 VNB N_A0_c_255_n 0.0117987f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_21 VNB N_A1_c_311_n 0.0222267f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=2.01
cc_22 VNB N_A1_M1005_g 0.0474113f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.77
cc_23 VNB A1 0.0108023f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=0.92
cc_24 VNB N_A1_c_314_n 0.0257125f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=2.775
cc_25 VNB N_VPWR_c_362_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=2.59
cc_26 VNB N_Y_c_409_n 0.00904014f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=2.295
cc_27 VNB N_VGND_c_462_n 0.00580638f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=0.45
cc_28 VNB N_VGND_c_463_n 0.0144502f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.625
cc_29 VNB N_VGND_c_464_n 0.0210785f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=2.775
cc_30 VNB N_VGND_c_465_n 0.049114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_466_n 0.0268595f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=2.675
cc_32 VNB N_VGND_c_467_n 0.193905f $X=-0.19 $Y=-0.245 $X2=3.005 $Y2=2.505
cc_33 VPB N_S_M1006_g 0.00134357f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.45
cc_34 VPB N_S_M1002_g 0.0429043f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.775
cc_35 VPB N_S_M1004_g 0.0212402f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=2.775
cc_36 VPB N_S_c_77_n 0.0126709f $X=-0.19 $Y=1.655 $X2=1.47 $Y2=2.127
cc_37 VPB N_S_c_78_n 0.00347051f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=2.905
cc_38 VPB N_S_c_79_n 0.00889853f $X=-0.19 $Y=1.655 $X2=2.87 $Y2=2.59
cc_39 VPB N_S_c_70_n 0.0091257f $X=-0.19 $Y=1.655 $X2=2.975 $Y2=1.79
cc_40 VPB N_S_c_71_n 0.0909798f $X=-0.19 $Y=1.655 $X2=2.975 $Y2=1.79
cc_41 VPB S 0.00292105f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_42 VPB N_S_c_83_n 0.0335339f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.845
cc_43 VPB N_S_c_84_n 0.00597513f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=2.01
cc_44 VPB N_A_47_48#_c_181_n 0.0193687f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=0.45
cc_45 VPB N_A_47_48#_M1007_g 0.0254055f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=2.295
cc_46 VPB N_A_47_48#_c_192_n 0.0231897f $X=-0.19 $Y=1.655 $X2=1.47 $Y2=2.127
cc_47 VPB N_A_47_48#_c_193_n 0.0430924f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_48 VPB N_A_47_48#_c_189_n 0.0406089f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_49 VPB N_A0_M1000_g 0.0311126f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.775
cc_50 VPB N_A0_c_257_n 0.0339764f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=2.127
cc_51 VPB N_A0_c_254_n 9.98064e-19 $X=-0.19 $Y=1.655 $X2=1.57 $Y2=2.245
cc_52 VPB N_A1_M1009_g 0.0442674f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.45
cc_53 VPB A1 0.00706168f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=0.92
cc_54 VPB N_A1_c_314_n 0.016768f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=2.775
cc_55 VPB N_VPWR_c_363_n 0.00883274f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=0.77
cc_56 VPB N_VPWR_c_364_n 0.0122366f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.625
cc_57 VPB N_VPWR_c_365_n 0.0114896f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=2.775
cc_58 VPB N_VPWR_c_366_n 0.0352477f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=2.775
cc_59 VPB N_VPWR_c_367_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_368_n 0.025192f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=0.845
cc_61 VPB N_VPWR_c_362_n 0.0523319f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=2.59
cc_62 VPB N_VPWR_c_370_n 0.00632158f $X=-0.19 $Y=1.655 $X2=3.005 $Y2=1.79
cc_63 VPB N_Y_c_410_n 0.0025188f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=0.77
cc_64 VPB N_Y_c_411_n 0.00890398f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=0.45
cc_65 VPB N_Y_c_412_n 0.00591428f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=0.92
cc_66 VPB N_Y_c_409_n 0.00397915f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=2.295
cc_67 N_S_M1006_g N_A_47_48#_c_181_n 0.00692556f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_68 N_S_c_77_n N_A_47_48#_c_181_n 0.00363332f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_69 S N_A_47_48#_c_181_n 0.00549894f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_70 N_S_c_83_n N_A_47_48#_c_181_n 0.0138047f $X=0.665 $Y=1.845 $X2=0 $Y2=0
cc_71 N_S_M1002_g N_A_47_48#_M1007_g 0.0195944f $X=0.755 $Y=2.775 $X2=0 $Y2=0
cc_72 N_S_c_77_n N_A_47_48#_M1007_g 0.00861831f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_73 N_S_c_78_n N_A_47_48#_M1007_g 0.00649812f $X=1.57 $Y=2.905 $X2=0 $Y2=0
cc_74 N_S_M1006_g N_A_47_48#_c_182_n 0.01593f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_75 N_S_c_77_n N_A_47_48#_c_184_n 0.00331809f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_76 N_S_M1002_g N_A_47_48#_c_192_n 0.0138047f $X=0.755 $Y=2.775 $X2=0 $Y2=0
cc_77 N_S_c_77_n N_A_47_48#_c_192_n 0.0155317f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_78 N_S_M1006_g N_A_47_48#_c_185_n 0.0104287f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_79 N_S_M1006_g N_A_47_48#_c_186_n 0.0177605f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_80 N_S_c_77_n N_A_47_48#_c_186_n 0.00488944f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_81 S N_A_47_48#_c_186_n 0.0316177f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_82 N_S_c_83_n N_A_47_48#_c_186_n 9.6352e-19 $X=0.665 $Y=1.845 $X2=0 $Y2=0
cc_83 N_S_M1006_g N_A_47_48#_c_187_n 0.0371579f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_84 N_S_M1006_g N_A_47_48#_c_188_n 0.0150582f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_85 N_S_M1002_g N_A_47_48#_c_193_n 0.00874167f $X=0.755 $Y=2.775 $X2=0 $Y2=0
cc_86 N_S_c_83_n N_A_47_48#_c_193_n 0.00196152f $X=0.665 $Y=1.845 $X2=0 $Y2=0
cc_87 N_S_c_84_n N_A_47_48#_c_193_n 0.0156054f $X=0.712 $Y=2.01 $X2=0 $Y2=0
cc_88 N_S_M1006_g N_A_47_48#_c_189_n 0.0153456f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_89 N_S_M1002_g N_A_47_48#_c_189_n 0.00495406f $X=0.755 $Y=2.775 $X2=0 $Y2=0
cc_90 S N_A_47_48#_c_189_n 0.037621f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_91 N_S_c_84_n N_A_47_48#_c_189_n 0.0205459f $X=0.712 $Y=2.01 $X2=0 $Y2=0
cc_92 N_S_c_77_n N_A0_M1000_g 4.99564e-19 $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_93 N_S_c_111_p N_A0_M1000_g 0.0115345f $X=2.385 $Y=2.99 $X2=0 $Y2=0
cc_94 N_S_c_112_p N_A0_M1000_g 0.00444742f $X=2.47 $Y=2.905 $X2=0 $Y2=0
cc_95 N_S_c_113_p N_A0_M1000_g 0.00150285f $X=2.555 $Y=2.59 $X2=0 $Y2=0
cc_96 N_S_c_71_n N_A0_M1000_g 0.0491507f $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_97 N_S_c_77_n N_A0_c_257_n 2.79128e-19 $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_98 N_S_c_71_n N_A0_c_257_n 0.0174333f $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_99 N_S_c_71_n N_A0_c_254_n 2.74778e-19 $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_100 N_S_c_73_n N_A0_c_254_n 0.00186061f $X=2.87 $Y=1.625 $X2=0 $Y2=0
cc_101 N_S_c_69_n N_A0_c_255_n 8.91099e-19 $X=2.675 $Y=0.845 $X2=0 $Y2=0
cc_102 N_S_c_73_n N_A0_c_255_n 0.00171058f $X=2.87 $Y=1.625 $X2=0 $Y2=0
cc_103 N_S_c_77_n N_A1_M1009_g 0.00586022f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_104 N_S_c_78_n N_A1_M1009_g 0.0030879f $X=1.57 $Y=2.905 $X2=0 $Y2=0
cc_105 N_S_c_111_p N_A1_M1009_g 0.0125941f $X=2.385 $Y=2.99 $X2=0 $Y2=0
cc_106 N_S_c_124_p N_A1_M1009_g 0.00113993f $X=1.67 $Y=2.99 $X2=0 $Y2=0
cc_107 N_S_c_68_n N_A1_M1005_g 0.0445426f $X=2.495 $Y=0.77 $X2=0 $Y2=0
cc_108 N_S_c_73_n N_A1_M1005_g 0.0147745f $X=2.87 $Y=1.625 $X2=0 $Y2=0
cc_109 N_S_M1006_g A1 3.32708e-19 $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_110 N_S_c_77_n A1 0.0492433f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_111 S A1 0.0256035f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_112 N_S_c_83_n A1 5.36148e-19 $X=0.665 $Y=1.845 $X2=0 $Y2=0
cc_113 N_S_c_77_n N_A1_c_314_n 0.00151689f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_114 N_S_c_79_n N_VPWR_M1004_d 0.00411434f $X=2.87 $Y=2.59 $X2=0 $Y2=0
cc_115 N_S_c_70_n N_VPWR_M1004_d 7.52137e-19 $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_116 N_S_M1002_g N_VPWR_c_363_n 0.0103081f $X=0.755 $Y=2.775 $X2=0 $Y2=0
cc_117 N_S_c_77_n N_VPWR_c_363_n 0.0261817f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_118 N_S_c_78_n N_VPWR_c_363_n 0.0152195f $X=1.57 $Y=2.905 $X2=0 $Y2=0
cc_119 N_S_M1004_g N_VPWR_c_364_n 0.00887148f $X=2.675 $Y=2.775 $X2=0 $Y2=0
cc_120 N_S_c_79_n N_VPWR_c_364_n 0.0220938f $X=2.87 $Y=2.59 $X2=0 $Y2=0
cc_121 N_S_c_71_n N_VPWR_c_364_n 7.47547e-19 $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_122 N_S_c_79_n N_VPWR_c_365_n 0.00164315f $X=2.87 $Y=2.59 $X2=0 $Y2=0
cc_123 N_S_M1004_g N_VPWR_c_366_n 0.00355956f $X=2.675 $Y=2.775 $X2=0 $Y2=0
cc_124 N_S_c_111_p N_VPWR_c_366_n 0.0512322f $X=2.385 $Y=2.99 $X2=0 $Y2=0
cc_125 N_S_c_124_p N_VPWR_c_366_n 0.01044f $X=1.67 $Y=2.99 $X2=0 $Y2=0
cc_126 N_S_c_79_n N_VPWR_c_366_n 0.00235807f $X=2.87 $Y=2.59 $X2=0 $Y2=0
cc_127 N_S_M1002_g N_VPWR_c_368_n 0.00549615f $X=0.755 $Y=2.775 $X2=0 $Y2=0
cc_128 N_S_M1002_g N_VPWR_c_362_n 0.0115192f $X=0.755 $Y=2.775 $X2=0 $Y2=0
cc_129 N_S_M1004_g N_VPWR_c_362_n 0.00424676f $X=2.675 $Y=2.775 $X2=0 $Y2=0
cc_130 N_S_c_111_p N_VPWR_c_362_n 0.0320806f $X=2.385 $Y=2.99 $X2=0 $Y2=0
cc_131 N_S_c_124_p N_VPWR_c_362_n 0.00776497f $X=1.67 $Y=2.99 $X2=0 $Y2=0
cc_132 N_S_c_79_n N_VPWR_c_362_n 0.00828415f $X=2.87 $Y=2.59 $X2=0 $Y2=0
cc_133 N_S_c_78_n A_292_491# 0.00143999f $X=1.57 $Y=2.905 $X2=-0.19 $Y2=-0.245
cc_134 N_S_c_124_p A_292_491# 9.38685e-19 $X=1.67 $Y=2.99 $X2=-0.19 $Y2=-0.245
cc_135 N_S_c_111_p N_Y_M1009_d 0.00482499f $X=2.385 $Y=2.99 $X2=0 $Y2=0
cc_136 N_S_c_78_n N_Y_c_410_n 0.00949835f $X=1.57 $Y=2.905 $X2=0 $Y2=0
cc_137 N_S_c_111_p N_Y_c_410_n 0.0180965f $X=2.385 $Y=2.99 $X2=0 $Y2=0
cc_138 N_S_M1004_g N_Y_c_411_n 0.00251186f $X=2.675 $Y=2.775 $X2=0 $Y2=0
cc_139 N_S_c_111_p N_Y_c_411_n 0.0047952f $X=2.385 $Y=2.99 $X2=0 $Y2=0
cc_140 N_S_c_79_n N_Y_c_411_n 0.0097169f $X=2.87 $Y=2.59 $X2=0 $Y2=0
cc_141 N_S_c_113_p N_Y_c_411_n 0.0134794f $X=2.555 $Y=2.59 $X2=0 $Y2=0
cc_142 N_S_c_70_n N_Y_c_411_n 0.0134931f $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_143 N_S_c_71_n N_Y_c_411_n 0.00463258f $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_144 N_S_c_77_n N_Y_c_412_n 0.00713124f $X=1.47 $Y=2.127 $X2=0 $Y2=0
cc_145 N_S_c_78_n N_Y_c_412_n 0.00764219f $X=1.57 $Y=2.905 $X2=0 $Y2=0
cc_146 N_S_c_68_n N_Y_c_409_n 0.0044405f $X=2.495 $Y=0.77 $X2=0 $Y2=0
cc_147 N_S_c_69_n N_Y_c_409_n 0.0139247f $X=2.675 $Y=0.845 $X2=0 $Y2=0
cc_148 N_S_c_70_n N_Y_c_409_n 0.0379154f $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_149 N_S_c_71_n N_Y_c_409_n 0.0159979f $X=2.975 $Y=1.79 $X2=0 $Y2=0
cc_150 N_S_c_73_n N_Y_c_409_n 0.039256f $X=2.87 $Y=1.625 $X2=0 $Y2=0
cc_151 N_S_c_68_n N_Y_c_430_n 0.0207554f $X=2.495 $Y=0.77 $X2=0 $Y2=0
cc_152 N_S_c_111_p A_465_491# 0.00189419f $X=2.385 $Y=2.99 $X2=-0.19 $Y2=-0.245
cc_153 N_S_c_112_p A_465_491# 0.00258422f $X=2.47 $Y=2.905 $X2=-0.19 $Y2=-0.245
cc_154 N_S_c_113_p A_465_491# 0.00363438f $X=2.555 $Y=2.59 $X2=-0.19 $Y2=-0.245
cc_155 N_S_M1006_g N_VGND_c_462_n 0.00528832f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_156 N_S_c_68_n N_VGND_c_464_n 0.00601189f $X=2.495 $Y=0.77 $X2=0 $Y2=0
cc_157 N_S_c_68_n N_VGND_c_465_n 0.00360601f $X=2.495 $Y=0.77 $X2=0 $Y2=0
cc_158 N_S_c_69_n N_VGND_c_465_n 0.00128799f $X=2.675 $Y=0.845 $X2=0 $Y2=0
cc_159 N_S_M1006_g N_VGND_c_466_n 0.00544432f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_160 N_S_M1006_g N_VGND_c_467_n 0.00744121f $X=0.575 $Y=0.45 $X2=0 $Y2=0
cc_161 N_S_c_68_n N_VGND_c_467_n 0.00664647f $X=2.495 $Y=0.77 $X2=0 $Y2=0
cc_162 N_S_c_69_n N_VGND_c_467_n 0.0013464f $X=2.675 $Y=0.845 $X2=0 $Y2=0
cc_163 N_A_47_48#_c_186_n N_A0_c_252_n 5.38951e-19 $X=1.055 $Y=0.935 $X2=0 $Y2=0
cc_164 N_A_47_48#_c_187_n N_A0_c_252_n 0.0268962f $X=1.055 $Y=0.935 $X2=0 $Y2=0
cc_165 N_A_47_48#_c_182_n N_A0_c_253_n 0.0268962f $X=1.055 $Y=0.77 $X2=0 $Y2=0
cc_166 N_A_47_48#_c_183_n N_A0_c_255_n 0.00185524f $X=1.055 $Y=1.275 $X2=0 $Y2=0
cc_167 N_A_47_48#_c_186_n N_A0_c_255_n 0.0361978f $X=1.055 $Y=0.935 $X2=0 $Y2=0
cc_168 N_A_47_48#_c_187_n N_A0_c_255_n 3.6596e-19 $X=1.055 $Y=0.935 $X2=0 $Y2=0
cc_169 N_A_47_48#_c_181_n N_A1_M1009_g 0.00721505f $X=1.145 $Y=2.05 $X2=0 $Y2=0
cc_170 N_A_47_48#_c_192_n N_A1_M1009_g 0.0669528f $X=1.385 $Y=2.125 $X2=0 $Y2=0
cc_171 N_A_47_48#_c_181_n A1 0.0126411f $X=1.145 $Y=2.05 $X2=0 $Y2=0
cc_172 N_A_47_48#_c_184_n A1 2.84752e-19 $X=1.055 $Y=1.44 $X2=0 $Y2=0
cc_173 N_A_47_48#_c_192_n A1 0.00157452f $X=1.385 $Y=2.125 $X2=0 $Y2=0
cc_174 N_A_47_48#_c_186_n A1 0.0114033f $X=1.055 $Y=0.935 $X2=0 $Y2=0
cc_175 N_A_47_48#_c_184_n N_A1_c_314_n 0.0273467f $X=1.055 $Y=1.44 $X2=0 $Y2=0
cc_176 N_A_47_48#_M1007_g N_VPWR_c_363_n 0.0101899f $X=1.385 $Y=2.775 $X2=0
+ $Y2=0
cc_177 N_A_47_48#_c_192_n N_VPWR_c_363_n 0.00109888f $X=1.385 $Y=2.125 $X2=0
+ $Y2=0
cc_178 N_A_47_48#_c_193_n N_VPWR_c_363_n 0.0454407f $X=0.54 $Y=2.6 $X2=0 $Y2=0
cc_179 N_A_47_48#_M1007_g N_VPWR_c_366_n 0.00585385f $X=1.385 $Y=2.775 $X2=0
+ $Y2=0
cc_180 N_A_47_48#_c_193_n N_VPWR_c_368_n 0.0370396f $X=0.54 $Y=2.6 $X2=0 $Y2=0
cc_181 N_A_47_48#_M1002_s N_VPWR_c_362_n 0.00215817f $X=0.415 $Y=2.455 $X2=0
+ $Y2=0
cc_182 N_A_47_48#_M1007_g N_VPWR_c_362_n 0.0112268f $X=1.385 $Y=2.775 $X2=0
+ $Y2=0
cc_183 N_A_47_48#_c_193_n N_VPWR_c_362_n 0.023589f $X=0.54 $Y=2.6 $X2=0 $Y2=0
cc_184 N_A_47_48#_c_182_n N_VGND_c_462_n 0.00550301f $X=1.055 $Y=0.77 $X2=0
+ $Y2=0
cc_185 N_A_47_48#_c_186_n N_VGND_c_462_n 0.02721f $X=1.055 $Y=0.935 $X2=0 $Y2=0
cc_186 N_A_47_48#_c_187_n N_VGND_c_462_n 0.00386685f $X=1.055 $Y=0.935 $X2=0
+ $Y2=0
cc_187 N_A_47_48#_c_182_n N_VGND_c_465_n 0.0058025f $X=1.055 $Y=0.77 $X2=0 $Y2=0
cc_188 N_A_47_48#_c_187_n N_VGND_c_465_n 6.77057e-19 $X=1.055 $Y=0.935 $X2=0
+ $Y2=0
cc_189 N_A_47_48#_c_185_n N_VGND_c_466_n 0.0272019f $X=0.36 $Y=0.45 $X2=0 $Y2=0
cc_190 N_A_47_48#_M1006_s N_VGND_c_467_n 0.00214782f $X=0.235 $Y=0.24 $X2=0
+ $Y2=0
cc_191 N_A_47_48#_c_182_n N_VGND_c_467_n 0.00642602f $X=1.055 $Y=0.77 $X2=0
+ $Y2=0
cc_192 N_A_47_48#_c_185_n N_VGND_c_467_n 0.0168268f $X=0.36 $Y=0.45 $X2=0 $Y2=0
cc_193 N_A_47_48#_c_186_n N_VGND_c_467_n 0.0137861f $X=1.055 $Y=0.935 $X2=0
+ $Y2=0
cc_194 N_A_47_48#_c_187_n N_VGND_c_467_n 9.23014e-19 $X=1.055 $Y=0.935 $X2=0
+ $Y2=0
cc_195 N_A0_M1000_g N_A1_M1009_g 0.0256436f $X=2.25 $Y=2.775 $X2=0 $Y2=0
cc_196 N_A0_c_254_n N_A1_M1009_g 9.73356e-19 $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_197 N_A0_c_257_n N_A1_c_311_n 0.00829656f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_198 N_A0_c_254_n N_A1_c_311_n 0.0101278f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_199 N_A0_c_255_n N_A1_c_311_n 0.0144244f $X=2.195 $Y=1.095 $X2=0 $Y2=0
cc_200 N_A0_c_252_n N_A1_M1005_g 0.0183783f $X=1.625 $Y=0.935 $X2=0 $Y2=0
cc_201 N_A0_c_253_n N_A1_M1005_g 0.0181708f $X=1.625 $Y=0.77 $X2=0 $Y2=0
cc_202 N_A0_c_255_n N_A1_M1005_g 0.0236851f $X=2.195 $Y=1.095 $X2=0 $Y2=0
cc_203 N_A0_c_257_n A1 6.37787e-19 $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_204 N_A0_c_254_n A1 0.0250451f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_205 N_A0_c_255_n A1 0.0311515f $X=2.195 $Y=1.095 $X2=0 $Y2=0
cc_206 N_A0_c_252_n N_A1_c_314_n 0.0177726f $X=1.625 $Y=0.935 $X2=0 $Y2=0
cc_207 N_A0_c_257_n N_A1_c_314_n 0.0211721f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_208 N_A0_c_254_n N_A1_c_314_n 0.00352882f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_209 N_A0_c_255_n N_A1_c_314_n 0.0106408f $X=2.195 $Y=1.095 $X2=0 $Y2=0
cc_210 N_A0_M1000_g N_VPWR_c_364_n 0.00128169f $X=2.25 $Y=2.775 $X2=0 $Y2=0
cc_211 N_A0_M1000_g N_VPWR_c_366_n 0.00357877f $X=2.25 $Y=2.775 $X2=0 $Y2=0
cc_212 N_A0_M1000_g N_VPWR_c_362_n 0.00564676f $X=2.25 $Y=2.775 $X2=0 $Y2=0
cc_213 N_A0_M1000_g N_Y_c_410_n 0.00354316f $X=2.25 $Y=2.775 $X2=0 $Y2=0
cc_214 N_A0_M1000_g N_Y_c_411_n 0.0125073f $X=2.25 $Y=2.775 $X2=0 $Y2=0
cc_215 N_A0_c_257_n N_Y_c_411_n 9.92475e-19 $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_216 N_A0_c_254_n N_Y_c_411_n 0.0137249f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_217 N_A0_c_257_n N_Y_c_412_n 0.00356932f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_218 N_A0_c_254_n N_Y_c_412_n 0.0116026f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_219 N_A0_M1000_g N_Y_c_409_n 0.00195709f $X=2.25 $Y=2.775 $X2=0 $Y2=0
cc_220 N_A0_c_257_n N_Y_c_409_n 0.00308377f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_221 N_A0_c_254_n N_Y_c_409_n 0.0469313f $X=2.195 $Y=1.9 $X2=0 $Y2=0
cc_222 N_A0_c_255_n N_Y_c_409_n 0.0475535f $X=2.195 $Y=1.095 $X2=0 $Y2=0
cc_223 N_A0_c_252_n N_Y_c_430_n 0.00309246f $X=1.625 $Y=0.935 $X2=0 $Y2=0
cc_224 N_A0_c_255_n N_Y_c_430_n 0.0518046f $X=2.195 $Y=1.095 $X2=0 $Y2=0
cc_225 N_A0_c_252_n N_VGND_c_465_n 9.42494e-19 $X=1.625 $Y=0.935 $X2=0 $Y2=0
cc_226 N_A0_c_253_n N_VGND_c_465_n 0.0058025f $X=1.625 $Y=0.77 $X2=0 $Y2=0
cc_227 N_A0_c_252_n N_VGND_c_467_n 0.0011812f $X=1.625 $Y=0.935 $X2=0 $Y2=0
cc_228 N_A0_c_253_n N_VGND_c_467_n 0.00666353f $X=1.625 $Y=0.77 $X2=0 $Y2=0
cc_229 N_A0_c_255_n N_VGND_c_467_n 0.00781162f $X=2.195 $Y=1.095 $X2=0 $Y2=0
cc_230 N_A1_M1009_g N_VPWR_c_366_n 0.00357877f $X=1.745 $Y=2.775 $X2=0 $Y2=0
cc_231 N_A1_M1009_g N_VPWR_c_362_n 0.00546467f $X=1.745 $Y=2.775 $X2=0 $Y2=0
cc_232 N_A1_M1009_g N_Y_c_410_n 0.00107829f $X=1.745 $Y=2.775 $X2=0 $Y2=0
cc_233 N_A1_M1009_g N_Y_c_412_n 0.00165185f $X=1.745 $Y=2.775 $X2=0 $Y2=0
cc_234 N_A1_c_311_n N_Y_c_412_n 0.00408181f $X=2.03 $Y=1.42 $X2=0 $Y2=0
cc_235 A1 N_Y_c_412_n 0.00110226f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_236 N_A1_c_311_n N_Y_c_409_n 2.62802e-19 $X=2.03 $Y=1.42 $X2=0 $Y2=0
cc_237 N_A1_M1005_g N_Y_c_409_n 0.00201886f $X=2.105 $Y=0.45 $X2=0 $Y2=0
cc_238 N_A1_M1005_g N_Y_c_430_n 0.0172168f $X=2.105 $Y=0.45 $X2=0 $Y2=0
cc_239 N_A1_M1005_g N_VGND_c_465_n 0.00360655f $X=2.105 $Y=0.45 $X2=0 $Y2=0
cc_240 N_A1_M1005_g N_VGND_c_467_n 0.00563499f $X=2.105 $Y=0.45 $X2=0 $Y2=0
cc_241 N_VPWR_c_362_n A_292_491# 0.00203663f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_242 N_VPWR_c_362_n N_Y_M1009_d 0.00285503f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_243 N_VPWR_c_362_n A_465_491# 0.00238596f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_244 N_Y_c_409_n N_VGND_M1003_d 7.24956e-19 $X=2.615 $Y=2.165 $X2=0 $Y2=0
cc_245 N_Y_c_430_n N_VGND_M1003_d 0.00555035f $X=2.53 $Y=0.462 $X2=0 $Y2=0
cc_246 N_Y_c_430_n N_VGND_c_464_n 0.0276755f $X=2.53 $Y=0.462 $X2=0 $Y2=0
cc_247 N_Y_c_430_n N_VGND_c_465_n 0.0518405f $X=2.53 $Y=0.462 $X2=0 $Y2=0
cc_248 N_Y_M1008_d N_VGND_c_467_n 0.00371499f $X=1.61 $Y=0.24 $X2=0 $Y2=0
cc_249 N_Y_c_430_n N_VGND_c_467_n 0.0378205f $X=2.53 $Y=0.462 $X2=0 $Y2=0
cc_250 N_Y_c_430_n A_436_48# 0.00263191f $X=2.53 $Y=0.462 $X2=-0.19 $Y2=-0.245
cc_251 N_VGND_c_467_n A_244_48# 0.010279f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_252 N_VGND_c_467_n A_436_48# 0.00194182f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
