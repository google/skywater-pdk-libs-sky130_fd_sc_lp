* File: sky130_fd_sc_lp__a21oi_4.pxi.spice
* Created: Fri Aug 28 09:51:51 2020
* 
x_PM_SKY130_FD_SC_LP__A21OI_4%A2 N_A2_M1000_g N_A2_M1008_g N_A2_M1007_g
+ N_A2_M1018_g N_A2_M1012_g N_A2_M1020_g N_A2_M1016_g N_A2_M1022_g N_A2_c_99_n
+ N_A2_c_100_n N_A2_c_101_n A2 A2 A2 A2 N_A2_c_103_n N_A2_c_104_n
+ PM_SKY130_FD_SC_LP__A21OI_4%A2
x_PM_SKY130_FD_SC_LP__A21OI_4%A1 N_A1_c_202_n N_A1_M1004_g N_A1_M1001_g
+ N_A1_c_204_n N_A1_M1005_g N_A1_M1003_g N_A1_c_206_n N_A1_M1013_g N_A1_M1015_g
+ N_A1_c_208_n N_A1_M1023_g N_A1_M1017_g A1 A1 A1 N_A1_c_211_n
+ PM_SKY130_FD_SC_LP__A21OI_4%A1
x_PM_SKY130_FD_SC_LP__A21OI_4%B1 N_B1_M1009_g N_B1_M1002_g N_B1_M1010_g
+ N_B1_M1006_g N_B1_M1014_g N_B1_M1011_g N_B1_M1021_g N_B1_M1019_g B1 B1 B1
+ N_B1_c_283_n N_B1_c_284_n PM_SKY130_FD_SC_LP__A21OI_4%B1
x_PM_SKY130_FD_SC_LP__A21OI_4%A_28_367# N_A_28_367#_M1008_d N_A_28_367#_M1018_d
+ N_A_28_367#_M1001_s N_A_28_367#_M1015_s N_A_28_367#_M1022_d
+ N_A_28_367#_M1006_d N_A_28_367#_M1019_d N_A_28_367#_c_354_n
+ N_A_28_367#_c_355_n N_A_28_367#_c_360_n N_A_28_367#_c_394_p
+ N_A_28_367#_c_364_n N_A_28_367#_c_395_p N_A_28_367#_c_366_n
+ N_A_28_367#_c_392_p N_A_28_367#_c_367_n N_A_28_367#_c_371_n
+ N_A_28_367#_c_397_p N_A_28_367#_c_381_n N_A_28_367#_c_419_p
+ N_A_28_367#_c_356_n N_A_28_367#_c_357_n N_A_28_367#_c_373_n
+ N_A_28_367#_c_375_n N_A_28_367#_c_376_n N_A_28_367#_c_400_p
+ PM_SKY130_FD_SC_LP__A21OI_4%A_28_367#
x_PM_SKY130_FD_SC_LP__A21OI_4%VPWR N_VPWR_M1008_s N_VPWR_M1020_s N_VPWR_M1003_d
+ N_VPWR_M1017_d N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_429_n
+ N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n
+ VPWR N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_425_n N_VPWR_c_438_n
+ N_VPWR_c_439_n PM_SKY130_FD_SC_LP__A21OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A21OI_4%Y N_Y_M1004_s N_Y_M1013_s N_Y_M1009_d N_Y_M1014_d
+ N_Y_M1002_s N_Y_M1011_s N_Y_c_570_p N_Y_c_511_n N_Y_c_531_n N_Y_c_535_n
+ N_Y_c_512_n N_Y_c_539_n N_Y_c_513_n N_Y_c_543_n N_Y_c_545_n N_Y_c_514_n Y Y Y
+ Y Y N_Y_c_517_n PM_SKY130_FD_SC_LP__A21OI_4%Y
x_PM_SKY130_FD_SC_LP__A21OI_4%VGND N_VGND_M1000_s N_VGND_M1007_s N_VGND_M1016_s
+ N_VGND_M1010_s N_VGND_M1021_s N_VGND_c_584_n N_VGND_c_585_n N_VGND_c_586_n
+ N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n VGND
+ N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n
+ N_VGND_c_596_n N_VGND_c_597_n N_VGND_c_598_n PM_SKY130_FD_SC_LP__A21OI_4%VGND
x_PM_SKY130_FD_SC_LP__A21OI_4%A_111_47# N_A_111_47#_M1000_d N_A_111_47#_M1012_d
+ N_A_111_47#_M1005_d N_A_111_47#_M1023_d N_A_111_47#_c_689_n
+ N_A_111_47#_c_666_n N_A_111_47#_c_667_n N_A_111_47#_c_694_n
+ N_A_111_47#_c_676_n PM_SKY130_FD_SC_LP__A21OI_4%A_111_47#
cc_1 VNB N_A2_M1000_g 0.0303725f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_2 VNB N_A2_M1008_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_3 VNB N_A2_M1007_g 0.0204793f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.655
cc_4 VNB N_A2_M1018_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_5 VNB N_A2_M1012_g 0.0206922f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.655
cc_6 VNB N_A2_M1020_g 0.00123444f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=2.465
cc_7 VNB N_A2_M1016_g 0.0256739f $X=-0.19 $Y=-0.245 $X2=3.49 $Y2=0.655
cc_8 VNB N_A2_c_99_n 0.0014593f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.51
cc_9 VNB N_A2_c_100_n 0.0259373f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.51
cc_10 VNB N_A2_c_101_n 0.0102309f $X=-0.19 $Y=-0.245 $X2=3.4 $Y2=1.7
cc_11 VNB A2 0.00256003f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_12 VNB N_A2_c_103_n 0.0920601f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.46
cc_13 VNB N_A2_c_104_n 0.0123312f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.58
cc_14 VNB N_A1_c_202_n 0.0164056f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.295
cc_15 VNB N_A1_M1001_g 0.00614581f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_16 VNB N_A1_c_204_n 0.0162004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_M1003_g 0.00671581f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.625
cc_18 VNB N_A1_c_206_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_19 VNB N_A1_M1015_g 0.00674202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_208_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=2.465
cc_21 VNB N_A1_M1017_g 0.00650228f $X=-0.19 $Y=-0.245 $X2=3.49 $Y2=0.655
cc_22 VNB A1 0.00396162f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_23 VNB N_A1_c_211_n 0.0744481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_M1009_g 0.0251491f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_25 VNB N_B1_M1010_g 0.0227f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.655
cc_26 VNB N_B1_M1014_g 0.0226795f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.655
cc_27 VNB N_B1_M1021_g 0.0279431f $X=-0.19 $Y=-0.245 $X2=3.49 $Y2=0.655
cc_28 VNB N_B1_c_283_n 0.00153206f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_29 VNB N_B1_c_284_n 0.0658776f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_30 VNB N_VPWR_c_425_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_31 VNB N_Y_c_511_n 0.0090711f $X=-0.19 $Y=-0.245 $X2=3.49 $Y2=1.345
cc_32 VNB N_Y_c_512_n 0.0131112f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.51
cc_33 VNB N_Y_c_513_n 0.0185189f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_Y_c_514_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB Y 0.00351834f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_36 VNB N_VGND_c_584_n 0.0109689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_585_n 0.0396934f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.655
cc_38 VNB N_VGND_c_586_n 4.06069e-19 $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=2.465
cc_39 VNB N_VGND_c_587_n 4.02668e-19 $X=-0.19 $Y=-0.245 $X2=3.49 $Y2=0.655
cc_40 VNB N_VGND_c_588_n 3.12649e-19 $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_41 VNB N_VGND_c_589_n 0.0114821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_590_n 0.0304238f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.51
cc_43 VNB N_VGND_c_591_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=3.4 $Y2=1.7
cc_44 VNB N_VGND_c_592_n 0.0515154f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_45 VNB N_VGND_c_593_n 0.0134822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_594_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.46
cc_47 VNB N_VGND_c_595_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_596_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.675
cc_49 VNB N_VGND_c_597_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_598_n 0.288746f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_51 VNB N_A_111_47#_c_666_n 0.00624544f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.295
cc_52 VNB N_A_111_47#_c_667_n 0.00352813f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.655
cc_53 VPB N_A2_M1008_g 0.024677f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_54 VPB N_A2_M1018_g 0.0185384f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_55 VPB N_A2_M1020_g 0.0186439f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=2.465
cc_56 VPB N_A2_M1022_g 0.0185582f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.465
cc_57 VPB N_A2_c_99_n 0.00219237f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=1.51
cc_58 VPB N_A2_c_100_n 0.00632276f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=1.51
cc_59 VPB N_A2_c_101_n 0.0103483f $X=-0.19 $Y=1.655 $X2=3.4 $Y2=1.7
cc_60 VPB A2 0.00125916f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_61 VPB N_A2_c_104_n 0.0146101f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=1.58
cc_62 VPB N_A1_M1001_g 0.0186439f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_63 VPB N_A1_M1003_g 0.0185384f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.625
cc_64 VPB N_A1_M1015_g 0.0185384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A1_M1017_g 0.0190283f $X=-0.19 $Y=1.655 $X2=3.49 $Y2=0.655
cc_66 VPB N_B1_M1002_g 0.0182176f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_67 VPB N_B1_M1006_g 0.0180539f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_68 VPB N_B1_M1011_g 0.0180517f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=2.465
cc_69 VPB N_B1_M1019_g 0.0216874f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.465
cc_70 VPB N_B1_c_283_n 0.00906084f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_71 VPB N_B1_c_284_n 0.0123406f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_72 VPB N_A_28_367#_c_354_n 0.00761272f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=2.465
cc_73 VPB N_A_28_367#_c_355_n 0.035973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_28_367#_c_356_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_75 VPB N_A_28_367#_c_357_n 0.0259042f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.46
cc_76 VPB N_VPWR_c_426_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_77 VPB N_VPWR_c_427_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.34 $Y2=0.655
cc_78 VPB N_VPWR_c_428_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.34 $Y2=2.465
cc_79 VPB N_VPWR_c_429_n 0.0129398f $X=-0.19 $Y=1.655 $X2=3.49 $Y2=1.345
cc_80 VPB N_VPWR_c_430_n 0.00274151f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=1.675
cc_81 VPB N_VPWR_c_431_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_432_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.537 $Y2=1.51
cc_83 VPB N_VPWR_c_433_n 0.0130339f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=1.51
cc_84 VPB N_VPWR_c_434_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=1.51
cc_85 VPB N_VPWR_c_435_n 0.0155214f $X=-0.19 $Y=1.655 $X2=3.4 $Y2=1.7
cc_86 VPB N_VPWR_c_436_n 0.0564562f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_87 VPB N_VPWR_c_425_n 0.0466438f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_88 VPB N_VPWR_c_438_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.46
cc_89 VPB N_VPWR_c_439_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_Y_c_513_n 0.00833994f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_91 N_A2_M1012_g N_A1_c_202_n 0.0209432f $X=1.34 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_92 N_A2_M1020_g N_A1_M1001_g 0.0398563f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_93 N_A2_c_101_n N_A1_M1001_g 0.00739945f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_94 A2 N_A1_M1001_g 0.00736792f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A2_c_101_n N_A1_M1003_g 0.0105539f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_96 A2 N_A1_M1003_g 5.21391e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A2_c_101_n N_A1_M1015_g 0.0105237f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_98 N_A2_M1016_g N_A1_c_208_n 0.0402569f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_99 N_A2_M1022_g N_A1_M1017_g 0.0317159f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A2_c_101_n N_A1_M1017_g 0.0102447f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_101 N_A2_M1012_g A1 3.33455e-19 $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_102 N_A2_M1016_g A1 0.00389254f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_103 N_A2_c_99_n A1 0.00741264f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A2_c_100_n A1 6.09783e-19 $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A2_c_101_n A1 0.0867491f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_106 A2 A1 0.00413847f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A2_c_103_n A1 3.84525e-19 $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_108 N_A2_c_99_n N_A1_c_211_n 0.00122077f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A2_c_100_n N_A1_c_211_n 0.0217117f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_110 N_A2_c_101_n N_A1_c_211_n 0.00753294f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_111 A2 N_A1_c_211_n 0.0109365f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A2_c_103_n N_A1_c_211_n 0.0193661f $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_113 N_A2_M1016_g N_B1_M1009_g 0.033074f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_114 N_A2_M1022_g N_B1_M1002_g 0.0191497f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A2_c_99_n N_B1_M1002_g 8.62125e-19 $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_116 N_A2_c_99_n N_B1_c_283_n 0.0224433f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_117 N_A2_c_100_n N_B1_c_283_n 8.65452e-19 $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A2_c_99_n N_B1_c_284_n 9.36698e-19 $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_119 N_A2_c_100_n N_B1_c_284_n 0.0215144f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_120 N_A2_c_103_n N_A_28_367#_c_354_n 0.00135497f $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_121 N_A2_c_104_n N_A_28_367#_c_354_n 0.021985f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_122 N_A2_M1008_g N_A_28_367#_c_360_n 0.0122595f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A2_M1018_g N_A_28_367#_c_360_n 0.0122595f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A2_c_103_n N_A_28_367#_c_360_n 4.78473e-19 $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_125 N_A2_c_104_n N_A_28_367#_c_360_n 0.0436835f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A2_M1020_g N_A_28_367#_c_364_n 0.0122129f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A2_c_104_n N_A_28_367#_c_364_n 0.0433494f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A2_c_101_n N_A_28_367#_c_366_n 0.0402256f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_129 N_A2_M1022_g N_A_28_367#_c_367_n 0.0131658f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A2_c_99_n N_A_28_367#_c_367_n 0.0135654f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A2_c_100_n N_A_28_367#_c_367_n 2.89632e-19 $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A2_c_101_n N_A_28_367#_c_367_n 0.029286f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_133 N_A2_c_99_n N_A_28_367#_c_371_n 0.00334932f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A2_c_100_n N_A_28_367#_c_371_n 2.57653e-19 $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A2_c_103_n N_A_28_367#_c_373_n 5.41908e-19 $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_136 N_A2_c_104_n N_A_28_367#_c_373_n 0.0156591f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A2_c_101_n N_A_28_367#_c_375_n 0.0142558f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_138 N_A2_c_101_n N_A_28_367#_c_376_n 0.0146339f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_139 N_A2_M1008_g N_VPWR_c_426_n 0.0158744f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A2_M1018_g N_VPWR_c_426_n 0.0140037f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A2_M1020_g N_VPWR_c_426_n 6.7059e-19 $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A2_M1018_g N_VPWR_c_427_n 6.7059e-19 $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A2_M1020_g N_VPWR_c_427_n 0.0139264f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A2_M1022_g N_VPWR_c_430_n 0.00397891f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A2_M1018_g N_VPWR_c_431_n 0.00486043f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A2_M1020_g N_VPWR_c_431_n 0.00486043f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A2_M1008_g N_VPWR_c_435_n 0.00486043f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A2_M1022_g N_VPWR_c_436_n 0.00585385f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A2_M1008_g N_VPWR_c_425_n 0.00918457f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A2_M1018_g N_VPWR_c_425_n 0.00824727f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A2_M1020_g N_VPWR_c_425_n 0.00824727f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A2_M1022_g N_VPWR_c_425_n 0.0106804f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A2_M1016_g N_Y_c_517_n 0.0144245f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_154 N_A2_c_99_n N_Y_c_517_n 0.0110112f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A2_c_100_n N_Y_c_517_n 0.0015512f $X=3.51 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A2_c_101_n N_Y_c_517_n 0.00817279f $X=3.4 $Y=1.7 $X2=0 $Y2=0
cc_157 N_A2_M1000_g N_VGND_c_585_n 0.00702716f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_158 N_A2_c_103_n N_VGND_c_585_n 0.00685402f $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_159 N_A2_c_104_n N_VGND_c_585_n 0.0167558f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A2_M1000_g N_VGND_c_586_n 6.3872e-19 $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A2_M1007_g N_VGND_c_586_n 0.0106924f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A2_M1012_g N_VGND_c_586_n 0.0117685f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A2_M1016_g N_VGND_c_587_n 0.00952448f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A2_M1000_g N_VGND_c_591_n 0.00585385f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_165 N_A2_M1007_g N_VGND_c_591_n 0.00486043f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A2_M1012_g N_VGND_c_592_n 0.00486043f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_167 N_A2_M1016_g N_VGND_c_592_n 0.00564095f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A2_M1000_g N_VGND_c_598_n 0.0114734f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A2_M1007_g N_VGND_c_598_n 0.00824727f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A2_M1012_g N_VGND_c_598_n 0.0082726f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_171 N_A2_M1016_g N_VGND_c_598_n 0.00524073f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_172 N_A2_M1007_g N_A_111_47#_c_666_n 0.0135173f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_173 N_A2_M1012_g N_A_111_47#_c_666_n 0.013425f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A2_c_103_n N_A_111_47#_c_666_n 0.00345061f $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_175 N_A2_c_104_n N_A_111_47#_c_666_n 0.0670587f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A2_M1000_g N_A_111_47#_c_667_n 0.00387885f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A2_c_103_n N_A_111_47#_c_667_n 0.00256759f $X=1.34 $Y=1.46 $X2=0 $Y2=0
cc_178 N_A2_c_104_n N_A_111_47#_c_667_n 0.0196911f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A1_M1001_g N_A_28_367#_c_364_n 0.0122129f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1003_g N_A_28_367#_c_366_n 0.0122595f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A1_M1015_g N_A_28_367#_c_366_n 0.0122595f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A1_M1017_g N_A_28_367#_c_367_n 0.012438f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A1_M1001_g N_VPWR_c_427_n 0.0141056f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A1_M1003_g N_VPWR_c_427_n 6.82688e-19 $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A1_M1001_g N_VPWR_c_428_n 6.7059e-19 $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A1_M1003_g N_VPWR_c_428_n 0.0140037f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A1_M1015_g N_VPWR_c_428_n 0.0140037f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A1_M1017_g N_VPWR_c_428_n 6.7059e-19 $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A1_M1015_g N_VPWR_c_429_n 0.00486043f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A1_M1017_g N_VPWR_c_429_n 0.00486043f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A1_M1015_g N_VPWR_c_430_n 6.7059e-19 $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A1_M1017_g N_VPWR_c_430_n 0.0138443f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A1_M1001_g N_VPWR_c_433_n 0.00486043f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A1_M1003_g N_VPWR_c_433_n 0.00486043f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A1_M1001_g N_VPWR_c_425_n 0.00824727f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A1_M1003_g N_VPWR_c_425_n 0.00824727f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A1_M1015_g N_VPWR_c_425_n 0.00824727f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A1_M1017_g N_VPWR_c_425_n 0.00824727f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A1_c_202_n N_Y_c_517_n 0.00310434f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_200 N_A1_c_204_n N_Y_c_517_n 0.00957371f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_201 N_A1_c_206_n N_Y_c_517_n 0.00957371f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_202 N_A1_c_208_n N_Y_c_517_n 0.00951606f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_203 A1 N_Y_c_517_n 0.0780805f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_204 N_A1_c_211_n N_Y_c_517_n 0.00706127f $X=3.06 $Y=1.35 $X2=0 $Y2=0
cc_205 N_A1_c_202_n N_VGND_c_586_n 0.00127727f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_206 N_A1_c_208_n N_VGND_c_587_n 0.00120867f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_207 N_A1_c_202_n N_VGND_c_592_n 0.00357877f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_208 N_A1_c_204_n N_VGND_c_592_n 0.00357877f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_209 N_A1_c_206_n N_VGND_c_592_n 0.00357877f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_210 N_A1_c_208_n N_VGND_c_592_n 0.00357877f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_211 N_A1_c_202_n N_VGND_c_598_n 0.00537654f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_212 N_A1_c_204_n N_VGND_c_598_n 0.00542194f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_213 N_A1_c_206_n N_VGND_c_598_n 0.00542194f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_214 N_A1_c_208_n N_VGND_c_598_n 0.00544922f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_215 N_A1_c_202_n N_A_111_47#_c_666_n 0.00416967f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A1_c_202_n N_A_111_47#_c_676_n 0.0178975f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_217 N_A1_c_204_n N_A_111_47#_c_676_n 0.0135994f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_218 N_A1_c_206_n N_A_111_47#_c_676_n 0.0135994f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_219 N_A1_c_208_n N_A_111_47#_c_676_n 0.0136458f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_220 N_B1_M1002_g N_A_28_367#_c_381_n 0.012237f $X=3.96 $Y=2.465 $X2=0 $Y2=0
cc_221 N_B1_M1006_g N_A_28_367#_c_381_n 0.0121905f $X=4.39 $Y=2.465 $X2=0 $Y2=0
cc_222 N_B1_M1011_g N_A_28_367#_c_356_n 0.012237f $X=4.82 $Y=2.465 $X2=0 $Y2=0
cc_223 N_B1_M1019_g N_A_28_367#_c_356_n 0.012237f $X=5.25 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B1_M1002_g N_VPWR_c_436_n 0.00357877f $X=3.96 $Y=2.465 $X2=0 $Y2=0
cc_225 N_B1_M1006_g N_VPWR_c_436_n 0.00357877f $X=4.39 $Y=2.465 $X2=0 $Y2=0
cc_226 N_B1_M1011_g N_VPWR_c_436_n 0.00357877f $X=4.82 $Y=2.465 $X2=0 $Y2=0
cc_227 N_B1_M1019_g N_VPWR_c_436_n 0.00357877f $X=5.25 $Y=2.465 $X2=0 $Y2=0
cc_228 N_B1_M1002_g N_VPWR_c_425_n 0.00537654f $X=3.96 $Y=2.465 $X2=0 $Y2=0
cc_229 N_B1_M1006_g N_VPWR_c_425_n 0.0053512f $X=4.39 $Y=2.465 $X2=0 $Y2=0
cc_230 N_B1_M1011_g N_VPWR_c_425_n 0.0053512f $X=4.82 $Y=2.465 $X2=0 $Y2=0
cc_231 N_B1_M1019_g N_VPWR_c_425_n 0.00631529f $X=5.25 $Y=2.465 $X2=0 $Y2=0
cc_232 N_B1_M1010_g N_Y_c_511_n 0.0139219f $X=4.39 $Y=0.655 $X2=0 $Y2=0
cc_233 N_B1_M1014_g N_Y_c_511_n 0.0142467f $X=4.82 $Y=0.655 $X2=0 $Y2=0
cc_234 N_B1_c_283_n N_Y_c_511_n 0.0499706f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_235 N_B1_c_284_n N_Y_c_511_n 0.00246472f $X=5.25 $Y=1.51 $X2=0 $Y2=0
cc_236 N_B1_M1006_g N_Y_c_531_n 0.0129934f $X=4.39 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1011_g N_Y_c_531_n 0.0129469f $X=4.82 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_c_283_n N_Y_c_531_n 0.0405553f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_239 N_B1_c_284_n N_Y_c_531_n 5.64665e-19 $X=5.25 $Y=1.51 $X2=0 $Y2=0
cc_240 N_B1_M1014_g N_Y_c_535_n 7.21728e-19 $X=4.82 $Y=0.655 $X2=0 $Y2=0
cc_241 N_B1_M1021_g N_Y_c_535_n 7.21728e-19 $X=5.25 $Y=0.655 $X2=0 $Y2=0
cc_242 N_B1_M1021_g N_Y_c_512_n 0.0169425f $X=5.25 $Y=0.655 $X2=0 $Y2=0
cc_243 N_B1_c_283_n N_Y_c_512_n 0.00763896f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_244 N_B1_M1019_g N_Y_c_539_n 0.0155962f $X=5.25 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_c_283_n N_Y_c_539_n 0.00509065f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_246 N_B1_M1021_g N_Y_c_513_n 0.0223553f $X=5.25 $Y=0.655 $X2=0 $Y2=0
cc_247 N_B1_c_283_n N_Y_c_513_n 0.0254362f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_248 N_B1_c_283_n N_Y_c_543_n 0.0175073f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_249 N_B1_c_284_n N_Y_c_543_n 6.37898e-19 $X=5.25 $Y=1.51 $X2=0 $Y2=0
cc_250 N_B1_c_283_n N_Y_c_545_n 0.0177168f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_251 N_B1_c_284_n N_Y_c_545_n 6.37898e-19 $X=5.25 $Y=1.51 $X2=0 $Y2=0
cc_252 N_B1_c_283_n N_Y_c_514_n 0.0160407f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_253 N_B1_c_284_n N_Y_c_514_n 0.00256759f $X=5.25 $Y=1.51 $X2=0 $Y2=0
cc_254 N_B1_M1009_g Y 0.00574401f $X=3.96 $Y=0.655 $X2=0 $Y2=0
cc_255 N_B1_M1010_g Y 2.24321e-19 $X=4.39 $Y=0.655 $X2=0 $Y2=0
cc_256 N_B1_c_283_n Y 0.0160407f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_257 N_B1_c_284_n Y 0.00256759f $X=5.25 $Y=1.51 $X2=0 $Y2=0
cc_258 N_B1_M1009_g N_Y_c_517_n 0.0123205f $X=3.96 $Y=0.655 $X2=0 $Y2=0
cc_259 N_B1_c_283_n N_Y_c_517_n 0.00598343f $X=5.07 $Y=1.51 $X2=0 $Y2=0
cc_260 N_B1_M1009_g N_VGND_c_587_n 0.00822115f $X=3.96 $Y=0.655 $X2=0 $Y2=0
cc_261 N_B1_M1010_g N_VGND_c_587_n 5.41941e-19 $X=4.39 $Y=0.655 $X2=0 $Y2=0
cc_262 N_B1_M1009_g N_VGND_c_588_n 6.26989e-19 $X=3.96 $Y=0.655 $X2=0 $Y2=0
cc_263 N_B1_M1010_g N_VGND_c_588_n 0.0118954f $X=4.39 $Y=0.655 $X2=0 $Y2=0
cc_264 N_B1_M1014_g N_VGND_c_588_n 0.0117077f $X=4.82 $Y=0.655 $X2=0 $Y2=0
cc_265 N_B1_M1021_g N_VGND_c_588_n 6.36641e-19 $X=5.25 $Y=0.655 $X2=0 $Y2=0
cc_266 N_B1_M1014_g N_VGND_c_590_n 6.36641e-19 $X=4.82 $Y=0.655 $X2=0 $Y2=0
cc_267 N_B1_M1021_g N_VGND_c_590_n 0.0132658f $X=5.25 $Y=0.655 $X2=0 $Y2=0
cc_268 N_B1_M1009_g N_VGND_c_593_n 0.00564095f $X=3.96 $Y=0.655 $X2=0 $Y2=0
cc_269 N_B1_M1010_g N_VGND_c_593_n 0.00486043f $X=4.39 $Y=0.655 $X2=0 $Y2=0
cc_270 N_B1_M1014_g N_VGND_c_594_n 0.00486043f $X=4.82 $Y=0.655 $X2=0 $Y2=0
cc_271 N_B1_M1021_g N_VGND_c_594_n 0.00486043f $X=5.25 $Y=0.655 $X2=0 $Y2=0
cc_272 N_B1_M1009_g N_VGND_c_598_n 0.00513564f $X=3.96 $Y=0.655 $X2=0 $Y2=0
cc_273 N_B1_M1010_g N_VGND_c_598_n 0.00824727f $X=4.39 $Y=0.655 $X2=0 $Y2=0
cc_274 N_B1_M1014_g N_VGND_c_598_n 0.00824727f $X=4.82 $Y=0.655 $X2=0 $Y2=0
cc_275 N_B1_M1021_g N_VGND_c_598_n 0.00824727f $X=5.25 $Y=0.655 $X2=0 $Y2=0
cc_276 N_A_28_367#_c_360_n N_VPWR_M1008_s 0.0033582f $X=1.03 $Y=2.04 $X2=-0.19
+ $Y2=1.655
cc_277 N_A_28_367#_c_364_n N_VPWR_M1020_s 0.00353353f $X=1.9 $Y=2.04 $X2=0 $Y2=0
cc_278 N_A_28_367#_c_366_n N_VPWR_M1003_d 0.00339614f $X=2.75 $Y=2.04 $X2=0
+ $Y2=0
cc_279 N_A_28_367#_c_367_n N_VPWR_M1017_d 0.00428266f $X=3.61 $Y=2.04 $X2=0
+ $Y2=0
cc_280 N_A_28_367#_c_360_n N_VPWR_c_426_n 0.0170777f $X=1.03 $Y=2.04 $X2=0 $Y2=0
cc_281 N_A_28_367#_c_364_n N_VPWR_c_427_n 0.0170777f $X=1.9 $Y=2.04 $X2=0 $Y2=0
cc_282 N_A_28_367#_c_366_n N_VPWR_c_428_n 0.0170777f $X=2.75 $Y=2.04 $X2=0 $Y2=0
cc_283 N_A_28_367#_c_392_p N_VPWR_c_429_n 0.0124525f $X=2.845 $Y=2.91 $X2=0
+ $Y2=0
cc_284 N_A_28_367#_c_367_n N_VPWR_c_430_n 0.0185459f $X=3.61 $Y=2.04 $X2=0 $Y2=0
cc_285 N_A_28_367#_c_394_p N_VPWR_c_431_n 0.0124525f $X=1.125 $Y=2.91 $X2=0
+ $Y2=0
cc_286 N_A_28_367#_c_395_p N_VPWR_c_433_n 0.0120977f $X=1.985 $Y=2.91 $X2=0
+ $Y2=0
cc_287 N_A_28_367#_c_355_n N_VPWR_c_435_n 0.0178111f $X=0.265 $Y=2.91 $X2=0
+ $Y2=0
cc_288 N_A_28_367#_c_397_p N_VPWR_c_436_n 0.0155393f $X=3.747 $Y=2.905 $X2=0
+ $Y2=0
cc_289 N_A_28_367#_c_381_n N_VPWR_c_436_n 0.0329427f $X=4.465 $Y=2.99 $X2=0
+ $Y2=0
cc_290 N_A_28_367#_c_356_n N_VPWR_c_436_n 0.052634f $X=5.325 $Y=2.99 $X2=0 $Y2=0
cc_291 N_A_28_367#_c_400_p N_VPWR_c_436_n 0.0155393f $X=4.602 $Y=2.99 $X2=0
+ $Y2=0
cc_292 N_A_28_367#_M1008_d N_VPWR_c_425_n 0.00371702f $X=0.14 $Y=1.835 $X2=0
+ $Y2=0
cc_293 N_A_28_367#_M1018_d N_VPWR_c_425_n 0.00536646f $X=0.985 $Y=1.835 $X2=0
+ $Y2=0
cc_294 N_A_28_367#_M1001_s N_VPWR_c_425_n 0.00571434f $X=1.845 $Y=1.835 $X2=0
+ $Y2=0
cc_295 N_A_28_367#_M1015_s N_VPWR_c_425_n 0.00536646f $X=2.705 $Y=1.835 $X2=0
+ $Y2=0
cc_296 N_A_28_367#_M1022_d N_VPWR_c_425_n 0.00220342f $X=3.605 $Y=1.835 $X2=0
+ $Y2=0
cc_297 N_A_28_367#_M1006_d N_VPWR_c_425_n 0.00220342f $X=4.465 $Y=1.835 $X2=0
+ $Y2=0
cc_298 N_A_28_367#_M1019_d N_VPWR_c_425_n 0.00215158f $X=5.325 $Y=1.835 $X2=0
+ $Y2=0
cc_299 N_A_28_367#_c_355_n N_VPWR_c_425_n 0.0100304f $X=0.265 $Y=2.91 $X2=0
+ $Y2=0
cc_300 N_A_28_367#_c_394_p N_VPWR_c_425_n 0.00730901f $X=1.125 $Y=2.91 $X2=0
+ $Y2=0
cc_301 N_A_28_367#_c_395_p N_VPWR_c_425_n 0.00691495f $X=1.985 $Y=2.91 $X2=0
+ $Y2=0
cc_302 N_A_28_367#_c_392_p N_VPWR_c_425_n 0.00730901f $X=2.845 $Y=2.91 $X2=0
+ $Y2=0
cc_303 N_A_28_367#_c_397_p N_VPWR_c_425_n 0.0106525f $X=3.747 $Y=2.905 $X2=0
+ $Y2=0
cc_304 N_A_28_367#_c_381_n N_VPWR_c_425_n 0.0203755f $X=4.465 $Y=2.99 $X2=0
+ $Y2=0
cc_305 N_A_28_367#_c_356_n N_VPWR_c_425_n 0.0323406f $X=5.325 $Y=2.99 $X2=0
+ $Y2=0
cc_306 N_A_28_367#_c_400_p N_VPWR_c_425_n 0.0106525f $X=4.602 $Y=2.99 $X2=0
+ $Y2=0
cc_307 N_A_28_367#_c_381_n N_Y_M1002_s 0.00332344f $X=4.465 $Y=2.99 $X2=0 $Y2=0
cc_308 N_A_28_367#_c_356_n N_Y_M1011_s 0.00332344f $X=5.325 $Y=2.99 $X2=0 $Y2=0
cc_309 N_A_28_367#_M1006_d N_Y_c_531_n 0.00333177f $X=4.465 $Y=1.835 $X2=0 $Y2=0
cc_310 N_A_28_367#_c_419_p N_Y_c_531_n 0.0135055f $X=4.605 $Y=2.47 $X2=0 $Y2=0
cc_311 N_A_28_367#_M1019_d N_Y_c_539_n 0.011265f $X=5.325 $Y=1.835 $X2=0 $Y2=0
cc_312 N_A_28_367#_c_357_n N_Y_c_539_n 0.0178857f $X=5.465 $Y=2.47 $X2=0 $Y2=0
cc_313 N_A_28_367#_M1019_d N_Y_c_513_n 0.00504205f $X=5.325 $Y=1.835 $X2=0 $Y2=0
cc_314 N_A_28_367#_c_381_n N_Y_c_543_n 0.0126348f $X=4.465 $Y=2.99 $X2=0 $Y2=0
cc_315 N_A_28_367#_c_356_n N_Y_c_545_n 0.0126348f $X=5.325 $Y=2.99 $X2=0 $Y2=0
cc_316 N_VPWR_c_425_n N_Y_M1002_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_425_n N_Y_M1011_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_318 N_Y_c_517_n N_VGND_M1016_s 0.00879689f $X=4.06 $Y=0.925 $X2=0 $Y2=0
cc_319 N_Y_c_517_n N_VGND_c_587_n 0.017112f $X=4.06 $Y=0.925 $X2=0 $Y2=0
cc_320 N_Y_c_511_n N_VGND_c_588_n 0.0216087f $X=4.94 $Y=1.17 $X2=0 $Y2=0
cc_321 N_Y_c_512_n N_VGND_c_590_n 0.0222601f $X=5.415 $Y=1.17 $X2=0 $Y2=0
cc_322 N_Y_c_570_p N_VGND_c_593_n 0.0128073f $X=4.175 $Y=0.42 $X2=0 $Y2=0
cc_323 N_Y_c_535_n N_VGND_c_594_n 0.0124525f $X=5.035 $Y=0.42 $X2=0 $Y2=0
cc_324 N_Y_M1004_s N_VGND_c_598_n 0.00225186f $X=1.845 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_M1013_s N_VGND_c_598_n 0.00225186f $X=2.705 $Y=0.235 $X2=0 $Y2=0
cc_326 N_Y_M1009_d N_VGND_c_598_n 0.00429287f $X=4.035 $Y=0.235 $X2=0 $Y2=0
cc_327 N_Y_M1014_d N_VGND_c_598_n 0.00536646f $X=4.895 $Y=0.235 $X2=0 $Y2=0
cc_328 N_Y_c_570_p N_VGND_c_598_n 0.0076925f $X=4.175 $Y=0.42 $X2=0 $Y2=0
cc_329 N_Y_c_535_n N_VGND_c_598_n 0.00730901f $X=5.035 $Y=0.42 $X2=0 $Y2=0
cc_330 N_Y_c_517_n N_VGND_c_598_n 0.0138337f $X=4.06 $Y=0.925 $X2=0 $Y2=0
cc_331 N_Y_c_517_n N_A_111_47#_M1005_d 0.00334119f $X=4.06 $Y=0.925 $X2=0 $Y2=0
cc_332 N_Y_c_517_n N_A_111_47#_M1023_d 0.00467463f $X=4.06 $Y=0.925 $X2=0 $Y2=0
cc_333 N_Y_M1004_s N_A_111_47#_c_676_n 0.00334419f $X=1.845 $Y=0.235 $X2=0 $Y2=0
cc_334 N_Y_M1013_s N_A_111_47#_c_676_n 0.00334419f $X=2.705 $Y=0.235 $X2=0 $Y2=0
cc_335 N_Y_c_517_n N_A_111_47#_c_676_n 0.0805471f $X=4.06 $Y=0.925 $X2=0 $Y2=0
cc_336 N_VGND_c_598_n N_A_111_47#_M1000_d 0.00397496f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_337 N_VGND_c_598_n N_A_111_47#_M1012_d 0.00376627f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_338 N_VGND_c_598_n N_A_111_47#_M1005_d 0.00225186f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_c_598_n N_A_111_47#_M1023_d 0.00247351f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_340 N_VGND_c_591_n N_A_111_47#_c_689_n 0.0138717f $X=0.96 $Y=0 $X2=0 $Y2=0
cc_341 N_VGND_c_598_n N_A_111_47#_c_689_n 0.00886411f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_M1007_s N_A_111_47#_c_666_n 0.00176461f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_343 N_VGND_c_586_n N_A_111_47#_c_666_n 0.0170777f $X=1.125 $Y=0.38 $X2=0
+ $Y2=0
cc_344 N_VGND_c_585_n N_A_111_47#_c_667_n 0.00166417f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_345 N_VGND_c_592_n N_A_111_47#_c_694_n 0.0125234f $X=3.56 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_598_n N_A_111_47#_c_694_n 0.00738676f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_347 N_VGND_c_592_n N_A_111_47#_c_676_n 0.0999294f $X=3.56 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_598_n N_A_111_47#_c_676_n 0.0634391f $X=5.52 $Y=0 $X2=0 $Y2=0
