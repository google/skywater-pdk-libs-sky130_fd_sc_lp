* File: sky130_fd_sc_lp__decapkapwr_6.pex.spice
* Created: Wed Sep  2 09:42:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_6%VGND 1 7 10 13 15 16 18 20 24 28 29 42
r30 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r31 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r32 36 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r33 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r35 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r36 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 30 38 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.25
+ $Y2=0
r38 30 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.72
+ $Y2=0
r39 29 41 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.665
+ $Y2=0
r40 29 35 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.16
+ $Y2=0
r41 24 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r42 24 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r43 20 22 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.615 $Y=0.405
+ $X2=2.615 $Y2=1.085
r44 18 41 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.665 $Y2=0
r45 18 20 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.405
r46 16 28 22.4154 $w=1.774e-06 $l=1.03959e-06 $layer=POLY_cond $X=0.915 $Y=1.77
+ $X2=1.4 $Y2=2.595
r47 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.915
+ $Y=1.77 $X2=0.915 $Y2=1.77
r48 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.5 $Y=1.77
+ $X2=0.915 $Y2=1.77
r49 10 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.335 $Y=0.38
+ $X2=0.335 $Y2=1.06
r50 8 13 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.5 $Y2=1.77
r51 8 12 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.335 $Y=1.605
+ $X2=0.335 $Y2=1.06
r52 7 38 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.25 $Y2=0
r53 7 10 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r54 1 22 121.333 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.615 $Y2=1.085
r55 1 20 121.333 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.615 $Y2=0.405
r56 1 12 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=0.335 $Y2=1.06
r57 1 10 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=0.335 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_6%KAPWR 1 7 9 11 13 16 22 24 25 28 36
r34 35 36 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.665 $Y=2.81
+ $X2=2.665 $Y2=2.81
r35 31 32 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.215 $Y=2.81
+ $X2=0.215 $Y2=2.81
r36 25 36 0.669526 $w=2.7e-07 $l=1.225e-06 $layer=MET1_cond $X=1.44 $Y=2.81
+ $X2=2.665 $Y2=2.81
r37 25 32 0.669526 $w=2.7e-07 $l=1.225e-06 $layer=MET1_cond $X=1.44 $Y=2.81
+ $X2=0.215 $Y2=2.81
r38 22 35 3.13952 $w=3.65e-07 $l=2e-07 $layer=LI1_cond $X=2.567 $Y=2.675
+ $X2=2.567 $Y2=2.875
r39 22 24 12.1559 $w=3.63e-07 $l=3.85e-07 $layer=LI1_cond $X=2.567 $Y=2.675
+ $X2=2.567 $Y2=2.29
r40 21 24 19.4179 $w=3.63e-07 $l=6.15e-07 $layer=LI1_cond $X=2.567 $Y=1.675
+ $X2=2.567 $Y2=2.29
r41 16 28 20.7068 $w=1.804e-06 $l=7.75e-07 $layer=POLY_cond $X=1.48 $Y=1.51
+ $X2=1.48 $Y2=0.735
r42 16 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.51 $X2=2.32 $Y2=1.51
r43 15 19 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=1.64 $Y=1.507
+ $X2=2.32 $Y2=1.507
r44 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.64
+ $Y=1.51 $X2=1.64 $Y2=1.51
r45 13 21 6.83279 $w=3.35e-07 $l=2.52389e-07 $layer=LI1_cond $X=2.385 $Y=1.507
+ $X2=2.567 $Y2=1.675
r46 13 19 2.23608 $w=3.33e-07 $l=6.5e-08 $layer=LI1_cond $X=2.385 $Y=1.507
+ $X2=2.32 $Y2=1.507
r47 12 31 3.69365 $w=2.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.425 $Y=2.81
+ $X2=0.26 $Y2=2.875
r48 11 35 3.8773 $w=2.7e-07 $l=2.12024e-07 $layer=LI1_cond $X=2.385 $Y=2.81
+ $X2=2.567 $Y2=2.875
r49 11 12 83.6588 $w=2.68e-07 $l=1.96e-06 $layer=LI1_cond $X=2.385 $Y=2.81
+ $X2=0.425 $Y2=2.81
r50 7 31 3.21187 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=0.26 $Y=2.675 $X2=0.26
+ $Y2=2.875
r51 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.26 $Y=2.675
+ $X2=0.26 $Y2=2.27
r52 1 35 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=2.55 $Y2=2.97
r53 1 31 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=0.26 $Y2=2.95
r54 1 24 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=2.55 $Y2=2.29
r55 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.095 $X2=0.26 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_6%VPWR 1 8 14
r14 5 14 0.00529514 $w=2.88e-06 $l=1.22e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.44 $Y2=3.208
r15 5 8 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33 $X2=2.64
+ $Y2=3.33
r16 4 8 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=2.64
+ $Y2=3.33
r17 4 5 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r18 1 14 4.34028e-05 $w=2.88e-06 $l=1e-09 $layer=MET1_cond $X=1.44 $Y=3.207
+ $X2=1.44 $Y2=3.208
.ends

