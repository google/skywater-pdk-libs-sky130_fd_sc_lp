* File: sky130_fd_sc_lp__nor3_1.pex.spice
* Created: Fri Aug 28 10:55:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3_1%A 3 6 8 9 13 15
c25 8 0 5.98877e-20 $X=0.24 $Y=1.295
r26 13 16 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.377 $Y=1.375
+ $X2=0.377 $Y2=1.54
r27 13 15 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.377 $Y=1.375
+ $X2=0.377 $Y2=1.21
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.375 $X2=0.37 $Y2=1.375
r29 9 14 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.375
r30 8 14 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.375
r31 6 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.54
r32 3 15 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.475 $Y=0.665
+ $X2=0.475 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_1%B 3 7 9 10 11 12 19 20 36
c44 20 0 1.47358e-19 $X=0.925 $Y=1.51
c45 7 0 5.98877e-20 $X=0.935 $Y=2.465
r46 36 37 1.32673 $w=3.83e-07 $l=1.5e-08 $layer=LI1_cond $X=0.817 $Y=1.665
+ $X2=0.817 $Y2=1.68
r47 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.675
r48 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.345
r49 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.51 $X2=0.925 $Y2=1.51
r50 11 12 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.405
+ $X2=0.765 $Y2=2.775
r51 10 11 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.035
+ $X2=0.765 $Y2=2.405
r52 9 36 1.04768 $w=3.83e-07 $l=3.5e-08 $layer=LI1_cond $X=0.817 $Y=1.63
+ $X2=0.817 $Y2=1.665
r53 9 20 3.59203 $w=3.83e-07 $l=1.2e-07 $layer=LI1_cond $X=0.817 $Y=1.63
+ $X2=0.817 $Y2=1.51
r54 9 10 13.1708 $w=2.78e-07 $l=3.2e-07 $layer=LI1_cond $X=0.765 $Y=1.715
+ $X2=0.765 $Y2=2.035
r55 9 37 1.44055 $w=2.78e-07 $l=3.5e-08 $layer=LI1_cond $X=0.765 $Y=1.715
+ $X2=0.765 $Y2=1.68
r56 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.935 $Y=2.465
+ $X2=0.935 $Y2=1.675
r57 3 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.905 $Y=0.665
+ $X2=0.905 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_1%C 3 7 9 14
r27 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.605
+ $Y=1.51 $X2=1.605 $Y2=1.51
r28 11 14 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.375 $Y=1.51
+ $X2=1.605 $Y2=1.51
r29 9 15 7.86588 $w=3.13e-07 $l=2.15e-07 $layer=LI1_cond $X=1.677 $Y=1.295
+ $X2=1.677 $Y2=1.51
r30 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=1.51
r31 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=2.465
r32 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.345
+ $X2=1.375 $Y2=1.51
r33 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.375 $Y=1.345
+ $X2=1.375 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_1%VPWR 1 4 6 10 17 18 28
r23 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r25 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 15 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 14 17 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r28 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 12 21 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r30 12 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 10 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 10 15 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 6 9 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.26 $Y=2.005
+ $X2=0.26 $Y2=2.95
r34 4 21 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r35 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r36 1 9 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r37 1 6 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_1%Y 1 2 3 12 14 15 17 18 20 25 26 27
r46 39 42 11.7045 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=1.265 $Y=2.005
+ $X2=1.59 $Y2=2.005
r47 31 42 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=1.63 $Y=2.005 $X2=1.59
+ $Y2=2.005
r48 27 37 3.79463 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.63 $Y=2.775
+ $X2=1.63 $Y2=2.91
r49 26 27 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=2.405
+ $X2=1.63 $Y2=2.775
r50 26 31 6.74601 $w=4.08e-07 $l=2.4e-07 $layer=LI1_cond $X=1.63 $Y=2.405
+ $X2=1.63 $Y2=2.165
r51 25 31 1.80069 $w=3.18e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=2.005 $X2=1.63
+ $Y2=2.005
r52 18 22 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.615 $Y=0.955
+ $X2=1.265 $Y2=0.955
r53 18 20 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=1.615 $Y=0.87
+ $X2=1.615 $Y2=0.42
r54 17 39 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.265 $Y=1.845
+ $X2=1.265 $Y2=2.005
r55 16 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=1.04
+ $X2=1.265 $Y2=0.955
r56 16 17 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.265 $Y=1.04
+ $X2=1.265 $Y2=1.845
r57 14 22 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.955
+ $X2=1.265 $Y2=0.955
r58 14 15 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.18 $Y=0.955
+ $X2=0.805 $Y2=0.955
r59 10 15 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.7 $Y=0.87
+ $X2=0.805 $Y2=0.955
r60 10 12 23.7662 $w=2.08e-07 $l=4.5e-07 $layer=LI1_cond $X=0.7 $Y=0.87 $X2=0.7
+ $Y2=0.42
r61 3 42 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=1.98
r62 3 37 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=2.91
r63 2 20 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.45
+ $Y=0.245 $X2=1.59 $Y2=0.42
r64 1 12 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.245 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_1%VGND 1 2 7 9 13 15 17 24 25 31 38
r30 31 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r31 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r32 25 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r33 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r34 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r35 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r36 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r37 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r38 18 28 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r39 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r40 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r41 17 20 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r42 15 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r43 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r44 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r45 11 13 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.57
r46 7 28 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r47 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r48 2 13 182 $w=1.7e-07 $l=3.9702e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.245 $X2=1.14 $Y2=0.57
r49 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.39
.ends

