* File: sky130_fd_sc_lp__a211o_2.spice
* Created: Wed Sep  2 09:17:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211o_2.pex.spice"
.subckt sky130_fd_sc_lp__a211o_2  VNB VPB A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 N_X_M1002_d N_A_80_21#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75003
+ A=0.126 P=1.98 MULT=1
MM1004 N_X_M1002_d N_A_80_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.336 PD=1.12 PS=1.64 NRD=0 NRS=49.284 M=1 R=5.6 SA=75000.6
+ SB=75002.6 A=0.126 P=1.98 MULT=1
MM1005 A_386_47# N_A2_M1005_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.336 PD=1.05 PS=1.64 NRD=7.14 NRS=49.284 M=1 R=5.6 SA=75001.6 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1007 N_A_80_21#_M1007_d N_A1_M1007_g A_386_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.21 AS=0.0882 PD=1.34 PS=1.05 NRD=14.28 NRS=7.14 M=1 R=5.6 SA=75001.9
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_B1_M1010_g N_A_80_21#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.21 PD=1.12 PS=1.34 NRD=0 NRS=17.136 M=1 R=5.6 SA=75002.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1001 N_A_80_21#_M1001_d N_C1_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_80_21#_M1011_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A2_M1009_g N_A_303_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.3339 PD=1.65 PS=3.05 NRD=8.5892 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 N_A_303_367#_M1000_d N_A1_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2079 AS=0.2457 PD=1.59 PS=1.65 NRD=2.3443 NRS=8.5892 M=1 R=8.4
+ SA=75000.7 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 A_590_367# N_B1_M1008_g N_A_303_367#_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1701 AS=0.2079 PD=1.53 PS=1.59 NRD=12.4898 NRS=5.4569 M=1 R=8.4
+ SA=75001.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_A_80_21#_M1006_d N_C1_M1006_g A_590_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1701 PD=3.05 PS=1.53 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75001.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a211o_2.pxi.spice"
*
.ends
*
*
