* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrbp_lp D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1028_23# a_778_49# a_1273_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_1614_74# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_455_49# a_272_419# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND GATE a_272_112# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1701_74# a_1028_23# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_778_49# a_455_49# a_955_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_1028_23# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 VPWR a_778_49# a_1028_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VGND a_1614_74# a_1859_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1614_74# a_1028_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_1614_74# a_1028_23# a_1701_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_455_49# a_272_419# a_542_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_944_49# a_1028_23# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR GATE a_272_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VPWR a_27_112# a_692_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_700_49# a_455_49# a_778_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_542_49# a_272_419# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_778_49# a_272_419# a_944_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1273_49# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_1028_23# a_1431_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_692_367# a_272_419# a_778_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 VGND a_27_112# a_700_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_114_112# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1431_49# a_1028_23# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_27_112# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_27_112# D a_114_112# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1859_74# a_1614_74# Q_N VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_272_112# GATE a_272_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR a_1028_23# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X29 a_955_367# a_1028_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
