* File: sky130_fd_sc_lp__o22a_4.pex.spice
* Created: Fri Aug 28 11:09:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22A_4%A_86_23# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 51 52 56 59 60 61 64 71 74 76 87
r148 84 85 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.795 $Y=1.49
+ $X2=2.03 $Y2=1.49
r149 83 84 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.6 $Y=1.49
+ $X2=1.795 $Y2=1.49
r150 82 83 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.365 $Y=1.49
+ $X2=1.6 $Y2=1.49
r151 81 82 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.17 $Y=1.49
+ $X2=1.365 $Y2=1.49
r152 77 79 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.505 $Y=1.49
+ $X2=0.935 $Y2=1.49
r153 70 87 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.3 $Y=1.49
+ $X2=2.46 $Y2=1.49
r154 70 85 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.3 $Y=1.49
+ $X2=2.03 $Y2=1.49
r155 69 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.3 $Y=1.49
+ $X2=2.595 $Y2=1.49
r156 69 70 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.3
+ $Y=1.49 $X2=2.3 $Y2=1.49
r157 65 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.775 $Y=2.015
+ $X2=3.61 $Y2=2.015
r158 64 76 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=2.015
+ $X2=5.48 $Y2=2.015
r159 64 65 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=5.315 $Y=2.015
+ $X2=3.775 $Y2=2.015
r160 60 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=2.015
+ $X2=3.61 $Y2=2.015
r161 60 61 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.445 $Y=2.015
+ $X2=2.68 $Y2=2.015
r162 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.595 $Y=1.93
+ $X2=2.68 $Y2=2.015
r163 58 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.575
+ $X2=2.595 $Y2=1.49
r164 58 59 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.595 $Y=1.575
+ $X2=2.595 $Y2=1.93
r165 54 56 38.1193 $w=2.58e-07 $l=8.6e-07 $layer=LI1_cond $X=3.18 $Y=0.385
+ $X2=4.04 $Y2=0.385
r166 52 54 31.6922 $w=2.58e-07 $l=7.15e-07 $layer=LI1_cond $X=2.465 $Y=0.385
+ $X2=3.18 $Y2=0.385
r167 51 69 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.38 $Y=1.405
+ $X2=2.3 $Y2=1.49
r168 50 52 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.38 $Y=0.515
+ $X2=2.465 $Y2=0.385
r169 50 51 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.38 $Y=0.515
+ $X2=2.38 $Y2=1.405
r170 48 81 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.94 $Y=1.49
+ $X2=1.17 $Y2=1.49
r171 48 79 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.94 $Y=1.49
+ $X2=0.935 $Y2=1.49
r172 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.94
+ $Y=1.49 $X2=0.94 $Y2=1.49
r173 45 69 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.295 $Y=1.49
+ $X2=2.3 $Y2=1.49
r174 45 47 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=2.295 $Y=1.49
+ $X2=0.94 $Y2=1.49
r175 41 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.655
+ $X2=2.46 $Y2=1.49
r176 41 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.46 $Y=1.655
+ $X2=2.46 $Y2=2.465
r177 37 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.655
+ $X2=2.03 $Y2=1.49
r178 37 39 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.03 $Y=1.655
+ $X2=2.03 $Y2=2.465
r179 33 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.325
+ $X2=1.795 $Y2=1.49
r180 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.795 $Y=1.325
+ $X2=1.795 $Y2=0.665
r181 29 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=1.655
+ $X2=1.6 $Y2=1.49
r182 29 31 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.6 $Y=1.655 $X2=1.6
+ $Y2=2.465
r183 25 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.49
r184 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=0.665
r185 21 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.655
+ $X2=1.17 $Y2=1.49
r186 21 23 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.17 $Y=1.655
+ $X2=1.17 $Y2=2.465
r187 17 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.325
+ $X2=0.935 $Y2=1.49
r188 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.935 $Y=1.325
+ $X2=0.935 $Y2=0.665
r189 13 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.505 $Y2=1.49
r190 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.505 $Y2=0.665
r191 4 76 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=5.34
+ $Y=1.835 $X2=5.48 $Y2=2.095
r192 3 74 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=3.47
+ $Y=1.835 $X2=3.61 $Y2=2.095
r193 2 56 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.04 $Y2=0.4
r194 1 54 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.04
+ $Y=0.235 $X2=3.18 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%B1 3 6 10 13 15 16 17 21 23 26 28 31
c81 26 0 8.07691e-20 $X=2.945 $Y=1.36
r82 26 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=1.36
+ $X2=2.945 $Y2=1.525
r83 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=1.36
+ $X2=2.945 $Y2=1.195
r84 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.945
+ $Y=1.36 $X2=2.945 $Y2=1.36
r85 23 27 5.3375 $w=4e-07 $l=1.75e-07 $layer=LI1_cond $X=3.12 $Y=1.3 $X2=2.945
+ $Y2=1.3
r86 21 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.275 $Y=1.35
+ $X2=4.275 $Y2=1.515
r87 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.275 $Y=1.35
+ $X2=4.275 $Y2=1.185
r88 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.275
+ $Y=1.35 $X2=4.275 $Y2=1.35
r89 17 20 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.275 $Y=1.16
+ $X2=4.275 $Y2=1.35
r90 16 23 9.15454 $w=4e-07 $l=2.24332e-07 $layer=LI1_cond $X=3.285 $Y=1.16
+ $X2=3.12 $Y2=1.3
r91 15 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.11 $Y=1.16
+ $X2=4.275 $Y2=1.16
r92 15 16 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.11 $Y=1.16
+ $X2=3.285 $Y2=1.16
r93 13 32 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.255 $Y=2.465
+ $X2=4.255 $Y2=1.515
r94 10 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.255 $Y=0.655
+ $X2=4.255 $Y2=1.185
r95 6 29 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.965 $Y=2.465 $X2=2.965
+ $Y2=1.525
r96 3 28 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.965 $Y=0.655
+ $X2=2.965 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%B2 3 7 11 15 17 23 24
c45 23 0 8.07691e-20 $X=3.735 $Y=1.51
r46 22 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.735 $Y=1.51
+ $X2=3.825 $Y2=1.51
r47 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.735
+ $Y=1.51 $X2=3.735 $Y2=1.51
r48 19 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.395 $Y=1.51
+ $X2=3.735 $Y2=1.51
r49 17 23 4.01413 $w=4.43e-07 $l=1.55e-07 $layer=LI1_cond $X=3.677 $Y=1.665
+ $X2=3.677 $Y2=1.51
r50 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.675
+ $X2=3.825 $Y2=1.51
r51 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.825 $Y=1.675
+ $X2=3.825 $Y2=2.465
r52 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.345
+ $X2=3.825 $Y2=1.51
r53 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.825 $Y=1.345
+ $X2=3.825 $Y2=0.655
r54 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.675
+ $X2=3.395 $Y2=1.51
r55 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.395 $Y=1.675
+ $X2=3.395 $Y2=2.465
r56 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.345
+ $X2=3.395 $Y2=1.51
r57 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.395 $Y=1.345
+ $X2=3.395 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%A1 3 6 10 13 15 17 21 23 25 32 35 37
c71 17 0 1.11629e-19 $X=4.815 $Y=1.16
r72 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.215 $Y=1.35
+ $X2=6.215 $Y2=1.515
r73 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.215 $Y=1.35
+ $X2=6.215 $Y2=1.185
r74 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.35 $X2=6.215 $Y2=1.35
r75 25 36 5.26547 $w=6.14e-07 $l=2.65e-07 $layer=LI1_cond $X=6.48 $Y=1.422
+ $X2=6.215 $Y2=1.422
r76 23 36 4.27199 $w=6.14e-07 $l=2.15e-07 $layer=LI1_cond $X=6 $Y=1.422
+ $X2=6.215 $Y2=1.422
r77 21 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.35
+ $X2=4.815 $Y2=1.515
r78 21 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.35
+ $X2=4.815 $Y2=1.185
r79 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.815
+ $Y=1.35 $X2=4.815 $Y2=1.35
r80 17 20 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.815 $Y=1.16
+ $X2=4.815 $Y2=1.35
r81 16 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.98 $Y=1.16
+ $X2=4.815 $Y2=1.16
r82 15 23 10.1543 $w=6.14e-07 $l=3.28548e-07 $layer=LI1_cond $X=5.85 $Y=1.16
+ $X2=6 $Y2=1.422
r83 15 16 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=5.85 $Y=1.16
+ $X2=4.98 $Y2=1.16
r84 13 38 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.125 $Y=2.465
+ $X2=6.125 $Y2=1.515
r85 10 37 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.125 $Y=0.655
+ $X2=6.125 $Y2=1.185
r86 6 33 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.835 $Y=2.465
+ $X2=4.835 $Y2=1.515
r87 3 32 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.765 $Y=0.655
+ $X2=4.765 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%A2 3 7 11 15 17 24
c47 24 0 1.11629e-19 $X=5.695 $Y=1.51
r48 22 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.355 $Y=1.51
+ $X2=5.695 $Y2=1.51
r49 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.355
+ $Y=1.51 $X2=5.355 $Y2=1.51
r50 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.265 $Y=1.51
+ $X2=5.355 $Y2=1.51
r51 17 23 5.67621 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=1.592
+ $X2=5.355 $Y2=1.592
r52 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.675
+ $X2=5.695 $Y2=1.51
r53 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.695 $Y=1.675
+ $X2=5.695 $Y2=2.465
r54 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.345
+ $X2=5.695 $Y2=1.51
r55 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.695 $Y=1.345
+ $X2=5.695 $Y2=0.655
r56 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.675
+ $X2=5.265 $Y2=1.51
r57 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.265 $Y=1.675
+ $X2=5.265 $Y2=2.465
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.345
+ $X2=5.265 $Y2=1.51
r59 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.265 $Y=1.345
+ $X2=5.265 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%VPWR 1 2 3 4 5 18 22 26 32 36 38 40 44 45 46
+ 52 57 65 74 77 80 84
r88 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r91 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 72 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r93 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r94 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r95 69 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 68 71 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r97 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r98 66 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.71 $Y=3.33
+ $X2=4.545 $Y2=3.33
r99 66 68 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.71 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 65 83 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.447 $Y2=3.33
r101 65 71 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6 $Y2=3.33
r102 64 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r104 61 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r106 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r107 58 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=2.71 $Y2=3.33
r108 58 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 57 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=3.33
+ $X2=4.545 $Y2=3.33
r110 57 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.38 $Y=3.33 $X2=4.08
+ $Y2=3.33
r111 56 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 56 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r113 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r114 53 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=3.33
+ $X2=1.815 $Y2=3.33
r115 53 55 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.98 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 52 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.71 $Y2=3.33
r117 52 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 50 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r119 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 46 64 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r121 46 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r122 44 49 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.79 $Y=3.33 $X2=0.72
+ $Y2=3.33
r123 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=3.33
+ $X2=0.955 $Y2=3.33
r124 40 43 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=6.34 $Y=2.025
+ $X2=6.34 $Y2=2.95
r125 38 83 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.34 $Y=3.245
+ $X2=6.447 $Y2=3.33
r126 38 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.34 $Y=3.245
+ $X2=6.34 $Y2=2.95
r127 34 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=3.245
+ $X2=4.545 $Y2=3.33
r128 34 36 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=4.545 $Y=3.245
+ $X2=4.545 $Y2=2.38
r129 30 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=3.33
r130 30 32 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=2.405
r131 26 29 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.815 $Y=2.19
+ $X2=1.815 $Y2=2.95
r132 24 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=3.245
+ $X2=1.815 $Y2=3.33
r133 24 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.815 $Y=3.245
+ $X2=1.815 $Y2=2.95
r134 23 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=3.33
+ $X2=0.955 $Y2=3.33
r135 22 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.815 $Y2=3.33
r136 22 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.12 $Y2=3.33
r137 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.955 $Y=2.18
+ $X2=0.955 $Y2=2.95
r138 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=3.245
+ $X2=0.955 $Y2=3.33
r139 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.955 $Y=3.245
+ $X2=0.955 $Y2=2.95
r140 5 43 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.2
+ $Y=1.835 $X2=6.34 $Y2=2.95
r141 5 40 400 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=6.2
+ $Y=1.835 $X2=6.34 $Y2=2.025
r142 4 36 300 $w=1.7e-07 $l=6.43584e-07 $layer=licon1_PDIFF $count=2 $X=4.33
+ $Y=1.835 $X2=4.545 $Y2=2.38
r143 3 32 300 $w=1.7e-07 $l=6.51652e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.835 $X2=2.71 $Y2=2.405
r144 2 29 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.675
+ $Y=1.835 $X2=1.815 $Y2=2.95
r145 2 26 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.675
+ $Y=1.835 $X2=1.815 $Y2=2.19
r146 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.83
+ $Y=1.835 $X2=0.955 $Y2=2.95
r147 1 18 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.83
+ $Y=1.835 $X2=0.955 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%X 1 2 3 4 13 14 17 19 20 23 27 31 35 40 41 42
+ 48
r54 46 55 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.295 $Y=1.14
+ $X2=0.72 $Y2=1.14
r55 46 48 1.92074 $w=4.18e-07 $l=7e-08 $layer=LI1_cond $X=0.295 $Y=1.225
+ $X2=0.295 $Y2=1.295
r56 41 46 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.24 $Y=1.14
+ $X2=0.295 $Y2=1.14
r57 41 42 9.9604 $w=4.18e-07 $l=3.63e-07 $layer=LI1_cond $X=0.295 $Y=1.302
+ $X2=0.295 $Y2=1.665
r58 41 48 0.192074 $w=4.18e-07 $l=7e-09 $layer=LI1_cond $X=0.295 $Y=1.302
+ $X2=0.295 $Y2=1.295
r59 39 42 2.46952 $w=4.18e-07 $l=9e-08 $layer=LI1_cond $X=0.295 $Y=1.755
+ $X2=0.295 $Y2=1.665
r60 35 37 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.245 $Y=1.98
+ $X2=2.245 $Y2=2.91
r61 33 35 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=2.245 $Y=1.925
+ $X2=2.245 $Y2=1.98
r62 29 31 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.6 $Y=1.055
+ $X2=1.6 $Y2=0.42
r63 28 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.48 $Y=1.84
+ $X2=1.385 $Y2=1.84
r64 27 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.15 $Y=1.84
+ $X2=2.245 $Y2=1.925
r65 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.15 $Y=1.84
+ $X2=1.48 $Y2=1.84
r66 23 25 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.385 $Y=1.98
+ $X2=1.385 $Y2=2.91
r67 21 40 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=1.925
+ $X2=1.385 $Y2=1.84
r68 21 23 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.385 $Y=1.925
+ $X2=1.385 $Y2=1.98
r69 20 55 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.815 $Y=1.14
+ $X2=0.72 $Y2=1.14
r70 19 29 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.485 $Y=1.14
+ $X2=1.6 $Y2=1.055
r71 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.485 $Y=1.14
+ $X2=0.815 $Y2=1.14
r72 15 55 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.055
+ $X2=0.72 $Y2=1.14
r73 15 17 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.72 $Y=1.055
+ $X2=0.72 $Y2=0.42
r74 14 39 8.54503 $w=1.7e-07 $l=2.48898e-07 $layer=LI1_cond $X=0.505 $Y=1.84
+ $X2=0.295 $Y2=1.755
r75 13 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.29 $Y=1.84
+ $X2=1.385 $Y2=1.84
r76 13 14 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.29 $Y=1.84
+ $X2=0.505 $Y2=1.84
r77 4 37 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.105
+ $Y=1.835 $X2=2.245 $Y2=2.91
r78 4 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.105
+ $Y=1.835 $X2=2.245 $Y2=1.98
r79 3 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.835 $X2=1.385 $Y2=2.91
r80 3 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.835 $X2=1.385 $Y2=1.98
r81 2 31 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.44
+ $Y=0.245 $X2=1.58 $Y2=0.42
r82 1 17 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.245 $X2=0.72 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%A_608_367# 1 2 9 11 12 15
r16 13 15 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=4.075 $Y=2.905
+ $X2=4.075 $Y2=2.435
r17 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.945 $Y=2.99
+ $X2=4.075 $Y2=2.905
r18 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.945 $Y=2.99
+ $X2=3.275 $Y2=2.99
r19 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.16 $Y=2.905
+ $X2=3.275 $Y2=2.99
r20 7 9 23.5499 $w=2.28e-07 $l=4.7e-07 $layer=LI1_cond $X=3.16 $Y=2.905 $X2=3.16
+ $Y2=2.435
r21 2 15 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=3.9
+ $Y=1.835 $X2=4.04 $Y2=2.435
r22 1 9 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=3.04
+ $Y=1.835 $X2=3.18 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%A_982_367# 1 2 9 11 12 13 15
r17 13 18 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=2.905
+ $X2=5.91 $Y2=2.99
r18 13 15 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=5.91 $Y=2.905 $X2=5.91
+ $Y2=2.105
r19 11 18 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.815 $Y=2.99
+ $X2=5.91 $Y2=2.99
r20 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.815 $Y=2.99
+ $X2=5.145 $Y2=2.99
r21 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.015 $Y=2.905
+ $X2=5.145 $Y2=2.99
r22 7 9 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=5.015 $Y=2.905
+ $X2=5.015 $Y2=2.435
r23 2 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.835 $X2=5.91 $Y2=2.91
r24 2 15 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.835 $X2=5.91 $Y2=2.105
r25 1 9 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=4.91
+ $Y=1.835 $X2=5.05 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 42 44 53 65 66 72 75
r99 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r100 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r101 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r102 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r103 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r104 63 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r105 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r106 60 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.01
+ $Y2=0
r107 60 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.52
+ $Y2=0
r108 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r109 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r110 55 58 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r111 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 53 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=0 $X2=5.01
+ $Y2=0
r113 53 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.845 $Y=0
+ $X2=4.56 $Y2=0
r114 52 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r115 52 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r116 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r117 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.15
+ $Y2=0
r118 49 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=0
+ $X2=1.68 $Y2=0
r119 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r120 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r121 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r122 45 69 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0
+ $X2=0.227 $Y2=0
r123 45 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0
+ $X2=0.72 $Y2=0
r124 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.15
+ $Y2=0
r125 44 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0
+ $X2=0.72 $Y2=0
r126 42 59 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.56
+ $Y2=0
r127 42 56 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.16
+ $Y2=0
r128 40 62 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.745 $Y=0
+ $X2=5.52 $Y2=0
r129 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=0 $X2=5.91
+ $Y2=0
r130 39 65 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=6.48 $Y2=0
r131 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0 $X2=5.91
+ $Y2=0
r132 37 51 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=0
+ $X2=1.68 $Y2=0
r133 37 38 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.005
+ $Y2=0
r134 36 55 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.16
+ $Y2=0
r135 36 38 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.005
+ $Y2=0
r136 32 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=0.085
+ $X2=5.91 $Y2=0
r137 32 34 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.91 $Y=0.085
+ $X2=5.91 $Y2=0.44
r138 28 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.085
+ $X2=5.01 $Y2=0
r139 28 30 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.01 $Y=0.085
+ $X2=5.01 $Y2=0.44
r140 24 38 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0
r141 24 26 14.6456 $w=2.38e-07 $l=3.05e-07 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0.39
r142 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r143 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.37
r144 16 69 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r145 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.29 $Y2=0.39
r146 5 34 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.77
+ $Y=0.235 $X2=5.91 $Y2=0.44
r147 4 30 182 $w=1.7e-07 $l=2.77263e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.235 $X2=5.01 $Y2=0.44
r148 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.245 $X2=2.01 $Y2=0.39
r149 2 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.245 $X2=1.15 $Y2=0.37
r150 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.245 $X2=0.29 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_4%A_525_47# 1 2 3 4 5 16 22 24 28 30 32 34 39
+ 41 43
r59 37 39 5.29958 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.75 $Y=0.85
+ $X2=2.865 $Y2=0.85
r60 32 45 3.13575 $w=2.6e-07 $l=1.44914e-07 $layer=LI1_cond $X=6.375 $Y=0.735
+ $X2=6.365 $Y2=0.875
r61 32 34 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=6.375 $Y=0.735
+ $X2=6.375 $Y2=0.42
r62 31 43 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.575 $Y=0.82
+ $X2=5.46 $Y2=0.82
r63 30 45 4.07647 $w=1.7e-07 $l=1.65227e-07 $layer=LI1_cond $X=6.225 $Y=0.82
+ $X2=6.365 $Y2=0.875
r64 30 31 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.225 $Y=0.82
+ $X2=5.575 $Y2=0.82
r65 26 43 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.46 $Y=0.735
+ $X2=5.46 $Y2=0.82
r66 26 28 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.46 $Y=0.735
+ $X2=5.46 $Y2=0.42
r67 25 41 7.08839 $w=1.95e-07 $l=1.57003e-07 $layer=LI1_cond $X=4.675 $Y=0.82
+ $X2=4.53 $Y2=0.795
r68 24 43 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.345 $Y=0.82
+ $X2=5.46 $Y2=0.82
r69 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.345 $Y=0.82
+ $X2=4.675 $Y2=0.82
r70 20 41 0.0392004 $w=2.9e-07 $l=1.1e-07 $layer=LI1_cond $X=4.53 $Y=0.685
+ $X2=4.53 $Y2=0.795
r71 20 22 10.5309 $w=2.88e-07 $l=2.65e-07 $layer=LI1_cond $X=4.53 $Y=0.685
+ $X2=4.53 $Y2=0.42
r72 19 39 39.0259 $w=2.18e-07 $l=7.45e-07 $layer=LI1_cond $X=3.61 $Y=0.795
+ $X2=2.865 $Y2=0.795
r73 16 41 7.08839 $w=1.95e-07 $l=1.45e-07 $layer=LI1_cond $X=4.385 $Y=0.795
+ $X2=4.53 $Y2=0.795
r74 16 19 40.5974 $w=2.18e-07 $l=7.75e-07 $layer=LI1_cond $X=4.385 $Y=0.795
+ $X2=3.61 $Y2=0.795
r75 5 45 182 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_NDIFF $count=1 $X=6.2
+ $Y=0.235 $X2=6.34 $Y2=0.85
r76 5 34 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.2
+ $Y=0.235 $X2=6.34 $Y2=0.42
r77 4 43 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.235 $X2=5.48 $Y2=0.82
r78 4 28 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.235 $X2=5.48 $Y2=0.42
r79 3 41 182 $w=1.7e-07 $l=6.8624e-07 $layer=licon1_NDIFF $count=1 $X=4.33
+ $Y=0.235 $X2=4.55 $Y2=0.82
r80 3 22 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=4.33
+ $Y=0.235 $X2=4.55 $Y2=0.42
r81 2 19 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=3.47
+ $Y=0.235 $X2=3.61 $Y2=0.79
r82 1 37 182 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.75 $Y2=0.85
.ends

