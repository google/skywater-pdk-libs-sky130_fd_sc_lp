* File: sky130_fd_sc_lp__and2_m.pxi.spice
* Created: Fri Aug 28 10:04:51 2020
* 
x_PM_SKY130_FD_SC_LP__AND2_M%A N_A_M1004_g N_A_c_37_n N_A_M1003_g A A
+ PM_SKY130_FD_SC_LP__AND2_M%A
x_PM_SKY130_FD_SC_LP__AND2_M%B N_B_M1001_g N_B_M1005_g N_B_c_62_n B B N_B_c_63_n
+ N_B_c_64_n PM_SKY130_FD_SC_LP__AND2_M%B
x_PM_SKY130_FD_SC_LP__AND2_M%A_34_141# N_A_34_141#_M1004_s N_A_34_141#_M1003_d
+ N_A_34_141#_c_92_n N_A_34_141#_M1002_g N_A_34_141#_M1000_g N_A_34_141#_c_90_n
+ N_A_34_141#_c_91_n N_A_34_141#_c_95_n PM_SKY130_FD_SC_LP__AND2_M%A_34_141#
x_PM_SKY130_FD_SC_LP__AND2_M%VPWR N_VPWR_M1003_s N_VPWR_M1005_d N_VPWR_c_137_n
+ N_VPWR_c_138_n N_VPWR_c_139_n N_VPWR_c_140_n VPWR N_VPWR_c_141_n
+ N_VPWR_c_136_n N_VPWR_c_143_n PM_SKY130_FD_SC_LP__AND2_M%VPWR
x_PM_SKY130_FD_SC_LP__AND2_M%X N_X_M1002_d N_X_M1000_d X X X X X X X
+ PM_SKY130_FD_SC_LP__AND2_M%X
x_PM_SKY130_FD_SC_LP__AND2_M%VGND N_VGND_M1001_d N_VGND_c_176_n N_VGND_c_177_n
+ N_VGND_c_178_n N_VGND_c_179_n VGND N_VGND_c_180_n N_VGND_c_181_n
+ PM_SKY130_FD_SC_LP__AND2_M%VGND
cc_1 VNB N_A_M1004_g 0.0242225f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.915
cc_2 VNB N_A_c_37_n 0.0424013f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.775
cc_3 VNB A 0.0194077f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B_M1001_g 0.0110295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_B_M1005_g 0.0136887f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.195
cc_6 VNB N_B_c_62_n 0.0175094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_63_n 0.0419192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_64_n 0.0290606f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.46
cc_9 VNB N_A_34_141#_M1002_g 0.0420768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_34_141#_c_90_n 0.0103949f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.46
cc_11 VNB N_A_34_141#_c_91_n 0.00328683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_136_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB X 0.0402804f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.195
cc_14 VNB N_VGND_c_176_n 0.00981171f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.195
cc_15 VNB N_VGND_c_177_n 0.0183219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_178_n 0.0329304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_179_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_180_n 0.0176897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_181_n 0.14844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VPB N_A_c_37_n 0.0241949f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.775
cc_21 VPB N_A_M1003_g 0.0274889f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.195
cc_22 VPB A 0.00423747f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_23 VPB N_B_M1005_g 0.0248645f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.195
cc_24 VPB N_A_34_141#_c_92_n 0.0422422f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.195
cc_25 VPB N_A_34_141#_M1002_g 0.0398132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_A_34_141#_c_91_n 0.0042121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_A_34_141#_c_95_n 0.044626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_137_n 0.0116371f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.195
cc_29 VPB N_VPWR_c_138_n 0.0401997f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_VPWR_c_139_n 0.0208198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_140_n 0.0188628f $X=-0.19 $Y=1.655 $X2=0.35 $Y2=1.46
cc_32 VPB N_VPWR_c_141_n 0.019599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_136_n 0.0662039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_143_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB X 0.0407654f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.195
cc_36 N_A_c_37_n N_B_M1001_g 0.0250751f $X=0.585 $Y=1.775 $X2=0 $Y2=0
cc_37 N_A_c_37_n N_B_M1005_g 0.0330239f $X=0.585 $Y=1.775 $X2=0 $Y2=0
cc_38 A N_B_M1005_g 2.33145e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_39 N_A_M1004_g N_B_c_63_n 0.0250751f $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_40 N_A_M1004_g N_B_c_64_n 0.00797344f $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_41 N_A_M1004_g N_A_34_141#_c_90_n 0.0136476f $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_42 N_A_c_37_n N_A_34_141#_c_90_n 0.0012985f $X=0.585 $Y=1.775 $X2=0 $Y2=0
cc_43 A N_A_34_141#_c_90_n 0.0200582f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_44 N_A_M1004_g N_A_34_141#_c_91_n 0.00639451f $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_45 N_A_c_37_n N_A_34_141#_c_91_n 0.00643393f $X=0.585 $Y=1.775 $X2=0 $Y2=0
cc_46 N_A_M1003_g N_A_34_141#_c_91_n 0.0257486f $X=0.585 $Y=2.195 $X2=0 $Y2=0
cc_47 A N_A_34_141#_c_91_n 0.0402781f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_48 N_A_M1003_g N_A_34_141#_c_95_n 0.00249837f $X=0.585 $Y=2.195 $X2=0 $Y2=0
cc_49 N_A_c_37_n N_VPWR_c_138_n 0.00448953f $X=0.585 $Y=1.775 $X2=0 $Y2=0
cc_50 N_A_M1003_g N_VPWR_c_138_n 0.00923921f $X=0.585 $Y=2.195 $X2=0 $Y2=0
cc_51 A N_VPWR_c_138_n 0.0104075f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_VPWR_c_136_n 0.00276198f $X=0.585 $Y=2.195 $X2=0 $Y2=0
cc_53 N_A_M1004_g N_VGND_c_178_n 4.61482e-19 $X=0.51 $Y=0.915 $X2=0 $Y2=0
cc_54 N_B_M1001_g N_A_34_141#_M1002_g 0.011069f $X=0.87 $Y=0.915 $X2=0 $Y2=0
cc_55 N_B_c_62_n N_A_34_141#_M1002_g 0.03918f $X=1.015 $Y=1.31 $X2=0 $Y2=0
cc_56 N_B_c_63_n N_A_34_141#_M1002_g 0.0010113f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_57 N_B_M1001_g N_A_34_141#_c_90_n 0.00707946f $X=0.87 $Y=0.915 $X2=0 $Y2=0
cc_58 N_B_c_64_n N_A_34_141#_c_90_n 0.0527213f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_59 N_B_M1001_g N_A_34_141#_c_91_n 0.00586534f $X=0.87 $Y=0.915 $X2=0 $Y2=0
cc_60 N_B_M1005_g N_A_34_141#_c_91_n 0.0261187f $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_61 N_B_c_62_n N_A_34_141#_c_91_n 0.009301f $X=1.015 $Y=1.31 $X2=0 $Y2=0
cc_62 N_B_M1005_g N_A_34_141#_c_95_n 0.00965003f $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_63 N_B_M1005_g N_VPWR_c_140_n 9.84115e-19 $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_64 N_B_M1001_g N_VGND_c_176_n 0.0016789f $X=0.87 $Y=0.915 $X2=0 $Y2=0
cc_65 N_B_M1001_g N_VGND_c_177_n 0.0036052f $X=0.87 $Y=0.915 $X2=0 $Y2=0
cc_66 N_B_c_63_n N_VGND_c_177_n 0.00773842f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_67 N_B_c_64_n N_VGND_c_177_n 0.0287387f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_68 N_B_c_63_n N_VGND_c_178_n 0.00870324f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_69 N_B_c_64_n N_VGND_c_178_n 0.0562652f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_70 N_B_c_63_n N_VGND_c_181_n 0.0111008f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_71 N_B_c_64_n N_VGND_c_181_n 0.0337313f $X=0.96 $Y=0.43 $X2=0 $Y2=0
cc_72 N_A_34_141#_c_91_n N_VPWR_c_138_n 0.0563274f $X=0.8 $Y=2.26 $X2=0 $Y2=0
cc_73 N_A_34_141#_c_95_n N_VPWR_c_138_n 0.00861359f $X=0.78 $Y=2.85 $X2=0 $Y2=0
cc_74 N_A_34_141#_c_92_n N_VPWR_c_139_n 0.00445258f $X=1.37 $Y=2.85 $X2=0 $Y2=0
cc_75 N_A_34_141#_c_91_n N_VPWR_c_139_n 0.0167839f $X=0.8 $Y=2.26 $X2=0 $Y2=0
cc_76 N_A_34_141#_c_95_n N_VPWR_c_139_n 0.0059602f $X=0.78 $Y=2.85 $X2=0 $Y2=0
cc_77 N_A_34_141#_c_92_n N_VPWR_c_140_n 0.018252f $X=1.37 $Y=2.85 $X2=0 $Y2=0
cc_78 N_A_34_141#_M1002_g N_VPWR_c_140_n 0.00678324f $X=1.445 $Y=0.915 $X2=0
+ $Y2=0
cc_79 N_A_34_141#_c_91_n N_VPWR_c_140_n 0.0568527f $X=0.8 $Y=2.26 $X2=0 $Y2=0
cc_80 N_A_34_141#_c_95_n N_VPWR_c_140_n 0.00508672f $X=0.78 $Y=2.85 $X2=0 $Y2=0
cc_81 N_A_34_141#_c_92_n N_VPWR_c_141_n 0.00550617f $X=1.37 $Y=2.85 $X2=0 $Y2=0
cc_82 N_A_34_141#_c_92_n N_VPWR_c_136_n 0.0106337f $X=1.37 $Y=2.85 $X2=0 $Y2=0
cc_83 N_A_34_141#_c_91_n N_VPWR_c_136_n 0.0108843f $X=0.8 $Y=2.26 $X2=0 $Y2=0
cc_84 N_A_34_141#_c_95_n N_VPWR_c_136_n 0.00806414f $X=0.78 $Y=2.85 $X2=0 $Y2=0
cc_85 N_A_34_141#_M1002_g X 0.0408638f $X=1.445 $Y=0.915 $X2=0 $Y2=0
cc_86 N_A_34_141#_c_91_n X 0.0244925f $X=0.8 $Y=2.26 $X2=0 $Y2=0
cc_87 N_A_34_141#_c_90_n A_117_141# 0.00107385f $X=0.615 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_34_141#_M1002_g N_VGND_c_176_n 0.00514587f $X=1.445 $Y=0.915 $X2=0
+ $Y2=0
cc_89 N_A_34_141#_c_90_n N_VGND_c_176_n 0.016313f $X=0.615 $Y=0.925 $X2=0 $Y2=0
cc_90 N_A_34_141#_c_91_n N_VGND_c_176_n 0.00877806f $X=0.8 $Y=2.26 $X2=0 $Y2=0
cc_91 N_A_34_141#_M1002_g N_VGND_c_177_n 0.00536689f $X=1.445 $Y=0.915 $X2=0
+ $Y2=0
cc_92 N_A_34_141#_M1002_g N_VGND_c_180_n 0.0031218f $X=1.445 $Y=0.915 $X2=0
+ $Y2=0
cc_93 N_A_34_141#_M1002_g N_VGND_c_181_n 0.00376215f $X=1.445 $Y=0.915 $X2=0
+ $Y2=0
cc_94 N_A_34_141#_c_90_n N_VGND_c_181_n 0.0015772f $X=0.615 $Y=0.925 $X2=0 $Y2=0
cc_95 N_VPWR_c_140_n X 0.0271668f $X=1.23 $Y=2.26 $X2=0 $Y2=0
cc_96 N_VPWR_c_141_n X 0.00563668f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_97 N_VPWR_c_136_n X 0.00642236f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_98 X N_VGND_c_177_n 0.0326503f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_99 X N_VGND_c_180_n 0.00563668f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_100 X N_VGND_c_181_n 0.00642236f $X=1.595 $Y=0.47 $X2=0 $Y2=0
