# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.840000 0.865000 1.790000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.160000 0.345000 6.630000 1.170000 ;
        RECT 6.260000 1.850000 6.630000 3.075000 ;
        RECT 6.450000 1.170000 6.630000 1.850000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.425000 0.345000 5.605000 1.345000 ;
        RECT 5.425000 1.345000 5.740000 2.130000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.035000 0.840000 1.375000 1.790000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.165000  0.390000 0.455000 1.960000 ;
      RECT 0.165000  1.960000 1.185000 2.130000 ;
      RECT 0.165000  2.130000 0.455000 2.980000 ;
      RECT 0.655000  2.300000 0.845000 3.245000 ;
      RECT 0.715000  0.085000 1.045000 0.670000 ;
      RECT 1.015000  2.130000 1.185000 2.905000 ;
      RECT 1.015000  2.905000 2.420000 3.075000 ;
      RECT 1.220000  0.330000 1.725000 0.670000 ;
      RECT 1.355000  2.405000 1.725000 2.735000 ;
      RECT 1.545000  0.670000 1.725000 2.405000 ;
      RECT 1.895000  0.255000 2.360000 0.535000 ;
      RECT 1.895000  0.535000 2.075000 1.195000 ;
      RECT 1.895000  1.195000 3.475000 1.365000 ;
      RECT 1.895000  1.365000 2.080000 2.735000 ;
      RECT 2.245000  0.705000 3.825000 0.875000 ;
      RECT 2.245000  0.875000 2.575000 1.025000 ;
      RECT 2.250000  1.535000 2.810000 2.175000 ;
      RECT 2.250000  2.175000 2.420000 2.905000 ;
      RECT 2.530000  0.085000 2.810000 0.535000 ;
      RECT 2.590000  2.345000 2.820000 3.245000 ;
      RECT 2.990000  1.365000 3.160000 2.905000 ;
      RECT 2.990000  2.905000 4.050000 3.075000 ;
      RECT 3.145000  1.045000 3.475000 1.195000 ;
      RECT 3.340000  1.605000 4.915000 1.775000 ;
      RECT 3.340000  1.775000 3.510000 2.405000 ;
      RECT 3.340000  2.405000 3.700000 2.735000 ;
      RECT 3.380000  0.315000 4.175000 0.535000 ;
      RECT 3.655000  0.875000 3.825000 1.175000 ;
      RECT 3.655000  1.175000 4.015000 1.435000 ;
      RECT 3.690000  1.945000 4.050000 2.205000 ;
      RECT 3.880000  2.205000 4.050000 2.905000 ;
      RECT 4.005000  0.535000 4.175000 0.725000 ;
      RECT 4.005000  0.725000 4.705000 0.895000 ;
      RECT 4.230000  1.945000 5.255000 2.205000 ;
      RECT 4.345000  0.085000 4.595000 0.555000 ;
      RECT 4.365000  2.400000 4.915000 2.640000 ;
      RECT 4.365000  2.640000 5.085000 3.245000 ;
      RECT 4.535000  0.895000 4.705000 1.335000 ;
      RECT 4.535000  1.335000 4.915000 1.605000 ;
      RECT 4.875000  0.345000 5.255000 1.165000 ;
      RECT 5.085000  1.165000 5.255000 1.945000 ;
      RECT 5.085000  2.205000 5.255000 2.300000 ;
      RECT 5.085000  2.300000 6.090000 2.470000 ;
      RECT 5.255000  2.470000 5.555000 3.075000 ;
      RECT 5.725000  2.640000 6.055000 3.245000 ;
      RECT 5.775000  0.085000 5.990000 1.170000 ;
      RECT 5.920000  1.340000 6.280000 1.670000 ;
      RECT 5.920000  1.670000 6.090000 2.300000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrtp_1
