* File: sky130_fd_sc_lp__o41ai_2.spice
* Created: Wed Sep  2 10:28:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41ai_2.pex.spice"
.subckt sky130_fd_sc_lp__o41ai_2  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_155_47#_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1008 N_Y_M1007_d N_B1_M1008_g N_A_155_47#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_A4_M1015_g N_A_155_47#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1869 AS=0.1176 PD=1.285 PS=1.12 NRD=10.704 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1015_d N_A4_M1016_g N_A_155_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1869 AS=0.1176 PD=1.285 PS=1.12 NRD=12.852 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A3_M1001_g N_A_155_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1428 AS=0.1176 PD=1.18 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1001_d N_A3_M1014_g N_A_155_47#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1428 AS=0.1176 PD=1.18 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_155_47#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1003_d N_A2_M1012_g N_A_155_47#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_A_155_47#_M1012_s N_A1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_A_155_47#_M1017_d N_A1_M1017_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75004.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_B1_M1018_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_A_313_365#_M1002_d N_A4_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1011 N_A_313_365#_M1011_d N_A4_M1011_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.32445 AS=0.1764 PD=1.775 PS=1.54 NRD=19.5424 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1013 N_A_313_365#_M1011_d N_A3_M1013_g N_A_615_365#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.32445 AS=0.1764 PD=1.775 PS=1.54 NRD=17.1981 NRS=0 M=1 R=8.4
+ SA=75001.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_A_313_365#_M1019_d N_A3_M1019_g N_A_615_365#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_808_367#_M1000_d N_A2_M1000_g N_A_615_365#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_A_808_367#_M1006_d N_A2_M1006_g N_A_615_365#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_A_808_367#_M1006_d N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_808_367#_M1010_d N_A1_M1010_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3719 P=16.99
*
.include "sky130_fd_sc_lp__o41ai_2.pxi.spice"
*
.ends
*
*
