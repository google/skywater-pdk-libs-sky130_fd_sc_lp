* File: sky130_fd_sc_lp__and4_1.pex.spice
* Created: Wed Sep  2 09:32:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4_1%A 2 5 9 11 12 13 14 19
c28 12 0 1.05412e-19 $X=0.24 $Y=0.925
r29 19 21 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.005
+ $X2=0.43 $Y2=0.84
r30 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.41
+ $Y=1.005 $X2=0.41 $Y2=1.005
r31 13 14 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r32 13 20 8.15143 $w=4.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.005
r33 12 20 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=0.29 $Y=0.925 $X2=0.29
+ $Y2=1.005
r34 9 11 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.54 $Y=2.045
+ $X2=0.54 $Y2=1.51
r35 5 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.54 $Y=0.445
+ $X2=0.54 $Y2=0.84
r36 2 11 49.8761 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=0.43 $Y=1.325
+ $X2=0.43 $Y2=1.51
r37 1 19 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=0.43 $Y=1.025 $X2=0.43
+ $Y2=1.005
r38 1 2 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=0.43 $Y=1.025 $X2=0.43
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_1%B 3 7 11 12 13 14 18
c34 7 0 1.05412e-19 $X=1.08 $Y=2.045
r35 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.11
+ $Y=0.97 $X2=1.11 $Y2=0.97
r36 14 19 11.7045 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=1.185 $Y=1.295
+ $X2=1.185 $Y2=0.97
r37 13 19 1.62062 $w=3.18e-07 $l=4.5e-08 $layer=LI1_cond $X=1.185 $Y=0.925
+ $X2=1.185 $Y2=0.97
r38 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.11 $Y=1.31
+ $X2=1.11 $Y2=0.97
r39 11 12 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.31
+ $X2=1.11 $Y2=1.475
r40 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=0.805
+ $X2=1.11 $Y2=0.97
r41 7 12 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.08 $Y=2.045
+ $X2=1.08 $Y2=1.475
r42 3 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.02 $Y=0.445
+ $X2=1.02 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_1%C 3 7 11 12 13 14 18
c30 12 0 1.60954e-19 $X=1.65 $Y=1.475
r31 13 14 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.67 $Y=0.925
+ $X2=1.67 $Y2=1.295
r32 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.65
+ $Y=0.97 $X2=1.65 $Y2=0.97
r33 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.65 $Y=1.31
+ $X2=1.65 $Y2=0.97
r34 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.31
+ $X2=1.65 $Y2=1.475
r35 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=0.805
+ $X2=1.65 $Y2=0.97
r36 7 12 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.67 $Y=2.045
+ $X2=1.67 $Y2=1.475
r37 3 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.56 $Y=0.445
+ $X2=1.56 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_1%D 3 7 9 12 13
c34 13 0 1.60954e-19 $X=2.19 $Y=1.51
r35 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.51
+ $X2=2.19 $Y2=1.675
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.51
+ $X2=2.19 $Y2=1.345
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.51 $X2=2.19 $Y2=1.51
r38 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.19 $Y=1.665
+ $X2=2.19 $Y2=1.51
r39 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.1 $Y=2.045 $X2=2.1
+ $Y2=1.675
r40 3 14 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.1 $Y=0.445 $X2=2.1
+ $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_1%A_40_47# 1 2 3 10 12 15 17 22 25 27 29 35 38
+ 46
c68 25 0 1.96611e-19 $X=0.805 $Y=2.045
r69 36 46 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.73 $Y=1.35
+ $X2=2.885 $Y2=1.35
r70 36 43 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.73 $Y=1.35 $X2=2.64
+ $Y2=1.35
r71 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.73
+ $Y=1.35 $X2=2.73 $Y2=1.35
r72 33 35 24.7562 $w=2.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.7 $Y=1.93 $X2=2.7
+ $Y2=1.35
r73 30 41 1.13371 $w=2.1e-07 $l=1.13e-07 $layer=LI1_cond $X=1.855 $Y=2.035
+ $X2=1.742 $Y2=2.035
r74 30 32 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=1.855 $Y=2.035
+ $X2=1.885 $Y2=2.035
r75 29 33 6.95594 $w=2.1e-07 $l=1.8e-07 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=2.7 $Y2=1.93
r76 29 32 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=1.885 $Y2=2.035
r77 28 38 2.49072 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.96 $Y=1.74
+ $X2=0.812 $Y2=1.74
r78 27 41 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.742 $Y=1.74
+ $X2=1.742 $Y2=2.035
r79 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.63 $Y=1.74
+ $X2=0.96 $Y2=1.74
r80 23 38 3.95216 $w=2.32e-07 $l=8.5e-08 $layer=LI1_cond $X=0.812 $Y=1.825
+ $X2=0.812 $Y2=1.74
r81 23 25 8.59449 $w=2.93e-07 $l=2.2e-07 $layer=LI1_cond $X=0.812 $Y=1.825
+ $X2=0.812 $Y2=2.045
r82 22 38 3.95216 $w=2.32e-07 $l=1.11781e-07 $layer=LI1_cond $X=0.75 $Y=1.655
+ $X2=0.812 $Y2=1.74
r83 21 22 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=0.75 $Y=0.61
+ $X2=0.75 $Y2=1.655
r84 17 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.665 $Y=0.445
+ $X2=0.75 $Y2=0.61
r85 17 19 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.665 $Y=0.445
+ $X2=0.325 $Y2=0.445
r86 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.515
+ $X2=2.885 $Y2=1.35
r87 13 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.885 $Y=1.515
+ $X2=2.885 $Y2=2.465
r88 10 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.185
+ $X2=2.64 $Y2=1.35
r89 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.64 $Y=1.185
+ $X2=2.64 $Y2=0.655
r90 3 32 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=1.835 $X2=1.885 $Y2=2.035
r91 2 25 600 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.835 $X2=0.805 $Y2=2.045
r92 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.235 $X2=0.325 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_1%VPWR 1 2 3 10 12 14 18 22 24 26 33 34 40 43
r29 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 34 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 31 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.67 $Y2=3.33
r36 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 30 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 27 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=3.33
+ $X2=1.295 $Y2=3.33
r40 27 29 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.46 $Y=3.33 $X2=2.16
+ $Y2=3.33
r41 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.67 $Y2=3.33
r42 26 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 20 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=3.33
r46 20 22 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=2.475
r47 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=3.245
+ $X2=1.295 $Y2=3.33
r48 16 18 39.6371 $w=3.28e-07 $l=1.135e-06 $layer=LI1_cond $X=1.295 $Y=3.245
+ $X2=1.295 $Y2=2.11
r49 15 37 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.245 $Y2=3.33
r50 14 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.13 $Y=3.33
+ $X2=1.295 $Y2=3.33
r51 14 15 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.13 $Y=3.33 $X2=0.49
+ $Y2=3.33
r52 10 37 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.325 $Y=3.245
+ $X2=0.245 $Y2=3.33
r53 10 12 41.907 $w=3.28e-07 $l=1.2e-06 $layer=LI1_cond $X=0.325 $Y=3.245
+ $X2=0.325 $Y2=2.045
r54 3 22 300 $w=1.7e-07 $l=8.52291e-07 $layer=licon1_PDIFF $count=2 $X=2.175
+ $Y=1.835 $X2=2.67 $Y2=2.475
r55 2 18 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.155
+ $Y=1.835 $X2=1.295 $Y2=2.11
r56 1 12 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.835 $X2=0.325 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_1%X 1 2 7 8 9 10 11 12 13 37
r15 13 34 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.14 $Y=2.775
+ $X2=3.14 $Y2=2.91
r16 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=2.405
+ $X2=3.14 $Y2=2.775
r17 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.14 $Y=1.98
+ $X2=3.14 $Y2=2.405
r18 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.14 $Y=1.665
+ $X2=3.14 $Y2=1.98
r19 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.665
r20 9 43 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.015
r21 8 43 5.33909 $w=5.83e-07 $l=9e-08 $layer=LI1_cond $X=2.982 $Y=0.925
+ $X2=2.982 $Y2=1.015
r22 7 8 7.56494 $w=5.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.982 $Y=0.555
+ $X2=2.982 $Y2=0.925
r23 7 37 3.47578 $w=5.83e-07 $l=1.7e-07 $layer=LI1_cond $X=2.982 $Y=0.555
+ $X2=2.982 $Y2=0.385
r24 2 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.91
r25 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=1.98
r26 1 37 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=2.715
+ $Y=0.235 $X2=2.855 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_1%VGND 1 6 11 12 13 23 24
r32 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r33 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r34 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 16 20 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r36 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 13 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r38 13 17 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r39 11 20 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.16
+ $Y2=0
r40 11 12 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.385
+ $Y2=0
r41 10 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.52 $Y=0 $X2=3.12
+ $Y2=0
r42 10 12 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.52 $Y=0 $X2=2.385
+ $Y2=0
r43 6 8 20.2745 $w=2.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.385 $Y=0.38
+ $X2=2.385 $Y2=0.855
r44 4 12 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0
r45 4 6 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0.38
r46 1 8 182 $w=1.7e-07 $l=7.30205e-07 $layer=licon1_NDIFF $count=1 $X=2.175
+ $Y=0.235 $X2=2.415 $Y2=0.855
r47 1 6 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.175
+ $Y=0.235 $X2=2.385 $Y2=0.38
.ends

