# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxtp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxtp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.820000 1.600000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 0.265000 8.035000 3.065000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.480000 0.905000 2.150000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.490000 0.445000 1.130000 ;
      RECT 0.115000  1.130000 1.545000 1.300000 ;
      RECT 0.115000  1.300000 0.365000 3.010000 ;
      RECT 0.905000  0.085000 1.235000 0.950000 ;
      RECT 0.935000  2.330000 1.265000 3.245000 ;
      RECT 1.375000  1.300000 1.545000 1.425000 ;
      RECT 1.375000  1.425000 3.310000 1.585000 ;
      RECT 1.375000  1.585000 4.270000 1.595000 ;
      RECT 1.725000  0.490000 2.055000 1.075000 ;
      RECT 1.725000  1.075000 3.880000 1.245000 ;
      RECT 1.725000  2.330000 2.055000 3.010000 ;
      RECT 1.885000  1.965000 3.730000 2.135000 ;
      RECT 1.885000  2.135000 2.055000 2.330000 ;
      RECT 2.295000  2.435000 2.625000 2.475000 ;
      RECT 2.295000  2.475000 4.895000 2.645000 ;
      RECT 2.295000  2.645000 2.625000 3.065000 ;
      RECT 2.465000  0.265000 2.795000 0.725000 ;
      RECT 2.465000  0.725000 4.275000 0.855000 ;
      RECT 2.465000  0.855000 4.620000 0.895000 ;
      RECT 2.980000  1.595000 4.270000 1.755000 ;
      RECT 3.195000  2.825000 3.525000 3.245000 ;
      RECT 3.285000  0.085000 3.615000 0.545000 ;
      RECT 3.400000  2.135000 3.730000 2.295000 ;
      RECT 3.550000  1.245000 3.880000 1.405000 ;
      RECT 3.940000  1.755000 4.270000 1.975000 ;
      RECT 4.095000  2.825000 5.245000 3.035000 ;
      RECT 4.105000  0.895000 4.620000 1.185000 ;
      RECT 4.450000  1.185000 4.620000 2.185000 ;
      RECT 4.450000  2.185000 4.895000 2.475000 ;
      RECT 4.455000  0.265000 4.785000 0.505000 ;
      RECT 4.455000  0.505000 4.970000 0.675000 ;
      RECT 4.800000  0.675000 4.970000 1.435000 ;
      RECT 4.800000  1.435000 6.170000 1.605000 ;
      RECT 5.075000  1.605000 5.245000 2.825000 ;
      RECT 5.150000  0.925000 6.685000 1.095000 ;
      RECT 5.150000  1.095000 5.480000 1.255000 ;
      RECT 5.280000  0.085000 5.610000 0.675000 ;
      RECT 5.565000  1.815000 5.895000 3.245000 ;
      RECT 5.840000  1.275000 6.170000 1.435000 ;
      RECT 6.355000  0.265000 6.685000 0.925000 ;
      RECT 6.355000  1.095000 6.685000 1.305000 ;
      RECT 6.355000  1.305000 7.525000 1.635000 ;
      RECT 6.355000  1.635000 6.685000 3.065000 ;
      RECT 6.915000  0.085000 7.245000 1.125000 ;
      RECT 6.915000  1.815000 7.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__dlxtp_lp
END LIBRARY
