* NGSPICE file created from sky130_fd_sc_lp__dlrtp_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlrtp_lp D GATE RESET_B VGND VNB VPB VPWR Q
M1000 VPWR a_638_73# a_800_343# VPB phighvt w=640000u l=150000u
+  ad=1.4461e+12p pd=1.238e+07u as=3.648e+11p ps=3.7e+06u
M1001 a_186_57# GATE a_114_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1002 VGND a_186_57# a_408_73# VNB nshort w=420000u l=150000u
+  ad=1.3923e+12p pd=8.44e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_1420_367# a_887_343# a_1208_75# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.182e+11p pd=6.18e+06u as=3.528e+11p ps=3.08e+06u
M1004 a_384_345# a_186_57# a_294_547# VPB phighvt w=640000u l=150000u
+  ad=2.304e+11p pd=2e+06u as=1.824e+11p ps=1.85e+06u
M1005 VPWR a_186_57# a_384_345# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_408_73# a_186_57# a_294_547# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.086e+11p ps=1.92e+06u
M1007 Q a_1208_75# a_1857_47# VNB nshort w=840000u l=150000u
+  ad=2.604e+11p pd=2.3e+06u as=1.764e+11p ps=2.1e+06u
M1008 a_617_345# D VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1009 a_996_343# a_1208_75# VPWR VPB phighvt w=420000u l=150000u
+  ad=2.394e+11p pd=2.82e+06u as=0p ps=0u
M1010 a_114_57# GATE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_638_73# D a_617_345# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1012 a_1593_367# RESET_B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1013 a_1208_75# RESET_B a_1593_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_638_73# a_1058_101# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1015 a_1510_47# a_887_343# a_1208_75# VNB nshort w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=2.394e+11p ps=2.25e+06u
M1016 a_1857_47# a_1208_75# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_887_343# a_186_57# a_800_343# VPB phighvt w=640000u l=150000u
+  ad=2.286e+11p pd=2.07e+06u as=0p ps=0u
M1018 a_186_57# GATE a_114_470# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.344e+11p ps=1.7e+06u
M1019 a_566_73# D VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1020 a_638_73# D a_566_73# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1021 VGND RESET_B a_1510_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_114_470# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1949_367# a_1208_75# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.024e+11p pd=3e+06u as=0p ps=0u
M1024 Q a_1208_75# a_1949_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1025 VPWR a_887_343# a_1420_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1058_101# a_294_547# a_887_343# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1027 a_996_343# a_294_547# a_887_343# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_887_343# a_186_57# a_862_101# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.877e+11p ps=3.05e+06u
M1029 a_862_101# a_1208_75# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

