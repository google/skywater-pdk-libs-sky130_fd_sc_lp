* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or2b_lp A B_N VGND VNB VPB VPWR X
X0 a_397_409# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_30_57# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_275_57# a_30_57# a_290_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_597_57# a_290_409# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_290_409# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_439_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_290_409# A a_439_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_117_57# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_30_57# B_N a_117_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_30_57# a_275_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_290_409# a_30_57# a_397_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VGND a_290_409# a_597_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
