* File: sky130_fd_sc_lp__nand2_1.pex.spice
* Created: Fri Aug 28 10:46:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_1%B 3 6 8 9 13 15
c22 8 0 1.75086e-19 $X=0.24 $Y=1.295
r23 13 16 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.46
+ $X2=0.362 $Y2=1.625
r24 13 15 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.46
+ $X2=0.362 $Y2=1.295
r25 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.46 $X2=0.33 $Y2=1.46
r26 9 14 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.46
r27 8 14 5.43295 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.46
r28 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.485 $Y=2.465
+ $X2=0.485 $Y2=1.625
r29 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.485 $Y=0.765
+ $X2=0.485 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_1%A 1 3 6 8 9 13
c24 1 0 1.75086e-19 $X=0.875 $Y=1.295
r25 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.46 $X2=1.07 $Y2=1.46
r26 13 15 23.869 $w=3.13e-07 $l=1.55e-07 $layer=POLY_cond $X=0.915 $Y=1.46
+ $X2=1.07 $Y2=1.46
r27 12 13 6.15974 $w=3.13e-07 $l=4e-08 $layer=POLY_cond $X=0.875 $Y=1.46
+ $X2=0.915 $Y2=1.46
r28 9 16 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.46
r29 8 16 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=1.295
+ $X2=1.17 $Y2=1.46
r30 4 13 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.625
+ $X2=0.915 $Y2=1.46
r31 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.915 $Y=1.625
+ $X2=0.915 $Y2=2.465
r32 1 12 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.875 $Y=1.295
+ $X2=0.875 $Y2=1.46
r33 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.875 $Y=1.295
+ $X2=0.875 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_1%VPWR 1 2 7 9 13 15 19 21 31
r22 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r23 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 22 27 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r25 22 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 21 30 4.49223 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.212 $Y2=3.33
r27 21 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 19 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r29 19 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 19 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 15 18 32.1569 $w=3.08e-07 $l=8.65e-07 $layer=LI1_cond $X=1.14 $Y=2.085
+ $X2=1.14 $Y2=2.95
r32 13 30 3.10696 $w=3.1e-07 $l=1.15521e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.212 $Y2=3.33
r33 13 18 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.95
r34 9 12 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.27 $Y=2.005
+ $X2=0.27 $Y2=2.95
r35 7 27 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r36 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.95
r37 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=2.95
r38 2 15 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=2.085
r39 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.95
r40 1 9 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_1%Y 1 2 7 8 9 10 11 12 13 37
c17 9 0 2.39113e-20 $X=0.72 $Y=1.295
r18 13 34 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.71 $Y=2.775
+ $X2=0.71 $Y2=2.91
r19 12 13 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.405
+ $X2=0.71 $Y2=2.775
r20 11 12 22.4459 $w=2.08e-07 $l=4.25e-07 $layer=LI1_cond $X=0.71 $Y=1.98
+ $X2=0.71 $Y2=2.405
r21 10 11 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.71 $Y2=1.98
r22 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.665
r23 9 43 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.04
r24 8 43 8.04582 $w=6.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.93 $Y=0.925
+ $X2=0.93 $Y2=1.04
r25 7 8 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.93 $Y=0.555 $X2=0.93
+ $Y2=0.925
r26 7 37 0.552036 $w=6.48e-07 $l=3e-08 $layer=LI1_cond $X=0.93 $Y=0.555 $X2=0.93
+ $Y2=0.525
r27 2 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.91
r28 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=1.98
r29 1 37 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=0.95 $Y=0.345
+ $X2=1.09 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_1%VGND 1 4 6 8 12 13
r14 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r15 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r16 10 16 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r17 10 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=1.2
+ $Y2=0
r18 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r19 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r20 4 16 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r21 4 6 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.49
r22 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.345 $X2=0.27 $Y2=0.49
.ends

