* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtp_lp2 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_658_47# a_413_47# a_736_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_122# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_500_47# a_256_405# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_736_47# a_256_405# a_850_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_898_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_1216_57# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_898_21# a_1380_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_413_47# a_256_405# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VPWR a_736_47# a_898_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VPWR a_898_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND a_27_122# a_658_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR GATE a_256_405# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_850_47# a_898_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_413_47# a_256_405# a_500_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_736_47# a_413_47# a_944_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_294_185# GATE a_256_405# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_898_21# a_736_47# a_1216_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_122# D a_114_122# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_740_419# a_256_405# a_736_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 VGND GATE a_294_185# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_944_419# a_898_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_1380_57# a_898_21# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR a_27_122# a_740_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X23 a_114_122# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
