* File: sky130_fd_sc_lp__o211a_4.pxi.spice
* Created: Wed Sep  2 10:14:00 2020
* 
x_PM_SKY130_FD_SC_LP__O211A_4%A_80_21# N_A_80_21#_M1016_d N_A_80_21#_M1005_s
+ N_A_80_21#_M1022_s N_A_80_21#_M1007_s N_A_80_21#_M1011_g N_A_80_21#_M1002_g
+ N_A_80_21#_M1014_g N_A_80_21#_M1009_g N_A_80_21#_M1015_g N_A_80_21#_M1012_g
+ N_A_80_21#_M1023_g N_A_80_21#_M1021_g N_A_80_21#_c_209_p N_A_80_21#_c_120_n
+ N_A_80_21#_c_121_n N_A_80_21#_c_122_n N_A_80_21#_c_123_n N_A_80_21#_c_134_p
+ N_A_80_21#_c_178_p N_A_80_21#_c_140_p N_A_80_21#_c_138_p N_A_80_21#_c_168_p
+ N_A_80_21#_c_124_n N_A_80_21#_c_150_p N_A_80_21#_c_125_n N_A_80_21#_c_142_p
+ N_A_80_21#_c_126_n PM_SKY130_FD_SC_LP__O211A_4%A_80_21#
x_PM_SKY130_FD_SC_LP__O211A_4%B1 N_B1_M1005_g N_B1_M1004_g N_B1_M1008_g
+ N_B1_M1017_g N_B1_c_280_n N_B1_c_263_n N_B1_c_264_n B1 B1 N_B1_c_265_n
+ N_B1_c_266_n PM_SKY130_FD_SC_LP__O211A_4%B1
x_PM_SKY130_FD_SC_LP__O211A_4%C1 N_C1_M1016_g N_C1_M1010_g N_C1_M1020_g
+ N_C1_M1022_g C1 N_C1_c_348_n N_C1_c_349_n PM_SKY130_FD_SC_LP__O211A_4%C1
x_PM_SKY130_FD_SC_LP__O211A_4%A1 N_A1_M1001_g N_A1_M1000_g N_A1_c_395_n
+ N_A1_M1003_g N_A1_M1019_g N_A1_c_397_n N_A1_c_398_n N_A1_c_399_n A1 A1
+ N_A1_c_400_n N_A1_c_401_n N_A1_c_402_n A1 PM_SKY130_FD_SC_LP__O211A_4%A1
x_PM_SKY130_FD_SC_LP__O211A_4%A2 N_A2_M1006_g N_A2_M1007_g N_A2_M1018_g
+ N_A2_M1013_g A2 A2 N_A2_c_468_n PM_SKY130_FD_SC_LP__O211A_4%A2
x_PM_SKY130_FD_SC_LP__O211A_4%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_M1021_d
+ N_VPWR_M1010_d N_VPWR_M1017_d N_VPWR_M1019_s N_VPWR_c_519_n N_VPWR_c_520_n
+ N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n
+ N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n VPWR
+ N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n
+ N_VPWR_c_535_n N_VPWR_c_536_n N_VPWR_c_518_n PM_SKY130_FD_SC_LP__O211A_4%VPWR
x_PM_SKY130_FD_SC_LP__O211A_4%X N_X_M1011_d N_X_M1015_d N_X_M1002_s N_X_M1012_s
+ N_X_c_614_n N_X_c_619_n N_X_c_620_n N_X_c_664_p N_X_c_615_n N_X_c_652_n
+ N_X_c_621_n N_X_c_663_p N_X_c_656_n N_X_c_616_n N_X_c_622_n X X N_X_c_617_n X
+ PM_SKY130_FD_SC_LP__O211A_4%X
x_PM_SKY130_FD_SC_LP__O211A_4%A_986_367# N_A_986_367#_M1000_d
+ N_A_986_367#_M1013_d N_A_986_367#_c_670_n N_A_986_367#_c_680_n
+ N_A_986_367#_c_675_n PM_SKY130_FD_SC_LP__O211A_4%A_986_367#
x_PM_SKY130_FD_SC_LP__O211A_4%VGND N_VGND_M1011_s N_VGND_M1014_s N_VGND_M1023_s
+ N_VGND_M1001_d N_VGND_M1018_s N_VGND_c_682_n N_VGND_c_683_n N_VGND_c_684_n
+ N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n N_VGND_c_689_n
+ N_VGND_c_690_n N_VGND_c_691_n VGND N_VGND_c_692_n N_VGND_c_693_n
+ N_VGND_c_694_n N_VGND_c_695_n N_VGND_c_696_n N_VGND_c_697_n
+ PM_SKY130_FD_SC_LP__O211A_4%VGND
x_PM_SKY130_FD_SC_LP__O211A_4%A_475_49# N_A_475_49#_M1004_d N_A_475_49#_M1008_d
+ N_A_475_49#_M1006_d N_A_475_49#_M1003_s N_A_475_49#_c_780_n
+ N_A_475_49#_c_781_n N_A_475_49#_c_787_n N_A_475_49#_c_828_n
+ N_A_475_49#_c_799_n N_A_475_49#_c_803_n N_A_475_49#_c_782_n
+ N_A_475_49#_c_783_n N_A_475_49#_c_793_n N_A_475_49#_c_810_n
+ PM_SKY130_FD_SC_LP__O211A_4%A_475_49#
x_PM_SKY130_FD_SC_LP__O211A_4%A_574_49# N_A_574_49#_M1004_s N_A_574_49#_M1020_s
+ N_A_574_49#_c_849_n PM_SKY130_FD_SC_LP__O211A_4%A_574_49#
cc_1 VNB N_A_80_21#_M1011_g 0.0258622f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_80_21#_M1002_g 5.40282e-19 $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.465
cc_3 VNB N_A_80_21#_M1014_g 0.0213903f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_4 VNB N_A_80_21#_M1009_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=2.465
cc_5 VNB N_A_80_21#_M1015_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_6 VNB N_A_80_21#_M1012_g 4.57047e-19 $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.465
cc_7 VNB N_A_80_21#_M1023_g 0.0273509f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_8 VNB N_A_80_21#_M1021_g 3.92279e-19 $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=2.465
cc_9 VNB N_A_80_21#_c_120_n 0.00246091f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.385
cc_10 VNB N_A_80_21#_c_121_n 3.99447e-19 $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=2.27
cc_11 VNB N_A_80_21#_c_122_n 0.0102249f $X=-0.19 $Y=-0.245 $X2=3.37 $Y2=1.15
cc_12 VNB N_A_80_21#_c_123_n 0.00796633f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=1.15
cc_13 VNB N_A_80_21#_c_124_n 0.00128591f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.485
cc_14 VNB N_A_80_21#_c_125_n 0.00482819f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=1.07
cc_15 VNB N_A_80_21#_c_126_n 0.114836f $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=1.48
cc_16 VNB N_B1_M1004_g 0.0285557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_M1008_g 0.0253654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_263_n 0.00243414f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.315
cc_19 VNB N_B1_c_264_n 0.0268304f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_20 VNB N_B1_c_265_n 0.0309123f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=1.645
cc_21 VNB N_B1_c_266_n 0.00258833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C1_M1016_g 0.0253344f $X=-0.19 $Y=-0.245 $X2=3.92 $Y2=1.835
cc_23 VNB N_C1_M1020_g 0.0268186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C1_c_348_n 0.00165536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_349_n 0.0405384f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.645
cc_26 VNB N_A1_M1000_g 0.00714672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_c_395_n 0.0196339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_M1019_g 0.00655341f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.315
cc_29 VNB N_A1_c_397_n 0.0199104f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_30 VNB N_A1_c_398_n 0.0136012f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.645
cc_31 VNB N_A1_c_399_n 0.0292611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_c_400_n 0.0179104f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=2.465
cc_33 VNB N_A1_c_401_n 0.0565587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_c_402_n 0.0117338f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.465
cc_35 VNB A1 0.0155807f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.315
cc_36 VNB N_A2_M1006_g 0.0230873f $X=-0.19 $Y=-0.245 $X2=3.92 $Y2=1.835
cc_37 VNB N_A2_M1018_g 0.0225714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB A2 0.00487676f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.465
cc_39 VNB N_A2_c_468_n 0.0301718f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=2.465
cc_40 VNB N_VPWR_c_518_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_614_n 7.8818e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.315
cc_42 VNB N_X_c_615_n 0.00615641f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.315
cc_43 VNB N_X_c_616_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=2.465
cc_44 VNB N_X_c_617_n 0.0084917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB X 0.0230986f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.48
cc_46 VNB N_VGND_c_682_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_683_n 0.0276525f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.465
cc_48 VNB N_VGND_c_684_n 3.15212e-19 $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_49 VNB N_VGND_c_685_n 0.00444657f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=2.465
cc_50 VNB N_VGND_c_686_n 0.00538269f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_51 VNB N_VGND_c_687_n 0.00450476f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.465
cc_52 VNB N_VGND_c_688_n 0.0150063f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.315
cc_53 VNB N_VGND_c_689_n 0.00452017f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_54 VNB N_VGND_c_690_n 0.0167176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_691_n 0.00362148f $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=1.645
cc_56 VNB N_VGND_c_692_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_693_n 0.0662037f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.235
cc_58 VNB N_VGND_c_694_n 0.020434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_695_n 0.342092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_696_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_697_n 0.00631724f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=2.435
cc_62 VNB N_A_475_49#_c_780_n 0.00290338f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.315
cc_63 VNB N_A_475_49#_c_781_n 0.00394846f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_64 VNB N_A_475_49#_c_782_n 0.00742799f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.315
cc_65 VNB N_A_475_49#_c_783_n 0.0192135f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=1.645
cc_66 VPB N_A_80_21#_M1002_g 0.0229919f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.465
cc_67 VPB N_A_80_21#_M1009_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=2.465
cc_68 VPB N_A_80_21#_M1012_g 0.0189066f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.465
cc_69 VPB N_A_80_21#_M1021_g 0.0187821f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=2.465
cc_70 VPB N_A_80_21#_c_121_n 0.00106148f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=2.27
cc_71 VPB N_B1_M1005_g 0.021201f $X=-0.19 $Y=1.655 $X2=3.92 $Y2=1.835
cc_72 VPB N_B1_M1017_g 0.0199923f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_73 VPB N_B1_c_263_n 0.00136973f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.315
cc_74 VPB N_B1_c_264_n 0.00656712f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.655
cc_75 VPB N_B1_c_265_n 0.00994084f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.645
cc_76 VPB N_B1_c_266_n 0.00131738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_C1_M1010_g 0.0215331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_C1_M1022_g 0.0191428f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_79 VPB N_C1_c_348_n 0.00334818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_C1_c_349_n 0.0103231f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=1.645
cc_81 VPB N_A1_M1000_g 0.0209526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A1_M1019_g 0.0239995f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.315
cc_83 VPB A1 0.011538f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.315
cc_84 VPB N_A2_M1007_g 0.0182425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A2_M1013_g 0.0182425f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_86 VPB A2 0.00905439f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.465
cc_87 VPB N_A2_c_468_n 0.00462236f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=2.465
cc_88 VPB N_VPWR_c_519_n 0.0415014f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.315
cc_89 VPB N_VPWR_c_520_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.295 $Y2=2.465
cc_90 VPB N_VPWR_c_521_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.645
cc_91 VPB N_VPWR_c_522_n 4.21859e-19 $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.315
cc_92 VPB N_VPWR_c_523_n 0.00468074f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=1.645
cc_93 VPB N_VPWR_c_524_n 0.0135296f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=2.465
cc_94 VPB N_VPWR_c_525_n 0.0479716f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=1.485
cc_95 VPB N_VPWR_c_526_n 0.0130339f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=1.485
cc_96 VPB N_VPWR_c_527_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=1.48
cc_97 VPB N_VPWR_c_528_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.235
cc_98 VPB N_VPWR_c_529_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.385
cc_99 VPB N_VPWR_c_530_n 0.017577f $X=-0.19 $Y=1.655 $X2=3.37 $Y2=1.15
cc_100 VPB N_VPWR_c_531_n 0.0219055f $X=-0.19 $Y=1.655 $X2=5.5 $Y2=2.27
cc_101 VPB N_VPWR_c_532_n 0.0172367f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.485
cc_102 VPB N_VPWR_c_533_n 0.0344653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_534_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.48
cc_104 VPB N_VPWR_c_535_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.48
cc_105 VPB N_VPWR_c_536_n 0.00506799f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=1.48
cc_106 VPB N_VPWR_c_518_n 0.0647765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_X_c_619_n 0.00879192f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_108 VPB N_X_c_620_n 0.0202382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_X_c_621_n 0.0051731f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.315
cc_110 VPB N_X_c_622_n 0.00135109f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=2.465
cc_111 VPB X 0.00588455f $X=-0.19 $Y=1.655 $X2=2.065 $Y2=1.48
cc_112 N_A_80_21#_M1021_g N_B1_M1005_g 0.049111f $X=2.155 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_121_n N_B1_M1005_g 0.00617979f $X=2.29 $Y=2.27 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_134_p N_B1_M1005_g 0.0132818f $X=2.705 $Y=2.355 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_120_n N_B1_M1004_g 0.00280505f $X=2.29 $Y=1.385 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_122_n N_B1_M1004_g 0.0127694f $X=3.37 $Y=1.15 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_126_n N_B1_M1004_g 5.56414e-19 $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_138_p N_B1_M1017_g 0.013108f $X=5.335 $Y=2.355 $X2=0 $Y2=0
cc_119 N_A_80_21#_M1022_s N_B1_c_280_n 0.00903518f $X=3.92 $Y=1.835 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_140_p N_B1_c_280_n 0.0323573f $X=3.965 $Y=2.355 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_138_p N_B1_c_280_n 0.0113161f $X=5.335 $Y=2.355 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_142_p N_B1_c_280_n 0.0234562f $X=4.13 $Y=2.435 $X2=0 $Y2=0
cc_123 N_A_80_21#_M1022_s N_B1_c_263_n 0.00121536f $X=3.92 $Y=1.835 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_142_p N_B1_c_264_n 4.96417e-19 $X=4.13 $Y=2.435 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_120_n N_B1_c_265_n 9.2064e-19 $X=2.29 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_121_n N_B1_c_265_n 6.06247e-19 $X=2.29 $Y=2.27 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_122_n N_B1_c_265_n 0.00917258f $X=3.37 $Y=1.15 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_134_p N_B1_c_265_n 0.00105558f $X=2.705 $Y=2.355 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_124_n N_B1_c_265_n 0.00205621f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_150_p N_B1_c_265_n 5.48245e-19 $X=3.2 $Y=2.435 $X2=0 $Y2=0
cc_131 N_A_80_21#_c_126_n N_B1_c_265_n 0.0208478f $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_132 N_A_80_21#_M1005_s N_B1_c_266_n 0.0117523f $X=2.66 $Y=1.835 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_121_n N_B1_c_266_n 0.0406477f $X=2.29 $Y=2.27 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_122_n N_B1_c_266_n 0.0583903f $X=3.37 $Y=1.15 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_134_p N_B1_c_266_n 0.00869878f $X=2.705 $Y=2.355 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_124_n N_B1_c_266_n 0.0159566f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_150_p N_B1_c_266_n 0.0507731f $X=3.2 $Y=2.435 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_126_n N_B1_c_266_n 6.16322e-19 $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_122_n N_C1_M1016_g 0.0111502f $X=3.37 $Y=1.15 $X2=0 $Y2=0
cc_140 N_A_80_21#_c_125_n N_C1_M1016_g 0.0030784f $X=3.535 $Y=1.07 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_140_p N_C1_M1010_g 0.0122595f $X=3.965 $Y=2.355 $X2=0 $Y2=0
cc_142 N_A_80_21#_c_125_n N_C1_M1020_g 0.00687255f $X=3.535 $Y=1.07 $X2=0 $Y2=0
cc_143 N_A_80_21#_c_140_p N_C1_M1022_g 0.0148598f $X=3.965 $Y=2.355 $X2=0 $Y2=0
cc_144 N_A_80_21#_c_125_n N_C1_c_348_n 0.019933f $X=3.535 $Y=1.07 $X2=0 $Y2=0
cc_145 N_A_80_21#_c_150_p N_C1_c_349_n 4.1502e-19 $X=3.2 $Y=2.435 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_125_n N_C1_c_349_n 0.00883401f $X=3.535 $Y=1.07 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_138_p N_A1_M1000_g 0.020011f $X=5.335 $Y=2.355 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_168_p N_A1_M1000_g 0.00165521f $X=5.5 $Y=2.035 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_138_p N_A2_M1007_g 0.0137596f $X=5.335 $Y=2.355 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_168_p N_A2_M1007_g 0.00699617f $X=5.5 $Y=2.035 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_138_p N_A2_M1013_g 0.00420364f $X=5.335 $Y=2.355 $X2=0 $Y2=0
cc_152 N_A_80_21#_c_168_p N_A2_M1013_g 0.00422842f $X=5.5 $Y=2.035 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_138_p A2 0.00363086f $X=5.335 $Y=2.355 $X2=0 $Y2=0
cc_154 N_A_80_21#_c_168_p A2 0.022935f $X=5.5 $Y=2.035 $X2=0 $Y2=0
cc_155 N_A_80_21#_c_168_p N_A2_c_468_n 6.34554e-19 $X=5.5 $Y=2.035 $X2=0 $Y2=0
cc_156 N_A_80_21#_c_121_n N_VPWR_M1021_d 0.00411051f $X=2.29 $Y=2.27 $X2=0 $Y2=0
cc_157 N_A_80_21#_c_134_p N_VPWR_M1021_d 0.00347755f $X=2.705 $Y=2.355 $X2=0
+ $Y2=0
cc_158 N_A_80_21#_c_178_p N_VPWR_M1021_d 9.62763e-19 $X=2.375 $Y=2.355 $X2=0
+ $Y2=0
cc_159 N_A_80_21#_c_140_p N_VPWR_M1010_d 0.00344105f $X=3.965 $Y=2.355 $X2=0
+ $Y2=0
cc_160 N_A_80_21#_c_138_p N_VPWR_M1017_d 0.0100499f $X=5.335 $Y=2.355 $X2=0
+ $Y2=0
cc_161 N_A_80_21#_M1002_g N_VPWR_c_519_n 0.0152824f $X=0.865 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_80_21#_M1009_g N_VPWR_c_519_n 7.27171e-19 $X=1.295 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_80_21#_M1002_g N_VPWR_c_520_n 7.42371e-19 $X=0.865 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_80_21#_M1009_g N_VPWR_c_520_n 0.0144441f $X=1.295 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_80_21#_M1012_g N_VPWR_c_520_n 0.0142189f $X=1.725 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_80_21#_M1021_g N_VPWR_c_520_n 7.27171e-19 $X=2.155 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_80_21#_M1012_g N_VPWR_c_521_n 5.81474e-19 $X=1.725 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_80_21#_M1021_g N_VPWR_c_521_n 0.0109892f $X=2.155 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_80_21#_c_134_p N_VPWR_c_521_n 0.00809557f $X=2.705 $Y=2.355 $X2=0
+ $Y2=0
cc_170 N_A_80_21#_c_178_p N_VPWR_c_521_n 0.00987845f $X=2.375 $Y=2.355 $X2=0
+ $Y2=0
cc_171 N_A_80_21#_c_140_p N_VPWR_c_522_n 0.0170777f $X=3.965 $Y=2.355 $X2=0
+ $Y2=0
cc_172 N_A_80_21#_c_138_p N_VPWR_c_523_n 0.0167599f $X=5.335 $Y=2.355 $X2=0
+ $Y2=0
cc_173 N_A_80_21#_M1002_g N_VPWR_c_526_n 0.00486043f $X=0.865 $Y=2.465 $X2=0
+ $Y2=0
cc_174 N_A_80_21#_M1009_g N_VPWR_c_526_n 0.00486043f $X=1.295 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_80_21#_M1012_g N_VPWR_c_528_n 0.00486043f $X=1.725 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_80_21#_M1021_g N_VPWR_c_528_n 0.00486043f $X=2.155 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_80_21#_c_150_p N_VPWR_c_531_n 0.0405775f $X=3.2 $Y=2.435 $X2=0 $Y2=0
cc_178 N_A_80_21#_c_142_p N_VPWR_c_532_n 0.0214287f $X=4.13 $Y=2.435 $X2=0 $Y2=0
cc_179 N_A_80_21#_M1005_s N_VPWR_c_518_n 0.00869072f $X=2.66 $Y=1.835 $X2=0
+ $Y2=0
cc_180 N_A_80_21#_M1022_s N_VPWR_c_518_n 0.0050864f $X=3.92 $Y=1.835 $X2=0 $Y2=0
cc_181 N_A_80_21#_M1007_s N_VPWR_c_518_n 0.00225186f $X=5.36 $Y=1.835 $X2=0
+ $Y2=0
cc_182 N_A_80_21#_M1002_g N_VPWR_c_518_n 0.00824727f $X=0.865 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_80_21#_M1009_g N_VPWR_c_518_n 0.00824727f $X=1.295 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_80_21#_M1012_g N_VPWR_c_518_n 0.00824727f $X=1.725 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_80_21#_M1021_g N_VPWR_c_518_n 0.00824727f $X=2.155 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_80_21#_c_150_p N_VPWR_c_518_n 0.0228601f $X=3.2 $Y=2.435 $X2=0 $Y2=0
cc_187 N_A_80_21#_c_142_p N_VPWR_c_518_n 0.0129463f $X=4.13 $Y=2.435 $X2=0 $Y2=0
cc_188 N_A_80_21#_M1011_g N_X_c_614_n 0.0166141f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A_80_21#_c_209_p N_X_c_614_n 0.00390667f $X=2.205 $Y=1.485 $X2=0 $Y2=0
cc_190 N_A_80_21#_M1002_g N_X_c_619_n 0.0152068f $X=0.865 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_80_21#_c_209_p N_X_c_619_n 0.0316102f $X=2.205 $Y=1.485 $X2=0 $Y2=0
cc_192 N_A_80_21#_c_126_n N_X_c_619_n 0.0112018f $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_193 N_A_80_21#_M1014_g N_X_c_615_n 0.0138879f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A_80_21#_M1015_g N_X_c_615_n 0.0135912f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_80_21#_M1023_g N_X_c_615_n 0.00214629f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A_80_21#_c_209_p N_X_c_615_n 0.0636118f $X=2.205 $Y=1.485 $X2=0 $Y2=0
cc_197 N_A_80_21#_c_123_n N_X_c_615_n 0.00591517f $X=2.375 $Y=1.15 $X2=0 $Y2=0
cc_198 N_A_80_21#_c_126_n N_X_c_615_n 0.00531191f $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_199 N_A_80_21#_M1009_g N_X_c_621_n 0.0131657f $X=1.295 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A_80_21#_M1012_g N_X_c_621_n 0.0130035f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A_80_21#_M1021_g N_X_c_621_n 6.55961e-19 $X=2.155 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A_80_21#_c_209_p N_X_c_621_n 0.0635203f $X=2.205 $Y=1.485 $X2=0 $Y2=0
cc_203 N_A_80_21#_c_121_n N_X_c_621_n 0.00947164f $X=2.29 $Y=2.27 $X2=0 $Y2=0
cc_204 N_A_80_21#_c_126_n N_X_c_621_n 0.00508005f $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_205 N_A_80_21#_c_209_p N_X_c_616_n 0.0154947f $X=2.205 $Y=1.485 $X2=0 $Y2=0
cc_206 N_A_80_21#_c_126_n N_X_c_616_n 0.00253619f $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_207 N_A_80_21#_c_209_p N_X_c_622_n 0.0146791f $X=2.205 $Y=1.485 $X2=0 $Y2=0
cc_208 N_A_80_21#_c_126_n N_X_c_622_n 0.00267368f $X=2.155 $Y=1.48 $X2=0 $Y2=0
cc_209 N_A_80_21#_M1011_g X 0.0171501f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A_80_21#_M1002_g X 0.00304876f $X=0.865 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_80_21#_c_209_p X 0.0164313f $X=2.205 $Y=1.485 $X2=0 $Y2=0
cc_212 N_A_80_21#_c_138_p N_A_986_367#_M1000_d 0.00878113f $X=5.335 $Y=2.355
+ $X2=-0.19 $Y2=-0.245
cc_213 N_A_80_21#_M1007_s N_A_986_367#_c_670_n 0.00338033f $X=5.36 $Y=1.835
+ $X2=0 $Y2=0
cc_214 N_A_80_21#_c_138_p N_A_986_367#_c_670_n 0.0307611f $X=5.335 $Y=2.355
+ $X2=0 $Y2=0
cc_215 N_A_80_21#_M1011_g N_VGND_c_683_n 0.0116447f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_216 N_A_80_21#_M1014_g N_VGND_c_683_n 6.25324e-19 $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_217 N_A_80_21#_M1011_g N_VGND_c_684_n 6.25324e-19 $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_218 N_A_80_21#_M1014_g N_VGND_c_684_n 0.0109423f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_219 N_A_80_21#_M1015_g N_VGND_c_684_n 0.0110229f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_220 N_A_80_21#_M1023_g N_VGND_c_684_n 6.39544e-19 $X=1.765 $Y=0.655 $X2=0
+ $Y2=0
cc_221 N_A_80_21#_M1023_g N_VGND_c_685_n 0.0034594f $X=1.765 $Y=0.655 $X2=0
+ $Y2=0
cc_222 N_A_80_21#_c_209_p N_VGND_c_685_n 0.00783521f $X=2.205 $Y=1.485 $X2=0
+ $Y2=0
cc_223 N_A_80_21#_c_126_n N_VGND_c_685_n 0.00514029f $X=2.155 $Y=1.48 $X2=0
+ $Y2=0
cc_224 N_A_80_21#_M1015_g N_VGND_c_688_n 0.00486043f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_A_80_21#_M1023_g N_VGND_c_688_n 0.00585385f $X=1.765 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_A_80_21#_M1011_g N_VGND_c_692_n 0.00486043f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_A_80_21#_M1014_g N_VGND_c_692_n 0.00486043f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_228 N_A_80_21#_M1016_d N_VGND_c_695_n 0.0037799f $X=3.3 $Y=0.245 $X2=0 $Y2=0
cc_229 N_A_80_21#_M1011_g N_VGND_c_695_n 0.00824727f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_A_80_21#_M1014_g N_VGND_c_695_n 0.00824727f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_231 N_A_80_21#_M1015_g N_VGND_c_695_n 0.00824727f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_232 N_A_80_21#_M1023_g N_VGND_c_695_n 0.0118221f $X=1.765 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_80_21#_c_122_n N_A_475_49#_M1004_d 0.00322334f $X=3.37 $Y=1.15
+ $X2=-0.19 $Y2=-0.245
cc_234 N_A_80_21#_c_122_n N_A_475_49#_c_780_n 0.0232791f $X=3.37 $Y=1.15 $X2=0
+ $Y2=0
cc_235 N_A_80_21#_c_123_n N_A_475_49#_c_780_n 0.00373133f $X=2.375 $Y=1.15 $X2=0
+ $Y2=0
cc_236 N_A_80_21#_M1016_d N_A_475_49#_c_787_n 0.00829257f $X=3.3 $Y=0.245 $X2=0
+ $Y2=0
cc_237 N_A_80_21#_c_122_n N_A_475_49#_c_787_n 0.0239892f $X=3.37 $Y=1.15 $X2=0
+ $Y2=0
cc_238 N_A_80_21#_c_125_n N_A_475_49#_c_787_n 0.0247293f $X=3.535 $Y=1.07 $X2=0
+ $Y2=0
cc_239 N_A_80_21#_c_122_n N_A_574_49#_M1004_s 0.00214083f $X=3.37 $Y=1.15
+ $X2=-0.19 $Y2=-0.245
cc_240 N_A_80_21#_M1016_d N_A_574_49#_c_849_n 0.00843896f $X=3.3 $Y=0.245 $X2=0
+ $Y2=0
cc_241 N_B1_M1004_g N_C1_M1016_g 0.0430691f $X=2.795 $Y=0.665 $X2=0 $Y2=0
cc_242 N_B1_M1005_g N_C1_M1010_g 0.0100484f $X=2.585 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_c_280_n N_C1_M1010_g 0.0150206f $X=4.13 $Y=2.015 $X2=0 $Y2=0
cc_244 N_B1_c_266_n N_C1_M1010_g 0.00711889f $X=3.275 $Y=1.752 $X2=0 $Y2=0
cc_245 N_B1_M1008_g N_C1_M1020_g 0.0426468f $X=4.275 $Y=0.665 $X2=0 $Y2=0
cc_246 N_B1_M1017_g N_C1_M1022_g 0.0324226f $X=4.385 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B1_c_280_n N_C1_M1022_g 0.0110126f $X=4.13 $Y=2.015 $X2=0 $Y2=0
cc_248 N_B1_c_263_n N_C1_M1022_g 0.00432908f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_249 N_B1_c_280_n N_C1_c_348_n 0.0318234f $X=4.13 $Y=2.015 $X2=0 $Y2=0
cc_250 N_B1_c_263_n N_C1_c_348_n 0.023426f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_251 N_B1_c_264_n N_C1_c_348_n 9.3672e-19 $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_252 N_B1_c_266_n N_C1_c_348_n 0.0294252f $X=3.275 $Y=1.752 $X2=0 $Y2=0
cc_253 N_B1_c_280_n N_C1_c_349_n 0.0021094f $X=4.13 $Y=2.015 $X2=0 $Y2=0
cc_254 N_B1_c_263_n N_C1_c_349_n 8.05589e-19 $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_255 N_B1_c_264_n N_C1_c_349_n 0.021349f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_256 N_B1_c_265_n N_C1_c_349_n 0.016404f $X=2.795 $Y=1.51 $X2=0 $Y2=0
cc_257 N_B1_c_266_n N_C1_c_349_n 0.0147615f $X=3.275 $Y=1.752 $X2=0 $Y2=0
cc_258 N_B1_c_280_n N_A1_M1000_g 0.00102491f $X=4.13 $Y=2.015 $X2=0 $Y2=0
cc_259 N_B1_c_263_n N_A1_M1000_g 0.002453f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_260 N_B1_c_264_n N_A1_M1000_g 0.051097f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_261 N_B1_M1008_g N_A1_c_398_n 9.07148e-19 $X=4.275 $Y=0.665 $X2=0 $Y2=0
cc_262 N_B1_c_263_n N_A1_c_398_n 0.0114561f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_263 N_B1_c_264_n N_A1_c_398_n 6.2784e-19 $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_264 N_B1_c_263_n N_A1_c_399_n 2.27356e-19 $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_265 N_B1_c_264_n N_A1_c_399_n 0.0113225f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_266 N_B1_M1008_g N_A1_c_400_n 0.0179325f $X=4.275 $Y=0.665 $X2=0 $Y2=0
cc_267 N_B1_c_280_n N_VPWR_M1010_d 0.00333608f $X=4.13 $Y=2.015 $X2=0 $Y2=0
cc_268 N_B1_M1005_g N_VPWR_c_521_n 0.0126883f $X=2.585 $Y=2.465 $X2=0 $Y2=0
cc_269 N_B1_M1017_g N_VPWR_c_522_n 5.38417e-19 $X=4.385 $Y=2.465 $X2=0 $Y2=0
cc_270 N_B1_M1017_g N_VPWR_c_523_n 0.00244436f $X=4.385 $Y=2.465 $X2=0 $Y2=0
cc_271 N_B1_M1005_g N_VPWR_c_531_n 0.00486043f $X=2.585 $Y=2.465 $X2=0 $Y2=0
cc_272 N_B1_M1017_g N_VPWR_c_532_n 0.00585385f $X=4.385 $Y=2.465 $X2=0 $Y2=0
cc_273 N_B1_M1005_g N_VPWR_c_518_n 0.00896275f $X=2.585 $Y=2.465 $X2=0 $Y2=0
cc_274 N_B1_M1017_g N_VPWR_c_518_n 0.0110254f $X=4.385 $Y=2.465 $X2=0 $Y2=0
cc_275 N_B1_M1004_g N_VGND_c_685_n 0.00406825f $X=2.795 $Y=0.665 $X2=0 $Y2=0
cc_276 N_B1_M1004_g N_VGND_c_693_n 0.00405838f $X=2.795 $Y=0.665 $X2=0 $Y2=0
cc_277 N_B1_M1008_g N_VGND_c_693_n 0.00405838f $X=4.275 $Y=0.665 $X2=0 $Y2=0
cc_278 N_B1_M1004_g N_VGND_c_695_n 0.00713027f $X=2.795 $Y=0.665 $X2=0 $Y2=0
cc_279 N_B1_M1008_g N_VGND_c_695_n 0.00593651f $X=4.275 $Y=0.665 $X2=0 $Y2=0
cc_280 N_B1_M1004_g N_A_475_49#_c_787_n 0.0136763f $X=2.795 $Y=0.665 $X2=0 $Y2=0
cc_281 N_B1_M1008_g N_A_475_49#_c_787_n 0.0116825f $X=4.275 $Y=0.665 $X2=0 $Y2=0
cc_282 N_B1_c_263_n N_A_475_49#_c_787_n 0.00595536f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_283 N_B1_c_263_n N_A_475_49#_c_793_n 0.00385354f $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_284 N_B1_c_264_n N_A_475_49#_c_793_n 5.10915e-19 $X=4.295 $Y=1.51 $X2=0 $Y2=0
cc_285 N_B1_M1004_g N_A_574_49#_c_849_n 0.00281111f $X=2.795 $Y=0.665 $X2=0
+ $Y2=0
cc_286 N_B1_M1008_g N_A_574_49#_c_849_n 0.00265785f $X=4.275 $Y=0.665 $X2=0
+ $Y2=0
cc_287 N_C1_M1010_g N_VPWR_c_522_n 0.0122298f $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_288 N_C1_M1022_g N_VPWR_c_522_n 0.0109317f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_289 N_C1_M1010_g N_VPWR_c_531_n 0.00486043f $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_290 N_C1_M1022_g N_VPWR_c_532_n 0.00486043f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_291 N_C1_M1010_g N_VPWR_c_518_n 0.00896275f $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_292 N_C1_M1022_g N_VPWR_c_518_n 0.00864313f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_293 N_C1_M1016_g N_VGND_c_693_n 0.00351226f $X=3.225 $Y=0.665 $X2=0 $Y2=0
cc_294 N_C1_M1020_g N_VGND_c_693_n 0.00351226f $X=3.845 $Y=0.665 $X2=0 $Y2=0
cc_295 N_C1_M1016_g N_VGND_c_695_n 0.00574421f $X=3.225 $Y=0.665 $X2=0 $Y2=0
cc_296 N_C1_M1020_g N_VGND_c_695_n 0.00574421f $X=3.845 $Y=0.665 $X2=0 $Y2=0
cc_297 N_C1_M1016_g N_A_475_49#_c_787_n 0.0118636f $X=3.225 $Y=0.665 $X2=0 $Y2=0
cc_298 N_C1_M1020_g N_A_475_49#_c_787_n 0.0133795f $X=3.845 $Y=0.665 $X2=0 $Y2=0
cc_299 N_C1_c_348_n N_A_475_49#_c_787_n 0.00494446f $X=3.755 $Y=1.51 $X2=0 $Y2=0
cc_300 N_C1_M1016_g N_A_574_49#_c_849_n 0.0098454f $X=3.225 $Y=0.665 $X2=0 $Y2=0
cc_301 N_C1_M1020_g N_A_574_49#_c_849_n 0.0098454f $X=3.845 $Y=0.665 $X2=0 $Y2=0
cc_302 N_A1_c_397_n N_A2_M1006_g 0.0105246f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_303 N_A1_c_398_n N_A2_M1006_g 0.00121025f $X=4.835 $Y=1.17 $X2=0 $Y2=0
cc_304 N_A1_c_399_n N_A2_M1006_g 0.0209616f $X=4.835 $Y=1.36 $X2=0 $Y2=0
cc_305 N_A1_c_400_n N_A2_M1006_g 0.025367f $X=4.835 $Y=1.195 $X2=0 $Y2=0
cc_306 N_A1_c_395_n N_A2_M1018_g 0.0251472f $X=6.145 $Y=1.195 $X2=0 $Y2=0
cc_307 N_A1_c_397_n N_A2_M1018_g 0.010445f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_308 A1 N_A2_M1018_g 7.21709e-19 $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_309 N_A1_M1019_g N_A2_M1013_g 0.0251472f $X=6.145 $Y=2.465 $X2=0 $Y2=0
cc_310 N_A1_M1000_g A2 0.00144725f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A1_M1019_g A2 0.00960015f $X=6.145 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A1_c_397_n A2 0.0701088f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_313 N_A1_c_398_n A2 0.00669589f $X=4.835 $Y=1.17 $X2=0 $Y2=0
cc_314 N_A1_c_401_n A2 0.00437034f $X=6.45 $Y=1.36 $X2=0 $Y2=0
cc_315 A1 A2 0.0274319f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_316 N_A1_M1000_g N_A2_c_468_n 0.0603109f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A1_c_397_n N_A2_c_468_n 0.00246472f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_318 N_A1_c_401_n N_A2_c_468_n 0.0251472f $X=6.45 $Y=1.36 $X2=0 $Y2=0
cc_319 N_A1_M1000_g N_VPWR_c_523_n 0.00355731f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A1_M1019_g N_VPWR_c_525_n 0.021641f $X=6.145 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A1_c_397_n N_VPWR_c_525_n 0.00216799f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_322 N_A1_c_401_n N_VPWR_c_525_n 0.00275697f $X=6.45 $Y=1.36 $X2=0 $Y2=0
cc_323 A1 N_VPWR_c_525_n 0.0191794f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_324 N_A1_M1000_g N_VPWR_c_533_n 0.00547467f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_325 N_A1_M1019_g N_VPWR_c_533_n 0.00486043f $X=6.145 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A1_M1000_g N_VPWR_c_518_n 0.0100622f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A1_M1019_g N_VPWR_c_518_n 0.0082726f $X=6.145 $Y=2.465 $X2=0 $Y2=0
cc_328 N_A1_M1000_g N_A_986_367#_c_670_n 0.00369163f $X=4.855 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_A1_c_398_n N_VGND_M1001_d 0.00186101f $X=4.835 $Y=1.17 $X2=0 $Y2=0
cc_330 N_A1_c_400_n N_VGND_c_686_n 0.00321818f $X=4.835 $Y=1.195 $X2=0 $Y2=0
cc_331 N_A1_c_395_n N_VGND_c_687_n 0.00271672f $X=6.145 $Y=1.195 $X2=0 $Y2=0
cc_332 N_A1_c_400_n N_VGND_c_693_n 0.00431866f $X=4.835 $Y=1.195 $X2=0 $Y2=0
cc_333 N_A1_c_395_n N_VGND_c_694_n 0.00419886f $X=6.145 $Y=1.195 $X2=0 $Y2=0
cc_334 N_A1_c_395_n N_VGND_c_695_n 0.00689946f $X=6.145 $Y=1.195 $X2=0 $Y2=0
cc_335 N_A1_c_400_n N_VGND_c_695_n 0.00631324f $X=4.835 $Y=1.195 $X2=0 $Y2=0
cc_336 N_A1_c_402_n N_A_475_49#_M1003_s 0.00186977f $X=6.475 $Y=1.255 $X2=0
+ $Y2=0
cc_337 N_A1_c_397_n N_A_475_49#_c_799_n 0.0218641f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_338 N_A1_c_398_n N_A_475_49#_c_799_n 0.0190828f $X=4.835 $Y=1.17 $X2=0 $Y2=0
cc_339 N_A1_c_399_n N_A_475_49#_c_799_n 8.14813e-19 $X=4.835 $Y=1.36 $X2=0 $Y2=0
cc_340 N_A1_c_400_n N_A_475_49#_c_799_n 0.0113869f $X=4.835 $Y=1.195 $X2=0 $Y2=0
cc_341 N_A1_c_395_n N_A_475_49#_c_803_n 5.25381e-19 $X=6.145 $Y=1.195 $X2=0
+ $Y2=0
cc_342 N_A1_c_400_n N_A_475_49#_c_803_n 4.56293e-19 $X=4.835 $Y=1.195 $X2=0
+ $Y2=0
cc_343 N_A1_c_395_n N_A_475_49#_c_782_n 0.00953162f $X=6.145 $Y=1.195 $X2=0
+ $Y2=0
cc_344 N_A1_c_397_n N_A_475_49#_c_782_n 0.0405578f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_345 N_A1_c_401_n N_A_475_49#_c_782_n 0.00169797f $X=6.45 $Y=1.36 $X2=0 $Y2=0
cc_346 N_A1_c_402_n N_A_475_49#_c_782_n 0.0190225f $X=6.475 $Y=1.255 $X2=0 $Y2=0
cc_347 N_A1_c_395_n N_A_475_49#_c_783_n 0.00637396f $X=6.145 $Y=1.195 $X2=0
+ $Y2=0
cc_348 N_A1_c_397_n N_A_475_49#_c_810_n 0.0217194f $X=6.315 $Y=1.17 $X2=0 $Y2=0
cc_349 N_A2_M1013_g N_VPWR_c_525_n 0.00109252f $X=5.715 $Y=2.465 $X2=0 $Y2=0
cc_350 N_A2_M1007_g N_VPWR_c_533_n 0.00357877f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_351 N_A2_M1013_g N_VPWR_c_533_n 0.00357877f $X=5.715 $Y=2.465 $X2=0 $Y2=0
cc_352 N_A2_M1007_g N_VPWR_c_518_n 0.00544922f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_353 N_A2_M1013_g N_VPWR_c_518_n 0.00537654f $X=5.715 $Y=2.465 $X2=0 $Y2=0
cc_354 N_A2_M1007_g N_A_986_367#_c_670_n 0.0117007f $X=5.285 $Y=2.465 $X2=0
+ $Y2=0
cc_355 N_A2_M1013_g N_A_986_367#_c_670_n 0.0150885f $X=5.715 $Y=2.465 $X2=0
+ $Y2=0
cc_356 A2 N_A_986_367#_c_675_n 0.0153284f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_357 N_A2_M1006_g N_VGND_c_686_n 0.0036092f $X=5.285 $Y=0.665 $X2=0 $Y2=0
cc_358 N_A2_M1018_g N_VGND_c_687_n 0.00149374f $X=5.715 $Y=0.665 $X2=0 $Y2=0
cc_359 N_A2_M1006_g N_VGND_c_690_n 0.00419886f $X=5.285 $Y=0.665 $X2=0 $Y2=0
cc_360 N_A2_M1018_g N_VGND_c_690_n 0.00419886f $X=5.715 $Y=0.665 $X2=0 $Y2=0
cc_361 N_A2_M1006_g N_VGND_c_695_n 0.00614215f $X=5.285 $Y=0.665 $X2=0 $Y2=0
cc_362 N_A2_M1018_g N_VGND_c_695_n 0.00588507f $X=5.715 $Y=0.665 $X2=0 $Y2=0
cc_363 N_A2_M1006_g N_A_475_49#_c_799_n 0.00938107f $X=5.285 $Y=0.665 $X2=0
+ $Y2=0
cc_364 N_A2_M1006_g N_A_475_49#_c_803_n 0.00689232f $X=5.285 $Y=0.665 $X2=0
+ $Y2=0
cc_365 N_A2_M1018_g N_A_475_49#_c_803_n 0.00637396f $X=5.715 $Y=0.665 $X2=0
+ $Y2=0
cc_366 N_A2_M1018_g N_A_475_49#_c_782_n 0.00881445f $X=5.715 $Y=0.665 $X2=0
+ $Y2=0
cc_367 N_A2_M1018_g N_A_475_49#_c_783_n 5.25381e-19 $X=5.715 $Y=0.665 $X2=0
+ $Y2=0
cc_368 N_A2_M1006_g N_A_475_49#_c_810_n 7.17169e-19 $X=5.285 $Y=0.665 $X2=0
+ $Y2=0
cc_369 N_A2_M1018_g N_A_475_49#_c_810_n 7.17169e-19 $X=5.715 $Y=0.665 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_518_n N_X_M1002_s 0.00571434f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_371 N_VPWR_c_518_n N_X_M1012_s 0.00536646f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_372 N_VPWR_M1002_d N_X_c_619_n 0.00262981f $X=0.525 $Y=1.835 $X2=0 $Y2=0
cc_373 N_VPWR_c_519_n N_X_c_619_n 0.0220026f $X=0.65 $Y=2.18 $X2=0 $Y2=0
cc_374 N_VPWR_c_526_n N_X_c_652_n 0.0120977f $X=1.345 $Y=3.33 $X2=0 $Y2=0
cc_375 N_VPWR_c_518_n N_X_c_652_n 0.00691495f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_M1009_d N_X_c_621_n 0.00176461f $X=1.37 $Y=1.835 $X2=0 $Y2=0
cc_377 N_VPWR_c_520_n N_X_c_621_n 0.0170777f $X=1.51 $Y=2.18 $X2=0 $Y2=0
cc_378 N_VPWR_c_528_n N_X_c_656_n 0.0124525f $X=2.205 $Y=3.33 $X2=0 $Y2=0
cc_379 N_VPWR_c_518_n N_X_c_656_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_c_518_n N_A_986_367#_M1000_d 0.00225186f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_381 N_VPWR_c_518_n N_A_986_367#_M1013_d 0.00376627f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_533_n N_A_986_367#_c_670_n 0.0521332f $X=6.195 $Y=3.33 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_518_n N_A_986_367#_c_670_n 0.0338183f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_533_n N_A_986_367#_c_680_n 0.0125234f $X=6.195 $Y=3.33 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_518_n N_A_986_367#_c_680_n 0.0073762f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_386 N_X_c_617_n N_VGND_M1011_s 0.00244292f $X=0.227 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_387 N_X_c_615_n N_VGND_M1014_s 0.00176461f $X=1.455 $Y=1.13 $X2=0 $Y2=0
cc_388 N_X_c_614_n N_VGND_c_683_n 0.00178608f $X=0.595 $Y=1.13 $X2=0 $Y2=0
cc_389 N_X_c_617_n N_VGND_c_683_n 0.0224079f $X=0.227 $Y=1.215 $X2=0 $Y2=0
cc_390 N_X_c_615_n N_VGND_c_684_n 0.0170777f $X=1.455 $Y=1.13 $X2=0 $Y2=0
cc_391 N_X_c_663_p N_VGND_c_688_n 0.0128073f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_392 N_X_c_664_p N_VGND_c_692_n 0.0124525f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_393 N_X_M1011_d N_VGND_c_695_n 0.00536646f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_394 N_X_M1015_d N_VGND_c_695_n 0.00501859f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_395 N_X_c_664_p N_VGND_c_695_n 0.00730901f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_396 N_X_c_663_p N_VGND_c_695_n 0.00769778f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_397 N_VGND_c_695_n N_A_475_49#_M1004_d 0.00296364f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_398 N_VGND_c_695_n N_A_475_49#_M1008_d 0.00266641f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_399 N_VGND_c_695_n N_A_475_49#_M1006_d 0.00223559f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_695_n N_A_475_49#_M1003_s 0.00212301f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_685_n N_A_475_49#_c_780_n 0.0164094f $X=1.98 $Y=0.38 $X2=0 $Y2=0
cc_402 N_VGND_c_685_n N_A_475_49#_c_781_n 0.0229633f $X=1.98 $Y=0.38 $X2=0 $Y2=0
cc_403 N_VGND_c_693_n N_A_475_49#_c_781_n 0.0229787f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_404 N_VGND_c_695_n N_A_475_49#_c_781_n 0.0127264f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_405 N_VGND_c_693_n N_A_475_49#_c_787_n 0.00476763f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_406 N_VGND_c_695_n N_A_475_49#_c_787_n 0.0104194f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_407 N_VGND_c_693_n N_A_475_49#_c_828_n 0.0166842f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_695_n N_A_475_49#_c_828_n 0.0104192f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_M1001_d N_A_475_49#_c_799_n 0.00584819f $X=4.82 $Y=0.245 $X2=0
+ $Y2=0
cc_410 N_VGND_c_686_n N_A_475_49#_c_799_n 0.0216986f $X=5 $Y=0.44 $X2=0 $Y2=0
cc_411 N_VGND_c_690_n N_A_475_49#_c_799_n 0.00191958f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_693_n N_A_475_49#_c_799_n 0.00205543f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_695_n N_A_475_49#_c_799_n 0.0086621f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_690_n N_A_475_49#_c_803_n 0.0188913f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_695_n N_A_475_49#_c_803_n 0.012376f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_M1018_s N_A_475_49#_c_782_n 0.00349386f $X=5.79 $Y=0.245 $X2=0
+ $Y2=0
cc_417 N_VGND_c_687_n N_A_475_49#_c_782_n 0.0130506f $X=5.93 $Y=0.41 $X2=0 $Y2=0
cc_418 N_VGND_c_690_n N_A_475_49#_c_782_n 0.00191958f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_c_694_n N_A_475_49#_c_782_n 0.00191958f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_695_n N_A_475_49#_c_782_n 0.00827851f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_694_n N_A_475_49#_c_783_n 0.0210049f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_695_n N_A_475_49#_c_783_n 0.0125589f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_695_n N_A_475_49#_c_793_n 8.87777e-19 $X=6.48 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_695_n N_A_574_49#_M1004_s 0.00223577f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_425 N_VGND_c_695_n N_A_574_49#_M1020_s 0.00223577f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_693_n N_A_574_49#_c_849_n 0.0780173f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_695_n N_A_574_49#_c_849_n 0.0502425f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_428 N_A_475_49#_c_787_n N_A_574_49#_M1004_s 0.00384083f $X=4.365 $Y=0.72
+ $X2=-0.19 $Y2=-0.245
cc_429 N_A_475_49#_c_787_n N_A_574_49#_M1020_s 0.00776805f $X=4.365 $Y=0.72
+ $X2=0 $Y2=0
cc_430 N_A_475_49#_c_787_n N_A_574_49#_c_849_n 0.0709297f $X=4.365 $Y=0.72 $X2=0
+ $Y2=0
