* File: sky130_fd_sc_lp__clkinv_1.pxi.spice
* Created: Fri Aug 28 10:17:44 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINV_1%A N_A_M1000_g N_A_M1001_g N_A_c_27_n N_A_M1002_g
+ A A A PM_SKY130_FD_SC_LP__CLKINV_1%A
x_PM_SKY130_FD_SC_LP__CLKINV_1%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_c_57_n
+ N_VPWR_c_58_n N_VPWR_c_59_n N_VPWR_c_60_n VPWR N_VPWR_c_61_n N_VPWR_c_56_n
+ PM_SKY130_FD_SC_LP__CLKINV_1%VPWR
x_PM_SKY130_FD_SC_LP__CLKINV_1%Y N_Y_M1001_s N_Y_M1000_s N_Y_c_77_n N_Y_c_81_n Y
+ Y Y PM_SKY130_FD_SC_LP__CLKINV_1%Y
x_PM_SKY130_FD_SC_LP__CLKINV_1%VGND N_VGND_M1001_d N_VGND_c_101_n N_VGND_c_102_n
+ VGND N_VGND_c_103_n N_VGND_c_104_n PM_SKY130_FD_SC_LP__CLKINV_1%VGND
cc_1 VNB N_A_M1001_g 0.0417082f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.56
cc_2 VNB N_A_c_27_n 0.102616f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.6
cc_3 VNB N_A_M1002_g 0.00312369f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.53
cc_4 VNB A 0.0438986f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_VPWR_c_56_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.27
cc_6 VNB N_Y_c_77_n 0.00194427f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.6
cc_7 VNB Y 0.019474f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB Y 0.0178819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB Y 0.00353325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_101_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_102_n 0.0228715f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.56
cc_12 VNB N_VGND_c_103_n 0.0327369f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.53
cc_13 VNB N_VGND_c_104_n 0.122328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VPB N_A_M1000_g 0.038271f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.53
cc_15 VPB N_A_c_27_n 0.0173042f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.6
cc_16 VPB N_A_M1002_g 0.0419935f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.53
cc_17 VPB A 0.0114762f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_18 VPB N_VPWR_c_57_n 0.0131663f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.56
cc_19 VPB N_VPWR_c_58_n 0.0400344f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.6
cc_20 VPB N_VPWR_c_59_n 0.0109759f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.53
cc_21 VPB N_VPWR_c_60_n 0.0437164f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_22 VPB N_VPWR_c_61_n 0.016185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_56_n 0.0546942f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.27
cc_24 VPB N_Y_c_81_n 0.00688915f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_25 VPB Y 0.0162053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 N_A_M1000_g N_VPWR_c_58_n 0.0133851f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_27 N_A_c_27_n N_VPWR_c_58_n 0.00138689f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_28 N_A_M1002_g N_VPWR_c_58_n 5.4051e-19 $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_29 A N_VPWR_c_58_n 0.0149329f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_30 N_A_M1002_g N_VPWR_c_60_n 0.00458933f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_31 N_A_M1000_g N_VPWR_c_61_n 0.00512473f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_32 N_A_M1002_g N_VPWR_c_61_n 0.00570944f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_33 N_A_M1000_g N_VPWR_c_56_n 0.00492022f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_34 N_A_M1002_g N_VPWR_c_56_n 0.00542671f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_35 N_A_M1001_g N_Y_c_77_n 0.00304928f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_36 A N_Y_c_77_n 0.0835948f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_37 N_A_M1000_g N_Y_c_81_n 0.00545505f $X=0.535 $Y=2.53 $X2=0 $Y2=0
cc_38 N_A_M1002_g N_Y_c_81_n 0.00606174f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_39 N_A_M1001_g Y 0.0176135f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_40 N_A_c_27_n Y 0.009494f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_41 N_A_c_27_n Y 0.0295942f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_42 N_A_c_27_n Y 0.00935938f $X=0.965 $Y=1.6 $X2=0 $Y2=0
cc_43 N_A_M1002_g Y 0.0205729f $X=0.965 $Y=2.53 $X2=0 $Y2=0
cc_44 N_A_M1001_g N_VGND_c_102_n 0.013725f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_45 N_A_M1001_g N_VGND_c_103_n 0.00396895f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_46 N_A_M1001_g N_VGND_c_104_n 0.00422451f $X=0.965 $Y=0.56 $X2=0 $Y2=0
cc_47 A N_VGND_c_104_n 0.0151652f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_48 N_VPWR_c_58_n N_Y_c_81_n 0.0302518f $X=0.32 $Y=2.345 $X2=0 $Y2=0
cc_49 N_VPWR_c_60_n N_Y_c_81_n 0.00152757f $X=1.18 $Y=2.345 $X2=0 $Y2=0
cc_50 N_VPWR_c_61_n N_Y_c_81_n 0.00978084f $X=1.045 $Y=3.33 $X2=0 $Y2=0
cc_51 N_VPWR_c_56_n N_Y_c_81_n 0.00836996f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_52 N_VPWR_c_60_n Y 0.0136765f $X=1.18 $Y=2.345 $X2=0 $Y2=0
cc_53 Y N_VGND_c_102_n 0.0212507f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_54 N_Y_c_77_n N_VGND_c_103_n 0.00706712f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_55 N_Y_c_77_n N_VGND_c_104_n 0.00711097f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_56 Y N_VGND_c_104_n 0.00673873f $X=1.115 $Y=0.84 $X2=0 $Y2=0
