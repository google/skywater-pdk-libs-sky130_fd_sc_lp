* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__invlp_4 A VGND VNB VPB VPWR Y
X0 a_118_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_118_367# A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR A a_118_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_114_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_114_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Y A a_118_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_114_53# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 Y A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_118_367# A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR A a_118_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y A a_118_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 Y A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_114_53# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_118_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
