* File: sky130_fd_sc_lp__or2_lp2.pex.spice
* Created: Wed Sep  2 10:29:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2_LP2%B 2 5 7 8 11 13 15 16 18 19 20 21 22 39
r45 39 41 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.78 $Y=1.345
+ $X2=0.78 $Y2=1.18
r46 21 22 5.4975 $w=8.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.527 $Y=2.405
+ $X2=0.527 $Y2=2.775
r47 20 21 5.4975 $w=8.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.527 $Y=2.035
+ $X2=0.527 $Y2=2.405
r48 19 20 5.4975 $w=8.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.527 $Y=1.665
+ $X2=0.527 $Y2=2.035
r49 18 19 5.4975 $w=8.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.527 $Y=1.295
+ $X2=0.527 $Y2=1.665
r50 18 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.765
+ $Y=1.345 $X2=0.765 $Y2=1.345
r51 13 16 69.4185 $w=1.84e-07 $l=2.65e-07 $layer=POLY_cond $X=1.54 $Y=1.837
+ $X2=1.275 $Y2=1.837
r52 13 15 109.896 $w=2.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.54 $Y=1.975
+ $X2=1.54 $Y2=2.545
r53 9 16 7.64856 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=1.275 $Y=1.7
+ $X2=1.275 $Y2=1.837
r54 9 11 617.883 $w=1.5e-07 $l=1.205e-06 $layer=POLY_cond $X=1.275 $Y=1.7
+ $X2=1.275 $Y2=0.495
r55 7 16 21.4346 $w=1.84e-07 $l=1.01366e-07 $layer=POLY_cond $X=1.2 $Y=1.775
+ $X2=1.275 $Y2=1.837
r56 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.2 $Y=1.775 $X2=0.96
+ $Y2=1.775
r57 5 41 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.885 $Y=0.495
+ $X2=0.885 $Y2=1.18
r58 2 8 33.3473 $w=1.5e-07 $l=2.14243e-07 $layer=POLY_cond $X=0.78 $Y=1.7
+ $X2=0.96 $Y2=1.775
r59 1 39 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=0.78 $Y=1.36 $X2=0.78
+ $Y2=1.345
r60 1 2 54.4984 $w=3.6e-07 $l=3.4e-07 $layer=POLY_cond $X=0.78 $Y=1.36 $X2=0.78
+ $Y2=1.7
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP2%A 3 7 11 17 19 20 23 24
c44 17 0 1.56547e-19 $X=2.065 $Y=0.98
r45 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.975
+ $Y=1.07 $X2=1.975 $Y2=1.07
r46 20 24 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.68 $Y=1.24
+ $X2=1.975 $Y2=1.24
r47 19 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.975 $Y=1.41
+ $X2=1.975 $Y2=1.07
r48 16 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.975 $Y=1.055
+ $X2=1.975 $Y2=1.07
r49 16 17 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.975 $Y=0.98
+ $X2=2.065 $Y2=0.98
r50 13 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.705 $Y=0.98
+ $X2=1.975 $Y2=0.98
r51 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.065 $Y=0.905
+ $X2=2.065 $Y2=0.98
r52 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.065 $Y=0.905
+ $X2=2.065 $Y2=0.495
r53 5 19 47.383 $w=2.95e-07 $l=3.16307e-07 $layer=POLY_cond $X=2.03 $Y=1.7
+ $X2=1.975 $Y2=1.41
r54 5 7 209.943 $w=2.5e-07 $l=8.45e-07 $layer=POLY_cond $X=2.03 $Y=1.7 $X2=2.03
+ $Y2=2.545
r55 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.705 $Y=0.905
+ $X2=1.705 $Y2=0.98
r56 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.705 $Y=0.905
+ $X2=1.705 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP2%A_226_409# 1 2 9 13 17 20 23 27 31 32 37 39
c71 32 0 1.60417e-19 $X=2.56 $Y=1.38
c72 20 0 1.56547e-19 $X=1.195 $Y=1.755
r73 34 37 7.6705 $w=4.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.195 $Y=0.495
+ $X2=1.49 $Y2=0.495
r74 32 41 65.7961 $w=5.35e-07 $l=5.05e-07 $layer=POLY_cond $X=2.662 $Y=1.38
+ $X2=2.662 $Y2=1.885
r75 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.56
+ $Y=1.38 $X2=2.56 $Y2=1.38
r76 29 31 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.56 $Y=1.755
+ $X2=2.56 $Y2=1.38
r77 28 39 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.44 $Y=1.84
+ $X2=1.275 $Y2=1.84
r78 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.395 $Y=1.84
+ $X2=2.56 $Y2=1.755
r79 27 28 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.395 $Y=1.84
+ $X2=1.44 $Y2=1.84
r80 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.275 $Y=2.19
+ $X2=1.275 $Y2=2.9
r81 21 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=1.925
+ $X2=1.275 $Y2=1.84
r82 21 23 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.275 $Y=1.925
+ $X2=1.275 $Y2=2.19
r83 20 39 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.195 $Y=1.755
+ $X2=1.275 $Y2=1.84
r84 19 34 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.195 $Y=0.725
+ $X2=1.195 $Y2=0.495
r85 19 20 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=1.195 $Y=0.725
+ $X2=1.195 $Y2=1.755
r86 15 32 31.8222 $w=2.67e-07 $l=2.62857e-07 $layer=POLY_cond $X=2.855 $Y=1.215
+ $X2=2.662 $Y2=1.38
r87 15 17 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.855 $Y=1.215
+ $X2=2.855 $Y2=0.495
r88 13 41 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.805 $Y=2.545
+ $X2=2.805 $Y2=1.885
r89 7 32 31.8222 $w=2.67e-07 $l=2.35465e-07 $layer=POLY_cond $X=2.495 $Y=1.215
+ $X2=2.662 $Y2=1.38
r90 7 9 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.495 $Y=1.215
+ $X2=2.495 $Y2=0.495
r91 2 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=2.045 $X2=1.275 $Y2=2.9
r92 2 23 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=2.045 $X2=1.275 $Y2=2.19
r93 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.35
+ $Y=0.285 $X2=1.49 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP2%VPWR 1 6 8 10 17 18 21
r24 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r25 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=3.33
+ $X2=2.295 $Y2=3.33
r28 15 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.46 $Y=3.33
+ $X2=3.12 $Y2=3.33
r29 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.13 $Y=3.33
+ $X2=2.295 $Y2=3.33
r31 10 12 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=2.13 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=3.245
+ $X2=2.295 $Y2=3.33
r35 4 6 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=2.295 $Y=3.245
+ $X2=2.295 $Y2=2.27
r36 1 6 300 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=2 $X=2.155
+ $Y=2.045 $X2=2.295 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP2%X 1 2 7 8 9 10 11 12 13
r14 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.07 $Y=2.775
+ $X2=3.07 $Y2=2.9
r15 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.07 $Y=2.405
+ $X2=3.07 $Y2=2.775
r16 12 34 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.07 $Y=2.405
+ $X2=3.07 $Y2=2.19
r17 11 34 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.07 $Y=2.035
+ $X2=3.07 $Y2=2.19
r18 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.07 $Y=1.665
+ $X2=3.07 $Y2=2.035
r19 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.07 $Y=1.295
+ $X2=3.07 $Y2=1.665
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.07 $Y=0.925 $X2=3.07
+ $Y2=1.295
r21 7 8 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.07 $Y=0.495 $X2=3.07
+ $Y2=0.925
r22 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=2.045 $X2=3.07 $Y2=2.9
r23 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=2.045 $X2=3.07 $Y2=2.19
r24 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.285 $X2=3.07 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP2%VGND 1 2 9 13 15 17 22 29 30 33 36
c37 13 0 1.60417e-19 $X=2.28 $Y=0.495
r38 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r41 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r43 27 29 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=3.12
+ $Y2=0
r44 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r45 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=0 $X2=0.67
+ $Y2=0
r47 23 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.835 $Y=0 $X2=1.2
+ $Y2=0
r48 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r49 22 25 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.2
+ $Y2=0
r50 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r51 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.505 $Y=0 $X2=0.67
+ $Y2=0
r53 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.505 $Y=0 $X2=0.24
+ $Y2=0
r54 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r55 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r56 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r57 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.495
r58 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085 $X2=0.67
+ $Y2=0
r59 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.67 $Y=0.085 $X2=0.67
+ $Y2=0.495
r60 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.285 $X2=2.28 $Y2=0.495
r61 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.525
+ $Y=0.285 $X2=0.67 $Y2=0.495
.ends

