* File: sky130_fd_sc_lp__a21bo_0.pex.spice
* Created: Wed Sep  2 09:18:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BO_0%A_72_212# 1 2 9 13 17 18 21 22 24 25 28 31
+ 33 38
c86 31 0 1.43696e-19 $X=2.29 $Y=1.56
r87 35 38 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.47
+ $X2=2.375 $Y2=0.47
r88 31 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=1.56
+ $X2=2.29 $Y2=1.645
r89 30 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=0.635
+ $X2=2.29 $Y2=0.47
r90 30 31 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.29 $Y=0.635
+ $X2=2.29 $Y2=1.56
r91 26 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.025 $Y=1.645
+ $X2=2.29 $Y2=1.645
r92 26 28 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=2.025 $Y=1.73
+ $X2=2.025 $Y2=2.435
r93 24 26 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.88 $Y=1.645
+ $X2=2.025 $Y2=1.645
r94 24 25 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=1.88 $Y=1.645
+ $X2=0.695 $Y2=1.645
r95 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.225 $X2=0.525 $Y2=1.225
r96 19 25 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.562 $Y=1.56
+ $X2=0.695 $Y2=1.645
r97 19 21 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=0.562 $Y=1.56
+ $X2=0.562 $Y2=1.225
r98 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=1.225
r99 17 18 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=1.73
r100 16 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.06
+ $X2=0.525 $Y2=1.225
r101 13 16 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.615 $Y=0.47
+ $X2=0.615 $Y2=1.06
r102 9 18 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=0.48 $Y=2.73 $X2=0.48
+ $Y2=1.73
r103 2 28 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=2.29 $X2=2.045 $Y2=2.435
r104 1 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.26 $X2=2.375 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%B1_N 3 7 9 10 11 12 13 17
r45 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.095
+ $Y=0.955 $X2=1.095 $Y2=0.955
r46 13 18 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.13 $Y=1.295
+ $X2=1.13 $Y2=0.955
r47 12 18 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=1.13 $Y=0.925
+ $X2=1.13 $Y2=0.955
r48 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=0.955
r49 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=1.46
r50 9 17 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=0.79
+ $X2=1.095 $Y2=0.955
r51 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.045 $Y=0.47
+ $X2=1.045 $Y2=0.79
r52 3 11 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=1.005 $Y=2.84
+ $X2=1.005 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%A_216_526# 1 2 9 10 11 13 15 18 22 23 26 30
+ 32 43 44 47 48 49 52
c81 26 0 3.98952e-20 $X=2.26 $Y=1.825
r82 47 49 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.955
+ $X2=1.665 $Y2=0.87
r83 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.665
+ $Y=0.955 $X2=1.665 $Y2=0.955
r84 44 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.995
+ $X2=1.485 $Y2=1.83
r85 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.485
+ $Y=1.995 $X2=1.485 $Y2=1.995
r86 36 49 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.585 $Y=0.635
+ $X2=1.585 $Y2=0.87
r87 32 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.5 $Y=0.47
+ $X2=1.585 $Y2=0.635
r88 32 34 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.5 $Y=0.47 $X2=1.26
+ $Y2=0.47
r89 28 43 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=1.22 $Y=2.03
+ $X2=1.485 $Y2=2.03
r90 28 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.22 $Y=2.16
+ $X2=1.22 $Y2=2.84
r91 24 26 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.16 $Y=1.825 $X2=2.26
+ $Y2=1.825
r92 22 52 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.575 $Y=1.46
+ $X2=1.575 $Y2=1.83
r93 21 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.665 $Y=1.295
+ $X2=1.665 $Y2=0.955
r94 21 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.295
+ $X2=1.665 $Y2=1.46
r95 20 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.665 $Y=0.94
+ $X2=1.665 $Y2=0.955
r96 16 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.26 $Y=1.9 $X2=2.26
+ $Y2=1.825
r97 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.26 $Y=1.9 $X2=2.26
+ $Y2=2.61
r98 15 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=1.75
+ $X2=2.16 $Y2=1.825
r99 14 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=0.94
+ $X2=2.16 $Y2=0.865
r100 14 15 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.16 $Y=0.94
+ $X2=2.16 $Y2=1.75
r101 11 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=0.79
+ $X2=2.16 $Y2=0.865
r102 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.16 $Y=0.79
+ $X2=2.16 $Y2=0.47
r103 10 20 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.83 $Y=0.865
+ $X2=1.665 $Y2=0.94
r104 9 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.085 $Y=0.865
+ $X2=2.16 $Y2=0.865
r105 9 10 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=2.085 $Y=0.865
+ $X2=1.83 $Y2=0.865
r106 2 30 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=2.63 $X2=1.22 $Y2=2.84
r107 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.26 $X2=1.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%A1 3 7 11 12 13 14 15 20
c47 13 0 1.43888e-19 $X=2.64 $Y=0.925
c48 7 0 1.43696e-19 $X=2.69 $Y=2.61
c49 3 0 1.00548e-19 $X=2.59 $Y=0.47
r50 14 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.665
r51 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=0.925
+ $X2=2.67 $Y2=1.295
r52 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.64
+ $Y=1.005 $X2=2.64 $Y2=1.005
r53 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.64 $Y=1.345
+ $X2=2.64 $Y2=1.005
r54 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.345
+ $X2=2.64 $Y2=1.51
r55 10 20 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=0.84
+ $X2=2.64 $Y2=1.005
r56 7 12 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=2.69 $Y=2.61 $X2=2.69
+ $Y2=1.51
r57 3 10 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.59 $Y=0.47 $X2=2.59
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%A2 3 7 11 12 13 14 15 20
c32 13 0 1.00548e-19 $X=3.12 $Y=0.925
c33 3 0 1.03993e-19 $X=3.12 $Y=0.47
r34 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.21
+ $Y=1.005 $X2=3.21 $Y2=1.005
r35 14 15 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.17 $Y=1.295
+ $X2=3.17 $Y2=1.665
r36 14 21 8.15143 $w=4.08e-07 $l=2.9e-07 $layer=LI1_cond $X=3.17 $Y=1.295
+ $X2=3.17 $Y2=1.005
r37 13 21 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=3.17 $Y=0.925 $X2=3.17
+ $Y2=1.005
r38 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.21 $Y=1.345
+ $X2=3.21 $Y2=1.005
r39 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.345
+ $X2=3.21 $Y2=1.51
r40 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.84
+ $X2=3.21 $Y2=1.005
r41 7 12 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=3.12 $Y=2.61 $X2=3.12
+ $Y2=1.51
r42 3 10 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.12 $Y=0.47 $X2=3.12
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%X 1 2 11 13 14 15 35
r20 21 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.255 $Y=2.115
+ $X2=0.255 $Y2=2.035
r21 15 26 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.255 $Y=2.775
+ $X2=0.255 $Y2=2.555
r22 14 26 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.255 $Y=2.405
+ $X2=0.255 $Y2=2.555
r23 13 35 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=0.255 $Y=2.032
+ $X2=0.255 $Y2=2.035
r24 13 14 10.0577 $w=3.28e-07 $l=2.88e-07 $layer=LI1_cond $X=0.255 $Y=2.117
+ $X2=0.255 $Y2=2.405
r25 13 21 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=0.255 $Y=2.117
+ $X2=0.255 $Y2=2.115
r26 8 13 56.3167 $w=2.73e-07 $l=1.315e-06 $layer=LI1_cond $X=0.175 $Y=0.635
+ $X2=0.175 $Y2=1.95
r27 7 11 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.175 $Y=0.47
+ $X2=0.4 $Y2=0.47
r28 7 8 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.175 $Y=0.47
+ $X2=0.175 $Y2=0.635
r29 2 26 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=2.41 $X2=0.265 $Y2=2.555
r30 1 11 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.26 $X2=0.4 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%VPWR 1 2 9 13 16 17 18 20 33 34 37
r41 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 25 37 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.737 $Y2=3.33
r49 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 20 37 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.737 $Y2=3.33
r53 20 22 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 16 30 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 16 17 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.902 $Y2=3.33
r58 15 33 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 15 17 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.902 $Y2=3.33
r60 11 17 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.902 $Y=3.245
+ $X2=2.902 $Y2=3.33
r61 11 13 34.7907 $w=2.63e-07 $l=8e-07 $layer=LI1_cond $X=2.902 $Y=3.245
+ $X2=2.902 $Y2=2.445
r62 7 37 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=3.245
+ $X2=0.737 $Y2=3.33
r63 7 9 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.737 $Y=3.245
+ $X2=0.737 $Y2=2.565
r64 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.765
+ $Y=2.29 $X2=2.905 $Y2=2.445
r65 1 9 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=2.41 $X2=0.695 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%A_467_458# 1 2 9 11 12 15
r26 13 15 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=3.352 $Y=2.1
+ $X2=3.352 $Y2=2.435
r27 11 13 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=3.205 $Y=2.015
+ $X2=3.352 $Y2=2.1
r28 11 12 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.205 $Y=2.015
+ $X2=2.6 $Y2=2.015
r29 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.47 $Y=2.1
+ $X2=2.6 $Y2=2.015
r30 7 9 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.47 $Y=2.1 $X2=2.47
+ $Y2=2.435
r31 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.195
+ $Y=2.29 $X2=3.335 $Y2=2.435
r32 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.335
+ $Y=2.29 $X2=2.475 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_0%VGND 1 2 3 14 18 22 25 26 28 29 30 43 44 47
r42 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 41 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r45 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r47 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r48 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 35 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r50 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 32 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.83
+ $Y2=0
r52 32 34 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.68
+ $Y2=0
r53 30 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r54 30 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r55 28 40 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.12
+ $Y2=0
r56 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.335
+ $Y2=0
r57 27 43 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.6 $Y2=0
r58 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.335
+ $Y2=0
r59 25 34 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.68
+ $Y2=0
r60 25 26 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.937
+ $Y2=0
r61 24 37 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.16
+ $Y2=0
r62 24 26 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.937
+ $Y2=0
r63 20 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0
r64 20 22 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0.47
r65 16 26 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.937 $Y=0.085
+ $X2=1.937 $Y2=0
r66 16 18 21.8974 $w=1.93e-07 $l=3.85e-07 $layer=LI1_cond $X=1.937 $Y=0.085
+ $X2=1.937 $Y2=0.47
r67 12 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0
r68 12 14 17.7476 $w=2.48e-07 $l=3.85e-07 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0.47
r69 3 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.26 $X2=3.335 $Y2=0.47
r70 2 18 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.26 $X2=1.945 $Y2=0.47
r71 1 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.26 $X2=0.83 $Y2=0.47
.ends

