* File: sky130_fd_sc_lp__einvn_m.pex.spice
* Created: Wed Sep  2 09:52:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVN_M%TE_B 4 5 7 8 10 12 13 14 15 19
r44 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.495
+ $X2=0.485 $Y2=0.66
r45 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=0.495 $X2=0.485 $Y2=0.495
r46 15 20 7.62885 $w=3.53e-07 $l=2.35e-07 $layer=LI1_cond $X=0.72 $Y=0.507
+ $X2=0.485 $Y2=0.507
r47 14 20 7.95348 $w=3.53e-07 $l=2.45e-07 $layer=LI1_cond $X=0.24 $Y=0.507
+ $X2=0.485 $Y2=0.507
r48 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.085 $Y=2.565
+ $X2=1.085 $Y2=2.885
r49 9 13 5.30422 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=0.73 $Y=2.49
+ $X2=0.615 $Y2=2.49
r50 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.01 $Y=2.49
+ $X2=1.085 $Y2=2.565
r51 8 9 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.01 $Y=2.49 $X2=0.73
+ $Y2=2.49
r52 5 13 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=0.655 $Y=2.565
+ $X2=0.615 $Y2=2.49
r53 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.655 $Y=2.565
+ $X2=0.655 $Y2=2.885
r54 4 22 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.575 $Y=0.98
+ $X2=0.575 $Y2=0.66
r55 2 13 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=0.575 $Y=2.415
+ $X2=0.615 $Y2=2.49
r56 2 4 735.819 $w=1.5e-07 $l=1.435e-06 $layer=POLY_cond $X=0.575 $Y=2.415
+ $X2=0.575 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_M%A_47_154# 1 2 9 15 19 21 25 27 28
c44 9 0 1.41744e-19 $X=1.015 $Y=0.98
r45 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.025
+ $Y=1.7 $X2=1.025 $Y2=1.7
r46 22 25 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=1.62
+ $X2=0.36 $Y2=1.62
r47 21 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=1.62
+ $X2=1.025 $Y2=1.62
r48 21 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.94 $Y=1.62
+ $X2=0.525 $Y2=1.62
r49 17 25 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.36 $Y=1.705
+ $X2=0.36 $Y2=1.62
r50 17 19 38.9386 $w=3.28e-07 $l=1.115e-06 $layer=LI1_cond $X=0.36 $Y=1.705
+ $X2=0.36 $Y2=2.82
r51 13 25 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.36 $Y=1.535
+ $X2=0.36 $Y2=1.62
r52 13 15 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=0.36 $Y=1.535
+ $X2=0.36 $Y2=1.02
r53 12 28 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=1.535
+ $X2=1.025 $Y2=1.7
r54 9 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.015 $Y=0.98
+ $X2=1.015 $Y2=1.535
r55 2 19 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=2.675 $X2=0.44 $Y2=2.82
r56 1 15 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.77 $X2=0.36 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_M%A 4 7 11 12 13 14 17
c32 14 0 1.41744e-19 $X=1.68 $Y=0.555
c33 13 0 7.59044e-20 $X=1.46 $Y=2.565
r34 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=0.42
+ $X2=1.465 $Y2=0.585
r35 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=0.42 $X2=1.465 $Y2=0.42
r36 14 18 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=0.47
+ $X2=1.465 $Y2=0.47
r37 12 13 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.46 $Y=2.415
+ $X2=1.46 $Y2=2.565
r38 11 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=1.475 $Y=1.415
+ $X2=1.475 $Y2=2.415
r39 10 11 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.46 $Y=1.265
+ $X2=1.46 $Y2=1.415
r40 7 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.445 $Y=2.885
+ $X2=1.445 $Y2=2.565
r41 4 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.445 $Y=0.98
+ $X2=1.445 $Y2=1.265
r42 4 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.445 $Y=0.98
+ $X2=1.445 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_M%VPWR 1 8 10 14 15 18
c27 14 0 7.59044e-20 $X=1.68 $Y=3.33
r28 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r30 12 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.87 $Y2=3.33
r31 12 14 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.68 $Y2=3.33
r32 10 15 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r33 10 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 6 18 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245 $X2=0.87
+ $Y2=3.33
r35 6 8 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=2.95
r36 1 8 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=2.675 $X2=0.87 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_M%Z 1 2 7 8 9 10 11 18
r18 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=2.405
+ $X2=1.66 $Y2=2.775
r19 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=2.035
+ $X2=1.66 $Y2=2.405
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.665 $X2=1.66
+ $Y2=2.035
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.295 $X2=1.66
+ $Y2=1.665
r22 7 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.66 $Y=1.295
+ $X2=1.66 $Y2=1.02
r23 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=2.675 $X2=1.66 $Y2=2.82
r24 1 18 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.77 $X2=1.66 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_M%VGND 1 5 9 12 13 14 21 22
r32 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r33 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 14 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r35 14 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r36 12 17 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r37 12 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.07
+ $Y2=0
r38 11 21 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.68
+ $Y2=0
r39 11 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.07
+ $Y2=0
r40 7 9 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.8 $Y=1.02 $X2=1.07
+ $Y2=1.02
r41 5 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0.855 $X2=1.07
+ $Y2=1.02
r42 4 13 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r43 4 5 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0.855
r44 1 7 182 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.77 $X2=0.8 $Y2=1.02
.ends

