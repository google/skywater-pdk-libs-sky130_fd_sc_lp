* NGSPICE file created from sky130_fd_sc_lp__o2bb2ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR A1_N a_804_39# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.0509e+12p pd=2.911e+07u as=1.4112e+12p ps=1.232e+07u
M1001 a_1235_65# A2_N a_804_39# VNB nshort w=840000u l=150000u
+  ad=1.218e+12p pd=1.13e+07u as=4.704e+11p ps=4.48e+06u
M1002 Y a_804_39# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.4112e+12p pd=1.232e+07u as=0p ps=0u
M1003 a_1235_65# A1_N VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.4784e+12p ps=1.36e+07u
M1004 a_1235_65# A1_N VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B2 a_132_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.449e+12p ps=1.238e+07u
M1006 VPWR A1_N a_804_39# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_804_39# A2_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_804_39# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B1 a_132_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_35_65# B2 VGND VNB nshort w=840000u l=150000u
+  ad=1.7388e+12p pd=1.59e+07u as=0p ps=0u
M1011 a_35_65# a_804_39# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=5.544e+11p ps=4.68e+06u
M1012 VPWR B1 a_132_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_804_39# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_804_39# A2_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_35_65# B2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_804_39# A2_N a_1235_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_35_65# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1235_65# A2_N a_804_39# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 a_35_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_804_39# A2_N a_1235_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_132_367# B2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_804_39# A1_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_804_39# a_35_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A1_N a_1235_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_804_39# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_804_39# A1_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y a_804_39# a_35_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR A2_N a_804_39# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND B2 a_35_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND B2 a_35_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_35_65# a_804_39# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_132_367# B2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR A2_N a_804_39# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND B1 a_35_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND A1_N a_1235_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_132_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y B2 a_132_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_132_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_35_65# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

