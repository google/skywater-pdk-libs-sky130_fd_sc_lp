# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a32oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.995000 1.210000 5.715000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.265000 1.210000 8.005000 1.435000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.315000 1.210000 10.455000 1.435000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.210000 3.815000 1.435000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.210000 1.845000 1.435000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 1.605000 6.095000 1.875000 ;
        RECT 0.600000 1.875000 0.930000 2.735000 ;
        RECT 1.460000 1.875000 1.790000 2.735000 ;
        RECT 2.250000 0.765000 6.095000 1.040000 ;
        RECT 2.320000 1.875000 2.650000 2.735000 ;
        RECT 3.180000 1.875000 3.510000 2.735000 ;
        RECT 5.885000 1.040000 6.095000 1.605000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.100000  0.255000  0.360000 0.870000 ;
      RECT 0.100000  0.870000  2.080000 1.040000 ;
      RECT 0.170000  1.825000  0.430000 2.905000 ;
      RECT 0.170000  2.905000  3.980000 3.075000 ;
      RECT 0.530000  0.085000  0.860000 0.700000 ;
      RECT 1.030000  0.255000  1.220000 0.870000 ;
      RECT 1.100000  2.045000  1.290000 2.905000 ;
      RECT 1.390000  0.085000  1.720000 0.700000 ;
      RECT 1.890000  0.255000  3.870000 0.595000 ;
      RECT 1.890000  0.595000  2.080000 0.870000 ;
      RECT 1.960000  2.045000  2.150000 2.905000 ;
      RECT 2.820000  2.045000  3.010000 2.905000 ;
      RECT 3.680000  2.045000  7.260000 2.225000 ;
      RECT 3.680000  2.225000  3.980000 2.905000 ;
      RECT 4.150000  2.395000  4.480000 3.245000 ;
      RECT 4.160000  0.265000  7.930000 0.595000 ;
      RECT 4.650000  2.225000  4.840000 3.075000 ;
      RECT 5.010000  2.445000  5.680000 3.245000 ;
      RECT 5.850000  2.225000  6.040000 3.075000 ;
      RECT 6.210000  2.395000  6.900000 3.245000 ;
      RECT 6.310000  0.765000  8.810000 0.815000 ;
      RECT 6.310000  0.815000  9.670000 1.040000 ;
      RECT 7.000000  1.605000  9.910000 1.775000 ;
      RECT 7.000000  1.775000  7.260000 2.045000 ;
      RECT 7.070000  2.225000  7.260000 3.075000 ;
      RECT 7.430000  1.945000  7.760000 3.245000 ;
      RECT 7.930000  1.775000  8.120000 3.075000 ;
      RECT 8.120000  0.085000  8.450000 0.595000 ;
      RECT 8.290000  1.945000  8.620000 3.245000 ;
      RECT 8.620000  0.255000  8.810000 0.765000 ;
      RECT 8.790000  1.775000  8.980000 3.075000 ;
      RECT 8.980000  0.085000  9.310000 0.595000 ;
      RECT 9.150000  1.945000  9.480000 3.245000 ;
      RECT 9.480000  0.255000  9.670000 0.815000 ;
      RECT 9.650000  1.775000  9.910000 3.075000 ;
      RECT 9.840000  0.085000 10.170000 1.040000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__a32oi_4
