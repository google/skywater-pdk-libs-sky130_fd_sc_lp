* File: sky130_fd_sc_lp__o2bb2a_1.spice
* Created: Wed Sep  2 10:21:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2a_1.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2a_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_80_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.21 AS=0.2226 PD=1.76667 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1010 A_237_131# N_A1_N_M1010_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.105 PD=0.66 PS=0.883333 NRD=18.564 NRS=55.704 M=1 R=2.8
+ SA=75000.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_286_492#_M1007_d N_A2_N_M1007_g A_237_131# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_506_47#_M1003_d N_A_286_492#_M1003_g N_A_80_21#_M1003_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_B2_M1006_g N_A_506_47#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_506_47#_M1000_d N_B1_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_80_21#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3969 AS=0.3339 PD=2.985 PS=3.05 NRD=17.1981 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_A_286_492#_M1009_d N_A1_N_M1009_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1323 PD=0.7 PS=0.995 NRD=0 NRS=228.658 M=1 R=2.8
+ SA=75001.1 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A2_N_M1004_g N_A_286_492#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0588 PD=0.94 PS=0.7 NRD=63.3158 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_80_21#_M1001_d N_A_286_492#_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1092 PD=0.7 PS=0.94 NRD=0 NRS=49.25 M=1 R=2.8 SA=75002.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_592_492# N_B2_M1008_g N_A_80_21#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g A_592_492# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o2bb2a_1.pxi.spice"
*
.ends
*
*
