* File: sky130_fd_sc_lp__fah_1.pex.spice
* Created: Wed Sep  2 09:53:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FAH_1%CI 3 7 9 12
r43 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.685
+ $X2=1.15 $Y2=1.85
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.685
+ $X2=1.15 $Y2=1.52
r45 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.685 $X2=1.15 $Y2=1.685
r46 7 15 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.195 $Y=2.595
+ $X2=1.195 $Y2=1.85
r47 3 14 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=1.12 $Y=0.995
+ $X2=1.12 $Y2=1.52
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_84_21# 1 2 9 11 13 14 16 18 21 24 25 26 27
+ 30 31 32 33 36 38 41 42 50 51
c156 51 0 2.59569e-20 $X=5.885 $Y=0.745
c157 50 0 1.67676e-19 $X=6.05 $Y=0.705
c158 42 0 1.37374e-19 $X=3.2 $Y=2.065
r159 50 51 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.05 $Y=0.745
+ $X2=5.885 $Y2=0.745
r160 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.2 $Y=2.065
+ $X2=3.2 $Y2=2.35
r161 41 53 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=2.03 $Y=1.985
+ $X2=1.75 $Y2=1.985
r162 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.985 $X2=2.03 $Y2=1.985
r163 38 51 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=4.19 $Y=0.7
+ $X2=5.885 $Y2=0.7
r164 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=0.615
+ $X2=4.19 $Y2=0.7
r165 35 36 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.105 $Y=0.435
+ $X2=4.105 $Y2=0.615
r166 34 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=2.35
+ $X2=3.2 $Y2=2.35
r167 33 48 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.32 $Y=2.35
+ $X2=4.32 $Y2=2.435
r168 33 34 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=4.195 $Y=2.35
+ $X2=3.285 $Y2=2.35
r169 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=0.35
+ $X2=4.105 $Y2=0.435
r170 31 32 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.02 $Y=0.35
+ $X2=2.79 $Y2=0.35
r171 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.705 $Y=0.435
+ $X2=2.79 $Y2=0.35
r172 29 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.705 $Y=0.435
+ $X2=2.705 $Y2=0.85
r173 28 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.065
+ $X2=2.03 $Y2=2.065
r174 27 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.065
+ $X2=3.2 $Y2=2.065
r175 27 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.115 $Y=2.065
+ $X2=2.195 $Y2=2.065
r176 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.62 $Y=0.935
+ $X2=2.705 $Y2=0.85
r177 25 26 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.62 $Y=0.935
+ $X2=2.195 $Y2=0.935
r178 24 40 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.98 $X2=2.03
+ $Y2=2.065
r179 23 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.03 $Y=1.02
+ $X2=2.195 $Y2=0.935
r180 23 24 33.5256 $w=3.28e-07 $l=9.6e-07 $layer=LI1_cond $X=2.03 $Y=1.02
+ $X2=2.03 $Y2=1.98
r181 19 21 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.63 $Y=1.29
+ $X2=1.75 $Y2=1.29
r182 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.82
+ $X2=1.75 $Y2=1.985
r183 17 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.365
+ $X2=1.75 $Y2=1.29
r184 17 18 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.75 $Y=1.365
+ $X2=1.75 $Y2=1.82
r185 16 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.63 $Y=1.215
+ $X2=1.63 $Y2=1.29
r186 15 16 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.63 $Y=0.255
+ $X2=1.63 $Y2=1.215
r187 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.555 $Y=0.18
+ $X2=1.63 $Y2=0.255
r188 13 14 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=1.555 $Y=0.18
+ $X2=0.57 $Y2=0.18
r189 9 11 805.043 $w=1.5e-07 $l=1.57e-06 $layer=POLY_cond $X=0.495 $Y=0.895
+ $X2=0.495 $Y2=2.465
r190 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.57 $Y2=0.18
r191 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.495 $Y2=0.895
r192 2 48 600 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=2.18 $X2=4.36 $Y2=2.435
r193 1 50 182 $w=1.7e-07 $l=2.8788e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.635 $X2=6.05 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_413_34# 1 2 7 9 12 14 15 16 19 20 21 23 24
+ 25 26 27 28 29 30 39
c135 39 0 9.39508e-20 $X=6.06 $Y=2.415
c136 27 0 2.88995e-19 $X=5.14 $Y=2.33
c137 26 0 1.27296e-19 $X=5.14 $Y=1.575
c138 14 0 1.7772e-20 $X=2.215 $Y=1.415
r139 39 42 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=6.06 $Y=2.415
+ $X2=6.06 $Y2=2.52
r140 36 38 4.22511 $w=2.31e-07 $l=8e-08 $layer=LI1_cond $X=5.067 $Y=1.05
+ $X2=5.067 $Y2=1.13
r141 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.415 $X2=2.54 $Y2=1.415
r142 30 33 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=1.285
+ $X2=2.54 $Y2=1.415
r143 28 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.895 $Y=2.415
+ $X2=6.06 $Y2=2.415
r144 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.895 $Y=2.415
+ $X2=5.225 $Y2=2.415
r145 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=2.33
+ $X2=5.225 $Y2=2.415
r146 26 38 24.3769 $w=2.31e-07 $l=4.80115e-07 $layer=LI1_cond $X=5.14 $Y=1.575
+ $X2=5.067 $Y2=1.13
r147 26 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.14 $Y=1.575
+ $X2=5.14 $Y2=2.33
r148 24 36 2.5345 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=4.91 $Y=1.05
+ $X2=5.067 $Y2=1.05
r149 24 25 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.91 $Y=1.05
+ $X2=3.84 $Y2=1.05
r150 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.755 $Y=0.965
+ $X2=3.84 $Y2=1.05
r151 22 23 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.755 $Y=0.785
+ $X2=3.755 $Y2=0.965
r152 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=0.7
+ $X2=3.755 $Y2=0.785
r153 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.67 $Y=0.7
+ $X2=3.14 $Y2=0.7
r154 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.055 $Y=0.785
+ $X2=3.14 $Y2=0.7
r155 18 19 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.055 $Y=0.785
+ $X2=3.055 $Y2=1.2
r156 17 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=1.285
+ $X2=2.54 $Y2=1.285
r157 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.97 $Y=1.285
+ $X2=3.055 $Y2=1.2
r158 16 17 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.97 $Y=1.285
+ $X2=2.705 $Y2=1.285
r159 15 34 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.64 $Y=1.415
+ $X2=2.54 $Y2=1.415
r160 14 34 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=2.215 $Y=1.415
+ $X2=2.54 $Y2=1.415
r161 10 15 21.1694 $w=3.64e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.715 $Y=1.58
+ $X2=2.64 $Y2=1.415
r162 10 12 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=2.715 $Y=1.58
+ $X2=2.715 $Y2=2.465
r163 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.14 $Y=1.25
+ $X2=2.215 $Y2=1.415
r164 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.14 $Y=1.25 $X2=2.14
+ $Y2=0.72
r165 2 42 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=1.895 $X2=6.06 $Y2=2.52
r166 1 38 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=4.935
+ $Y=0.635 $X2=5.075 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_239_135# 1 2 3 4 15 17 18 21 24 25 31 33 35
+ 37 40 42 45 46 48 50 53 54 55 57 59 60 63 67 75 77 83
c223 60 0 1.7772e-20 $X=1.495 $Y=2.075
c224 55 0 1.59085e-19 $X=6.215 $Y=2.045
c225 53 0 1.89042e-19 $X=6.13 $Y=1.96
c226 37 0 3.54844e-19 $X=4.16 $Y=1.515
c227 21 0 1.116e-19 $X=3.485 $Y=2.355
r228 82 83 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=2.872
+ $X2=5.68 $Y2=2.872
r229 77 79 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=1.055
+ $X2=5.505 $Y2=1.14
r230 67 69 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.44 $Y=2.7
+ $X2=3.44 $Y2=2.98
r231 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.85 $Y=2.415
+ $X2=2.85 $Y2=2.7
r232 59 61 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=1.495 $Y=2.395
+ $X2=1.495 $Y2=2.415
r233 59 60 13.7257 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=1.495 $Y=2.395
+ $X2=1.495 $Y2=2.075
r234 56 57 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.49 $Y=2.13
+ $X2=6.49 $Y2=2.895
r235 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.405 $Y=2.045
+ $X2=6.49 $Y2=2.13
r236 54 55 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.405 $Y=2.045
+ $X2=6.215 $Y2=2.045
r237 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.13 $Y=1.96
+ $X2=6.215 $Y2=2.045
r238 52 53 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=6.13 $Y=1.225
+ $X2=6.13 $Y2=1.96
r239 50 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.405 $Y=2.98
+ $X2=6.49 $Y2=2.895
r240 50 83 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.405 $Y=2.98
+ $X2=5.68 $Y2=2.98
r241 49 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.67 $Y=1.14
+ $X2=5.505 $Y2=1.14
r242 48 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.045 $Y=1.14
+ $X2=6.13 $Y2=1.225
r243 48 49 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.045 $Y=1.14
+ $X2=5.67 $Y2=1.14
r244 47 75 3.37808 $w=2.77e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=2.872
+ $X2=4.79 $Y2=2.872
r245 46 82 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=5.488 $Y=2.872
+ $X2=5.515 $Y2=2.872
r246 46 47 18.3493 $w=3.83e-07 $l=6.13e-07 $layer=LI1_cond $X=5.488 $Y=2.872
+ $X2=4.875 $Y2=2.872
r247 45 75 3.15366 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=4.79 $Y=2.68
+ $X2=4.79 $Y2=2.872
r248 44 45 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.79 $Y=1.98 $X2=4.79
+ $Y2=2.68
r249 43 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.33 $Y=1.895
+ $X2=4.245 $Y2=1.895
r250 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.705 $Y=1.895
+ $X2=4.79 $Y2=1.98
r251 42 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.705 $Y=1.895
+ $X2=4.33 $Y2=1.895
r252 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.98
+ $Y=1.515 $X2=3.98 $Y2=1.515
r253 37 73 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.245 $Y=1.515
+ $X2=4.245 $Y2=1.895
r254 37 39 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.16 $Y=1.515
+ $X2=3.98 $Y2=1.515
r255 36 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.98
+ $X2=3.44 $Y2=2.98
r256 35 75 3.37808 $w=2.77e-07 $l=1.44375e-07 $layer=LI1_cond $X=4.705 $Y=2.98
+ $X2=4.79 $Y2=2.872
r257 35 36 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=4.705 $Y=2.98
+ $X2=3.525 $Y2=2.98
r258 34 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=2.7
+ $X2=2.85 $Y2=2.7
r259 33 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=2.7
+ $X2=3.44 $Y2=2.7
r260 33 34 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.355 $Y=2.7
+ $X2=2.935 $Y2=2.7
r261 32 61 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.665 $Y=2.415
+ $X2=1.495 $Y2=2.415
r262 31 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=2.415
+ $X2=2.85 $Y2=2.415
r263 31 32 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.765 $Y=2.415
+ $X2=1.665 $Y2=2.415
r264 29 60 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.58 $Y=1.34
+ $X2=1.58 $Y2=2.075
r265 25 29 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.495 $Y=1.215
+ $X2=1.58 $Y2=1.34
r266 25 27 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=1.495 $Y=1.215
+ $X2=1.335 $Y2=1.215
r267 23 40 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.56 $Y=1.515
+ $X2=3.98 $Y2=1.515
r268 23 24 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.515
+ $X2=3.485 $Y2=1.515
r269 19 24 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.68
+ $X2=3.485 $Y2=1.515
r270 19 21 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.485 $Y=1.68
+ $X2=3.485 $Y2=2.355
r271 17 24 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.41 $Y=1.425
+ $X2=3.485 $Y2=1.515
r272 17 18 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.41 $Y=1.425
+ $X2=3.15 $Y2=1.425
r273 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.075 $Y=1.35
+ $X2=3.15 $Y2=1.425
r274 13 15 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.075 $Y=1.35
+ $X2=3.075 $Y2=0.82
r275 4 82 600 $w=1.7e-07 $l=8.12558e-07 $layer=licon1_PDIFF $count=1 $X=5.26
+ $Y=2.07 $X2=5.515 $Y2=2.765
r276 3 59 600 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=1 $X=1.27
+ $Y=2.095 $X2=1.41 $Y2=2.395
r277 2 77 182 $w=1.7e-07 $l=4.84974e-07 $layer=licon1_NDIFF $count=1 $X=5.365
+ $Y=0.635 $X2=5.505 $Y2=1.055
r278 1 27 182 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.675 $X2=1.335 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_814_384# 1 2 7 9 10 11 13 14 15 19 20 21 25
+ 28 31 32 33 34 36 38 40 41 47 51 52
c186 52 0 2.09421e-19 $X=5.74 $Y=1.57
c187 51 0 3.02499e-19 $X=5.74 $Y=1.57
c188 47 0 3.59697e-19 $X=9.36 $Y=2.035
c189 41 0 3.48127e-19 $X=5.665 $Y=2.035
c190 40 0 2.76112e-20 $X=9.215 $Y=2.035
c191 36 0 1.35512e-19 $X=10.495 $Y=0.935
c192 34 0 1.87437e-19 $X=10.495 $Y=1.09
c193 25 0 5.84493e-20 $X=5.72 $Y=0.955
c194 10 0 1.13792e-19 $X=4.385 $Y=1.995
r195 51 54 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=5.747 $Y=1.57
+ $X2=5.747 $Y2=1.735
r196 51 53 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=5.747 $Y=1.57
+ $X2=5.747 $Y2=1.405
r197 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.74
+ $Y=1.57 $X2=5.74 $Y2=1.57
r198 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=2.035
+ $X2=9.36 $Y2=2.035
r199 44 52 12.0908 $w=4.58e-07 $l=4.65e-07 $layer=LI1_cond $X=5.635 $Y=2.035
+ $X2=5.635 $Y2=1.57
r200 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r201 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r202 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=2.035
+ $X2=9.36 $Y2=2.035
r203 40 41 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=9.215 $Y=2.035
+ $X2=5.665 $Y2=2.035
r204 38 48 20.5974 $w=2.08e-07 $l=3.9e-07 $layer=LI1_cond $X=9.75 $Y=2.045
+ $X2=9.36 $Y2=2.045
r205 34 39 10.2261 $w=3.3e-07 $l=2.55e-07 $layer=LI1_cond $X=10.495 $Y=1.09
+ $X2=10.495 $Y2=1.345
r206 34 36 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.495 $Y=1.09
+ $X2=10.495 $Y2=0.935
r207 32 39 2.92482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.33 $Y=1.345
+ $X2=10.495 $Y2=1.345
r208 32 33 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=10.33 $Y=1.345
+ $X2=9.92 $Y2=1.345
r209 31 38 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.835 $Y=1.94
+ $X2=9.75 $Y2=2.045
r210 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.835 $Y=1.43
+ $X2=9.92 $Y2=1.345
r211 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.835 $Y=1.43
+ $X2=9.835 $Y2=1.94
r212 28 54 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.845 $Y=2.315
+ $X2=5.845 $Y2=1.735
r213 25 53 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.72 $Y=0.955
+ $X2=5.72 $Y2=1.405
r214 22 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.72 $Y=0.265
+ $X2=5.72 $Y2=0.955
r215 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.645 $Y=0.19
+ $X2=5.72 $Y2=0.265
r216 20 21 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.645 $Y=0.19
+ $X2=4.935 $Y2=0.19
r217 17 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.86 $Y=1.385
+ $X2=4.86 $Y2=0.955
r218 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.86 $Y=0.265
+ $X2=4.935 $Y2=0.19
r219 16 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.86 $Y=0.265
+ $X2=4.86 $Y2=0.955
r220 14 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.785 $Y=1.46
+ $X2=4.86 $Y2=1.385
r221 14 15 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.785 $Y=1.46
+ $X2=4.535 $Y2=1.46
r222 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.46 $Y=1.535
+ $X2=4.535 $Y2=1.46
r223 12 13 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=4.46 $Y=1.535
+ $X2=4.46 $Y2=1.92
r224 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.385 $Y=1.995
+ $X2=4.46 $Y2=1.92
r225 10 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.385 $Y=1.995
+ $X2=4.22 $Y2=1.995
r226 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.145 $Y=2.07
+ $X2=4.22 $Y2=1.995
r227 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.145 $Y=2.07
+ $X2=4.145 $Y2=2.6
r228 2 48 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.835 $X2=9.36 $Y2=2.045
r229 1 36 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=10.355
+ $Y=0.595 $X2=10.495 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_1022_362# 1 2 10 11 13 15 16 19 23 24 26 27
+ 30 32 34 35 36 37 46 50 51 58
c197 58 0 1.63712e-19 $X=9.405 $Y=0.78
c198 46 0 1.14729e-19 $X=10.8 $Y=1.665
c199 26 0 9.39508e-20 $X=6.387 $Y=1.26
c200 24 0 4.13992e-20 $X=6.755 $Y=1.26
c201 23 0 1.83464e-19 $X=6.51 $Y=2.315
r202 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.92
+ $Y=0.83 $X2=6.92 $Y2=0.83
r203 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=1.665
+ $X2=10.8 $Y2=1.665
r204 44 58 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=9.405 $Y=1.665
+ $X2=9.405 $Y2=0.78
r205 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.665
r206 40 51 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=6.92 $Y=1.665
+ $X2=6.92 $Y2=0.83
r207 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.665
r208 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.505 $Y=1.665
+ $X2=9.36 $Y2=1.665
r209 36 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=1.665
+ $X2=10.8 $Y2=1.665
r210 36 37 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=10.655 $Y=1.665
+ $X2=9.505 $Y2=1.665
r211 35 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=1.665
+ $X2=6.96 $Y2=1.665
r212 34 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=9.36 $Y2=1.665
r213 34 35 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=7.105 $Y2=1.665
r214 30 47 24.7211 $w=1.9e-07 $l=3.85e-07 $layer=LI1_cond $X=10.415 $Y=1.665
+ $X2=10.8 $Y2=1.665
r215 30 32 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=10.415 $Y=1.78
+ $X2=10.415 $Y2=1.98
r216 29 50 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.92 $Y=1.185
+ $X2=6.92 $Y2=0.83
r217 26 28 82.1715 $w=3.95e-07 $l=4.25e-07 $layer=POLY_cond $X=6.387 $Y=1.26
+ $X2=6.387 $Y2=1.685
r218 26 27 32.8921 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=6.387 $Y=1.26
+ $X2=6.387 $Y2=1.185
r219 25 26 25.5547 $w=1.5e-07 $l=1.98e-07 $layer=POLY_cond $X=6.585 $Y=1.26
+ $X2=6.387 $Y2=1.26
r220 24 29 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.755 $Y=1.26
+ $X2=6.92 $Y2=1.185
r221 24 25 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.755 $Y=1.26
+ $X2=6.585 $Y2=1.26
r222 23 28 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=6.51 $Y=2.315
+ $X2=6.51 $Y2=1.685
r223 21 23 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.51 $Y=3.075
+ $X2=6.51 $Y2=2.315
r224 19 27 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.265 $Y=0.79
+ $X2=6.265 $Y2=1.185
r225 15 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.435 $Y=3.15
+ $X2=6.51 $Y2=3.075
r226 15 16 602.5 $w=1.5e-07 $l=1.175e-06 $layer=POLY_cond $X=6.435 $Y=3.15
+ $X2=5.26 $Y2=3.15
r227 11 13 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=5.29 $Y=1.67
+ $X2=5.29 $Y2=0.955
r228 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.185 $Y=3.075
+ $X2=5.26 $Y2=3.15
r229 8 10 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=5.185 $Y=3.075
+ $X2=5.185 $Y2=2.49
r230 7 11 68.5196 $w=2.04e-07 $l=3.38452e-07 $layer=POLY_cond $X=5.185 $Y=1.96
+ $X2=5.29 $Y2=1.67
r231 7 10 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.185 $Y=1.96
+ $X2=5.185 $Y2=2.49
r232 2 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.275
+ $Y=1.835 $X2=10.415 $Y2=1.98
r233 1 58 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=9.265
+ $Y=0.625 $X2=9.405 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_878_41# 1 2 3 10 11 14 19 20 24 29 32 33 36
+ 38 42 44 46 48 49 51 52 56 57 63
c151 46 0 4.13992e-20 $X=7.265 $Y=2.045
c152 36 0 1.63712e-19 $X=10.28 $Y=1.42
c153 14 0 1.79467e-19 $X=9.145 $Y=2.255
r154 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.2
+ $Y=0.555 $X2=8.2 $Y2=0.555
r155 54 56 12.2561 $w=3.13e-07 $l=3.35e-07 $layer=LI1_cond $X=8.202 $Y=0.89
+ $X2=8.202 $Y2=0.555
r156 53 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=0.975
+ $X2=7.35 $Y2=0.975
r157 52 54 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=8.045 $Y=0.975
+ $X2=8.202 $Y2=0.89
r158 52 53 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.045 $Y=0.975
+ $X2=7.435 $Y2=0.975
r159 50 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=1.06
+ $X2=7.35 $Y2=0.975
r160 50 51 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.35 $Y=1.06 $X2=7.35
+ $Y2=1.96
r161 49 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=0.89
+ $X2=7.35 $Y2=0.975
r162 48 62 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=0.435
+ $X2=7.35 $Y2=0.35
r163 48 49 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=7.35 $Y=0.435
+ $X2=7.35 $Y2=0.89
r164 47 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=2.045
+ $X2=6.84 $Y2=2.045
r165 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.265 $Y=2.045
+ $X2=7.35 $Y2=1.96
r166 46 47 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.265 $Y=2.045
+ $X2=6.925 $Y2=2.045
r167 42 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.13
+ $X2=6.84 $Y2=2.045
r168 42 44 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.84 $Y=2.13
+ $X2=6.84 $Y2=2.9
r169 38 62 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.265 $Y=0.35
+ $X2=7.35 $Y2=0.35
r170 38 40 178.107 $w=1.68e-07 $l=2.73e-06 $layer=LI1_cond $X=7.265 $Y=0.35
+ $X2=4.535 $Y2=0.35
r171 34 36 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=10.2 $Y=1.42
+ $X2=10.28 $Y2=1.42
r172 31 32 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=9.167 $Y=1.375
+ $X2=9.167 $Y2=1.525
r173 30 57 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=8.2 $Y=0.255 $X2=8.2
+ $Y2=0.555
r174 27 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.28 $Y=1.345
+ $X2=10.28 $Y2=1.42
r175 27 29 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.28 $Y=1.345
+ $X2=10.28 $Y2=0.915
r176 26 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.28 $Y=0.255
+ $X2=10.28 $Y2=0.915
r177 22 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.2 $Y=1.495
+ $X2=10.2 $Y2=1.42
r178 22 24 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=10.2 $Y=1.495
+ $X2=10.2 $Y2=2.255
r179 21 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.265 $Y=0.18
+ $X2=9.19 $Y2=0.18
r180 20 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.205 $Y=0.18
+ $X2=10.28 $Y2=0.255
r181 20 21 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=10.205 $Y=0.18
+ $X2=9.265 $Y2=0.18
r182 19 31 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.19 $Y=0.945
+ $X2=9.19 $Y2=1.375
r183 16 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.19 $Y=0.255
+ $X2=9.19 $Y2=0.18
r184 16 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.19 $Y=0.255
+ $X2=9.19 $Y2=0.945
r185 14 32 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=9.145 $Y=2.255
+ $X2=9.145 $Y2=1.525
r186 11 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.365 $Y=0.18
+ $X2=8.2 $Y2=0.255
r187 10 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.115 $Y=0.18
+ $X2=9.19 $Y2=0.18
r188 10 11 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=9.115 $Y=0.18
+ $X2=8.365 $Y2=0.18
r189 3 60 400 $w=1.7e-07 $l=3.51675e-07 $layer=licon1_PDIFF $count=1 $X=6.585
+ $Y=1.895 $X2=6.84 $Y2=2.125
r190 3 44 400 $w=1.7e-07 $l=1.1253e-06 $layer=licon1_PDIFF $count=1 $X=6.585
+ $Y=1.895 $X2=6.84 $Y2=2.9
r191 2 62 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=7.205
+ $Y=0.235 $X2=7.35 $Y2=0.43
r192 1 40 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.205 $X2=4.535 $Y2=0.35
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%B 1 3 4 5 8 12 17 20 22 26 29 31 34 35 38 39
+ 40 41 45
c127 45 0 2.76112e-20 $X=7.87 $Y=2.455
c128 26 0 3.65352e-20 $X=10.71 $Y=0.915
c129 20 0 1.35512e-19 $X=9.62 $Y=0.945
c130 17 0 1.80229e-19 $X=9.575 $Y=2.255
r131 40 41 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.87 $Y=2.405
+ $X2=7.87 $Y2=2.775
r132 40 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.87
+ $Y=2.455 $X2=7.87 $Y2=2.455
r133 37 38 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=9.597 $Y=1.575
+ $X2=9.597 $Y2=1.725
r134 35 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.87 $Y=2.795
+ $X2=7.87 $Y2=2.455
r135 35 36 52.4708 $w=3.3e-07 $l=3.32415e-07 $layer=POLY_cond $X=7.87 $Y=2.795
+ $X2=7.885 $Y2=3.12
r136 34 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.87 $Y=2.29
+ $X2=7.87 $Y2=2.455
r137 30 31 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=7.565 $Y=1.65
+ $X2=7.78 $Y2=1.65
r138 26 29 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=10.71 $Y=0.915
+ $X2=10.71 $Y2=2.255
r139 24 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.71 $Y=3.045
+ $X2=10.71 $Y2=2.255
r140 23 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.65 $Y=3.12
+ $X2=9.575 $Y2=3.12
r141 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.635 $Y=3.12
+ $X2=10.71 $Y2=3.045
r142 22 23 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=10.635 $Y=3.12
+ $X2=9.65 $Y2=3.12
r143 20 37 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=9.62 $Y=0.945
+ $X2=9.62 $Y2=1.575
r144 17 38 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.575 $Y=2.255
+ $X2=9.575 $Y2=1.725
r145 15 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.575 $Y=3.045
+ $X2=9.575 $Y2=3.12
r146 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.575 $Y=3.045
+ $X2=9.575 $Y2=2.255
r147 13 36 12.1867 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=8.035 $Y=3.12
+ $X2=7.885 $Y2=3.12
r148 12 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.5 $Y=3.12
+ $X2=9.575 $Y2=3.12
r149 12 13 751.202 $w=1.5e-07 $l=1.465e-06 $layer=POLY_cond $X=9.5 $Y=3.12
+ $X2=8.035 $Y2=3.12
r150 10 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.78 $Y=1.725
+ $X2=7.78 $Y2=1.65
r151 10 34 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=7.78 $Y=1.725
+ $X2=7.78 $Y2=2.29
r152 6 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.565 $Y=1.575
+ $X2=7.565 $Y2=1.65
r153 6 8 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=7.565 $Y=1.575
+ $X2=7.565 $Y2=0.655
r154 4 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.49 $Y=1.65
+ $X2=7.565 $Y2=1.65
r155 4 5 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.49 $Y=1.65 $X2=7.13
+ $Y2=1.65
r156 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.055 $Y=1.725
+ $X2=7.13 $Y2=1.65
r157 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.055 $Y=1.725
+ $X2=7.055 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_2229_269# 1 2 9 11 13 15 16 20 24 28 32 34
c69 28 0 1.6374e-19 $X=11.61 $Y=1.285
c70 11 0 7.27084e-20 $X=11.255 $Y=1.345
r71 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.61
+ $Y=1.51 $X2=11.61 $Y2=1.51
r72 28 31 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=11.61 $Y=1.285
+ $X2=11.61 $Y2=1.51
r73 24 26 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=13.16 $Y=2.19
+ $X2=13.16 $Y2=2.9
r74 22 34 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.16 $Y=1.37
+ $X2=13.16 $Y2=1.285
r75 22 24 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=13.16 $Y=1.37
+ $X2=13.16 $Y2=2.19
r76 18 34 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.16 $Y=1.2
+ $X2=13.16 $Y2=1.285
r77 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=13.16 $Y=1.2
+ $X2=13.16 $Y2=0.505
r78 17 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.775 $Y=1.285
+ $X2=11.61 $Y2=1.285
r79 16 34 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.995 $Y=1.285
+ $X2=13.16 $Y2=1.285
r80 16 17 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=12.995 $Y=1.285
+ $X2=11.775 $Y2=1.285
r81 14 32 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=11.33 $Y=1.51
+ $X2=11.61 $Y2=1.51
r82 14 15 5.03009 $w=3.3e-07 $l=9.3e-08 $layer=POLY_cond $X=11.33 $Y=1.51
+ $X2=11.237 $Y2=1.51
r83 11 15 37.0704 $w=1.5e-07 $l=1.73767e-07 $layer=POLY_cond $X=11.255 $Y=1.345
+ $X2=11.237 $Y2=1.51
r84 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.255 $Y=1.345
+ $X2=11.255 $Y2=0.815
r85 7 15 37.0704 $w=1.5e-07 $l=1.73292e-07 $layer=POLY_cond $X=11.22 $Y=1.675
+ $X2=11.237 $Y2=1.51
r86 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.22 $Y=1.675
+ $X2=11.22 $Y2=2.465
r87 2 26 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=2.045 $X2=13.16 $Y2=2.9
r88 2 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=2.045 $X2=13.16 $Y2=2.19
r89 1 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.02
+ $Y=0.36 $X2=13.16 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A 3 7 9 13 17 19 20 22 26
c53 22 0 1.27205e-19 $X=12.425 $Y=1.625
r54 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.425 $Y=1.715
+ $X2=12.425 $Y2=1.88
r55 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.425
+ $Y=1.715 $X2=12.425 $Y2=1.715
r56 22 25 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.425 $Y=1.625
+ $X2=12.425 $Y2=1.715
r57 22 23 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.425 $Y=1.625
+ $X2=12.425 $Y2=1.55
r58 20 26 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=12.24 $Y=1.715
+ $X2=12.425 $Y2=1.715
r59 15 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.945 $Y=1.7
+ $X2=12.945 $Y2=1.625
r60 15 17 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=12.945 $Y=1.7
+ $X2=12.945 $Y2=2.545
r61 11 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.945 $Y=1.55
+ $X2=12.945 $Y2=1.625
r62 11 13 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=12.945 $Y=1.55
+ $X2=12.945 $Y2=0.68
r63 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.59 $Y=1.625
+ $X2=12.425 $Y2=1.625
r64 9 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.87 $Y=1.625
+ $X2=12.945 $Y2=1.625
r65 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.87 $Y=1.625
+ $X2=12.59 $Y2=1.625
r66 7 27 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=12.515 $Y=2.545
+ $X2=12.515 $Y2=1.88
r67 3 23 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=12.515 $Y=0.68
+ $X2=12.515 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%SUM 1 2 7 8 9 10 11 12 13
r15 13 39 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.28 $Y=2.775
+ $X2=0.28 $Y2=2.9
r16 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.775
r17 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.28 $Y=1.98
+ $X2=0.28 $Y2=2.405
r18 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=1.98
r19 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.295
+ $X2=0.28 $Y2=1.665
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=0.925 $X2=0.28
+ $Y2=1.295
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=0.555 $X2=0.28
+ $Y2=0.925
r22 2 39 400 $w=1.7e-07 $l=1.13519e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.9
r23 2 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.98
r24 1 7 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.475 $X2=0.28 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%VPWR 1 2 3 4 5 18 22 26 28 32 35 36 37 39 44
+ 53 62 63 66 69 76 79
c131 69 0 7.74056e-20 $X=3.01 $Y=3.05
c132 63 0 3.41944e-20 $X=13.2 $Y=3.33
r133 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r134 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r135 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r136 72 73 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r137 69 72 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.01 $Y=3.05
+ $X2=3.01 $Y2=3.33
r138 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r140 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r141 60 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.815 $Y=3.33
+ $X2=12.73 $Y2=3.33
r142 60 62 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.815 $Y=3.33
+ $X2=13.2 $Y2=3.33
r143 59 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r144 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r145 56 59 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=11.28 $Y2=3.33
r146 55 58 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=11.28 $Y2=3.33
r147 55 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r148 53 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.62 $Y=3.33
+ $X2=11.745 $Y2=3.33
r149 53 58 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.62 $Y=3.33
+ $X2=11.28 $Y2=3.33
r150 52 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r151 51 52 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r152 49 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.01 $Y2=3.33
r153 49 51 246.936 $w=1.68e-07 $l=3.785e-06 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=6.96 $Y2=3.33
r154 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r155 48 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=0.72 $Y2=3.33
r156 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r157 45 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.71 $Y2=3.33
r158 45 47 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=2.64 $Y2=3.33
r159 44 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.01 $Y2=3.33
r160 44 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.64 $Y2=3.33
r161 42 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r162 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r163 39 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.71 $Y2=3.33
r164 39 41 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r165 37 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r166 37 73 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=3.12 $Y2=3.33
r167 35 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=6.96 $Y2=3.33
r168 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=7.27 $Y2=3.33
r169 34 55 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.435 $Y=3.33
+ $X2=7.44 $Y2=3.33
r170 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=3.33
+ $X2=7.27 $Y2=3.33
r171 30 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.73 $Y=3.245
+ $X2=12.73 $Y2=3.33
r172 30 32 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=12.73 $Y=3.245
+ $X2=12.73 $Y2=2.225
r173 29 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.87 $Y=3.33
+ $X2=11.745 $Y2=3.33
r174 28 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.645 $Y=3.33
+ $X2=12.73 $Y2=3.33
r175 28 29 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=12.645 $Y=3.33
+ $X2=11.87 $Y2=3.33
r176 24 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.745 $Y=3.245
+ $X2=11.745 $Y2=3.33
r177 24 26 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=11.745 $Y=3.245
+ $X2=11.745 $Y2=3.025
r178 20 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.27 $Y=3.245
+ $X2=7.27 $Y2=3.33
r179 20 22 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=7.27 $Y=3.245
+ $X2=7.27 $Y2=2.475
r180 16 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=3.33
r181 16 18 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=2.545
r182 5 32 300 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=2 $X=12.59
+ $Y=2.045 $X2=12.73 $Y2=2.225
r183 4 26 600 $w=1.7e-07 $l=1.37986e-06 $layer=licon1_PDIFF $count=1 $X=11.295
+ $Y=1.835 $X2=11.705 $Y2=3.025
r184 3 22 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=7.13
+ $Y=1.835 $X2=7.27 $Y2=2.475
r185 2 69 600 $w=1.7e-07 $l=1.32043e-06 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.835 $X2=3.01 $Y2=3.05
r186 1 18 300 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%COUT 1 2 8 9 10 12 13 14 17 20 24
r77 24 27 2.72626 $w=3.58e-07 $l=8e-08 $layer=LI1_cond $X=1.802 $Y=0.555
+ $X2=1.802 $Y2=0.475
r78 20 22 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=2.46 $Y=2.87
+ $X2=2.46 $Y2=2.98
r79 15 17 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.72 $Y=2.115
+ $X2=1.06 $Y2=2.115
r80 13 22 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.335 $Y=2.98
+ $X2=2.46 $Y2=2.98
r81 13 14 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.335 $Y=2.98
+ $X2=1.145 $Y2=2.98
r82 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.895
+ $X2=1.145 $Y2=2.98
r83 11 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=2.2 $X2=1.06
+ $Y2=2.115
r84 11 12 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.06 $Y=2.2
+ $X2=1.06 $Y2=2.895
r85 9 24 9.20112 $w=3.58e-07 $l=3.99824e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.802 $Y2=0.555
r86 9 10 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=0.805 $Y2=0.825
r87 8 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.03 $X2=0.72
+ $Y2=2.115
r88 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=0.91
+ $X2=0.805 $Y2=0.825
r89 7 8 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=0.72 $Y=0.91 $X2=0.72
+ $Y2=2.03
r90 2 20 600 $w=1.7e-07 $l=1.10512e-06 $layer=licon1_PDIFF $count=1 $X=2.355
+ $Y=1.835 $X2=2.5 $Y2=2.87
r91 1 27 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=1.78
+ $Y=0.3 $X2=1.925 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_630_100# 1 2 3 12 16 18 19 21 22 28 34
c94 34 0 5.84493e-20 $X=6.48 $Y=0.87
c95 22 0 1.99242e-19 $X=3.265 $Y=1.665
c96 21 0 1.37374e-19 $X=6.335 $Y=1.665
c97 12 0 2.52136e-20 $X=3.405 $Y=1.13
r98 29 34 48.9848 $w=1.78e-07 $l=7.95e-07 $layer=LI1_cond $X=6.485 $Y=1.665
+ $X2=6.485 $Y2=0.87
r99 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r100 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r101 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r102 21 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r103 21 22 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=3.265 $Y2=1.665
r104 19 25 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=3.32 $Y=1.665
+ $X2=3.12 $Y2=1.665
r105 18 20 18.9213 $w=2.16e-07 $l=3.35e-07 $layer=LI1_cond $X=3.477 $Y=1.665
+ $X2=3.477 $Y2=2
r106 18 19 0.329861 $w=2.3e-07 $l=1.57e-07 $layer=LI1_cond $X=3.477 $Y=1.665
+ $X2=3.32 $Y2=1.665
r107 14 20 2.14224 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=3.635 $Y=2
+ $X2=3.477 $Y2=2
r108 14 16 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.635 $Y=2
+ $X2=3.815 $Y2=2
r109 10 18 7.08249 $w=2.16e-07 $l=1.46646e-07 $layer=LI1_cond $X=3.405 $Y=1.55
+ $X2=3.477 $Y2=1.665
r110 10 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.405 $Y=1.55
+ $X2=3.405 $Y2=1.13
r111 3 16 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.855 $X2=3.815 $Y2=2
r112 2 34 182 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.47 $X2=6.48 $Y2=0.87
r113 1 12 182 $w=1.7e-07 $l=7.46693e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.5 $X2=3.405 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_1741_367# 1 2 3 4 16 19 21 26 29 32 34 35 41
+ 45
r78 35 37 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.85 $Y=2.415
+ $X2=8.85 $Y2=2.53
r79 33 34 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.872 $Y=1.59
+ $X2=8.872 $Y2=1.76
r80 32 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.18 $Y=1.96
+ $X2=11.18 $Y2=2.045
r81 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.18 $Y=1.37
+ $X2=11.18 $Y2=1.285
r82 31 32 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.18 $Y=1.37
+ $X2=11.18 $Y2=1.96
r83 27 45 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=11 $Y=1.285
+ $X2=11.18 $Y2=1.285
r84 27 29 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=11 $Y=1.2 $X2=11
+ $Y2=0.935
r85 24 26 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=10.925 $Y=2.33
+ $X2=10.925 $Y2=2.23
r86 23 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.925 $Y=2.045
+ $X2=11.18 $Y2=2.045
r87 23 26 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=10.925 $Y=2.13
+ $X2=10.925 $Y2=2.23
r88 22 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=2.415
+ $X2=8.85 $Y2=2.415
r89 21 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.76 $Y=2.415
+ $X2=10.925 $Y2=2.33
r90 21 22 113.845 $w=1.68e-07 $l=1.745e-06 $layer=LI1_cond $X=10.76 $Y=2.415
+ $X2=9.015 $Y2=2.415
r91 19 33 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=8.975 $Y=0.78
+ $X2=8.975 $Y2=1.59
r92 16 34 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=8.85 $Y=1.98
+ $X2=8.85 $Y2=1.76
r93 14 35 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=2.33
+ $X2=8.85 $Y2=2.415
r94 14 16 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.85 $Y=2.33
+ $X2=8.85 $Y2=1.98
r95 4 26 600 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=10.785
+ $Y=1.835 $X2=10.925 $Y2=2.23
r96 3 37 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.835 $X2=8.85 $Y2=2.53
r97 3 16 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.835 $X2=8.85 $Y2=1.98
r98 2 29 182 $w=1.7e-07 $l=4.49778e-07 $layer=licon1_NDIFF $count=1 $X=10.785
+ $Y=0.595 $X2=11.04 $Y2=0.935
r99 1 19 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=8.83
+ $Y=0.625 $X2=8.975 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%A_1930_367# 1 2 3 4 14 15 16 18 19 20 23 25 27
+ 30 31 33 34 37 41 47 50 54 55 59
c147 59 0 1.25754e-19 $X=12.3 $Y=2.595
r148 55 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.355 $Y=2.595
+ $X2=11.355 $Y2=2.765
r149 50 52 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=9.905 $Y=2.765
+ $X2=9.905 $Y2=2.96
r150 45 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.42 $Y=1.325
+ $X2=8.625 $Y2=1.325
r151 39 59 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.3 $Y=2.51
+ $X2=12.3 $Y2=2.595
r152 39 41 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=12.3 $Y=2.51
+ $X2=12.3 $Y2=2.225
r153 35 37 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=12.3 $Y=0.85
+ $X2=12.3 $Y2=0.505
r154 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.135 $Y=0.935
+ $X2=12.3 $Y2=0.85
r155 33 34 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=12.135 $Y=0.935
+ $X2=11.475 $Y2=0.935
r156 32 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.44 $Y=2.595
+ $X2=11.355 $Y2=2.595
r157 31 59 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.135 $Y=2.595
+ $X2=12.3 $Y2=2.595
r158 31 32 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=12.135 $Y=2.595
+ $X2=11.44 $Y2=2.595
r159 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.39 $Y=0.85
+ $X2=11.475 $Y2=0.935
r160 29 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=11.39 $Y=0.435
+ $X2=11.39 $Y2=0.85
r161 28 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.115 $Y=0.35
+ $X2=9.95 $Y2=0.35
r162 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.305 $Y=0.35
+ $X2=11.39 $Y2=0.435
r163 27 28 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=11.305 $Y=0.35
+ $X2=10.115 $Y2=0.35
r164 26 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.07 $Y=2.765
+ $X2=9.905 $Y2=2.765
r165 25 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.27 $Y=2.765
+ $X2=11.355 $Y2=2.765
r166 25 26 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=11.27 $Y=2.765
+ $X2=10.07 $Y2=2.765
r167 21 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=0.435
+ $X2=9.95 $Y2=0.35
r168 21 23 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=9.95 $Y=0.435
+ $X2=9.95 $Y2=0.825
r169 19 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.785 $Y=0.35
+ $X2=9.95 $Y2=0.35
r170 19 20 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=9.785 $Y=0.35
+ $X2=8.71 $Y2=0.35
r171 18 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.625 $Y=1.24
+ $X2=8.625 $Y2=1.325
r172 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.625 $Y=0.435
+ $X2=8.71 $Y2=0.35
r173 17 18 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.625 $Y=0.435
+ $X2=8.625 $Y2=1.24
r174 15 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.74 $Y=2.96
+ $X2=9.905 $Y2=2.96
r175 15 16 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=9.74 $Y=2.96
+ $X2=8.505 $Y2=2.96
r176 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=2.875
+ $X2=8.505 $Y2=2.96
r177 13 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=1.41
+ $X2=8.42 $Y2=1.325
r178 13 14 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=8.42 $Y=1.41
+ $X2=8.42 $Y2=2.875
r179 4 41 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=12.155
+ $Y=2.045 $X2=12.3 $Y2=2.225
r180 3 50 600 $w=1.7e-07 $l=1.04979e-06 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.835 $X2=9.905 $Y2=2.765
r181 2 37 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.155
+ $Y=0.36 $X2=12.3 $Y2=0.505
r182 1 23 182 $w=1.7e-07 $l=3.40624e-07 $layer=licon1_NDIFF $count=1 $X=9.695
+ $Y=0.625 $X2=9.95 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__FAH_1%VGND 1 2 3 4 5 20 24 28 32 34 38 41 42 44 45
+ 46 61 70 71 74 77 80
r122 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r123 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r124 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r125 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 71 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r127 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r128 68 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=12.73 $Y2=0
r129 68 70 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=13.2 $Y2=0
r130 67 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r131 66 67 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r132 64 67 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=11.28 $Y2=0
r133 63 66 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=11.28 $Y2=0
r134 63 64 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r135 61 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.655 $Y=0
+ $X2=11.78 $Y2=0
r136 61 66 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.655 $Y=0
+ $X2=11.28 $Y2=0
r137 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r138 59 60 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r139 56 59 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=7.44
+ $Y2=0
r140 56 57 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r141 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r142 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r143 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r144 51 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r145 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r146 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r147 48 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.825
+ $Y2=0
r148 48 50 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r149 46 60 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.72 $Y=0 $X2=7.44
+ $Y2=0
r150 46 57 1.13724 $w=4.9e-07 $l=4.08e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=2.64
+ $Y2=0
r151 44 59 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.615 $Y=0
+ $X2=7.44 $Y2=0
r152 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.74
+ $Y2=0
r153 43 63 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.865 $Y=0 $X2=7.92
+ $Y2=0
r154 43 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.865 $Y=0 $X2=7.74
+ $Y2=0
r155 41 53 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.16
+ $Y2=0
r156 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.355
+ $Y2=0
r157 40 56 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.44 $Y=0 $X2=2.64
+ $Y2=0
r158 40 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0 $X2=2.355
+ $Y2=0
r159 36 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.73 $Y=0.085
+ $X2=12.73 $Y2=0
r160 36 38 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=12.73 $Y=0.085
+ $X2=12.73 $Y2=0.505
r161 35 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=11.78 $Y2=0
r162 34 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.645 $Y=0
+ $X2=12.73 $Y2=0
r163 34 35 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=12.645 $Y=0
+ $X2=11.905 $Y2=0
r164 30 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.78 $Y=0.085
+ $X2=11.78 $Y2=0
r165 30 32 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=11.78 $Y=0.085
+ $X2=11.78 $Y2=0.505
r166 26 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.74 $Y=0.085
+ $X2=7.74 $Y2=0
r167 26 28 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=7.74 $Y=0.085
+ $X2=7.74 $Y2=0.46
r168 22 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=0.085
+ $X2=2.355 $Y2=0
r169 22 24 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.355 $Y=0.085
+ $X2=2.355 $Y2=0.475
r170 18 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r171 18 20 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.475
r172 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.59
+ $Y=0.36 $X2=12.73 $Y2=0.505
r173 4 32 182 $w=1.7e-07 $l=4.61736e-07 $layer=licon1_NDIFF $count=1 $X=11.33
+ $Y=0.395 $X2=11.74 $Y2=0.505
r174 3 28 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=7.64
+ $Y=0.235 $X2=7.78 $Y2=0.46
r175 2 24 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.3 $X2=2.355 $Y2=0.475
r176 1 20 182 $w=1.7e-07 $l=2.55e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.475 $X2=0.825 $Y2=0.475
.ends

