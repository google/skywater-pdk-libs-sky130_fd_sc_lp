* NGSPICE file created from sky130_fd_sc_lp__sdfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 a_1445_324# a_1295_379# a_1752_60# VNB nshort w=640000u l=150000u
+  ad=3.70575e+11p pd=2.82e+06u as=3.648e+11p ps=3.7e+06u
M1001 a_1996_379# a_1295_379# a_1445_324# VPB phighvt w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=8.358e+11p ps=3.67e+06u
M1002 VPWR a_2449_137# a_3279_367# VPB phighvt w=640000u l=150000u
+  ad=3.7737e+12p pd=2.813e+07u as=1.824e+11p ps=1.85e+06u
M1003 VPWR a_1926_21# a_1996_379# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Q a_3279_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1005 a_1295_379# a_995_66# a_200_119# VNB nshort w=420000u l=150000u
+  ad=2.6775e+11p pd=2.18e+06u as=2.961e+11p ps=3.09e+06u
M1006 VGND RESET_B a_1926_21# VNB nshort w=420000u l=150000u
+  ad=2.3603e+12p pd=1.951e+07u as=1.197e+11p ps=1.41e+06u
M1007 a_314_119# D a_200_119# VNB nshort w=420000u l=150000u
+  ad=2.058e+11p pd=1.82e+06u as=0p ps=0u
M1008 a_1752_60# a_1926_21# a_1445_324# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_1445_324# a_1397_379# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 a_328_429# SCE VGND VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
M1011 a_2449_137# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1012 a_200_119# SCE a_122_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 VGND a_328_429# a_314_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2401_163# a_995_66# a_2299_119# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.139e+11p ps=2e+06u
M1015 a_838_50# CLK_N VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1016 a_2299_119# a_838_50# a_2198_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.272e+11p ps=1.99e+06u
M1017 a_2636_119# a_1926_21# a_2449_137# VNB nshort w=640000u l=150000u
+  ad=5.3795e+11p pd=4.52e+06u as=3.5265e+11p ps=2.65e+06u
M1018 VPWR a_838_50# a_995_66# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1019 VPWR RESET_B a_1926_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1020 Q_N a_2449_137# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1021 Q_N a_2449_137# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1022 a_2636_119# SET_B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_3279_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1024 VPWR SCD a_27_474# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.616e+11p ps=3.69e+06u
M1025 VGND a_2449_137# a_2401_163# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_2401_506# a_838_50# a_2299_119# VPB phighvt w=420000u l=150000u
+  ad=2.793e+11p pd=2.17e+06u as=2.6985e+11p ps=2.4e+06u
M1027 a_2198_119# a_1445_324# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1439_104# a_838_50# a_1295_379# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=0p ps=0u
M1029 a_838_50# CLK_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1030 a_1445_324# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_474# a_328_429# a_200_119# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.968e+11p ps=3.24e+06u
M1032 a_122_119# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1295_379# a_838_50# a_200_119# VPB phighvt w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1034 a_1397_379# a_995_66# a_1295_379# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1752_60# SET_B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_2449_137# a_2299_119# a_2636_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_2449_137# a_2401_506# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_2299_119# a_995_66# a_2198_379# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=3.33725e+11p ps=2.88e+06u
M1039 VGND a_838_50# a_995_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.239e+11p ps=1.43e+06u
M1040 VGND a_1445_324# a_1439_104# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_2449_137# a_3279_367# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1042 a_200_474# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1043 a_2198_379# a_1445_324# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR a_1926_21# a_2798_451# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1045 a_2798_451# a_2299_119# a_2449_137# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_200_119# D a_200_474# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_328_429# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
.ends

