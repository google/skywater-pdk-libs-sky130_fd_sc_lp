* File: sky130_fd_sc_lp__busdriver2_20.pex.spice
* Created: Fri Aug 28 10:13:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%TE_B 1 3 6 8 10 12 15 17 18 25
c40 15 0 5.76855e-20 $X=0.925 $Y=2.465
r41 24 25 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.57 $Y2=1.35
r42 21 24 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.28 $Y=1.35
+ $X2=0.495 $Y2=1.35
r43 18 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.35 $X2=0.28 $Y2=1.35
r44 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.925 $Y=1.335
+ $X2=0.925 $Y2=1.26
r45 13 15 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=0.925 $Y=1.335
+ $X2=0.925 $Y2=2.465
r46 10 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=1.26
r47 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=0.655
r48 8 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.85 $Y=1.26
+ $X2=0.925 $Y2=1.26
r49 8 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.85 $Y=1.26 $X2=0.57
+ $Y2=1.26
r50 4 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.495 $Y2=1.35
r51 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.495 $Y2=2.465
r52 1 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.35
r53 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_114_47# 1 2 9 13 17 19 20 23 27 29
+ 33 35 37 38 39 40 42 43 45 46 48 49 51 52 53 54 56 57 59 60 62 64 65 67 69 70
+ 72 74 75 77 79 80 82 84 85 87 89 90 92 94 99 104 105 106 107 108 109 112 116
+ 122 125 126 131 141
c275 141 0 1.98224e-19 $X=6.15 $Y=1.16
c276 72 0 7.60313e-20 $X=7.47 $Y=0.985
c277 33 0 1.19111e-20 $X=2.645 $Y=2.465
c278 27 0 1.023e-19 $X=2.215 $Y=2.465
c279 19 0 1.91375e-19 $X=2.1 $Y=1.41
r280 140 141 40.661 $w=3.5e-07 $l=1.3e-07 $layer=POLY_cond $X=6.02 $Y=1.16
+ $X2=6.15 $Y2=1.16
r281 132 140 5.77042 $w=3.5e-07 $l=3.5e-08 $layer=POLY_cond $X=5.985 $Y=1.16
+ $X2=6.02 $Y2=1.16
r282 132 138 65.1233 $w=3.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.985 $Y=1.16
+ $X2=5.59 $Y2=1.16
r283 131 132 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=5.985
+ $Y=1.17 $X2=5.985 $Y2=1.17
r284 129 137 51.8515 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.925 $Y=1.235
+ $X2=3.28 $Y2=1.235
r285 129 135 40.897 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=2.925 $Y=1.235
+ $X2=2.645 $Y2=1.235
r286 128 131 106.863 $w=3.28e-07 $l=3.06e-06 $layer=LI1_cond $X=2.925 $Y=1.17
+ $X2=5.985 $Y2=1.17
r287 128 129 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=2.925
+ $Y=1.17 $X2=2.925 $Y2=1.17
r288 126 128 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=2.36 $Y=1.17
+ $X2=2.925 $Y2=1.17
r289 125 126 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.275 $Y=1.005
+ $X2=2.36 $Y2=1.17
r290 124 125 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.275 $Y=0.795
+ $X2=2.275 $Y2=1.005
r291 123 134 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.71
+ $X2=0.71 $Y2=0.71
r292 122 124 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=0.71
+ $X2=2.275 $Y2=0.795
r293 122 123 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.19 $Y=0.71
+ $X2=0.795 $Y2=0.71
r294 118 120 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.71 $Y=1.98
+ $X2=0.71 $Y2=2.9
r295 116 118 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=0.71 $Y=0.93
+ $X2=0.71 $Y2=1.98
r296 114 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.795
+ $X2=0.71 $Y2=0.71
r297 114 116 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.71 $Y=0.795
+ $X2=0.71 $Y2=0.93
r298 110 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.625
+ $X2=0.71 $Y2=0.71
r299 110 112 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.71 $Y=0.625
+ $X2=0.71 $Y2=0.43
r300 102 103 70.8938 $w=3.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.65 $Y=1.16
+ $X2=5.08 $Y2=1.16
r301 101 102 70.8938 $w=3.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.22 $Y=1.16
+ $X2=4.65 $Y2=1.16
r302 100 101 70.8938 $w=3.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.79 $Y=1.16
+ $X2=4.22 $Y2=1.16
r303 97 98 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.515 $Y=1.41
+ $X2=1.785 $Y2=1.41
r304 95 97 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.355 $Y=1.41
+ $X2=1.515 $Y2=1.41
r305 92 94 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.19 $Y=0.985
+ $X2=9.19 $Y2=0.555
r306 91 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.835 $Y=1.06
+ $X2=8.76 $Y2=1.06
r307 90 92 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.115 $Y=1.06
+ $X2=9.19 $Y2=0.985
r308 90 91 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.115 $Y=1.06
+ $X2=8.835 $Y2=1.06
r309 87 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.76 $Y=0.985
+ $X2=8.76 $Y2=1.06
r310 87 89 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.76 $Y=0.985
+ $X2=8.76 $Y2=0.555
r311 86 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.405 $Y=1.06
+ $X2=8.33 $Y2=1.06
r312 85 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.685 $Y=1.06
+ $X2=8.76 $Y2=1.06
r313 85 86 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.685 $Y=1.06
+ $X2=8.405 $Y2=1.06
r314 82 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.33 $Y=0.985
+ $X2=8.33 $Y2=1.06
r315 82 84 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.33 $Y=0.985
+ $X2=8.33 $Y2=0.555
r316 81 107 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.975 $Y=1.06
+ $X2=7.9 $Y2=1.06
r317 80 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.255 $Y=1.06
+ $X2=8.33 $Y2=1.06
r318 80 81 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.255 $Y=1.06
+ $X2=7.975 $Y2=1.06
r319 77 107 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.9 $Y=0.985
+ $X2=7.9 $Y2=1.06
r320 77 79 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.9 $Y=0.985
+ $X2=7.9 $Y2=0.555
r321 76 106 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.545 $Y=1.06
+ $X2=7.47 $Y2=1.06
r322 75 107 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.825 $Y=1.06
+ $X2=7.9 $Y2=1.06
r323 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.825 $Y=1.06
+ $X2=7.545 $Y2=1.06
r324 72 106 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.47 $Y=0.985
+ $X2=7.47 $Y2=1.06
r325 72 74 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.47 $Y=0.985
+ $X2=7.47 $Y2=0.555
r326 71 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.115 $Y=1.06
+ $X2=7.04 $Y2=1.06
r327 70 106 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.395 $Y=1.06
+ $X2=7.47 $Y2=1.06
r328 70 71 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.395 $Y=1.06
+ $X2=7.115 $Y2=1.06
r329 67 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.04 $Y=0.985
+ $X2=7.04 $Y2=1.06
r330 67 69 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.04 $Y=0.985
+ $X2=7.04 $Y2=0.555
r331 66 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.685 $Y=1.06
+ $X2=6.61 $Y2=1.06
r332 65 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.965 $Y=1.06
+ $X2=7.04 $Y2=1.06
r333 65 66 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.965 $Y=1.06
+ $X2=6.685 $Y2=1.06
r334 62 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.61 $Y=0.985
+ $X2=6.61 $Y2=1.06
r335 62 64 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.61 $Y=0.985
+ $X2=6.61 $Y2=0.555
r336 60 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.535 $Y=1.06
+ $X2=6.61 $Y2=1.06
r337 60 141 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.535 $Y=1.06
+ $X2=6.15 $Y2=1.06
r338 57 140 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.02 $Y=0.985
+ $X2=6.02 $Y2=1.16
r339 57 59 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.02 $Y=0.985
+ $X2=6.02 $Y2=0.555
r340 54 138 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.59 $Y=0.985
+ $X2=5.59 $Y2=1.16
r341 54 56 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.59 $Y=0.985
+ $X2=5.59 $Y2=0.555
r342 53 103 12.3652 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.155 $Y=1.16
+ $X2=5.08 $Y2=1.16
r343 52 138 12.3652 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.515 $Y=1.16
+ $X2=5.59 $Y2=1.16
r344 52 53 59.3529 $w=3.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.515 $Y=1.16
+ $X2=5.155 $Y2=1.16
r345 49 103 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.08 $Y=0.985
+ $X2=5.08 $Y2=1.16
r346 49 51 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.08 $Y=0.985
+ $X2=5.08 $Y2=0.555
r347 46 102 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.65 $Y=0.985
+ $X2=4.65 $Y2=1.16
r348 46 48 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.65 $Y=0.985
+ $X2=4.65 $Y2=0.555
r349 43 101 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.22 $Y=0.985
+ $X2=4.22 $Y2=1.16
r350 43 45 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.22 $Y=0.985
+ $X2=4.22 $Y2=0.555
r351 40 100 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.79 $Y=0.985
+ $X2=3.79 $Y2=1.16
r352 40 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.79 $Y=0.985
+ $X2=3.79 $Y2=0.555
r353 39 137 10.5425 $w=3.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.355 $Y=1.16
+ $X2=3.28 $Y2=1.235
r354 38 100 12.3652 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.715 $Y=1.16
+ $X2=3.79 $Y2=1.16
r355 38 39 59.3529 $w=3.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.715 $Y=1.16
+ $X2=3.355 $Y2=1.16
r356 35 137 21.2229 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.28 $Y=0.985
+ $X2=3.28 $Y2=1.235
r357 35 37 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.28 $Y=0.985
+ $X2=3.28 $Y2=0.555
r358 31 135 21.2229 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.645 $Y=1.485
+ $X2=2.645 $Y2=1.235
r359 31 33 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.645 $Y=1.485
+ $X2=2.645 $Y2=2.465
r360 30 99 12.05 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.29 $Y=1.41
+ $X2=2.195 $Y2=1.41
r361 29 135 25.4547 $w=3.3e-07 $l=2.09165e-07 $layer=POLY_cond $X=2.57 $Y=1.41
+ $X2=2.645 $Y2=1.235
r362 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.57 $Y=1.41
+ $X2=2.29 $Y2=1.41
r363 25 99 12.05 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.215 $Y=1.485
+ $X2=2.195 $Y2=1.41
r364 25 27 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.215 $Y=1.485
+ $X2=2.215 $Y2=2.465
r365 21 99 12.05 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.175 $Y=1.335
+ $X2=2.195 $Y2=1.41
r366 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.175 $Y=1.335
+ $X2=2.175 $Y2=0.655
r367 20 98 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.86 $Y=1.41
+ $X2=1.785 $Y2=1.41
r368 19 99 12.05 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.1 $Y=1.41 $X2=2.195
+ $Y2=1.41
r369 19 20 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.1 $Y=1.41
+ $X2=1.86 $Y2=1.41
r370 15 98 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.785 $Y=1.485
+ $X2=1.785 $Y2=1.41
r371 15 17 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.785 $Y=1.485
+ $X2=1.785 $Y2=2.465
r372 11 97 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.515 $Y=1.335
+ $X2=1.515 $Y2=1.41
r373 11 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.515 $Y=1.335
+ $X2=1.515 $Y2=0.655
r374 7 95 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.355 $Y=1.485
+ $X2=1.355 $Y2=1.41
r375 7 9 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.355 $Y=1.485
+ $X2=1.355 $Y2=2.465
r376 2 120 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.9
r377 2 118 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=1.98
r378 1 116 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.93
r379 1 112 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_286_367# 1 2 3 10 12 13 14 15 17 18
+ 20 22 23 25 27 28 30 32 33 35 37 38 40 42 43 45 47 48 50 52 53 55 56 58 59 61
+ 62 64 65 67 68 70 71 73 74 76 77 78 79 81 82 84 86 87 89 91 92 93 94 95 96 97
+ 98 99 100 103 107 109 110 113 117 119 126 134
c329 134 0 1.023e-19 $X=6.39 $Y=1.515
c330 110 0 2.49061e-19 $X=2.01 $Y=1.9
c331 109 0 1.19111e-20 $X=2.265 $Y=1.9
c332 84 0 4.06089e-20 $X=10.835 $Y=1.725
r333 142 143 57.0964 $w=3.63e-07 $l=4.3e-07 $layer=POLY_cond $X=9.115 $Y=1.535
+ $X2=9.545 $Y2=1.535
r334 141 142 57.0964 $w=3.63e-07 $l=4.3e-07 $layer=POLY_cond $X=8.685 $Y=1.535
+ $X2=9.115 $Y2=1.535
r335 140 141 57.0964 $w=3.63e-07 $l=4.3e-07 $layer=POLY_cond $X=8.255 $Y=1.535
+ $X2=8.685 $Y2=1.535
r336 139 140 59.7521 $w=3.63e-07 $l=4.5e-07 $layer=POLY_cond $X=7.805 $Y=1.535
+ $X2=8.255 $Y2=1.535
r337 138 139 57.0964 $w=3.63e-07 $l=4.3e-07 $layer=POLY_cond $X=7.375 $Y=1.535
+ $X2=7.805 $Y2=1.535
r338 137 138 57.0964 $w=3.63e-07 $l=4.3e-07 $layer=POLY_cond $X=6.945 $Y=1.535
+ $X2=7.375 $Y2=1.535
r339 133 137 51.7851 $w=3.63e-07 $l=3.9e-07 $layer=POLY_cond $X=6.555 $Y=1.535
+ $X2=6.945 $Y2=1.535
r340 133 135 5.31129 $w=3.63e-07 $l=4e-08 $layer=POLY_cond $X=6.555 $Y=1.535
+ $X2=6.515 $Y2=1.535
r341 132 134 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=1.515
+ $X2=6.39 $Y2=1.515
r342 132 133 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=6.555
+ $Y=1.51 $X2=6.555 $Y2=1.51
r343 128 130 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.43 $Y=1.9 $X2=2.43
+ $Y2=1.98
r344 126 128 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.43 $Y=1.6
+ $X2=2.43 $Y2=1.9
r345 120 143 9.29477 $w=3.63e-07 $l=7e-08 $layer=POLY_cond $X=9.615 $Y=1.535
+ $X2=9.545 $Y2=1.535
r346 119 120 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=9.615
+ $Y=1.51 $X2=9.615 $Y2=1.51
r347 117 132 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=6.56 $Y=1.515
+ $X2=6.555 $Y2=1.515
r348 117 119 103.55 $w=3.38e-07 $l=3.055e-06 $layer=LI1_cond $X=6.56 $Y=1.515
+ $X2=9.615 $Y2=1.515
r349 116 126 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=1.6
+ $X2=2.43 $Y2=1.6
r350 116 134 247.588 $w=1.68e-07 $l=3.795e-06 $layer=LI1_cond $X=2.595 $Y=1.6
+ $X2=6.39 $Y2=1.6
r351 111 130 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.43 $Y=1.985
+ $X2=2.43 $Y2=1.98
r352 111 113 31.9541 $w=3.28e-07 $l=9.15e-07 $layer=LI1_cond $X=2.43 $Y=1.985
+ $X2=2.43 $Y2=2.9
r353 109 128 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.9
+ $X2=2.43 $Y2=1.9
r354 109 110 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.265 $Y=1.9
+ $X2=2.01 $Y2=1.9
r355 105 110 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=1.9
+ $X2=2.01 $Y2=1.9
r356 105 123 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.845 $Y=1.9
+ $X2=1.57 $Y2=1.9
r357 105 107 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=1.845 $Y=1.815
+ $X2=1.845 $Y2=1.06
r358 103 123 31.9541 $w=3.28e-07 $l=9.15e-07 $layer=LI1_cond $X=1.57 $Y=2.9
+ $X2=1.57 $Y2=1.985
r359 89 91 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=11.265 $Y=1.725
+ $X2=11.265 $Y2=2.465
r360 88 100 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.91 $Y=1.65
+ $X2=10.835 $Y2=1.65
r361 87 89 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.19 $Y=1.65
+ $X2=11.265 $Y2=1.725
r362 87 88 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=11.19 $Y=1.65
+ $X2=10.91 $Y2=1.65
r363 84 100 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.835 $Y=1.725
+ $X2=10.835 $Y2=1.65
r364 84 86 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=10.835 $Y=1.725
+ $X2=10.835 $Y2=2.465
r365 83 99 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.48 $Y=1.65
+ $X2=10.405 $Y2=1.65
r366 82 100 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.76 $Y=1.65
+ $X2=10.835 $Y2=1.65
r367 82 83 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.76 $Y=1.65
+ $X2=10.48 $Y2=1.65
r368 79 99 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.405 $Y=1.725
+ $X2=10.405 $Y2=1.65
r369 79 81 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=10.405 $Y=1.725
+ $X2=10.405 $Y2=2.465
r370 77 99 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.33 $Y=1.65
+ $X2=10.405 $Y2=1.65
r371 77 78 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.33 $Y=1.65
+ $X2=10.05 $Y2=1.65
r372 74 78 27.0016 $w=3.63e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.975 $Y=1.725
+ $X2=10.05 $Y2=1.65
r373 74 120 47.8017 $w=3.63e-07 $l=4.44972e-07 $layer=POLY_cond $X=9.975
+ $Y=1.725 $X2=9.615 $Y2=1.535
r374 74 76 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.975 $Y=1.725
+ $X2=9.975 $Y2=2.465
r375 71 143 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.545 $Y=1.725
+ $X2=9.545 $Y2=1.535
r376 71 73 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.545 $Y=1.725
+ $X2=9.545 $Y2=2.465
r377 68 142 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.115 $Y=1.725
+ $X2=9.115 $Y2=1.535
r378 68 70 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.115 $Y=1.725
+ $X2=9.115 $Y2=2.465
r379 65 141 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.685 $Y=1.725
+ $X2=8.685 $Y2=1.535
r380 65 67 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.685 $Y=1.725
+ $X2=8.685 $Y2=2.465
r381 62 140 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.255 $Y=1.725
+ $X2=8.255 $Y2=1.535
r382 62 64 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.255 $Y=1.725
+ $X2=8.255 $Y2=2.465
r383 59 139 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.805 $Y=1.725
+ $X2=7.805 $Y2=1.535
r384 59 61 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.805 $Y=1.725
+ $X2=7.805 $Y2=2.465
r385 56 138 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.375 $Y=1.725
+ $X2=7.375 $Y2=1.535
r386 56 58 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.375 $Y=1.725
+ $X2=7.375 $Y2=2.465
r387 53 137 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.945 $Y=1.725
+ $X2=6.945 $Y2=1.535
r388 53 55 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.945 $Y=1.725
+ $X2=6.945 $Y2=2.465
r389 50 135 23.5056 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.515 $Y=1.725
+ $X2=6.515 $Y2=1.535
r390 50 52 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.515 $Y=1.725
+ $X2=6.515 $Y2=2.465
r391 49 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.16 $Y=1.65
+ $X2=6.085 $Y2=1.65
r392 48 135 33.6407 $w=3.63e-07 $l=1.73205e-07 $layer=POLY_cond $X=6.39 $Y=1.65
+ $X2=6.515 $Y2=1.535
r393 48 49 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.39 $Y=1.65
+ $X2=6.16 $Y2=1.65
r394 45 98 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=1.725
+ $X2=6.085 $Y2=1.65
r395 45 47 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.085 $Y=1.725
+ $X2=6.085 $Y2=2.465
r396 44 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.73 $Y=1.65
+ $X2=5.655 $Y2=1.65
r397 43 98 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.01 $Y=1.65
+ $X2=6.085 $Y2=1.65
r398 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.01 $Y=1.65
+ $X2=5.73 $Y2=1.65
r399 40 97 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.655 $Y=1.725
+ $X2=5.655 $Y2=1.65
r400 40 42 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.655 $Y=1.725
+ $X2=5.655 $Y2=2.465
r401 39 96 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.3 $Y=1.65
+ $X2=5.225 $Y2=1.65
r402 38 97 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.58 $Y=1.65
+ $X2=5.655 $Y2=1.65
r403 38 39 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.58 $Y=1.65
+ $X2=5.3 $Y2=1.65
r404 35 96 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.225 $Y=1.725
+ $X2=5.225 $Y2=1.65
r405 35 37 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.225 $Y=1.725
+ $X2=5.225 $Y2=2.465
r406 34 95 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.87 $Y=1.65
+ $X2=4.795 $Y2=1.65
r407 33 96 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.15 $Y=1.65
+ $X2=5.225 $Y2=1.65
r408 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.15 $Y=1.65
+ $X2=4.87 $Y2=1.65
r409 30 95 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.795 $Y=1.725
+ $X2=4.795 $Y2=1.65
r410 30 32 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.795 $Y=1.725
+ $X2=4.795 $Y2=2.465
r411 29 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.44 $Y=1.65
+ $X2=4.365 $Y2=1.65
r412 28 95 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.72 $Y=1.65
+ $X2=4.795 $Y2=1.65
r413 28 29 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.72 $Y=1.65
+ $X2=4.44 $Y2=1.65
r414 25 94 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.365 $Y=1.725
+ $X2=4.365 $Y2=1.65
r415 25 27 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.365 $Y=1.725
+ $X2=4.365 $Y2=2.465
r416 24 93 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.01 $Y=1.65
+ $X2=3.935 $Y2=1.65
r417 23 94 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=1.65
+ $X2=4.365 $Y2=1.65
r418 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.29 $Y=1.65
+ $X2=4.01 $Y2=1.65
r419 20 93 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.935 $Y=1.725
+ $X2=3.935 $Y2=1.65
r420 20 22 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.935 $Y=1.725
+ $X2=3.935 $Y2=2.465
r421 19 92 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.58 $Y=1.65
+ $X2=3.505 $Y2=1.65
r422 18 93 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.86 $Y=1.65
+ $X2=3.935 $Y2=1.65
r423 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.86 $Y=1.65
+ $X2=3.58 $Y2=1.65
r424 15 92 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=1.725
+ $X2=3.505 $Y2=1.65
r425 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.505 $Y=1.725
+ $X2=3.505 $Y2=2.465
r426 13 92 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.43 $Y=1.65
+ $X2=3.505 $Y2=1.65
r427 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.43 $Y=1.65
+ $X2=3.15 $Y2=1.65
r428 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.075 $Y=1.725
+ $X2=3.15 $Y2=1.65
r429 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.075 $Y=1.725
+ $X2=3.075 $Y2=2.465
r430 3 130 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=1.98
r431 3 113 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=2.9
r432 2 123 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=1.98
r433 2 103 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.9
r434 1 107 182 $w=1.7e-07 $l=9.43928e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.235 $X2=1.845 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_1909_21# 1 2 3 4 5 6 19 21 22 23 24
+ 26 27 29 31 32 34 36 37 39 41 42 44 46 49 51 53 56 58 60 63 65 67 70 72 74 77
+ 79 81 84 86 88 91 93 95 98 100 102 105 109 113 117 121 125 129 133 137 141 145
+ 149 151 152 153 154 155 163 170 172 175 179 181 185 189 193 195 199 203 207
+ 211 215 216 217 218 219 220
c446 170 0 1.20079e-19 $X=21.265 $Y=1.15
r447 249 250 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=18.29 $Y=1.155
+ $X2=18.72 $Y2=1.155
r448 248 249 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=17.86 $Y=1.155
+ $X2=18.29 $Y2=1.155
r449 247 248 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=17.43 $Y=1.155
+ $X2=17.86 $Y2=1.155
r450 246 247 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=17 $Y=1.155
+ $X2=17.43 $Y2=1.155
r451 245 246 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=16.57 $Y=1.155
+ $X2=17 $Y2=1.155
r452 244 245 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=16.14 $Y=1.155
+ $X2=16.57 $Y2=1.155
r453 241 242 37.747 $w=3.32e-07 $l=2.6e-07 $layer=POLY_cond $X=15.45 $Y=1.155
+ $X2=15.71 $Y2=1.155
r454 238 239 37.747 $w=3.32e-07 $l=2.6e-07 $layer=POLY_cond $X=15.02 $Y=1.155
+ $X2=15.28 $Y2=1.155
r455 237 238 24.6807 $w=3.32e-07 $l=1.7e-07 $layer=POLY_cond $X=14.85 $Y=1.155
+ $X2=15.02 $Y2=1.155
r456 236 237 37.747 $w=3.32e-07 $l=2.6e-07 $layer=POLY_cond $X=14.59 $Y=1.155
+ $X2=14.85 $Y2=1.155
r457 235 236 24.6807 $w=3.32e-07 $l=1.7e-07 $layer=POLY_cond $X=14.42 $Y=1.155
+ $X2=14.59 $Y2=1.155
r458 234 235 37.747 $w=3.32e-07 $l=2.6e-07 $layer=POLY_cond $X=14.16 $Y=1.155
+ $X2=14.42 $Y2=1.155
r459 233 234 24.6807 $w=3.32e-07 $l=1.7e-07 $layer=POLY_cond $X=13.99 $Y=1.155
+ $X2=14.16 $Y2=1.155
r460 232 233 37.747 $w=3.32e-07 $l=2.6e-07 $layer=POLY_cond $X=13.73 $Y=1.155
+ $X2=13.99 $Y2=1.155
r461 231 232 24.6807 $w=3.32e-07 $l=1.7e-07 $layer=POLY_cond $X=13.56 $Y=1.155
+ $X2=13.73 $Y2=1.155
r462 230 231 37.747 $w=3.32e-07 $l=2.6e-07 $layer=POLY_cond $X=13.3 $Y=1.155
+ $X2=13.56 $Y2=1.155
r463 229 230 24.6807 $w=3.32e-07 $l=1.7e-07 $layer=POLY_cond $X=13.13 $Y=1.155
+ $X2=13.3 $Y2=1.155
r464 228 229 37.747 $w=3.32e-07 $l=2.6e-07 $layer=POLY_cond $X=12.87 $Y=1.155
+ $X2=13.13 $Y2=1.155
r465 227 228 24.6807 $w=3.32e-07 $l=1.7e-07 $layer=POLY_cond $X=12.7 $Y=1.155
+ $X2=12.87 $Y2=1.155
r466 211 213 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=24.25 $Y=1.98
+ $X2=24.25 $Y2=2.9
r467 209 211 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=24.25 $Y=1.865
+ $X2=24.25 $Y2=1.98
r468 208 219 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.53 $Y=1.78
+ $X2=23.365 $Y2=1.78
r469 207 209 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=24.085 $Y=1.78
+ $X2=24.25 $Y2=1.865
r470 207 208 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=24.085 $Y=1.78
+ $X2=23.53 $Y2=1.78
r471 203 205 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=23.365 $Y=1.98
+ $X2=23.365 $Y2=2.9
r472 201 219 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=23.365 $Y=1.865
+ $X2=23.365 $Y2=1.78
r473 201 203 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=23.365 $Y=1.865
+ $X2=23.365 $Y2=1.98
r474 197 199 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=23.215 $Y=0.83
+ $X2=23.215 $Y2=0.43
r475 196 218 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.67 $Y=1.78
+ $X2=22.505 $Y2=1.78
r476 195 219 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.2 $Y=1.78
+ $X2=23.365 $Y2=1.78
r477 195 196 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=23.2 $Y=1.78
+ $X2=22.67 $Y2=1.78
r478 194 217 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.36 $Y=0.915
+ $X2=22.195 $Y2=0.915
r479 193 197 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=23.05 $Y=0.915
+ $X2=23.215 $Y2=0.83
r480 193 194 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=23.05 $Y=0.915
+ $X2=22.36 $Y2=0.915
r481 189 191 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=22.505 $Y=1.98
+ $X2=22.505 $Y2=2.9
r482 187 218 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=22.505 $Y=1.865
+ $X2=22.505 $Y2=1.78
r483 187 189 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=22.505 $Y=1.865
+ $X2=22.505 $Y2=1.98
r484 183 217 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=22.195 $Y=0.83
+ $X2=22.195 $Y2=0.915
r485 183 185 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=22.195 $Y=0.83
+ $X2=22.195 $Y2=0.38
r486 182 216 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=21.81 $Y=1.78
+ $X2=21.645 $Y2=1.78
r487 181 218 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.34 $Y=1.78
+ $X2=22.505 $Y2=1.78
r488 181 182 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=22.34 $Y=1.78
+ $X2=21.81 $Y2=1.78
r489 180 215 3.70735 $w=2.5e-07 $l=1.94921e-07 $layer=LI1_cond $X=21.65 $Y=0.915
+ $X2=21.565 $Y2=1.072
r490 179 217 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.03 $Y=0.915
+ $X2=22.195 $Y2=0.915
r491 179 180 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=22.03 $Y=0.915
+ $X2=21.65 $Y2=0.915
r492 175 177 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=21.645 $Y=1.98
+ $X2=21.645 $Y2=2.9
r493 173 216 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=21.645 $Y=1.865
+ $X2=21.645 $Y2=1.78
r494 173 175 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=21.645 $Y=1.865
+ $X2=21.645 $Y2=1.98
r495 172 216 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=21.565
+ $Y=1.695 $X2=21.645 $Y2=1.78
r496 171 215 2.76166 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=21.565 $Y=1.315
+ $X2=21.565 $Y2=1.072
r497 171 172 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=21.565 $Y=1.315
+ $X2=21.565 $Y2=1.695
r498 170 220 131.146 $w=3.3e-07 $l=7.5e-07 $layer=POLY_cond $X=21.265 $Y=1.15
+ $X2=20.515 $Y2=1.15
r499 169 170 17.0918 $w=1.7e-07 $l=1.445e-06 $layer=licon1_POLY $count=8
+ $X=21.265 $Y=1.15 $X2=21.265 $Y2=1.15
r500 167 244 45.7319 $w=3.32e-07 $l=3.15e-07 $layer=POLY_cond $X=15.825 $Y=1.155
+ $X2=16.14 $Y2=1.155
r501 167 242 16.6958 $w=3.32e-07 $l=1.15e-07 $layer=POLY_cond $X=15.825 $Y=1.155
+ $X2=15.71 $Y2=1.155
r502 166 169 189.978 $w=3.28e-07 $l=5.44e-06 $layer=LI1_cond $X=15.825 $Y=1.15
+ $X2=21.265 $Y2=1.15
r503 166 167 17.0918 $w=1.7e-07 $l=1.445e-06 $layer=licon1_POLY $count=8
+ $X=15.825 $Y=1.15 $X2=15.825 $Y2=1.15
r504 163 215 3.70735 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=21.48 $Y=1.15
+ $X2=21.565 $Y2=1.072
r505 163 169 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=21.48 $Y=1.15
+ $X2=21.265 $Y2=1.15
r506 162 241 23.2289 $w=3.32e-07 $l=1.6e-07 $layer=POLY_cond $X=15.29 $Y=1.155
+ $X2=15.45 $Y2=1.155
r507 162 239 1.45181 $w=3.32e-07 $l=1e-08 $layer=POLY_cond $X=15.29 $Y=1.155
+ $X2=15.28 $Y2=1.155
r508 161 162 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=15.29
+ $Y=1.16 $X2=15.29 $Y2=1.16
r509 158 227 18.8735 $w=3.32e-07 $l=1.3e-07 $layer=POLY_cond $X=12.57 $Y=1.155
+ $X2=12.7 $Y2=1.155
r510 158 225 18.8735 $w=3.32e-07 $l=1.3e-07 $layer=POLY_cond $X=12.57 $Y=1.155
+ $X2=12.44 $Y2=1.155
r511 157 161 125.386 $w=2.48e-07 $l=2.72e-06 $layer=LI1_cond $X=12.57 $Y=1.2
+ $X2=15.29 $Y2=1.2
r512 157 158 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=12.57
+ $Y=1.16 $X2=12.57 $Y2=1.16
r513 155 166 22.2022 $w=2.72e-07 $l=5.19399e-07 $layer=LI1_cond $X=15.33 $Y=1.2
+ $X2=15.825 $Y2=1.15
r514 155 161 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=15.33 $Y=1.2
+ $X2=15.29 $Y2=1.2
r515 147 220 10.8886 $w=3.32e-07 $l=7.74597e-08 $layer=POLY_cond $X=20.44
+ $Y=1.155 $X2=20.515 $Y2=1.15
r516 147 149 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=20.44 $Y=1.315
+ $X2=20.44 $Y2=2.155
r517 143 147 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=20.01 $Y=1.155
+ $X2=20.44 $Y2=1.155
r518 143 145 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=20.01 $Y=1.315
+ $X2=20.01 $Y2=2.155
r519 139 143 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=19.58 $Y=1.155
+ $X2=20.01 $Y2=1.155
r520 139 141 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=19.58 $Y=1.315
+ $X2=19.58 $Y2=2.155
r521 135 139 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=19.15 $Y=1.155
+ $X2=19.58 $Y2=1.155
r522 135 250 62.4277 $w=3.32e-07 $l=4.3e-07 $layer=POLY_cond $X=19.15 $Y=1.155
+ $X2=18.72 $Y2=1.155
r523 135 137 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=19.15 $Y=1.315
+ $X2=19.15 $Y2=2.155
r524 131 250 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=18.72 $Y=1.325
+ $X2=18.72 $Y2=1.155
r525 131 133 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=18.72 $Y=1.325
+ $X2=18.72 $Y2=2.155
r526 127 249 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=18.29 $Y=1.325
+ $X2=18.29 $Y2=1.155
r527 127 129 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=18.29 $Y=1.325
+ $X2=18.29 $Y2=2.155
r528 123 248 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=17.86 $Y=1.325
+ $X2=17.86 $Y2=1.155
r529 123 125 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=17.86 $Y=1.325
+ $X2=17.86 $Y2=2.155
r530 119 247 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=17.43 $Y=1.325
+ $X2=17.43 $Y2=1.155
r531 119 121 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=17.43 $Y=1.325
+ $X2=17.43 $Y2=2.155
r532 115 246 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=17 $Y=1.325
+ $X2=17 $Y2=1.155
r533 115 117 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=17 $Y=1.325
+ $X2=17 $Y2=2.155
r534 111 245 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=16.57 $Y=1.325
+ $X2=16.57 $Y2=1.155
r535 111 113 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=16.57 $Y=1.325
+ $X2=16.57 $Y2=2.155
r536 107 244 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=16.14 $Y=1.325
+ $X2=16.14 $Y2=1.155
r537 107 109 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=16.14 $Y=1.325
+ $X2=16.14 $Y2=2.155
r538 103 242 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=15.71 $Y=1.325
+ $X2=15.71 $Y2=1.155
r539 103 105 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=15.71 $Y=1.325
+ $X2=15.71 $Y2=2.155
r540 100 241 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=15.45 $Y=0.985
+ $X2=15.45 $Y2=1.155
r541 100 102 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=15.45 $Y=0.985
+ $X2=15.45 $Y2=0.555
r542 96 239 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=15.28 $Y=1.325
+ $X2=15.28 $Y2=1.155
r543 96 98 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=15.28 $Y=1.325
+ $X2=15.28 $Y2=2.155
r544 93 238 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=15.02 $Y=0.985
+ $X2=15.02 $Y2=1.155
r545 93 95 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=15.02 $Y=0.985
+ $X2=15.02 $Y2=0.555
r546 89 237 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=14.85 $Y=1.325
+ $X2=14.85 $Y2=1.155
r547 89 91 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=14.85 $Y=1.325
+ $X2=14.85 $Y2=2.155
r548 86 236 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=14.59 $Y=0.985
+ $X2=14.59 $Y2=1.155
r549 86 88 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=14.59 $Y=0.985
+ $X2=14.59 $Y2=0.555
r550 82 235 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=14.42 $Y=1.325
+ $X2=14.42 $Y2=1.155
r551 82 84 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=14.42 $Y=1.325
+ $X2=14.42 $Y2=2.155
r552 79 234 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=14.16 $Y=0.985
+ $X2=14.16 $Y2=1.155
r553 79 81 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=14.16 $Y=0.985
+ $X2=14.16 $Y2=0.555
r554 75 233 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=13.99 $Y=1.325
+ $X2=13.99 $Y2=1.155
r555 75 77 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=13.99 $Y=1.325
+ $X2=13.99 $Y2=2.155
r556 72 232 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=13.73 $Y=0.985
+ $X2=13.73 $Y2=1.155
r557 72 74 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.73 $Y=0.985
+ $X2=13.73 $Y2=0.555
r558 68 231 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=13.56 $Y=1.325
+ $X2=13.56 $Y2=1.155
r559 68 70 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=13.56 $Y=1.325
+ $X2=13.56 $Y2=2.155
r560 65 230 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=13.3 $Y=0.985
+ $X2=13.3 $Y2=1.155
r561 65 67 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.3 $Y=0.985
+ $X2=13.3 $Y2=0.555
r562 61 229 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=13.13 $Y=1.325
+ $X2=13.13 $Y2=1.155
r563 61 63 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=13.13 $Y=1.325
+ $X2=13.13 $Y2=2.155
r564 58 228 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.87 $Y=0.985
+ $X2=12.87 $Y2=1.155
r565 58 60 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.87 $Y=0.985
+ $X2=12.87 $Y2=0.555
r566 54 227 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.7 $Y=1.325
+ $X2=12.7 $Y2=1.155
r567 54 56 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=12.7 $Y=1.325
+ $X2=12.7 $Y2=2.155
r568 51 225 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.44 $Y=0.985
+ $X2=12.44 $Y2=1.155
r569 51 53 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.44 $Y=0.985
+ $X2=12.44 $Y2=0.555
r570 47 225 24.6807 $w=3.32e-07 $l=2.40416e-07 $layer=POLY_cond $X=12.27
+ $Y=1.325 $X2=12.44 $Y2=1.155
r571 47 223 37.747 $w=3.32e-07 $l=3.34365e-07 $layer=POLY_cond $X=12.27 $Y=1.325
+ $X2=12.01 $Y2=1.155
r572 47 49 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=12.27 $Y=1.325
+ $X2=12.27 $Y2=2.155
r573 44 223 21.3668 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.01 $Y=0.985
+ $X2=12.01 $Y2=1.155
r574 44 46 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.01 $Y=0.985
+ $X2=12.01 $Y2=0.555
r575 43 154 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.655 $Y=1.06
+ $X2=11.58 $Y2=1.06
r576 42 223 25.5476 $w=3.32e-07 $l=1.27083e-07 $layer=POLY_cond $X=11.935
+ $Y=1.06 $X2=12.01 $Y2=1.155
r577 42 43 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=11.935 $Y=1.06
+ $X2=11.655 $Y2=1.06
r578 39 154 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.58 $Y=0.985
+ $X2=11.58 $Y2=1.06
r579 39 41 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.58 $Y=0.985
+ $X2=11.58 $Y2=0.555
r580 38 153 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.225 $Y=1.06
+ $X2=11.15 $Y2=1.06
r581 37 154 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.505 $Y=1.06
+ $X2=11.58 $Y2=1.06
r582 37 38 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=11.505 $Y=1.06
+ $X2=11.225 $Y2=1.06
r583 34 153 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.15 $Y=0.985
+ $X2=11.15 $Y2=1.06
r584 34 36 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.15 $Y=0.985
+ $X2=11.15 $Y2=0.555
r585 33 152 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=1.06
+ $X2=10.64 $Y2=1.06
r586 32 153 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.075 $Y=1.06
+ $X2=11.15 $Y2=1.06
r587 32 33 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=11.075 $Y=1.06
+ $X2=10.715 $Y2=1.06
r588 29 152 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.64 $Y=0.985
+ $X2=10.64 $Y2=1.06
r589 29 31 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.64 $Y=0.985
+ $X2=10.64 $Y2=0.555
r590 28 151 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.205 $Y=1.06
+ $X2=10.13 $Y2=1.06
r591 27 152 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.565 $Y=1.06
+ $X2=10.64 $Y2=1.06
r592 27 28 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.565 $Y=1.06
+ $X2=10.205 $Y2=1.06
r593 24 151 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.13 $Y=0.985
+ $X2=10.13 $Y2=1.06
r594 24 26 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.13 $Y=0.985
+ $X2=10.13 $Y2=0.555
r595 22 151 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.055 $Y=1.06
+ $X2=10.13 $Y2=1.06
r596 22 23 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.055 $Y=1.06
+ $X2=9.695 $Y2=1.06
r597 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.62 $Y=0.985
+ $X2=9.695 $Y2=1.06
r598 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.62 $Y=0.985
+ $X2=9.62 $Y2=0.555
r599 6 213 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=24.11
+ $Y=1.835 $X2=24.25 $Y2=2.9
r600 6 211 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=24.11
+ $Y=1.835 $X2=24.25 $Y2=1.98
r601 5 205 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=23.225
+ $Y=1.835 $X2=23.365 $Y2=2.9
r602 5 203 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=23.225
+ $Y=1.835 $X2=23.365 $Y2=1.98
r603 4 191 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=22.365
+ $Y=1.835 $X2=22.505 $Y2=2.9
r604 4 189 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=22.365
+ $Y=1.835 $X2=22.505 $Y2=1.98
r605 3 177 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=21.505
+ $Y=1.835 $X2=21.645 $Y2=2.9
r606 3 175 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=21.505
+ $Y=1.835 $X2=21.645 $Y2=1.98
r607 2 199 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=23.075
+ $Y=0.235 $X2=23.215 $Y2=0.43
r608 1 185 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=21.98
+ $Y=0.235 $X2=22.195 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A 3 5 6 9 11 13 16 18 20 23 25 27 30
+ 32 34 37 41 45 47 48 49 50 51 52 82
c133 52 0 1.20079e-19 $X=24.72 $Y=1.295
r134 82 83 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=24.375
+ $Y=1.35 $X2=24.375 $Y2=1.35
r135 73 75 10.727 $w=3.37e-07 $l=7.5e-08 $layer=POLY_cond $X=23.355 $Y=1.445
+ $X2=23.43 $Y2=1.445
r136 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.675
+ $Y=1.35 $X2=22.675 $Y2=1.35
r137 65 67 37.9021 $w=3.37e-07 $l=2.65e-07 $layer=POLY_cond $X=22.41 $Y=1.445
+ $X2=22.675 $Y2=1.445
r138 63 65 10.727 $w=3.37e-07 $l=7.5e-08 $layer=POLY_cond $X=22.335 $Y=1.445
+ $X2=22.41 $Y2=1.445
r139 59 60 6.4362 $w=3.37e-07 $l=4.5e-08 $layer=POLY_cond $X=21.86 $Y=1.445
+ $X2=21.905 $Y2=1.445
r140 52 83 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=24.72 $Y=1.347
+ $X2=24.375 $Y2=1.347
r141 51 83 4.64417 $w=3.33e-07 $l=1.35e-07 $layer=LI1_cond $X=24.24 $Y=1.347
+ $X2=24.375 $Y2=1.347
r142 50 51 18.7487 $w=3.33e-07 $l=5.45e-07 $layer=LI1_cond $X=23.695 $Y=1.347
+ $X2=24.24 $Y2=1.347
r143 50 78 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=23.695
+ $Y=1.35 $X2=23.695 $Y2=1.35
r144 49 50 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=23.28 $Y=1.347
+ $X2=23.695 $Y2=1.347
r145 49 73 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=23.355
+ $Y=1.35 $X2=23.355 $Y2=1.35
r146 48 49 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=22.8 $Y=1.347
+ $X2=23.28 $Y2=1.347
r147 48 68 4.30016 $w=3.33e-07 $l=1.25e-07 $layer=LI1_cond $X=22.8 $Y=1.347
+ $X2=22.675 $Y2=1.347
r148 47 68 12.2125 $w=3.33e-07 $l=3.55e-07 $layer=LI1_cond $X=22.32 $Y=1.347
+ $X2=22.675 $Y2=1.347
r149 47 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=22.335
+ $Y=1.35 $X2=22.335 $Y2=1.35
r150 43 82 12.8724 $w=3.37e-07 $l=9e-08 $layer=POLY_cond $X=24.465 $Y=1.445
+ $X2=24.375 $Y2=1.445
r151 43 45 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=24.465 $Y=1.515
+ $X2=24.465 $Y2=2.465
r152 39 82 48.6291 $w=3.37e-07 $l=3.4e-07 $layer=POLY_cond $X=24.035 $Y=1.445
+ $X2=24.375 $Y2=1.445
r153 39 78 48.6291 $w=3.37e-07 $l=3.4e-07 $layer=POLY_cond $X=24.035 $Y=1.445
+ $X2=23.695 $Y2=1.445
r154 39 41 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=24.035 $Y=1.515
+ $X2=24.035 $Y2=2.465
r155 35 78 16.4481 $w=3.37e-07 $l=1.15e-07 $layer=POLY_cond $X=23.58 $Y=1.445
+ $X2=23.695 $Y2=1.445
r156 35 75 21.454 $w=3.37e-07 $l=1.5e-07 $layer=POLY_cond $X=23.58 $Y=1.445
+ $X2=23.43 $Y2=1.445
r157 35 37 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=23.58 $Y=1.515
+ $X2=23.58 $Y2=2.465
r158 32 75 21.7231 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=23.43 $Y=1.185
+ $X2=23.43 $Y2=1.445
r159 32 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=23.43 $Y=1.185
+ $X2=23.43 $Y2=0.655
r160 28 73 29.3205 $w=3.37e-07 $l=2.05e-07 $layer=POLY_cond $X=23.15 $Y=1.445
+ $X2=23.355 $Y2=1.445
r161 28 70 21.454 $w=3.37e-07 $l=1.5e-07 $layer=POLY_cond $X=23.15 $Y=1.445
+ $X2=23 $Y2=1.445
r162 28 30 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=23.15 $Y=1.515
+ $X2=23.15 $Y2=2.465
r163 25 70 21.7231 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=23 $Y=1.185 $X2=23
+ $Y2=1.445
r164 25 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=23 $Y=1.185 $X2=23
+ $Y2=0.655
r165 21 70 40.0475 $w=3.37e-07 $l=2.8e-07 $layer=POLY_cond $X=22.72 $Y=1.445
+ $X2=23 $Y2=1.445
r166 21 67 6.4362 $w=3.37e-07 $l=4.5e-08 $layer=POLY_cond $X=22.72 $Y=1.445
+ $X2=22.675 $Y2=1.445
r167 21 23 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=22.72 $Y=1.515
+ $X2=22.72 $Y2=2.465
r168 18 65 21.7231 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=22.41 $Y=1.185
+ $X2=22.41 $Y2=1.445
r169 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=22.41 $Y=1.185
+ $X2=22.41 $Y2=0.655
r170 14 63 6.4362 $w=3.37e-07 $l=4.5e-08 $layer=POLY_cond $X=22.29 $Y=1.445
+ $X2=22.335 $Y2=1.445
r171 14 60 55.0653 $w=3.37e-07 $l=3.85e-07 $layer=POLY_cond $X=22.29 $Y=1.445
+ $X2=21.905 $Y2=1.445
r172 14 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=22.29 $Y=1.515
+ $X2=22.29 $Y2=2.465
r173 11 60 21.7231 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=21.905 $Y=1.185
+ $X2=21.905 $Y2=1.445
r174 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=21.905 $Y=1.185
+ $X2=21.905 $Y2=0.655
r175 7 59 21.7231 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=21.86 $Y=1.705
+ $X2=21.86 $Y2=1.445
r176 7 9 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=21.86 $Y=1.705
+ $X2=21.86 $Y2=2.465
r177 5 59 25.7805 $w=3.37e-07 $l=2.19317e-07 $layer=POLY_cond $X=21.785 $Y=1.63
+ $X2=21.86 $Y2=1.445
r178 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=21.785 $Y=1.63
+ $X2=21.505 $Y2=1.63
r179 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.43 $Y=1.705
+ $X2=21.505 $Y2=1.63
r180 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=21.43 $Y=1.705
+ $X2=21.43 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 58 60 66 72 76 82 84 88 92 96 100 104 106 110 114 118 124 128
+ 134 138 142 146 150 152 157 158 160 161 163 164 165 166 168 169 171 172 174
+ 175 176 177 179 180 182 183 185 186 188 189 191 192 193 194 195 245 254 257
+ 260 264
r325 263 264 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.72 $Y=3.33
+ $X2=24.72 $Y2=3.33
r326 260 261 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=23.76 $Y=3.33
+ $X2=23.76 $Y2=3.33
r327 257 258 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r328 254 255 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r329 251 252 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r330 249 264 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=24.24 $Y=3.33
+ $X2=24.72 $Y2=3.33
r331 249 261 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=24.24 $Y=3.33
+ $X2=23.76 $Y2=3.33
r332 248 249 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.24 $Y=3.33
+ $X2=24.24 $Y2=3.33
r333 246 260 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=23.88 $Y=3.33
+ $X2=23.795 $Y2=3.33
r334 246 248 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=23.88 $Y=3.33
+ $X2=24.24 $Y2=3.33
r335 245 263 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=24.595 $Y=3.33
+ $X2=24.777 $Y2=3.33
r336 245 248 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=24.595 $Y=3.33
+ $X2=24.24 $Y2=3.33
r337 244 261 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=22.8 $Y=3.33
+ $X2=23.76 $Y2=3.33
r338 243 244 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=22.8 $Y=3.33
+ $X2=22.8 $Y2=3.33
r339 241 244 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=21.84 $Y=3.33
+ $X2=22.8 $Y2=3.33
r340 240 241 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=21.84 $Y=3.33
+ $X2=21.84 $Y2=3.33
r341 238 241 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=20.88 $Y=3.33
+ $X2=21.84 $Y2=3.33
r342 237 238 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=20.88 $Y=3.33
+ $X2=20.88 $Y2=3.33
r343 234 237 594.995 $w=1.68e-07 $l=9.12e-06 $layer=LI1_cond $X=11.76 $Y=3.33
+ $X2=20.88 $Y2=3.33
r344 234 235 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r345 232 235 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r346 231 232 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r347 229 232 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r348 228 229 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r349 226 229 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r350 226 258 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r351 225 226 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r352 223 257 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.995 $Y=3.33
+ $X2=8.9 $Y2=3.33
r353 223 225 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.995 $Y=3.33
+ $X2=9.36 $Y2=3.33
r354 222 258 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r355 221 222 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r356 219 222 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r357 218 219 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r358 216 219 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r359 215 216 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r360 213 216 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r361 213 255 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r362 212 213 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r363 210 254 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=4.58 $Y2=3.33
r364 210 212 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=5.04 $Y2=3.33
r365 209 255 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r366 208 209 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r367 206 209 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r368 205 206 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r369 203 206 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r370 202 203 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r371 200 203 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r372 200 252 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r373 199 200 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r374 197 251 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r375 197 199 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r376 195 238 2.34137 $w=4.9e-07 $l=8.4e-06 $layer=MET1_cond $X=12.48 $Y=3.33
+ $X2=20.88 $Y2=3.33
r377 195 235 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=12.48 $Y=3.33
+ $X2=11.76 $Y2=3.33
r378 193 243 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=22.85 $Y=3.33
+ $X2=22.8 $Y2=3.33
r379 193 194 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.85 $Y=3.33
+ $X2=22.935 $Y2=3.33
r380 191 240 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=21.99 $Y=3.33
+ $X2=21.84 $Y2=3.33
r381 191 192 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.99 $Y=3.33
+ $X2=22.075 $Y2=3.33
r382 190 243 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=22.16 $Y=3.33
+ $X2=22.8 $Y2=3.33
r383 190 192 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.16 $Y=3.33
+ $X2=22.075 $Y2=3.33
r384 188 237 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=21.05 $Y=3.33
+ $X2=20.88 $Y2=3.33
r385 188 189 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=21.05 $Y=3.33
+ $X2=21.175 $Y2=3.33
r386 187 240 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=21.3 $Y=3.33
+ $X2=21.84 $Y2=3.33
r387 187 189 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=21.3 $Y=3.33
+ $X2=21.175 $Y2=3.33
r388 185 231 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=11.315 $Y=3.33
+ $X2=11.28 $Y2=3.33
r389 185 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.315 $Y=3.33
+ $X2=11.48 $Y2=3.33
r390 184 234 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=11.645 $Y=3.33
+ $X2=11.76 $Y2=3.33
r391 184 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.645 $Y=3.33
+ $X2=11.48 $Y2=3.33
r392 182 228 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.32 $Y2=3.33
r393 182 183 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.62 $Y2=3.33
r394 181 231 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=10.705 $Y=3.33
+ $X2=11.28 $Y2=3.33
r395 181 183 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.705 $Y=3.33
+ $X2=10.62 $Y2=3.33
r396 179 225 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.665 $Y=3.33
+ $X2=9.36 $Y2=3.33
r397 179 180 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.665 $Y=3.33
+ $X2=9.76 $Y2=3.33
r398 178 228 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=9.855 $Y=3.33
+ $X2=10.32 $Y2=3.33
r399 178 180 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.855 $Y=3.33
+ $X2=9.76 $Y2=3.33
r400 176 221 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=7.92 $Y2=3.33
r401 176 177 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=8.02 $Y2=3.33
r402 174 218 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.065 $Y=3.33
+ $X2=6.96 $Y2=3.33
r403 174 175 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.065 $Y=3.33
+ $X2=7.16 $Y2=3.33
r404 173 221 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.255 $Y=3.33
+ $X2=7.92 $Y2=3.33
r405 173 175 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.255 $Y=3.33
+ $X2=7.16 $Y2=3.33
r406 171 215 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.205 $Y=3.33
+ $X2=6 $Y2=3.33
r407 171 172 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.205 $Y=3.33
+ $X2=6.3 $Y2=3.33
r408 170 218 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.395 $Y=3.33
+ $X2=6.96 $Y2=3.33
r409 170 172 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.395 $Y=3.33
+ $X2=6.3 $Y2=3.33
r410 168 212 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.345 $Y=3.33
+ $X2=5.04 $Y2=3.33
r411 168 169 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.345 $Y=3.33
+ $X2=5.44 $Y2=3.33
r412 167 215 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.535 $Y=3.33
+ $X2=6 $Y2=3.33
r413 167 169 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.535 $Y=3.33
+ $X2=5.44 $Y2=3.33
r414 165 208 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=3.6 $Y2=3.33
r415 165 166 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=3.72 $Y2=3.33
r416 163 205 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.64 $Y2=3.33
r417 163 164 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.86 $Y2=3.33
r418 162 208 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r419 162 164 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.86 $Y2=3.33
r420 160 202 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r421 160 161 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2 $Y2=3.33
r422 159 205 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.64 $Y2=3.33
r423 159 161 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2 $Y2=3.33
r424 157 199 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r425 157 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.1 $Y2=3.33
r426 156 202 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.68 $Y2=3.33
r427 156 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.1 $Y2=3.33
r428 152 155 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=24.72 $Y=1.98
+ $X2=24.72 $Y2=2.95
r429 150 263 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=24.72 $Y=3.245
+ $X2=24.777 $Y2=3.33
r430 150 155 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=24.72 $Y=3.245
+ $X2=24.72 $Y2=2.95
r431 146 149 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=23.795 $Y=2.21
+ $X2=23.795 $Y2=2.95
r432 144 260 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=23.795 $Y=3.245
+ $X2=23.795 $Y2=3.33
r433 144 149 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=23.795 $Y=3.245
+ $X2=23.795 $Y2=2.95
r434 143 194 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=23.02 $Y=3.33
+ $X2=22.935 $Y2=3.33
r435 142 260 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=23.71 $Y=3.33
+ $X2=23.795 $Y2=3.33
r436 142 143 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=23.71 $Y=3.33
+ $X2=23.02 $Y2=3.33
r437 138 141 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=22.935 $Y=2.21
+ $X2=22.935 $Y2=2.95
r438 136 194 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.935 $Y=3.245
+ $X2=22.935 $Y2=3.33
r439 136 141 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=22.935 $Y=3.245
+ $X2=22.935 $Y2=2.95
r440 132 192 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.075 $Y=3.245
+ $X2=22.075 $Y2=3.33
r441 132 134 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=22.075 $Y=3.245
+ $X2=22.075 $Y2=2.33
r442 128 131 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=21.175 $Y=1.98
+ $X2=21.175 $Y2=2.95
r443 126 189 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=21.175 $Y=3.245
+ $X2=21.175 $Y2=3.33
r444 126 131 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=21.175 $Y=3.245
+ $X2=21.175 $Y2=2.95
r445 122 186 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.48 $Y=3.245
+ $X2=11.48 $Y2=3.33
r446 122 124 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=11.48 $Y=3.245
+ $X2=11.48 $Y2=2.53
r447 118 121 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=10.62 $Y=1.98
+ $X2=10.62 $Y2=2.95
r448 116 183 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.62 $Y=3.245
+ $X2=10.62 $Y2=3.33
r449 116 121 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.62 $Y=3.245
+ $X2=10.62 $Y2=2.95
r450 112 180 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=3.245
+ $X2=9.76 $Y2=3.33
r451 112 114 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=9.76 $Y=3.245
+ $X2=9.76 $Y2=2.37
r452 108 257 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=3.245
+ $X2=8.9 $Y2=3.33
r453 108 110 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=8.9 $Y=3.245
+ $X2=8.9 $Y2=2.37
r454 107 177 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.115 $Y=3.33
+ $X2=8.02 $Y2=3.33
r455 106 257 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=8.9 $Y2=3.33
r456 106 107 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=8.115 $Y2=3.33
r457 102 177 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=3.245
+ $X2=8.02 $Y2=3.33
r458 102 104 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=8.02 $Y=3.245
+ $X2=8.02 $Y2=2.37
r459 98 175 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.16 $Y=3.245
+ $X2=7.16 $Y2=3.33
r460 98 100 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=7.16 $Y=3.245
+ $X2=7.16 $Y2=2.37
r461 94 172 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=3.245
+ $X2=6.3 $Y2=3.33
r462 94 96 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=6.3 $Y=3.245
+ $X2=6.3 $Y2=2.37
r463 90 169 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=3.33
r464 90 92 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=2.37
r465 86 254 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=3.245
+ $X2=4.58 $Y2=3.33
r466 86 88 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=4.58 $Y=3.245
+ $X2=4.58 $Y2=2.37
r467 85 166 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.72 $Y2=3.33
r468 84 254 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.485 $Y=3.33
+ $X2=4.58 $Y2=3.33
r469 84 85 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.485 $Y=3.33
+ $X2=3.815 $Y2=3.33
r470 80 166 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=3.245
+ $X2=3.72 $Y2=3.33
r471 80 82 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=3.72 $Y=3.245
+ $X2=3.72 $Y2=2.37
r472 76 79 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.86 $Y=2.02
+ $X2=2.86 $Y2=2.95
r473 74 164 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=3.245
+ $X2=2.86 $Y2=3.33
r474 74 79 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.86 $Y=3.245
+ $X2=2.86 $Y2=2.95
r475 70 161 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=3.33
r476 70 72 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=2.33
r477 66 69 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=1.1 $Y=1.98 $X2=1.1
+ $Y2=2.95
r478 64 158 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=3.245
+ $X2=1.1 $Y2=3.33
r479 64 69 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=3.245
+ $X2=1.1 $Y2=2.95
r480 60 63 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=0.28 $Y=1.98
+ $X2=0.28 $Y2=2.95
r481 58 251 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r482 58 63 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.95
r483 19 155 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=24.54
+ $Y=1.835 $X2=24.68 $Y2=2.95
r484 19 152 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=24.54
+ $Y=1.835 $X2=24.68 $Y2=1.98
r485 18 149 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=23.655
+ $Y=1.835 $X2=23.795 $Y2=2.95
r486 18 146 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=23.655
+ $Y=1.835 $X2=23.795 $Y2=2.21
r487 17 141 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=22.795
+ $Y=1.835 $X2=22.935 $Y2=2.95
r488 17 138 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=22.795
+ $Y=1.835 $X2=22.935 $Y2=2.21
r489 16 134 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=21.935
+ $Y=1.835 $X2=22.075 $Y2=2.33
r490 15 131 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=21.07
+ $Y=1.835 $X2=21.215 $Y2=2.95
r491 15 128 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=21.07
+ $Y=1.835 $X2=21.215 $Y2=1.98
r492 14 124 300 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=2 $X=11.34
+ $Y=1.835 $X2=11.48 $Y2=2.53
r493 13 121 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.48
+ $Y=1.835 $X2=10.62 $Y2=2.95
r494 13 118 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.48
+ $Y=1.835 $X2=10.62 $Y2=1.98
r495 12 114 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=9.62
+ $Y=1.835 $X2=9.76 $Y2=2.37
r496 11 110 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=8.76
+ $Y=1.835 $X2=8.9 $Y2=2.37
r497 10 104 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=7.88
+ $Y=1.835 $X2=8.02 $Y2=2.37
r498 9 100 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=7.02
+ $Y=1.835 $X2=7.16 $Y2=2.37
r499 8 96 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=6.16
+ $Y=1.835 $X2=6.3 $Y2=2.37
r500 7 92 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=5.3
+ $Y=1.835 $X2=5.44 $Y2=2.37
r501 6 88 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=1.835 $X2=4.58 $Y2=2.37
r502 5 82 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=2.37
r503 4 79 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.95
r504 4 76 400 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.02
r505 3 72 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.33
r506 2 69 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.95
r507 2 66 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=1.98
r508 1 63 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.95
r509 1 60 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_630_367# 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 17 18 19 20 63 67 71 75 79 83 87 91 94 97 99 100 102 105 107 109
+ 110 111 112 115 119 123 127 131 135 139 143 147 151 155 159 163 167 171 175
+ 179 184 186 188 190 192 194 196 198 200 202 205 206 207 208 209 210 211 212
r342 179 182 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=20.225 $Y=1.98
+ $X2=20.225 $Y2=2.66
r343 177 182 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=20.225 $Y=2.885
+ $X2=20.225 $Y2=2.66
r344 176 212 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=19.53 $Y=2.975
+ $X2=19.365 $Y2=2.975
r345 175 177 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=20.06 $Y=2.975
+ $X2=20.225 $Y2=2.885
r346 175 176 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=20.06 $Y=2.975
+ $X2=19.53 $Y2=2.975
r347 171 174 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=19.365 $Y=1.98
+ $X2=19.365 $Y2=2.66
r348 169 212 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=19.365 $Y=2.885
+ $X2=19.365 $Y2=2.975
r349 169 174 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=19.365 $Y=2.885
+ $X2=19.365 $Y2=2.66
r350 168 211 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=18.67 $Y=2.975
+ $X2=18.505 $Y2=2.975
r351 167 212 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=19.2 $Y=2.975
+ $X2=19.365 $Y2=2.975
r352 167 168 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=19.2 $Y=2.975
+ $X2=18.67 $Y2=2.975
r353 163 166 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=18.505 $Y=1.98
+ $X2=18.505 $Y2=2.66
r354 161 211 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=18.505 $Y=2.885
+ $X2=18.505 $Y2=2.975
r355 161 166 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=18.505 $Y=2.885
+ $X2=18.505 $Y2=2.66
r356 160 210 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=17.81 $Y=2.975
+ $X2=17.645 $Y2=2.975
r357 159 211 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=18.34 $Y=2.975
+ $X2=18.505 $Y2=2.975
r358 159 160 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=18.34 $Y=2.975
+ $X2=17.81 $Y2=2.975
r359 155 158 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=17.645 $Y=1.98
+ $X2=17.645 $Y2=2.66
r360 153 210 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=17.645 $Y=2.885
+ $X2=17.645 $Y2=2.975
r361 153 158 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=17.645 $Y=2.885
+ $X2=17.645 $Y2=2.66
r362 152 209 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=16.95 $Y=2.975
+ $X2=16.785 $Y2=2.975
r363 151 210 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=17.48 $Y=2.975
+ $X2=17.645 $Y2=2.975
r364 151 152 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=17.48 $Y=2.975
+ $X2=16.95 $Y2=2.975
r365 147 150 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.785 $Y=1.98
+ $X2=16.785 $Y2=2.66
r366 145 209 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=16.785 $Y=2.885
+ $X2=16.785 $Y2=2.975
r367 145 150 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=16.785 $Y=2.885
+ $X2=16.785 $Y2=2.66
r368 144 208 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=16.09 $Y=2.975
+ $X2=15.925 $Y2=2.975
r369 143 209 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=16.62 $Y=2.975
+ $X2=16.785 $Y2=2.975
r370 143 144 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=16.62 $Y=2.975
+ $X2=16.09 $Y2=2.975
r371 139 142 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=15.925 $Y=1.98
+ $X2=15.925 $Y2=2.66
r372 137 208 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=15.925 $Y=2.885
+ $X2=15.925 $Y2=2.975
r373 137 142 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=15.925 $Y=2.885
+ $X2=15.925 $Y2=2.66
r374 136 207 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=15.23 $Y=2.975
+ $X2=15.065 $Y2=2.975
r375 135 208 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=15.76 $Y=2.975
+ $X2=15.925 $Y2=2.975
r376 135 136 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=15.76 $Y=2.975
+ $X2=15.23 $Y2=2.975
r377 131 134 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=15.065 $Y=1.98
+ $X2=15.065 $Y2=2.66
r378 129 207 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=15.065 $Y=2.885
+ $X2=15.065 $Y2=2.975
r379 129 134 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=15.065 $Y=2.885
+ $X2=15.065 $Y2=2.66
r380 128 206 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.37 $Y=2.975
+ $X2=14.205 $Y2=2.975
r381 127 207 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.9 $Y=2.975
+ $X2=15.065 $Y2=2.975
r382 127 128 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=14.9 $Y=2.975
+ $X2=14.37 $Y2=2.975
r383 123 126 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=14.205 $Y=1.98
+ $X2=14.205 $Y2=2.66
r384 121 206 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=14.205 $Y=2.885
+ $X2=14.205 $Y2=2.975
r385 121 126 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=14.205 $Y=2.885
+ $X2=14.205 $Y2=2.66
r386 120 205 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.51 $Y=2.975
+ $X2=13.345 $Y2=2.975
r387 119 206 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.04 $Y=2.975
+ $X2=14.205 $Y2=2.975
r388 119 120 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=14.04 $Y=2.975
+ $X2=13.51 $Y2=2.975
r389 115 118 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.345 $Y=1.98
+ $X2=13.345 $Y2=2.66
r390 113 205 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=13.345 $Y=2.885
+ $X2=13.345 $Y2=2.975
r391 113 118 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=13.345 $Y=2.885
+ $X2=13.345 $Y2=2.66
r392 111 205 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.18 $Y=2.975
+ $X2=13.345 $Y2=2.975
r393 111 112 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=13.18 $Y=2.975
+ $X2=12.65 $Y2=2.975
r394 110 112 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=12.485
+ $Y=2.885 $X2=12.65 $Y2=2.975
r395 109 204 2.9017 $w=3.3e-07 $l=1.13e-07 $layer=LI1_cond $X=12.485 $Y=2.185
+ $X2=12.485 $Y2=2.072
r396 109 110 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=12.485 $Y=2.185
+ $X2=12.485 $Y2=2.885
r397 108 202 1.72457 $w=2.25e-07 $l=1.25e-07 $layer=LI1_cond $X=11.135 $Y=2.072
+ $X2=11.01 $Y2=2.072
r398 107 204 4.237 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=12.32 $Y=2.072
+ $X2=12.485 $Y2=2.072
r399 107 108 60.6953 $w=2.23e-07 $l=1.185e-06 $layer=LI1_cond $X=12.32 $Y=2.072
+ $X2=11.135 $Y2=2.072
r400 103 202 4.72821 $w=2.5e-07 $l=1.13e-07 $layer=LI1_cond $X=11.01 $Y=2.185
+ $X2=11.01 $Y2=2.072
r401 103 105 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=11.01 $Y=2.185
+ $X2=11.01 $Y2=2.44
r402 102 202 4.72821 $w=2.5e-07 $l=1.12e-07 $layer=LI1_cond $X=11.01 $Y=1.96
+ $X2=11.01 $Y2=2.072
r403 101 102 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=11.01 $Y=1.635
+ $X2=11.01 $Y2=1.96
r404 99 101 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.885 $Y=1.55
+ $X2=11.01 $Y2=1.635
r405 99 100 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.885 $Y=1.55
+ $X2=10.355 $Y2=1.55
r406 95 200 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.19 $Y=2.035
+ $X2=10.19 $Y2=1.95
r407 95 97 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=10.19 $Y=2.035
+ $X2=10.19 $Y2=2.9
r408 94 200 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.19 $Y=1.865
+ $X2=10.19 $Y2=1.95
r409 93 100 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.19 $Y=1.635
+ $X2=10.355 $Y2=1.55
r410 93 94 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=10.19 $Y=1.635
+ $X2=10.19 $Y2=1.865
r411 92 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=1.95
+ $X2=9.33 $Y2=1.95
r412 91 200 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.025 $Y=1.95
+ $X2=10.19 $Y2=1.95
r413 91 92 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.025 $Y=1.95
+ $X2=9.495 $Y2=1.95
r414 88 196 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.635 $Y=1.95
+ $X2=8.47 $Y2=1.95
r415 87 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.165 $Y=1.95
+ $X2=9.33 $Y2=1.95
r416 87 88 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.165 $Y=1.95
+ $X2=8.635 $Y2=1.95
r417 84 194 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=1.95
+ $X2=7.59 $Y2=1.95
r418 83 196 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.305 $Y=1.95
+ $X2=8.47 $Y2=1.95
r419 83 84 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.305 $Y=1.95
+ $X2=7.755 $Y2=1.95
r420 80 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.895 $Y=1.95
+ $X2=6.73 $Y2=1.95
r421 79 194 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.425 $Y=1.95
+ $X2=7.59 $Y2=1.95
r422 79 80 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.425 $Y=1.95
+ $X2=6.895 $Y2=1.95
r423 76 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.035 $Y=1.95
+ $X2=5.87 $Y2=1.95
r424 75 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.565 $Y=1.95
+ $X2=6.73 $Y2=1.95
r425 75 76 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.565 $Y=1.95
+ $X2=6.035 $Y2=1.95
r426 72 188 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=1.95
+ $X2=5.01 $Y2=1.95
r427 71 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.705 $Y=1.95
+ $X2=5.87 $Y2=1.95
r428 71 72 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.705 $Y=1.95
+ $X2=5.175 $Y2=1.95
r429 68 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=1.95
+ $X2=4.15 $Y2=1.95
r430 67 188 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=1.95
+ $X2=5.01 $Y2=1.95
r431 67 68 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.845 $Y=1.95
+ $X2=4.315 $Y2=1.95
r432 64 184 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=1.95
+ $X2=3.29 $Y2=1.95
r433 63 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=1.95
+ $X2=4.15 $Y2=1.95
r434 63 64 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.985 $Y=1.95
+ $X2=3.455 $Y2=1.95
r435 20 182 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=20.085
+ $Y=1.525 $X2=20.225 $Y2=2.66
r436 20 179 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=20.085
+ $Y=1.525 $X2=20.225 $Y2=1.98
r437 19 174 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=19.225
+ $Y=1.525 $X2=19.365 $Y2=2.66
r438 19 171 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=19.225
+ $Y=1.525 $X2=19.365 $Y2=1.98
r439 18 166 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=18.365
+ $Y=1.525 $X2=18.505 $Y2=2.66
r440 18 163 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=18.365
+ $Y=1.525 $X2=18.505 $Y2=1.98
r441 17 158 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=17.505
+ $Y=1.525 $X2=17.645 $Y2=2.66
r442 17 155 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=17.505
+ $Y=1.525 $X2=17.645 $Y2=1.98
r443 16 150 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=16.645
+ $Y=1.525 $X2=16.785 $Y2=2.66
r444 16 147 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=16.645
+ $Y=1.525 $X2=16.785 $Y2=1.98
r445 15 142 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=15.785
+ $Y=1.525 $X2=15.925 $Y2=2.66
r446 15 139 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=15.785
+ $Y=1.525 $X2=15.925 $Y2=1.98
r447 14 134 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=14.925
+ $Y=1.525 $X2=15.065 $Y2=2.66
r448 14 131 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=14.925
+ $Y=1.525 $X2=15.065 $Y2=1.98
r449 13 126 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=14.065
+ $Y=1.525 $X2=14.205 $Y2=2.66
r450 13 123 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=14.065
+ $Y=1.525 $X2=14.205 $Y2=1.98
r451 12 118 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=13.205
+ $Y=1.525 $X2=13.345 $Y2=2.66
r452 12 115 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=13.205
+ $Y=1.525 $X2=13.345 $Y2=1.98
r453 11 204 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=12.345
+ $Y=1.525 $X2=12.485 $Y2=2.125
r454 10 202 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.91
+ $Y=1.835 $X2=11.05 $Y2=1.98
r455 10 105 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=10.91
+ $Y=1.835 $X2=11.05 $Y2=2.44
r456 9 200 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.05
+ $Y=1.835 $X2=10.19 $Y2=1.98
r457 9 97 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=10.05
+ $Y=1.835 $X2=10.19 $Y2=2.9
r458 8 198 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=9.19
+ $Y=1.835 $X2=9.33 $Y2=2.03
r459 7 196 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=8.33
+ $Y=1.835 $X2=8.47 $Y2=2.03
r460 6 194 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=7.45
+ $Y=1.835 $X2=7.59 $Y2=2.03
r461 5 192 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=6.59
+ $Y=1.835 $X2=6.73 $Y2=2.03
r462 4 190 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=5.73
+ $Y=1.835 $X2=5.87 $Y2=2.03
r463 3 188 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=4.87
+ $Y=1.835 $X2=5.01 $Y2=2.03
r464 2 186 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=4.01
+ $Y=1.835 $X2=4.15 $Y2=2.03
r465 1 184 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=2.03
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 55 69 71 75 77 81 83 87 89 93 95 99 101 105 107 111 113 117 119 123
+ 125 127 129 132 134 136 138 140 142 144 146 148 151 152 153 159 161
c200 161 0 1.47022e-19 $X=11.76 $Y=0.925
c201 159 0 4.06089e-20 $X=11.77 $Y=1.505
r202 158 161 0.393548 $w=9.28e-07 $l=3e-08 $layer=LI1_cond $X=11.77 $Y=0.895
+ $X2=11.77 $Y2=0.925
r203 153 159 2.24069 $w=9.3e-07 $l=1.37e-07 $layer=LI1_cond $X=11.77 $Y=1.642
+ $X2=11.77 $Y2=1.505
r204 152 159 2.75484 $w=9.28e-07 $l=2.1e-07 $layer=LI1_cond $X=11.77 $Y=1.295
+ $X2=11.77 $Y2=1.505
r205 151 158 2.64086 $w=9.3e-07 $l=1.25e-07 $layer=LI1_cond $X=11.77 $Y=0.77
+ $X2=11.77 $Y2=0.895
r206 151 152 4.49957 $w=9.28e-07 $l=3.43e-07 $layer=LI1_cond $X=11.77 $Y=0.952
+ $X2=11.77 $Y2=1.295
r207 151 161 0.354194 $w=9.28e-07 $l=2.7e-08 $layer=LI1_cond $X=11.77 $Y=0.952
+ $X2=11.77 $Y2=0.925
r208 127 150 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=20.695 $Y=1.725
+ $X2=20.695 $Y2=1.61
r209 127 129 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=20.695 $Y=1.725
+ $X2=20.695 $Y2=2.64
r210 126 148 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=19.89 $Y=1.61
+ $X2=19.795 $Y2=1.61
r211 125 150 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=20.57 $Y=1.61
+ $X2=20.695 $Y2=1.61
r212 125 126 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=20.57 $Y=1.61
+ $X2=19.89 $Y2=1.61
r213 121 148 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=19.795 $Y=1.725
+ $X2=19.795 $Y2=1.61
r214 121 123 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=19.795 $Y=1.725
+ $X2=19.795 $Y2=2.55
r215 120 146 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=19.03 $Y=1.61
+ $X2=18.935 $Y2=1.61
r216 119 148 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=19.7 $Y=1.61
+ $X2=19.795 $Y2=1.61
r217 119 120 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=19.7 $Y=1.61
+ $X2=19.03 $Y2=1.61
r218 115 146 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=18.935 $Y=1.725
+ $X2=18.935 $Y2=1.61
r219 115 117 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=18.935 $Y=1.725
+ $X2=18.935 $Y2=2.55
r220 114 144 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=18.17 $Y=1.61
+ $X2=18.075 $Y2=1.61
r221 113 146 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=18.84 $Y=1.61
+ $X2=18.935 $Y2=1.61
r222 113 114 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=18.84 $Y=1.61
+ $X2=18.17 $Y2=1.61
r223 109 144 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=18.075 $Y=1.725
+ $X2=18.075 $Y2=1.61
r224 109 111 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=18.075 $Y=1.725
+ $X2=18.075 $Y2=2.55
r225 108 142 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=17.31 $Y=1.61
+ $X2=17.215 $Y2=1.61
r226 107 144 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=17.98 $Y=1.61
+ $X2=18.075 $Y2=1.61
r227 107 108 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=17.98 $Y=1.61
+ $X2=17.31 $Y2=1.61
r228 103 142 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=17.215 $Y=1.725
+ $X2=17.215 $Y2=1.61
r229 103 105 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=17.215 $Y=1.725
+ $X2=17.215 $Y2=2.55
r230 102 140 4.47804 $w=2.25e-07 $l=2.36749e-07 $layer=LI1_cond $X=16.45 $Y=1.61
+ $X2=16.26 $Y2=1.505
r231 101 142 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=17.12 $Y=1.61
+ $X2=17.215 $Y2=1.61
r232 101 102 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=17.12 $Y=1.61
+ $X2=16.45 $Y2=1.61
r233 97 140 1.9579 $w=1.9e-07 $l=2.63249e-07 $layer=LI1_cond $X=16.355 $Y=1.725
+ $X2=16.26 $Y2=1.505
r234 97 99 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=16.355 $Y=1.725
+ $X2=16.355 $Y2=2.55
r235 96 138 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=15.59 $Y=1.615
+ $X2=15.495 $Y2=1.615
r236 95 140 4.47804 $w=2.25e-07 $l=1.1e-07 $layer=LI1_cond $X=16.26 $Y=1.615
+ $X2=16.26 $Y2=1.505
r237 95 96 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=16.26 $Y=1.615
+ $X2=15.59 $Y2=1.615
r238 91 138 1.87542 $w=1.9e-07 $l=1.1e-07 $layer=LI1_cond $X=15.495 $Y=1.725
+ $X2=15.495 $Y2=1.615
r239 91 93 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=15.495 $Y=1.725
+ $X2=15.495 $Y2=2.55
r240 90 136 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=14.73 $Y=1.615
+ $X2=14.635 $Y2=1.615
r241 89 138 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=15.4 $Y=1.615
+ $X2=15.495 $Y2=1.615
r242 89 90 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=15.4 $Y=1.615
+ $X2=14.73 $Y2=1.615
r243 85 136 1.87542 $w=1.9e-07 $l=1.1e-07 $layer=LI1_cond $X=14.635 $Y=1.725
+ $X2=14.635 $Y2=1.615
r244 85 87 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=14.635 $Y=1.725
+ $X2=14.635 $Y2=2.55
r245 84 134 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=13.87 $Y=1.615
+ $X2=13.775 $Y2=1.615
r246 83 136 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=14.54 $Y=1.615
+ $X2=14.635 $Y2=1.615
r247 83 84 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=14.54 $Y=1.615
+ $X2=13.87 $Y2=1.615
r248 79 134 1.87542 $w=1.9e-07 $l=1.1e-07 $layer=LI1_cond $X=13.775 $Y=1.725
+ $X2=13.775 $Y2=1.615
r249 79 81 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=13.775 $Y=1.725
+ $X2=13.775 $Y2=2.55
r250 78 132 4.12396 $w=2.47e-07 $l=1.07657e-07 $layer=LI1_cond $X=13.01 $Y=1.615
+ $X2=12.915 $Y2=1.642
r251 77 134 4.56504 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=13.68 $Y=1.615
+ $X2=13.775 $Y2=1.615
r252 77 78 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=13.68 $Y=1.615
+ $X2=13.01 $Y2=1.615
r253 73 132 2.30976 $w=1.9e-07 $l=1.38e-07 $layer=LI1_cond $X=12.915 $Y=1.78
+ $X2=12.915 $Y2=1.642
r254 73 75 19.2632 $w=1.88e-07 $l=3.3e-07 $layer=LI1_cond $X=12.915 $Y=1.78
+ $X2=12.915 $Y2=2.11
r255 72 153 7.60527 $w=2.75e-07 $l=4.65e-07 $layer=LI1_cond $X=12.235 $Y=1.642
+ $X2=11.77 $Y2=1.642
r256 71 132 4.12396 $w=2.47e-07 $l=9.5e-08 $layer=LI1_cond $X=12.82 $Y=1.642
+ $X2=12.915 $Y2=1.642
r257 71 72 24.5156 $w=2.73e-07 $l=5.85e-07 $layer=LI1_cond $X=12.82 $Y=1.642
+ $X2=12.235 $Y2=1.642
r258 67 69 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=14.375 $Y=0.77
+ $X2=15.235 $Y2=0.77
r259 65 67 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=13.515 $Y=0.77
+ $X2=14.375 $Y2=0.77
r260 63 65 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=12.655 $Y=0.77
+ $X2=13.515 $Y2=0.77
r261 61 151 12.9322 $w=2.5e-07 $l=4.65e-07 $layer=LI1_cond $X=12.235 $Y=0.77
+ $X2=11.77 $Y2=0.77
r262 61 63 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=12.235 $Y=0.77
+ $X2=12.655 $Y2=0.77
r263 57 60 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=9.915 $Y=0.77
+ $X2=10.935 $Y2=0.77
r264 55 151 12.9322 $w=2.5e-07 $l=4.65e-07 $layer=LI1_cond $X=11.305 $Y=0.77
+ $X2=11.77 $Y2=0.77
r265 55 60 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=11.305 $Y=0.77
+ $X2=10.935 $Y2=0.77
r266 18 150 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=20.515
+ $Y=1.525 $X2=20.655 $Y2=1.67
r267 18 129 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=20.515
+ $Y=1.525 $X2=20.655 $Y2=2.64
r268 17 148 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=19.655
+ $Y=1.525 $X2=19.795 $Y2=1.67
r269 17 123 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=19.655
+ $Y=1.525 $X2=19.795 $Y2=2.55
r270 16 146 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=18.795
+ $Y=1.525 $X2=18.935 $Y2=1.67
r271 16 117 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=18.795
+ $Y=1.525 $X2=18.935 $Y2=2.55
r272 15 144 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=17.935
+ $Y=1.525 $X2=18.075 $Y2=1.67
r273 15 111 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=17.935
+ $Y=1.525 $X2=18.075 $Y2=2.55
r274 14 142 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=17.075
+ $Y=1.525 $X2=17.215 $Y2=1.67
r275 14 105 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=17.075
+ $Y=1.525 $X2=17.215 $Y2=2.55
r276 13 140 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=16.215
+ $Y=1.525 $X2=16.355 $Y2=1.67
r277 13 99 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=16.215
+ $Y=1.525 $X2=16.355 $Y2=2.55
r278 12 138 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.355
+ $Y=1.525 $X2=15.495 $Y2=1.67
r279 12 93 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=15.355
+ $Y=1.525 $X2=15.495 $Y2=2.55
r280 11 136 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.495
+ $Y=1.525 $X2=14.635 $Y2=1.67
r281 11 87 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=14.495
+ $Y=1.525 $X2=14.635 $Y2=2.55
r282 10 134 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.635
+ $Y=1.525 $X2=13.775 $Y2=1.67
r283 10 81 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=13.635
+ $Y=1.525 $X2=13.775 $Y2=2.55
r284 9 132 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.775
+ $Y=1.525 $X2=12.915 $Y2=1.67
r285 9 75 300 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_PDIFF $count=2 $X=12.775
+ $Y=1.525 $X2=12.915 $Y2=2.11
r286 8 153 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.91
+ $Y=1.525 $X2=12.055 $Y2=1.67
r287 7 69 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=15.095
+ $Y=0.235 $X2=15.235 $Y2=0.73
r288 6 67 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=14.235
+ $Y=0.235 $X2=14.375 $Y2=0.73
r289 5 65 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=13.375
+ $Y=0.235 $X2=13.515 $Y2=0.73
r290 4 63 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=12.515
+ $Y=0.235 $X2=12.655 $Y2=0.73
r291 3 151 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=11.655
+ $Y=0.235 $X2=11.795 $Y2=0.73
r292 2 60 182 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_NDIFF $count=1 $X=10.715
+ $Y=0.235 $X2=10.935 $Y2=0.75
r293 1 57 182 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_NDIFF $count=1 $X=9.695
+ $Y=0.235 $X2=9.915 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 40
+ 42 46 50 54 58 62 66 70 74 78 82 86 90 93 94 96 97 99 100 102 103 105 106 108
+ 109 111 112 114 115 117 118 119 121 130 162 168 169 175 178 181
r243 181 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.76 $Y=0
+ $X2=23.76 $Y2=0
r244 178 179 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r245 175 176 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r246 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r247 169 182 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=24.72 $Y=0
+ $X2=23.76 $Y2=0
r248 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.72 $Y=0
+ $X2=24.72 $Y2=0
r249 166 181 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.89 $Y=0
+ $X2=23.725 $Y2=0
r250 166 168 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=23.89 $Y=0
+ $X2=24.72 $Y2=0
r251 165 182 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=23.28 $Y=0
+ $X2=23.76 $Y2=0
r252 164 165 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=23.28 $Y=0
+ $X2=23.28 $Y2=0
r253 162 181 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.56 $Y=0
+ $X2=23.725 $Y2=0
r254 162 164 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=23.56 $Y=0
+ $X2=23.28 $Y2=0
r255 161 165 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=22.32 $Y=0
+ $X2=23.28 $Y2=0
r256 160 161 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=22.32 $Y=0
+ $X2=22.32 $Y2=0
r257 158 161 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=21.36 $Y=0
+ $X2=22.32 $Y2=0
r258 157 158 0.715385 $w=1.7e-07 $l=2.21e-06 $layer=mcon $count=13 $X=21.36 $Y=0
+ $X2=21.36 $Y2=0
r259 154 157 782.888 $w=1.68e-07 $l=1.2e-05 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=21.36 $Y2=0
r260 154 155 0.715385 $w=1.7e-07 $l=2.21e-06 $layer=mcon $count=13 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r261 152 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r262 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r263 149 152 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.88 $Y2=0
r264 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r265 146 149 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.92 $Y2=0
r266 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r267 143 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r268 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r269 140 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r270 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r271 137 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r272 137 179 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=3.6 $Y2=0
r273 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r274 134 178 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0
+ $X2=3.575 $Y2=0
r275 134 136 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.74 $Y=0
+ $X2=4.08 $Y2=0
r276 133 179 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=3.6 $Y2=0
r277 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r278 130 178 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=0
+ $X2=3.575 $Y2=0
r279 130 132 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.41 $Y=0
+ $X2=3.12 $Y2=0
r280 129 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.12 $Y2=0
r281 129 176 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.2 $Y2=0
r282 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r283 126 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.22 $Y2=0
r284 126 128 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=2.16 $Y2=0
r285 125 176 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.2 $Y2=0
r286 125 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r287 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r288 122 172 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r289 122 124 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r290 121 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=1.22 $Y2=0
r291 121 124 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r292 119 158 2.47516 $w=4.9e-07 $l=8.88e-06 $layer=MET1_cond $X=12.48 $Y=0
+ $X2=21.36 $Y2=0
r293 119 155 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=12.48 $Y=0
+ $X2=9.36 $Y2=0
r294 117 160 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=22.54 $Y=0
+ $X2=22.32 $Y2=0
r295 117 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.54 $Y=0
+ $X2=22.705 $Y2=0
r296 116 164 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=22.87 $Y=0
+ $X2=23.28 $Y2=0
r297 116 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.87 $Y=0
+ $X2=22.705 $Y2=0
r298 114 157 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=21.52 $Y=0
+ $X2=21.36 $Y2=0
r299 114 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=21.52 $Y=0
+ $X2=21.685 $Y2=0
r300 113 160 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=21.85 $Y=0
+ $X2=22.32 $Y2=0
r301 113 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=21.85 $Y=0
+ $X2=21.685 $Y2=0
r302 111 151 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.89 $Y=0 $X2=8.88
+ $Y2=0
r303 111 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=0
+ $X2=8.975 $Y2=0
r304 110 154 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.06 $Y=0 $X2=9.36
+ $Y2=0
r305 110 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.06 $Y=0
+ $X2=8.975 $Y2=0
r306 108 148 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.03 $Y=0
+ $X2=7.92 $Y2=0
r307 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.03 $Y=0
+ $X2=8.115 $Y2=0
r308 107 151 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.2 $Y=0 $X2=8.88
+ $Y2=0
r309 107 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.2 $Y=0 $X2=8.115
+ $Y2=0
r310 105 145 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=0
+ $X2=6.96 $Y2=0
r311 105 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=0
+ $X2=7.255 $Y2=0
r312 104 148 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.34 $Y=0
+ $X2=7.92 $Y2=0
r313 104 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.34 $Y=0
+ $X2=7.255 $Y2=0
r314 102 142 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.15 $Y=0 $X2=6
+ $Y2=0
r315 102 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.15 $Y=0
+ $X2=6.315 $Y2=0
r316 101 145 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r317 101 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0
+ $X2=6.315 $Y2=0
r318 99 139 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.13 $Y=0 $X2=5.04
+ $Y2=0
r319 99 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=0
+ $X2=5.295 $Y2=0
r320 98 142 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.46 $Y=0 $X2=6
+ $Y2=0
r321 98 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=0
+ $X2=5.295 $Y2=0
r322 96 136 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.08
+ $Y2=0
r323 96 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.435
+ $Y2=0
r324 95 139 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=5.04
+ $Y2=0
r325 95 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.435
+ $Y2=0
r326 93 128 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.16
+ $Y2=0
r327 93 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.505
+ $Y2=0
r328 92 132 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=3.12
+ $Y2=0
r329 92 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.505
+ $Y2=0
r330 88 181 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=23.725 $Y=0.085
+ $X2=23.725 $Y2=0
r331 88 90 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=23.725 $Y=0.085
+ $X2=23.725 $Y2=0.38
r332 84 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=22.705 $Y=0.085
+ $X2=22.705 $Y2=0
r333 84 86 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=22.705 $Y=0.085
+ $X2=22.705 $Y2=0.43
r334 80 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=21.685 $Y=0.085
+ $X2=21.685 $Y2=0
r335 80 82 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=21.685 $Y=0.085
+ $X2=21.685 $Y2=0.43
r336 76 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.975 $Y=0.085
+ $X2=8.975 $Y2=0
r337 76 78 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.975 $Y=0.085
+ $X2=8.975 $Y2=0.515
r338 72 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0
r339 72 74 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0.515
r340 68 106 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.255 $Y=0.085
+ $X2=7.255 $Y2=0
r341 68 70 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.255 $Y=0.085
+ $X2=7.255 $Y2=0.515
r342 64 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.315 $Y=0.085
+ $X2=6.315 $Y2=0
r343 64 66 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=6.315 $Y=0.085
+ $X2=6.315 $Y2=0.385
r344 60 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.295 $Y=0.085
+ $X2=5.295 $Y2=0
r345 60 62 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=5.295 $Y=0.085
+ $X2=5.295 $Y2=0.385
r346 56 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0
r347 56 58 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0.385
r348 52 178 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0
r349 52 54 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0.385
r350 48 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0
r351 48 50 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0.28
r352 44 175 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r353 44 46 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.36
r354 40 172 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r355 40 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.38
r356 13 90 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=23.505
+ $Y=0.235 $X2=23.725 $Y2=0.38
r357 12 86 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=22.485
+ $Y=0.235 $X2=22.705 $Y2=0.43
r358 11 82 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=21.54
+ $Y=0.235 $X2=21.685 $Y2=0.43
r359 10 78 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=8.835
+ $Y=0.235 $X2=8.975 $Y2=0.515
r360 9 74 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.235 $X2=8.115 $Y2=0.515
r361 8 70 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=7.115
+ $Y=0.235 $X2=7.255 $Y2=0.515
r362 7 66 182 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_NDIFF $count=1 $X=6.095
+ $Y=0.235 $X2=6.315 $Y2=0.385
r363 6 62 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=5.155
+ $Y=0.235 $X2=5.295 $Y2=0.385
r364 5 58 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.295
+ $Y=0.235 $X2=4.435 $Y2=0.385
r365 4 54 182 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.235 $X2=3.575 $Y2=0.385
r366 3 50 182 $w=1.7e-07 $l=2.76586e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.235 $X2=2.505 $Y2=0.28
r367 2 46 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.235
+ $X2=1.22 $Y2=0.36
r368 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_584_47# 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 48 50 51 54 56 60 62 66 68 70 74 75 76 79 81 85 87 92 93 94 107 108
+ 109 110 111 112 113
c212 110 0 7.60313e-20 $X=6.825 $Y=0.74
c213 76 0 1.98224e-19 $X=6.99 $Y=1.08
r214 113 116 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=15.745 $Y=0.37
+ $X2=15.745 $Y2=0.535
r215 104 106 45.4199 $w=2.08e-07 $l=8.6e-07 $layer=LI1_cond $X=13.945 $Y=0.37
+ $X2=14.805 $Y2=0.37
r216 102 104 45.4199 $w=2.08e-07 $l=8.6e-07 $layer=LI1_cond $X=13.085 $Y=0.37
+ $X2=13.945 $Y2=0.37
r217 100 102 45.4199 $w=2.08e-07 $l=8.6e-07 $layer=LI1_cond $X=12.225 $Y=0.37
+ $X2=13.085 $Y2=0.37
r218 98 100 45.4199 $w=2.08e-07 $l=8.6e-07 $layer=LI1_cond $X=11.365 $Y=0.37
+ $X2=12.225 $Y2=0.37
r219 96 98 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=10.425 $Y=0.37
+ $X2=11.365 $Y2=0.37
r220 94 96 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=9.57 $Y=0.37
+ $X2=10.425 $Y2=0.37
r221 93 113 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=15.58 $Y=0.37
+ $X2=15.745 $Y2=0.37
r222 93 106 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=15.58 $Y=0.37
+ $X2=14.805 $Y2=0.37
r223 90 92 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=9.405 $Y=0.995
+ $X2=9.405 $Y2=0.58
r224 89 94 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=9.405 $Y=0.475
+ $X2=9.57 $Y2=0.37
r225 89 92 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=9.405 $Y=0.475
+ $X2=9.405 $Y2=0.58
r226 88 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.71 $Y=1.08
+ $X2=8.545 $Y2=1.08
r227 87 90 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.24 $Y=1.08
+ $X2=9.405 $Y2=0.995
r228 87 88 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.24 $Y=1.08
+ $X2=8.71 $Y2=1.08
r229 83 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=0.995
+ $X2=8.545 $Y2=1.08
r230 83 85 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=8.545 $Y=0.995
+ $X2=8.545 $Y2=0.58
r231 82 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.85 $Y=1.08
+ $X2=7.685 $Y2=1.08
r232 81 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.38 $Y=1.08
+ $X2=8.545 $Y2=1.08
r233 81 82 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.38 $Y=1.08
+ $X2=7.85 $Y2=1.08
r234 77 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=0.995
+ $X2=7.685 $Y2=1.08
r235 77 79 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=7.685 $Y=0.995
+ $X2=7.685 $Y2=0.58
r236 75 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.52 $Y=1.08
+ $X2=7.685 $Y2=1.08
r237 75 76 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.52 $Y=1.08
+ $X2=6.99 $Y2=1.08
r238 74 76 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.825 $Y=0.995
+ $X2=6.99 $Y2=1.08
r239 73 110 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.825 $Y=0.825
+ $X2=6.825 $Y2=0.74
r240 73 74 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.825 $Y=0.825
+ $X2=6.825 $Y2=0.995
r241 70 110 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.825 $Y=0.655
+ $X2=6.825 $Y2=0.74
r242 70 72 2.77273 $w=3.3e-07 $l=7.5e-08 $layer=LI1_cond $X=6.825 $Y=0.655
+ $X2=6.825 $Y2=0.58
r243 69 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=0.74
+ $X2=5.805 $Y2=0.74
r244 68 110 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.66 $Y=0.74
+ $X2=6.825 $Y2=0.74
r245 68 69 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.66 $Y=0.74
+ $X2=5.97 $Y2=0.74
r246 64 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=0.655
+ $X2=5.805 $Y2=0.74
r247 64 66 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.805 $Y=0.655
+ $X2=5.805 $Y2=0.545
r248 63 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=0.74
+ $X2=4.865 $Y2=0.74
r249 62 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.64 $Y=0.74
+ $X2=5.805 $Y2=0.74
r250 62 63 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.64 $Y=0.74
+ $X2=4.95 $Y2=0.74
r251 58 108 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=0.655
+ $X2=4.865 $Y2=0.74
r252 58 60 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.865 $Y=0.655
+ $X2=4.865 $Y2=0.545
r253 57 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=0.74
+ $X2=4.005 $Y2=0.74
r254 56 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=0.74
+ $X2=4.865 $Y2=0.74
r255 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.78 $Y=0.74
+ $X2=4.09 $Y2=0.74
r256 52 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.005 $Y=0.655
+ $X2=4.005 $Y2=0.74
r257 52 54 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.005 $Y=0.655
+ $X2=4.005 $Y2=0.545
r258 50 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=0.74
+ $X2=4.005 $Y2=0.74
r259 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.92 $Y=0.74
+ $X2=3.23 $Y2=0.74
r260 46 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.065 $Y=0.655
+ $X2=3.23 $Y2=0.74
r261 46 48 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.065 $Y=0.655
+ $X2=3.065 $Y2=0.545
r262 15 116 182 $w=1.7e-07 $l=3.94968e-07 $layer=licon1_NDIFF $count=1 $X=15.525
+ $Y=0.235 $X2=15.745 $Y2=0.535
r263 14 106 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=14.665
+ $Y=0.235 $X2=14.805 $Y2=0.38
r264 13 104 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=13.805
+ $Y=0.235 $X2=13.945 $Y2=0.38
r265 12 102 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=12.945
+ $Y=0.235 $X2=13.085 $Y2=0.38
r266 11 100 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=12.085
+ $Y=0.235 $X2=12.225 $Y2=0.38
r267 10 98 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.225
+ $Y=0.235 $X2=11.365 $Y2=0.38
r268 9 96 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=10.205
+ $Y=0.235 $X2=10.425 $Y2=0.38
r269 8 92 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=9.265
+ $Y=0.235 $X2=9.405 $Y2=0.58
r270 7 85 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=8.405
+ $Y=0.235 $X2=8.545 $Y2=0.58
r271 6 79 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=7.545
+ $Y=0.235 $X2=7.685 $Y2=0.58
r272 5 72 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=6.685
+ $Y=0.235 $X2=6.825 $Y2=0.58
r273 4 66 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=5.665
+ $Y=0.235 $X2=5.805 $Y2=0.545
r274 3 60 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=4.725
+ $Y=0.235 $X2=4.865 $Y2=0.545
r275 2 54 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=3.865
+ $Y=0.235 $X2=4.005 $Y2=0.545
r276 1 48 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=2.92
+ $Y=0.235 $X2=3.065 $Y2=0.545
.ends

