* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32a_m A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_249_403# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.36e+11p ps=3.28e+06u
M1001 a_86_55# A3 a_321_403# VPB phighvt w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=1.638e+11p ps=1.62e+06u
M1002 VGND A2 a_249_81# VNB nshort w=420000u l=150000u
+  ad=4.263e+11p pd=3.71e+06u as=3.633e+11p ps=4.25e+06u
M1003 VPWR B1 a_566_403# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.029e+11p ps=1.33e+06u
M1004 a_249_81# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_86_55# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 a_321_403# A2 a_249_403# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_249_81# B1 a_86_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1008 a_86_55# B2 a_249_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_249_81# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_566_403# B2 a_86_55# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_86_55# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends
