* File: sky130_fd_sc_lp__dfrbp_1.pex.spice
* Created: Wed Sep  2 09:43:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFRBP_1%CLK 3 7 9 10 14
c34 7 0 1.3822e-19 $X=0.48 $Y=2.68
c35 3 0 4.07885e-20 $X=0.48 $Y=0.75
r36 14 17 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.592 $Y=1.805
+ $X2=0.592 $Y2=1.97
r37 14 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.592 $Y=1.805
+ $X2=0.592 $Y2=1.64
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.615
+ $Y=1.805 $X2=0.615 $Y2=1.805
r39 10 15 6.88472 $w=3.83e-07 $l=2.3e-07 $layer=LI1_cond $X=0.722 $Y=2.035
+ $X2=0.722 $Y2=1.805
r40 9 15 4.1907 $w=3.83e-07 $l=1.4e-07 $layer=LI1_cond $X=0.722 $Y=1.665
+ $X2=0.722 $Y2=1.805
r41 7 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.48 $Y=2.68 $X2=0.48
+ $Y2=1.97
r42 3 16 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.48 $Y=0.75 $X2=0.48
+ $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%D 3 6 9 10 11 12 13 17
c47 17 0 1.27153e-19 $X=2.49 $Y=1.65
c48 13 0 1.36523e-19 $X=2.16 $Y=1.665
r49 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.49
+ $Y=1.65 $X2=2.49 $Y2=1.65
r50 13 18 0.369697 $w=4.95e-07 $l=1.5e-08 $layer=LI1_cond $X=2.302 $Y=1.665
+ $X2=2.302 $Y2=1.65
r51 12 18 8.74949 $w=4.95e-07 $l=3.55e-07 $layer=LI1_cond $X=2.302 $Y=1.295
+ $X2=2.302 $Y2=1.65
r52 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.49 $Y=1.99
+ $X2=2.49 $Y2=1.65
r53 10 11 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.99
+ $X2=2.49 $Y2=2.155
r54 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.485
+ $X2=2.49 $Y2=1.65
r55 6 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.43 $Y=2.525
+ $X2=2.43 $Y2=2.155
r56 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.4 $Y=1.165 $X2=2.4
+ $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_197_108# 1 2 7 9 11 13 14 16 17 21 23 25
+ 27 28 31 33 35 38 39 41 45 51 52 53 54 58 62 73
c192 53 0 1.3822e-19 $X=1.252 $Y=2.1
c193 35 0 1.27153e-19 $X=3.095 $Y=0.715
c194 27 0 1.05547e-19 $X=1.252 $Y=1.722
c195 7 0 1.278e-20 $X=3.44 $Y=1.945
r196 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.405
+ $Y=1.78 $X2=3.405 $Y2=1.78
r197 59 62 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.18 $Y=1.78
+ $X2=3.405 $Y2=1.78
r198 54 56 12.6753 $w=2.08e-07 $l=2.4e-07 $layer=LI1_cond $X=2.15 $Y=0.715
+ $X2=2.15 $Y2=0.955
r199 51 53 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=1.23 $Y=2.35
+ $X2=1.23 $Y2=2.1
r200 46 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.555
+ $X2=6.53 $Y2=1.555
r201 46 70 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.365 $Y=1.555
+ $X2=6.15 $Y2=1.555
r202 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=1.555 $X2=6.365 $Y2=1.555
r203 43 45 40.9747 $w=1.78e-07 $l=6.65e-07 $layer=LI1_cond $X=6.36 $Y=0.89
+ $X2=6.36 $Y2=1.555
r204 42 67 2.11506 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=4.755 $Y=0.805
+ $X2=4.647 $Y2=0.805
r205 41 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.27 $Y=0.805
+ $X2=6.36 $Y2=0.89
r206 41 42 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=6.27 $Y=0.805
+ $X2=4.755 $Y2=0.805
r207 40 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=0.715
+ $X2=3.18 $Y2=0.715
r208 39 67 4.82418 $w=2.13e-07 $l=9e-08 $layer=LI1_cond $X=4.647 $Y=0.715
+ $X2=4.647 $Y2=0.805
r209 39 40 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=4.54 $Y=0.715
+ $X2=3.265 $Y2=0.715
r210 38 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.615
+ $X2=3.18 $Y2=1.78
r211 37 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=0.8 $X2=3.18
+ $Y2=0.715
r212 37 38 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.18 $Y=0.8
+ $X2=3.18 $Y2=1.615
r213 36 54 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.255 $Y=0.715
+ $X2=2.15 $Y2=0.715
r214 35 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.715
+ $X2=3.18 $Y2=0.715
r215 35 36 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.095 $Y=0.715
+ $X2=2.255 $Y2=0.715
r216 34 49 7.51051 $w=3.33e-07 $l=2.93094e-07 $layer=LI1_cond $X=1.395 $Y=0.955
+ $X2=1.187 $Y2=0.75
r217 33 56 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.045 $Y=0.955
+ $X2=2.15 $Y2=0.955
r218 33 34 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.045 $Y=0.955
+ $X2=1.395 $Y2=0.955
r219 31 34 5.34516 $w=3.33e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.3 $Y=1.04
+ $X2=1.395 $Y2=0.955
r220 31 52 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=1.3 $Y=1.04 $X2=1.3
+ $Y2=1.58
r221 28 53 6.0629 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=1.252 $Y=1.958
+ $X2=1.252 $Y2=2.1
r222 27 52 7.02549 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=1.252 $Y=1.722
+ $X2=1.252 $Y2=1.58
r223 27 28 9.54304 $w=2.83e-07 $l=2.36e-07 $layer=LI1_cond $X=1.252 $Y=1.722
+ $X2=1.252 $Y2=1.958
r224 23 51 6.50835 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=1.19 $Y=2.51
+ $X2=1.19 $Y2=2.35
r225 23 25 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=1.19 $Y=2.51
+ $X2=1.19 $Y2=2.515
r226 19 21 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=6.915 $Y=1.72
+ $X2=6.915 $Y2=2.57
r227 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.84 $Y=1.645
+ $X2=6.915 $Y2=1.72
r228 17 73 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.84 $Y=1.645
+ $X2=6.53 $Y2=1.645
r229 14 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.15 $Y=1.39
+ $X2=6.15 $Y2=1.555
r230 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.15 $Y=1.39
+ $X2=6.15 $Y2=0.96
r231 11 63 59.1843 $w=4.1e-07 $l=4.22137e-07 $layer=POLY_cond $X=3.735 $Y=1.45
+ $X2=3.525 $Y2=1.78
r232 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.735 $Y=1.45
+ $X2=3.735 $Y2=1.165
r233 7 63 39.7867 $w=4.1e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.44 $Y=1.945
+ $X2=3.525 $Y2=1.78
r234 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.44 $Y=1.945
+ $X2=3.44 $Y2=2.525
r235 2 25 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=2.36 $X2=1.125 $Y2=2.515
r236 1 49 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.54 $X2=1.145 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_804_328# 1 2 9 13 17 18 20 21 23 24 25 27
+ 30 33 37
c109 18 0 1.04851e-19 $X=4.185 $Y=1.805
c110 17 0 1.278e-20 $X=4.185 $Y=1.805
r111 33 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.935 $Y=1.155
+ $X2=5.935 $Y2=1.32
r112 28 37 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=6.037 $Y=2.07
+ $X2=6.037 $Y2=1.985
r113 28 30 36.1814 $w=2.13e-07 $l=6.75e-07 $layer=LI1_cond $X=6.037 $Y=2.07
+ $X2=6.037 $Y2=2.745
r114 27 37 4.65272 $w=1.92e-07 $l=9.53677e-08 $layer=LI1_cond $X=6.015 $Y=1.9
+ $X2=6.037 $Y2=1.985
r115 27 35 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.015 $Y=1.9
+ $X2=6.015 $Y2=1.32
r116 24 37 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.93 $Y=1.985
+ $X2=6.037 $Y2=1.985
r117 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.93 $Y=1.985
+ $X2=5.24 $Y2=1.985
r118 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.155 $Y=1.9
+ $X2=5.24 $Y2=1.985
r119 22 23 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.155 $Y=1.61
+ $X2=5.155 $Y2=1.9
r120 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.07 $Y=1.525
+ $X2=5.155 $Y2=1.61
r121 20 21 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=5.07 $Y=1.525
+ $X2=4.295 $Y2=1.525
r122 18 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.185 $Y=1.805
+ $X2=4.185 $Y2=1.97
r123 18 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.185 $Y=1.805
+ $X2=4.185 $Y2=1.64
r124 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.185
+ $Y=1.805 $X2=4.185 $Y2=1.805
r125 15 21 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=4.167 $Y=1.61
+ $X2=4.295 $Y2=1.525
r126 15 17 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=4.167 $Y=1.61
+ $X2=4.167 $Y2=1.805
r127 13 40 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.23 $Y=2.525
+ $X2=4.23 $Y2=1.97
r128 9 39 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.165 $Y=1.165
+ $X2=4.165 $Y2=1.64
r129 2 37 400 $w=1.7e-07 $l=3.08504e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.895 $X2=6.04 $Y2=2.065
r130 2 30 400 $w=1.7e-07 $l=9.60339e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.895 $X2=6.04 $Y2=2.745
r131 1 33 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.64 $X2=5.935 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%RESET_B 3 8 9 10 14 17 21 25 30 33 34 35 36
+ 37 45 48 49 51 52 59 60
c199 59 0 4.9151e-20 $X=7.905 $Y=2.035
c200 45 0 1.14348e-19 $X=7.92 $Y=2.035
c201 9 0 1.36523e-19 $X=4.56 $Y=0.54
r202 58 60 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.905 $Y=2.035
+ $X2=8.055 $Y2=2.035
r203 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.905
+ $Y=2.035 $X2=7.905 $Y2=2.035
r204 55 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.815 $Y=2.035
+ $X2=7.905 $Y2=2.035
r205 51 54 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=4.765 $Y=1.955
+ $X2=4.765 $Y2=2.12
r206 51 53 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=4.765 $Y=1.955
+ $X2=4.765 $Y2=1.79
r207 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.805
+ $Y=1.955 $X2=4.805 $Y2=1.955
r208 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.775
+ $Y=1.65 $X2=1.775 $Y2=1.65
r209 45 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r210 44 52 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=4.56 $Y=1.955
+ $X2=4.805 $Y2=1.955
r211 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.035
+ $X2=4.56 $Y2=2.035
r212 40 49 16.743 $w=2.63e-07 $l=3.85e-07 $layer=LI1_cond $X=1.727 $Y=2.035
+ $X2=1.727 $Y2=1.65
r213 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.035
r214 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.035
+ $X2=4.56 $Y2=2.035
r215 36 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r216 36 37 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.705 $Y2=2.035
r217 35 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=2.035
+ $X2=1.68 $Y2=2.035
r218 34 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=4.56 $Y2=2.035
r219 34 35 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=1.825 $Y2=2.035
r220 32 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.775 $Y=1.99
+ $X2=1.775 $Y2=1.65
r221 32 33 45.2978 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.99
+ $X2=1.775 $Y2=2.155
r222 28 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.775 $Y=1.635
+ $X2=1.775 $Y2=1.65
r223 28 30 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.775 $Y=1.56
+ $X2=2.04 $Y2=1.56
r224 23 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=2.2
+ $X2=8.055 $Y2=2.035
r225 23 25 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.055 $Y=2.2
+ $X2=8.055 $Y2=2.57
r226 19 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.815 $Y=1.87
+ $X2=7.815 $Y2=2.035
r227 19 21 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=7.815 $Y=1.87
+ $X2=7.815 $Y2=0.85
r228 17 54 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.78 $Y=2.525
+ $X2=4.78 $Y2=2.12
r229 14 53 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=4.635 $Y=1.165
+ $X2=4.635 $Y2=1.79
r230 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.635 $Y=0.615
+ $X2=4.635 $Y2=1.165
r231 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.56 $Y=0.54
+ $X2=4.635 $Y2=0.615
r232 9 10 1253.71 $w=1.5e-07 $l=2.445e-06 $layer=POLY_cond $X=4.56 $Y=0.54
+ $X2=2.115 $Y2=0.54
r233 6 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.04 $Y=1.485
+ $X2=2.04 $Y2=1.56
r234 6 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.04 $Y=1.485
+ $X2=2.04 $Y2=1.165
r235 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.04 $Y=0.615
+ $X2=2.115 $Y2=0.54
r236 5 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.04 $Y=0.615
+ $X2=2.04 $Y2=1.165
r237 3 33 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.86 $Y=2.525
+ $X2=1.86 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_603_191# 1 2 3 10 12 15 18 19 21 22 23 27
+ 34 38 47
c100 23 0 1.04851e-19 $X=5.41 $Y=1.16
c101 22 0 1.60894e-19 $X=3.965 $Y=2.385
r102 46 47 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.72 $Y=1.555
+ $X2=5.73 $Y2=1.555
r103 36 37 3.43032 $w=4.09e-07 $l=1.15e-07 $layer=LI1_cond $X=3.655 $Y=2.517
+ $X2=3.77 $Y2=2.517
r104 33 34 3.34173 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.77 $Y=1.135
+ $X2=3.86 $Y2=1.135
r105 31 33 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.52 $Y=1.135
+ $X2=3.77 $Y2=1.135
r106 28 46 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.505 $Y=1.555
+ $X2=5.72 $Y2=1.555
r107 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.505
+ $Y=1.555 $X2=5.505 $Y2=1.555
r108 25 27 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=5.505 $Y=1.26
+ $X2=5.505 $Y2=1.555
r109 23 25 6.82232 $w=2e-07 $l=1.39642e-07 $layer=LI1_cond $X=5.41 $Y=1.16
+ $X2=5.505 $Y2=1.26
r110 23 38 66.2682 $w=1.98e-07 $l=1.195e-06 $layer=LI1_cond $X=5.41 $Y=1.16
+ $X2=4.215 $Y2=1.16
r111 22 37 10.0903 $w=4.09e-07 $l=2.52517e-07 $layer=LI1_cond $X=3.965 $Y=2.385
+ $X2=3.77 $Y2=2.517
r112 21 42 6.82058 $w=2.43e-07 $l=1.45e-07 $layer=LI1_cond $X=4.972 $Y=2.385
+ $X2=4.972 $Y2=2.53
r113 21 22 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.85 $Y=2.385
+ $X2=3.965 $Y2=2.385
r114 19 38 6.88214 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=4.07 $Y=1.115
+ $X2=4.215 $Y2=1.115
r115 19 34 8.34528 $w=2.88e-07 $l=2.1e-07 $layer=LI1_cond $X=4.07 $Y=1.115
+ $X2=3.86 $Y2=1.115
r116 18 37 5.56675 $w=1.8e-07 $l=2.17e-07 $layer=LI1_cond $X=3.77 $Y=2.3
+ $X2=3.77 $Y2=2.517
r117 17 33 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.77 $Y=1.3
+ $X2=3.77 $Y2=1.135
r118 17 18 61.6162 $w=1.78e-07 $l=1e-06 $layer=LI1_cond $X=3.77 $Y=1.3 $X2=3.77
+ $Y2=2.3
r119 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=1.72
+ $X2=5.73 $Y2=1.555
r120 13 15 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.73 $Y=1.72
+ $X2=5.73 $Y2=2.315
r121 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.72 $Y=1.39
+ $X2=5.72 $Y2=1.555
r122 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.72 $Y=1.39
+ $X2=5.72 $Y2=0.96
r123 3 42 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=2.315 $X2=4.995 $Y2=2.53
r124 2 36 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=2.315 $X2=3.655 $Y2=2.535
r125 1 31 182 $w=1.7e-07 $l=5.88154e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.955 $X2=3.52 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_28_108# 1 2 10 14 15 16 17 18 20 23 25 29
+ 31 35 39 41 43 44 47 51 55 56 58
c151 23 0 1.60894e-19 $X=2.94 $Y=1.165
r152 56 61 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.952 $Y=1.235
+ $X2=0.952 $Y2=1.4
r153 56 60 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.952 $Y=1.235
+ $X2=0.952 $Y2=1.07
r154 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=1.235 $X2=0.93 $Y2=1.235
r155 53 58 0.94211 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.43 $Y=1.235
+ $X2=0.265 $Y2=1.235
r156 53 55 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.43 $Y=1.235
+ $X2=0.93 $Y2=1.235
r157 49 58 5.66538 $w=2.95e-07 $l=1.81659e-07 $layer=LI1_cond $X=0.23 $Y=1.4
+ $X2=0.265 $Y2=1.235
r158 49 51 49.4221 $w=2.58e-07 $l=1.115e-06 $layer=LI1_cond $X=0.23 $Y=1.4
+ $X2=0.23 $Y2=2.515
r159 45 58 5.66538 $w=2.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=1.07
+ $X2=0.265 $Y2=1.235
r160 45 47 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.265 $Y=1.07
+ $X2=0.265 $Y2=0.75
r161 41 42 49.1513 $w=1.52e-07 $l=1.55e-07 $layer=POLY_cond $X=0.91 $Y=2.202
+ $X2=1.065 $Y2=2.202
r162 37 39 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=7.025 $Y=0.255
+ $X2=7.025 $Y2=0.85
r163 33 35 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=6.39 $Y=3.075
+ $X2=6.39 $Y2=2.48
r164 32 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.945 $Y=3.15
+ $X2=3.87 $Y2=3.15
r165 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.315 $Y=3.15
+ $X2=6.39 $Y2=3.075
r166 31 32 1215.26 $w=1.5e-07 $l=2.37e-06 $layer=POLY_cond $X=6.315 $Y=3.15
+ $X2=3.945 $Y2=3.15
r167 27 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.87 $Y=3.075
+ $X2=3.87 $Y2=3.15
r168 27 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.87 $Y=3.075
+ $X2=3.87 $Y2=2.525
r169 26 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=3.15
+ $X2=2.94 $Y2=3.15
r170 25 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.795 $Y=3.15
+ $X2=3.87 $Y2=3.15
r171 25 26 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.795 $Y=3.15
+ $X2=3.015 $Y2=3.15
r172 21 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=3.075
+ $X2=2.94 $Y2=3.15
r173 21 23 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=2.94 $Y=3.075
+ $X2=2.94 $Y2=1.165
r174 20 42 3.14937 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=1.065 $Y=2.12
+ $X2=1.065 $Y2=2.202
r175 20 61 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.065 $Y=2.12
+ $X2=1.065 $Y2=1.4
r176 17 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=3.15
+ $X2=2.94 $Y2=3.15
r177 17 18 964 $w=1.5e-07 $l=1.88e-06 $layer=POLY_cond $X=2.865 $Y=3.15
+ $X2=0.985 $Y2=3.15
r178 15 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.95 $Y=0.18
+ $X2=7.025 $Y2=0.255
r179 15 16 3058.65 $w=1.5e-07 $l=5.965e-06 $layer=POLY_cond $X=6.95 $Y=0.18
+ $X2=0.985 $Y2=0.18
r180 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=3.075
+ $X2=0.985 $Y2=3.15
r181 12 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.91 $Y=3.075
+ $X2=0.91 $Y2=2.68
r182 11 41 3.14937 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=0.91 $Y=2.285
+ $X2=0.91 $Y2=2.202
r183 11 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.91 $Y=2.285
+ $X2=0.91 $Y2=2.68
r184 10 60 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.91 $Y=0.75
+ $X2=0.91 $Y2=1.07
r185 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.985 $Y2=0.18
r186 7 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.91 $Y2=0.75
r187 2 51 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=2.36 $X2=0.265 $Y2=2.515
r188 1 47 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.54 $X2=0.265 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_1440_304# 1 2 9 13 17 18 23 30 32 33 35 36
+ 39 40
c95 17 0 1.14348e-19 $X=7.365 $Y=2.025
c96 9 0 4.9151e-20 $X=7.275 $Y=2.57
r97 38 40 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.335 $Y=1.785
+ $X2=8.7 $Y2=1.785
r98 38 39 6.04704 $w=3.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=1.785
+ $X2=8.25 $Y2=1.785
r99 35 36 11.4521 $w=2.53e-07 $l=2.25e-07 $layer=LI1_cond $X=8.292 $Y=2.57
+ $X2=8.292 $Y2=2.345
r100 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.365
+ $Y=1.685 $X2=7.365 $Y2=1.685
r101 30 40 4.96451 $w=1.8e-07 $l=1.85e-07 $layer=LI1_cond $X=8.7 $Y=1.6 $X2=8.7
+ $Y2=1.785
r102 29 30 36.0455 $w=1.78e-07 $l=5.85e-07 $layer=LI1_cond $X=8.7 $Y=1.015
+ $X2=8.7 $Y2=1.6
r103 27 38 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.335 $Y=1.97
+ $X2=8.335 $Y2=1.785
r104 27 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.335 $Y=1.97
+ $X2=8.335 $Y2=2.345
r105 23 29 7.61292 $w=3.3e-07 $l=2.05122e-07 $layer=LI1_cond $X=8.61 $Y=0.85
+ $X2=8.7 $Y2=1.015
r106 23 25 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=8.61 $Y=0.85
+ $X2=8.39 $Y2=0.85
r107 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.53 $Y=1.685
+ $X2=7.365 $Y2=1.685
r108 22 39 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.53 $Y=1.685
+ $X2=8.25 $Y2=1.685
r109 17 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.365 $Y=2.025
+ $X2=7.365 $Y2=1.685
r110 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.365 $Y=2.025
+ $X2=7.365 $Y2=2.19
r111 16 33 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.365 $Y=1.52
+ $X2=7.365 $Y2=1.685
r112 13 16 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.385 $Y=0.85
+ $X2=7.385 $Y2=1.52
r113 9 18 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=7.275 $Y=2.57
+ $X2=7.275 $Y2=2.19
r114 2 35 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.13
+ $Y=2.36 $X2=8.27 $Y2=2.57
r115 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.25
+ $Y=0.64 $X2=8.39 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_1245_128# 1 2 7 9 12 16 20 24 28 31 32 33
+ 35 41 45 48 49 50 53 56 58 60 61 65 69 70 71 72 76 77 79 80 81 87 90
c201 90 0 9.16501e-20 $X=10.942 $Y=1.185
c202 16 0 1.83812e-19 $X=9.455 $Y=0.905
r203 80 91 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=10.942 $Y=1.35
+ $X2=10.942 $Y2=1.515
r204 80 90 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=10.942 $Y=1.35
+ $X2=10.942 $Y2=1.185
r205 79 81 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=10.92 $Y=1.35
+ $X2=10.92 $Y2=1.185
r206 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.93
+ $Y=1.35 $X2=10.93 $Y2=1.35
r207 72 74 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=9.045 $Y=0.43
+ $X2=9.045 $Y2=0.71
r208 67 81 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.91 $Y=0.795
+ $X2=10.91 $Y2=1.185
r209 66 77 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.64 $Y=0.71 $X2=9.55
+ $Y2=0.71
r210 65 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.825 $Y=0.71
+ $X2=10.91 $Y2=0.795
r211 65 66 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=10.825 $Y=0.71
+ $X2=9.64 $Y2=0.71
r212 63 77 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.55 $Y=0.795
+ $X2=9.55 $Y2=0.71
r213 63 76 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=9.55 $Y=0.795
+ $X2=9.55 $Y2=1.325
r214 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.43
+ $Y=1.49 $X2=9.43 $Y2=1.49
r215 58 76 7.48172 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=9.492 $Y=1.472
+ $X2=9.492 $Y2=1.325
r216 58 60 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=9.492 $Y=1.472
+ $X2=9.492 $Y2=1.49
r217 57 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.13 $Y=0.71
+ $X2=9.045 $Y2=0.71
r218 56 77 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.46 $Y=0.71 $X2=9.55
+ $Y2=0.71
r219 56 57 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.46 $Y=0.71
+ $X2=9.13 $Y2=0.71
r220 54 87 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=8.265 $Y=1.335
+ $X2=8.485 $Y2=1.335
r221 54 84 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.265 $Y=1.335
+ $X2=8.175 $Y2=1.335
r222 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.265
+ $Y=1.335 $X2=8.265 $Y2=1.335
r223 51 71 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.045 $Y=1.31
+ $X2=7.96 $Y2=1.31
r224 51 53 10.5641 $w=2.38e-07 $l=2.2e-07 $layer=LI1_cond $X=8.045 $Y=1.31
+ $X2=8.265 $Y2=1.31
r225 49 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=0.43
+ $X2=9.045 $Y2=0.43
r226 49 50 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=8.96 $Y=0.43
+ $X2=8.045 $Y2=0.43
r227 48 71 2.11342 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.96 $Y=1.19
+ $X2=7.96 $Y2=1.31
r228 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.96 $Y=0.515
+ $X2=8.045 $Y2=0.43
r229 47 48 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.96 $Y=0.515
+ $X2=7.96 $Y2=1.19
r230 46 70 1.72457 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=6.82 $Y=1.34 $X2=6.72
+ $Y2=1.34
r231 45 71 4.3182 $w=2.1e-07 $l=9.88686e-08 $layer=LI1_cond $X=7.875 $Y=1.34
+ $X2=7.96 $Y2=1.31
r232 45 46 65.0051 $w=1.78e-07 $l=1.055e-06 $layer=LI1_cond $X=7.875 $Y=1.34
+ $X2=6.82 $Y2=1.34
r233 43 70 4.72821 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=6.72 $Y=1.43 $X2=6.72
+ $Y2=1.34
r234 43 69 33.8273 $w=1.98e-07 $l=6.1e-07 $layer=LI1_cond $X=6.72 $Y=1.43
+ $X2=6.72 $Y2=2.04
r235 39 70 4.72821 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=6.72 $Y=1.25 $X2=6.72
+ $Y2=1.34
r236 39 41 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=6.72 $Y=1.25
+ $X2=6.72 $Y2=0.795
r237 35 37 19.6275 $w=3.18e-07 $l=5.45e-07 $layer=LI1_cond $X=6.66 $Y=2.205
+ $X2=6.66 $Y2=2.75
r238 33 69 7.37399 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=6.66 $Y=2.2
+ $X2=6.66 $Y2=2.04
r239 33 35 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=6.66 $Y=2.2 $X2=6.66
+ $Y2=2.205
r240 31 61 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.43 $Y=1.83
+ $X2=9.43 $Y2=1.49
r241 31 32 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.43 $Y=1.83
+ $X2=9.43 $Y2=1.995
r242 30 61 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.43 $Y=1.325
+ $X2=9.43 $Y2=1.49
r243 28 90 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.045 $Y=0.655
+ $X2=11.045 $Y2=1.185
r244 24 91 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=10.965 $Y=2.465
+ $X2=10.965 $Y2=1.515
r245 20 32 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.455 $Y=2.755
+ $X2=9.455 $Y2=1.995
r246 16 30 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=9.455 $Y=0.905
+ $X2=9.455 $Y2=1.325
r247 10 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.485 $Y=1.5
+ $X2=8.485 $Y2=1.335
r248 10 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=8.485 $Y=1.5
+ $X2=8.485 $Y2=2.57
r249 7 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.175 $Y=1.17
+ $X2=8.175 $Y2=1.335
r250 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.175 $Y=1.17
+ $X2=8.175 $Y2=0.85
r251 2 37 600 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=2.06 $X2=6.605 $Y2=2.75
r252 2 35 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=2.06 $X2=6.605 $Y2=2.205
r253 1 41 91 $w=1.7e-07 $l=5.52087e-07 $layer=licon1_NDIFF $count=2 $X=6.225
+ $Y=0.64 $X2=6.705 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_1796_139# 1 2 9 11 15 17 18 21 23 26 29 31
+ 32
r83 32 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.97 $Y=1.51 $X2=9.97
+ $Y2=1.6
r84 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.97 $Y=1.51
+ $X2=9.97 $Y2=1.345
r85 31 34 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=9.942 $Y=1.51
+ $X2=9.942 $Y2=1.675
r86 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.97
+ $Y=1.51 $X2=9.97 $Y2=1.51
r87 26 34 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=9.915 $Y=2.165
+ $X2=9.915 $Y2=1.675
r88 24 29 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.325 $Y=2.25
+ $X2=9.16 $Y2=2.25
r89 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.83 $Y=2.25
+ $X2=9.915 $Y2=2.165
r90 23 24 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=9.83 $Y=2.25
+ $X2=9.325 $Y2=2.25
r91 19 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.16 $Y=2.335
+ $X2=9.16 $Y2=2.25
r92 19 21 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=9.16 $Y=2.335
+ $X2=9.16 $Y2=2.56
r93 18 29 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=9.08 $Y=2.165
+ $X2=9.16 $Y2=2.25
r94 17 28 10.1209 $w=2.83e-07 $l=2.11305e-07 $layer=LI1_cond $X=9.08 $Y=1.25
+ $X2=9.125 $Y2=1.06
r95 17 18 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=9.08 $Y=1.25
+ $X2=9.08 $Y2=2.165
r96 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.48 $Y=1.675
+ $X2=10.48 $Y2=2.465
r97 12 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.135 $Y=1.6
+ $X2=9.97 $Y2=1.6
r98 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.405 $Y=1.6
+ $X2=10.48 $Y2=1.675
r99 11 12 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.405 $Y=1.6
+ $X2=10.135 $Y2=1.6
r100 9 36 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.04 $Y=0.765
+ $X2=10.04 $Y2=1.345
r101 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.095
+ $Y=2.435 $X2=9.24 $Y2=2.56
r102 1 28 182 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_NDIFF $count=1 $X=8.98
+ $Y=0.695 $X2=9.125 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 55
+ 60 61 63 64 66 67 68 70 75 80 88 93 112 113 116 119 122 125 128
r142 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r143 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r144 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r145 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r146 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r148 110 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r149 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r150 107 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r151 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r152 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r153 104 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 101 128 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.995 $Y=3.33
+ $X2=7.66 $Y2=3.33
r156 101 103 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.995 $Y=3.33
+ $X2=8.4 $Y2=3.33
r157 100 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r158 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r159 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r160 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r161 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r162 94 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=3.33
+ $X2=5.515 $Y2=3.33
r163 94 96 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.68 $Y=3.33 $X2=6
+ $Y2=3.33
r164 93 128 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.325 $Y=3.33
+ $X2=7.66 $Y2=3.33
r165 93 99 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.325 $Y=3.33
+ $X2=6.96 $Y2=3.33
r166 92 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r167 92 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r168 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r169 89 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.505 $Y2=3.33
r170 89 91 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=5.04 $Y2=3.33
r171 88 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=3.33
+ $X2=5.515 $Y2=3.33
r172 88 91 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.35 $Y=3.33
+ $X2=5.04 $Y2=3.33
r173 87 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r174 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 84 87 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r176 84 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r177 83 86 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r178 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r179 81 119 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.145 $Y2=3.33
r180 81 83 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.64 $Y2=3.33
r181 80 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.34 $Y=3.33
+ $X2=4.505 $Y2=3.33
r182 80 86 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.34 $Y=3.33
+ $X2=4.08 $Y2=3.33
r183 79 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r184 79 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r185 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r186 76 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=3.33
+ $X2=0.695 $Y2=3.33
r187 76 78 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.86 $Y=3.33
+ $X2=1.68 $Y2=3.33
r188 75 119 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=2.145 $Y2=3.33
r189 75 78 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 73 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r191 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r192 70 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.695 $Y2=3.33
r193 70 72 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.24 $Y2=3.33
r194 68 97 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r195 68 126 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r196 66 109 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.6 $Y=3.33
+ $X2=10.32 $Y2=3.33
r197 66 67 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=10.6 $Y=3.33
+ $X2=10.732 $Y2=3.33
r198 65 112 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=11.28 $Y2=3.33
r199 65 67 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=10.732 $Y2=3.33
r200 63 106 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=9.505 $Y=3.33
+ $X2=9.36 $Y2=3.33
r201 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.505 $Y=3.33
+ $X2=9.67 $Y2=3.33
r202 62 109 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=9.835 $Y=3.33
+ $X2=10.32 $Y2=3.33
r203 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.835 $Y=3.33
+ $X2=9.67 $Y2=3.33
r204 60 103 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=8.59 $Y=3.33
+ $X2=8.4 $Y2=3.33
r205 60 61 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=8.59 $Y=3.33
+ $X2=8.707 $Y2=3.33
r206 59 106 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.825 $Y=3.33
+ $X2=9.36 $Y2=3.33
r207 59 61 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=8.825 $Y=3.33
+ $X2=8.707 $Y2=3.33
r208 55 58 41.9663 $w=2.63e-07 $l=9.65e-07 $layer=LI1_cond $X=10.732 $Y=1.985
+ $X2=10.732 $Y2=2.95
r209 53 67 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=10.732 $Y=3.245
+ $X2=10.732 $Y2=3.33
r210 53 58 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=10.732 $Y=3.245
+ $X2=10.732 $Y2=2.95
r211 49 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=3.245
+ $X2=9.67 $Y2=3.33
r212 49 51 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=9.67 $Y=3.245
+ $X2=9.67 $Y2=2.59
r213 45 61 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.707 $Y=3.245
+ $X2=8.707 $Y2=3.33
r214 45 47 33.1021 $w=2.33e-07 $l=6.75e-07 $layer=LI1_cond $X=8.707 $Y=3.245
+ $X2=8.707 $Y2=2.57
r215 41 128 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.66 $Y=3.245
+ $X2=7.66 $Y2=3.33
r216 41 43 12.05 $w=6.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.66 $Y=3.245
+ $X2=7.66 $Y2=2.57
r217 37 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=3.245
+ $X2=5.515 $Y2=3.33
r218 37 39 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=5.515 $Y=3.245
+ $X2=5.515 $Y2=2.405
r219 33 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.505 $Y=3.245
+ $X2=4.505 $Y2=3.33
r220 33 35 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.505 $Y=3.245
+ $X2=4.505 $Y2=2.75
r221 29 119 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=3.245
+ $X2=2.145 $Y2=3.33
r222 29 31 16.2988 $w=3.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.145 $Y=3.245
+ $X2=2.145 $Y2=2.75
r223 25 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r224 25 27 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.515
r225 8 58 400 $w=1.7e-07 $l=1.19931e-06 $layer=licon1_PDIFF $count=1 $X=10.555
+ $Y=1.835 $X2=10.73 $Y2=2.95
r226 8 55 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=10.555
+ $Y=1.835 $X2=10.73 $Y2=1.985
r227 7 51 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=9.53
+ $Y=2.435 $X2=9.67 $Y2=2.59
r228 6 47 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=2.36 $X2=8.7 $Y2=2.57
r229 5 43 300 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_PDIFF $count=2 $X=7.35
+ $Y=2.36 $X2=7.84 $Y2=2.57
r230 4 39 600 $w=1.7e-07 $l=5.69078e-07 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.895 $X2=5.515 $Y2=2.405
r231 3 35 600 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=2.315 $X2=4.505 $Y2=2.75
r232 2 31 600 $w=1.7e-07 $l=5.29693e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=2.315 $X2=2.145 $Y2=2.75
r233 1 27 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=2.36 $X2=0.695 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%A_304_463# 1 2 3 4 13 16 19 24 28
r50 28 30 9.0501 $w=5.19e-07 $l=3.85e-07 $layer=LI1_cond $X=2.84 $Y=2.425
+ $X2=3.225 $Y2=2.425
r51 27 28 4.58382 $w=5.19e-07 $l=1.95e-07 $layer=LI1_cond $X=2.645 $Y=2.425
+ $X2=2.84 $Y2=2.425
r52 22 24 7.92305 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=1.1
+ $X2=2.84 $Y2=1.1
r53 16 28 7.39147 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=2.84 $Y=2.115
+ $X2=2.84 $Y2=2.425
r54 15 24 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.84 $Y=1.22 $X2=2.84
+ $Y2=1.1
r55 15 16 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.84 $Y=1.22
+ $X2=2.84 $Y2=2.115
r56 14 19 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.73 $Y=2.41
+ $X2=1.625 $Y2=2.41
r57 13 27 8.41732 $w=5.19e-07 $l=1.1225e-07 $layer=LI1_cond $X=2.54 $Y=2.41
+ $X2=2.645 $Y2=2.425
r58 13 14 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.54 $Y=2.41
+ $X2=1.73 $Y2=2.41
r59 4 30 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=2.315 $X2=3.225 $Y2=2.52
r60 3 27 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=2.315 $X2=2.645 $Y2=2.52
r61 2 19 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=2.315 $X2=1.645 $Y2=2.49
r62 1 22 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.955 $X2=2.675 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%Q 1 2 10 13 14 15 16 17 32
c31 13 0 9.16501e-20 $X=10.32 $Y=1.295
c32 10 0 1.83812e-19 $X=10.327 $Y=1.065
r33 29 32 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=10.3 $Y=1.975
+ $X2=10.3 $Y2=2.02
r34 17 39 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=10.3 $Y=2.775
+ $X2=10.3 $Y2=2.91
r35 16 17 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=10.3 $Y=2.405
+ $X2=10.3 $Y2=2.775
r36 15 29 0.576222 $w=2.58e-07 $l=1.3e-08 $layer=LI1_cond $X=10.3 $Y=1.962
+ $X2=10.3 $Y2=1.975
r37 15 42 5.73379 $w=2.58e-07 $l=1.17e-07 $layer=LI1_cond $X=10.3 $Y=1.962
+ $X2=10.3 $Y2=1.845
r38 15 16 15.8683 $w=2.58e-07 $l=3.58e-07 $layer=LI1_cond $X=10.3 $Y=2.047
+ $X2=10.3 $Y2=2.405
r39 15 32 1.19677 $w=2.58e-07 $l=2.7e-08 $layer=LI1_cond $X=10.3 $Y=2.047
+ $X2=10.3 $Y2=2.02
r40 14 42 9.73836 $w=2.03e-07 $l=1.8e-07 $layer=LI1_cond $X=10.327 $Y=1.665
+ $X2=10.327 $Y2=1.845
r41 13 14 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=10.327 $Y=1.295
+ $X2=10.327 $Y2=1.665
r42 11 13 7.03326 $w=2.03e-07 $l=1.3e-07 $layer=LI1_cond $X=10.327 $Y=1.165
+ $X2=10.327 $Y2=1.295
r43 10 11 0.595843 $w=2.05e-07 $l=1e-07 $layer=LI1_cond $X=10.327 $Y=1.065
+ $X2=10.327 $Y2=1.165
r44 8 10 3.99273 $w=1.98e-07 $l=7.2e-08 $layer=LI1_cond $X=10.255 $Y=1.065
+ $X2=10.327 $Y2=1.065
r45 2 39 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.835 $X2=10.265 $Y2=2.91
r46 2 32 400 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.835 $X2=10.265 $Y2=2.02
r47 1 8 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=10.115
+ $Y=0.345 $X2=10.255 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%Q_N 1 2 7 8 9 10 11 12 13 25 31 40
r22 38 40 0.432166 $w=3.98e-07 $l=1.5e-08 $layer=LI1_cond $X=11.235 $Y=2.02
+ $X2=11.235 $Y2=2.035
r23 23 31 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=11.3 $Y=0.96
+ $X2=11.3 $Y2=0.925
r24 13 47 3.8895 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=11.235 $Y=2.775
+ $X2=11.235 $Y2=2.91
r25 12 13 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=11.235 $Y=2.405
+ $X2=11.235 $Y2=2.775
r26 11 38 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=11.235 $Y=1.985
+ $X2=11.235 $Y2=2.02
r27 11 53 6.36561 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=11.235 $Y=1.985
+ $X2=11.235 $Y2=1.82
r28 11 12 9.65171 $w=3.98e-07 $l=3.35e-07 $layer=LI1_cond $X=11.235 $Y=2.07
+ $X2=11.235 $Y2=2.405
r29 11 40 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=11.235 $Y=2.07
+ $X2=11.235 $Y2=2.035
r30 10 53 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=11.31 $Y=1.665
+ $X2=11.31 $Y2=1.82
r31 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=11.31 $Y=1.295
+ $X2=11.31 $Y2=1.665
r32 9 50 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=11.31 $Y=1.295
+ $X2=11.31 $Y2=1.095
r33 8 50 4.77682 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=11.3 $Y=0.985
+ $X2=11.3 $Y2=1.095
r34 8 23 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=11.3 $Y=0.985
+ $X2=11.3 $Y2=0.96
r35 8 31 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=11.3 $Y=0.9 $X2=11.3
+ $Y2=0.925
r36 7 8 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.3 $Y=0.555
+ $X2=11.3 $Y2=0.9
r37 7 25 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=11.3 $Y=0.555
+ $X2=11.3 $Y2=0.42
r38 2 11 400 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=11.04
+ $Y=1.835 $X2=11.2 $Y2=1.985
r39 2 47 400 $w=1.7e-07 $l=1.15223e-06 $layer=licon1_PDIFF $count=1 $X=11.04
+ $Y=1.835 $X2=11.2 $Y2=2.91
r40 1 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=11.12
+ $Y=0.235 $X2=11.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45 46
+ 48 53 58 70 77 84 85 88 91 94 97 100
r109 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r110 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r111 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r112 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r113 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r114 85 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r115 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r116 82 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.995 $Y=0
+ $X2=10.83 $Y2=0
r117 82 84 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.995 $Y=0
+ $X2=11.28 $Y2=0
r118 81 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r119 81 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r120 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r121 78 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.93 $Y=0 $X2=9.765
+ $Y2=0
r122 78 80 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.93 $Y=0 $X2=10.32
+ $Y2=0
r123 77 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=10.83 $Y2=0
r124 77 80 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=10.32 $Y2=0
r125 76 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r126 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r127 73 76 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.36 $Y2=0
r128 72 75 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.36
+ $Y2=0
r129 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r130 70 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.6 $Y=0 $X2=9.765
+ $Y2=0
r131 70 75 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.6 $Y=0 $X2=9.36
+ $Y2=0
r132 69 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r133 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r134 66 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.555 $Y=0 $X2=5.39
+ $Y2=0
r135 66 68 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=5.555 $Y=0
+ $X2=7.44 $Y2=0
r136 65 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r137 64 65 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r138 62 65 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=5.04 $Y2=0
r139 62 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r140 61 64 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=5.04
+ $Y2=0
r141 61 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r142 59 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r143 59 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.16 $Y2=0
r144 58 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.39
+ $Y2=0
r145 58 64 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.04 $Y2=0
r146 57 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r147 57 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r148 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r149 54 88 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.705
+ $Y2=0
r150 54 56 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=1.2
+ $Y2=0
r151 53 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r152 53 56 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r153 51 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r154 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r155 48 88 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.705
+ $Y2=0
r156 48 50 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.24
+ $Y2=0
r157 46 69 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r158 46 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r159 44 68 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.495 $Y=0 $X2=7.44
+ $Y2=0
r160 44 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.495 $Y=0 $X2=7.59
+ $Y2=0
r161 43 72 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.685 $Y=0
+ $X2=7.92 $Y2=0
r162 43 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.685 $Y=0 $X2=7.59
+ $Y2=0
r163 39 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.83 $Y=0.085
+ $X2=10.83 $Y2=0
r164 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=10.83 $Y=0.085
+ $X2=10.83 $Y2=0.36
r165 35 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.765 $Y=0.085
+ $X2=9.765 $Y2=0
r166 35 37 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.765 $Y=0.085
+ $X2=9.765 $Y2=0.36
r167 31 45 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=0.085
+ $X2=7.59 $Y2=0
r168 31 33 40.8612 $w=1.88e-07 $l=7e-07 $layer=LI1_cond $X=7.59 $Y=0.085
+ $X2=7.59 $Y2=0.785
r169 27 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.39 $Y=0.085
+ $X2=5.39 $Y2=0
r170 27 29 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.39 $Y=0.085
+ $X2=5.39 $Y2=0.455
r171 23 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r172 23 25 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.59
r173 19 88 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r174 19 21 34.329 $w=2.08e-07 $l=6.5e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.735
r175 6 41 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=10.685
+ $Y=0.235 $X2=10.83 $Y2=0.36
r176 5 37 182 $w=1.7e-07 $l=4.36978e-07 $layer=licon1_NDIFF $count=1 $X=9.53
+ $Y=0.695 $X2=9.765 $Y2=0.36
r177 4 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.64 $X2=7.6 $Y2=0.785
r178 3 29 182 $w=1.7e-07 $l=8.95768e-07 $layer=licon1_NDIFF $count=1 $X=4.71
+ $Y=0.955 $X2=5.39 $Y2=0.455
r179 2 25 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.43 $X2=1.71 $Y2=0.59
r180 1 21 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.54 $X2=0.695 $Y2=0.735
.ends

