* File: sky130_fd_sc_lp__dfxtp_4.spice
* Created: Fri Aug 28 10:24:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfxtp_4.pex.spice"
.subckt sky130_fd_sc_lp__dfxtp_4  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1004 N_A_110_70#_M1004_d N_CLK_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_110_70#_M1011_g N_A_217_413#_M1011_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1019 N_A_431_119#_M1019_d N_D_M1019_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0819 PD=0.8 PS=0.81 NRD=25.704 NRS=14.28 M=1 R=2.8 SA=75000.7
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_526_413#_M1000_d N_A_110_70#_M1000_g N_A_431_119#_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.07875 AS=0.0798 PD=0.795 PS=0.8 NRD=17.136 NRS=2.856 M=1
+ R=2.8 SA=75001.3 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1005 A_642_119# N_A_217_413#_M1005_g N_A_526_413#_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.07875 PD=0.63 PS=0.795 NRD=14.28 NRS=9.996 M=1 R=2.8
+ SA=75001.8 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_684_93#_M1001_g A_642_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.119621 AS=0.0441 PD=0.966792 PS=0.63 NRD=45.708 NRS=14.28 M=1 R=2.8
+ SA=75002.1 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1016 N_A_684_93#_M1016_d N_A_526_413#_M1016_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.64 AD=0.135185 AS=0.182279 PD=1.24981 PS=1.47321 NRD=2.808 NRS=26.244 M=1
+ R=4.26667 SA=75002 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1007 N_A_941_379#_M1007_d N_A_217_413#_M1007_g N_A_684_93#_M1016_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.07455 AS=0.0887151 PD=0.775 PS=0.820189 NRD=21.42 NRS=28.56
+ M=1 R=2.8 SA=75003.4 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1017 A_1070_119# N_A_110_70#_M1017_g N_A_941_379#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.07455 PD=0.63 PS=0.775 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75003.9 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1112_93#_M1010_g A_1070_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1071 AS=0.0441 PD=0.853333 PS=0.63 NRD=28.56 NRS=14.28 M=1 R=2.8
+ SA=75004.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1026 N_A_1112_93#_M1026_d N_A_941_379#_M1026_g N_VGND_M1010_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.2142 PD=2.25 PS=1.70667 NRD=2.856 NRS=8.568 M=1
+ R=5.6 SA=75002.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_Q_M1013_d N_A_1112_93#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1014 N_Q_M1013_d N_A_1112_93#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1020 N_Q_M1020_d N_A_1112_93#_M1020_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1029 N_Q_M1020_d N_A_1112_93#_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1023 N_A_110_70#_M1023_d N_CLK_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VPWR_M1015_d N_A_110_70#_M1015_g N_A_217_413#_M1015_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.174672 AS=0.1696 PD=1.43698 PS=1.81 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1027 N_A_431_119#_M1027_d N_D_M1027_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.114628 PD=0.7 PS=0.943019 NRD=0 NRS=102.204 M=1 R=2.8
+ SA=75000.9 SB=75004 A=0.063 P=1.14 MULT=1
MM1008 N_A_526_413#_M1008_d N_A_217_413#_M1008_g N_A_431_119#_M1027_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=0.97 PS=0.7 NRD=121.943 NRS=0 M=1
+ R=2.8 SA=75001.3 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1022 A_666_413# N_A_110_70#_M1022_g N_A_526_413#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1155 PD=0.63 PS=0.97 NRD=23.443 NRS=4.6886 M=1 R=2.8
+ SA=75002 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_684_93#_M1024_g A_666_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.117233 AS=0.0441 PD=0.936667 PS=0.63 NRD=105.119 NRS=23.443 M=1 R=2.8
+ SA=75002.4 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1003 N_A_684_93#_M1003_d N_A_526_413#_M1003_g N_VPWR_M1024_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.234467 PD=1.12 PS=1.87333 NRD=0 NRS=15.2281 M=1
+ R=5.6 SA=75001.6 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1021 N_A_941_379#_M1021_d N_A_110_70#_M1021_g N_A_684_93#_M1003_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.337483 AS=0.1176 PD=2.08667 PS=1.12 NRD=82.0702 NRS=0 M=1
+ R=5.6 SA=75002 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1006 A_1116_441# N_A_217_413#_M1006_g N_A_941_379#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.168742 PD=0.63 PS=1.04333 NRD=23.443 NRS=45.7237 M=1
+ R=2.8 SA=75003.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_1112_93#_M1012_g A_1116_441# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0441 PD=0.8175 PS=0.63 NRD=45.7237 NRS=23.443 M=1 R=2.8
+ SA=75003.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1028 N_A_1112_93#_M1028_d N_A_941_379#_M1028_g N_VPWR_M1012_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_1112_93#_M1002_g N_Q_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_1112_93#_M1009_g N_Q_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1009_d N_A_1112_93#_M1018_g N_Q_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_A_1112_93#_M1025_g N_Q_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX30_noxref VNB VPB NWDIODE A=17.8319 P=22.95
c_100 VNB 0 4.11139e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfxtp_4.pxi.spice"
*
.ends
*
*
