* File: sky130_fd_sc_lp__xnor2_4.spice
* Created: Fri Aug 28 11:35:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor2_4.pex.spice"
.subckt sky130_fd_sc_lp__xnor2_4  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_A_31_65#_M1006_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1512 PD=2.25 PS=1.2 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.2
+ SB=75005.2 A=0.126 P=1.98 MULT=1
MM1017 N_A_31_65#_M1017_d N_A_M1017_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=1.428 M=1 R=5.6 SA=75000.7
+ SB=75004.7 A=0.126 P=1.98 MULT=1
MM1024 N_A_31_65#_M1017_d N_A_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1000 N_A_31_65#_M1000_d N_B_M1000_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1003 N_A_31_65#_M1000_d N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75003.4
+ A=0.126 P=1.98 MULT=1
MM1011 N_A_31_65#_M1011_d N_B_M1011_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4 SB=75003
+ A=0.126 P=1.98 MULT=1
MM1023 N_A_31_65#_M1011_d N_B_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9 SB=75002.6
+ A=0.126 P=1.98 MULT=1
MM1027 N_A_31_65#_M1027_d N_A_M1027_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75003.4
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_A_808_39#_M1001_g N_A_31_65#_M1027_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.8
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1001_d N_A_808_39#_M1009_g N_A_31_65#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1218 PD=1.12 PS=1.13 NRD=0 NRS=1.428 M=1 R=5.6
+ SA=75004.2 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1010 N_Y_M1010_d N_A_808_39#_M1010_g N_A_31_65#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1218 PD=1.19 PS=1.13 NRD=9.996 NRS=0 M=1 R=5.6 SA=75004.7
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1029 N_Y_M1010_d N_A_808_39#_M1029_g N_A_31_65#_M1029_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.2898 PD=1.19 PS=2.37 NRD=0 NRS=9.996 M=1 R=5.6 SA=75005.2
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_1235_65#_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.2226 PD=1.2 PS=2.21 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1030 N_VGND_M1018_d N_A_M1030_g N_A_1235_65#_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=1.428 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1032 N_VGND_M1032_d N_A_M1032_g N_A_1235_65#_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1034 N_VGND_M1032_d N_A_M1034_g N_A_1235_65#_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1004 N_A_808_39#_M1004_d N_B_M1004_g N_A_1235_65#_M1034_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1015 N_A_808_39#_M1004_d N_B_M1015_g N_A_1235_65#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1025 N_A_808_39#_M1025_d N_B_M1025_g N_A_1235_65#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1028 N_A_808_39#_M1025_d N_B_M1028_g N_A_1235_65#_M1028_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1019 N_VPWR_M1019_d N_A_M1019_g N_A_110_367#_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75009.3 A=0.189 P=2.82 MULT=1
MM1031 N_VPWR_M1031_d N_A_M1031_g N_A_110_367#_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.290975 AS=0.1764 PD=1.795 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75008.9 A=0.189 P=2.82 MULT=1
MM1036 N_VPWR_M1031_d N_A_M1036_g N_A_110_367#_M1036_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.290975 AS=0.1764 PD=1.795 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4 SA=75001.2
+ SB=75008.3 A=0.189 P=2.82 MULT=1
MM1002 N_A_110_367#_M1036_s N_B_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75007.8 A=0.189 P=2.82 MULT=1
MM1012 N_A_110_367#_M1012_d N_B_M1012_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75007.4 A=0.189 P=2.82 MULT=1
MM1013 N_A_110_367#_M1012_d N_B_M1013_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5 SB=75007
+ A=0.189 P=2.82 MULT=1
MM1022 N_A_110_367#_M1022_d N_B_M1022_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75006.5 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1037_d N_A_M1037_g N_A_110_367#_M1022_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75006.1 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1037_d N_A_808_39#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1020 N_VPWR_M1020_d N_A_808_39#_M1020_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.63315 AS=0.1764 PD=2.265 PS=1.54 NRD=21.8867 NRS=0 M=1 R=8.4 SA=75004.3
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1033 N_VPWR_M1020_d N_A_808_39#_M1033_g N_Y_M1033_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.63315 AS=0.1764 PD=2.265 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1038 N_VPWR_M1038_d N_A_808_39#_M1038_g N_Y_M1033_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1038_d N_A_M1008_g N_A_808_39#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.3
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_808_39#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.7
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1014_d N_A_M1026_g N_A_808_39#_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1039 N_VPWR_M1039_d N_A_M1039_g N_A_808_39#_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_A_808_39#_M1007_d N_B_M1007_g N_VPWR_M1039_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008 SB=75001.5
+ A=0.189 P=2.82 MULT=1
MM1016 N_A_808_39#_M1007_d N_B_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1021 N_A_808_39#_M1021_d N_B_M1021_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1035 N_A_808_39#_M1021_d N_B_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75009.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.5079 P=24.65
*
.include "sky130_fd_sc_lp__xnor2_4.pxi.spice"
*
.ends
*
*
