* File: sky130_fd_sc_lp__nand4bb_lp.pex.spice
* Created: Wed Sep  2 10:07:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%A_N 3 7 11 15 16 17 20 21
c44 7 0 1.06129e-19 $X=0.725 $Y=2.595
r45 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.02 $X2=0.63 $Y2=1.02
r46 17 21 8.56545 $w=3.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.02
r47 16 20 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=0.607 $Y=1.338
+ $X2=0.607 $Y2=1.02
r48 15 20 5.19077 $w=3.75e-07 $l=3.5e-08 $layer=POLY_cond $X=0.607 $Y=0.985
+ $X2=0.607 $Y2=1.02
r49 5 16 46.4148 $w=3.24e-07 $l=3.66279e-07 $layer=POLY_cond $X=0.725 $Y=1.65
+ $X2=0.607 $Y2=1.338
r50 5 7 234.789 $w=2.5e-07 $l=9.45e-07 $layer=POLY_cond $X=0.725 $Y=1.65
+ $X2=0.725 $Y2=2.595
r51 1 15 24.6308 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=0.835
+ $X2=0.675 $Y2=0.985
r52 1 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.855 $Y=0.835
+ $X2=0.855 $Y2=0.445
r53 1 3 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.495 $Y=0.835
+ $X2=0.495 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%A_27_47# 1 2 7 9 13 14 15 17 19 20 22 25
+ 27 31 32 35 38
c81 27 0 1.85715e-19 $X=1.09 $Y=1.81
r82 35 37 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.28 $Y=0.47
+ $X2=0.28 $Y2=0.675
r83 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.255
+ $Y=1.39 $X2=1.255 $Y2=1.39
r84 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.255 $Y=1.725
+ $X2=1.255 $Y2=1.39
r85 28 38 3.9231 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.625 $Y=1.81
+ $X2=0.37 $Y2=1.81
r86 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.09 $Y=1.81
+ $X2=1.255 $Y2=1.725
r87 27 28 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.09 $Y=1.81
+ $X2=0.625 $Y2=1.81
r88 23 38 2.80976 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.37 $Y=1.895
+ $X2=0.37 $Y2=1.81
r89 23 25 8.09112 $w=5.08e-07 $l=3.45e-07 $layer=LI1_cond $X=0.37 $Y=1.895
+ $X2=0.37 $Y2=2.24
r90 22 38 2.80976 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.2 $Y=1.725
+ $X2=0.37 $Y2=1.81
r91 22 37 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=0.2 $Y=1.725
+ $X2=0.2 $Y2=0.675
r92 20 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.255 $Y=1.73
+ $X2=1.255 $Y2=1.39
r93 19 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.255 $Y=1.225
+ $X2=1.255 $Y2=1.39
r94 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.845 $Y=0.73
+ $X2=1.845 $Y2=0.445
r95 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.77 $Y=0.805
+ $X2=1.845 $Y2=0.73
r96 13 14 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.77 $Y=0.805
+ $X2=1.42 $Y2=0.805
r97 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.345 $Y=0.88
+ $X2=1.42 $Y2=0.805
r98 11 19 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.345 $Y=0.88
+ $X2=1.345 $Y2=1.225
r99 7 20 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.255 $Y=1.895
+ $X2=1.255 $Y2=1.73
r100 7 9 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.255 $Y=1.895
+ $X2=1.255 $Y2=2.595
r101 2 25 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.315
+ $Y=2.095 $X2=0.46 $Y2=2.24
r102 1 35 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%A_332_352# 1 2 7 9 13 15 19 22 24 29 31
c74 7 0 3.05353e-19 $X=1.785 $Y=1.885
r75 31 33 9.16063 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.04 $Y=0.4
+ $X2=4.04 $Y2=0.585
r76 24 27 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.115 $Y=1.255
+ $X2=2.115 $Y2=1.35
r77 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.115
+ $Y=1.255 $X2=2.115 $Y2=1.255
r78 22 29 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.12 $Y=1.265
+ $X2=4.015 $Y2=1.35
r79 22 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.12 $Y=1.265
+ $X2=4.12 $Y2=0.585
r80 17 29 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=1.435
+ $X2=4.015 $Y2=1.35
r81 17 19 24.4136 $w=3.78e-07 $l=8.05e-07 $layer=LI1_cond $X=4.015 $Y=1.435
+ $X2=4.015 $Y2=2.24
r82 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=1.35
+ $X2=2.115 $Y2=1.35
r83 15 29 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.825 $Y=1.35
+ $X2=4.015 $Y2=1.35
r84 15 16 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=3.825 $Y=1.35
+ $X2=2.28 $Y2=1.35
r85 11 25 41.3402 $w=4.77e-07 $l=3.06594e-07 $layer=POLY_cond $X=2.205 $Y=1.09
+ $X2=1.97 $Y2=1.255
r86 11 13 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.205 $Y=1.09
+ $X2=2.205 $Y2=0.445
r87 7 25 74.5248 $w=4.77e-07 $l=7.16554e-07 $layer=POLY_cond $X=1.785 $Y=1.885
+ $X2=1.97 $Y2=1.255
r88 7 9 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.785 $Y=1.885
+ $X2=1.785 $Y2=2.595
r89 2 19 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.85
+ $Y=2.095 $X2=3.99 $Y2=2.24
r90 1 31 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.04 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%C 3 7 9 12 13
r42 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.77
+ $X2=2.655 $Y2=1.935
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.77
+ $X2=2.655 $Y2=1.605
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.77 $X2=2.655 $Y2=1.77
r45 9 13 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.655 $Y=2.035
+ $X2=2.655 $Y2=1.77
r46 7 14 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=2.595 $Y=0.445
+ $X2=2.595 $Y2=1.605
r47 3 15 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.625 $Y=2.595
+ $X2=2.625 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%D 1 3 8 12 14 17 18 19
r46 17 20 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.77
+ $X2=3.195 $Y2=1.935
r47 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.77
+ $X2=3.195 $Y2=1.605
r48 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=1.77 $X2=3.195 $Y2=1.77
r49 14 18 8.60274 $w=3.53e-07 $l=2.65e-07 $layer=LI1_cond $X=3.182 $Y=2.035
+ $X2=3.182 $Y2=1.77
r50 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.985 $Y=0.805
+ $X2=3.105 $Y2=0.805
r51 8 20 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.155 $Y=2.595
+ $X2=3.155 $Y2=1.935
r52 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=0.88
+ $X2=3.105 $Y2=0.805
r53 4 19 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=3.105 $Y=0.88
+ $X2=3.105 $Y2=1.605
r54 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.985 $Y=0.73
+ $X2=2.985 $Y2=0.805
r55 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.985 $Y=0.73 $X2=2.985
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%B_N 1 3 6 8 10 11 12 13 23
r40 22 23 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.725 $Y=0.93
+ $X2=3.825 $Y2=0.93
r41 20 22 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=3.555 $Y=0.93
+ $X2=3.725 $Y2=0.93
r42 17 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.465 $Y=0.93
+ $X2=3.555 $Y2=0.93
r43 13 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.555
+ $Y=0.93 $X2=3.555 $Y2=0.93
r44 12 13 15.666 $w=3.18e-07 $l=4.35e-07 $layer=LI1_cond $X=3.12 $Y=0.925
+ $X2=3.555 $Y2=0.925
r45 11 12 17.2866 $w=3.18e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0.925
+ $X2=3.12 $Y2=0.925
r46 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=0.765
+ $X2=3.825 $Y2=0.93
r47 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.825 $Y=0.765
+ $X2=3.825 $Y2=0.445
r48 4 22 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.725 $Y=1.095
+ $X2=3.725 $Y2=0.93
r49 4 6 372.68 $w=2.5e-07 $l=1.5e-06 $layer=POLY_cond $X=3.725 $Y=1.095
+ $X2=3.725 $Y2=2.595
r50 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.465 $Y=0.765
+ $X2=3.465 $Y2=0.93
r51 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.465 $Y=0.765
+ $X2=3.465 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%VPWR 1 2 3 12 18 22 25 26 28 29 30 36 45
+ 46 49
r65 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.05 $Y2=3.33
r69 40 42 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.05 $Y2=3.33
r72 36 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 34 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 30 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r76 30 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 30 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 28 42 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=3.42 $Y2=3.33
r80 27 45 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=4.08 $Y2=3.33
r81 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=3.42 $Y2=3.33
r82 25 33 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.99 $Y2=3.33
r84 24 38 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.99 $Y2=3.33
r86 20 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=3.245
+ $X2=3.42 $Y2=3.33
r87 20 22 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.42 $Y=3.245
+ $X2=3.42 $Y2=2.495
r88 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=3.33
r89 16 18 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=2.905
r90 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.99 $Y=2.24 $X2=0.99
+ $Y2=2.95
r91 10 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=3.245
+ $X2=0.99 $Y2=3.33
r92 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.99 $Y=3.245
+ $X2=0.99 $Y2=2.95
r93 3 22 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=2.095 $X2=3.42 $Y2=2.495
r94 2 18 600 $w=1.7e-07 $l=8.77211e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=2.095 $X2=2.05 $Y2=2.905
r95 1 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.85
+ $Y=2.095 $X2=0.99 $Y2=2.95
r96 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.85
+ $Y=2.095 $X2=0.99 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%Y 1 2 3 13 14 16 17 18 23 25 30 31
c66 25 0 1.19638e-19 $X=1.63 $Y=0.47
r67 31 34 0.664496 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.16 $Y=2.425
+ $X2=2.16 $Y2=2.33
r68 31 34 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=2.16 $Y=2.325
+ $X2=2.16 $Y2=2.33
r69 28 31 10.7728 $w=2.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.16 $Y=2.11
+ $X2=2.16 $Y2=2.325
r70 25 27 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.63 $Y=0.47
+ $X2=1.63 $Y2=0.675
r71 19 31 6.03773 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.275 $Y=2.425
+ $X2=2.16 $Y2=2.425
r72 18 30 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=2.425
+ $X2=2.89 $Y2=2.425
r73 18 19 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=2.725 $Y=2.425
+ $X2=2.275 $Y2=2.425
r74 16 28 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.045 $Y=2.025
+ $X2=2.16 $Y2=2.11
r75 16 17 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.045 $Y=2.025
+ $X2=1.77 $Y2=2.025
r76 15 23 4.61244 $w=1.9e-07 $l=1.74714e-07 $layer=LI1_cond $X=1.685 $Y=2.425
+ $X2=1.52 $Y2=2.405
r77 14 31 6.03773 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=2.425
+ $X2=2.16 $Y2=2.425
r78 14 15 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=2.045 $Y=2.425
+ $X2=1.685 $Y2=2.425
r79 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.685 $Y=1.94
+ $X2=1.77 $Y2=2.025
r80 13 27 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=1.685 $Y=1.94
+ $X2=1.685 $Y2=0.675
r81 3 30 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=2.75
+ $Y=2.095 $X2=2.89 $Y2=2.495
r82 2 23 300 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_PDIFF $count=2 $X=1.38
+ $Y=2.095 $X2=1.52 $Y2=2.455
r83 1 25 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.63 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r58 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r59 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r60 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r61 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r62 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.2
+ $Y2=0
r63 27 29 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=4.08
+ $Y2=0
r64 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r65 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r67 23 25 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=2.64 $Y2=0
r68 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=3.2
+ $Y2=0
r69 22 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=2.64
+ $Y2=0
r70 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r71 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r72 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r73 17 19 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r74 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r75 15 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r76 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.085 $X2=3.2
+ $Y2=0
r77 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.2 $Y=0.085
+ $X2=3.2 $Y2=0.4
r78 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r79 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0.445
r80 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.235 $X2=3.2 $Y2=0.4
r81 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.445
.ends

