* File: sky130_fd_sc_lp__a211oi_m.pxi.spice
* Created: Wed Sep  2 09:18:28 2020
* 
x_PM_SKY130_FD_SC_LP__A211OI_M%A2 N_A2_M1005_g N_A2_M1004_g N_A2_c_48_n
+ N_A2_c_49_n N_A2_c_50_n A2 A2 N_A2_c_51_n PM_SKY130_FD_SC_LP__A211OI_M%A2
x_PM_SKY130_FD_SC_LP__A211OI_M%A1 N_A1_M1001_g N_A1_M1006_g N_A1_c_77_n
+ N_A1_c_78_n A1 N_A1_c_79_n N_A1_c_80_n PM_SKY130_FD_SC_LP__A211OI_M%A1
x_PM_SKY130_FD_SC_LP__A211OI_M%B1 N_B1_M1003_g N_B1_M1002_g N_B1_c_114_n
+ N_B1_c_115_n B1 N_B1_c_117_n PM_SKY130_FD_SC_LP__A211OI_M%B1
x_PM_SKY130_FD_SC_LP__A211OI_M%C1 N_C1_M1007_g N_C1_M1000_g N_C1_c_150_n C1 C1
+ C1 PM_SKY130_FD_SC_LP__A211OI_M%C1
x_PM_SKY130_FD_SC_LP__A211OI_M%A_27_369# N_A_27_369#_M1004_s N_A_27_369#_M1006_d
+ N_A_27_369#_c_177_n N_A_27_369#_c_178_n N_A_27_369#_c_190_n
+ PM_SKY130_FD_SC_LP__A211OI_M%A_27_369#
x_PM_SKY130_FD_SC_LP__A211OI_M%VPWR N_VPWR_M1004_d N_VPWR_c_197_n VPWR
+ N_VPWR_c_198_n N_VPWR_c_199_n N_VPWR_c_196_n N_VPWR_c_201_n
+ PM_SKY130_FD_SC_LP__A211OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A211OI_M%Y N_Y_M1001_d N_Y_M1007_d N_Y_M1000_d N_Y_c_220_n
+ N_Y_c_214_n N_Y_c_215_n N_Y_c_216_n N_Y_c_217_n Y Y Y Y
+ PM_SKY130_FD_SC_LP__A211OI_M%Y
x_PM_SKY130_FD_SC_LP__A211OI_M%VGND N_VGND_M1005_s N_VGND_M1003_d N_VGND_c_252_n
+ N_VGND_c_253_n N_VGND_c_254_n VGND N_VGND_c_255_n N_VGND_c_256_n
+ N_VGND_c_257_n N_VGND_c_258_n PM_SKY130_FD_SC_LP__A211OI_M%VGND
cc_1 VNB N_A2_M1004_g 0.0178397f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.055
cc_2 VNB N_A2_c_48_n 0.0207565f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.765
cc_3 VNB N_A2_c_49_n 0.0268221f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.915
cc_4 VNB N_A2_c_50_n 0.0274561f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.435
cc_5 VNB N_A2_c_51_n 0.0391509f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.93
cc_6 VNB N_A1_M1001_g 0.0251381f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_7 VNB N_A1_M1006_g 0.004142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A1_c_77_n 0.0195623f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.285
cc_9 VNB N_A1_c_78_n 0.0147491f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.285
cc_10 VNB N_A1_c_79_n 0.0197317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_80_n 0.0131186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_M1003_g 0.0256982f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_13 VNB N_B1_M1002_g 0.00383951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_114_n 0.0187158f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.285
cc_15 VNB N_B1_c_115_n 0.019069f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.285
cc_16 VNB B1 0.0131054f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.435
cc_17 VNB N_B1_c_117_n 0.014738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C1_M1007_g 0.075604f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_19 VNB N_VPWR_c_196_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.925
cc_20 VNB N_Y_c_214_n 0.00625652f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_21 VNB N_Y_c_215_n 0.00915587f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_Y_c_216_n 0.0116356f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.93
cc_23 VNB N_Y_c_217_n 0.0076782f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.925
cc_24 VNB Y 0.0351163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_252_n 0.0103338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_253_n 0.0135112f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.765
cc_27 VNB N_VGND_c_254_n 0.00295613f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.435
cc_28 VNB N_VGND_c_255_n 0.0278679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_256_n 0.01882f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_30 VNB N_VGND_c_257_n 0.148363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_258_n 0.00521963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_A2_M1004_g 0.0309303f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.055
cc_33 VPB N_A1_M1006_g 0.0255315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_B1_M1002_g 0.0202709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_C1_M1007_g 0.0404006f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_36 VPB N_C1_c_150_n 0.0826154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB C1 0.0316098f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=0.765
cc_38 VPB C1 0.00473343f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=0.915
cc_39 VPB N_A_27_369#_c_177_n 0.0156387f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.285
cc_40 VPB N_A_27_369#_c_178_n 0.00851175f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.285
cc_41 VPB N_VPWR_c_197_n 0.0573696f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.055
cc_42 VPB N_VPWR_c_198_n 0.0194863f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=0.915
cc_43 VPB N_VPWR_c_199_n 0.0439346f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=0.93
cc_44 VPB N_VPWR_c_196_n 0.0915004f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=0.925
cc_45 VPB N_VPWR_c_201_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.295
cc_46 VPB Y 0.0201863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 N_A2_c_48_n N_A1_M1001_g 0.0517074f $X=0.337 $Y=0.765 $X2=0 $Y2=0
cc_48 A2 N_A1_M1001_g 9.37765e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_49 N_A2_M1004_g N_A1_M1006_g 0.0181708f $X=0.475 $Y=2.055 $X2=0 $Y2=0
cc_50 N_A2_c_50_n N_A1_c_77_n 0.00955724f $X=0.337 $Y=1.435 $X2=0 $Y2=0
cc_51 N_A2_M1004_g N_A1_c_78_n 0.00955724f $X=0.475 $Y=2.055 $X2=0 $Y2=0
cc_52 A2 N_A1_c_79_n 3.7954e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_53 N_A2_c_51_n N_A1_c_79_n 0.0147495f $X=0.29 $Y=0.93 $X2=0 $Y2=0
cc_54 N_A2_c_50_n N_A1_c_80_n 0.00408086f $X=0.337 $Y=1.435 $X2=0 $Y2=0
cc_55 A2 N_A1_c_80_n 0.0299746f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_56 N_A2_c_51_n N_A1_c_80_n 0.00204066f $X=0.29 $Y=0.93 $X2=0 $Y2=0
cc_57 N_A2_M1004_g N_A_27_369#_c_177_n 0.0189388f $X=0.475 $Y=2.055 $X2=0 $Y2=0
cc_58 N_A2_c_50_n N_A_27_369#_c_177_n 8.71842e-19 $X=0.337 $Y=1.435 $X2=0 $Y2=0
cc_59 A2 N_A_27_369#_c_177_n 0.00426754f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_60 N_A2_c_50_n N_A_27_369#_c_178_n 0.00543181f $X=0.337 $Y=1.435 $X2=0 $Y2=0
cc_61 A2 N_A_27_369#_c_178_n 0.0115333f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_62 N_A2_M1004_g N_VPWR_c_197_n 0.0128552f $X=0.475 $Y=2.055 $X2=0 $Y2=0
cc_63 N_A2_c_48_n N_VGND_c_253_n 0.010878f $X=0.337 $Y=0.765 $X2=0 $Y2=0
cc_64 N_A2_c_49_n N_VGND_c_253_n 0.0068247f $X=0.337 $Y=0.915 $X2=0 $Y2=0
cc_65 A2 N_VGND_c_253_n 0.0111987f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_A2_c_48_n N_VGND_c_255_n 0.00486043f $X=0.337 $Y=0.765 $X2=0 $Y2=0
cc_67 N_A2_c_48_n N_VGND_c_257_n 0.00729715f $X=0.337 $Y=0.765 $X2=0 $Y2=0
cc_68 A2 N_VGND_c_257_n 0.00229955f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_69 N_A1_M1001_g N_B1_M1003_g 0.0187209f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A1_M1006_g N_B1_M1002_g 0.0184997f $X=1.015 $Y=2.055 $X2=0 $Y2=0
cc_71 N_A1_c_77_n N_B1_c_114_n 0.0149567f $X=0.925 $Y=1.42 $X2=0 $Y2=0
cc_72 N_A1_c_78_n N_B1_c_115_n 0.0149567f $X=0.925 $Y=1.585 $X2=0 $Y2=0
cc_73 N_A1_c_79_n B1 6.37378e-19 $X=0.925 $Y=1.08 $X2=0 $Y2=0
cc_74 N_A1_c_80_n B1 0.0340191f $X=0.925 $Y=1.08 $X2=0 $Y2=0
cc_75 N_A1_c_79_n N_B1_c_117_n 0.0149567f $X=0.925 $Y=1.08 $X2=0 $Y2=0
cc_76 N_A1_c_80_n N_B1_c_117_n 6.37551e-19 $X=0.925 $Y=1.08 $X2=0 $Y2=0
cc_77 N_A1_M1006_g N_A_27_369#_c_177_n 0.0149512f $X=1.015 $Y=2.055 $X2=0 $Y2=0
cc_78 N_A1_c_78_n N_A_27_369#_c_177_n 0.00516074f $X=0.925 $Y=1.585 $X2=0 $Y2=0
cc_79 N_A1_c_80_n N_A_27_369#_c_177_n 0.0338618f $X=0.925 $Y=1.08 $X2=0 $Y2=0
cc_80 N_A1_M1006_g N_VPWR_c_197_n 0.00831167f $X=1.015 $Y=2.055 $X2=0 $Y2=0
cc_81 N_A1_M1001_g N_Y_c_220_n 0.00542452f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A1_M1001_g N_Y_c_215_n 0.00502338f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A1_c_79_n N_Y_c_215_n 0.00103161f $X=0.925 $Y=1.08 $X2=0 $Y2=0
cc_84 N_A1_c_80_n N_Y_c_215_n 0.00283146f $X=0.925 $Y=1.08 $X2=0 $Y2=0
cc_85 N_A1_M1001_g N_VGND_c_253_n 0.00209922f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A1_M1001_g N_VGND_c_254_n 0.00136958f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A1_M1001_g N_VGND_c_255_n 0.00585385f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A1_M1001_g N_VGND_c_257_n 0.011101f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_89 N_B1_M1003_g N_C1_M1007_g 0.0185814f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_90 N_B1_M1002_g N_C1_M1007_g 0.037419f $X=1.495 $Y=2.055 $X2=0 $Y2=0
cc_91 B1 N_C1_M1007_g 0.00356249f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_92 N_B1_c_117_n N_C1_M1007_g 0.0401688f $X=1.465 $Y=1.08 $X2=0 $Y2=0
cc_93 N_B1_M1002_g N_C1_c_150_n 0.010741f $X=1.495 $Y=2.055 $X2=0 $Y2=0
cc_94 N_B1_M1002_g C1 4.62255e-19 $X=1.495 $Y=2.055 $X2=0 $Y2=0
cc_95 N_B1_M1002_g C1 0.00115303f $X=1.495 $Y=2.055 $X2=0 $Y2=0
cc_96 N_B1_M1002_g N_A_27_369#_c_177_n 0.00261962f $X=1.495 $Y=2.055 $X2=0 $Y2=0
cc_97 N_B1_c_115_n N_A_27_369#_c_177_n 0.00103048f $X=1.465 $Y=1.585 $X2=0 $Y2=0
cc_98 B1 N_A_27_369#_c_177_n 0.00282208f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B1_M1003_g N_Y_c_214_n 0.0121491f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_100 B1 N_Y_c_214_n 0.0346505f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B1_c_117_n N_Y_c_214_n 0.00514801f $X=1.465 $Y=1.08 $X2=0 $Y2=0
cc_102 N_B1_M1003_g Y 4.58782e-19 $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_103 N_B1_M1002_g Y 0.00181585f $X=1.495 $Y=2.055 $X2=0 $Y2=0
cc_104 N_B1_c_115_n Y 4.36259e-19 $X=1.465 $Y=1.585 $X2=0 $Y2=0
cc_105 B1 Y 0.0367409f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B1_c_117_n Y 8.49423e-19 $X=1.465 $Y=1.08 $X2=0 $Y2=0
cc_107 N_B1_M1003_g N_VGND_c_254_n 0.00742704f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B1_M1003_g N_VGND_c_255_n 0.00411627f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_109 N_B1_M1003_g N_VGND_c_257_n 0.00507831f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_110 N_C1_c_150_n N_A_27_369#_c_190_n 2.63493e-19 $X=1.84 $Y=2.775 $X2=0 $Y2=0
cc_111 C1 N_A_27_369#_c_190_n 5.09399e-19 $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_112 N_C1_c_150_n N_VPWR_c_197_n 0.00206959f $X=1.84 $Y=2.775 $X2=0 $Y2=0
cc_113 C1 N_VPWR_c_197_n 0.0135142f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_114 N_C1_c_150_n N_VPWR_c_199_n 0.011282f $X=1.84 $Y=2.775 $X2=0 $Y2=0
cc_115 C1 N_VPWR_c_199_n 0.0148879f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_116 C1 N_VPWR_c_199_n 0.0182867f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_117 N_C1_c_150_n N_VPWR_c_196_n 0.015816f $X=1.84 $Y=2.775 $X2=0 $Y2=0
cc_118 C1 N_VPWR_c_196_n 0.014039f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_119 C1 N_VPWR_c_196_n 0.0182294f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_120 N_C1_M1007_g N_Y_c_214_n 0.0128434f $X=1.915 $Y=0.445 $X2=0 $Y2=0
cc_121 N_C1_M1007_g N_Y_c_217_n 0.00416651f $X=1.915 $Y=0.445 $X2=0 $Y2=0
cc_122 N_C1_M1007_g Y 0.0414252f $X=1.915 $Y=0.445 $X2=0 $Y2=0
cc_123 C1 Y 0.0200637f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_124 N_C1_M1007_g N_VGND_c_254_n 0.00716165f $X=1.915 $Y=0.445 $X2=0 $Y2=0
cc_125 N_C1_M1007_g N_VGND_c_256_n 0.0042654f $X=1.915 $Y=0.445 $X2=0 $Y2=0
cc_126 N_C1_M1007_g N_VGND_c_257_n 0.00725794f $X=1.915 $Y=0.445 $X2=0 $Y2=0
cc_127 N_A_27_369#_c_177_n N_VPWR_M1004_d 0.00326552f $X=1.125 $Y=1.77 $X2=-0.19
+ $Y2=1.655
cc_128 N_A_27_369#_c_177_n N_VPWR_c_197_n 0.0210643f $X=1.125 $Y=1.77 $X2=0
+ $Y2=0
cc_129 N_A_27_369#_c_177_n Y 0.00525052f $X=1.125 $Y=1.77 $X2=0 $Y2=0
cc_130 N_A_27_369#_c_190_n Y 0.00701414f $X=1.23 $Y=1.97 $X2=0 $Y2=0
cc_131 N_Y_c_214_n N_VGND_M1003_d 0.00295242f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_132 N_Y_c_220_n N_VGND_c_253_n 0.00371471f $X=1.16 $Y=0.51 $X2=0 $Y2=0
cc_133 N_Y_c_214_n N_VGND_c_254_n 0.0196407f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_134 N_Y_c_220_n N_VGND_c_255_n 0.00857019f $X=1.16 $Y=0.51 $X2=0 $Y2=0
cc_135 N_Y_c_214_n N_VGND_c_255_n 0.00263146f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_136 N_Y_c_214_n N_VGND_c_256_n 0.00265869f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_137 N_Y_c_216_n N_VGND_c_256_n 0.0114859f $X=2.13 $Y=0.51 $X2=0 $Y2=0
cc_138 N_Y_c_217_n N_VGND_c_256_n 7.64527e-19 $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_139 N_Y_M1001_d N_VGND_c_257_n 0.00841067f $X=0.91 $Y=0.235 $X2=0 $Y2=0
cc_140 N_Y_M1007_d N_VGND_c_257_n 0.0023508f $X=1.99 $Y=0.235 $X2=0 $Y2=0
cc_141 N_Y_c_220_n N_VGND_c_257_n 0.00761208f $X=1.16 $Y=0.51 $X2=0 $Y2=0
cc_142 N_Y_c_214_n N_VGND_c_257_n 0.0106691f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_143 N_Y_c_216_n N_VGND_c_257_n 0.00992777f $X=2.13 $Y=0.51 $X2=0 $Y2=0
cc_144 N_Y_c_217_n N_VGND_c_257_n 0.00166523f $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_145 N_VGND_c_257_n A_110_47# 0.00899413f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
