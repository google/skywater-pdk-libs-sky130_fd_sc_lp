* File: sky130_fd_sc_lp__buf_0.pex.spice
* Created: Fri Aug 28 10:09:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUF_0%A_70_157# 1 2 9 12 15 16 17 18 19 21 22 24 25
+ 28 32 36 37
r63 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.515
+ $Y=0.95 $X2=0.515 $Y2=0.95
r64 30 32 12.9397 $w=2.83e-07 $l=3.2e-07 $layer=LI1_cond $X=1.202 $Y=0.785
+ $X2=1.202 $Y2=0.465
r65 26 28 20.4147 $w=3.48e-07 $l=6.2e-07 $layer=LI1_cond $X=1.17 $Y=2.225
+ $X2=1.17 $Y2=2.845
r66 24 26 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.995 $Y=2.14
+ $X2=1.17 $Y2=2.225
r67 24 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.995 $Y=2.14
+ $X2=0.68 $Y2=2.14
r68 23 35 4.02313 $w=1.85e-07 $l=1.25e-07 $layer=LI1_cond $X=0.68 $Y=0.877
+ $X2=0.555 $Y2=0.877
r69 22 30 7.22568 $w=1.85e-07 $l=1.82285e-07 $layer=LI1_cond $X=1.06 $Y=0.877
+ $X2=1.202 $Y2=0.785
r70 22 23 22.7813 $w=1.83e-07 $l=3.8e-07 $layer=LI1_cond $X=1.06 $Y=0.877
+ $X2=0.68 $Y2=0.877
r71 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.595 $Y=2.055
+ $X2=0.68 $Y2=2.14
r72 21 37 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.595 $Y=2.055
+ $X2=0.595 $Y2=1.455
r73 19 37 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=1.33
+ $X2=0.555 $Y2=1.455
r74 18 35 2.99321 $w=2.5e-07 $l=9.3e-08 $layer=LI1_cond $X=0.555 $Y=0.97
+ $X2=0.555 $Y2=0.877
r75 18 19 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=0.555 $Y=0.97
+ $X2=0.555 $Y2=1.33
r76 16 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.515 $Y=1.29
+ $X2=0.515 $Y2=0.95
r77 16 17 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.29
+ $X2=0.515 $Y2=1.455
r78 15 36 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=0.785
+ $X2=0.515 $Y2=0.95
r79 12 17 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=0.475 $Y=2.735
+ $X2=0.475 $Y2=1.455
r80 9 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.465
+ $X2=0.475 $Y2=0.785
r81 2 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=2.635 $X2=1.18 $Y2=2.845
r82 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.255 $X2=1.18 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_0%A 3 7 11 12 13 14 18
r33 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.055
+ $Y=1.38 $X2=1.055 $Y2=1.38
r34 14 19 7.49192 $w=4.53e-07 $l=2.85e-07 $layer=LI1_cond $X=1.117 $Y=1.665
+ $X2=1.117 $Y2=1.38
r35 13 19 2.23443 $w=4.53e-07 $l=8.5e-08 $layer=LI1_cond $X=1.117 $Y=1.295
+ $X2=1.117 $Y2=1.38
r36 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.055 $Y=1.72
+ $X2=1.055 $Y2=1.38
r37 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.72
+ $X2=1.055 $Y2=1.885
r38 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.215
+ $X2=1.055 $Y2=1.38
r39 7 12 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=0.965 $Y=2.845
+ $X2=0.965 $Y2=1.885
r40 3 10 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.965 $Y=0.465
+ $X2=0.965 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_0%X 1 2 12 14 15 16 17 18 29 34
r23 34 35 0.83707 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=0.245 $Y=2.405
+ $X2=0.245 $Y2=2.395
r24 27 29 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=0.245 $Y=2.55
+ $X2=0.245 $Y2=2.56
r25 18 29 7.99275 $w=3.08e-07 $l=2.15e-07 $layer=LI1_cond $X=0.245 $Y=2.775
+ $X2=0.245 $Y2=2.56
r26 17 27 4.01496 $w=3.08e-07 $l=1.08e-07 $layer=LI1_cond $X=0.245 $Y=2.442
+ $X2=0.245 $Y2=2.55
r27 17 34 1.3755 $w=3.08e-07 $l=3.7e-08 $layer=LI1_cond $X=0.245 $Y=2.442
+ $X2=0.245 $Y2=2.405
r28 17 35 1.75171 $w=2.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.215 $Y=2.357
+ $X2=0.215 $Y2=2.395
r29 16 17 14.8435 $w=2.48e-07 $l=3.22e-07 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=2.357
r30 14 16 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.215 $Y=1.73
+ $X2=0.215 $Y2=2.035
r31 14 15 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=1.73
+ $X2=0.215 $Y2=1.605
r32 9 12 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=0.45
+ $X2=0.26 $Y2=0.45
r33 7 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.175 $Y=0.615
+ $X2=0.175 $Y2=0.45
r34 7 15 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=0.175 $Y=0.615
+ $X2=0.175 $Y2=1.605
r35 2 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.415 $X2=0.26 $Y2=2.56
r36 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.255 $X2=0.26 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_0%VPWR 1 6 10 12 19 20 23
r20 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r21 17 23 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.697 $Y2=3.33
r22 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=1.2 $Y2=3.33
r23 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 12 23 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.697 $Y2=3.33
r25 12 14 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r26 10 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r27 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 10 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 6 9 15.8178 $w=2.53e-07 $l=3.5e-07 $layer=LI1_cond $X=0.697 $Y=2.56
+ $X2=0.697 $Y2=2.91
r30 4 23 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.697 $Y=3.245
+ $X2=0.697 $Y2=3.33
r31 4 9 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=0.697 $Y=3.245
+ $X2=0.697 $Y2=2.91
r32 1 9 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.415 $X2=0.69 $Y2=2.91
r33 1 6 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.415 $X2=0.69 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_0%VGND 1 6 8 10 17 18 21
r21 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r22 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.725
+ $Y2=0
r23 15 17 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r24 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r25 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.725
+ $Y2=0
r26 10 12 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r27 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r28 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r29 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r31 4 6 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.465
r32 1 6 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.255 $X2=0.725 $Y2=0.465
.ends

