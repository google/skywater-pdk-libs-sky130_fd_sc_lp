* File: sky130_fd_sc_lp__o32ai_2.pex.spice
* Created: Fri Aug 28 11:18:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32AI_2%B2 3 7 11 15 17 18 19 28
r44 26 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.625 $Y=1.51
+ $X2=0.965 $Y2=1.51
r45 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.51 $X2=0.625 $Y2=1.51
r46 23 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.535 $Y=1.51
+ $X2=0.625 $Y2=1.51
r47 18 19 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=1.2 $Y2=1.587
r48 18 27 3.36868 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=0.625 $Y2=1.587
r49 17 27 13.652 $w=3.23e-07 $l=3.85e-07 $layer=LI1_cond $X=0.24 $Y=1.587
+ $X2=0.625 $Y2=1.587
r50 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.675
+ $X2=0.965 $Y2=1.51
r51 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.965 $Y=1.675
+ $X2=0.965 $Y2=2.465
r52 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.345
+ $X2=0.965 $Y2=1.51
r53 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.965 $Y=1.345 $X2=0.965
+ $Y2=0.745
r54 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.675
+ $X2=0.535 $Y2=1.51
r55 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.535 $Y=1.675
+ $X2=0.535 $Y2=2.465
r56 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.345
+ $X2=0.535 $Y2=1.51
r57 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.535 $Y=1.345 $X2=0.535
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%B1 3 7 11 15 17 23 24
c49 23 0 1.26527e-19 $X=1.63 $Y=1.51
c50 3 0 2.33755e-21 $X=1.395 $Y=2.465
r51 24 25 23.2289 $w=3.32e-07 $l=1.6e-07 $layer=POLY_cond $X=1.825 $Y=1.512
+ $X2=1.985 $Y2=1.512
r52 22 24 28.3102 $w=3.32e-07 $l=1.95e-07 $layer=POLY_cond $X=1.63 $Y=1.512
+ $X2=1.825 $Y2=1.512
r53 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.51 $X2=1.63 $Y2=1.51
r54 20 22 22.503 $w=3.32e-07 $l=1.55e-07 $layer=POLY_cond $X=1.475 $Y=1.512
+ $X2=1.63 $Y2=1.512
r55 17 23 4.89394 $w=3.63e-07 $l=1.55e-07 $layer=LI1_cond $X=1.647 $Y=1.665
+ $X2=1.647 $Y2=1.51
r56 13 25 21.3668 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=1.985 $Y=1.345
+ $X2=1.985 $Y2=1.512
r57 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.985 $Y=1.345
+ $X2=1.985 $Y2=0.745
r58 9 24 21.3668 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=1.825 $Y=1.68
+ $X2=1.825 $Y2=1.512
r59 9 11 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.825 $Y=1.68
+ $X2=1.825 $Y2=2.465
r60 5 20 21.3668 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=1.475 $Y=1.345
+ $X2=1.475 $Y2=1.512
r61 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.475 $Y=1.345 $X2=1.475
+ $Y2=0.745
r62 1 20 11.6145 $w=3.32e-07 $l=8e-08 $layer=POLY_cond $X=1.395 $Y=1.512
+ $X2=1.475 $Y2=1.512
r63 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.395 $Y=1.675
+ $X2=1.395 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%A3 3 7 11 15 17 18 28
c59 28 0 1.26527e-19 $X=3.455 $Y=1.5
c60 18 0 2.33755e-21 $X=2.64 $Y=1.665
r61 27 28 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.385 $Y=1.5 $X2=3.455
+ $Y2=1.5
r62 26 27 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.955 $Y=1.5
+ $X2=3.385 $Y2=1.5
r63 24 26 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.585 $Y=1.5
+ $X2=2.955 $Y2=1.5
r64 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=1.5 $X2=2.585 $Y2=1.5
r65 21 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.495 $Y=1.5 $X2=2.585
+ $Y2=1.5
r66 18 25 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=2.64 $Y=1.582
+ $X2=2.585 $Y2=1.582
r67 17 25 14.6205 $w=3.33e-07 $l=4.25e-07 $layer=LI1_cond $X=2.16 $Y=1.582
+ $X2=2.585 $Y2=1.582
r68 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.455 $Y=1.335
+ $X2=3.455 $Y2=1.5
r69 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.455 $Y=1.335
+ $X2=3.455 $Y2=0.745
r70 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.385 $Y=1.665
+ $X2=3.385 $Y2=1.5
r71 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.385 $Y=1.665
+ $X2=3.385 $Y2=2.455
r72 5 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.665
+ $X2=2.955 $Y2=1.5
r73 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.955 $Y=1.665
+ $X2=2.955 $Y2=2.455
r74 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.335
+ $X2=2.495 $Y2=1.5
r75 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.495 $Y=1.335
+ $X2=2.495 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%A2 3 5 7 10 12 14 15 16 17 28
c55 28 0 5.67181e-19 $X=4.355 $Y=1.44
c56 12 0 4.85921e-20 $X=4.355 $Y=1.275
r57 26 28 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.335 $Y=1.44
+ $X2=4.355 $Y2=1.44
r58 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.335
+ $Y=1.44 $X2=4.335 $Y2=1.44
r59 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.245 $Y=1.44
+ $X2=4.335 $Y2=1.44
r60 23 24 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.895 $Y=1.44
+ $X2=4.245 $Y2=1.44
r61 21 23 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.815 $Y=1.44
+ $X2=3.895 $Y2=1.44
r62 17 27 8.23174 $w=3.13e-07 $l=2.25e-07 $layer=LI1_cond $X=4.56 $Y=1.367
+ $X2=4.335 $Y2=1.367
r63 16 27 9.3293 $w=3.13e-07 $l=2.55e-07 $layer=LI1_cond $X=4.08 $Y=1.367
+ $X2=4.335 $Y2=1.367
r64 15 16 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.367 $X2=4.08
+ $Y2=1.367
r65 12 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.275
+ $X2=4.355 $Y2=1.44
r66 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.355 $Y=1.275
+ $X2=4.355 $Y2=0.745
r67 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.605
+ $X2=4.245 $Y2=1.44
r68 8 10 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=4.245 $Y=1.605
+ $X2=4.245 $Y2=2.455
r69 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.895 $Y=1.275
+ $X2=3.895 $Y2=1.44
r70 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.895 $Y=1.275
+ $X2=3.895 $Y2=0.745
r71 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.605
+ $X2=3.815 $Y2=1.44
r72 1 3 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=3.815 $Y=1.605
+ $X2=3.815 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%A1 1 3 6 8 10 13 15 16 17 31
c39 17 0 2.4547e-19 $X=6 $Y=1.295
r40 29 31 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.535 $Y=1.44
+ $X2=5.625 $Y2=1.44
r41 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.535
+ $Y=1.44 $X2=5.535 $Y2=1.44
r42 27 29 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=5.215 $Y=1.44
+ $X2=5.535 $Y2=1.44
r43 26 27 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.195 $Y=1.44
+ $X2=5.215 $Y2=1.44
r44 24 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.98 $Y=1.44
+ $X2=5.195 $Y2=1.44
r45 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.98
+ $Y=1.44 $X2=4.98 $Y2=1.44
r46 21 24 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.785 $Y=1.44
+ $X2=4.98 $Y2=1.44
r47 17 30 17.0123 $w=3.13e-07 $l=4.65e-07 $layer=LI1_cond $X=6 $Y=1.367
+ $X2=5.535 $Y2=1.367
r48 16 30 0.548782 $w=3.13e-07 $l=1.5e-08 $layer=LI1_cond $X=5.52 $Y=1.367
+ $X2=5.535 $Y2=1.367
r49 15 16 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.367
+ $X2=5.52 $Y2=1.367
r50 15 25 2.19513 $w=3.13e-07 $l=6e-08 $layer=LI1_cond $X=5.04 $Y=1.367 $X2=4.98
+ $Y2=1.367
r51 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.625 $Y=1.605
+ $X2=5.625 $Y2=1.44
r52 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.625 $Y=1.605
+ $X2=5.625 $Y2=2.465
r53 8 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.215 $Y=1.275
+ $X2=5.215 $Y2=1.44
r54 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.215 $Y=1.275
+ $X2=5.215 $Y2=0.745
r55 4 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.195 $Y=1.605
+ $X2=5.195 $Y2=1.44
r56 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.195 $Y=1.605
+ $X2=5.195 $Y2=2.465
r57 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.275
+ $X2=4.785 $Y2=1.44
r58 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.785 $Y=1.275
+ $X2=4.785 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%A_39_367# 1 2 3 10 12 14 16 18 20 22
r30 20 29 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=2.075 $Y=2.45
+ $X2=2.075 $Y2=2.355
r31 20 22 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=2.075 $Y=2.45
+ $X2=2.075 $Y2=2.91
r32 19 27 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.275 $Y=2.355
+ $X2=1.18 $Y2=2.355
r33 18 29 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=1.945 $Y=2.355
+ $X2=2.075 $Y2=2.355
r34 18 19 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.945 $Y=2.355
+ $X2=1.275 $Y2=2.355
r35 16 27 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.18 $Y=2.45 $X2=1.18
+ $Y2=2.355
r36 16 17 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=1.18 $Y=2.45
+ $X2=1.18 $Y2=2.905
r37 15 25 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.415 $Y=2.99
+ $X2=0.285 $Y2=2.99
r38 14 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.18 $Y2=2.905
r39 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.415 $Y2=2.99
r40 10 25 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.905
+ $X2=0.285 $Y2=2.99
r41 10 12 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.285 $Y=2.905
+ $X2=0.285 $Y2=2.085
r42 3 29 600 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.835 $X2=2.04 $Y2=2.345
r43 3 22 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.835 $X2=2.04 $Y2=2.91
r44 2 27 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=1.835 $X2=1.18 $Y2=2.425
r45 1 25 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.32 $Y2=2.91
r46 1 12 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.32 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%Y 1 2 3 4 15 19 20 21 25 27 30 31 32 33 34
+ 35 42 45
r86 42 45 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=1.245 $X2=3.17
+ $Y2=1.295
r87 35 54 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.17 $Y=2.405
+ $X2=3.17 $Y2=2.65
r88 34 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=2.005
+ $X2=3.17 $Y2=1.92
r89 34 49 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=2.005
+ $X2=3.17 $Y2=2.09
r90 34 35 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.17 $Y=2.105 $X2=3.17
+ $Y2=2.405
r91 34 49 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.17 $Y=2.105
+ $X2=3.17 $Y2=2.09
r92 33 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.17 $Y=1.665
+ $X2=3.17 $Y2=1.92
r93 32 42 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=1.16 $X2=3.17
+ $Y2=1.245
r94 32 33 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=3.17 $Y=1.312
+ $X2=3.17 $Y2=1.665
r95 32 45 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=3.17 $Y=1.312
+ $X2=3.17 $Y2=1.295
r96 28 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=1.16
+ $X2=1.77 $Y2=1.16
r97 27 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=1.16
+ $X2=3.17 $Y2=1.16
r98 27 28 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.005 $Y=1.16
+ $X2=1.935 $Y2=1.16
r99 23 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=1.075
+ $X2=1.77 $Y2=1.16
r100 23 25 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.77 $Y=1.075
+ $X2=1.77 $Y2=0.68
r101 22 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=2.005
+ $X2=0.75 $Y2=2.005
r102 21 34 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=2.005
+ $X2=3.17 $Y2=2.005
r103 21 22 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=3.005 $Y=2.005
+ $X2=0.915 $Y2=2.005
r104 19 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=1.16
+ $X2=1.77 $Y2=1.16
r105 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.605 $Y=1.16
+ $X2=0.915 $Y2=1.16
r106 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.75 $Y=1.075
+ $X2=0.915 $Y2=1.16
r107 13 15 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.75 $Y=1.075
+ $X2=0.75 $Y2=0.68
r108 4 34 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.825 $X2=3.17 $Y2=1.95
r109 4 54 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.825 $X2=3.17 $Y2=2.65
r110 3 30 300 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.835 $X2=0.75 $Y2=2.015
r111 2 25 91 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.325 $X2=1.77 $Y2=0.68
r112 1 15 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=0.61
+ $Y=0.325 $X2=0.75 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%VPWR 1 2 3 12 16 20 22 26 28 36 44 50 53 57
r75 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r76 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 48 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r79 48 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r80 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 45 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=3.33
+ $X2=4.98 $Y2=3.33
r82 45 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.145 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 44 56 4.23407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.975 $Y2=3.33
r84 44 47 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r88 39 42 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r89 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r90 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=3.33
+ $X2=1.61 $Y2=3.33
r91 37 39 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.775 $Y=3.33
+ $X2=2.16 $Y2=3.33
r92 36 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=3.33
+ $X2=4.98 $Y2=3.33
r93 36 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.815 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r96 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r97 30 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r98 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 28 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.61 $Y2=3.33
r100 28 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r101 26 43 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r102 26 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 22 25 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=5.857 $Y=1.98
+ $X2=5.857 $Y2=2.95
r104 20 56 3.24346 $w=2.95e-07 $l=1.54771e-07 $layer=LI1_cond $X=5.857 $Y=3.245
+ $X2=5.975 $Y2=3.33
r105 20 25 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=5.857 $Y=3.245
+ $X2=5.857 $Y2=2.95
r106 16 19 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.98 $Y=2.13
+ $X2=4.98 $Y2=2.95
r107 14 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=3.245
+ $X2=4.98 $Y2=3.33
r108 14 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.98 $Y=3.245
+ $X2=4.98 $Y2=2.95
r109 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=3.245
+ $X2=1.61 $Y2=3.33
r110 10 12 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.61 $Y=3.245
+ $X2=1.61 $Y2=2.745
r111 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.835 $X2=5.84 $Y2=2.95
r112 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.835 $X2=5.84 $Y2=1.98
r113 2 19 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.835 $X2=4.98 $Y2=2.95
r114 2 16 400 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.835 $X2=4.98 $Y2=2.13
r115 1 12 600 $w=1.7e-07 $l=9.77497e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.835 $X2=1.61 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%A_519_365# 1 2 3 12 14 15 18 20 22 24 27
r42 22 29 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.905
+ $X2=4.495 $Y2=2.99
r43 22 24 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=4.495 $Y=2.905
+ $X2=4.495 $Y2=2.21
r44 21 27 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.695 $Y=2.99 $X2=3.6
+ $Y2=2.99
r45 20 29 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.365 $Y=2.99
+ $X2=4.495 $Y2=2.99
r46 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.365 $Y=2.99
+ $X2=3.695 $Y2=2.99
r47 16 27 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.905 $X2=3.6
+ $Y2=2.99
r48 16 18 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=3.6 $Y=2.905
+ $X2=3.6 $Y2=1.98
r49 14 27 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.505 $Y=2.99 $X2=3.6
+ $Y2=2.99
r50 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.505 $Y=2.99
+ $X2=2.825 $Y2=2.99
r51 10 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.69 $Y=2.905
+ $X2=2.825 $Y2=2.99
r52 10 12 20.4879 $w=2.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.69 $Y=2.905
+ $X2=2.69 $Y2=2.425
r53 3 29 400 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.825 $X2=4.46 $Y2=2.91
r54 3 24 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.825 $X2=4.46 $Y2=2.21
r55 2 27 400 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=3.46
+ $Y=1.825 $X2=3.6 $Y2=2.91
r56 2 18 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=3.46
+ $Y=1.825 $X2=3.6 $Y2=1.98
r57 1 12 300 $w=1.7e-07 $l=6.59545e-07 $layer=licon1_PDIFF $count=2 $X=2.595
+ $Y=1.825 $X2=2.72 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%A_778_365# 1 2 9 13 14 17
r31 17 19 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=5.427 $Y=1.98
+ $X2=5.427 $Y2=2.91
r32 15 17 5.37807 $w=2.23e-07 $l=1.05e-07 $layer=LI1_cond $X=5.427 $Y=1.875
+ $X2=5.427 $Y2=1.98
r33 13 15 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=5.315 $Y=1.79
+ $X2=5.427 $Y2=1.875
r34 13 14 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=5.315 $Y=1.79
+ $X2=4.195 $Y2=1.79
r35 9 11 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.03 $Y=1.95 $X2=4.03
+ $Y2=2.65
r36 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.03 $Y=1.875
+ $X2=4.195 $Y2=1.79
r37 7 9 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=4.03 $Y=1.875 $X2=4.03
+ $Y2=1.95
r38 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.835 $X2=5.41 $Y2=2.91
r39 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.835 $X2=5.41 $Y2=1.98
r40 1 11 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.825 $X2=4.03 $Y2=2.65
r41 1 9 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.825 $X2=4.03 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%A_39_65# 1 2 3 4 5 6 21 23 24 27 29 34 35 36
+ 39 41 45 47 49 51 53 54 60
c89 60 0 1.75061e-19 $X=4.57 $Y=0.955
c90 54 0 1.95243e-19 $X=3.64 $Y=0.82
r91 54 57 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.64 $Y=0.82
+ $X2=3.64 $Y2=0.955
r92 54 55 4.4265 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.82 $X2=3.64
+ $Y2=0.735
r93 49 62 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=0.87
+ $X2=5.465 $Y2=0.955
r94 49 51 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=5.465 $Y=0.87
+ $X2=5.465 $Y2=0.48
r95 48 60 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.665 $Y=0.955
+ $X2=4.565 $Y2=0.955
r96 47 62 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.335 $Y=0.955
+ $X2=5.465 $Y2=0.955
r97 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.335 $Y=0.955
+ $X2=4.665 $Y2=0.955
r98 43 60 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0.87
+ $X2=4.565 $Y2=0.955
r99 43 45 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=4.565 $Y=0.87
+ $X2=4.565 $Y2=0.48
r100 42 57 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.775 $Y=0.955
+ $X2=3.64 $Y2=0.955
r101 41 60 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.465 $Y=0.955
+ $X2=4.565 $Y2=0.955
r102 41 42 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.465 $Y=0.955
+ $X2=3.775 $Y2=0.955
r103 39 55 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.675 $Y=0.48
+ $X2=3.675 $Y2=0.735
r104 35 54 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.505 $Y=0.82
+ $X2=3.64 $Y2=0.82
r105 35 36 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.505 $Y=0.82
+ $X2=2.445 $Y2=0.82
r106 32 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.28 $Y=0.735
+ $X2=2.445 $Y2=0.82
r107 32 34 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.28 $Y=0.735
+ $X2=2.28 $Y2=0.45
r108 31 34 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.28 $Y=0.425
+ $X2=2.28 $Y2=0.45
r109 30 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=0.34
+ $X2=1.26 $Y2=0.34
r110 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.115 $Y=0.34
+ $X2=2.28 $Y2=0.425
r111 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.115 $Y=0.34
+ $X2=1.425 $Y2=0.34
r112 25 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=0.425
+ $X2=1.26 $Y2=0.34
r113 25 27 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.26 $Y=0.425
+ $X2=1.26 $Y2=0.45
r114 23 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=0.34
+ $X2=1.26 $Y2=0.34
r115 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.095 $Y=0.34
+ $X2=0.415 $Y2=0.34
r116 19 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.285 $Y=0.425
+ $X2=0.415 $Y2=0.34
r117 19 21 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.285 $Y=0.425
+ $X2=0.285 $Y2=0.47
r118 6 62 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.325 $X2=5.43 $Y2=0.955
r119 6 51 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.325 $X2=5.43 $Y2=0.48
r120 5 60 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.325 $X2=4.57 $Y2=0.955
r121 5 45 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.325 $X2=4.57 $Y2=0.48
r122 4 57 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=3.53
+ $Y=0.325 $X2=3.67 $Y2=0.955
r123 4 39 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.53
+ $Y=0.325 $X2=3.67 $Y2=0.48
r124 3 34 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.325 $X2=2.28 $Y2=0.45
r125 2 27 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=1.04
+ $Y=0.325 $X2=1.26 $Y2=0.45
r126 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.195
+ $Y=0.325 $X2=0.32 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_2%VGND 1 2 3 12 16 18 25 30 37 38 43 49 51 54
r72 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r73 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r74 48 49 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0.24
+ $X2=3.405 $Y2=0.24
r75 45 48 2.20814 $w=6.48e-07 $l=1.2e-07 $layer=LI1_cond $X=3.12 $Y=0.24
+ $X2=3.24 $Y2=0.24
r76 41 45 8.83258 $w=6.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0.24
+ $X2=3.12 $Y2=0.24
r77 41 43 7.90576 $w=6.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.64 $Y=0.24
+ $X2=2.615 $Y2=0.24
r78 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r79 38 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r80 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r81 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r82 35 37 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=6
+ $Y2=0
r83 34 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r84 34 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r85 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r86 31 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=0 $X2=4.11
+ $Y2=0
r87 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=0 $X2=4.56
+ $Y2=0
r88 30 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r89 30 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.56
+ $Y2=0
r90 29 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r91 28 49 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.405
+ $Y2=0
r92 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r93 25 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=4.11
+ $Y2=0
r94 25 28 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=3.6
+ $Y2=0
r95 23 42 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r96 22 43 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=0.24 $Y=0
+ $X2=2.615 $Y2=0
r97 22 23 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r98 18 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r99 18 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r100 18 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r101 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r102 14 16 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.575
r103 10 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0
r104 10 12 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0.575
r105 3 16 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.325 $X2=5 $Y2=0.575
r106 2 12 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.97
+ $Y=0.325 $X2=4.11 $Y2=0.575
r107 1 48 91 $w=1.7e-07 $l=7.38952e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.325 $X2=3.24 $Y2=0.47
.ends

