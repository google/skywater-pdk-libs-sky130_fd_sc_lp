* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__clkbuflp_4 A VGND VNB VPB VPWR X
X0 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_110_47# A a_130_417# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 VPWR A a_130_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_372_47# a_130_417# X VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X6 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 X a_130_417# a_530_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X8 a_530_47# a_130_417# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X9 a_130_417# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND a_130_417# a_372_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X11 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
