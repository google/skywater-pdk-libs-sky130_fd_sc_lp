# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a32oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a32oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.425000 2.765000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.425000 4.655000 1.750000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.755000 1.195000 6.155000 1.525000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 1.425000 2.265000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.485000 1.275000 ;
        RECT 0.085000 1.275000 1.060000 1.525000 ;
        RECT 0.085000 1.525000 0.435000 1.760000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.695000 1.725000 1.865000 ;
        RECT 0.605000 1.865000 0.935000 2.735000 ;
        RECT 1.465000 0.605000 1.795000 1.075000 ;
        RECT 1.465000 1.075000 3.335000 1.245000 ;
        RECT 1.465000 1.865000 1.725000 1.920000 ;
        RECT 1.465000 1.920000 3.335000 2.120000 ;
        RECT 1.465000 2.120000 1.795000 2.735000 ;
        RECT 3.005000 0.605000 3.335000 1.075000 ;
        RECT 3.005000 1.245000 3.335000 1.920000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.240000 0.085000 ;
        RECT 0.605000  0.085000 0.935000 0.700000 ;
        RECT 4.895000  0.085000 5.225000 0.905000 ;
        RECT 5.755000  0.085000 6.085000 1.025000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.240000 3.415000 ;
        RECT 2.560000 2.630000 3.335000 3.245000 ;
        RECT 3.945000 2.260000 4.645000 3.245000 ;
        RECT 5.175000 2.095000 5.505000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.315000 0.435000 0.870000 ;
      RECT 0.175000 0.870000 1.295000 1.040000 ;
      RECT 0.175000 1.930000 0.435000 2.905000 ;
      RECT 0.175000 2.905000 2.345000 3.075000 ;
      RECT 1.105000 0.265000 2.295000 0.435000 ;
      RECT 1.105000 0.435000 1.295000 0.870000 ;
      RECT 1.105000 2.035000 1.295000 2.905000 ;
      RECT 1.965000 0.435000 2.295000 0.905000 ;
      RECT 2.015000 2.290000 3.775000 2.460000 ;
      RECT 2.015000 2.460000 2.345000 2.905000 ;
      RECT 2.505000 0.265000 4.695000 0.435000 ;
      RECT 2.505000 0.435000 2.835000 0.905000 ;
      RECT 3.505000 0.435000 3.695000 1.205000 ;
      RECT 3.505000 2.460000 3.775000 3.075000 ;
      RECT 3.515000 1.920000 5.935000 1.925000 ;
      RECT 3.515000 1.925000 5.005000 2.090000 ;
      RECT 3.515000 2.090000 3.775000 2.290000 ;
      RECT 3.865000 0.605000 4.195000 1.075000 ;
      RECT 3.865000 1.075000 5.585000 1.245000 ;
      RECT 4.365000 0.435000 4.695000 0.905000 ;
      RECT 4.815000 2.090000 5.005000 3.075000 ;
      RECT 4.825000 1.755000 5.935000 1.920000 ;
      RECT 5.395000 0.255000 5.585000 1.075000 ;
      RECT 5.675000 1.925000 5.935000 3.075000 ;
  END
END sky130_fd_sc_lp__a32oi_2
