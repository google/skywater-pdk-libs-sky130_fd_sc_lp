* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4b_lp A_N B C D VGND VNB VPB VPWR Y
X0 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR A_N a_87_231# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_251_47# C a_329_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Y a_87_231# a_173_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_509_47# A_N a_87_231# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_87_231# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_329_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_173_47# B a_251_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND A_N a_509_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
