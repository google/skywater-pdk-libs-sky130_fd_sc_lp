* File: sky130_fd_sc_lp__nor4_lp.pxi.spice
* Created: Fri Aug 28 10:57:49 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4_LP%C N_C_M1005_g N_C_M1007_g N_C_c_72_n N_C_M1001_g
+ N_C_c_74_n N_C_c_75_n C C N_C_c_77_n PM_SKY130_FD_SC_LP__NOR4_LP%C
x_PM_SKY130_FD_SC_LP__NOR4_LP%D N_D_M1008_g N_D_M1000_g N_D_M1009_g D D
+ N_D_c_116_n PM_SKY130_FD_SC_LP__NOR4_LP%D
x_PM_SKY130_FD_SC_LP__NOR4_LP%B N_B_c_155_n N_B_M1002_g N_B_c_156_n N_B_c_157_n
+ N_B_c_158_n N_B_M1010_g N_B_c_159_n N_B_M1006_g N_B_c_160_n N_B_c_165_n B B
+ N_B_c_162_n N_B_c_163_n PM_SKY130_FD_SC_LP__NOR4_LP%B
x_PM_SKY130_FD_SC_LP__NOR4_LP%A N_A_c_212_n N_A_M1003_g N_A_M1011_g N_A_c_213_n
+ N_A_M1004_g N_A_c_214_n N_A_c_215_n A A N_A_c_216_n N_A_c_217_n
+ PM_SKY130_FD_SC_LP__NOR4_LP%A
x_PM_SKY130_FD_SC_LP__NOR4_LP%A_27_409# N_A_27_409#_M1005_s N_A_27_409#_M1000_d
+ N_A_27_409#_c_253_n N_A_27_409#_c_254_n N_A_27_409#_c_255_n
+ N_A_27_409#_c_256_n N_A_27_409#_c_257_n N_A_27_409#_c_258_n
+ PM_SKY130_FD_SC_LP__NOR4_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__NOR4_LP%A_134_409# N_A_134_409#_M1005_d
+ N_A_134_409#_M1006_s N_A_134_409#_c_288_n N_A_134_409#_c_289_n
+ N_A_134_409#_c_290_n N_A_134_409#_c_291_n N_A_134_409#_c_292_n
+ PM_SKY130_FD_SC_LP__NOR4_LP%A_134_409#
x_PM_SKY130_FD_SC_LP__NOR4_LP%Y N_Y_M1001_d N_Y_M1010_d N_Y_M1000_s N_Y_c_319_n
+ N_Y_c_320_n N_Y_c_321_n Y Y Y N_Y_c_324_n PM_SKY130_FD_SC_LP__NOR4_LP%Y
x_PM_SKY130_FD_SC_LP__NOR4_LP%VPWR N_VPWR_M1011_d N_VPWR_c_376_n N_VPWR_c_377_n
+ VPWR N_VPWR_c_378_n N_VPWR_c_375_n PM_SKY130_FD_SC_LP__NOR4_LP%VPWR
x_PM_SKY130_FD_SC_LP__NOR4_LP%VGND N_VGND_M1007_s N_VGND_M1009_d N_VGND_M1004_d
+ N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n
+ N_VGND_c_403_n N_VGND_c_404_n VGND N_VGND_c_405_n N_VGND_c_406_n
+ PM_SKY130_FD_SC_LP__NOR4_LP%VGND
cc_1 VNB N_C_M1007_g 0.0430624f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.495
cc_2 VNB N_C_c_72_n 0.0243931f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.185
cc_3 VNB N_C_M1001_g 0.0281687f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.495
cc_4 VNB N_C_c_74_n 0.0149722f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.185
cc_5 VNB N_C_c_75_n 0.00365942f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.78
cc_6 VNB C 0.0327333f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_C_c_77_n 0.0324668f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.275
cc_8 VNB N_D_M1008_g 0.02906f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_9 VNB N_D_M1000_g 0.0015747f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.495
cc_10 VNB N_D_M1009_g 0.0312851f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.11
cc_11 VNB D 0.0208795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_D_c_116_n 0.03839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_155_n 0.0137751f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.78
cc_14 VNB N_B_c_156_n 0.00999536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_157_n 0.00866592f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.11
cc_16 VNB N_B_c_158_n 0.0136612f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.495
cc_17 VNB N_B_c_159_n 0.0269561f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.495
cc_18 VNB N_B_c_160_n 0.00438508f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.615
cc_19 VNB B 0.00187286f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_B_c_162_n 0.0229871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_163_n 0.0176472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_212_n 0.0139219f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.78
cc_23 VNB N_A_c_213_n 0.0179135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_214_n 0.0348663f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.26
cc_25 VNB N_A_c_215_n 0.0279772f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.615
cc_26 VNB N_A_c_216_n 0.0420548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_217_n 0.0318274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_319_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.495
cc_29 VNB N_Y_c_320_n 0.0282352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_321_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.78
cc_31 VNB Y 0.00868308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_375_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_398_n 0.0152105f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.185
cc_34 VNB N_VGND_c_399_n 0.0254175f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.495
cc_35 VNB N_VGND_c_400_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.185
cc_36 VNB N_VGND_c_401_n 0.0113827f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.78
cc_37 VNB N_VGND_c_402_n 0.0249862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_403_n 0.0352526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_404_n 0.00497896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_405_n 0.0352526f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.445
cc_41 VNB N_VGND_c_406_n 0.238962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_C_M1005_g 0.0496714f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_43 VPB N_C_c_75_n 0.0137024f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.78
cc_44 VPB C 0.0107254f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_45 VPB N_D_M1000_g 0.032414f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.495
cc_46 VPB N_B_M1006_g 0.03317f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.26
cc_47 VPB N_B_c_165_n 0.0199171f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.78
cc_48 VPB B 0.00113701f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_49 VPB N_A_M1011_g 0.0474898f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.495
cc_50 VPB N_A_c_215_n 0.00327929f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.615
cc_51 VPB N_A_c_217_n 0.0112757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_27_409#_c_253_n 0.0150561f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.495
cc_53 VPB N_A_27_409#_c_254_n 0.0307705f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.185
cc_54 VPB N_A_27_409#_c_255_n 0.0100264f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.11
cc_55 VPB N_A_27_409#_c_256_n 0.00865023f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.26
cc_56 VPB N_A_27_409#_c_257_n 0.00606349f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_57 VPB N_A_27_409#_c_258_n 0.00152567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_134_409#_c_288_n 0.00868814f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.185
cc_59 VPB N_A_134_409#_c_289_n 0.0392396f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.11
cc_60 VPB N_A_134_409#_c_290_n 0.00244893f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.495
cc_61 VPB N_A_134_409#_c_291_n 0.00246318f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.495
cc_62 VPB N_A_134_409#_c_292_n 0.019902f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.26
cc_63 VPB Y 0.00402901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_Y_c_324_n 0.0111573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_376_n 0.0139087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_377_n 0.0469276f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.495
cc_67 VPB N_VPWR_c_378_n 0.0856465f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.495
cc_68 VPB N_VPWR_c_375_n 0.0766244f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 N_C_M1001_g N_D_M1008_g 0.0158364f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_70 C N_D_M1000_g 5.0219e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_C_c_72_n N_D_c_116_n 0.0158364f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_72 N_C_M1005_g N_A_27_409#_c_253_n 0.00657138f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_73 N_C_c_75_n N_A_27_409#_c_253_n 0.00153853f $X=0.525 $Y=1.78 $X2=0 $Y2=0
cc_74 C N_A_27_409#_c_253_n 0.0225633f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_C_M1005_g N_A_27_409#_c_254_n 0.0185198f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_76 N_C_M1005_g N_A_27_409#_c_255_n 0.0214874f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_77 C N_A_27_409#_c_255_n 0.0158542f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_78 N_C_M1005_g N_A_134_409#_c_288_n 0.00916508f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_79 N_C_M1005_g N_A_134_409#_c_290_n 0.00546325f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_80 N_C_M1007_g N_Y_c_319_n 0.00149969f $X=0.615 $Y=0.495 $X2=0 $Y2=0
cc_81 N_C_M1001_g N_Y_c_319_n 0.00975774f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_82 N_C_M1007_g Y 0.00166508f $X=0.615 $Y=0.495 $X2=0 $Y2=0
cc_83 N_C_c_72_n Y 0.00451298f $X=0.9 $Y=1.185 $X2=0 $Y2=0
cc_84 N_C_M1001_g Y 0.00957333f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_85 C Y 0.0412965f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_86 N_C_c_77_n Y 0.00188972f $X=0.525 $Y=1.275 $X2=0 $Y2=0
cc_87 N_C_M1005_g N_Y_c_324_n 0.00623693f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_88 N_C_c_75_n N_Y_c_324_n 7.73575e-19 $X=0.525 $Y=1.78 $X2=0 $Y2=0
cc_89 C N_Y_c_324_n 0.0121562f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_C_M1005_g N_VPWR_c_378_n 0.00825264f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_91 N_C_M1005_g N_VPWR_c_375_n 0.0164048f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_92 N_C_M1007_g N_VGND_c_399_n 0.0142556f $X=0.615 $Y=0.495 $X2=0 $Y2=0
cc_93 N_C_M1001_g N_VGND_c_399_n 0.002112f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_94 N_C_c_74_n N_VGND_c_399_n 0.00421792f $X=0.525 $Y=1.185 $X2=0 $Y2=0
cc_95 C N_VGND_c_399_n 0.0162621f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_96 N_C_M1007_g N_VGND_c_403_n 0.00445056f $X=0.615 $Y=0.495 $X2=0 $Y2=0
cc_97 N_C_M1001_g N_VGND_c_403_n 0.00502664f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_98 N_C_M1007_g N_VGND_c_406_n 0.00796275f $X=0.615 $Y=0.495 $X2=0 $Y2=0
cc_99 N_C_M1001_g N_VGND_c_406_n 0.00942073f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_100 N_D_M1009_g N_B_c_155_n 0.0204765f $X=1.765 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_101 D N_B_c_157_n 0.00107498f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_102 N_D_M1000_g N_B_c_159_n 0.00548046f $X=1.635 $Y=2.155 $X2=0 $Y2=0
cc_103 D B 0.0204149f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_104 N_D_c_116_n N_B_c_162_n 0.00415374f $X=1.675 $Y=1.29 $X2=0 $Y2=0
cc_105 N_D_M1009_g N_B_c_163_n 0.00415374f $X=1.765 $Y=0.495 $X2=0 $Y2=0
cc_106 D N_B_c_163_n 0.00453211f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_107 N_D_M1000_g N_A_27_409#_c_255_n 0.0221672f $X=1.635 $Y=2.155 $X2=0 $Y2=0
cc_108 N_D_M1000_g N_A_27_409#_c_256_n 0.0144366f $X=1.635 $Y=2.155 $X2=0 $Y2=0
cc_109 D N_A_27_409#_c_256_n 0.0273201f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_110 N_D_c_116_n N_A_27_409#_c_256_n 0.00216661f $X=1.675 $Y=1.29 $X2=0 $Y2=0
cc_111 N_D_M1000_g N_A_27_409#_c_257_n 0.0166032f $X=1.635 $Y=2.155 $X2=0 $Y2=0
cc_112 N_D_M1000_g N_A_27_409#_c_258_n 3.84191e-19 $X=1.635 $Y=2.155 $X2=0 $Y2=0
cc_113 N_D_M1000_g N_A_134_409#_c_288_n 0.00776016f $X=1.635 $Y=2.155 $X2=0
+ $Y2=0
cc_114 N_D_M1000_g N_A_134_409#_c_289_n 0.00814521f $X=1.635 $Y=2.155 $X2=0
+ $Y2=0
cc_115 N_D_M1000_g N_A_134_409#_c_292_n 0.00411381f $X=1.635 $Y=2.155 $X2=0
+ $Y2=0
cc_116 N_D_M1008_g N_Y_c_319_n 0.0099359f $X=1.405 $Y=0.495 $X2=0 $Y2=0
cc_117 N_D_M1009_g N_Y_c_319_n 0.00179788f $X=1.765 $Y=0.495 $X2=0 $Y2=0
cc_118 N_D_M1008_g N_Y_c_320_n 0.0112099f $X=1.405 $Y=0.495 $X2=0 $Y2=0
cc_119 N_D_M1009_g N_Y_c_320_n 0.0111421f $X=1.765 $Y=0.495 $X2=0 $Y2=0
cc_120 D N_Y_c_320_n 0.0563172f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_121 N_D_c_116_n N_Y_c_320_n 7.85225e-19 $X=1.675 $Y=1.29 $X2=0 $Y2=0
cc_122 N_D_M1008_g Y 0.0100883f $X=1.405 $Y=0.495 $X2=0 $Y2=0
cc_123 D Y 0.0245674f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_124 N_D_c_116_n Y 0.00806277f $X=1.675 $Y=1.29 $X2=0 $Y2=0
cc_125 N_D_M1000_g N_Y_c_324_n 0.00697148f $X=1.635 $Y=2.155 $X2=0 $Y2=0
cc_126 D N_Y_c_324_n 0.00179207f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_127 N_D_c_116_n N_Y_c_324_n 0.00652578f $X=1.675 $Y=1.29 $X2=0 $Y2=0
cc_128 N_D_M1008_g N_VGND_c_400_n 0.00175817f $X=1.405 $Y=0.495 $X2=0 $Y2=0
cc_129 N_D_M1009_g N_VGND_c_400_n 0.00984956f $X=1.765 $Y=0.495 $X2=0 $Y2=0
cc_130 N_D_M1008_g N_VGND_c_403_n 0.00502664f $X=1.405 $Y=0.495 $X2=0 $Y2=0
cc_131 N_D_M1009_g N_VGND_c_403_n 0.00445056f $X=1.765 $Y=0.495 $X2=0 $Y2=0
cc_132 N_D_M1008_g N_VGND_c_406_n 0.00553313f $X=1.405 $Y=0.495 $X2=0 $Y2=0
cc_133 N_D_M1009_g N_VGND_c_406_n 0.00409056f $X=1.765 $Y=0.495 $X2=0 $Y2=0
cc_134 N_B_c_158_n N_A_c_212_n 0.00909f $X=2.555 $Y=0.78 $X2=-0.19 $Y2=-0.245
cc_135 N_B_c_165_n N_A_M1011_g 0.0445774f $X=2.665 $Y=1.845 $X2=0 $Y2=0
cc_136 N_B_c_160_n N_A_c_214_n 0.00909f $X=2.555 $Y=0.855 $X2=0 $Y2=0
cc_137 N_B_c_159_n N_A_c_215_n 0.0514503f $X=2.665 $Y=1.66 $X2=0 $Y2=0
cc_138 B N_A_c_215_n 0.00111521f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_139 B N_A_c_216_n 0.00153647f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B_c_162_n N_A_c_216_n 0.00687292f $X=2.645 $Y=1.34 $X2=0 $Y2=0
cc_141 N_B_c_163_n N_A_c_216_n 0.00552324f $X=2.665 $Y=1.175 $X2=0 $Y2=0
cc_142 B N_A_c_217_n 0.0245681f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_143 N_B_c_162_n N_A_c_217_n 0.00236464f $X=2.645 $Y=1.34 $X2=0 $Y2=0
cc_144 N_B_c_163_n N_A_c_217_n 0.00117149f $X=2.665 $Y=1.175 $X2=0 $Y2=0
cc_145 N_B_c_159_n N_A_27_409#_c_256_n 0.00198937f $X=2.665 $Y=1.66 $X2=0 $Y2=0
cc_146 N_B_M1006_g N_A_27_409#_c_256_n 0.00505346f $X=2.725 $Y=2.545 $X2=0 $Y2=0
cc_147 B N_A_27_409#_c_256_n 0.00853202f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_148 N_B_M1006_g N_A_134_409#_c_291_n 0.00427649f $X=2.725 $Y=2.545 $X2=0
+ $Y2=0
cc_149 N_B_M1006_g N_A_134_409#_c_292_n 0.0178221f $X=2.725 $Y=2.545 $X2=0 $Y2=0
cc_150 N_B_c_165_n N_A_134_409#_c_292_n 9.23979e-19 $X=2.665 $Y=1.845 $X2=0
+ $Y2=0
cc_151 B N_A_134_409#_c_292_n 0.0120847f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B_c_155_n N_Y_c_320_n 0.00313643f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_153 N_B_c_156_n N_Y_c_320_n 0.00622831f $X=2.48 $Y=0.855 $X2=0 $Y2=0
cc_154 N_B_c_157_n N_Y_c_320_n 0.00601707f $X=2.27 $Y=0.855 $X2=0 $Y2=0
cc_155 N_B_c_158_n N_Y_c_320_n 0.00274956f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_156 N_B_c_160_n N_Y_c_320_n 0.0038886f $X=2.555 $Y=0.855 $X2=0 $Y2=0
cc_157 B N_Y_c_320_n 0.0217209f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_158 N_B_c_162_n N_Y_c_320_n 0.00319065f $X=2.645 $Y=1.34 $X2=0 $Y2=0
cc_159 N_B_c_163_n N_Y_c_320_n 0.00297679f $X=2.665 $Y=1.175 $X2=0 $Y2=0
cc_160 N_B_c_155_n N_Y_c_321_n 0.00179788f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_161 N_B_c_158_n N_Y_c_321_n 0.0099359f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_162 N_B_M1006_g N_VPWR_c_377_n 0.00519241f $X=2.725 $Y=2.545 $X2=0 $Y2=0
cc_163 N_B_M1006_g N_VPWR_c_378_n 0.0085862f $X=2.725 $Y=2.545 $X2=0 $Y2=0
cc_164 N_B_M1006_g N_VPWR_c_375_n 0.0165862f $X=2.725 $Y=2.545 $X2=0 $Y2=0
cc_165 N_B_c_155_n N_VGND_c_400_n 0.00984956f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_166 N_B_c_158_n N_VGND_c_400_n 0.00175817f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_167 N_B_c_155_n N_VGND_c_405_n 0.00445056f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_168 N_B_c_156_n N_VGND_c_405_n 2.13211e-19 $X=2.48 $Y=0.855 $X2=0 $Y2=0
cc_169 N_B_c_158_n N_VGND_c_405_n 0.00502664f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_170 N_B_c_155_n N_VGND_c_406_n 0.00409056f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_171 N_B_c_158_n N_VGND_c_406_n 0.00553313f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_172 N_A_M1011_g N_A_134_409#_c_291_n 7.28154e-19 $X=3.215 $Y=2.545 $X2=0
+ $Y2=0
cc_173 N_A_M1011_g N_A_134_409#_c_292_n 0.00375854f $X=3.215 $Y=2.545 $X2=0
+ $Y2=0
cc_174 N_A_c_212_n N_Y_c_320_n 2.06353e-19 $X=2.985 $Y=0.785 $X2=0 $Y2=0
cc_175 N_A_c_214_n N_Y_c_320_n 0.00896552f $X=3.355 $Y=0.935 $X2=0 $Y2=0
cc_176 N_A_c_217_n N_Y_c_320_n 0.00240354f $X=3.355 $Y=1.07 $X2=0 $Y2=0
cc_177 N_A_c_212_n N_Y_c_321_n 0.00975774f $X=2.985 $Y=0.785 $X2=0 $Y2=0
cc_178 N_A_c_213_n N_Y_c_321_n 0.00149969f $X=3.345 $Y=0.785 $X2=0 $Y2=0
cc_179 N_A_M1011_g N_VPWR_c_377_n 0.0267797f $X=3.215 $Y=2.545 $X2=0 $Y2=0
cc_180 N_A_c_215_n N_VPWR_c_377_n 8.96377e-19 $X=3.355 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_c_217_n N_VPWR_c_377_n 0.0235305f $X=3.355 $Y=1.07 $X2=0 $Y2=0
cc_182 N_A_M1011_g N_VPWR_c_378_n 0.00802402f $X=3.215 $Y=2.545 $X2=0 $Y2=0
cc_183 N_A_M1011_g N_VPWR_c_375_n 0.0142664f $X=3.215 $Y=2.545 $X2=0 $Y2=0
cc_184 N_A_c_212_n N_VGND_c_402_n 0.002112f $X=2.985 $Y=0.785 $X2=0 $Y2=0
cc_185 N_A_c_213_n N_VGND_c_402_n 0.0140665f $X=3.345 $Y=0.785 $X2=0 $Y2=0
cc_186 N_A_c_214_n N_VGND_c_402_n 0.00312804f $X=3.355 $Y=0.935 $X2=0 $Y2=0
cc_187 N_A_c_217_n N_VGND_c_402_n 0.0279252f $X=3.355 $Y=1.07 $X2=0 $Y2=0
cc_188 N_A_c_212_n N_VGND_c_405_n 0.00502664f $X=2.985 $Y=0.785 $X2=0 $Y2=0
cc_189 N_A_c_213_n N_VGND_c_405_n 0.00445056f $X=3.345 $Y=0.785 $X2=0 $Y2=0
cc_190 N_A_c_212_n N_VGND_c_406_n 0.00942073f $X=2.985 $Y=0.785 $X2=0 $Y2=0
cc_191 N_A_c_213_n N_VGND_c_406_n 0.00796275f $X=3.345 $Y=0.785 $X2=0 $Y2=0
cc_192 N_A_c_214_n N_VGND_c_406_n 6.31283e-19 $X=3.355 $Y=0.935 $X2=0 $Y2=0
cc_193 N_A_27_409#_c_255_n N_A_134_409#_M1005_d 0.00968926f $X=1.735 $Y=2.23
+ $X2=-0.19 $Y2=1.655
cc_194 N_A_27_409#_c_254_n N_A_134_409#_c_288_n 0.0263233f $X=0.28 $Y=2.9 $X2=0
+ $Y2=0
cc_195 N_A_27_409#_c_255_n N_A_134_409#_c_288_n 0.0207591f $X=1.735 $Y=2.23
+ $X2=0 $Y2=0
cc_196 N_A_27_409#_c_255_n N_A_134_409#_c_289_n 0.0222266f $X=1.735 $Y=2.23
+ $X2=0 $Y2=0
cc_197 N_A_27_409#_c_257_n N_A_134_409#_c_289_n 0.0209306f $X=1.9 $Y=2.51 $X2=0
+ $Y2=0
cc_198 N_A_27_409#_c_254_n N_A_134_409#_c_290_n 0.0119061f $X=0.28 $Y=2.9 $X2=0
+ $Y2=0
cc_199 N_A_27_409#_c_256_n N_A_134_409#_c_292_n 0.00805651f $X=1.9 $Y=1.8 $X2=0
+ $Y2=0
cc_200 N_A_27_409#_c_257_n N_A_134_409#_c_292_n 0.0242369f $X=1.9 $Y=2.51 $X2=0
+ $Y2=0
cc_201 N_A_27_409#_c_258_n N_A_134_409#_c_292_n 0.0121616f $X=1.9 $Y=2.23 $X2=0
+ $Y2=0
cc_202 N_A_27_409#_c_255_n N_Y_M1000_s 0.0079226f $X=1.735 $Y=2.23 $X2=0 $Y2=0
cc_203 N_A_27_409#_c_255_n N_Y_c_324_n 0.0335998f $X=1.735 $Y=2.23 $X2=0 $Y2=0
cc_204 N_A_27_409#_c_256_n N_Y_c_324_n 0.0224526f $X=1.9 $Y=1.8 $X2=0 $Y2=0
cc_205 N_A_27_409#_c_254_n N_VPWR_c_378_n 0.0220321f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_206 N_A_27_409#_c_254_n N_VPWR_c_375_n 0.0125808f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_207 N_A_134_409#_c_289_n N_VPWR_c_378_n 0.079983f $X=2.295 $Y=2.98 $X2=0
+ $Y2=0
cc_208 N_A_134_409#_c_290_n N_VPWR_c_378_n 0.0218741f $X=0.975 $Y=2.98 $X2=0
+ $Y2=0
cc_209 N_A_134_409#_c_291_n N_VPWR_c_378_n 0.0221635f $X=2.46 $Y=2.895 $X2=0
+ $Y2=0
cc_210 N_A_134_409#_c_289_n N_VPWR_c_375_n 0.0493242f $X=2.295 $Y=2.98 $X2=0
+ $Y2=0
cc_211 N_A_134_409#_c_290_n N_VPWR_c_375_n 0.0125933f $X=0.975 $Y=2.98 $X2=0
+ $Y2=0
cc_212 N_A_134_409#_c_291_n N_VPWR_c_375_n 0.0126536f $X=2.46 $Y=2.895 $X2=0
+ $Y2=0
cc_213 N_Y_c_319_n N_VGND_c_399_n 0.0153904f $X=1.19 $Y=0.495 $X2=0 $Y2=0
cc_214 N_Y_c_319_n N_VGND_c_400_n 0.0110409f $X=1.19 $Y=0.495 $X2=0 $Y2=0
cc_215 N_Y_c_320_n N_VGND_c_400_n 0.0198622f $X=2.605 $Y=0.86 $X2=0 $Y2=0
cc_216 N_Y_c_321_n N_VGND_c_400_n 0.0110409f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_217 N_Y_c_321_n N_VGND_c_402_n 0.0153904f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_218 N_Y_c_319_n N_VGND_c_403_n 0.021949f $X=1.19 $Y=0.495 $X2=0 $Y2=0
cc_219 N_Y_c_321_n N_VGND_c_405_n 0.021949f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_220 N_Y_c_319_n N_VGND_c_406_n 0.0124703f $X=1.19 $Y=0.495 $X2=0 $Y2=0
cc_221 N_Y_c_320_n N_VGND_c_406_n 0.0312393f $X=2.605 $Y=0.86 $X2=0 $Y2=0
cc_222 N_Y_c_321_n N_VGND_c_406_n 0.0124703f $X=2.77 $Y=0.495 $X2=0 $Y2=0
