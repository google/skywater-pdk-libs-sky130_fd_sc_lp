* NGSPICE file created from sky130_fd_sc_lp__iso0p_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__iso0p_lp2 A SLEEP KAPWR VGND VNB VPB VPWR X
M1000 a_342_417# A a_340_93# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_602_93# a_342_417# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.759e+11p ps=3.47e+06u
M1002 X a_342_417# a_602_93# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 VGND SLEEP a_112_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 a_340_93# a_27_93# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 KAPWR A a_342_417# VPB phighvt w=1e+06u l=250000u
+  ad=1.66e+12p pd=7.32e+06u as=3e+11p ps=2.6e+06u
M1006 X a_342_417# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1007 KAPWR SLEEP a_27_93# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1008 a_112_93# SLEEP a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1009 a_342_417# a_27_93# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

