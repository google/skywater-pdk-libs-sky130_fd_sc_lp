* File: sky130_fd_sc_lp__einvp_0.pxi.spice
* Created: Fri Aug 28 10:33:35 2020
* 
x_PM_SKY130_FD_SC_LP__EINVP_0%TE N_TE_c_38_n N_TE_M1003_g N_TE_M1000_g
+ N_TE_M1004_g N_TE_c_40_n N_TE_c_41_n TE TE TE N_TE_c_43_n
+ PM_SKY130_FD_SC_LP__EINVP_0%TE
x_PM_SKY130_FD_SC_LP__EINVP_0%A_32_70# N_A_32_70#_M1003_s N_A_32_70#_M1000_s
+ N_A_32_70#_M1002_g N_A_32_70#_c_77_n N_A_32_70#_c_80_n N_A_32_70#_c_81_n
+ N_A_32_70#_c_82_n N_A_32_70#_c_83_n PM_SKY130_FD_SC_LP__EINVP_0%A_32_70#
x_PM_SKY130_FD_SC_LP__EINVP_0%A N_A_M1005_g N_A_M1001_g A A A A N_A_c_115_n
+ N_A_c_116_n PM_SKY130_FD_SC_LP__EINVP_0%A
x_PM_SKY130_FD_SC_LP__EINVP_0%VPWR N_VPWR_M1000_d N_VPWR_c_145_n VPWR
+ N_VPWR_c_146_n N_VPWR_c_147_n N_VPWR_c_144_n N_VPWR_c_149_n
+ PM_SKY130_FD_SC_LP__EINVP_0%VPWR
x_PM_SKY130_FD_SC_LP__EINVP_0%Z N_Z_M1005_d N_Z_M1001_d N_Z_c_170_n N_Z_c_171_n
+ Z Z N_Z_c_174_n PM_SKY130_FD_SC_LP__EINVP_0%Z
x_PM_SKY130_FD_SC_LP__EINVP_0%VGND N_VGND_M1003_d N_VGND_c_204_n VGND
+ N_VGND_c_205_n N_VGND_c_206_n N_VGND_c_207_n N_VGND_c_208_n
+ PM_SKY130_FD_SC_LP__EINVP_0%VGND
cc_1 VNB N_TE_c_38_n 0.0365372f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.88
cc_2 VNB N_TE_M1000_g 0.00684225f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.85
cc_3 VNB N_TE_c_40_n 0.0259053f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.03
cc_4 VNB N_TE_c_41_n 0.0230613f $X=-0.19 $Y=-0.245 $X2=0.622 $Y2=1.55
cc_5 VNB TE 0.00741257f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_TE_c_43_n 0.0268465f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.045
cc_7 VNB N_A_32_70#_c_77_n 0.0604144f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.03
cc_8 VNB N_A_M1001_g 0.00685791f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.85
cc_9 VNB A 0.0344399f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.88
cc_10 VNB N_A_c_115_n 0.0965592f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_A_c_116_n 0.0219716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_144_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_Z_c_170_n 0.00715071f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.88
cc_14 VNB N_Z_c_171_n 0.0165509f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.88
cc_15 VNB N_VGND_c_204_n 0.00344978f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.85
cc_16 VNB N_VGND_c_205_n 0.0175105f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.56
cc_17 VNB N_VGND_c_206_n 0.0310079f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_18 VNB N_VGND_c_207_n 0.144886f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_19 VNB N_VGND_c_208_n 0.00579822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VPB N_TE_M1000_g 0.0760796f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.85
cc_21 VPB TE 0.00379041f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_22 VPB N_A_32_70#_M1002_g 0.0197405f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.56
cc_23 VPB N_A_32_70#_c_77_n 0.0139164f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.03
cc_24 VPB N_A_32_70#_c_80_n 0.0306948f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_25 VPB N_A_32_70#_c_81_n 0.00468694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_A_32_70#_c_82_n 0.039012f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.045
cc_27 VPB N_A_32_70#_c_83_n 0.0167985f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.045
cc_28 VPB N_A_M1001_g 0.0604245f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.85
cc_29 VPB A 0.026022f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.88
cc_30 VPB N_VPWR_c_145_n 0.00619582f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.85
cc_31 VPB N_VPWR_c_146_n 0.0191288f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.56
cc_32 VPB N_VPWR_c_147_n 0.0278089f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_33 VPB N_VPWR_c_144_n 0.0569614f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_34 VPB N_VPWR_c_149_n 0.00585466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_Z_c_170_n 0.00603309f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.88
cc_36 VPB Z 0.016003f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.353
cc_37 VPB N_Z_c_174_n 0.0261107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 N_TE_M1000_g N_A_32_70#_M1002_g 0.0161622f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_39 N_TE_c_38_n N_A_32_70#_c_77_n 0.034645f $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_40 TE N_A_32_70#_c_77_n 0.0680504f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_41 N_TE_M1000_g N_A_32_70#_c_80_n 0.0175572f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_42 N_TE_M1000_g N_A_32_70#_c_81_n 0.0181449f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_43 N_TE_c_41_n N_A_32_70#_c_81_n 9.99002e-19 $X=0.622 $Y=1.55 $X2=0 $Y2=0
cc_44 TE N_A_32_70#_c_81_n 0.030134f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_45 N_TE_M1000_g N_A_32_70#_c_82_n 0.0213328f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_46 N_TE_c_41_n N_A_32_70#_c_82_n 9.88495e-19 $X=0.622 $Y=1.55 $X2=0 $Y2=0
cc_47 TE N_A_32_70#_c_82_n 0.00270081f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_48 N_TE_M1000_g N_A_32_70#_c_83_n 0.00874187f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_49 TE N_A_M1001_g 0.00106334f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_50 N_TE_c_40_n N_A_c_115_n 0.020887f $X=0.715 $Y=1.03 $X2=0 $Y2=0
cc_51 TE N_A_c_115_n 0.00203146f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_52 N_TE_c_43_n N_A_c_115_n 0.013234f $X=0.655 $Y=1.045 $X2=0 $Y2=0
cc_53 N_TE_c_38_n N_A_c_116_n 0.020887f $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_54 N_TE_M1000_g N_VPWR_c_145_n 0.0073464f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_55 N_TE_M1000_g N_VPWR_c_146_n 0.00517695f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_56 N_TE_M1000_g N_VPWR_c_144_n 0.0105249f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_57 N_TE_c_38_n N_Z_c_170_n 0.00293284f $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_58 N_TE_M1000_g N_Z_c_170_n 0.00453826f $X=0.5 $Y=2.85 $X2=0 $Y2=0
cc_59 TE N_Z_c_170_n 0.0507761f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_60 N_TE_c_43_n N_Z_c_170_n 0.00156975f $X=0.655 $Y=1.045 $X2=0 $Y2=0
cc_61 N_TE_c_38_n N_Z_c_171_n 9.38751e-19 $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_62 N_TE_c_38_n N_VGND_c_204_n 0.0217259f $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_63 N_TE_c_40_n N_VGND_c_204_n 7.02505e-19 $X=0.715 $Y=1.03 $X2=0 $Y2=0
cc_64 TE N_VGND_c_204_n 0.0230233f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_65 N_TE_c_38_n N_VGND_c_205_n 0.00396895f $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_66 N_TE_c_38_n N_VGND_c_206_n 0.00396895f $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_67 N_TE_c_38_n N_VGND_c_207_n 0.0142591f $X=0.5 $Y=0.88 $X2=0 $Y2=0
cc_68 TE N_VGND_c_207_n 0.00257162f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_69 N_A_32_70#_M1002_g N_A_M1001_g 0.0464487f $X=1.025 $Y=2.74 $X2=0 $Y2=0
cc_70 N_A_32_70#_c_81_n N_A_M1001_g 2.84118e-19 $X=0.95 $Y=2.095 $X2=0 $Y2=0
cc_71 N_A_32_70#_c_82_n N_A_M1001_g 0.0186135f $X=0.95 $Y=2.095 $X2=0 $Y2=0
cc_72 N_A_32_70#_M1002_g N_VPWR_c_145_n 0.0152622f $X=1.025 $Y=2.74 $X2=0 $Y2=0
cc_73 N_A_32_70#_c_80_n N_VPWR_c_145_n 0.0307426f $X=0.285 $Y=2.85 $X2=0 $Y2=0
cc_74 N_A_32_70#_c_81_n N_VPWR_c_145_n 0.0272719f $X=0.95 $Y=2.095 $X2=0 $Y2=0
cc_75 N_A_32_70#_c_82_n N_VPWR_c_145_n 0.0036701f $X=0.95 $Y=2.095 $X2=0 $Y2=0
cc_76 N_A_32_70#_c_80_n N_VPWR_c_146_n 0.0151997f $X=0.285 $Y=2.85 $X2=0 $Y2=0
cc_77 N_A_32_70#_M1002_g N_VPWR_c_147_n 0.00456975f $X=1.025 $Y=2.74 $X2=0 $Y2=0
cc_78 N_A_32_70#_M1002_g N_VPWR_c_144_n 0.00811515f $X=1.025 $Y=2.74 $X2=0 $Y2=0
cc_79 N_A_32_70#_c_80_n N_VPWR_c_144_n 0.0122376f $X=0.285 $Y=2.85 $X2=0 $Y2=0
cc_80 N_A_32_70#_M1002_g N_Z_c_170_n 6.61652e-19 $X=1.025 $Y=2.74 $X2=0 $Y2=0
cc_81 N_A_32_70#_c_81_n N_Z_c_170_n 0.0263181f $X=0.95 $Y=2.095 $X2=0 $Y2=0
cc_82 N_A_32_70#_c_82_n N_Z_c_170_n 0.0021636f $X=0.95 $Y=2.095 $X2=0 $Y2=0
cc_83 N_A_32_70#_M1002_g Z 0.00441959f $X=1.025 $Y=2.74 $X2=0 $Y2=0
cc_84 N_A_32_70#_M1002_g N_Z_c_174_n 0.00165448f $X=1.025 $Y=2.74 $X2=0 $Y2=0
cc_85 N_A_32_70#_c_77_n N_VGND_c_205_n 0.00930971f $X=0.285 $Y=0.56 $X2=0 $Y2=0
cc_86 N_A_32_70#_c_77_n N_VGND_c_207_n 0.00926582f $X=0.285 $Y=0.56 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_VPWR_c_145_n 0.00261767f $X=1.415 $Y=2.74 $X2=0 $Y2=0
cc_88 N_A_M1001_g N_VPWR_c_147_n 0.00515911f $X=1.415 $Y=2.74 $X2=0 $Y2=0
cc_89 N_A_M1001_g N_VPWR_c_144_n 0.00668383f $X=1.415 $Y=2.74 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_Z_c_170_n 0.0228428f $X=1.415 $Y=2.74 $X2=0 $Y2=0
cc_91 A N_Z_c_170_n 0.0886707f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A_c_115_n N_Z_c_170_n 0.0248281f $X=1.65 $Y=1.045 $X2=0 $Y2=0
cc_93 N_A_c_116_n N_Z_c_170_n 0.0107368f $X=1.53 $Y=0.88 $X2=0 $Y2=0
cc_94 A N_Z_c_171_n 0.011403f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_95 N_A_c_115_n N_Z_c_171_n 0.00701437f $X=1.65 $Y=1.045 $X2=0 $Y2=0
cc_96 N_A_c_116_n N_Z_c_171_n 0.00823877f $X=1.53 $Y=0.88 $X2=0 $Y2=0
cc_97 N_A_M1001_g Z 0.0147305f $X=1.415 $Y=2.74 $X2=0 $Y2=0
cc_98 A Z 0.0228888f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_99 N_A_M1001_g N_Z_c_174_n 0.0102489f $X=1.415 $Y=2.74 $X2=0 $Y2=0
cc_100 N_A_c_116_n N_VGND_c_204_n 0.00101031f $X=1.53 $Y=0.88 $X2=0 $Y2=0
cc_101 N_A_c_116_n N_VGND_c_206_n 0.00301434f $X=1.53 $Y=0.88 $X2=0 $Y2=0
cc_102 A N_VGND_c_207_n 0.00553089f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A_c_116_n N_VGND_c_207_n 0.00412668f $X=1.53 $Y=0.88 $X2=0 $Y2=0
cc_104 N_VPWR_c_145_n Z 0.0038559f $X=0.81 $Y=2.575 $X2=0 $Y2=0
cc_105 N_VPWR_c_144_n Z 0.00826198f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_106 N_VPWR_c_145_n N_Z_c_174_n 0.018801f $X=0.81 $Y=2.575 $X2=0 $Y2=0
cc_107 N_VPWR_c_147_n N_Z_c_174_n 0.026f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_108 N_VPWR_c_144_n N_Z_c_174_n 0.0141411f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_109 A_220_484# Z 0.00229738f $X=1.1 $Y=2.42 $X2=1.595 $Y2=2.32
cc_110 N_Z_c_171_n N_VGND_c_204_n 0.00756955f $X=1.535 $Y=0.505 $X2=0 $Y2=0
cc_111 N_Z_c_171_n N_VGND_c_206_n 0.0213423f $X=1.535 $Y=0.505 $X2=0 $Y2=0
cc_112 N_Z_c_171_n N_VGND_c_207_n 0.0172435f $X=1.535 $Y=0.505 $X2=0 $Y2=0
