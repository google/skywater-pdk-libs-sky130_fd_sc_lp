# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2111o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a2111o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.695000 1.210000 5.170000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.340000 1.210000 5.850000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.335000 4.165000 1.535000 ;
        RECT 3.375000 1.535000 4.165000 1.785000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.425000 2.795000 1.770000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.425000 0.535000 1.750000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.390000 0.255000 6.580000 1.065000 ;
        RECT 6.390000 1.065000 8.075000 1.235000 ;
        RECT 6.390000 1.745000 8.075000 1.925000 ;
        RECT 6.390000 1.925000 6.580000 3.075000 ;
        RECT 7.250000 0.255000 7.440000 1.065000 ;
        RECT 7.250000 1.925000 7.440000 3.075000 ;
        RECT 7.715000 1.235000 8.075000 1.745000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.775000  0.085000 1.105000 0.885000 ;
        RECT 1.675000  0.085000 2.005000 0.815000 ;
        RECT 2.575000  0.085000 3.510000 0.815000 ;
        RECT 5.030000  0.085000 5.360000 0.590000 ;
        RECT 5.890000  0.085000 6.220000 1.040000 ;
        RECT 6.750000  0.085000 7.080000 0.895000 ;
        RECT 7.610000  0.085000 7.940000 0.895000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 4.040000 2.295000 4.370000 3.245000 ;
        RECT 5.030000 2.295000 5.360000 3.245000 ;
        RECT 5.890000 1.955000 6.220000 3.245000 ;
        RECT 6.750000 2.095000 7.080000 3.245000 ;
        RECT 7.610000 2.105000 7.940000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.275000 1.920000 0.535000 2.905000 ;
      RECT 0.275000 2.905000 2.325000 3.075000 ;
      RECT 0.345000 0.255000 0.605000 1.065000 ;
      RECT 0.345000 1.065000 4.515000 1.155000 ;
      RECT 0.345000 1.155000 1.455000 1.235000 ;
      RECT 0.705000 1.235000 0.935000 1.930000 ;
      RECT 0.705000 1.930000 1.035000 2.735000 ;
      RECT 1.205000 1.940000 1.395000 2.905000 ;
      RECT 1.275000 0.255000 1.505000 0.985000 ;
      RECT 1.275000 0.985000 4.515000 1.065000 ;
      RECT 1.565000 1.940000 3.205000 2.110000 ;
      RECT 1.565000 2.110000 1.895000 2.735000 ;
      RECT 2.065000 2.280000 2.325000 2.905000 ;
      RECT 2.175000 0.255000 2.405000 0.985000 ;
      RECT 2.515000 2.280000 2.845000 2.905000 ;
      RECT 2.515000 2.905000 3.825000 3.075000 ;
      RECT 2.965000 1.705000 3.205000 1.940000 ;
      RECT 3.015000 2.110000 3.205000 2.735000 ;
      RECT 3.495000 1.955000 5.720000 2.125000 ;
      RECT 3.495000 2.125000 3.825000 2.905000 ;
      RECT 3.680000 0.255000 4.800000 0.465000 ;
      RECT 3.680000 0.465000 3.870000 0.985000 ;
      RECT 4.040000 0.635000 4.860000 0.760000 ;
      RECT 4.040000 0.760000 5.720000 0.815000 ;
      RECT 4.345000 1.155000 4.515000 1.615000 ;
      RECT 4.345000 1.615000 6.200000 1.785000 ;
      RECT 4.540000 2.125000 4.800000 3.025000 ;
      RECT 4.685000 0.815000 5.720000 1.040000 ;
      RECT 5.530000 0.255000 5.720000 0.760000 ;
      RECT 5.530000 2.125000 5.720000 3.075000 ;
      RECT 6.020000 1.405000 7.545000 1.575000 ;
      RECT 6.020000 1.575000 6.200000 1.615000 ;
  END
END sky130_fd_sc_lp__a2111o_4
