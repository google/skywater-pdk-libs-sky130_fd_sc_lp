* File: sky130_fd_sc_lp__busreceiver_0.spice
* Created: Fri Aug 28 10:14:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__busreceiver_0.pex.spice"
.subckt sky130_fd_sc_lp__busreceiver_0  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_70_157#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0714 AS=0.1113 PD=0.76 PS=1.37 NRD=9.996 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_70_157#_M1000_d N_A_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0714 PD=1.37 PS=0.76 NRD=0 NRS=7.14 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_70_157#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.121419 AS=0.1696 PD=1.1834 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.5 A=0.096 P=1.58 MULT=1
MM1002 N_A_70_157#_M1002_d N_A_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0796811 PD=1.37 PS=0.776604 NRD=0 NRS=29.3136 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__busreceiver_0.pxi.spice"
*
.ends
*
*
