* NGSPICE file created from sky130_fd_sc_lp__a41o_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a41o_m A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_300_508# VPB phighvt w=420000u l=150000u
+  ad=3.465e+11p pd=4.17e+06u as=3.465e+11p ps=4.17e+06u
M1001 a_335_47# A1 a_80_153# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.407e+11p ps=1.51e+06u
M1002 a_300_508# B1 a_80_153# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VPWR A3 a_300_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_80_153# B1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1005 VGND A4 a_551_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_443_47# A2 a_335_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1007 a_300_508# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_551_47# A3 a_443_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_80_153# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1010 VGND a_80_153# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 a_300_508# A4 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

