* File: sky130_fd_sc_lp__nor3b_4.spice
* Created: Fri Aug 28 10:56:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor3b_4.pex.spice"
.subckt sky130_fd_sc_lp__nor3b_4  VNB VPB C_N A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_C_N_M1007_g N_A_38_367#_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.2226 PD=1.2 PS=2.21 NRD=6.42 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005.6 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=4.992 M=1 R=5.6 SA=75000.7 SB=75005.1
+ A=0.126 P=1.98 MULT=1
MM1016 N_Y_M1005_d N_A_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=5.712 M=1 R=5.6 SA=75001.1 SB=75004.7
+ A=0.126 P=1.98 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=5.712 M=1 R=5.6 SA=75001.6 SB=75004.2
+ A=0.126 P=1.98 MULT=1
MM1025 N_Y_M1017_d N_A_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1 SB=75003.8 A=0.126
+ P=1.98 MULT=1
MM1002 N_VGND_M1025_s N_A_38_367#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A_38_367#_M1003_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1003_d N_A_38_367#_M1015_g N_Y_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.4
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1022_d N_A_38_367#_M1022_g N_Y_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1722 AS=0.1176 PD=1.25 PS=1.12 NRD=9.276 NRS=0 M=1 R=5.6 SA=75003.8
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1722 PD=1.12 PS=1.25 NRD=0 NRS=9.276 M=1 R=5.6 SA=75004.3 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1004_d N_B_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.8 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1010 N_Y_M1010_d N_B_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.2 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1019 N_Y_M1010_d N_B_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75005.6 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_C_N_M1013_g N_A_38_367#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75000.2 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1001 N_A_211_367#_M1001_d N_A_M1001_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1014 N_A_211_367#_M1001_d N_A_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1020 N_A_211_367#_M1020_d N_A_M1020_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1021 N_A_211_367#_M1020_d N_A_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A_38_367#_M1006_g N_A_576_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1006_d N_A_38_367#_M1011_g N_A_576_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1018 N_Y_M1018_d N_A_38_367#_M1018_g N_A_576_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1023 N_Y_M1018_d N_A_38_367#_M1023_g N_A_576_367#_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1000 N_A_576_367#_M1023_s N_B_M1000_g N_A_211_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_A_576_367#_M1008_d N_B_M1008_g N_A_211_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1012 N_A_576_367#_M1008_d N_B_M1012_g N_A_211_367#_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1024 N_A_576_367#_M1024_d N_B_M1024_g N_A_211_367#_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__nor3b_4.pxi.spice"
*
.ends
*
*
