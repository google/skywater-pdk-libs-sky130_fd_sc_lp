* File: sky130_fd_sc_lp__fa_2.pxi.spice
* Created: Fri Aug 28 10:34:52 2020
* 
x_PM_SKY130_FD_SC_LP__FA_2%A_84_21# N_A_84_21#_M1019_d N_A_84_21#_M1017_d
+ N_A_84_21#_M1007_g N_A_84_21#_M1020_g N_A_84_21#_c_177_n N_A_84_21#_M1008_g
+ N_A_84_21#_M1030_g N_A_84_21#_c_179_n N_A_84_21#_c_180_n N_A_84_21#_c_181_n
+ N_A_84_21#_c_182_n N_A_84_21#_c_183_n N_A_84_21#_c_191_n N_A_84_21#_c_192_n
+ N_A_84_21#_c_184_n N_A_84_21#_c_212_p N_A_84_21#_c_193_n N_A_84_21#_c_185_n
+ N_A_84_21#_c_186_n N_A_84_21#_c_194_n N_A_84_21#_c_195_n
+ PM_SKY130_FD_SC_LP__FA_2%A_84_21#
x_PM_SKY130_FD_SC_LP__FA_2%A N_A_M1012_g N_A_M1001_g N_A_M1002_g N_A_M1010_g
+ N_A_M1021_g N_A_M1026_g N_A_M1009_g N_A_M1025_g N_A_c_330_n N_A_c_331_n
+ N_A_c_332_n N_A_c_343_n N_A_c_344_n N_A_c_345_n N_A_c_387_p N_A_c_346_n
+ N_A_c_389_p N_A_c_333_n N_A_c_334_n N_A_c_348_n N_A_c_349_n A N_A_c_335_n
+ N_A_c_336_n N_A_c_337_n PM_SKY130_FD_SC_LP__FA_2%A
x_PM_SKY130_FD_SC_LP__FA_2%A_395_398# N_A_395_398#_M1018_d N_A_395_398#_M1006_d
+ N_A_395_398#_M1011_d N_A_395_398#_M1014_d N_A_395_398#_M1022_g
+ N_A_395_398#_M1031_g N_A_395_398#_c_537_n N_A_395_398#_M1004_g
+ N_A_395_398#_M1003_g N_A_395_398#_c_539_n N_A_395_398#_M1016_g
+ N_A_395_398#_M1028_g N_A_395_398#_c_541_n N_A_395_398#_c_542_n
+ N_A_395_398#_c_543_n N_A_395_398#_c_576_n N_A_395_398#_c_577_n
+ N_A_395_398#_c_544_n N_A_395_398#_c_545_n N_A_395_398#_c_546_n
+ N_A_395_398#_c_547_n N_A_395_398#_c_580_n N_A_395_398#_c_548_n
+ N_A_395_398#_c_558_n N_A_395_398#_c_559_n N_A_395_398#_c_549_n
+ N_A_395_398#_c_550_n N_A_395_398#_c_560_n N_A_395_398#_c_601_n
+ N_A_395_398#_c_561_n N_A_395_398#_c_562_n N_A_395_398#_c_563_n
+ N_A_395_398#_c_551_n N_A_395_398#_c_565_n N_A_395_398#_c_552_n
+ N_A_395_398#_c_553_n PM_SKY130_FD_SC_LP__FA_2%A_395_398#
x_PM_SKY130_FD_SC_LP__FA_2%CIN N_CIN_M1011_g N_CIN_M1018_g N_CIN_c_814_n
+ N_CIN_c_815_n N_CIN_c_816_n N_CIN_M1019_g N_CIN_M1017_g N_CIN_c_818_n
+ N_CIN_M1015_g N_CIN_M1005_g N_CIN_c_820_n N_CIN_c_810_n CIN N_CIN_c_812_n
+ PM_SKY130_FD_SC_LP__FA_2%CIN
x_PM_SKY130_FD_SC_LP__FA_2%B N_B_M1023_g N_B_M1027_g N_B_c_917_n N_B_c_918_n
+ N_B_M1029_g N_B_M1013_g N_B_c_920_n N_B_c_921_n N_B_M1000_g N_B_M1024_g
+ N_B_M1006_g N_B_M1014_g N_B_c_925_n N_B_c_926_n N_B_c_927_n N_B_c_928_n
+ N_B_c_975_n N_B_c_929_n B N_B_c_931_n N_B_c_932_n PM_SKY130_FD_SC_LP__FA_2%B
x_PM_SKY130_FD_SC_LP__FA_2%VPWR N_VPWR_M1020_s N_VPWR_M1030_s N_VPWR_M1012_d
+ N_VPWR_M1005_d N_VPWR_M1021_d N_VPWR_M1028_s N_VPWR_c_1084_n N_VPWR_c_1085_n
+ N_VPWR_c_1086_n N_VPWR_c_1087_n N_VPWR_c_1088_n N_VPWR_c_1121_n
+ N_VPWR_c_1089_n N_VPWR_c_1090_n N_VPWR_c_1091_n VPWR N_VPWR_c_1092_n
+ N_VPWR_c_1093_n N_VPWR_c_1094_n N_VPWR_c_1095_n N_VPWR_c_1096_n
+ N_VPWR_c_1083_n N_VPWR_c_1098_n N_VPWR_c_1099_n N_VPWR_c_1100_n
+ N_VPWR_c_1101_n PM_SKY130_FD_SC_LP__FA_2%VPWR
x_PM_SKY130_FD_SC_LP__FA_2%SUM N_SUM_M1007_s N_SUM_M1020_d N_SUM_c_1216_n
+ N_SUM_c_1219_n N_SUM_c_1220_n N_SUM_c_1232_n SUM SUM SUM SUM SUM
+ N_SUM_c_1212_n SUM PM_SKY130_FD_SC_LP__FA_2%SUM
x_PM_SKY130_FD_SC_LP__FA_2%A_309_398# N_A_309_398#_M1027_d N_A_309_398#_M1012_s
+ N_A_309_398#_c_1262_n N_A_309_398#_c_1263_n N_A_309_398#_c_1264_n
+ N_A_309_398#_c_1265_n PM_SKY130_FD_SC_LP__FA_2%A_309_398#
x_PM_SKY130_FD_SC_LP__FA_2%A_941_419# N_A_941_419#_M1031_d N_A_941_419#_M1000_d
+ N_A_941_419#_c_1301_n N_A_941_419#_c_1297_n N_A_941_419#_c_1298_n
+ N_A_941_419#_c_1299_n PM_SKY130_FD_SC_LP__FA_2%A_941_419#
x_PM_SKY130_FD_SC_LP__FA_2%COUT N_COUT_M1004_d N_COUT_M1003_d COUT COUT
+ N_COUT_c_1333_n COUT PM_SKY130_FD_SC_LP__FA_2%COUT
x_PM_SKY130_FD_SC_LP__FA_2%VGND N_VGND_M1007_d N_VGND_M1008_d N_VGND_M1001_d
+ N_VGND_M1015_d N_VGND_M1026_d N_VGND_M1016_s N_VGND_c_1366_n N_VGND_c_1367_n
+ N_VGND_c_1368_n N_VGND_c_1369_n N_VGND_c_1370_n N_VGND_c_1371_n
+ N_VGND_c_1372_n N_VGND_c_1373_n N_VGND_c_1374_n N_VGND_c_1375_n VGND
+ N_VGND_c_1376_n N_VGND_c_1377_n N_VGND_c_1378_n N_VGND_c_1379_n
+ N_VGND_c_1380_n N_VGND_c_1381_n N_VGND_c_1382_n PM_SKY130_FD_SC_LP__FA_2%VGND
x_PM_SKY130_FD_SC_LP__FA_2%A_309_131# N_A_309_131#_M1023_d N_A_309_131#_M1001_s
+ N_A_309_131#_c_1473_n N_A_309_131#_c_1474_n N_A_309_131#_c_1475_n
+ PM_SKY130_FD_SC_LP__FA_2%A_309_131#
x_PM_SKY130_FD_SC_LP__FA_2%A_940_119# N_A_940_119#_M1022_d N_A_940_119#_M1024_d
+ N_A_940_119#_c_1509_n N_A_940_119#_c_1501_n N_A_940_119#_c_1502_n
+ N_A_940_119#_c_1519_n PM_SKY130_FD_SC_LP__FA_2%A_940_119#
cc_1 VNB N_A_84_21#_M1007_g 0.0268962f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_A_84_21#_M1020_g 0.00805423f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_A_84_21#_c_177_n 0.0316066f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.42
cc_4 VNB N_A_84_21#_M1008_g 0.0246956f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_5 VNB N_A_84_21#_c_179_n 0.00616449f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.42
cc_6 VNB N_A_84_21#_c_180_n 0.00466715f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.51
cc_7 VNB N_A_84_21#_c_181_n 0.0294639f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=1.315
cc_8 VNB N_A_84_21#_c_182_n 0.00490696f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.785
cc_9 VNB N_A_84_21#_c_183_n 0.00701348f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=1.17
cc_10 VNB N_A_84_21#_c_184_n 0.00372363f $X=-0.19 $Y=-0.245 $X2=3.715 $Y2=0.805
cc_11 VNB N_A_84_21#_c_185_n 0.00458615f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.315
cc_12 VNB N_A_84_21#_c_186_n 0.00642311f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.17
cc_13 VNB N_A_M1001_g 0.0312956f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_14 VNB N_A_M1002_g 0.0236472f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.495
cc_15 VNB N_A_M1026_g 0.0466359f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_16 VNB N_A_M1009_g 0.0229012f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.51
cc_17 VNB N_A_c_330_n 0.0110273f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.4
cc_18 VNB N_A_c_331_n 0.0108472f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.87
cc_19 VNB N_A_c_332_n 8.71732e-19 $X=-0.19 $Y=-0.245 $X2=4.41 $Y2=0.805
cc_20 VNB N_A_c_333_n 0.00666738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_334_n 0.00827158f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=1.17
cc_22 VNB N_A_c_335_n 0.0356948f $X=-0.19 $Y=-0.245 $X2=1.017 $Y2=1.675
cc_23 VNB N_A_c_336_n 0.023246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_337_n 0.00502186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_395_398#_M1022_g 0.041981f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.42
cc_26 VNB N_A_395_398#_c_537_n 0.0190105f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.675
cc_27 VNB N_A_395_398#_M1003_g 0.0138665f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.51
cc_28 VNB N_A_395_398#_c_539_n 0.019495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_395_398#_M1028_g 0.00627073f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=1.17
cc_30 VNB N_A_395_398#_c_541_n 0.00957461f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=1.87
cc_31 VNB N_A_395_398#_c_542_n 0.00213435f $X=-0.19 $Y=-0.245 $X2=3.715
+ $Y2=0.805
cc_32 VNB N_A_395_398#_c_543_n 0.00588479f $X=-0.19 $Y=-0.245 $X2=4.41 $Y2=0.805
cc_33 VNB N_A_395_398#_c_544_n 0.00253172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_395_398#_c_545_n 0.0428223f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.51
cc_35 VNB N_A_395_398#_c_546_n 0.0138506f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.17
cc_36 VNB N_A_395_398#_c_547_n 6.43948e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_395_398#_c_548_n 0.00327046f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=0.805
cc_38 VNB N_A_395_398#_c_549_n 0.00442974f $X=-0.19 $Y=-0.245 $X2=4.375 $Y2=2.16
cc_39 VNB N_A_395_398#_c_550_n 0.0161719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_395_398#_c_551_n 0.0112182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_395_398#_c_552_n 0.0121213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_395_398#_c_553_n 0.0230931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_CIN_M1018_g 0.0425412f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_44 VNB N_CIN_M1019_g 0.0399556f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.42
cc_45 VNB N_CIN_M1015_g 0.0209054f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_46 VNB N_CIN_M1005_g 0.0120675f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.51
cc_47 VNB N_CIN_c_810_n 0.0238819f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.315
cc_48 VNB CIN 0.00146022f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.785
cc_49 VNB N_CIN_c_812_n 0.029891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_B_M1023_g 0.0583565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_B_c_917_n 0.154681f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_52 VNB N_B_c_918_n 0.0102351f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_53 VNB N_B_M1029_g 0.0537657f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.495
cc_54 VNB N_B_c_920_n 0.144464f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.42
cc_55 VNB N_B_c_921_n 0.0411915f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.345
cc_56 VNB N_B_M1024_g 0.0305325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_B_M1006_g 0.0118276f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.51
cc_58 VNB N_B_M1014_g 0.0154476f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=1.315
cc_59 VNB N_B_c_925_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.4
cc_60 VNB N_B_c_926_n 0.0103654f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=1.17
cc_61 VNB N_B_c_927_n 0.0172651f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.17
cc_62 VNB N_B_c_928_n 0.0046517f $X=-0.19 $Y=-0.245 $X2=3.715 $Y2=0.805
cc_63 VNB N_B_c_929_n 0.00101098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB B 0.0195169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_B_c_931_n 0.0534397f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=0.805
cc_66 VNB N_B_c_932_n 0.00844734f $X=-0.19 $Y=-0.245 $X2=3.69 $Y2=1.87
cc_67 VNB N_VPWR_c_1083_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_SUM_c_1212_n 0.00857636f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=1.315
cc_69 VNB SUM 0.035907f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.785
cc_70 VNB N_COUT_c_1333_n 0.0014272f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_71 VNB COUT 0.00263891f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_72 VNB N_VGND_c_1366_n 0.0107277f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_73 VNB N_VGND_c_1367_n 0.0168434f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.675
cc_74 VNB N_VGND_c_1368_n 0.00876047f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.42
cc_75 VNB N_VGND_c_1369_n 0.0109825f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.51
cc_76 VNB N_VGND_c_1370_n 0.0107524f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.4
cc_77 VNB N_VGND_c_1371_n 0.0186799f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=1.17
cc_78 VNB N_VGND_c_1372_n 0.047239f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.87
cc_79 VNB N_VGND_c_1373_n 0.00279655f $X=-0.19 $Y=-0.245 $X2=3.715 $Y2=0.805
cc_80 VNB N_VGND_c_1374_n 0.013424f $X=-0.19 $Y=-0.245 $X2=4.41 $Y2=0.805
cc_81 VNB N_VGND_c_1375_n 0.0181447f $X=-0.19 $Y=-0.245 $X2=4.41 $Y2=0.805
cc_82 VNB N_VGND_c_1376_n 0.0173087f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.51
cc_83 VNB N_VGND_c_1377_n 0.0474958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1378_n 0.0350474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1379_n 0.454191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1380_n 0.0053824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1381_n 0.00938842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1382_n 0.0127902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_309_131#_c_1473_n 0.0195634f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.345
cc_90 VNB N_A_309_131#_c_1474_n 0.00505032f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.495
cc_91 VNB N_A_309_131#_c_1475_n 0.00647189f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=2.465
cc_92 VNB N_A_940_119#_c_1501_n 0.012382f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.495
cc_93 VNB N_A_940_119#_c_1502_n 0.00369837f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=2.465
cc_94 VPB N_A_84_21#_M1020_g 0.0215411f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_95 VPB N_A_84_21#_c_177_n 0.00608107f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.42
cc_96 VPB N_A_84_21#_M1030_g 0.0214105f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_97 VPB N_A_84_21#_c_182_n 0.00117245f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.785
cc_98 VPB N_A_84_21#_c_191_n 0.00737751f $X=-0.19 $Y=1.655 $X2=3.605 $Y2=1.87
cc_99 VPB N_A_84_21#_c_192_n 0.00237367f $X=-0.19 $Y=1.655 $X2=3.04 $Y2=1.87
cc_100 VPB N_A_84_21#_c_193_n 0.00157353f $X=-0.19 $Y=1.655 $X2=4.245 $Y2=2.16
cc_101 VPB N_A_84_21#_c_194_n 0.00349326f $X=-0.19 $Y=1.655 $X2=3.69 $Y2=1.87
cc_102 VPB N_A_84_21#_c_195_n 0.00424488f $X=-0.19 $Y=1.655 $X2=4.41 $Y2=2.24
cc_103 VPB N_A_M1012_g 0.0303359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_M1010_g 0.0272525f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.42
cc_105 VPB N_A_M1021_g 0.0281043f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_106 VPB N_A_M1025_g 0.0222135f $X=-0.19 $Y=1.655 $X2=2.87 $Y2=1.315
cc_107 VPB N_A_c_332_n 0.00166748f $X=-0.19 $Y=1.655 $X2=4.41 $Y2=0.805
cc_108 VPB N_A_c_343_n 0.0096922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_c_344_n 5.64283e-19 $X=-0.19 $Y=1.655 $X2=4.245 $Y2=2.16
cc_110 VPB N_A_c_345_n 0.00307567f $X=-0.19 $Y=1.655 $X2=3.775 $Y2=2.16
cc_111 VPB N_A_c_346_n 0.00492652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_c_334_n 0.0242241f $X=-0.19 $Y=1.655 $X2=3.63 $Y2=1.17
cc_113 VPB N_A_c_348_n 0.00599105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_c_349_n 0.00212794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_c_335_n 0.00750534f $X=-0.19 $Y=1.655 $X2=1.017 $Y2=1.675
cc_116 VPB N_A_c_336_n 0.00642647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_c_337_n 0.00358702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_395_398#_M1031_g 0.0186213f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_119 VPB N_A_395_398#_M1003_g 0.0220162f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=1.51
cc_120 VPB N_A_395_398#_M1028_g 0.0234832f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=1.17
cc_121 VPB N_A_395_398#_c_542_n 0.001734f $X=-0.19 $Y=1.655 $X2=3.715 $Y2=0.805
cc_122 VPB N_A_395_398#_c_558_n 0.00576199f $X=-0.19 $Y=1.655 $X2=3.69 $Y2=1.87
cc_123 VPB N_A_395_398#_c_559_n 0.0111283f $X=-0.19 $Y=1.655 $X2=3.69 $Y2=2.16
cc_124 VPB N_A_395_398#_c_560_n 0.0172351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_395_398#_c_561_n 0.00656256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_395_398#_c_562_n 0.00213323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_395_398#_c_563_n 0.0091049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_395_398#_c_551_n 0.0308111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_395_398#_c_565_n 0.0040097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_395_398#_c_553_n 0.0397783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_CIN_M1011_g 0.0183817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_CIN_c_814_n 0.0775359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_CIN_c_815_n 0.120305f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.495
cc_134 VPB N_CIN_c_816_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_135 VPB N_CIN_M1019_g 0.0471661f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.42
cc_136 VPB N_CIN_c_818_n 0.0787005f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_137 VPB N_CIN_M1005_g 0.0422613f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=1.51
cc_138 VPB N_CIN_c_820_n 0.00749069f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=1.51
cc_139 VPB CIN 0.00174635f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.785
cc_140 VPB N_CIN_c_812_n 0.0237896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_B_M1023_g 0.0300601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_B_M1029_g 0.0275904f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.495
cc_143 VPB N_B_c_921_n 0.00549294f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.345
cc_144 VPB N_B_M1000_g 0.0390096f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_145 VPB N_B_M1014_g 0.024859f $X=-0.19 $Y=1.655 $X2=2.87 $Y2=1.315
cc_146 VPB N_B_c_929_n 8.80119e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_1084_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_148 VPB N_VPWR_c_1085_n 0.0197167f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.675
cc_149 VPB N_VPWR_c_1086_n 0.0109785f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.42
cc_150 VPB N_VPWR_c_1087_n 0.00768785f $X=-0.19 $Y=1.655 $X2=2.87 $Y2=1.315
cc_151 VPB N_VPWR_c_1088_n 0.00581176f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=1.17
cc_152 VPB N_VPWR_c_1089_n 0.0195032f $X=-0.19 $Y=1.655 $X2=4.245 $Y2=2.16
cc_153 VPB N_VPWR_c_1090_n 0.0147344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_1091_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.575 $Y2=1.315
cc_155 VPB N_VPWR_c_1092_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_1093_n 0.0433074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_1094_n 0.0558436f $X=-0.19 $Y=1.655 $X2=3.69 $Y2=2.16
cc_158 VPB N_VPWR_c_1095_n 0.0162889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_1096_n 0.0443074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1083_n 0.0927393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1098_n 0.00597398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1099_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1100_n 0.00519718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1101_n 0.017051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB SUM 0.00837207f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_166 VPB SUM 0.0278035f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.785
cc_167 VPB N_A_309_398#_c_1262_n 0.00124188f $X=-0.19 $Y=1.655 $X2=0.495
+ $Y2=0.655
cc_168 VPB N_A_309_398#_c_1263_n 0.0187623f $X=-0.19 $Y=1.655 $X2=0.495
+ $Y2=1.495
cc_169 VPB N_A_309_398#_c_1264_n 0.00463264f $X=-0.19 $Y=1.655 $X2=0.495
+ $Y2=2.465
cc_170 VPB N_A_309_398#_c_1265_n 0.00664198f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.42
cc_171 VPB N_A_941_419#_c_1297_n 0.00187308f $X=-0.19 $Y=1.655 $X2=0.495
+ $Y2=1.495
cc_172 VPB N_A_941_419#_c_1298_n 0.00237027f $X=-0.19 $Y=1.655 $X2=0.495
+ $Y2=2.465
cc_173 VPB N_A_941_419#_c_1299_n 0.0043335f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.42
cc_174 VPB COUT 0.00471054f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_175 N_A_84_21#_c_182_n N_A_M1012_g 0.00331308f $X=2.955 $Y=1.785 $X2=0 $Y2=0
cc_176 N_A_84_21#_c_192_n N_A_M1012_g 0.00826977f $X=3.04 $Y=1.87 $X2=0 $Y2=0
cc_177 N_A_84_21#_c_181_n N_A_M1001_g 8.24058e-19 $X=2.87 $Y=1.315 $X2=0 $Y2=0
cc_178 N_A_84_21#_c_183_n N_A_M1001_g 0.00919437f $X=3.545 $Y=1.17 $X2=0 $Y2=0
cc_179 N_A_84_21#_c_184_n N_A_M1001_g 8.94209e-19 $X=3.715 $Y=0.805 $X2=0 $Y2=0
cc_180 N_A_84_21#_c_186_n N_A_M1001_g 0.0105421f $X=2.955 $Y=1.17 $X2=0 $Y2=0
cc_181 N_A_84_21#_c_183_n N_A_M1002_g 0.0130092f $X=3.545 $Y=1.17 $X2=0 $Y2=0
cc_182 N_A_84_21#_c_184_n N_A_M1002_g 0.00933558f $X=3.715 $Y=0.805 $X2=0 $Y2=0
cc_183 N_A_84_21#_c_186_n N_A_M1002_g 6.20981e-19 $X=2.955 $Y=1.17 $X2=0 $Y2=0
cc_184 N_A_84_21#_c_182_n N_A_M1010_g 5.86732e-19 $X=2.955 $Y=1.785 $X2=0 $Y2=0
cc_185 N_A_84_21#_c_191_n N_A_M1010_g 0.00937122f $X=3.605 $Y=1.87 $X2=0 $Y2=0
cc_186 N_A_84_21#_c_194_n N_A_M1010_g 0.00360429f $X=3.69 $Y=1.87 $X2=0 $Y2=0
cc_187 N_A_84_21#_c_182_n N_A_c_330_n 0.0129482f $X=2.955 $Y=1.785 $X2=0 $Y2=0
cc_188 N_A_84_21#_c_183_n N_A_c_330_n 0.021815f $X=3.545 $Y=1.17 $X2=0 $Y2=0
cc_189 N_A_84_21#_c_191_n N_A_c_330_n 0.0257233f $X=3.605 $Y=1.87 $X2=0 $Y2=0
cc_190 N_A_84_21#_c_184_n N_A_c_330_n 0.0135328f $X=3.715 $Y=0.805 $X2=0 $Y2=0
cc_191 N_A_84_21#_c_212_p N_A_c_330_n 0.0171935f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_192 N_A_84_21#_c_193_n N_A_c_330_n 0.00931724f $X=4.245 $Y=2.16 $X2=0 $Y2=0
cc_193 N_A_84_21#_c_194_n N_A_c_330_n 0.012944f $X=3.69 $Y=1.87 $X2=0 $Y2=0
cc_194 N_A_84_21#_c_195_n N_A_c_330_n 0.00173318f $X=4.41 $Y=2.24 $X2=0 $Y2=0
cc_195 N_A_84_21#_c_212_p N_A_c_333_n 0.00783928f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_196 N_A_84_21#_c_195_n N_A_c_333_n 0.00409129f $X=4.41 $Y=2.24 $X2=0 $Y2=0
cc_197 N_A_84_21#_c_181_n N_A_c_335_n 2.98617e-19 $X=2.87 $Y=1.315 $X2=0 $Y2=0
cc_198 N_A_84_21#_c_182_n N_A_c_335_n 0.0130849f $X=2.955 $Y=1.785 $X2=0 $Y2=0
cc_199 N_A_84_21#_c_183_n N_A_c_335_n 0.00249007f $X=3.545 $Y=1.17 $X2=0 $Y2=0
cc_200 N_A_84_21#_c_191_n N_A_c_335_n 0.00510554f $X=3.605 $Y=1.87 $X2=0 $Y2=0
cc_201 N_A_84_21#_c_186_n N_A_c_335_n 0.00454622f $X=2.955 $Y=1.17 $X2=0 $Y2=0
cc_202 N_A_84_21#_M1007_g N_A_395_398#_c_542_n 0.00195325f $X=0.495 $Y=0.655
+ $X2=0 $Y2=0
cc_203 N_A_84_21#_M1020_g N_A_395_398#_c_542_n 0.00843086f $X=0.495 $Y=2.465
+ $X2=0 $Y2=0
cc_204 N_A_84_21#_c_177_n N_A_395_398#_c_542_n 0.014497f $X=0.85 $Y=1.42 $X2=0
+ $Y2=0
cc_205 N_A_84_21#_M1008_g N_A_395_398#_c_542_n 0.00208272f $X=0.925 $Y=0.655
+ $X2=0 $Y2=0
cc_206 N_A_84_21#_c_179_n N_A_395_398#_c_542_n 0.00201611f $X=0.495 $Y=1.42
+ $X2=0 $Y2=0
cc_207 N_A_84_21#_c_180_n N_A_395_398#_c_542_n 0.0131478f $X=1.49 $Y=1.51 $X2=0
+ $Y2=0
cc_208 N_A_84_21#_c_177_n N_A_395_398#_c_543_n 0.00331717f $X=0.85 $Y=1.42 $X2=0
+ $Y2=0
cc_209 N_A_84_21#_M1008_g N_A_395_398#_c_543_n 0.0136273f $X=0.925 $Y=0.655
+ $X2=0 $Y2=0
cc_210 N_A_84_21#_c_180_n N_A_395_398#_c_543_n 0.0131559f $X=1.49 $Y=1.51 $X2=0
+ $Y2=0
cc_211 N_A_84_21#_M1007_g N_A_395_398#_c_576_n 0.00517822f $X=0.495 $Y=0.655
+ $X2=0 $Y2=0
cc_212 N_A_84_21#_c_180_n N_A_395_398#_c_577_n 0.00940804f $X=1.49 $Y=1.51 $X2=0
+ $Y2=0
cc_213 N_A_84_21#_c_181_n N_A_395_398#_c_577_n 0.0316581f $X=2.87 $Y=1.315 $X2=0
+ $Y2=0
cc_214 N_A_84_21#_c_185_n N_A_395_398#_c_577_n 0.010375f $X=1.575 $Y=1.315 $X2=0
+ $Y2=0
cc_215 N_A_84_21#_M1020_g N_A_395_398#_c_580_n 0.0067755f $X=0.495 $Y=2.465
+ $X2=0 $Y2=0
cc_216 N_A_84_21#_c_177_n N_A_395_398#_c_548_n 0.00322764f $X=0.85 $Y=1.42 $X2=0
+ $Y2=0
cc_217 N_A_84_21#_M1008_g N_A_395_398#_c_548_n 4.4635e-19 $X=0.925 $Y=0.655
+ $X2=0 $Y2=0
cc_218 N_A_84_21#_c_180_n N_A_395_398#_c_548_n 0.0124611f $X=1.49 $Y=1.51 $X2=0
+ $Y2=0
cc_219 N_A_84_21#_c_185_n N_A_395_398#_c_548_n 7.70754e-19 $X=1.575 $Y=1.315
+ $X2=0 $Y2=0
cc_220 N_A_84_21#_c_177_n N_A_395_398#_c_558_n 0.00512044f $X=0.85 $Y=1.42 $X2=0
+ $Y2=0
cc_221 N_A_84_21#_M1030_g N_A_395_398#_c_558_n 0.0180791f $X=0.925 $Y=2.465
+ $X2=0 $Y2=0
cc_222 N_A_84_21#_c_180_n N_A_395_398#_c_558_n 0.022529f $X=1.49 $Y=1.51 $X2=0
+ $Y2=0
cc_223 N_A_84_21#_c_181_n N_A_395_398#_c_558_n 0.00488163f $X=2.87 $Y=1.315
+ $X2=0 $Y2=0
cc_224 N_A_84_21#_c_185_n N_A_395_398#_c_558_n 0.00698117f $X=1.575 $Y=1.315
+ $X2=0 $Y2=0
cc_225 N_A_84_21#_c_192_n N_A_395_398#_c_559_n 0.00135985f $X=3.04 $Y=1.87 $X2=0
+ $Y2=0
cc_226 N_A_84_21#_c_181_n N_A_395_398#_c_549_n 0.022295f $X=2.87 $Y=1.315 $X2=0
+ $Y2=0
cc_227 N_A_84_21#_M1017_d N_A_395_398#_c_560_n 0.00182568f $X=4.27 $Y=2.095
+ $X2=0 $Y2=0
cc_228 N_A_84_21#_c_180_n N_A_395_398#_c_560_n 0.00380091f $X=1.49 $Y=1.51 $X2=0
+ $Y2=0
cc_229 N_A_84_21#_c_181_n N_A_395_398#_c_560_n 0.0114629f $X=2.87 $Y=1.315 $X2=0
+ $Y2=0
cc_230 N_A_84_21#_c_191_n N_A_395_398#_c_560_n 0.0216877f $X=3.605 $Y=1.87 $X2=0
+ $Y2=0
cc_231 N_A_84_21#_c_192_n N_A_395_398#_c_560_n 0.00811848f $X=3.04 $Y=1.87 $X2=0
+ $Y2=0
cc_232 N_A_84_21#_c_193_n N_A_395_398#_c_560_n 0.0278652f $X=4.245 $Y=2.16 $X2=0
+ $Y2=0
cc_233 N_A_84_21#_c_185_n N_A_395_398#_c_560_n 0.00116063f $X=1.575 $Y=1.315
+ $X2=0 $Y2=0
cc_234 N_A_84_21#_c_194_n N_A_395_398#_c_560_n 0.0201589f $X=3.69 $Y=1.87 $X2=0
+ $Y2=0
cc_235 N_A_84_21#_c_195_n N_A_395_398#_c_560_n 0.0181448f $X=4.41 $Y=2.24 $X2=0
+ $Y2=0
cc_236 N_A_84_21#_c_177_n N_A_395_398#_c_601_n 0.00148918f $X=0.85 $Y=1.42 $X2=0
+ $Y2=0
cc_237 N_A_84_21#_M1030_g N_A_395_398#_c_601_n 9.73171e-19 $X=0.925 $Y=2.465
+ $X2=0 $Y2=0
cc_238 N_A_84_21#_c_180_n N_A_395_398#_c_601_n 2.06085e-19 $X=1.49 $Y=1.51 $X2=0
+ $Y2=0
cc_239 N_A_84_21#_c_195_n N_A_395_398#_c_562_n 0.00143583f $X=4.41 $Y=2.24 $X2=0
+ $Y2=0
cc_240 N_A_84_21#_c_195_n N_A_395_398#_c_565_n 0.00248883f $X=4.41 $Y=2.24 $X2=0
+ $Y2=0
cc_241 N_A_84_21#_c_181_n N_CIN_M1018_g 0.0129118f $X=2.87 $Y=1.315 $X2=0 $Y2=0
cc_242 N_A_84_21#_c_185_n N_CIN_M1018_g 0.00194358f $X=1.575 $Y=1.315 $X2=0
+ $Y2=0
cc_243 N_A_84_21#_c_212_p N_CIN_M1019_g 0.0135558f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_244 N_A_84_21#_c_193_n N_CIN_M1019_g 0.0110449f $X=4.245 $Y=2.16 $X2=0 $Y2=0
cc_245 N_A_84_21#_c_194_n N_CIN_M1019_g 0.00183749f $X=3.69 $Y=1.87 $X2=0 $Y2=0
cc_246 N_A_84_21#_c_195_n N_CIN_M1019_g 0.00998383f $X=4.41 $Y=2.24 $X2=0 $Y2=0
cc_247 N_A_84_21#_c_195_n N_CIN_c_818_n 0.00288899f $X=4.41 $Y=2.24 $X2=0 $Y2=0
cc_248 N_A_84_21#_c_181_n CIN 0.0513884f $X=2.87 $Y=1.315 $X2=0 $Y2=0
cc_249 N_A_84_21#_c_182_n CIN 0.0101157f $X=2.955 $Y=1.785 $X2=0 $Y2=0
cc_250 N_A_84_21#_c_185_n CIN 0.00191797f $X=1.575 $Y=1.315 $X2=0 $Y2=0
cc_251 N_A_84_21#_c_181_n N_CIN_c_812_n 0.0142907f $X=2.87 $Y=1.315 $X2=0 $Y2=0
cc_252 N_A_84_21#_c_182_n N_CIN_c_812_n 0.00248146f $X=2.955 $Y=1.785 $X2=0
+ $Y2=0
cc_253 N_A_84_21#_c_192_n N_CIN_c_812_n 0.00339859f $X=3.04 $Y=1.87 $X2=0 $Y2=0
cc_254 N_A_84_21#_c_185_n N_CIN_c_812_n 0.00173991f $X=1.575 $Y=1.315 $X2=0
+ $Y2=0
cc_255 N_A_84_21#_c_177_n N_B_M1023_g 0.0219211f $X=0.85 $Y=1.42 $X2=0 $Y2=0
cc_256 N_A_84_21#_M1030_g N_B_M1023_g 0.0267369f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A_84_21#_c_180_n N_B_M1023_g 0.00732362f $X=1.49 $Y=1.51 $X2=0 $Y2=0
cc_258 N_A_84_21#_c_181_n N_B_M1023_g 3.4364e-19 $X=2.87 $Y=1.315 $X2=0 $Y2=0
cc_259 N_A_84_21#_c_185_n N_B_M1023_g 0.0103892f $X=1.575 $Y=1.315 $X2=0 $Y2=0
cc_260 N_A_84_21#_c_184_n N_B_c_917_n 0.00197128f $X=3.715 $Y=0.805 $X2=0 $Y2=0
cc_261 N_A_84_21#_M1008_g N_B_c_918_n 0.0278772f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A_84_21#_c_184_n N_B_M1029_g 0.00569994f $X=3.715 $Y=0.805 $X2=0 $Y2=0
cc_263 N_A_84_21#_c_212_p N_B_M1029_g 0.0155727f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_264 N_A_84_21#_c_193_n N_B_M1029_g 0.0120753f $X=4.245 $Y=2.16 $X2=0 $Y2=0
cc_265 N_A_84_21#_c_194_n N_B_M1029_g 0.0092359f $X=3.69 $Y=1.87 $X2=0 $Y2=0
cc_266 N_A_84_21#_c_195_n N_B_M1029_g 0.00251411f $X=4.41 $Y=2.24 $X2=0 $Y2=0
cc_267 N_A_84_21#_c_212_p N_B_c_920_n 0.00668326f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_268 N_A_84_21#_M1020_g N_VPWR_c_1085_n 0.0111146f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_269 N_A_84_21#_M1030_g N_VPWR_c_1085_n 5.67328e-19 $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_84_21#_M1020_g N_VPWR_c_1086_n 6.18119e-19 $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_84_21#_M1030_g N_VPWR_c_1086_n 0.0149036f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_A_84_21#_c_191_n N_VPWR_c_1087_n 0.0165714f $X=3.605 $Y=1.87 $X2=0
+ $Y2=0
cc_273 N_A_84_21#_M1020_g N_VPWR_c_1092_n 0.00486043f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_274 N_A_84_21#_M1030_g N_VPWR_c_1092_n 0.00486043f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_275 N_A_84_21#_c_195_n N_VPWR_c_1094_n 0.00574841f $X=4.41 $Y=2.24 $X2=0
+ $Y2=0
cc_276 N_A_84_21#_M1020_g N_VPWR_c_1083_n 0.00454119f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_A_84_21#_M1030_g N_VPWR_c_1083_n 0.00824727f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_A_84_21#_c_195_n N_VPWR_c_1083_n 0.00704652f $X=4.41 $Y=2.24 $X2=0
+ $Y2=0
cc_279 N_A_84_21#_M1007_g N_SUM_c_1216_n 0.0139502f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_280 N_A_84_21#_c_177_n N_SUM_c_1216_n 2.54341e-19 $X=0.85 $Y=1.42 $X2=0 $Y2=0
cc_281 N_A_84_21#_M1008_g N_SUM_c_1216_n 0.00388351f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_282 N_A_84_21#_M1020_g N_SUM_c_1219_n 0.0137789f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_84_21#_M1007_g N_SUM_c_1220_n 0.0109581f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_284 N_A_84_21#_M1008_g N_SUM_c_1220_n 0.00539566f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_285 N_A_84_21#_M1007_g SUM 0.0374699f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_286 N_A_84_21#_c_192_n N_A_309_398#_c_1265_n 0.00195553f $X=3.04 $Y=1.87
+ $X2=0 $Y2=0
cc_287 N_A_84_21#_c_194_n A_710_419# 0.00413256f $X=3.69 $Y=1.87 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_84_21#_c_193_n A_782_419# 0.00366293f $X=4.245 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_84_21#_c_195_n N_A_941_419#_c_1299_n 0.00768023f $X=4.41 $Y=2.24
+ $X2=0 $Y2=0
cc_290 N_A_84_21#_M1007_g N_VGND_c_1367_n 0.00327088f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_291 N_A_84_21#_M1008_g N_VGND_c_1368_n 0.00240658f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_292 N_A_84_21#_c_183_n N_VGND_c_1369_n 0.0153144f $X=3.545 $Y=1.17 $X2=0
+ $Y2=0
cc_293 N_A_84_21#_M1007_g N_VGND_c_1376_n 0.00426006f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_294 N_A_84_21#_M1008_g N_VGND_c_1376_n 0.0054895f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_295 N_A_84_21#_c_184_n N_VGND_c_1377_n 0.0025454f $X=3.715 $Y=0.805 $X2=0
+ $Y2=0
cc_296 N_A_84_21#_c_212_p N_VGND_c_1377_n 0.0122663f $X=4.41 $Y=0.805 $X2=0
+ $Y2=0
cc_297 N_A_84_21#_M1007_g N_VGND_c_1379_n 0.00675648f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_298 N_A_84_21#_M1008_g N_VGND_c_1379_n 0.0101718f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_299 N_A_84_21#_c_184_n N_VGND_c_1379_n 0.00439046f $X=3.715 $Y=0.805 $X2=0
+ $Y2=0
cc_300 N_A_84_21#_c_212_p N_VGND_c_1379_n 0.0203621f $X=4.41 $Y=0.805 $X2=0
+ $Y2=0
cc_301 N_A_84_21#_c_181_n N_A_309_131#_c_1474_n 0.010712f $X=2.87 $Y=1.315 $X2=0
+ $Y2=0
cc_302 N_A_84_21#_c_186_n N_A_309_131#_c_1474_n 0.00842735f $X=2.955 $Y=1.17
+ $X2=0 $Y2=0
cc_303 N_A_84_21#_c_184_n A_710_119# 0.00151919f $X=3.715 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_304 N_A_84_21#_c_212_p A_782_119# 0.00319459f $X=4.41 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_305 N_A_c_331_n N_A_395_398#_M1022_g 0.0161821f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_306 N_A_c_332_n N_A_395_398#_M1022_g 4.56102e-19 $X=5.39 $Y=1.845 $X2=0 $Y2=0
cc_307 N_A_c_333_n N_A_395_398#_M1022_g 0.00298981f $X=4.41 $Y=1.42 $X2=0 $Y2=0
cc_308 N_A_M1026_g N_A_395_398#_c_537_n 0.0162793f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_309 N_A_M1021_g N_A_395_398#_M1003_g 0.00674694f $X=6.19 $Y=2.54 $X2=0 $Y2=0
cc_310 N_A_M1026_g N_A_395_398#_M1003_g 0.00393116f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_311 N_A_c_345_n N_A_395_398#_M1003_g 0.00506379f $X=6.765 $Y=2.015 $X2=0
+ $Y2=0
cc_312 N_A_c_387_p N_A_395_398#_M1003_g 0.0064631f $X=6.85 $Y=2.325 $X2=0 $Y2=0
cc_313 N_A_c_346_n N_A_395_398#_M1003_g 0.00994449f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_314 N_A_c_389_p N_A_395_398#_M1003_g 0.00300833f $X=6.935 $Y=2.41 $X2=0 $Y2=0
cc_315 N_A_c_334_n N_A_395_398#_M1003_g 0.00712159f $X=6.28 $Y=1.77 $X2=0 $Y2=0
cc_316 N_A_c_348_n N_A_395_398#_M1003_g 7.84818e-19 $X=6.28 $Y=1.93 $X2=0 $Y2=0
cc_317 N_A_M1009_g N_A_395_398#_c_539_n 0.0109455f $X=8.19 $Y=0.895 $X2=0 $Y2=0
cc_318 N_A_M1025_g N_A_395_398#_M1028_g 0.0126001f $X=8.19 $Y=2.155 $X2=0 $Y2=0
cc_319 N_A_c_387_p N_A_395_398#_M1028_g 8.33057e-19 $X=6.85 $Y=2.325 $X2=0 $Y2=0
cc_320 N_A_c_346_n N_A_395_398#_M1028_g 0.0132779f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_321 N_A_c_349_n N_A_395_398#_M1028_g 0.00693451f $X=7.91 $Y=2.325 $X2=0 $Y2=0
cc_322 N_A_c_336_n N_A_395_398#_M1028_g 0.00282104f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_323 N_A_c_337_n N_A_395_398#_M1028_g 0.00197837f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_324 N_A_c_345_n N_A_395_398#_c_541_n 6.13969e-19 $X=6.765 $Y=2.015 $X2=0
+ $Y2=0
cc_325 N_A_M1009_g N_A_395_398#_c_544_n 4.99325e-19 $X=8.19 $Y=0.895 $X2=0 $Y2=0
cc_326 N_A_c_336_n N_A_395_398#_c_544_n 5.37243e-19 $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_327 N_A_c_337_n N_A_395_398#_c_544_n 0.0100838f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_328 N_A_M1009_g N_A_395_398#_c_545_n 0.00458665f $X=8.19 $Y=0.895 $X2=0 $Y2=0
cc_329 N_A_c_336_n N_A_395_398#_c_545_n 0.0132256f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_330 N_A_c_337_n N_A_395_398#_c_545_n 9.19045e-19 $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_331 N_A_M1009_g N_A_395_398#_c_546_n 0.0123831f $X=8.19 $Y=0.895 $X2=0 $Y2=0
cc_332 N_A_c_336_n N_A_395_398#_c_546_n 0.00438376f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_333 N_A_c_337_n N_A_395_398#_c_546_n 0.033793f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_334 N_A_M1001_g N_A_395_398#_c_549_n 0.00253981f $X=3.045 $Y=0.805 $X2=0
+ $Y2=0
cc_335 N_A_M1012_g N_A_395_398#_c_560_n 0.00967645f $X=2.965 $Y=2.415 $X2=0
+ $Y2=0
cc_336 N_A_M1010_g N_A_395_398#_c_560_n 0.00892077f $X=3.475 $Y=2.415 $X2=0
+ $Y2=0
cc_337 N_A_c_330_n N_A_395_398#_c_560_n 0.0134742f $X=4.325 $Y=1.525 $X2=0 $Y2=0
cc_338 N_A_c_331_n N_A_395_398#_c_560_n 0.0061373f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_339 N_A_c_333_n N_A_395_398#_c_560_n 0.0040975f $X=4.41 $Y=1.42 $X2=0 $Y2=0
cc_340 N_A_M1021_g N_A_395_398#_c_561_n 0.00697542f $X=6.19 $Y=2.54 $X2=0 $Y2=0
cc_341 N_A_M1025_g N_A_395_398#_c_561_n 0.0101902f $X=8.19 $Y=2.155 $X2=0 $Y2=0
cc_342 N_A_c_331_n N_A_395_398#_c_561_n 0.00346562f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_343 N_A_c_343_n N_A_395_398#_c_561_n 0.0207852f $X=6.115 $Y=1.93 $X2=0 $Y2=0
cc_344 N_A_c_344_n N_A_395_398#_c_561_n 0.0117657f $X=5.475 $Y=1.93 $X2=0 $Y2=0
cc_345 N_A_c_345_n N_A_395_398#_c_561_n 0.0215904f $X=6.765 $Y=2.015 $X2=0 $Y2=0
cc_346 N_A_c_387_p N_A_395_398#_c_561_n 0.00322544f $X=6.85 $Y=2.325 $X2=0 $Y2=0
cc_347 N_A_c_346_n N_A_395_398#_c_561_n 0.0266853f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_348 N_A_c_348_n N_A_395_398#_c_561_n 0.0141718f $X=6.28 $Y=1.93 $X2=0 $Y2=0
cc_349 N_A_c_349_n N_A_395_398#_c_561_n 0.0207327f $X=7.91 $Y=2.325 $X2=0 $Y2=0
cc_350 N_A_c_337_n N_A_395_398#_c_561_n 0.0118131f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_351 N_A_c_331_n N_A_395_398#_c_562_n 0.00330344f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_352 N_A_c_344_n N_A_395_398#_c_562_n 0.00139236f $X=5.475 $Y=1.93 $X2=0 $Y2=0
cc_353 N_A_c_331_n N_A_395_398#_c_551_n 0.00699956f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_354 N_A_c_332_n N_A_395_398#_c_551_n 5.69846e-19 $X=5.39 $Y=1.845 $X2=0 $Y2=0
cc_355 N_A_c_331_n N_A_395_398#_c_565_n 0.0335688f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_356 N_A_c_332_n N_A_395_398#_c_565_n 0.0125905f $X=5.39 $Y=1.845 $X2=0 $Y2=0
cc_357 N_A_c_344_n N_A_395_398#_c_565_n 0.0124072f $X=5.475 $Y=1.93 $X2=0 $Y2=0
cc_358 N_A_c_346_n N_A_395_398#_c_553_n 0.00299164f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_359 N_A_c_349_n N_A_395_398#_c_553_n 0.00835838f $X=7.91 $Y=2.325 $X2=0 $Y2=0
cc_360 N_A_c_337_n N_A_395_398#_c_553_n 0.0138707f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_361 N_A_c_335_n N_CIN_M1018_g 0.00192431f $X=3.475 $Y=1.52 $X2=0 $Y2=0
cc_362 N_A_M1012_g N_CIN_c_814_n 0.0135816f $X=2.965 $Y=2.415 $X2=0 $Y2=0
cc_363 N_A_M1012_g N_CIN_c_815_n 0.0101508f $X=2.965 $Y=2.415 $X2=0 $Y2=0
cc_364 N_A_M1010_g N_CIN_c_815_n 0.0103107f $X=3.475 $Y=2.415 $X2=0 $Y2=0
cc_365 N_A_c_330_n N_CIN_M1019_g 0.0119375f $X=4.325 $Y=1.525 $X2=0 $Y2=0
cc_366 N_A_c_333_n N_CIN_M1019_g 0.00276305f $X=4.41 $Y=1.42 $X2=0 $Y2=0
cc_367 N_A_c_331_n N_CIN_M1005_g 0.00534782f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_368 N_A_c_332_n N_CIN_M1005_g 0.00777661f $X=5.39 $Y=1.845 $X2=0 $Y2=0
cc_369 N_A_c_344_n N_CIN_M1005_g 0.0049046f $X=5.475 $Y=1.93 $X2=0 $Y2=0
cc_370 N_A_c_331_n N_CIN_c_810_n 0.00928826f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_371 N_A_c_335_n CIN 8.24094e-19 $X=3.475 $Y=1.52 $X2=0 $Y2=0
cc_372 N_A_c_335_n N_CIN_c_812_n 0.0135816f $X=3.475 $Y=1.52 $X2=0 $Y2=0
cc_373 N_A_M1001_g N_B_c_917_n 0.0101549f $X=3.045 $Y=0.805 $X2=0 $Y2=0
cc_374 N_A_M1002_g N_B_c_917_n 0.0104164f $X=3.475 $Y=0.805 $X2=0 $Y2=0
cc_375 N_A_M1002_g N_B_M1029_g 0.1507f $X=3.475 $Y=0.805 $X2=0 $Y2=0
cc_376 N_A_c_330_n N_B_M1029_g 0.0125375f $X=4.325 $Y=1.525 $X2=0 $Y2=0
cc_377 N_A_M1026_g N_B_c_921_n 0.0135831f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_378 N_A_c_331_n N_B_c_921_n 0.00120117f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_379 N_A_c_332_n N_B_c_921_n 9.69406e-19 $X=5.39 $Y=1.845 $X2=0 $Y2=0
cc_380 N_A_c_343_n N_B_c_921_n 0.00338421f $X=6.115 $Y=1.93 $X2=0 $Y2=0
cc_381 N_A_c_334_n N_B_c_921_n 0.0040574f $X=6.28 $Y=1.77 $X2=0 $Y2=0
cc_382 N_A_c_332_n N_B_M1000_g 0.00186823f $X=5.39 $Y=1.845 $X2=0 $Y2=0
cc_383 N_A_c_343_n N_B_M1000_g 0.0103119f $X=6.115 $Y=1.93 $X2=0 $Y2=0
cc_384 N_A_c_334_n N_B_M1000_g 0.0306019f $X=6.28 $Y=1.77 $X2=0 $Y2=0
cc_385 N_A_c_348_n N_B_M1000_g 6.83184e-19 $X=6.28 $Y=1.93 $X2=0 $Y2=0
cc_386 N_A_M1026_g N_B_M1024_g 0.0202763f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_387 N_A_c_336_n N_B_M1006_g 0.0424542f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_388 N_A_c_337_n N_B_M1014_g 0.00117654f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_389 N_A_M1025_g N_B_c_926_n 0.0424542f $X=8.19 $Y=2.155 $X2=0 $Y2=0
cc_390 N_A_M1026_g N_B_c_927_n 0.0157639f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_391 N_A_c_343_n N_B_c_927_n 0.00837813f $X=6.115 $Y=1.93 $X2=0 $Y2=0
cc_392 N_A_c_345_n N_B_c_927_n 0.00860592f $X=6.765 $Y=2.015 $X2=0 $Y2=0
cc_393 N_A_c_334_n N_B_c_927_n 0.00480643f $X=6.28 $Y=1.77 $X2=0 $Y2=0
cc_394 N_A_c_348_n N_B_c_927_n 0.0236827f $X=6.28 $Y=1.93 $X2=0 $Y2=0
cc_395 N_A_M1026_g N_B_c_928_n 0.0084959f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_396 N_A_M1026_g N_B_c_975_n 0.00507176f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_397 N_A_M1026_g N_B_c_929_n 7.27889e-19 $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_398 N_A_c_331_n N_B_c_929_n 0.0141053f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_399 N_A_c_332_n N_B_c_929_n 0.011771f $X=5.39 $Y=1.845 $X2=0 $Y2=0
cc_400 N_A_c_343_n N_B_c_929_n 0.0166816f $X=6.115 $Y=1.93 $X2=0 $Y2=0
cc_401 N_A_c_334_n N_B_c_929_n 4.29681e-19 $X=6.28 $Y=1.77 $X2=0 $Y2=0
cc_402 N_A_M1009_g N_B_c_931_n 0.0424542f $X=8.19 $Y=0.895 $X2=0 $Y2=0
cc_403 N_A_M1009_g N_B_c_932_n 0.0114351f $X=8.19 $Y=0.895 $X2=0 $Y2=0
cc_404 N_A_c_345_n N_VPWR_M1021_d 0.0103497f $X=6.765 $Y=2.015 $X2=0 $Y2=0
cc_405 N_A_c_387_p N_VPWR_M1021_d 0.0030818f $X=6.85 $Y=2.325 $X2=0 $Y2=0
cc_406 N_A_c_389_p N_VPWR_M1021_d 0.00272549f $X=6.935 $Y=2.41 $X2=0 $Y2=0
cc_407 N_A_c_348_n N_VPWR_M1021_d 3.28668e-19 $X=6.28 $Y=1.93 $X2=0 $Y2=0
cc_408 N_A_c_346_n N_VPWR_M1028_s 0.0109605f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_409 N_A_c_349_n N_VPWR_M1028_s 0.0179381f $X=7.91 $Y=2.325 $X2=0 $Y2=0
cc_410 N_A_M1012_g N_VPWR_c_1087_n 0.00420576f $X=2.965 $Y=2.415 $X2=0 $Y2=0
cc_411 N_A_M1010_g N_VPWR_c_1087_n 0.0138718f $X=3.475 $Y=2.415 $X2=0 $Y2=0
cc_412 N_A_M1021_g N_VPWR_c_1121_n 0.00436921f $X=6.19 $Y=2.54 $X2=0 $Y2=0
cc_413 N_A_c_345_n N_VPWR_c_1121_n 0.00877343f $X=6.765 $Y=2.015 $X2=0 $Y2=0
cc_414 N_A_c_387_p N_VPWR_c_1121_n 0.00376375f $X=6.85 $Y=2.325 $X2=0 $Y2=0
cc_415 N_A_c_389_p N_VPWR_c_1121_n 0.0130694f $X=6.935 $Y=2.41 $X2=0 $Y2=0
cc_416 N_A_c_334_n N_VPWR_c_1121_n 8.31313e-19 $X=6.28 $Y=1.77 $X2=0 $Y2=0
cc_417 N_A_c_348_n N_VPWR_c_1121_n 0.0118774f $X=6.28 $Y=1.93 $X2=0 $Y2=0
cc_418 N_A_c_346_n N_VPWR_c_1089_n 0.0208314f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_419 N_A_M1021_g N_VPWR_c_1095_n 0.00422593f $X=6.19 $Y=2.54 $X2=0 $Y2=0
cc_420 N_A_M1025_g N_VPWR_c_1096_n 0.00312414f $X=8.19 $Y=2.155 $X2=0 $Y2=0
cc_421 N_A_M1012_g N_VPWR_c_1083_n 7.82699e-19 $X=2.965 $Y=2.415 $X2=0 $Y2=0
cc_422 N_A_M1010_g N_VPWR_c_1083_n 7.88961e-19 $X=3.475 $Y=2.415 $X2=0 $Y2=0
cc_423 N_A_M1021_g N_VPWR_c_1083_n 0.00432128f $X=6.19 $Y=2.54 $X2=0 $Y2=0
cc_424 N_A_M1025_g N_VPWR_c_1083_n 0.00410284f $X=8.19 $Y=2.155 $X2=0 $Y2=0
cc_425 N_A_c_346_n N_VPWR_c_1083_n 0.0259067f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_426 N_A_c_389_p N_VPWR_c_1083_n 6.00243e-19 $X=6.935 $Y=2.41 $X2=0 $Y2=0
cc_427 N_A_M1021_g N_VPWR_c_1101_n 0.00732418f $X=6.19 $Y=2.54 $X2=0 $Y2=0
cc_428 N_A_c_345_n N_VPWR_c_1101_n 0.00363973f $X=6.765 $Y=2.015 $X2=0 $Y2=0
cc_429 N_A_c_389_p N_VPWR_c_1101_n 0.00927754f $X=6.935 $Y=2.41 $X2=0 $Y2=0
cc_430 N_A_M1012_g N_A_309_398#_c_1263_n 0.00129728f $X=2.965 $Y=2.415 $X2=0
+ $Y2=0
cc_431 N_A_M1012_g N_A_309_398#_c_1265_n 0.00847976f $X=2.965 $Y=2.415 $X2=0
+ $Y2=0
cc_432 N_A_M1010_g N_A_309_398#_c_1265_n 2.03017e-19 $X=3.475 $Y=2.415 $X2=0
+ $Y2=0
cc_433 N_A_c_343_n N_A_941_419#_c_1301_n 0.011389f $X=6.115 $Y=1.93 $X2=0 $Y2=0
cc_434 N_A_c_344_n N_A_941_419#_c_1301_n 0.00548895f $X=5.475 $Y=1.93 $X2=0
+ $Y2=0
cc_435 N_A_M1021_g N_A_941_419#_c_1297_n 5.03748e-19 $X=6.19 $Y=2.54 $X2=0 $Y2=0
cc_436 N_A_c_343_n N_A_941_419#_c_1297_n 0.0168007f $X=6.115 $Y=1.93 $X2=0 $Y2=0
cc_437 N_A_c_346_n N_COUT_M1003_d 0.00498542f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_438 N_A_M1026_g N_COUT_c_1333_n 9.67293e-19 $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_439 N_A_M1026_g COUT 0.00129388f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_440 N_A_c_345_n COUT 0.0113577f $X=6.765 $Y=2.015 $X2=0 $Y2=0
cc_441 N_A_c_387_p COUT 0.00150729f $X=6.85 $Y=2.325 $X2=0 $Y2=0
cc_442 N_A_c_346_n COUT 0.0137335f $X=7.815 $Y=2.41 $X2=0 $Y2=0
cc_443 N_A_c_334_n COUT 0.00177283f $X=6.28 $Y=1.77 $X2=0 $Y2=0
cc_444 N_A_c_348_n COUT 0.00658313f $X=6.28 $Y=1.93 $X2=0 $Y2=0
cc_445 N_A_c_349_n COUT 0.00785465f $X=7.91 $Y=2.325 $X2=0 $Y2=0
cc_446 N_A_c_337_n COUT 0.00814639f $X=8.1 $Y=1.51 $X2=0 $Y2=0
cc_447 N_A_M1001_g N_VGND_c_1369_n 9.41818e-19 $X=3.045 $Y=0.805 $X2=0 $Y2=0
cc_448 N_A_M1002_g N_VGND_c_1369_n 0.00333437f $X=3.475 $Y=0.805 $X2=0 $Y2=0
cc_449 N_A_M1026_g N_VGND_c_1370_n 0.00112647f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_450 N_A_M1026_g N_VGND_c_1371_n 0.00431487f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_451 N_A_M1009_g N_VGND_c_1378_n 6.37941e-19 $X=8.19 $Y=0.895 $X2=0 $Y2=0
cc_452 N_A_M1001_g N_VGND_c_1379_n 7.82699e-19 $X=3.045 $Y=0.805 $X2=0 $Y2=0
cc_453 N_A_M1002_g N_VGND_c_1379_n 9.39239e-19 $X=3.475 $Y=0.805 $X2=0 $Y2=0
cc_454 N_A_M1026_g N_VGND_c_1379_n 0.00477801f $X=6.29 $Y=0.805 $X2=0 $Y2=0
cc_455 N_A_M1001_g N_A_309_131#_c_1473_n 0.00268017f $X=3.045 $Y=0.805 $X2=0
+ $Y2=0
cc_456 N_A_M1001_g N_A_309_131#_c_1474_n 0.00550791f $X=3.045 $Y=0.805 $X2=0
+ $Y2=0
cc_457 N_A_c_335_n N_A_309_131#_c_1474_n 2.39079e-19 $X=3.475 $Y=1.52 $X2=0
+ $Y2=0
cc_458 N_A_M1026_g N_A_940_119#_c_1501_n 0.00178478f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_459 N_A_c_331_n N_A_940_119#_c_1501_n 0.0400839f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_460 N_A_c_331_n N_A_940_119#_c_1502_n 0.0190198f $X=5.305 $Y=1.42 $X2=0 $Y2=0
cc_461 N_A_395_398#_c_558_n N_CIN_M1011_g 0.012468f $X=2.02 $Y=2.035 $X2=0 $Y2=0
cc_462 N_A_395_398#_c_577_n N_CIN_M1018_g 0.00952021f $X=2.145 $Y=0.965 $X2=0
+ $Y2=0
cc_463 N_A_395_398#_c_549_n N_CIN_M1018_g 0.00514581f $X=2.31 $Y=0.875 $X2=0
+ $Y2=0
cc_464 N_A_395_398#_c_559_n N_CIN_c_814_n 0.010789f $X=2.115 $Y=2.135 $X2=0
+ $Y2=0
cc_465 N_A_395_398#_c_560_n N_CIN_c_814_n 0.0103394f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_466 N_A_395_398#_M1022_g N_CIN_M1019_g 0.0515262f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_467 N_A_395_398#_M1031_g N_CIN_M1019_g 0.0135701f $X=4.63 $Y=2.415 $X2=0
+ $Y2=0
cc_468 N_A_395_398#_c_560_n N_CIN_M1019_g 0.00298515f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_469 N_A_395_398#_c_565_n N_CIN_M1019_g 0.00231057f $X=4.84 $Y=1.77 $X2=0
+ $Y2=0
cc_470 N_A_395_398#_M1031_g N_CIN_c_818_n 0.0104164f $X=4.63 $Y=2.415 $X2=0
+ $Y2=0
cc_471 N_A_395_398#_M1022_g N_CIN_M1015_g 0.0236465f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_472 N_A_395_398#_M1022_g N_CIN_M1005_g 0.00333394f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_473 N_A_395_398#_M1031_g N_CIN_M1005_g 0.0169736f $X=4.63 $Y=2.415 $X2=0
+ $Y2=0
cc_474 N_A_395_398#_c_561_n N_CIN_M1005_g 0.00451377f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_475 N_A_395_398#_c_562_n N_CIN_M1005_g 0.00163808f $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_476 N_A_395_398#_c_551_n N_CIN_M1005_g 0.0198828f $X=4.84 $Y=1.77 $X2=0 $Y2=0
cc_477 N_A_395_398#_c_565_n N_CIN_M1005_g 0.00477826f $X=4.84 $Y=1.77 $X2=0
+ $Y2=0
cc_478 N_A_395_398#_c_551_n N_CIN_c_810_n 0.00130959f $X=4.84 $Y=1.77 $X2=0
+ $Y2=0
cc_479 N_A_395_398#_c_565_n N_CIN_c_810_n 6.57557e-19 $X=4.84 $Y=1.77 $X2=0
+ $Y2=0
cc_480 N_A_395_398#_c_558_n CIN 0.0122627f $X=2.02 $Y=2.035 $X2=0 $Y2=0
cc_481 N_A_395_398#_c_559_n CIN 0.0196416f $X=2.115 $Y=2.135 $X2=0 $Y2=0
cc_482 N_A_395_398#_c_560_n CIN 0.0142557f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_483 N_A_395_398#_c_559_n N_CIN_c_812_n 0.00507346f $X=2.115 $Y=2.135 $X2=0
+ $Y2=0
cc_484 N_A_395_398#_c_577_n N_B_M1023_g 0.016366f $X=2.145 $Y=0.965 $X2=0 $Y2=0
cc_485 N_A_395_398#_c_548_n N_B_M1023_g 0.00429712f $X=1.14 $Y=0.965 $X2=0 $Y2=0
cc_486 N_A_395_398#_c_558_n N_B_M1023_g 0.0181505f $X=2.02 $Y=2.035 $X2=0 $Y2=0
cc_487 N_A_395_398#_c_549_n N_B_M1023_g 8.33984e-19 $X=2.31 $Y=0.875 $X2=0 $Y2=0
cc_488 N_A_395_398#_c_577_n N_B_c_917_n 3.46599e-19 $X=2.145 $Y=0.965 $X2=0
+ $Y2=0
cc_489 N_A_395_398#_c_560_n N_B_M1029_g 0.00207426f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_490 N_A_395_398#_M1022_g N_B_c_920_n 0.0104164f $X=4.625 $Y=0.805 $X2=0 $Y2=0
cc_491 N_A_395_398#_c_561_n N_B_M1000_g 0.00255335f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_492 N_A_395_398#_c_546_n N_B_M1006_g 0.0084664f $X=8.68 $Y=1.16 $X2=0 $Y2=0
cc_493 N_A_395_398#_c_550_n N_B_M1006_g 0.00123567f $X=8.86 $Y=0.96 $X2=0 $Y2=0
cc_494 N_A_395_398#_c_561_n N_B_M1014_g 0.0130348f $X=8.735 $Y=2.035 $X2=0 $Y2=0
cc_495 N_A_395_398#_c_553_n N_B_M1014_g 0.0145952f $X=8.785 $Y=1.99 $X2=0 $Y2=0
cc_496 N_A_395_398#_c_546_n N_B_c_926_n 0.00933848f $X=8.68 $Y=1.16 $X2=0 $Y2=0
cc_497 N_A_395_398#_c_550_n N_B_c_926_n 0.00573763f $X=8.86 $Y=0.96 $X2=0 $Y2=0
cc_498 N_A_395_398#_c_561_n N_B_c_926_n 4.86074e-19 $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_499 N_A_395_398#_M1003_g N_B_c_927_n 5.92827e-19 $X=6.985 $Y=2.465 $X2=0
+ $Y2=0
cc_500 N_A_395_398#_c_541_n N_B_c_927_n 3.3355e-19 $X=6.95 $Y=1.29 $X2=0 $Y2=0
cc_501 N_A_395_398#_c_561_n N_B_c_927_n 0.00434472f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_502 N_A_395_398#_c_537_n N_B_c_928_n 0.00790707f $X=6.915 $Y=1.215 $X2=0
+ $Y2=0
cc_503 N_A_395_398#_c_561_n N_B_c_929_n 0.00145669f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_504 N_A_395_398#_M1006_d B 0.00331651f $X=8.625 $Y=0.685 $X2=0 $Y2=0
cc_505 N_A_395_398#_c_550_n B 0.0291748f $X=8.86 $Y=0.96 $X2=0 $Y2=0
cc_506 N_A_395_398#_c_550_n N_B_c_931_n 8.76264e-19 $X=8.86 $Y=0.96 $X2=0 $Y2=0
cc_507 N_A_395_398#_c_537_n N_B_c_932_n 0.0124573f $X=6.915 $Y=1.215 $X2=0 $Y2=0
cc_508 N_A_395_398#_c_539_n N_B_c_932_n 0.016695f $X=7.345 $Y=1.215 $X2=0 $Y2=0
cc_509 N_A_395_398#_c_545_n N_B_c_932_n 0.00118015f $X=7.56 $Y=1.38 $X2=0 $Y2=0
cc_510 N_A_395_398#_c_546_n N_B_c_932_n 0.0314202f $X=8.68 $Y=1.16 $X2=0 $Y2=0
cc_511 N_A_395_398#_c_547_n N_B_c_932_n 0.00732531f $X=7.645 $Y=1.16 $X2=0 $Y2=0
cc_512 N_A_395_398#_c_552_n N_B_c_932_n 3.39151e-19 $X=7.27 $Y=1.38 $X2=0 $Y2=0
cc_513 N_A_395_398#_c_558_n N_VPWR_M1030_s 0.00607417f $X=2.02 $Y=2.035 $X2=0
+ $Y2=0
cc_514 N_A_395_398#_c_560_n N_VPWR_M1012_d 0.0043064f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_515 N_A_395_398#_c_561_n N_VPWR_M1021_d 0.0039827f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_516 N_A_395_398#_c_561_n N_VPWR_M1028_s 0.0145575f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_517 N_A_395_398#_c_558_n N_VPWR_c_1086_n 0.0228478f $X=2.02 $Y=2.035 $X2=0
+ $Y2=0
cc_518 N_A_395_398#_c_560_n N_VPWR_c_1086_n 0.00286643f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_519 N_A_395_398#_c_560_n N_VPWR_c_1087_n 0.0100009f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_520 N_A_395_398#_M1003_g N_VPWR_c_1121_n 0.00426989f $X=6.985 $Y=2.465 $X2=0
+ $Y2=0
cc_521 N_A_395_398#_c_561_n N_VPWR_c_1121_n 0.00856429f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_522 N_A_395_398#_M1003_g N_VPWR_c_1089_n 0.00169308f $X=6.985 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A_395_398#_M1028_g N_VPWR_c_1089_n 0.0147834f $X=7.415 $Y=2.465 $X2=0
+ $Y2=0
cc_524 N_A_395_398#_M1003_g N_VPWR_c_1090_n 0.00487821f $X=6.985 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A_395_398#_M1028_g N_VPWR_c_1090_n 0.00486043f $X=7.415 $Y=2.465 $X2=0
+ $Y2=0
cc_526 N_A_395_398#_M1031_g N_VPWR_c_1083_n 9.39239e-19 $X=4.63 $Y=2.415 $X2=0
+ $Y2=0
cc_527 N_A_395_398#_M1003_g N_VPWR_c_1083_n 0.00459249f $X=6.985 $Y=2.465 $X2=0
+ $Y2=0
cc_528 N_A_395_398#_M1028_g N_VPWR_c_1083_n 0.00460886f $X=7.415 $Y=2.465 $X2=0
+ $Y2=0
cc_529 N_A_395_398#_c_553_n N_VPWR_c_1083_n 0.0135839f $X=8.785 $Y=1.99 $X2=0
+ $Y2=0
cc_530 N_A_395_398#_M1003_g N_VPWR_c_1101_n 0.014664f $X=6.985 $Y=2.465 $X2=0
+ $Y2=0
cc_531 N_A_395_398#_M1028_g N_VPWR_c_1101_n 0.001705f $X=7.415 $Y=2.465 $X2=0
+ $Y2=0
cc_532 N_A_395_398#_c_561_n N_VPWR_c_1101_n 0.00481536f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_533 N_A_395_398#_c_576_n N_SUM_M1007_s 0.00127262f $X=0.685 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_534 N_A_395_398#_c_542_n N_SUM_M1020_d 9.77818e-19 $X=0.595 $Y=1.92 $X2=0
+ $Y2=0
cc_535 N_A_395_398#_c_580_n N_SUM_M1020_d 2.67944e-19 $X=0.685 $Y=2.035 $X2=0
+ $Y2=0
cc_536 N_A_395_398#_c_558_n N_SUM_M1020_d 0.00192134f $X=2.02 $Y=2.035 $X2=0
+ $Y2=0
cc_537 N_A_395_398#_c_601_n N_SUM_M1020_d 0.00402378f $X=0.865 $Y=2.035 $X2=0
+ $Y2=0
cc_538 N_A_395_398#_c_543_n N_SUM_c_1216_n 0.012871f $X=1.055 $Y=1.16 $X2=0
+ $Y2=0
cc_539 N_A_395_398#_c_576_n N_SUM_c_1216_n 0.0128735f $X=0.685 $Y=1.16 $X2=0
+ $Y2=0
cc_540 N_A_395_398#_c_580_n N_SUM_c_1219_n 0.00561649f $X=0.685 $Y=2.035 $X2=0
+ $Y2=0
cc_541 N_A_395_398#_c_601_n N_SUM_c_1219_n 3.03435e-19 $X=0.865 $Y=2.035 $X2=0
+ $Y2=0
cc_542 N_A_395_398#_c_580_n N_SUM_c_1232_n 0.00442791f $X=0.685 $Y=2.035 $X2=0
+ $Y2=0
cc_543 N_A_395_398#_c_558_n N_SUM_c_1232_n 0.00788103f $X=2.02 $Y=2.035 $X2=0
+ $Y2=0
cc_544 N_A_395_398#_c_601_n N_SUM_c_1232_n 0.00400967f $X=0.865 $Y=2.035 $X2=0
+ $Y2=0
cc_545 N_A_395_398#_c_542_n SUM 0.0497497f $X=0.595 $Y=1.92 $X2=0 $Y2=0
cc_546 N_A_395_398#_c_576_n SUM 0.0137469f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_547 N_A_395_398#_c_580_n SUM 0.0171556f $X=0.685 $Y=2.035 $X2=0 $Y2=0
cc_548 N_A_395_398#_c_601_n SUM 0.0014554f $X=0.865 $Y=2.035 $X2=0 $Y2=0
cc_549 N_A_395_398#_c_558_n N_A_309_398#_M1027_d 0.00178113f $X=2.02 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_550 N_A_395_398#_c_560_n N_A_309_398#_M1012_s 0.00191144f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_551 N_A_395_398#_c_558_n N_A_309_398#_c_1262_n 0.0158193f $X=2.02 $Y=2.035
+ $X2=0 $Y2=0
cc_552 N_A_395_398#_c_559_n N_A_309_398#_c_1262_n 0.0123683f $X=2.115 $Y=2.135
+ $X2=0 $Y2=0
cc_553 N_A_395_398#_c_560_n N_A_309_398#_c_1262_n 0.00249677f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_554 N_A_395_398#_c_558_n N_A_309_398#_c_1263_n 0.00380171f $X=2.02 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_A_395_398#_c_559_n N_A_309_398#_c_1263_n 0.0198879f $X=2.115 $Y=2.135
+ $X2=0 $Y2=0
cc_556 N_A_395_398#_c_559_n N_A_309_398#_c_1265_n 0.0269231f $X=2.115 $Y=2.135
+ $X2=0 $Y2=0
cc_557 N_A_395_398#_c_560_n N_A_309_398#_c_1265_n 0.0182998f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_558 N_A_395_398#_c_560_n A_710_419# 0.00205389f $X=4.895 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_559 N_A_395_398#_c_562_n N_A_941_419#_M1031_d 0.00201707f $X=5.185 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_560 N_A_395_398#_c_565_n N_A_941_419#_M1031_d 0.00352405f $X=4.84 $Y=1.77
+ $X2=-0.19 $Y2=-0.245
cc_561 N_A_395_398#_c_561_n N_A_941_419#_c_1301_n 0.0172304f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_562 N_A_395_398#_c_562_n N_A_941_419#_c_1301_n 0.00294066f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_563 N_A_395_398#_c_561_n N_A_941_419#_c_1297_n 0.00736521f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_564 N_A_395_398#_M1031_g N_A_941_419#_c_1299_n 0.00876277f $X=4.63 $Y=2.415
+ $X2=0 $Y2=0
cc_565 N_A_395_398#_c_560_n N_A_941_419#_c_1299_n 8.23155e-19 $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_566 N_A_395_398#_c_562_n N_A_941_419#_c_1299_n 0.00676212f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_567 N_A_395_398#_c_551_n N_A_941_419#_c_1299_n 0.00106129f $X=4.84 $Y=1.77
+ $X2=0 $Y2=0
cc_568 N_A_395_398#_c_565_n N_A_941_419#_c_1299_n 0.0241561f $X=4.84 $Y=1.77
+ $X2=0 $Y2=0
cc_569 N_A_395_398#_c_561_n N_COUT_M1003_d 0.00171758f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_570 N_A_395_398#_c_537_n N_COUT_c_1333_n 0.00898441f $X=6.915 $Y=1.215 $X2=0
+ $Y2=0
cc_571 N_A_395_398#_M1003_g N_COUT_c_1333_n 0.00545094f $X=6.985 $Y=2.465 $X2=0
+ $Y2=0
cc_572 N_A_395_398#_c_539_n N_COUT_c_1333_n 0.0124834f $X=7.345 $Y=1.215 $X2=0
+ $Y2=0
cc_573 N_A_395_398#_c_541_n N_COUT_c_1333_n 0.00447255f $X=6.95 $Y=1.29 $X2=0
+ $Y2=0
cc_574 N_A_395_398#_c_544_n N_COUT_c_1333_n 0.0211729f $X=7.56 $Y=1.38 $X2=0
+ $Y2=0
cc_575 N_A_395_398#_c_545_n N_COUT_c_1333_n 0.00671667f $X=7.56 $Y=1.38 $X2=0
+ $Y2=0
cc_576 N_A_395_398#_c_547_n N_COUT_c_1333_n 0.01298f $X=7.645 $Y=1.16 $X2=0
+ $Y2=0
cc_577 N_A_395_398#_c_552_n N_COUT_c_1333_n 0.00997715f $X=7.27 $Y=1.38 $X2=0
+ $Y2=0
cc_578 N_A_395_398#_M1003_g COUT 0.0117103f $X=6.985 $Y=2.465 $X2=0 $Y2=0
cc_579 N_A_395_398#_M1028_g COUT 0.00423882f $X=7.415 $Y=2.465 $X2=0 $Y2=0
cc_580 N_A_395_398#_c_544_n COUT 7.36385e-19 $X=7.56 $Y=1.38 $X2=0 $Y2=0
cc_581 N_A_395_398#_c_545_n COUT 0.00123382f $X=7.56 $Y=1.38 $X2=0 $Y2=0
cc_582 N_A_395_398#_c_561_n COUT 0.0207307f $X=8.735 $Y=2.035 $X2=0 $Y2=0
cc_583 N_A_395_398#_c_561_n A_1653_367# 0.0159747f $X=8.735 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_584 N_A_395_398#_c_577_n N_VGND_M1008_d 0.00375252f $X=2.145 $Y=0.965 $X2=0
+ $Y2=0
cc_585 N_A_395_398#_c_548_n N_VGND_M1008_d 0.00300767f $X=1.14 $Y=0.965 $X2=0
+ $Y2=0
cc_586 N_A_395_398#_c_546_n N_VGND_M1016_s 0.00648266f $X=8.68 $Y=1.16 $X2=0
+ $Y2=0
cc_587 N_A_395_398#_c_547_n N_VGND_M1016_s 0.00269369f $X=7.645 $Y=1.16 $X2=0
+ $Y2=0
cc_588 N_A_395_398#_c_577_n N_VGND_c_1368_n 0.0080545f $X=2.145 $Y=0.965 $X2=0
+ $Y2=0
cc_589 N_A_395_398#_c_548_n N_VGND_c_1368_n 0.0143934f $X=1.14 $Y=0.965 $X2=0
+ $Y2=0
cc_590 N_A_395_398#_M1022_g N_VGND_c_1370_n 8.30893e-19 $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_591 N_A_395_398#_c_539_n N_VGND_c_1374_n 0.0063503f $X=7.345 $Y=1.215 $X2=0
+ $Y2=0
cc_592 N_A_395_398#_c_537_n N_VGND_c_1375_n 0.00384695f $X=6.915 $Y=1.215 $X2=0
+ $Y2=0
cc_593 N_A_395_398#_c_539_n N_VGND_c_1375_n 0.00384695f $X=7.345 $Y=1.215 $X2=0
+ $Y2=0
cc_594 N_A_395_398#_M1022_g N_VGND_c_1379_n 9.39239e-19 $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_595 N_A_395_398#_c_537_n N_VGND_c_1379_n 0.00642093f $X=6.915 $Y=1.215 $X2=0
+ $Y2=0
cc_596 N_A_395_398#_c_539_n N_VGND_c_1379_n 0.00642093f $X=7.345 $Y=1.215 $X2=0
+ $Y2=0
cc_597 N_A_395_398#_c_537_n N_VGND_c_1382_n 0.0063503f $X=6.915 $Y=1.215 $X2=0
+ $Y2=0
cc_598 N_A_395_398#_c_577_n N_A_309_131#_M1023_d 0.00921918f $X=2.145 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_599 N_A_395_398#_c_577_n N_A_309_131#_c_1473_n 0.00614315f $X=2.145 $Y=0.965
+ $X2=0 $Y2=0
cc_600 N_A_395_398#_c_549_n N_A_309_131#_c_1473_n 0.022378f $X=2.31 $Y=0.875
+ $X2=0 $Y2=0
cc_601 N_A_395_398#_c_549_n N_A_309_131#_c_1474_n 0.0157855f $X=2.31 $Y=0.875
+ $X2=0 $Y2=0
cc_602 N_A_395_398#_c_577_n N_A_309_131#_c_1475_n 0.0251704f $X=2.145 $Y=0.965
+ $X2=0 $Y2=0
cc_603 N_A_395_398#_M1022_g N_A_940_119#_c_1502_n 0.0050915f $X=4.625 $Y=0.805
+ $X2=0 $Y2=0
cc_604 N_A_395_398#_c_546_n A_1653_137# 0.0014993f $X=8.68 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_605 N_CIN_M1018_g N_B_M1023_g 0.0222335f $X=2.095 $Y=0.865 $X2=0 $Y2=0
cc_606 CIN N_B_M1023_g 9.71165e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_607 N_CIN_c_812_n N_B_M1023_g 0.0416577f $X=2.41 $Y=1.665 $X2=0 $Y2=0
cc_608 N_CIN_M1018_g N_B_c_917_n 0.00639096f $X=2.095 $Y=0.865 $X2=0 $Y2=0
cc_609 N_CIN_c_815_n N_B_M1029_g 0.0104164f $X=4.12 $Y=3.15 $X2=0 $Y2=0
cc_610 N_CIN_M1019_g N_B_M1029_g 0.151805f $X=4.195 $Y=0.805 $X2=0 $Y2=0
cc_611 N_CIN_M1019_g N_B_c_920_n 0.00979198f $X=4.195 $Y=0.805 $X2=0 $Y2=0
cc_612 N_CIN_M1015_g N_B_c_920_n 0.0103107f $X=5.055 $Y=0.805 $X2=0 $Y2=0
cc_613 N_CIN_M1015_g N_B_c_921_n 0.00172689f $X=5.055 $Y=0.805 $X2=0 $Y2=0
cc_614 N_CIN_c_810_n N_B_c_921_n 0.0252723f $X=5.29 $Y=1.29 $X2=0 $Y2=0
cc_615 N_CIN_M1005_g N_B_M1000_g 0.0378647f $X=5.29 $Y=2.54 $X2=0 $Y2=0
cc_616 N_CIN_M1015_g N_B_M1024_g 0.00431453f $X=5.055 $Y=0.805 $X2=0 $Y2=0
cc_617 N_CIN_c_810_n N_B_c_929_n 3.00385e-19 $X=5.29 $Y=1.29 $X2=0 $Y2=0
cc_618 N_CIN_c_814_n N_VPWR_c_1087_n 0.00240653f $X=2.41 $Y=3.075 $X2=0 $Y2=0
cc_619 N_CIN_c_815_n N_VPWR_c_1087_n 0.025796f $X=4.12 $Y=3.15 $X2=0 $Y2=0
cc_620 N_CIN_M1019_g N_VPWR_c_1087_n 0.00453189f $X=4.195 $Y=0.805 $X2=0 $Y2=0
cc_621 N_CIN_c_818_n N_VPWR_c_1088_n 0.00718254f $X=5.215 $Y=3.15 $X2=0 $Y2=0
cc_622 N_CIN_M1005_g N_VPWR_c_1088_n 0.0143866f $X=5.29 $Y=2.54 $X2=0 $Y2=0
cc_623 N_CIN_M1011_g N_VPWR_c_1093_n 2.40582e-19 $X=1.9 $Y=2.31 $X2=0 $Y2=0
cc_624 N_CIN_c_816_n N_VPWR_c_1093_n 0.0195441f $X=2.485 $Y=3.15 $X2=0 $Y2=0
cc_625 N_CIN_c_815_n N_VPWR_c_1094_n 0.0630258f $X=4.12 $Y=3.15 $X2=0 $Y2=0
cc_626 N_CIN_c_815_n N_VPWR_c_1083_n 0.0493564f $X=4.12 $Y=3.15 $X2=0 $Y2=0
cc_627 N_CIN_c_816_n N_VPWR_c_1083_n 0.00609198f $X=2.485 $Y=3.15 $X2=0 $Y2=0
cc_628 N_CIN_c_818_n N_VPWR_c_1083_n 0.034068f $X=5.215 $Y=3.15 $X2=0 $Y2=0
cc_629 N_CIN_c_820_n N_VPWR_c_1083_n 0.00845505f $X=4.195 $Y=3.15 $X2=0 $Y2=0
cc_630 N_CIN_M1011_g N_A_309_398#_c_1262_n 0.00797644f $X=1.9 $Y=2.31 $X2=0
+ $Y2=0
cc_631 N_CIN_c_814_n N_A_309_398#_c_1262_n 0.00222235f $X=2.41 $Y=3.075 $X2=0
+ $Y2=0
cc_632 N_CIN_M1011_g N_A_309_398#_c_1263_n 0.00448896f $X=1.9 $Y=2.31 $X2=0
+ $Y2=0
cc_633 N_CIN_c_814_n N_A_309_398#_c_1263_n 0.0182906f $X=2.41 $Y=3.075 $X2=0
+ $Y2=0
cc_634 N_CIN_c_815_n N_A_309_398#_c_1263_n 0.00768299f $X=4.12 $Y=3.15 $X2=0
+ $Y2=0
cc_635 N_CIN_c_814_n N_A_309_398#_c_1265_n 0.00992844f $X=2.41 $Y=3.075 $X2=0
+ $Y2=0
cc_636 N_CIN_M1005_g N_A_941_419#_c_1301_n 0.0137708f $X=5.29 $Y=2.54 $X2=0
+ $Y2=0
cc_637 N_CIN_M1005_g N_A_941_419#_c_1297_n 4.33356e-19 $X=5.29 $Y=2.54 $X2=0
+ $Y2=0
cc_638 N_CIN_M1019_g N_A_941_419#_c_1299_n 8.54173e-19 $X=4.195 $Y=0.805 $X2=0
+ $Y2=0
cc_639 N_CIN_c_818_n N_A_941_419#_c_1299_n 0.00726673f $X=5.215 $Y=3.15 $X2=0
+ $Y2=0
cc_640 N_CIN_M1005_g N_A_941_419#_c_1299_n 0.00774283f $X=5.29 $Y=2.54 $X2=0
+ $Y2=0
cc_641 N_CIN_M1015_g N_VGND_c_1370_n 0.00847923f $X=5.055 $Y=0.805 $X2=0 $Y2=0
cc_642 N_CIN_M1019_g N_VGND_c_1379_n 9.39239e-19 $X=4.195 $Y=0.805 $X2=0 $Y2=0
cc_643 N_CIN_M1015_g N_VGND_c_1379_n 7.88961e-19 $X=5.055 $Y=0.805 $X2=0 $Y2=0
cc_644 N_CIN_M1018_g N_A_309_131#_c_1473_n 0.00457109f $X=2.095 $Y=0.865 $X2=0
+ $Y2=0
cc_645 N_CIN_M1018_g N_A_309_131#_c_1474_n 0.00410955f $X=2.095 $Y=0.865 $X2=0
+ $Y2=0
cc_646 N_CIN_M1018_g N_A_309_131#_c_1475_n 0.00380175f $X=2.095 $Y=0.865 $X2=0
+ $Y2=0
cc_647 N_CIN_M1015_g N_A_940_119#_c_1501_n 0.014981f $X=5.055 $Y=0.805 $X2=0
+ $Y2=0
cc_648 N_CIN_c_810_n N_A_940_119#_c_1501_n 0.00642828f $X=5.29 $Y=1.29 $X2=0
+ $Y2=0
cc_649 N_B_M1023_g N_VPWR_c_1086_n 0.00297902f $X=1.47 $Y=0.865 $X2=0 $Y2=0
cc_650 N_B_M1029_g N_VPWR_c_1087_n 0.00318847f $X=3.835 $Y=0.805 $X2=0 $Y2=0
cc_651 N_B_M1000_g N_VPWR_c_1088_n 0.00191011f $X=5.76 $Y=2.54 $X2=0 $Y2=0
cc_652 N_B_M1000_g N_VPWR_c_1121_n 4.6693e-19 $X=5.76 $Y=2.54 $X2=0 $Y2=0
cc_653 N_B_M1023_g N_VPWR_c_1093_n 0.00324954f $X=1.47 $Y=0.865 $X2=0 $Y2=0
cc_654 N_B_M1000_g N_VPWR_c_1095_n 0.00505936f $X=5.76 $Y=2.54 $X2=0 $Y2=0
cc_655 N_B_M1014_g N_VPWR_c_1096_n 0.00312414f $X=8.55 $Y=2.155 $X2=0 $Y2=0
cc_656 N_B_M1023_g N_VPWR_c_1083_n 0.00375911f $X=1.47 $Y=0.865 $X2=0 $Y2=0
cc_657 N_B_M1029_g N_VPWR_c_1083_n 9.39239e-19 $X=3.835 $Y=0.805 $X2=0 $Y2=0
cc_658 N_B_M1000_g N_VPWR_c_1083_n 0.00514438f $X=5.76 $Y=2.54 $X2=0 $Y2=0
cc_659 N_B_M1014_g N_VPWR_c_1083_n 0.00410284f $X=8.55 $Y=2.155 $X2=0 $Y2=0
cc_660 N_B_M1023_g N_SUM_c_1216_n 7.13672e-19 $X=1.47 $Y=0.865 $X2=0 $Y2=0
cc_661 N_B_M1023_g N_A_309_398#_c_1262_n 0.00694783f $X=1.47 $Y=0.865 $X2=0
+ $Y2=0
cc_662 N_B_M1000_g N_A_941_419#_c_1301_n 0.00937766f $X=5.76 $Y=2.54 $X2=0 $Y2=0
cc_663 N_B_M1000_g N_A_941_419#_c_1297_n 0.00317937f $X=5.76 $Y=2.54 $X2=0 $Y2=0
cc_664 N_B_c_932_n N_COUT_M1004_d 0.00416244f $X=8.5 $Y=0.475 $X2=-0.19
+ $Y2=-0.245
cc_665 N_B_c_927_n N_COUT_c_1333_n 0.0151981f $X=6.525 $Y=1.42 $X2=0 $Y2=0
cc_666 N_B_c_928_n N_COUT_c_1333_n 0.0356585f $X=6.61 $Y=1.335 $X2=0 $Y2=0
cc_667 N_B_c_932_n N_COUT_c_1333_n 0.0240891f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_668 N_B_c_928_n N_VGND_M1026_d 0.0118428f $X=6.61 $Y=1.335 $X2=0 $Y2=0
cc_669 N_B_c_975_n N_VGND_M1026_d 0.00534743f $X=6.695 $Y=0.61 $X2=0 $Y2=0
cc_670 N_B_c_932_n N_VGND_M1026_d 0.00418611f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_671 N_B_c_932_n N_VGND_M1016_s 0.0132276f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_672 N_B_c_918_n N_VGND_c_1368_n 0.0102548f $X=1.545 $Y=0.18 $X2=0 $Y2=0
cc_673 N_B_c_917_n N_VGND_c_1369_n 0.0192621f $X=3.76 $Y=0.18 $X2=0 $Y2=0
cc_674 N_B_M1029_g N_VGND_c_1369_n 0.00615763f $X=3.835 $Y=0.805 $X2=0 $Y2=0
cc_675 N_B_c_920_n N_VGND_c_1370_n 0.0417382f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_676 N_B_M1024_g N_VGND_c_1370_n 0.0212207f $X=5.86 $Y=0.805 $X2=0 $Y2=0
cc_677 N_B_c_920_n N_VGND_c_1371_n 0.00486043f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_678 N_B_c_918_n N_VGND_c_1372_n 0.0448001f $X=1.545 $Y=0.18 $X2=0 $Y2=0
cc_679 N_B_c_931_n N_VGND_c_1374_n 0.00267868f $X=8.665 $Y=0.41 $X2=0 $Y2=0
cc_680 N_B_c_932_n N_VGND_c_1374_n 0.0240258f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_681 N_B_c_932_n N_VGND_c_1375_n 0.0131559f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_682 N_B_c_917_n N_VGND_c_1377_n 0.0492803f $X=3.76 $Y=0.18 $X2=0 $Y2=0
cc_683 B N_VGND_c_1378_n 0.035099f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_684 N_B_c_931_n N_VGND_c_1378_n 0.00627223f $X=8.665 $Y=0.41 $X2=0 $Y2=0
cc_685 N_B_c_932_n N_VGND_c_1378_n 0.0162603f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_686 N_B_c_917_n N_VGND_c_1379_n 0.0558311f $X=3.76 $Y=0.18 $X2=0 $Y2=0
cc_687 N_B_c_918_n N_VGND_c_1379_n 0.0103645f $X=1.545 $Y=0.18 $X2=0 $Y2=0
cc_688 N_B_c_920_n N_VGND_c_1379_n 0.0452207f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_689 N_B_c_925_n N_VGND_c_1379_n 0.00432325f $X=3.835 $Y=0.18 $X2=0 $Y2=0
cc_690 N_B_c_975_n N_VGND_c_1379_n 0.00107416f $X=6.695 $Y=0.61 $X2=0 $Y2=0
cc_691 B N_VGND_c_1379_n 0.0186639f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_692 N_B_c_931_n N_VGND_c_1379_n 0.0120379f $X=8.665 $Y=0.41 $X2=0 $Y2=0
cc_693 N_B_c_932_n N_VGND_c_1379_n 0.0439196f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_694 N_B_c_920_n N_VGND_c_1382_n 0.00339966f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_695 N_B_c_975_n N_VGND_c_1382_n 0.013757f $X=6.695 $Y=0.61 $X2=0 $Y2=0
cc_696 N_B_c_932_n N_VGND_c_1382_n 0.00642031f $X=8.5 $Y=0.475 $X2=0 $Y2=0
cc_697 N_B_c_917_n N_A_309_131#_c_1473_n 0.0203698f $X=3.76 $Y=0.18 $X2=0 $Y2=0
cc_698 N_B_M1023_g N_A_309_131#_c_1475_n 0.00574428f $X=1.47 $Y=0.865 $X2=0
+ $Y2=0
cc_699 N_B_c_917_n N_A_309_131#_c_1475_n 0.00739275f $X=3.76 $Y=0.18 $X2=0 $Y2=0
cc_700 N_B_c_920_n N_A_940_119#_c_1509_n 0.00397333f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_701 N_B_c_921_n N_A_940_119#_c_1501_n 0.00801231f $X=5.76 $Y=1.665 $X2=0
+ $Y2=0
cc_702 N_B_M1024_g N_A_940_119#_c_1501_n 0.0112562f $X=5.86 $Y=0.805 $X2=0 $Y2=0
cc_703 N_B_c_927_n N_A_940_119#_c_1501_n 0.0218611f $X=6.525 $Y=1.42 $X2=0 $Y2=0
cc_704 N_B_c_928_n N_A_940_119#_c_1501_n 0.00799556f $X=6.61 $Y=1.335 $X2=0
+ $Y2=0
cc_705 N_B_c_929_n N_A_940_119#_c_1501_n 0.0189287f $X=5.775 $Y=1.42 $X2=0 $Y2=0
cc_706 N_B_c_932_n A_1653_137# 0.0014993f $X=8.5 $Y=0.475 $X2=-0.19 $Y2=-0.245
cc_707 N_VPWR_c_1083_n N_SUM_M1020_d 0.00408483f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_708 N_VPWR_M1020_s N_SUM_c_1219_n 0.00131332f $X=0.155 $Y=1.835 $X2=0 $Y2=0
cc_709 N_VPWR_c_1085_n N_SUM_c_1219_n 0.00393958f $X=0.28 $Y=2.825 $X2=0 $Y2=0
cc_710 N_VPWR_c_1083_n N_SUM_c_1219_n 0.00526949f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_711 N_VPWR_c_1092_n N_SUM_c_1232_n 0.0124525f $X=0.975 $Y=3.33 $X2=0 $Y2=0
cc_712 N_VPWR_c_1083_n N_SUM_c_1232_n 0.00730901f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_713 N_VPWR_M1020_s SUM 0.00275377f $X=0.155 $Y=1.835 $X2=0 $Y2=0
cc_714 N_VPWR_c_1085_n SUM 0.0193613f $X=0.28 $Y=2.825 $X2=0 $Y2=0
cc_715 N_VPWR_c_1083_n SUM 0.00199722f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_716 N_VPWR_M1020_s SUM 0.00812813f $X=0.155 $Y=1.835 $X2=0 $Y2=0
cc_717 N_VPWR_c_1086_n N_A_309_398#_c_1262_n 0.026985f $X=1.185 $Y=2.425 $X2=0
+ $Y2=0
cc_718 N_VPWR_c_1087_n N_A_309_398#_c_1263_n 0.0142338f $X=3.26 $Y=2.25 $X2=0
+ $Y2=0
cc_719 N_VPWR_c_1093_n N_A_309_398#_c_1263_n 0.0457931f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_720 N_VPWR_c_1083_n N_A_309_398#_c_1263_n 0.0359575f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_721 N_VPWR_c_1086_n N_A_309_398#_c_1264_n 0.0151771f $X=1.185 $Y=2.425 $X2=0
+ $Y2=0
cc_722 N_VPWR_c_1093_n N_A_309_398#_c_1264_n 0.0153232f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_723 N_VPWR_c_1083_n N_A_309_398#_c_1264_n 0.0122547f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_724 N_VPWR_c_1087_n N_A_309_398#_c_1265_n 0.0275136f $X=3.26 $Y=2.25 $X2=0
+ $Y2=0
cc_725 N_VPWR_M1005_d N_A_941_419#_c_1301_n 0.00455106f $X=5.365 $Y=2.22 $X2=0
+ $Y2=0
cc_726 N_VPWR_c_1088_n N_A_941_419#_c_1301_n 0.0165244f $X=5.52 $Y=2.735 $X2=0
+ $Y2=0
cc_727 N_VPWR_c_1083_n N_A_941_419#_c_1301_n 0.0113958f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_728 N_VPWR_c_1083_n N_A_941_419#_c_1297_n 0.00147737f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_729 N_VPWR_c_1088_n N_A_941_419#_c_1298_n 0.00987822f $X=5.52 $Y=2.735 $X2=0
+ $Y2=0
cc_730 N_VPWR_c_1121_n N_A_941_419#_c_1298_n 0.0162497f $X=6.405 $Y=2.355 $X2=0
+ $Y2=0
cc_731 N_VPWR_c_1095_n N_A_941_419#_c_1298_n 0.00656181f $X=6.24 $Y=3.33 $X2=0
+ $Y2=0
cc_732 N_VPWR_c_1083_n N_A_941_419#_c_1298_n 0.00732212f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_733 N_VPWR_c_1088_n N_A_941_419#_c_1299_n 0.015434f $X=5.52 $Y=2.735 $X2=0
+ $Y2=0
cc_734 N_VPWR_c_1094_n N_A_941_419#_c_1299_n 0.0106152f $X=5.355 $Y=3.33 $X2=0
+ $Y2=0
cc_735 N_VPWR_c_1083_n N_A_941_419#_c_1299_n 0.0100662f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_736 N_VPWR_c_1083_n N_COUT_M1003_d 0.00408795f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_737 N_SUM_c_1216_n N_VGND_M1007_d 0.00131772f $X=0.545 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_738 N_SUM_c_1212_n N_VGND_M1007_d 0.00278905f $X=0.21 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_739 SUM N_VGND_M1007_d 0.00275868f $X=0.24 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_740 N_SUM_c_1212_n N_VGND_c_1366_n 5.10683e-19 $X=0.21 $Y=0.905 $X2=0 $Y2=0
cc_741 N_SUM_c_1216_n N_VGND_c_1367_n 0.00216437f $X=0.545 $Y=0.815 $X2=0 $Y2=0
cc_742 N_SUM_c_1212_n N_VGND_c_1367_n 0.0190579f $X=0.21 $Y=0.905 $X2=0 $Y2=0
cc_743 N_SUM_c_1216_n N_VGND_c_1376_n 0.00201199f $X=0.545 $Y=0.815 $X2=0 $Y2=0
cc_744 N_SUM_c_1220_n N_VGND_c_1376_n 0.0188748f $X=0.71 $Y=0.38 $X2=0 $Y2=0
cc_745 N_SUM_M1007_s N_VGND_c_1379_n 0.00223559f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_746 N_SUM_c_1216_n N_VGND_c_1379_n 0.00401697f $X=0.545 $Y=0.815 $X2=0 $Y2=0
cc_747 N_SUM_c_1220_n N_VGND_c_1379_n 0.012371f $X=0.71 $Y=0.38 $X2=0 $Y2=0
cc_748 N_SUM_c_1212_n N_VGND_c_1379_n 0.00184834f $X=0.21 $Y=0.905 $X2=0 $Y2=0
cc_749 N_VGND_c_1369_n N_A_309_131#_c_1473_n 0.0142263f $X=3.26 $Y=0.75 $X2=0
+ $Y2=0
cc_750 N_VGND_c_1372_n N_A_309_131#_c_1473_n 0.0395237f $X=3.165 $Y=0 $X2=0
+ $Y2=0
cc_751 N_VGND_c_1379_n N_A_309_131#_c_1473_n 0.0322225f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_752 N_VGND_c_1369_n N_A_309_131#_c_1474_n 0.0161313f $X=3.26 $Y=0.75 $X2=0
+ $Y2=0
cc_753 N_VGND_c_1368_n N_A_309_131#_c_1475_n 0.0182158f $X=1.16 $Y=0.545 $X2=0
+ $Y2=0
cc_754 N_VGND_c_1372_n N_A_309_131#_c_1475_n 0.0128859f $X=3.165 $Y=0 $X2=0
+ $Y2=0
cc_755 N_VGND_c_1379_n N_A_309_131#_c_1475_n 0.0103756f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_756 N_VGND_c_1377_n N_A_940_119#_c_1509_n 0.00370526f $X=5.105 $Y=0 $X2=0
+ $Y2=0
cc_757 N_VGND_c_1379_n N_A_940_119#_c_1509_n 0.00591522f $X=8.88 $Y=0 $X2=0
+ $Y2=0
cc_758 N_VGND_M1015_d N_A_940_119#_c_1501_n 0.00602962f $X=5.13 $Y=0.595 $X2=0
+ $Y2=0
cc_759 N_VGND_c_1370_n N_A_940_119#_c_1501_n 0.0475871f $X=5.645 $Y=0.74 $X2=0
+ $Y2=0
cc_760 N_VGND_c_1371_n N_A_940_119#_c_1519_n 0.00294932f $X=6.455 $Y=0 $X2=0
+ $Y2=0
cc_761 N_VGND_c_1379_n N_A_940_119#_c_1519_n 0.00559992f $X=8.88 $Y=0 $X2=0
+ $Y2=0
