* File: sky130_fd_sc_lp__nor4bb_lp.pxi.spice
* Created: Fri Aug 28 10:59:20 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%C_N N_C_N_c_102_n N_C_N_M1005_g N_C_N_c_103_n
+ N_C_N_M1007_g N_C_N_c_104_n N_C_N_c_105_n N_C_N_M1001_g N_C_N_c_111_n
+ N_C_N_c_106_n C_N C_N N_C_N_c_108_n N_C_N_c_109_n
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%C_N
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%A_27_409# N_A_27_409#_M1007_s
+ N_A_27_409#_M1005_s N_A_27_409#_M1008_g N_A_27_409#_M1016_g
+ N_A_27_409#_M1009_g N_A_27_409#_c_157_n N_A_27_409#_c_164_n
+ N_A_27_409#_c_165_n N_A_27_409#_c_158_n N_A_27_409#_c_159_n
+ N_A_27_409#_c_160_n N_A_27_409#_c_161_n N_A_27_409#_c_162_n
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%A_430_21# N_A_430_21#_M1017_d
+ N_A_430_21#_M1006_d N_A_430_21#_M1013_g N_A_430_21#_c_238_n
+ N_A_430_21#_c_239_n N_A_430_21#_M1014_g N_A_430_21#_M1000_g
+ N_A_430_21#_c_242_n N_A_430_21#_c_249_n N_A_430_21#_c_285_p
+ N_A_430_21#_c_250_n N_A_430_21#_c_243_n N_A_430_21#_c_244_n
+ N_A_430_21#_c_252_n N_A_430_21#_c_245_n N_A_430_21#_c_246_n
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%A_430_21#
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%B N_B_c_323_n N_B_M1002_g N_B_c_324_n
+ N_B_c_325_n N_B_c_326_n N_B_M1004_g N_B_c_327_n N_B_M1003_g N_B_c_329_n B
+ N_B_c_330_n PM_SKY130_FD_SC_LP__NOR4BB_LP%B
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%A N_A_c_373_n N_A_M1010_g N_A_c_374_n
+ N_A_c_375_n N_A_c_376_n N_A_M1012_g N_A_M1011_g N_A_c_378_n N_A_c_379_n A A
+ N_A_c_381_n PM_SKY130_FD_SC_LP__NOR4BB_LP%A
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%D_N N_D_N_M1015_g N_D_N_M1006_g N_D_N_M1017_g
+ D_N N_D_N_c_428_n N_D_N_c_429_n PM_SKY130_FD_SC_LP__NOR4BB_LP%D_N
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%VPWR N_VPWR_M1005_d N_VPWR_M1011_d
+ N_VPWR_c_458_n N_VPWR_c_459_n VPWR N_VPWR_c_460_n N_VPWR_c_461_n
+ N_VPWR_c_457_n N_VPWR_c_463_n N_VPWR_c_464_n
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%VPWR
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%A_245_409# N_A_245_409#_M1016_s
+ N_A_245_409#_M1000_d N_A_245_409#_c_499_n N_A_245_409#_c_500_n
+ N_A_245_409#_c_501_n N_A_245_409#_c_502_n
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%A_245_409#
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%A_352_409# N_A_352_409#_M1016_d
+ N_A_352_409#_M1003_s N_A_352_409#_c_532_n N_A_352_409#_c_533_n
+ N_A_352_409#_c_534_n N_A_352_409#_c_535_n N_A_352_409#_c_536_n
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%A_352_409#
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%Y N_Y_M1009_d N_Y_M1004_d N_Y_M1000_s
+ N_Y_c_560_n N_Y_c_563_n N_Y_c_602_n N_Y_c_561_n Y Y N_Y_c_565_n Y
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%Y
x_PM_SKY130_FD_SC_LP__NOR4BB_LP%VGND N_VGND_M1001_d N_VGND_M1014_d
+ N_VGND_M1012_d N_VGND_c_626_n N_VGND_c_627_n N_VGND_c_628_n VGND
+ N_VGND_c_629_n N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n
+ N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n
+ PM_SKY130_FD_SC_LP__NOR4BB_LP%VGND
cc_1 VNB N_C_N_c_102_n 0.0222849f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.658
cc_2 VNB N_C_N_c_103_n 0.0172366f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.73
cc_3 VNB N_C_N_c_104_n 0.0179281f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.805
cc_4 VNB N_C_N_c_105_n 0.013722f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.73
cc_5 VNB N_C_N_c_106_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.805
cc_6 VNB C_N 0.00500328f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_C_N_c_108_n 0.0194926f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.34
cc_8 VNB N_C_N_c_109_n 0.0196215f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.175
cc_9 VNB N_A_27_409#_M1008_g 0.0335127f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.445
cc_10 VNB N_A_27_409#_M1009_g 0.0284956f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.845
cc_11 VNB N_A_27_409#_c_157_n 0.0272131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_409#_c_158_n 0.0109159f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.665
cc_13 VNB N_A_27_409#_c_159_n 0.00148114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_409#_c_160_n 0.0153292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_409#_c_161_n 0.0315082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_409#_c_162_n 0.0769976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_430_21#_M1013_g 0.0317926f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.445
cc_18 VNB N_A_430_21#_c_238_n 0.0100692f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.175
cc_19 VNB N_A_430_21#_c_239_n 0.0086695f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.805
cc_20 VNB N_A_430_21#_M1014_g 0.0370598f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_21 VNB N_A_430_21#_M1000_g 0.00154414f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_A_430_21#_c_242_n 0.00104111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_430_21#_c_243_n 0.0483223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_430_21#_c_244_n 0.004557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_430_21#_c_245_n 0.0145699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_430_21#_c_246_n 0.0310763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_323_n 0.0142027f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.362
cc_28 VNB N_B_c_324_n 0.0101813f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_29 VNB N_B_c_325_n 0.00940486f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_30 VNB N_B_c_326_n 0.0135266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_c_327_n 0.0204828f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.88
cc_32 VNB N_B_M1003_g 0.0149455f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.805
cc_33 VNB N_B_c_329_n 0.00437176f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_34 VNB N_B_c_330_n 0.0556594f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.34
cc_35 VNB N_A_c_373_n 0.0140729f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.362
cc_36 VNB N_A_c_374_n 0.0151447f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_37 VNB N_A_c_375_n 0.00723986f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_38 VNB N_A_c_376_n 0.0152541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_M1011_g 0.0103916f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.175
cc_40 VNB N_A_c_378_n 0.0111627f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.73
cc_41 VNB N_A_c_379_n 0.0116736f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_42 VNB A 0.0158754f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.805
cc_43 VNB N_A_c_381_n 0.0295264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_D_N_M1015_g 0.0205446f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.845
cc_45 VNB N_D_N_M1006_g 0.0126755f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.73
cc_46 VNB N_D_N_M1017_g 0.0231466f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.175
cc_47 VNB N_D_N_c_428_n 0.0768822f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_48 VNB N_D_N_c_429_n 0.00296462f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.845
cc_49 VNB N_VPWR_c_457_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Y_c_560_n 0.0303342f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.88
cc_51 VNB N_Y_c_561_n 0.00275823f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_52 VNB Y 0.00289937f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.34
cc_53 VNB N_VGND_c_626_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.805
cc_54 VNB N_VGND_c_627_n 0.00283116f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_55 VNB N_VGND_c_628_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_56 VNB N_VGND_c_629_n 0.0302588f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.34
cc_57 VNB N_VGND_c_630_n 0.0319926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_631_n 0.0384538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_632_n 0.034917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_633_n 0.293059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_634_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_635_n 0.00511034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_636_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_C_N_M1005_g 0.039241f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_65 VPB N_C_N_c_111_n 0.0184705f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.845
cc_66 VPB C_N 0.00338093f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_67 VPB N_A_27_409#_M1016_g 0.0463352f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.805
cc_68 VPB N_A_27_409#_c_164_n 0.00810785f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.34
cc_69 VPB N_A_27_409#_c_165_n 0.0357032f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.295
cc_70 VPB N_A_27_409#_c_159_n 0.00795773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_27_409#_c_161_n 0.0177946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_27_409#_c_162_n 0.034231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_430_21#_M1000_g 0.0321265f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_74 VPB N_A_430_21#_c_242_n 0.00546222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_430_21#_c_249_n 0.0470551f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.34
cc_76 VPB N_A_430_21#_c_250_n 0.0682556f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.295
cc_77 VPB N_A_430_21#_c_243_n 8.91883e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_430_21#_c_252_n 0.0173977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_B_M1003_g 0.0499702f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.805
cc_80 VPB N_A_M1011_g 0.0387666f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.175
cc_81 VPB N_D_N_M1006_g 0.0477496f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.73
cc_82 VPB N_VPWR_c_458_n 0.020253f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.175
cc_83 VPB N_VPWR_c_459_n 0.00712932f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.845
cc_84 VPB N_VPWR_c_460_n 0.0870991f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.34
cc_85 VPB N_VPWR_c_461_n 0.0290594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_457_n 0.094948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_463_n 0.0251504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_464_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_245_409#_c_499_n 0.00578548f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.73
cc_90 VPB N_A_245_409#_c_500_n 0.00860266f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.445
cc_91 VPB N_A_245_409#_c_501_n 0.00835883f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.175
cc_92 VPB N_A_245_409#_c_502_n 0.00896709f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.805
cc_93 VPB N_A_352_409#_c_532_n 0.00716906f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.445
cc_94 VPB N_A_352_409#_c_533_n 0.0386413f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.175
cc_95 VPB N_A_352_409#_c_534_n 0.00244612f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.805
cc_96 VPB N_A_352_409#_c_535_n 0.00246318f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.805
cc_97 VPB N_A_352_409#_c_536_n 0.0127542f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.445
cc_98 VPB N_Y_c_563_n 0.00437887f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.73
cc_99 VPB Y 0.00249981f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.34
cc_100 VPB N_Y_c_565_n 0.00990818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 N_C_N_c_105_n N_A_27_409#_M1008_g 0.0179709f $X=1.005 $Y=0.73 $X2=0 $Y2=0
cc_102 N_C_N_c_109_n N_A_27_409#_M1008_g 0.00279816f $X=0.607 $Y=1.175 $X2=0
+ $Y2=0
cc_103 N_C_N_c_111_n N_A_27_409#_M1016_g 6.07098e-19 $X=0.607 $Y=1.845 $X2=0
+ $Y2=0
cc_104 C_N N_A_27_409#_M1016_g 8.69183e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_105 N_C_N_c_103_n N_A_27_409#_c_157_n 0.00961612f $X=0.645 $Y=0.73 $X2=0
+ $Y2=0
cc_106 N_C_N_c_105_n N_A_27_409#_c_157_n 0.00145013f $X=1.005 $Y=0.73 $X2=0
+ $Y2=0
cc_107 N_C_N_c_106_n N_A_27_409#_c_157_n 0.00668784f $X=0.645 $Y=0.805 $X2=0
+ $Y2=0
cc_108 N_C_N_M1005_g N_A_27_409#_c_164_n 0.00104139f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_109 N_C_N_c_104_n N_A_27_409#_c_158_n 0.0156514f $X=0.93 $Y=0.805 $X2=0 $Y2=0
cc_110 N_C_N_c_106_n N_A_27_409#_c_158_n 0.00357648f $X=0.645 $Y=0.805 $X2=0
+ $Y2=0
cc_111 C_N N_A_27_409#_c_158_n 0.0179397f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_112 N_C_N_c_108_n N_A_27_409#_c_158_n 2.40353e-19 $X=0.63 $Y=1.34 $X2=0 $Y2=0
cc_113 N_C_N_c_109_n N_A_27_409#_c_158_n 0.00531063f $X=0.607 $Y=1.175 $X2=0
+ $Y2=0
cc_114 C_N N_A_27_409#_c_159_n 0.0405176f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_C_N_c_108_n N_A_27_409#_c_159_n 7.32632e-19 $X=0.63 $Y=1.34 $X2=0 $Y2=0
cc_116 N_C_N_c_109_n N_A_27_409#_c_159_n 0.00305204f $X=0.607 $Y=1.175 $X2=0
+ $Y2=0
cc_117 N_C_N_c_106_n N_A_27_409#_c_160_n 0.00134476f $X=0.645 $Y=0.805 $X2=0
+ $Y2=0
cc_118 C_N N_A_27_409#_c_160_n 0.0108863f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_119 N_C_N_c_108_n N_A_27_409#_c_160_n 0.00300934f $X=0.63 $Y=1.34 $X2=0 $Y2=0
cc_120 N_C_N_c_109_n N_A_27_409#_c_160_n 0.00315954f $X=0.607 $Y=1.175 $X2=0
+ $Y2=0
cc_121 C_N N_A_27_409#_c_161_n 0.0485802f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_122 N_C_N_c_108_n N_A_27_409#_c_161_n 0.0228214f $X=0.63 $Y=1.34 $X2=0 $Y2=0
cc_123 N_C_N_c_109_n N_A_27_409#_c_161_n 0.00541891f $X=0.607 $Y=1.175 $X2=0
+ $Y2=0
cc_124 N_C_N_c_104_n N_A_27_409#_c_162_n 0.00139458f $X=0.93 $Y=0.805 $X2=0
+ $Y2=0
cc_125 C_N N_A_27_409#_c_162_n 0.00434786f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_126 N_C_N_c_108_n N_A_27_409#_c_162_n 0.0312331f $X=0.63 $Y=1.34 $X2=0 $Y2=0
cc_127 N_C_N_c_109_n N_A_27_409#_c_162_n 0.00232995f $X=0.607 $Y=1.175 $X2=0
+ $Y2=0
cc_128 N_C_N_M1005_g N_VPWR_c_458_n 0.0231779f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_129 N_C_N_c_111_n N_VPWR_c_458_n 9.71192e-19 $X=0.607 $Y=1.845 $X2=0 $Y2=0
cc_130 C_N N_VPWR_c_458_n 0.0161006f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_131 N_C_N_M1005_g N_VPWR_c_457_n 0.0149742f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_132 N_C_N_M1005_g N_VPWR_c_463_n 0.00802402f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_133 N_C_N_M1005_g N_A_245_409#_c_499_n 6.72974e-19 $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_134 N_C_N_M1005_g N_A_245_409#_c_500_n 0.0012739f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_135 N_C_N_c_103_n N_VGND_c_626_n 0.00231629f $X=0.645 $Y=0.73 $X2=0 $Y2=0
cc_136 N_C_N_c_105_n N_VGND_c_626_n 0.011926f $X=1.005 $Y=0.73 $X2=0 $Y2=0
cc_137 N_C_N_c_103_n N_VGND_c_629_n 0.00549284f $X=0.645 $Y=0.73 $X2=0 $Y2=0
cc_138 N_C_N_c_104_n N_VGND_c_629_n 4.87571e-19 $X=0.93 $Y=0.805 $X2=0 $Y2=0
cc_139 N_C_N_c_105_n N_VGND_c_629_n 0.00486043f $X=1.005 $Y=0.73 $X2=0 $Y2=0
cc_140 N_C_N_c_103_n N_VGND_c_633_n 0.0072374f $X=0.645 $Y=0.73 $X2=0 $Y2=0
cc_141 N_C_N_c_104_n N_VGND_c_633_n 6.51792e-19 $X=0.93 $Y=0.805 $X2=0 $Y2=0
cc_142 N_C_N_c_105_n N_VGND_c_633_n 0.00436085f $X=1.005 $Y=0.73 $X2=0 $Y2=0
cc_143 N_A_27_409#_M1009_g N_A_430_21#_M1013_g 0.0191545f $X=1.795 $Y=0.445
+ $X2=0 $Y2=0
cc_144 N_A_27_409#_c_162_n N_A_430_21#_c_239_n 0.0191545f $X=1.795 $Y=1.455
+ $X2=0 $Y2=0
cc_145 N_A_27_409#_c_162_n N_A_430_21#_c_246_n 0.00213773f $X=1.795 $Y=1.455
+ $X2=0 $Y2=0
cc_146 N_A_27_409#_M1016_g N_VPWR_c_458_n 0.00380322f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_147 N_A_27_409#_c_164_n N_VPWR_c_458_n 0.0272606f $X=0.24 $Y=2.15 $X2=0 $Y2=0
cc_148 N_A_27_409#_M1016_g N_VPWR_c_460_n 0.00825264f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_149 N_A_27_409#_M1016_g N_VPWR_c_457_n 0.0166629f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_150 N_A_27_409#_c_165_n N_VPWR_c_457_n 0.0095959f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_151 N_A_27_409#_c_165_n N_VPWR_c_463_n 0.0167213f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_152 N_A_27_409#_M1016_g N_A_245_409#_c_499_n 0.00921512f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_153 N_A_27_409#_c_159_n N_A_245_409#_c_499_n 0.0125024f $X=1.22 $Y=1.285
+ $X2=0 $Y2=0
cc_154 N_A_27_409#_c_162_n N_A_245_409#_c_499_n 0.00703416f $X=1.795 $Y=1.455
+ $X2=0 $Y2=0
cc_155 N_A_27_409#_M1016_g N_A_245_409#_c_500_n 0.0178196f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_156 N_A_27_409#_M1016_g N_A_245_409#_c_501_n 0.0210588f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_157 N_A_27_409#_c_162_n N_A_245_409#_c_501_n 0.00226141f $X=1.795 $Y=1.455
+ $X2=0 $Y2=0
cc_158 N_A_27_409#_M1016_g N_A_352_409#_c_532_n 0.00805817f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_159 N_A_27_409#_M1016_g N_A_352_409#_c_534_n 0.00497284f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_160 N_A_27_409#_M1008_g N_Y_c_561_n 0.0074673f $X=1.435 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_27_409#_M1009_g N_Y_c_561_n 0.019602f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_27_409#_c_158_n N_Y_c_561_n 0.0136557f $X=1.055 $Y=0.91 $X2=0 $Y2=0
cc_163 N_A_27_409#_M1008_g Y 9.80258e-19 $X=1.435 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_27_409#_M1009_g Y 0.0041955f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_27_409#_c_158_n Y 8.07588e-19 $X=1.055 $Y=0.91 $X2=0 $Y2=0
cc_166 N_A_27_409#_c_159_n Y 0.0522305f $X=1.22 $Y=1.285 $X2=0 $Y2=0
cc_167 N_A_27_409#_c_162_n Y 0.0342675f $X=1.795 $Y=1.455 $X2=0 $Y2=0
cc_168 N_A_27_409#_M1016_g N_Y_c_565_n 0.00738618f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_169 N_A_27_409#_c_159_n N_Y_c_565_n 0.00800389f $X=1.22 $Y=1.285 $X2=0 $Y2=0
cc_170 N_A_27_409#_c_162_n N_Y_c_565_n 0.013968f $X=1.795 $Y=1.455 $X2=0 $Y2=0
cc_171 N_A_27_409#_M1008_g N_VGND_c_626_n 0.00976273f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_172 N_A_27_409#_M1009_g N_VGND_c_626_n 0.00158064f $X=1.795 $Y=0.445 $X2=0
+ $Y2=0
cc_173 N_A_27_409#_c_157_n N_VGND_c_626_n 0.0130887f $X=0.43 $Y=0.47 $X2=0 $Y2=0
cc_174 N_A_27_409#_c_158_n N_VGND_c_626_n 0.0227656f $X=1.055 $Y=0.91 $X2=0
+ $Y2=0
cc_175 N_A_27_409#_c_162_n N_VGND_c_626_n 9.7121e-19 $X=1.795 $Y=1.455 $X2=0
+ $Y2=0
cc_176 N_A_27_409#_c_157_n N_VGND_c_629_n 0.0299021f $X=0.43 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A_27_409#_M1008_g N_VGND_c_630_n 0.00486043f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A_27_409#_M1009_g N_VGND_c_630_n 0.00359757f $X=1.795 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_27_409#_M1007_s N_VGND_c_633_n 0.00232985f $X=0.285 $Y=0.235 $X2=0
+ $Y2=0
cc_180 N_A_27_409#_M1008_g N_VGND_c_633_n 0.00814425f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_27_409#_M1009_g N_VGND_c_633_n 0.00523988f $X=1.795 $Y=0.445 $X2=0
+ $Y2=0
cc_182 N_A_27_409#_c_157_n N_VGND_c_633_n 0.0183848f $X=0.43 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A_27_409#_c_158_n N_VGND_c_633_n 0.0147838f $X=1.055 $Y=0.91 $X2=0
+ $Y2=0
cc_184 N_A_430_21#_M1014_g N_B_c_323_n 0.0173235f $X=2.585 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_430_21#_M1014_g N_B_c_327_n 0.00518129f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A_430_21#_c_249_n N_B_M1003_g 0.0298834f $X=4.975 $Y=1.76 $X2=0 $Y2=0
cc_187 N_A_430_21#_c_249_n B 0.0236618f $X=4.975 $Y=1.76 $X2=0 $Y2=0
cc_188 N_A_430_21#_c_244_n B 0.0139054f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_189 N_A_430_21#_c_246_n B 3.19059e-19 $X=2.68 $Y=1.24 $X2=0 $Y2=0
cc_190 N_A_430_21#_c_249_n N_B_c_330_n 0.00942295f $X=4.975 $Y=1.76 $X2=0 $Y2=0
cc_191 N_A_430_21#_c_244_n N_B_c_330_n 0.0031225f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_192 N_A_430_21#_c_246_n N_B_c_330_n 0.00717526f $X=2.68 $Y=1.24 $X2=0 $Y2=0
cc_193 N_A_430_21#_c_249_n N_A_M1011_g 0.0217391f $X=4.975 $Y=1.76 $X2=0 $Y2=0
cc_194 N_A_430_21#_c_250_n N_A_M1011_g 0.00105557f $X=5.14 $Y=2.19 $X2=0 $Y2=0
cc_195 N_A_430_21#_c_249_n N_A_c_379_n 0.00206279f $X=4.975 $Y=1.76 $X2=0 $Y2=0
cc_196 N_A_430_21#_c_249_n A 0.0548185f $X=4.975 $Y=1.76 $X2=0 $Y2=0
cc_197 N_A_430_21#_c_245_n N_D_N_M1015_g 0.00114698f $X=5.43 $Y=0.455 $X2=0
+ $Y2=0
cc_198 N_A_430_21#_c_249_n N_D_N_M1006_g 0.0220008f $X=4.975 $Y=1.76 $X2=0 $Y2=0
cc_199 N_A_430_21#_c_250_n N_D_N_M1006_g 0.0239601f $X=5.14 $Y=2.19 $X2=0 $Y2=0
cc_200 N_A_430_21#_c_243_n N_D_N_M1006_g 0.00359279f $X=5.51 $Y=1.675 $X2=0
+ $Y2=0
cc_201 N_A_430_21#_c_252_n N_D_N_M1006_g 0.00472289f $X=5.285 $Y=1.76 $X2=0
+ $Y2=0
cc_202 N_A_430_21#_c_243_n N_D_N_M1017_g 0.0225129f $X=5.51 $Y=1.675 $X2=0 $Y2=0
cc_203 N_A_430_21#_c_245_n N_D_N_M1017_g 0.00844626f $X=5.43 $Y=0.455 $X2=0
+ $Y2=0
cc_204 N_A_430_21#_c_252_n N_D_N_c_428_n 0.00650287f $X=5.285 $Y=1.76 $X2=0
+ $Y2=0
cc_205 N_A_430_21#_c_249_n N_D_N_c_429_n 0.00861307f $X=4.975 $Y=1.76 $X2=0
+ $Y2=0
cc_206 N_A_430_21#_c_243_n N_D_N_c_429_n 0.0388942f $X=5.51 $Y=1.675 $X2=0 $Y2=0
cc_207 N_A_430_21#_c_252_n N_D_N_c_429_n 0.0177081f $X=5.285 $Y=1.76 $X2=0 $Y2=0
cc_208 N_A_430_21#_c_249_n N_VPWR_c_459_n 0.0264018f $X=4.975 $Y=1.76 $X2=0
+ $Y2=0
cc_209 N_A_430_21#_c_250_n N_VPWR_c_459_n 0.0338651f $X=5.14 $Y=2.19 $X2=0 $Y2=0
cc_210 N_A_430_21#_c_250_n N_VPWR_c_461_n 0.0415852f $X=5.14 $Y=2.19 $X2=0 $Y2=0
cc_211 N_A_430_21#_c_250_n N_VPWR_c_457_n 0.0238018f $X=5.14 $Y=2.19 $X2=0 $Y2=0
cc_212 N_A_430_21#_c_249_n N_A_245_409#_M1000_d 0.0025972f $X=4.975 $Y=1.76
+ $X2=0 $Y2=0
cc_213 N_A_430_21#_c_285_p N_A_245_409#_M1000_d 7.44328e-19 $X=2.975 $Y=1.76
+ $X2=0 $Y2=0
cc_214 N_A_430_21#_M1000_g N_A_245_409#_c_501_n 0.0198224f $X=2.725 $Y=2.195
+ $X2=0 $Y2=0
cc_215 N_A_430_21#_M1000_g N_A_245_409#_c_502_n 0.0244525f $X=2.725 $Y=2.195
+ $X2=0 $Y2=0
cc_216 N_A_430_21#_c_249_n N_A_245_409#_c_502_n 0.0140765f $X=4.975 $Y=1.76
+ $X2=0 $Y2=0
cc_217 N_A_430_21#_c_285_p N_A_245_409#_c_502_n 0.0074927f $X=2.975 $Y=1.76
+ $X2=0 $Y2=0
cc_218 N_A_430_21#_M1000_g N_A_352_409#_c_532_n 0.00776016f $X=2.725 $Y=2.195
+ $X2=0 $Y2=0
cc_219 N_A_430_21#_M1000_g N_A_352_409#_c_533_n 0.00846208f $X=2.725 $Y=2.195
+ $X2=0 $Y2=0
cc_220 N_A_430_21#_M1000_g N_A_352_409#_c_536_n 0.00418213f $X=2.725 $Y=2.195
+ $X2=0 $Y2=0
cc_221 N_A_430_21#_c_249_n N_A_352_409#_c_536_n 0.0264016f $X=4.975 $Y=1.76
+ $X2=0 $Y2=0
cc_222 N_A_430_21#_M1013_g N_Y_c_560_n 0.0034451f $X=2.225 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A_430_21#_c_238_n N_Y_c_560_n 0.00101607f $X=2.51 $Y=1.24 $X2=0 $Y2=0
cc_224 N_A_430_21#_M1014_g N_Y_c_560_n 0.0125233f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_430_21#_c_244_n N_Y_c_560_n 0.032747f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_226 N_A_430_21#_c_246_n N_Y_c_560_n 0.00497309f $X=2.68 $Y=1.24 $X2=0 $Y2=0
cc_227 N_A_430_21#_c_239_n N_Y_c_563_n 0.00828554f $X=2.3 $Y=1.24 $X2=0 $Y2=0
cc_228 N_A_430_21#_M1000_g N_Y_c_563_n 0.011505f $X=2.725 $Y=2.195 $X2=0 $Y2=0
cc_229 N_A_430_21#_c_285_p N_Y_c_563_n 0.0135525f $X=2.975 $Y=1.76 $X2=0 $Y2=0
cc_230 N_A_430_21#_c_244_n N_Y_c_563_n 0.00785717f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_231 N_A_430_21#_c_246_n N_Y_c_563_n 0.00256273f $X=2.68 $Y=1.24 $X2=0 $Y2=0
cc_232 N_A_430_21#_M1013_g N_Y_c_561_n 0.0181986f $X=2.225 $Y=0.445 $X2=0 $Y2=0
cc_233 N_A_430_21#_M1014_g N_Y_c_561_n 0.00189981f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_234 N_A_430_21#_M1013_g Y 0.00677065f $X=2.225 $Y=0.445 $X2=0 $Y2=0
cc_235 N_A_430_21#_c_239_n Y 0.00912225f $X=2.3 $Y=1.24 $X2=0 $Y2=0
cc_236 N_A_430_21#_M1014_g Y 0.00110327f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A_430_21#_M1000_g Y 0.00399373f $X=2.725 $Y=2.195 $X2=0 $Y2=0
cc_238 N_A_430_21#_c_242_n Y 0.00616868f $X=2.89 $Y=1.675 $X2=0 $Y2=0
cc_239 N_A_430_21#_c_244_n Y 0.0208997f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_240 N_A_430_21#_c_246_n Y 0.00197975f $X=2.68 $Y=1.24 $X2=0 $Y2=0
cc_241 N_A_430_21#_M1013_g N_VGND_c_627_n 0.00228849f $X=2.225 $Y=0.445 $X2=0
+ $Y2=0
cc_242 N_A_430_21#_M1014_g N_VGND_c_627_n 0.011648f $X=2.585 $Y=0.445 $X2=0
+ $Y2=0
cc_243 N_A_430_21#_c_245_n N_VGND_c_628_n 0.0104495f $X=5.43 $Y=0.455 $X2=0
+ $Y2=0
cc_244 N_A_430_21#_M1013_g N_VGND_c_630_n 0.0054778f $X=2.225 $Y=0.445 $X2=0
+ $Y2=0
cc_245 N_A_430_21#_M1014_g N_VGND_c_630_n 0.00486043f $X=2.585 $Y=0.445 $X2=0
+ $Y2=0
cc_246 N_A_430_21#_c_245_n N_VGND_c_632_n 0.0194886f $X=5.43 $Y=0.455 $X2=0
+ $Y2=0
cc_247 N_A_430_21#_M1017_d N_VGND_c_633_n 0.00232985f $X=5.29 $Y=0.235 $X2=0
+ $Y2=0
cc_248 N_A_430_21#_M1013_g N_VGND_c_633_n 0.00611135f $X=2.225 $Y=0.445 $X2=0
+ $Y2=0
cc_249 N_A_430_21#_M1014_g N_VGND_c_633_n 0.00435613f $X=2.585 $Y=0.445 $X2=0
+ $Y2=0
cc_250 N_A_430_21#_c_245_n N_VGND_c_633_n 0.0124792f $X=5.43 $Y=0.455 $X2=0
+ $Y2=0
cc_251 N_B_c_326_n N_A_c_373_n 0.00935182f $X=3.405 $Y=0.73 $X2=-0.19 $Y2=-0.245
cc_252 N_B_c_329_n N_A_c_375_n 0.00935182f $X=3.405 $Y=0.805 $X2=0 $Y2=0
cc_253 N_B_c_330_n N_A_c_375_n 0.010912f $X=3.815 $Y=1.33 $X2=0 $Y2=0
cc_254 N_B_M1003_g N_A_c_379_n 0.0565688f $X=3.815 $Y=2.545 $X2=0 $Y2=0
cc_255 N_B_c_327_n A 0.00413803f $X=3.405 $Y=1.165 $X2=0 $Y2=0
cc_256 B A 0.0208786f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_257 N_B_c_330_n A 0.00370257f $X=3.815 $Y=1.33 $X2=0 $Y2=0
cc_258 N_B_c_327_n N_A_c_381_n 0.00285432f $X=3.405 $Y=1.165 $X2=0 $Y2=0
cc_259 B N_A_c_381_n 2.21262e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_260 N_B_c_330_n N_A_c_381_n 0.0565688f $X=3.815 $Y=1.33 $X2=0 $Y2=0
cc_261 N_B_M1003_g N_VPWR_c_459_n 0.00519241f $X=3.815 $Y=2.545 $X2=0 $Y2=0
cc_262 N_B_M1003_g N_VPWR_c_460_n 0.0085862f $X=3.815 $Y=2.545 $X2=0 $Y2=0
cc_263 N_B_M1003_g N_VPWR_c_457_n 0.0165862f $X=3.815 $Y=2.545 $X2=0 $Y2=0
cc_264 N_B_M1003_g N_A_245_409#_c_502_n 6.72974e-19 $X=3.815 $Y=2.545 $X2=0
+ $Y2=0
cc_265 N_B_M1003_g N_A_352_409#_c_535_n 0.00427649f $X=3.815 $Y=2.545 $X2=0
+ $Y2=0
cc_266 N_B_M1003_g N_A_352_409#_c_536_n 0.0178231f $X=3.815 $Y=2.545 $X2=0 $Y2=0
cc_267 N_B_c_324_n N_Y_c_560_n 0.00944489f $X=3.33 $Y=0.805 $X2=0 $Y2=0
cc_268 N_B_c_325_n N_Y_c_560_n 0.00771533f $X=3.12 $Y=0.805 $X2=0 $Y2=0
cc_269 N_B_c_327_n N_Y_c_560_n 0.00893692f $X=3.405 $Y=1.165 $X2=0 $Y2=0
cc_270 N_B_c_329_n N_Y_c_560_n 0.00459419f $X=3.405 $Y=0.805 $X2=0 $Y2=0
cc_271 B N_Y_c_560_n 0.0257309f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_272 N_B_c_330_n N_Y_c_560_n 0.00841653f $X=3.815 $Y=1.33 $X2=0 $Y2=0
cc_273 N_B_c_323_n N_Y_c_602_n 0.00149562f $X=3.045 $Y=0.73 $X2=0 $Y2=0
cc_274 N_B_c_326_n N_Y_c_602_n 0.0088976f $X=3.405 $Y=0.73 $X2=0 $Y2=0
cc_275 N_B_c_329_n N_Y_c_602_n 0.00495788f $X=3.405 $Y=0.805 $X2=0 $Y2=0
cc_276 N_B_c_323_n N_VGND_c_627_n 0.00333146f $X=3.045 $Y=0.73 $X2=0 $Y2=0
cc_277 N_B_c_323_n N_VGND_c_631_n 0.00585385f $X=3.045 $Y=0.73 $X2=0 $Y2=0
cc_278 N_B_c_324_n N_VGND_c_631_n 4.87571e-19 $X=3.33 $Y=0.805 $X2=0 $Y2=0
cc_279 N_B_c_326_n N_VGND_c_631_n 0.00549284f $X=3.405 $Y=0.73 $X2=0 $Y2=0
cc_280 N_B_c_323_n N_VGND_c_633_n 0.00602236f $X=3.045 $Y=0.73 $X2=0 $Y2=0
cc_281 N_B_c_324_n N_VGND_c_633_n 6.51792e-19 $X=3.33 $Y=0.805 $X2=0 $Y2=0
cc_282 N_B_c_326_n N_VGND_c_633_n 0.00610391f $X=3.405 $Y=0.73 $X2=0 $Y2=0
cc_283 N_A_c_376_n N_D_N_M1015_g 0.0146702f $X=4.255 $Y=0.73 $X2=0 $Y2=0
cc_284 N_A_M1011_g N_D_N_M1006_g 0.0288697f $X=4.305 $Y=2.545 $X2=0 $Y2=0
cc_285 N_A_c_378_n N_D_N_c_428_n 0.0361179f $X=4.18 $Y=0.73 $X2=0 $Y2=0
cc_286 A N_D_N_c_428_n 0.00575307f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_287 N_A_c_378_n N_D_N_c_429_n 5.38516e-19 $X=4.18 $Y=0.73 $X2=0 $Y2=0
cc_288 A N_D_N_c_429_n 0.0541474f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_289 N_A_M1011_g N_VPWR_c_459_n 0.025411f $X=4.305 $Y=2.545 $X2=0 $Y2=0
cc_290 N_A_M1011_g N_VPWR_c_460_n 0.00802402f $X=4.305 $Y=2.545 $X2=0 $Y2=0
cc_291 N_A_M1011_g N_VPWR_c_457_n 0.0142664f $X=4.305 $Y=2.545 $X2=0 $Y2=0
cc_292 N_A_M1011_g N_A_352_409#_c_535_n 7.28154e-19 $X=4.305 $Y=2.545 $X2=0
+ $Y2=0
cc_293 N_A_M1011_g N_A_352_409#_c_536_n 0.00375854f $X=4.305 $Y=2.545 $X2=0
+ $Y2=0
cc_294 N_A_c_375_n N_Y_c_560_n 0.00238434f $X=3.91 $Y=0.805 $X2=0 $Y2=0
cc_295 A N_Y_c_560_n 0.0138537f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_296 N_A_c_381_n N_Y_c_560_n 3.24343e-19 $X=4.345 $Y=0.99 $X2=0 $Y2=0
cc_297 N_A_c_373_n N_Y_c_602_n 0.00926343f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_298 N_A_c_375_n N_Y_c_602_n 0.00499729f $X=3.91 $Y=0.805 $X2=0 $Y2=0
cc_299 N_A_c_376_n N_Y_c_602_n 0.0015204f $X=4.255 $Y=0.73 $X2=0 $Y2=0
cc_300 N_A_c_373_n N_VGND_c_628_n 0.00230093f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_301 N_A_c_376_n N_VGND_c_628_n 0.0127075f $X=4.255 $Y=0.73 $X2=0 $Y2=0
cc_302 N_A_c_378_n N_VGND_c_628_n 0.00466416f $X=4.18 $Y=0.73 $X2=0 $Y2=0
cc_303 A N_VGND_c_628_n 0.0244748f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_304 N_A_c_373_n N_VGND_c_631_n 0.00549284f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_305 N_A_c_374_n N_VGND_c_631_n 0.00146271f $X=4.18 $Y=0.805 $X2=0 $Y2=0
cc_306 N_A_c_376_n N_VGND_c_631_n 0.00486043f $X=4.255 $Y=0.73 $X2=0 $Y2=0
cc_307 N_A_c_373_n N_VGND_c_633_n 0.0100905f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_308 N_A_c_374_n N_VGND_c_633_n 0.00195537f $X=4.18 $Y=0.805 $X2=0 $Y2=0
cc_309 N_A_c_376_n N_VGND_c_633_n 0.0045595f $X=4.255 $Y=0.73 $X2=0 $Y2=0
cc_310 A N_VGND_c_633_n 0.0145667f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_311 N_D_N_M1006_g N_VPWR_c_459_n 0.00319461f $X=4.875 $Y=2.545 $X2=0 $Y2=0
cc_312 N_D_N_M1006_g N_VPWR_c_461_n 0.0086001f $X=4.875 $Y=2.545 $X2=0 $Y2=0
cc_313 N_D_N_M1006_g N_VPWR_c_457_n 0.0165291f $X=4.875 $Y=2.545 $X2=0 $Y2=0
cc_314 N_D_N_M1015_g N_VGND_c_628_n 0.00876879f $X=4.825 $Y=0.445 $X2=0 $Y2=0
cc_315 N_D_N_M1015_g N_VGND_c_632_n 0.00585385f $X=4.825 $Y=0.445 $X2=0 $Y2=0
cc_316 N_D_N_M1017_g N_VGND_c_632_n 0.00549284f $X=5.215 $Y=0.445 $X2=0 $Y2=0
cc_317 N_D_N_M1015_g N_VGND_c_633_n 0.00989822f $X=4.825 $Y=0.445 $X2=0 $Y2=0
cc_318 N_D_N_M1017_g N_VGND_c_633_n 0.00972717f $X=5.215 $Y=0.445 $X2=0 $Y2=0
cc_319 N_D_N_c_429_n N_VGND_c_633_n 0.0114645f $X=5.02 $Y=0.99 $X2=0 $Y2=0
cc_320 N_VPWR_c_458_n N_A_245_409#_c_499_n 0.0229861f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_458_n N_A_245_409#_c_500_n 0.0478334f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_460_n N_A_245_409#_c_500_n 0.0220321f $X=4.405 $Y=3.33 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_457_n N_A_245_409#_c_500_n 0.0125808f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_460_n N_A_352_409#_c_533_n 0.079983f $X=4.405 $Y=3.33 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_457_n N_A_352_409#_c_533_n 0.0493242f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_460_n N_A_352_409#_c_534_n 0.021757f $X=4.405 $Y=3.33 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_457_n N_A_352_409#_c_534_n 0.0125691f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_460_n N_A_352_409#_c_535_n 0.0221635f $X=4.405 $Y=3.33 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_457_n N_A_352_409#_c_535_n 0.0126536f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_A_245_409#_c_501_n N_A_352_409#_M1016_d 0.006983f $X=2.825 $Y=2.27
+ $X2=-0.19 $Y2=1.655
cc_331 N_A_245_409#_c_500_n N_A_352_409#_c_532_n 0.0236877f $X=1.37 $Y=2.9 $X2=0
+ $Y2=0
cc_332 N_A_245_409#_c_501_n N_A_352_409#_c_532_n 0.0206372f $X=2.825 $Y=2.27
+ $X2=0 $Y2=0
cc_333 N_A_245_409#_c_501_n N_A_352_409#_c_533_n 0.0236107f $X=2.825 $Y=2.27
+ $X2=0 $Y2=0
cc_334 N_A_245_409#_c_502_n N_A_352_409#_c_533_n 0.0247135f $X=2.99 $Y=2.19
+ $X2=0 $Y2=0
cc_335 N_A_245_409#_c_500_n N_A_352_409#_c_534_n 0.0119061f $X=1.37 $Y=2.9 $X2=0
+ $Y2=0
cc_336 N_A_245_409#_c_502_n N_A_352_409#_c_536_n 0.047223f $X=2.99 $Y=2.19 $X2=0
+ $Y2=0
cc_337 N_A_245_409#_c_501_n N_Y_M1000_s 0.00773144f $X=2.825 $Y=2.27 $X2=0 $Y2=0
cc_338 N_A_245_409#_c_501_n N_Y_c_563_n 0.021375f $X=2.825 $Y=2.27 $X2=0 $Y2=0
cc_339 N_A_245_409#_c_501_n N_Y_c_565_n 0.0342666f $X=2.825 $Y=2.27 $X2=0 $Y2=0
cc_340 N_Y_c_560_n N_VGND_c_627_n 0.0205453f $X=3.455 $Y=0.9 $X2=0 $Y2=0
cc_341 N_Y_c_561_n N_VGND_c_627_n 0.0130164f $X=1.92 $Y=0.985 $X2=0 $Y2=0
cc_342 N_Y_c_602_n N_VGND_c_628_n 0.0114276f $X=3.62 $Y=0.47 $X2=0 $Y2=0
cc_343 N_Y_c_561_n N_VGND_c_630_n 0.034298f $X=1.92 $Y=0.985 $X2=0 $Y2=0
cc_344 N_Y_c_602_n N_VGND_c_631_n 0.0179149f $X=3.62 $Y=0.47 $X2=0 $Y2=0
cc_345 N_Y_M1009_d N_VGND_c_633_n 0.0022543f $X=1.87 $Y=0.235 $X2=0 $Y2=0
cc_346 N_Y_M1004_d N_VGND_c_633_n 0.0022543f $X=3.48 $Y=0.235 $X2=0 $Y2=0
cc_347 N_Y_c_560_n N_VGND_c_633_n 0.027296f $X=3.455 $Y=0.9 $X2=0 $Y2=0
cc_348 N_Y_c_602_n N_VGND_c_633_n 0.0124902f $X=3.62 $Y=0.47 $X2=0 $Y2=0
cc_349 N_Y_c_561_n N_VGND_c_633_n 0.0260422f $X=1.92 $Y=0.985 $X2=0 $Y2=0
cc_350 N_Y_c_561_n A_302_47# 9.59731e-19 $X=1.92 $Y=0.985 $X2=-0.19 $Y2=-0.245
cc_351 A_144_47# N_VGND_c_633_n 0.00303453f $X=0.72 $Y=0.235 $X2=5.52 $Y2=0
cc_352 N_VGND_c_633_n A_302_47# 0.00360352f $X=5.52 $Y=0 $X2=-0.19 $Y2=-0.245
cc_353 N_VGND_c_633_n A_460_47# 0.00300307f $X=5.52 $Y=0 $X2=-0.19 $Y2=-0.245
cc_354 N_VGND_c_633_n A_624_47# 0.00300307f $X=5.52 $Y=0 $X2=-0.19 $Y2=-0.245
cc_355 N_VGND_c_633_n A_782_47# 0.00546239f $X=5.52 $Y=0 $X2=-0.19 $Y2=-0.245
cc_356 N_VGND_c_633_n A_980_47# 0.00346444f $X=5.52 $Y=0 $X2=-0.19 $Y2=-0.245
