# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__srsdfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.590000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.475000 0.265000 13.835000 1.145000 ;
        RECT 13.475000 1.815000 13.835000 3.075000 ;
        RECT 13.665000 1.145000 13.835000 1.815000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.750000 2.490000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.985000 1.965000 1.010000 ;
        RECT 0.425000 1.010000 0.755000 1.315000 ;
        RECT 0.585000 0.840000 1.965000 0.985000 ;
        RECT 1.795000 1.010000 1.965000 1.180000 ;
        RECT 1.795000 1.180000 2.275000 1.510000 ;
    END
  END SCE
  PIN SLEEP_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.805000 0.255000 11.850000 0.425000 ;
        RECT  9.805000 0.425000 10.135000 0.575000 ;
        RECT 11.520000 0.425000 11.850000 0.650000 ;
    END
  END SLEEP_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 9.725000 1.500000 11.010000 1.830000 ;
    END
  END CLK
  PIN KAPWR
    ANTENNADIFFAREA  0.710800 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 13.850000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.085000  0.255000  0.415000 0.675000 ;
      RECT  0.085000  0.675000  0.255000 1.910000 ;
      RECT  0.085000  1.910000  1.905000 2.080000 ;
      RECT  0.085000  2.080000  0.385000 3.045000 ;
      RECT  0.565000  2.365000  0.895000 3.245000 ;
      RECT  0.585000  1.555000  0.915000 1.750000 ;
      RECT  0.585000  1.750000  1.905000 1.910000 ;
      RECT  0.595000  0.085000  0.925000 0.670000 ;
      RECT  1.385000  2.320000  2.990000 2.490000 ;
      RECT  1.385000  2.490000  1.715000 3.045000 ;
      RECT  1.525000  0.255000  1.855000 0.500000 ;
      RECT  1.525000  0.500000  2.305000 0.670000 ;
      RECT  2.135000  0.670000  2.305000 0.840000 ;
      RECT  2.135000  0.840000  2.655000 1.010000 ;
      RECT  2.400000  2.660000  2.650000 3.245000 ;
      RECT  2.475000  0.085000  2.645000 0.670000 ;
      RECT  2.485000  1.010000  2.830000 1.180000 ;
      RECT  2.660000  1.180000  2.830000 2.320000 ;
      RECT  2.820000  2.490000  2.990000 2.905000 ;
      RECT  2.820000  2.905000  4.425000 3.075000 ;
      RECT  2.825000  0.255000  4.575000 0.425000 ;
      RECT  2.825000  0.425000  3.570000 0.585000 ;
      RECT  2.825000  0.585000  3.170000 0.675000 ;
      RECT  3.000000  0.675000  3.170000 1.980000 ;
      RECT  3.000000  1.980000  3.455000 2.150000 ;
      RECT  3.205000  2.150000  3.455000 2.405000 ;
      RECT  3.205000  2.405000  3.925000 2.735000 ;
      RECT  3.475000  0.755000  3.805000 1.135000 ;
      RECT  3.635000  1.135000  3.805000 2.065000 ;
      RECT  3.635000  2.065000  4.425000 2.235000 ;
      RECT  3.985000  0.675000  4.235000 1.725000 ;
      RECT  3.985000  1.725000  5.440000 1.895000 ;
      RECT  4.095000  2.235000  4.425000 2.905000 ;
      RECT  4.405000  0.425000  4.575000 0.615000 ;
      RECT  4.405000  0.615000  5.440000 0.785000 ;
      RECT  4.570000  0.955000  5.780000 1.125000 ;
      RECT  4.570000  1.125000  4.900000 1.555000 ;
      RECT  4.595000  1.895000  4.925000 2.625000 ;
      RECT  4.595000  2.625000  6.165000 2.795000 ;
      RECT  4.595000  2.795000  4.925000 3.075000 ;
      RECT  4.805000  0.085000  5.055000 0.445000 ;
      RECT  5.110000  1.295000  5.440000 1.725000 ;
      RECT  5.270000  0.255000  7.780000 0.425000 ;
      RECT  5.270000  0.425000  5.440000 0.615000 ;
      RECT  5.290000  2.105000  6.665000 2.455000 ;
      RECT  5.495000  2.965000  5.825000 3.245000 ;
      RECT  5.610000  0.595000  5.780000 0.955000 ;
      RECT  5.610000  1.125000  5.780000 2.105000 ;
      RECT  5.950000  0.425000  6.120000 1.095000 ;
      RECT  5.950000  1.095000  6.540000 1.425000 ;
      RECT  5.995000  2.795000  6.165000 2.905000 ;
      RECT  5.995000  2.905000  8.340000 3.075000 ;
      RECT  6.335000  2.455000  6.665000 2.735000 ;
      RECT  6.880000  0.595000  7.210000 0.925000 ;
      RECT  7.040000  0.925000  7.210000 1.425000 ;
      RECT  7.040000  1.425000  8.880000 1.595000 ;
      RECT  7.195000  1.595000  7.525000 2.265000 ;
      RECT  7.195000  2.265000  9.065000 2.340000 ;
      RECT  7.195000  2.340000 10.345000 2.435000 ;
      RECT  7.195000  2.435000  7.525000 2.735000 ;
      RECT  7.380000  0.425000  7.780000 1.085000 ;
      RECT  7.380000  1.085000  9.420000 1.255000 ;
      RECT  7.950000  0.085000  8.280000 0.915000 ;
      RECT  8.010000  1.765000  8.340000 1.925000 ;
      RECT  8.010000  1.925000  9.405000 2.000000 ;
      RECT  8.010000  2.000000 11.350000 2.095000 ;
      RECT  8.010000  2.745000  8.340000 2.905000 ;
      RECT  8.550000  1.595000  8.880000 1.755000 ;
      RECT  8.735000  2.435000 10.345000 2.510000 ;
      RECT  8.735000  2.510000  9.065000 3.075000 ;
      RECT  8.970000  0.585000  9.300000 0.745000 ;
      RECT  8.970000  0.745000 11.315000 0.765000 ;
      RECT  8.970000  0.765000 10.475000 0.915000 ;
      RECT  9.090000  1.255000  9.420000 1.725000 ;
      RECT  9.235000  2.095000 11.350000 2.170000 ;
      RECT  9.590000  0.915000  9.920000 1.120000 ;
      RECT  9.725000  2.680000 10.005000 3.075000 ;
      RECT 10.175000  2.510000 10.345000 2.905000 ;
      RECT 10.175000  2.905000 11.025000 3.075000 ;
      RECT 10.305000  0.595000 11.315000 0.745000 ;
      RECT 10.515000  2.170000 10.685000 2.735000 ;
      RECT 10.645000  0.935000 10.975000 1.160000 ;
      RECT 10.645000  1.160000 11.350000 1.330000 ;
      RECT 10.855000  2.340000 11.705000 2.510000 ;
      RECT 10.855000  2.510000 11.025000 2.905000 ;
      RECT 11.145000  0.765000 11.315000 0.820000 ;
      RECT 11.145000  0.820000 11.690000 0.990000 ;
      RECT 11.180000  1.330000 11.350000 2.000000 ;
      RECT 11.195000  2.680000 11.365000 3.075000 ;
      RECT 11.520000  0.990000 11.690000 2.000000 ;
      RECT 11.520000  2.000000 12.125000 2.170000 ;
      RECT 11.535000  2.510000 11.705000 2.745000 ;
      RECT 11.535000  2.745000 12.595000 3.075000 ;
      RECT 11.875000  2.170000 12.125000 2.575000 ;
      RECT 12.020000  0.085000 12.270000 1.330000 ;
      RECT 12.500000  0.265000 12.830000 1.315000 ;
      RECT 12.500000  1.315000 13.495000 1.645000 ;
      RECT 12.500000  1.645000 12.830000 2.495000 ;
      RECT 13.045000  0.085000 13.295000 1.145000 ;
      RECT 13.045000  1.815000 13.295000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  2.735000  9.925000 2.905000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  2.735000 11.365000 2.905000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_lp__srsdfxtp_1
