* File: sky130_fd_sc_lp__or2_lp2.pxi.spice
* Created: Fri Aug 28 11:21:44 2020
* 
x_PM_SKY130_FD_SC_LP__OR2_LP2%B N_B_c_49_n N_B_M1007_g N_B_c_55_n N_B_c_56_n
+ N_B_M1008_g N_B_c_58_n N_B_M1001_g N_B_c_59_n B B B B B N_B_c_53_n
+ PM_SKY130_FD_SC_LP__OR2_LP2%B
x_PM_SKY130_FD_SC_LP__OR2_LP2%A N_A_M1002_g N_A_M1005_g N_A_M1000_g N_A_c_96_n
+ N_A_c_97_n A N_A_c_98_n N_A_c_99_n PM_SKY130_FD_SC_LP__OR2_LP2%A
x_PM_SKY130_FD_SC_LP__OR2_LP2%A_226_409# N_A_226_409#_M1008_d
+ N_A_226_409#_M1001_s N_A_226_409#_M1003_g N_A_226_409#_M1006_g
+ N_A_226_409#_M1004_g N_A_226_409#_c_140_n N_A_226_409#_c_146_n
+ N_A_226_409#_c_147_n N_A_226_409#_c_141_n N_A_226_409#_c_142_n
+ N_A_226_409#_c_143_n N_A_226_409#_c_149_n
+ PM_SKY130_FD_SC_LP__OR2_LP2%A_226_409#
x_PM_SKY130_FD_SC_LP__OR2_LP2%VPWR N_VPWR_M1005_d N_VPWR_c_210_n VPWR
+ N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_209_n N_VPWR_c_214_n
+ PM_SKY130_FD_SC_LP__OR2_LP2%VPWR
x_PM_SKY130_FD_SC_LP__OR2_LP2%X N_X_M1004_d N_X_M1006_d X X X X X X X
+ PM_SKY130_FD_SC_LP__OR2_LP2%X
x_PM_SKY130_FD_SC_LP__OR2_LP2%VGND N_VGND_M1007_s N_VGND_M1000_d N_VGND_c_247_n
+ N_VGND_c_248_n VGND N_VGND_c_249_n N_VGND_c_250_n N_VGND_c_251_n
+ N_VGND_c_252_n N_VGND_c_253_n N_VGND_c_254_n PM_SKY130_FD_SC_LP__OR2_LP2%VGND
cc_1 VNB N_B_c_49_n 0.024217f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.7
cc_2 VNB N_B_M1007_g 0.0492118f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.495
cc_3 VNB N_B_M1008_g 0.0582257f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=0.495
cc_4 VNB B 0.0443091f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_B_c_53_n 0.0208209f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.345
cc_6 VNB N_A_M1002_g 0.0202463f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.18
cc_7 VNB N_A_M1000_g 0.0199512f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=0.495
cc_8 VNB N_A_c_96_n 0.0188696f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.837
cc_9 VNB N_A_c_97_n 0.0200708f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A_c_98_n 0.0236468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_99_n 0.0148227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_226_409#_M1003_g 0.0352042f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.7
cc_13 VNB N_A_226_409#_M1004_g 0.0431902f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.837
cc_14 VNB N_A_226_409#_c_140_n 0.00742849f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_15 VNB N_A_226_409#_c_141_n 0.00158268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_226_409#_c_142_n 0.0472655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_226_409#_c_143_n 0.0122165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_209_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB X 0.0587996f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.775
cc_20 VNB N_VGND_c_247_n 0.0256276f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.7
cc_21 VNB N_VGND_c_248_n 0.0124633f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.975
cc_22 VNB N_VGND_c_249_n 0.0182134f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.837
cc_23 VNB N_VGND_c_250_n 0.0342115f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.69
cc_24 VNB N_VGND_c_251_n 0.0275168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_252_n 0.233447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_253_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_254_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_B_c_49_n 0.00362432f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.7
cc_29 VPB N_B_c_55_n 0.0168983f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.775
cc_30 VPB N_B_c_56_n 0.0211155f $X=-0.19 $Y=1.655 $X2=0.96 $Y2=1.775
cc_31 VPB N_B_M1008_g 0.00243952f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=0.495
cc_32 VPB N_B_c_58_n 0.0233468f $X=-0.19 $Y=1.655 $X2=1.54 $Y2=1.975
cc_33 VPB N_B_c_59_n 0.0375091f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.837
cc_34 VPB B 0.095633f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_35 VPB N_A_M1005_g 0.0376391f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.775
cc_36 VPB N_A_c_97_n 0.00326474f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_37 VPB N_A_226_409#_M1006_g 0.0324079f $X=-0.19 $Y=1.655 $X2=1.54 $Y2=1.975
cc_38 VPB N_A_226_409#_c_140_n 2.72658e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_39 VPB N_A_226_409#_c_146_n 0.0187707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_226_409#_c_147_n 0.031218f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_226_409#_c_142_n 0.0310915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_226_409#_c_149_n 7.18167e-19 $X=-0.19 $Y=1.655 $X2=0.765 $Y2=1.345
cc_43 VPB N_VPWR_c_210_n 0.00423941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_211_n 0.0609238f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=0.495
cc_45 VPB N_VPWR_c_212_n 0.0277571f $X=-0.19 $Y=1.655 $X2=1.54 $Y2=1.837
cc_46 VPB N_VPWR_c_209_n 0.0846194f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_47 VPB N_VPWR_c_214_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_48 VPB X 0.0573842f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.775
cc_49 N_B_M1008_g N_A_M1002_g 0.022993f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_50 N_B_c_59_n N_A_M1005_g 0.0794349f $X=1.275 $Y=1.837 $X2=0 $Y2=0
cc_51 N_B_M1008_g N_A_c_97_n 0.00286218f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_52 N_B_M1008_g N_A_c_98_n 0.0103846f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_53 N_B_M1008_g N_A_c_99_n 0.00574589f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_54 N_B_c_59_n N_A_c_99_n 6.11703e-19 $X=1.275 $Y=1.837 $X2=0 $Y2=0
cc_55 N_B_M1007_g N_A_226_409#_c_140_n 0.0125991f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_56 N_B_c_55_n N_A_226_409#_c_140_n 0.00120871f $X=1.2 $Y=1.775 $X2=0 $Y2=0
cc_57 N_B_M1008_g N_A_226_409#_c_140_n 0.0233567f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_58 N_B_c_59_n N_A_226_409#_c_140_n 0.00141685f $X=1.275 $Y=1.837 $X2=0 $Y2=0
cc_59 B N_A_226_409#_c_140_n 0.0434897f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_B_c_58_n N_A_226_409#_c_146_n 0.023356f $X=1.54 $Y=1.975 $X2=0 $Y2=0
cc_61 N_B_c_59_n N_A_226_409#_c_146_n 0.00195687f $X=1.275 $Y=1.837 $X2=0 $Y2=0
cc_62 B N_A_226_409#_c_146_n 0.0816127f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_B_c_59_n N_A_226_409#_c_147_n 0.020861f $X=1.275 $Y=1.837 $X2=0 $Y2=0
cc_64 N_B_M1007_g N_A_226_409#_c_143_n 0.00349982f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_65 N_B_M1008_g N_A_226_409#_c_143_n 0.0143981f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_66 N_B_c_55_n N_A_226_409#_c_149_n 0.00445197f $X=1.2 $Y=1.775 $X2=0 $Y2=0
cc_67 N_B_c_59_n N_A_226_409#_c_149_n 0.0167516f $X=1.275 $Y=1.837 $X2=0 $Y2=0
cc_68 B N_A_226_409#_c_149_n 0.0143628f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_B_c_58_n N_VPWR_c_210_n 0.00484657f $X=1.54 $Y=1.975 $X2=0 $Y2=0
cc_70 N_B_c_58_n N_VPWR_c_211_n 0.0086001f $X=1.54 $Y=1.975 $X2=0 $Y2=0
cc_71 B N_VPWR_c_211_n 0.0262577f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_B_c_58_n N_VPWR_c_209_n 0.0166232f $X=1.54 $Y=1.975 $X2=0 $Y2=0
cc_73 B N_VPWR_c_209_n 0.0279979f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B_M1007_g N_VGND_c_247_n 0.0126777f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_75 N_B_M1008_g N_VGND_c_247_n 0.00126144f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_76 B N_VGND_c_247_n 0.0142766f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_B_c_53_n N_VGND_c_247_n 0.00142984f $X=0.765 $Y=1.345 $X2=0 $Y2=0
cc_78 N_B_M1007_g N_VGND_c_250_n 0.00445056f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_79 N_B_M1008_g N_VGND_c_250_n 0.00327726f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_80 N_B_M1007_g N_VGND_c_252_n 0.00802306f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_81 N_B_M1008_g N_VGND_c_252_n 0.00481302f $X=1.275 $Y=0.495 $X2=0 $Y2=0
cc_82 N_A_M1000_g N_A_226_409#_M1003_g 0.0301347f $X=2.065 $Y=0.495 $X2=0 $Y2=0
cc_83 N_A_c_99_n N_A_226_409#_M1003_g 0.00191919f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_84 N_A_M1005_g N_A_226_409#_M1006_g 0.017721f $X=2.03 $Y=2.545 $X2=0 $Y2=0
cc_85 N_A_M1002_g N_A_226_409#_c_140_n 9.88678e-19 $X=1.705 $Y=0.495 $X2=0 $Y2=0
cc_86 N_A_c_97_n N_A_226_409#_c_140_n 8.29939e-19 $X=1.975 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_98_n N_A_226_409#_c_140_n 4.37796e-19 $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_88 N_A_c_99_n N_A_226_409#_c_140_n 0.0361877f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_89 N_A_M1005_g N_A_226_409#_c_146_n 0.0049233f $X=2.03 $Y=2.545 $X2=0 $Y2=0
cc_90 N_A_M1005_g N_A_226_409#_c_147_n 0.0222664f $X=2.03 $Y=2.545 $X2=0 $Y2=0
cc_91 N_A_c_97_n N_A_226_409#_c_147_n 0.00247487f $X=1.975 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_99_n N_A_226_409#_c_147_n 0.0439839f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_93 N_A_c_97_n N_A_226_409#_c_141_n 0.001216f $X=1.975 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_98_n N_A_226_409#_c_141_n 4.59979e-19 $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_95 N_A_c_99_n N_A_226_409#_c_141_n 0.0203894f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_96 N_A_c_97_n N_A_226_409#_c_142_n 0.0179764f $X=1.975 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_98_n N_A_226_409#_c_142_n 0.0184735f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_98 N_A_c_99_n N_A_226_409#_c_142_n 0.00148106f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_99 N_A_M1002_g N_A_226_409#_c_143_n 0.00867914f $X=1.705 $Y=0.495 $X2=0 $Y2=0
cc_100 N_A_M1000_g N_A_226_409#_c_143_n 0.0012437f $X=2.065 $Y=0.495 $X2=0 $Y2=0
cc_101 N_A_c_99_n N_A_226_409#_c_143_n 0.00756724f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_102 N_A_M1005_g N_VPWR_c_210_n 0.0276765f $X=2.03 $Y=2.545 $X2=0 $Y2=0
cc_103 N_A_M1005_g N_VPWR_c_211_n 0.00802402f $X=2.03 $Y=2.545 $X2=0 $Y2=0
cc_104 N_A_M1005_g N_VPWR_c_209_n 0.0142664f $X=2.03 $Y=2.545 $X2=0 $Y2=0
cc_105 N_A_M1002_g N_VGND_c_248_n 0.00211588f $X=1.705 $Y=0.495 $X2=0 $Y2=0
cc_106 N_A_M1000_g N_VGND_c_248_n 0.0125133f $X=2.065 $Y=0.495 $X2=0 $Y2=0
cc_107 N_A_c_99_n N_VGND_c_248_n 0.00192823f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_108 N_A_M1002_g N_VGND_c_250_n 0.00501304f $X=1.705 $Y=0.495 $X2=0 $Y2=0
cc_109 N_A_M1000_g N_VGND_c_250_n 0.00445056f $X=2.065 $Y=0.495 $X2=0 $Y2=0
cc_110 N_A_M1002_g N_VGND_c_252_n 0.00938372f $X=1.705 $Y=0.495 $X2=0 $Y2=0
cc_111 N_A_M1000_g N_VGND_c_252_n 0.00796275f $X=2.065 $Y=0.495 $X2=0 $Y2=0
cc_112 N_A_226_409#_M1006_g N_VPWR_c_210_n 0.0129585f $X=2.805 $Y=2.545 $X2=0
+ $Y2=0
cc_113 N_A_226_409#_c_147_n N_VPWR_c_210_n 0.0239129f $X=2.395 $Y=1.84 $X2=0
+ $Y2=0
cc_114 N_A_226_409#_c_142_n N_VPWR_c_210_n 4.4776e-19 $X=2.56 $Y=1.38 $X2=0
+ $Y2=0
cc_115 N_A_226_409#_c_146_n N_VPWR_c_211_n 0.0220321f $X=1.275 $Y=2.19 $X2=0
+ $Y2=0
cc_116 N_A_226_409#_M1006_g N_VPWR_c_212_n 0.0086001f $X=2.805 $Y=2.545 $X2=0
+ $Y2=0
cc_117 N_A_226_409#_M1006_g N_VPWR_c_209_n 0.0167763f $X=2.805 $Y=2.545 $X2=0
+ $Y2=0
cc_118 N_A_226_409#_c_146_n N_VPWR_c_209_n 0.0125808f $X=1.275 $Y=2.19 $X2=0
+ $Y2=0
cc_119 N_A_226_409#_M1003_g X 0.00370468f $X=2.495 $Y=0.495 $X2=0 $Y2=0
cc_120 N_A_226_409#_M1006_g X 0.0314276f $X=2.805 $Y=2.545 $X2=0 $Y2=0
cc_121 N_A_226_409#_M1004_g X 0.0273034f $X=2.855 $Y=0.495 $X2=0 $Y2=0
cc_122 N_A_226_409#_c_147_n X 0.0128825f $X=2.395 $Y=1.84 $X2=0 $Y2=0
cc_123 N_A_226_409#_c_141_n X 0.0386728f $X=2.56 $Y=1.38 $X2=0 $Y2=0
cc_124 N_A_226_409#_c_142_n X 0.024757f $X=2.56 $Y=1.38 $X2=0 $Y2=0
cc_125 N_A_226_409#_c_143_n N_VGND_c_247_n 0.025737f $X=1.49 $Y=0.495 $X2=0
+ $Y2=0
cc_126 N_A_226_409#_M1003_g N_VGND_c_248_n 0.0128002f $X=2.495 $Y=0.495 $X2=0
+ $Y2=0
cc_127 N_A_226_409#_M1004_g N_VGND_c_248_n 0.002112f $X=2.855 $Y=0.495 $X2=0
+ $Y2=0
cc_128 N_A_226_409#_c_141_n N_VGND_c_248_n 0.00182217f $X=2.56 $Y=1.38 $X2=0
+ $Y2=0
cc_129 N_A_226_409#_c_143_n N_VGND_c_248_n 0.0159687f $X=1.49 $Y=0.495 $X2=0
+ $Y2=0
cc_130 N_A_226_409#_c_143_n N_VGND_c_250_n 0.0348952f $X=1.49 $Y=0.495 $X2=0
+ $Y2=0
cc_131 N_A_226_409#_M1003_g N_VGND_c_251_n 0.00445056f $X=2.495 $Y=0.495 $X2=0
+ $Y2=0
cc_132 N_A_226_409#_M1004_g N_VGND_c_251_n 0.00502664f $X=2.855 $Y=0.495 $X2=0
+ $Y2=0
cc_133 N_A_226_409#_M1003_g N_VGND_c_252_n 0.00796275f $X=2.495 $Y=0.495 $X2=0
+ $Y2=0
cc_134 N_A_226_409#_M1004_g N_VGND_c_252_n 0.0100677f $X=2.855 $Y=0.495 $X2=0
+ $Y2=0
cc_135 N_A_226_409#_c_143_n N_VGND_c_252_n 0.0200515f $X=1.49 $Y=0.495 $X2=0
+ $Y2=0
cc_136 N_A_226_409#_c_143_n A_192_57# 0.0043889f $X=1.49 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_137 N_VPWR_c_210_n X 0.035459f $X=2.295 $Y=2.27 $X2=0 $Y2=0
cc_138 N_VPWR_c_212_n X 0.0220321f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_139 N_VPWR_c_209_n X 0.0125808f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_140 X N_VGND_c_248_n 0.0153904f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_141 X N_VGND_c_251_n 0.0220321f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_142 X N_VGND_c_252_n 0.0125808f $X=3.035 $Y=0.47 $X2=0 $Y2=0
