# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.810000 1.820000 1.820000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.315000 0.265000 17.670000 1.125000 ;
        RECT 17.315000 1.815000 17.670000 3.065000 ;
        RECT 17.500000 1.125000 17.670000 1.815000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.592200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.850000 0.265000 16.255000 1.145000 ;
        RECT 15.900000 1.835000 16.255000 3.065000 ;
        RECT 16.085000 1.145000 16.255000 1.835000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.005000 1.345000 15.365000 1.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.215000 0.550000 1.885000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.850000 1.215000 1.310000 1.780000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  8.735000 1.180000  9.025000 1.225000 ;
        RECT  8.735000 1.225000 13.345000 1.365000 ;
        RECT  8.735000 1.365000  9.025000 1.410000 ;
        RECT 13.055000 1.180000 13.345000 1.225000 ;
        RECT 13.055000 1.365000 13.345000 1.410000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.860000 0.870000 4.195000 1.540000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 17.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 17.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.760000 0.085000 ;
      RECT  0.000000  3.245000 17.760000 3.415000 ;
      RECT  0.115000  2.065000  1.145000 2.235000 ;
      RECT  0.115000  2.235000  0.365000 3.030000 ;
      RECT  0.155000  0.085000  0.485000 1.035000 ;
      RECT  0.545000  2.415000  0.795000 3.245000 ;
      RECT  0.975000  2.235000  1.145000 2.895000 ;
      RECT  0.975000  2.895000  2.095000 3.065000 ;
      RECT  0.980000  0.460000  2.170000 0.630000 ;
      RECT  0.980000  0.630000  1.310000 1.035000 ;
      RECT  1.335000  2.000000  2.170000 2.170000 ;
      RECT  1.335000  2.170000  1.585000 2.715000 ;
      RECT  1.765000  2.350000  2.095000 2.895000 ;
      RECT  2.000000  0.630000  2.170000 1.685000 ;
      RECT  2.000000  1.685000  2.915000 1.855000 ;
      RECT  2.000000  1.855000  2.170000 2.000000 ;
      RECT  2.350000  0.085000  2.680000 0.995000 ;
      RECT  2.350000  1.175000  3.265000 1.505000 ;
      RECT  2.395000  2.035000  2.565000 3.245000 ;
      RECT  2.745000  1.855000  2.915000 2.895000 ;
      RECT  2.745000  2.895000  3.615000 3.065000 ;
      RECT  3.095000  0.575000  3.425000 1.035000 ;
      RECT  3.095000  1.035000  3.265000 1.175000 ;
      RECT  3.095000  1.505000  3.265000 2.715000 ;
      RECT  3.445000  1.720000  4.315000 1.890000 ;
      RECT  3.445000  1.890000  3.615000 2.895000 ;
      RECT  3.655000  0.085000  3.985000 0.690000 ;
      RECT  3.795000  2.070000  3.965000 3.245000 ;
      RECT  4.145000  1.890000  4.315000 2.895000 ;
      RECT  4.145000  2.895000  5.290000 3.065000 ;
      RECT  4.165000  0.265000  4.545000 0.690000 ;
      RECT  4.375000  0.690000  4.545000 0.870000 ;
      RECT  4.375000  0.870000  4.760000 1.540000 ;
      RECT  4.495000  1.540000  4.760000 2.715000 ;
      RECT  4.955000  0.310000  5.285000 1.345000 ;
      RECT  4.955000  1.345000  6.000000 1.675000 ;
      RECT  4.955000  1.675000  5.295000 2.145000 ;
      RECT  5.120000  2.325000  6.350000 2.495000 ;
      RECT  5.120000  2.495000  5.290000 2.895000 ;
      RECT  5.465000  0.085000  5.795000 0.770000 ;
      RECT  5.470000  2.675000  5.800000 3.245000 ;
      RECT  6.020000  1.875000  6.350000 2.325000 ;
      RECT  6.025000  0.605000  6.355000 1.065000 ;
      RECT  6.180000  1.065000  6.350000 1.875000 ;
      RECT  6.530000  1.875000  7.660000 2.045000 ;
      RECT  6.530000  2.045000  6.865000 2.335000 ;
      RECT  6.535000  0.500000  6.865000 1.875000 ;
      RECT  7.045000  0.705000  8.555000 0.875000 ;
      RECT  7.045000  0.875000  7.310000 1.380000 ;
      RECT  7.490000  1.055000  8.390000 1.225000 ;
      RECT  7.490000  1.225000  7.660000 1.875000 ;
      RECT  7.840000  1.405000  8.040000 1.940000 ;
      RECT  7.840000  1.940000  9.855000 2.110000 ;
      RECT  7.875000  0.085000  8.205000 0.525000 ;
      RECT  8.220000  1.225000  8.390000 1.590000 ;
      RECT  8.220000  1.590000  9.505000 1.735000 ;
      RECT  8.220000  1.735000  9.345000 1.760000 ;
      RECT  8.300000  2.290000  8.630000 3.245000 ;
      RECT  8.385000  0.265000 10.435000 0.435000 ;
      RECT  8.385000  0.435000  8.555000 0.705000 ;
      RECT  8.570000  1.080000  8.995000 1.410000 ;
      RECT  8.735000  0.615000 10.085000 0.785000 ;
      RECT  8.735000  0.785000  9.065000 0.900000 ;
      RECT  9.175000  1.405000  9.505000 1.590000 ;
      RECT  9.245000  0.965000  9.575000 1.055000 ;
      RECT  9.245000  1.055000  9.855000 1.225000 ;
      RECT  9.525000  1.915000  9.855000 1.940000 ;
      RECT  9.525000  2.110000  9.855000 2.755000 ;
      RECT  9.685000  1.225000  9.855000 1.435000 ;
      RECT  9.685000  1.435000 10.940000 1.725000 ;
      RECT  9.685000  1.725000  9.855000 1.915000 ;
      RECT  9.755000  0.785000 10.085000 0.875000 ;
      RECT 10.265000  0.435000 10.435000 1.085000 ;
      RECT 10.265000  1.085000 11.290000 1.255000 ;
      RECT 10.345000  1.905000 10.675000 3.245000 ;
      RECT 10.615000  0.085000 10.865000 0.905000 ;
      RECT 11.120000  1.255000 11.290000 1.345000 ;
      RECT 11.120000  1.345000 11.530000 1.675000 ;
      RECT 11.120000  1.675000 11.290000 2.895000 ;
      RECT 11.120000  2.895000 12.430000 3.065000 ;
      RECT 11.470000  0.575000 11.880000 0.830000 ;
      RECT 11.470000  0.830000 13.710000 1.000000 ;
      RECT 11.470000  1.000000 11.880000 1.165000 ;
      RECT 11.470000  2.120000 11.880000 2.715000 ;
      RECT 11.710000  1.165000 11.880000 2.120000 ;
      RECT 12.100000  1.700000 12.430000 2.895000 ;
      RECT 12.640000  1.960000 13.865000 2.290000 ;
      RECT 12.645000  0.085000 12.975000 0.650000 ;
      RECT 13.000000  1.180000 13.330000 1.780000 ;
      RECT 13.105000  2.470000 13.355000 3.245000 ;
      RECT 13.235000  0.265000 14.665000 0.435000 ;
      RECT 13.235000  0.435000 13.565000 0.650000 ;
      RECT 13.535000  2.290000 13.865000 2.470000 ;
      RECT 13.535000  2.470000 15.720000 2.640000 ;
      RECT 13.535000  2.640000 13.865000 3.065000 ;
      RECT 13.540000  1.000000 13.710000 1.435000 ;
      RECT 13.540000  1.435000 13.870000 1.765000 ;
      RECT 13.905000  0.615000 14.155000 1.085000 ;
      RECT 13.905000  1.085000 14.220000 1.255000 ;
      RECT 14.050000  1.255000 14.220000 2.470000 ;
      RECT 14.325000  2.820000 14.655000 3.245000 ;
      RECT 14.335000  0.435000 14.665000 0.815000 ;
      RECT 14.400000  0.995000 15.240000 1.165000 ;
      RECT 14.400000  1.165000 14.730000 1.960000 ;
      RECT 14.400000  1.960000 15.210000 2.290000 ;
      RECT 14.910000  0.265000 15.240000 0.995000 ;
      RECT 15.390000  2.820000 15.720000 3.245000 ;
      RECT 15.420000  0.085000 15.670000 1.145000 ;
      RECT 15.550000  1.325000 15.905000 1.655000 ;
      RECT 15.550000  1.655000 15.720000 2.470000 ;
      RECT 16.455000  0.265000 16.660000 1.305000 ;
      RECT 16.455000  1.305000 17.320000 1.635000 ;
      RECT 16.455000  1.635000 16.705000 2.495000 ;
      RECT 16.840000  0.085000 17.090000 0.725000 ;
      RECT 16.885000  1.815000 17.135000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.210000  8.965000 1.380000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  1.210000 13.285000 1.380000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfbbn_1
END LIBRARY
