* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__iso0n_lp2 A SLEEP_B KAGND VGND VNB VPB VPWR X
X0 VPWR A a_65_65# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_65_65# A a_152_65# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_316_65# a_65_65# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_65_65# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 KAGND a_65_65# a_316_65# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_65_65# SLEEP_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_152_65# SLEEP_B KAGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
