* File: sky130_fd_sc_lp__sdfsbp_lp.pxi.spice
* Created: Wed Sep  2 10:35:29 2020
* 
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%SCE N_SCE_M1010_g N_SCE_M1023_g N_SCE_c_333_n
+ N_SCE_M1007_g N_SCE_M1032_g N_SCE_M1046_g N_SCE_c_335_n N_SCE_c_336_n
+ N_SCE_c_337_n N_SCE_c_338_n N_SCE_c_339_n N_SCE_c_340_n N_SCE_c_341_n
+ N_SCE_c_342_n N_SCE_c_343_n N_SCE_c_344_n N_SCE_c_351_n N_SCE_c_345_n SCE SCE
+ N_SCE_c_346_n N_SCE_c_347_n PM_SKY130_FD_SC_LP__SDFSBP_LP%SCE
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_27_409# N_A_27_409#_M1023_s
+ N_A_27_409#_M1010_s N_A_27_409#_M1045_g N_A_27_409#_c_440_n
+ N_A_27_409#_c_441_n N_A_27_409#_M1015_g N_A_27_409#_c_442_n
+ N_A_27_409#_c_443_n N_A_27_409#_c_444_n N_A_27_409#_c_445_n
+ N_A_27_409#_c_451_n N_A_27_409#_c_446_n N_A_27_409#_c_447_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%D N_D_M1031_g N_D_M1016_g D D N_D_c_509_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%D
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%SCD N_SCD_c_550_n N_SCD_M1033_g N_SCD_M1024_g
+ N_SCD_c_551_n SCD SCD N_SCD_c_553_n N_SCD_c_554_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%SCD
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%CLK N_CLK_M1042_g N_CLK_c_604_n N_CLK_M1047_g
+ N_CLK_M1006_g N_CLK_c_606_n CLK N_CLK_c_608_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%CLK
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_987_409# N_A_987_409#_M1039_d
+ N_A_987_409#_M1034_d N_A_987_409#_M1008_g N_A_987_409#_M1018_g
+ N_A_987_409#_M1022_g N_A_987_409#_M1035_g N_A_987_409#_c_671_n
+ N_A_987_409#_c_672_n N_A_987_409#_c_673_n N_A_987_409#_c_657_n
+ N_A_987_409#_c_674_n N_A_987_409#_c_658_n N_A_987_409#_c_659_n
+ N_A_987_409#_c_684_p N_A_987_409#_c_685_p N_A_987_409#_c_681_p
+ N_A_987_409#_c_686_p N_A_987_409#_c_660_n N_A_987_409#_c_661_n
+ N_A_987_409#_c_675_n N_A_987_409#_c_662_n N_A_987_409#_c_663_n
+ N_A_987_409#_c_664_n N_A_987_409#_c_665_n N_A_987_409#_c_695_p
+ N_A_987_409#_c_666_n N_A_987_409#_c_667_n N_A_987_409#_c_668_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_987_409#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_1423_99# N_A_1423_99#_M1001_s
+ N_A_1423_99#_M1026_d N_A_1423_99#_M1011_g N_A_1423_99#_M1004_g
+ N_A_1423_99#_c_869_n N_A_1423_99#_c_870_n N_A_1423_99#_c_871_n
+ N_A_1423_99#_c_872_n N_A_1423_99#_c_888_n N_A_1423_99#_c_878_n
+ N_A_1423_99#_c_873_n N_A_1423_99#_c_874_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_1423_99#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_1201_419# N_A_1201_419#_M1043_d
+ N_A_1201_419#_M1008_d N_A_1201_419#_M1026_g N_A_1201_419#_c_949_n
+ N_A_1201_419#_c_950_n N_A_1201_419#_c_951_n N_A_1201_419#_M1001_g
+ N_A_1201_419#_M1025_g N_A_1201_419#_M1002_g N_A_1201_419#_c_953_n
+ N_A_1201_419#_c_972_n N_A_1201_419#_c_992_n N_A_1201_419#_c_973_n
+ N_A_1201_419#_c_974_n N_A_1201_419#_c_1001_n N_A_1201_419#_c_954_n
+ N_A_1201_419#_c_955_n N_A_1201_419#_c_956_n N_A_1201_419#_c_957_n
+ N_A_1201_419#_c_958_n N_A_1201_419#_c_959_n N_A_1201_419#_c_960_n
+ N_A_1201_419#_c_961_n N_A_1201_419#_c_962_n N_A_1201_419#_c_963_n
+ N_A_1201_419#_c_964_n N_A_1201_419#_c_965_n N_A_1201_419#_c_1062_n
+ N_A_1201_419#_c_966_n N_A_1201_419#_c_967_n N_A_1201_419#_c_968_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_1201_419#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%SET_B N_SET_B_M1005_g N_SET_B_M1037_g
+ N_SET_B_c_1148_n N_SET_B_M1048_g N_SET_B_c_1149_n N_SET_B_c_1150_n
+ N_SET_B_M1027_g N_SET_B_c_1151_n N_SET_B_c_1152_n N_SET_B_c_1153_n SET_B
+ N_SET_B_c_1155_n N_SET_B_c_1156_n N_SET_B_c_1157_n N_SET_B_c_1158_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%SET_B
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_761_113# N_A_761_113#_M1042_s
+ N_A_761_113#_M1047_s N_A_761_113#_M1034_g N_A_761_113#_c_1276_n
+ N_A_761_113#_M1040_g N_A_761_113#_c_1277_n N_A_761_113#_c_1278_n
+ N_A_761_113#_c_1279_n N_A_761_113#_M1039_g N_A_761_113#_c_1280_n
+ N_A_761_113#_c_1281_n N_A_761_113#_c_1282_n N_A_761_113#_M1043_g
+ N_A_761_113#_c_1298_n N_A_761_113#_c_1299_n N_A_761_113#_c_1284_n
+ N_A_761_113#_c_1285_n N_A_761_113#_c_1300_n N_A_761_113#_M1020_g
+ N_A_761_113#_M1000_g N_A_761_113#_c_1302_n N_A_761_113#_c_1303_n
+ N_A_761_113#_c_1286_n N_A_761_113#_c_1287_n N_A_761_113#_c_1288_n
+ N_A_761_113#_M1028_g N_A_761_113#_c_1290_n N_A_761_113#_c_1291_n
+ N_A_761_113#_c_1305_n N_A_761_113#_c_1292_n N_A_761_113#_c_1307_n
+ N_A_761_113#_c_1293_n N_A_761_113#_c_1294_n N_A_761_113#_c_1310_n
+ N_A_761_113#_c_1295_n PM_SKY130_FD_SC_LP__SDFSBP_LP%A_761_113#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2220_40# N_A_2220_40#_M1013_s
+ N_A_2220_40#_M1012_s N_A_2220_40#_M1029_g N_A_2220_40#_c_1488_n
+ N_A_2220_40#_M1021_g N_A_2220_40#_c_1496_n N_A_2220_40#_c_1489_n
+ N_A_2220_40#_c_1490_n N_A_2220_40#_c_1491_n N_A_2220_40#_c_1492_n
+ N_A_2220_40#_c_1497_n N_A_2220_40#_c_1493_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2220_40#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2019_419# N_A_2019_419#_M1022_d
+ N_A_2019_419#_M1000_d N_A_2019_419#_M1027_d N_A_2019_419#_M1013_g
+ N_A_2019_419#_c_1575_n N_A_2019_419#_c_1576_n N_A_2019_419#_M1014_g
+ N_A_2019_419#_M1012_g N_A_2019_419#_c_1578_n N_A_2019_419#_M1036_g
+ N_A_2019_419#_c_1579_n N_A_2019_419#_c_1580_n N_A_2019_419#_c_1581_n
+ N_A_2019_419#_c_1582_n N_A_2019_419#_M1038_g N_A_2019_419#_c_1583_n
+ N_A_2019_419#_M1017_g N_A_2019_419#_c_1585_n N_A_2019_419#_c_1586_n
+ N_A_2019_419#_M1044_g N_A_2019_419#_M1009_g N_A_2019_419#_c_1588_n
+ N_A_2019_419#_M1030_g N_A_2019_419#_c_1589_n N_A_2019_419#_c_1590_n
+ N_A_2019_419#_c_1591_n N_A_2019_419#_c_1592_n N_A_2019_419#_c_1609_n
+ N_A_2019_419#_c_1593_n N_A_2019_419#_c_1594_n N_A_2019_419#_c_1595_n
+ N_A_2019_419#_c_1633_n N_A_2019_419#_c_1603_n N_A_2019_419#_c_1641_n
+ N_A_2019_419#_c_1604_n N_A_2019_419#_c_1642_n N_A_2019_419#_c_1596_n
+ N_A_2019_419#_c_1597_n N_A_2019_419#_c_1605_n N_A_2019_419#_c_1606_n
+ N_A_2019_419#_c_1685_n N_A_2019_419#_c_1607_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2019_419#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2865_74# N_A_2865_74#_M1044_s
+ N_A_2865_74#_M1009_s N_A_2865_74#_c_1794_n N_A_2865_74#_M1019_g
+ N_A_2865_74#_M1003_g N_A_2865_74#_M1041_g N_A_2865_74#_c_1786_n
+ N_A_2865_74#_c_1787_n N_A_2865_74#_c_1788_n N_A_2865_74#_c_1796_n
+ N_A_2865_74#_c_1789_n N_A_2865_74#_c_1790_n N_A_2865_74#_c_1791_n
+ N_A_2865_74#_c_1792_n N_A_2865_74#_c_1793_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2865_74#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%VPWR N_VPWR_M1010_d N_VPWR_M1046_d
+ N_VPWR_M1047_d N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_M1021_d N_VPWR_M1012_d
+ N_VPWR_M1009_d N_VPWR_c_1854_n N_VPWR_c_1855_n N_VPWR_c_1856_n N_VPWR_c_1857_n
+ N_VPWR_c_1858_n N_VPWR_c_1859_n N_VPWR_c_1860_n N_VPWR_c_1861_n
+ N_VPWR_c_1862_n N_VPWR_c_1863_n N_VPWR_c_1864_n VPWR N_VPWR_c_1865_n
+ N_VPWR_c_1866_n N_VPWR_c_1867_n N_VPWR_c_1868_n N_VPWR_c_1869_n
+ N_VPWR_c_1870_n N_VPWR_c_1853_n N_VPWR_c_1872_n N_VPWR_c_1873_n
+ N_VPWR_c_1874_n N_VPWR_c_1875_n N_VPWR_c_1876_n N_VPWR_c_1877_n
+ N_VPWR_c_1878_n PM_SKY130_FD_SC_LP__SDFSBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_245_409# N_A_245_409#_M1045_s
+ N_A_245_409#_M1024_d N_A_245_409#_c_2022_n N_A_245_409#_c_2023_n
+ N_A_245_409#_c_2024_n N_A_245_409#_c_2029_n N_A_245_409#_c_2030_n
+ N_A_245_409#_c_2031_n N_A_245_409#_c_2025_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%A_245_409#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%A_352_409# N_A_352_409#_M1016_d
+ N_A_352_409#_M1043_s N_A_352_409#_M1045_d N_A_352_409#_M1008_s
+ N_A_352_409#_c_2096_n N_A_352_409#_c_2090_n N_A_352_409#_c_2091_n
+ N_A_352_409#_c_2074_n N_A_352_409#_c_2075_n N_A_352_409#_c_2076_n
+ N_A_352_409#_c_2077_n N_A_352_409#_c_2078_n N_A_352_409#_c_2079_n
+ N_A_352_409#_c_2080_n N_A_352_409#_c_2081_n N_A_352_409#_c_2082_n
+ N_A_352_409#_c_2083_n N_A_352_409#_c_2084_n N_A_352_409#_c_2085_n
+ N_A_352_409#_c_2093_n N_A_352_409#_c_2086_n N_A_352_409#_c_2087_n
+ N_A_352_409#_c_2139_n N_A_352_409#_c_2088_n N_A_352_409#_c_2089_n
+ N_A_352_409#_c_2095_n PM_SKY130_FD_SC_LP__SDFSBP_LP%A_352_409#
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%Q_N N_Q_N_M1038_d N_Q_N_M1017_d N_Q_N_c_2268_n
+ N_Q_N_c_2273_n Q_N Q_N Q_N Q_N N_Q_N_c_2270_n N_Q_N_c_2271_n
+ PM_SKY130_FD_SC_LP__SDFSBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%Q N_Q_M1041_d N_Q_M1019_d N_Q_c_2311_n Q Q Q
+ N_Q_c_2314_n N_Q_c_2312_n PM_SKY130_FD_SC_LP__SDFSBP_LP%Q
x_PM_SKY130_FD_SC_LP__SDFSBP_LP%VGND N_VGND_M1007_d N_VGND_M1033_d
+ N_VGND_M1006_d N_VGND_M1011_d N_VGND_M1037_d N_VGND_M1048_d N_VGND_M1014_d
+ N_VGND_M1030_d N_VGND_c_2335_n N_VGND_c_2336_n N_VGND_c_2337_n N_VGND_c_2338_n
+ N_VGND_c_2339_n N_VGND_c_2340_n N_VGND_c_2341_n N_VGND_c_2342_n
+ N_VGND_c_2343_n N_VGND_c_2344_n VGND N_VGND_c_2345_n N_VGND_c_2346_n
+ N_VGND_c_2347_n N_VGND_c_2348_n N_VGND_c_2349_n N_VGND_c_2350_n
+ N_VGND_c_2351_n N_VGND_c_2352_n N_VGND_c_2353_n N_VGND_c_2354_n
+ N_VGND_c_2355_n N_VGND_c_2356_n N_VGND_c_2357_n N_VGND_c_2358_n
+ N_VGND_c_2359_n N_VGND_c_2360_n PM_SKY130_FD_SC_LP__SDFSBP_LP%VGND
cc_1 VNB N_SCE_M1010_g 0.0416063f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_2 VNB N_SCE_M1023_g 0.0358922f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.445
cc_3 VNB N_SCE_c_333_n 0.0128837f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.11
cc_4 VNB N_SCE_M1007_g 0.0229033f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_5 VNB N_SCE_c_335_n 0.012551f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.11
cc_6 VNB N_SCE_c_336_n 0.0139924f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=0.73
cc_7 VNB N_SCE_c_337_n 0.00854036f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=0.88
cc_8 VNB N_SCE_c_338_n 0.0135498f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.12
cc_9 VNB N_SCE_c_339_n 0.0238997f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.625
cc_10 VNB N_SCE_c_340_n 0.00205846f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.79
cc_11 VNB N_SCE_c_341_n 0.0299599f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.02
cc_12 VNB N_SCE_c_342_n 0.006395f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.045
cc_13 VNB N_SCE_c_343_n 0.00543481f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_14 VNB N_SCE_c_344_n 0.0120135f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.195
cc_15 VNB N_SCE_c_345_n 0.0161348f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_16 VNB N_SCE_c_346_n 0.00886132f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.045
cc_17 VNB N_SCE_c_347_n 0.00430375f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=1.045
cc_18 VNB N_A_27_409#_c_440_n 0.0316342f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_19 VNB N_A_27_409#_c_441_n 0.0163133f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_20 VNB N_A_27_409#_c_442_n 0.0249404f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.445
cc_21 VNB N_A_27_409#_c_443_n 0.0114478f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.445
cc_22 VNB N_A_27_409#_c_444_n 0.0142885f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_23 VNB N_A_27_409#_c_445_n 0.0523146f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.11
cc_24 VNB N_A_27_409#_c_446_n 0.00394592f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.02
cc_25 VNB N_A_27_409#_c_447_n 0.0104307f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_26 VNB N_D_M1016_g 0.0498011f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.445
cc_27 VNB D 0.00319663f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.11
cc_28 VNB N_D_c_509_n 0.0153543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_SCD_c_550_n 0.0168176f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.185
cc_30 VNB N_SCD_c_551_n 0.0224492f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_31 VNB SCD 0.00311164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_SCD_c_553_n 0.0684031f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_33 VNB N_SCD_c_554_n 0.0146821f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=2.545
cc_34 VNB N_CLK_M1042_g 0.0204989f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_35 VNB N_CLK_c_604_n 0.0228399f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.445
cc_36 VNB N_CLK_M1006_g 0.0178711f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_37 VNB N_CLK_c_606_n 0.0179947f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.445
cc_38 VNB CLK 0.00287673f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.445
cc_39 VNB N_CLK_c_608_n 0.00498413f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_40 VNB N_A_987_409#_M1018_g 0.0235177f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_41 VNB N_A_987_409#_c_657_n 0.00362479f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.625
cc_42 VNB N_A_987_409#_c_658_n 0.0119592f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.02
cc_43 VNB N_A_987_409#_c_659_n 0.0292866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_987_409#_c_660_n 0.00929646f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.84
cc_45 VNB N_A_987_409#_c_661_n 0.0340604f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=0.84
cc_46 VNB N_A_987_409#_c_662_n 0.00619271f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.02
cc_47 VNB N_A_987_409#_c_663_n 0.00905831f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.045
cc_48 VNB N_A_987_409#_c_664_n 0.0175712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_987_409#_c_665_n 0.00617082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_987_409#_c_666_n 2.06456e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_987_409#_c_667_n 0.0100917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_987_409#_c_668_n 0.0192932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1423_99#_M1011_g 0.0365611f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.11
cc_54 VNB N_A_1423_99#_c_869_n 0.00217892f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.88
cc_55 VNB N_A_1423_99#_c_870_n 0.0297966f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_56 VNB N_A_1423_99#_c_871_n 0.0179156f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_57 VNB N_A_1423_99#_c_872_n 0.00550319f $X=-0.19 $Y=-0.245 $X2=2.655
+ $Y2=2.545
cc_58 VNB N_A_1423_99#_c_873_n 0.00770186f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_59 VNB N_A_1423_99#_c_874_n 0.00810752f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.02
cc_60 VNB N_A_1201_419#_c_949_n 0.0174032f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.445
cc_61 VNB N_A_1201_419#_c_950_n 0.0107278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1201_419#_c_951_n 0.0173062f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.73
cc_63 VNB N_A_1201_419#_M1002_g 0.0200402f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.11
cc_64 VNB N_A_1201_419#_c_953_n 0.0214232f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.12
cc_65 VNB N_A_1201_419#_c_954_n 0.00529599f $X=-0.19 $Y=-0.245 $X2=2.275
+ $Y2=1.195
cc_66 VNB N_A_1201_419#_c_955_n 0.00723397f $X=-0.19 $Y=-0.245 $X2=2.672
+ $Y2=1.28
cc_67 VNB N_A_1201_419#_c_956_n 0.0126151f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_68 VNB N_A_1201_419#_c_957_n 0.0249251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1201_419#_c_958_n 0.00348498f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=0.84
cc_70 VNB N_A_1201_419#_c_959_n 0.00163489f $X=-0.19 $Y=-0.245 $X2=2.075
+ $Y2=0.84
cc_71 VNB N_A_1201_419#_c_960_n 0.00929075f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_72 VNB N_A_1201_419#_c_961_n 0.0038168f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.11
cc_73 VNB N_A_1201_419#_c_962_n 0.00861335f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=1.045
cc_74 VNB N_A_1201_419#_c_963_n 0.0057805f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.045
cc_75 VNB N_A_1201_419#_c_964_n 0.0049364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1201_419#_c_965_n 0.00579562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1201_419#_c_966_n 0.00513707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1201_419#_c_967_n 0.0145087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1201_419#_c_968_n 0.0179362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_SET_B_M1037_g 0.036722f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.445
cc_81 VNB N_SET_B_c_1148_n 0.017129f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.11
cc_82 VNB N_SET_B_c_1149_n 0.0342178f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_83 VNB N_SET_B_c_1150_n 0.00771918f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_84 VNB N_SET_B_c_1151_n 0.0237848f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_85 VNB N_SET_B_c_1152_n 0.00109121f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=2.545
cc_86 VNB N_SET_B_c_1153_n 5.93655e-19 $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.11
cc_87 VNB SET_B 0.00270455f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=0.88
cc_88 VNB N_SET_B_c_1155_n 0.0169015f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.02
cc_89 VNB N_SET_B_c_1156_n 0.0113848f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.045
cc_90 VNB N_SET_B_c_1157_n 0.00187773f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_91 VNB N_SET_B_c_1158_n 0.0347167f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.195
cc_92 VNB N_A_761_113#_c_1276_n 0.0135195f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.855
cc_93 VNB N_A_761_113#_c_1277_n 0.0221339f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.73
cc_94 VNB N_A_761_113#_c_1278_n 0.00724822f $X=-0.19 $Y=-0.245 $X2=2.555
+ $Y2=0.445
cc_95 VNB N_A_761_113#_c_1279_n 0.015684f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.88
cc_96 VNB N_A_761_113#_c_1280_n 0.052887f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=2.545
cc_97 VNB N_A_761_113#_c_1281_n 0.0175779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_761_113#_c_1282_n 0.022435f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.11
cc_99 VNB N_A_761_113#_M1043_g 0.0194388f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.12
cc_100 VNB N_A_761_113#_c_1284_n 0.334181f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.02
cc_101 VNB N_A_761_113#_c_1285_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.02
cc_102 VNB N_A_761_113#_c_1286_n 0.0187734f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_103 VNB N_A_761_113#_c_1287_n 0.0201998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_761_113#_c_1288_n 0.00866264f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=0.84
cc_105 VNB N_A_761_113#_M1028_g 0.0265219f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_106 VNB N_A_761_113#_c_1290_n 0.0046367f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=1.02
cc_107 VNB N_A_761_113#_c_1291_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=0.855
cc_108 VNB N_A_761_113#_c_1292_n 0.0126431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_761_113#_c_1293_n 0.00164109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_761_113#_c_1294_n 0.0177347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_761_113#_c_1295_n 0.00242811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2220_40#_M1029_g 0.0360294f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.11
cc_113 VNB N_A_2220_40#_c_1488_n 0.061624f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.855
cc_114 VNB N_A_2220_40#_c_1489_n 0.00546287f $X=-0.19 $Y=-0.245 $X2=2.655
+ $Y2=1.79
cc_115 VNB N_A_2220_40#_c_1490_n 0.00265771f $X=-0.19 $Y=-0.245 $X2=2.655
+ $Y2=2.545
cc_116 VNB N_A_2220_40#_c_1491_n 0.0135141f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=1.11
cc_117 VNB N_A_2220_40#_c_1492_n 0.011827f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.02
cc_118 VNB N_A_2220_40#_c_1493_n 0.00593972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2019_419#_M1013_g 0.0356483f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.445
cc_120 VNB N_A_2019_419#_c_1575_n 0.0108061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_2019_419#_c_1576_n 0.00896356f $X=-0.19 $Y=-0.245 $X2=2.555
+ $Y2=0.73
cc_122 VNB N_A_2019_419#_M1014_g 0.0351977f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=0.88
cc_123 VNB N_A_2019_419#_c_1578_n 0.0136473f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=1.11
cc_124 VNB N_A_2019_419#_c_1579_n 0.0166386f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_125 VNB N_A_2019_419#_c_1580_n 0.00964834f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.625
cc_126 VNB N_A_2019_419#_c_1581_n 0.00735986f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.79
cc_127 VNB N_A_2019_419#_c_1582_n 0.0170358f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.02
cc_128 VNB N_A_2019_419#_c_1583_n 0.0398726f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=1.02
cc_129 VNB N_A_2019_419#_M1017_g 0.0247057f $X=-0.19 $Y=-0.245 $X2=2.04
+ $Y2=1.045
cc_130 VNB N_A_2019_419#_c_1585_n 0.0423767f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.195
cc_131 VNB N_A_2019_419#_c_1586_n 0.0174274f $X=-0.19 $Y=-0.245 $X2=2.672
+ $Y2=1.28
cc_132 VNB N_A_2019_419#_M1009_g 0.0446898f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=0.84
cc_133 VNB N_A_2019_419#_c_1588_n 0.01411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_2019_419#_c_1589_n 0.0139138f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=0.855
cc_135 VNB N_A_2019_419#_c_1590_n 0.00580226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_2019_419#_c_1591_n 0.0178063f $X=-0.19 $Y=-0.245 $X2=2.275
+ $Y2=1.045
cc_137 VNB N_A_2019_419#_c_1592_n 0.0126933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_2019_419#_c_1593_n 0.0188831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_2019_419#_c_1594_n 0.00407158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_2019_419#_c_1595_n 0.00493733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_2019_419#_c_1596_n 0.00624999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_2019_419#_c_1597_n 0.0274823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_2865_74#_M1003_g 0.0203009f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.445
cc_144 VNB N_A_2865_74#_M1041_g 0.0264335f $X=-0.19 $Y=-0.245 $X2=2.555
+ $Y2=0.445
cc_145 VNB N_A_2865_74#_c_1786_n 0.0123434f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=0.88
cc_146 VNB N_A_2865_74#_c_1787_n 0.0256476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_2865_74#_c_1788_n 0.0128113f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=0.88
cc_148 VNB N_A_2865_74#_c_1789_n 0.0115614f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=1.02
cc_149 VNB N_A_2865_74#_c_1790_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=1.8
+ $Y2=1.045
cc_150 VNB N_A_2865_74#_c_1791_n 0.0285864f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.195
cc_151 VNB N_A_2865_74#_c_1792_n 0.00856748f $X=-0.19 $Y=-0.245 $X2=2.672
+ $Y2=1.285
cc_152 VNB N_A_2865_74#_c_1793_n 0.00887229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VPWR_c_1853_n 0.681144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_352_409#_c_2074_n 0.0102129f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=1.12
cc_155 VNB N_A_352_409#_c_2075_n 0.00535067f $X=-0.19 $Y=-0.245 $X2=2.655
+ $Y2=2.545
cc_156 VNB N_A_352_409#_c_2076_n 0.00958083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_A_352_409#_c_2077_n 0.00805858f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=0.88
cc_158 VNB N_A_352_409#_c_2078_n 0.0225539f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_159 VNB N_A_352_409#_c_2079_n 0.00358581f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.12
cc_160 VNB N_A_352_409#_c_2080_n 0.00179493f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.79
cc_161 VNB N_A_352_409#_c_2081_n 0.00910579f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.02
cc_162 VNB N_A_352_409#_c_2082_n 4.42176e-19 $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=1.02
cc_163 VNB N_A_352_409#_c_2083_n 0.00173012f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=1.02
cc_164 VNB N_A_352_409#_c_2084_n 0.0212329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_A_352_409#_c_2085_n 0.00291864f $X=-0.19 $Y=-0.245 $X2=2.04
+ $Y2=1.045
cc_166 VNB N_A_352_409#_c_2086_n 0.00214722f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=0.84
cc_167 VNB N_A_352_409#_c_2087_n 0.00298693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_A_352_409#_c_2088_n 0.00842906f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=0.855
cc_169 VNB N_A_352_409#_c_2089_n 0.0065073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_Q_N_c_2268_n 0.0063437f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.445
cc_171 VNB Q_N 0.00813609f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=0.445
cc_172 VNB N_Q_N_c_2270_n 3.43398e-19 $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=0.73
cc_173 VNB N_Q_N_c_2271_n 0.0125023f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.02
cc_174 VNB N_Q_c_2311_n 0.0255421f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.11
cc_175 VNB N_Q_c_2312_n 0.0406949f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.625
cc_176 VNB N_VGND_c_2335_n 0.00548094f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_177 VNB N_VGND_c_2336_n 0.00708737f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.02
cc_178 VNB N_VGND_c_2337_n 0.0132052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2338_n 0.0120044f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=1.195
cc_180 VNB N_VGND_c_2339_n 0.0163182f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_181 VNB N_VGND_c_2340_n 0.0120509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2341_n 0.00526739f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.855
cc_183 VNB N_VGND_c_2342_n 0.0153684f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.045
cc_184 VNB N_VGND_c_2343_n 0.0327909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2344_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=1.045
cc_186 VNB N_VGND_c_2345_n 0.0305356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2346_n 0.0446941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2347_n 0.0650097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_VGND_c_2348_n 0.0347337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_VGND_c_2349_n 0.0660237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_191 VNB N_VGND_c_2350_n 0.0291285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_192 VNB N_VGND_c_2351_n 0.0492505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_193 VNB N_VGND_c_2352_n 0.0280628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_194 VNB N_VGND_c_2353_n 0.827466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_195 VNB N_VGND_c_2354_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_196 VNB N_VGND_c_2355_n 0.00510766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_197 VNB N_VGND_c_2356_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_198 VNB N_VGND_c_2357_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_199 VNB N_VGND_c_2358_n 0.00585462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_200 VNB N_VGND_c_2359_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_201 VNB N_VGND_c_2360_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_202 VPB N_SCE_M1010_g 0.0571298f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_203 VPB N_SCE_M1046_g 0.0303663f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=2.545
cc_204 VPB N_SCE_c_340_n 0.0114869f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.79
cc_205 VPB N_SCE_c_351_n 6.99016e-19 $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_206 VPB N_A_27_409#_M1045_g 0.0443959f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.11
cc_207 VPB N_A_27_409#_c_442_n 0.0220293f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=0.445
cc_208 VPB N_A_27_409#_c_443_n 0.00366841f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=0.445
cc_209 VPB N_A_27_409#_c_451_n 0.0531568f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.12
cc_210 VPB N_A_27_409#_c_446_n 0.00646656f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.02
cc_211 VPB N_A_27_409#_c_447_n 0.00453508f $X=-0.19 $Y=1.655 $X2=1.8 $Y2=1.045
cc_212 VPB N_D_M1031_g 0.0307404f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_213 VPB D 0.00288225f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.11
cc_214 VPB N_D_c_509_n 0.0093985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_SCD_M1024_g 0.0366762f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.445
cc_216 VPB SCD 0.00666349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_SCD_c_553_n 0.023946f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=1.12
cc_218 VPB N_CLK_M1047_g 0.0361437f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.11
cc_219 VPB CLK 0.00234957f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=0.445
cc_220 VPB N_CLK_c_608_n 0.0128414f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=1.79
cc_221 VPB N_A_987_409#_M1008_g 0.0405391f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.11
cc_222 VPB N_A_987_409#_M1035_g 0.0293041f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=1.79
cc_223 VPB N_A_987_409#_c_671_n 0.0074982f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.11
cc_224 VPB N_A_987_409#_c_672_n 0.010702f $X=-0.19 $Y=1.655 $X2=2.57 $Y2=0.88
cc_225 VPB N_A_987_409#_c_673_n 0.00251866f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.285
cc_226 VPB N_A_987_409#_c_674_n 0.00332444f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.02
cc_227 VPB N_A_987_409#_c_675_n 0.00282811f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.285
cc_228 VPB N_A_987_409#_c_662_n 0.00251445f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.02
cc_229 VPB N_A_987_409#_c_664_n 0.0101687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_987_409#_c_665_n 0.00261578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_987_409#_c_666_n 5.97937e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_987_409#_c_667_n 0.0207726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1423_99#_M1004_g 0.0347232f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.445
cc_234 VPB N_A_1423_99#_c_869_n 0.00470401f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.88
cc_235 VPB N_A_1423_99#_c_870_n 0.0330447f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=1.12
cc_236 VPB N_A_1423_99#_c_878_n 0.0113971f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.11
cc_237 VPB N_A_1201_419#_M1026_g 0.0306599f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.11
cc_238 VPB N_A_1201_419#_M1025_g 0.0324088f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=1.79
cc_239 VPB N_A_1201_419#_c_953_n 0.00390768f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.12
cc_240 VPB N_A_1201_419#_c_972_n 0.0138055f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.625
cc_241 VPB N_A_1201_419#_c_973_n 0.00654541f $X=-0.19 $Y=1.655 $X2=1.095
+ $Y2=1.02
cc_242 VPB N_A_1201_419#_c_974_n 0.00276195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1201_419#_c_954_n 0.00941752f $X=-0.19 $Y=1.655 $X2=2.275
+ $Y2=1.195
cc_244 VPB N_A_1201_419#_c_959_n 0.00412877f $X=-0.19 $Y=1.655 $X2=2.075
+ $Y2=0.84
cc_245 VPB N_A_1201_419#_c_960_n 0.0172475f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.285
cc_246 VPB N_A_1201_419#_c_966_n 0.00134312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_SET_B_M1005_g 0.0317962f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_248 VPB N_SET_B_M1027_g 0.0351313f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.88
cc_249 VPB N_SET_B_c_1151_n 0.0178545f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=1.79
cc_250 VPB N_SET_B_c_1153_n 0.00396468f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.11
cc_251 VPB SET_B 0.00130979f $X=-0.19 $Y=1.655 $X2=2.57 $Y2=0.88
cc_252 VPB N_SET_B_c_1155_n 0.0244663f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.02
cc_253 VPB N_SET_B_c_1156_n 0.0177182f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.045
cc_254 VPB N_SET_B_c_1157_n 0.00343611f $X=-0.19 $Y=1.655 $X2=1.8 $Y2=1.045
cc_255 VPB N_A_761_113#_M1034_g 0.0293162f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.11
cc_256 VPB N_A_761_113#_c_1282_n 0.0169276f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.11
cc_257 VPB N_A_761_113#_c_1298_n 0.0262822f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.625
cc_258 VPB N_A_761_113#_c_1299_n 0.0115398f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.79
cc_259 VPB N_A_761_113#_c_1300_n 0.0220437f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.02
cc_260 VPB N_A_761_113#_M1000_g 0.0315059f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.195
cc_261 VPB N_A_761_113#_c_1302_n 0.0277013f $X=-0.19 $Y=1.655 $X2=2.672 $Y2=1.28
cc_262 VPB N_A_761_113#_c_1303_n 0.00859771f $X=-0.19 $Y=1.655 $X2=2.672
+ $Y2=1.285
cc_263 VPB N_A_761_113#_c_1286_n 0.00377826f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.285
cc_264 VPB N_A_761_113#_c_1305_n 0.0118214f $X=-0.19 $Y=1.655 $X2=1.565
+ $Y2=1.045
cc_265 VPB N_A_761_113#_c_1292_n 0.00707126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_761_113#_c_1307_n 0.00386474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_761_113#_c_1293_n 5.74637e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_761_113#_c_1294_n 0.0278062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_761_113#_c_1310_n 0.00621098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_2220_40#_c_1488_n 0.0260955f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=0.855
cc_271 VPB N_A_2220_40#_M1021_g 0.0300127f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.445
cc_272 VPB N_A_2220_40#_c_1496_n 0.0025059f $X=-0.19 $Y=1.655 $X2=2.555
+ $Y2=0.445
cc_273 VPB N_A_2220_40#_c_1497_n 0.0102983f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.02
cc_274 VPB N_A_2220_40#_c_1493_n 0.00783433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_2019_419#_M1012_g 0.0300153f $X=-0.19 $Y=1.655 $X2=2.655
+ $Y2=2.545
cc_276 VPB N_A_2019_419#_M1017_g 0.045923f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.045
cc_277 VPB N_A_2019_419#_M1009_g 0.0318444f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.84
cc_278 VPB N_A_2019_419#_c_1590_n 0.0245563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_2019_419#_c_1595_n 0.00302646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_2019_419#_c_1603_n 0.00445816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_A_2019_419#_c_1604_n 0.0122288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_A_2019_419#_c_1605_n 0.00167999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_2019_419#_c_1606_n 0.00279664f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_2019_419#_c_1607_n 0.00408534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_A_2865_74#_c_1794_n 0.0251587f $X=-0.19 $Y=1.655 $X2=0.615
+ $Y2=0.445
cc_286 VPB N_A_2865_74#_c_1786_n 0.0121354f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.88
cc_287 VPB N_A_2865_74#_c_1796_n 0.0194066f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.625
cc_288 VPB N_A_2865_74#_c_1789_n 0.00354496f $X=-0.19 $Y=1.655 $X2=1.095
+ $Y2=1.02
cc_289 VPB N_VPWR_c_1854_n 0.0167989f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.625
cc_290 VPB N_VPWR_c_1855_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1856_n 0.00177638f $X=-0.19 $Y=1.655 $X2=2.275 $Y2=1.195
cc_292 VPB N_VPWR_c_1857_n 0.00284591f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_293 VPB N_VPWR_c_1858_n 0.017902f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.84
cc_294 VPB N_VPWR_c_1859_n 0.00284591f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_295 VPB N_VPWR_c_1860_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1861_n 0.0068482f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.045
cc_297 VPB N_VPWR_c_1862_n 0.0139381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_1863_n 0.0432384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1864_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_1865_n 0.0336586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_1866_n 0.0704474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_1867_n 0.0678789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_1868_n 0.0435469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1869_n 0.0356754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_1870_n 0.0270602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_1853_n 0.123833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_1872_n 0.0243996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_1873_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_1874_n 0.00510127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_1875_n 0.00510127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_1876_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_1877_n 0.00428995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_1878_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_314 VPB N_A_245_409#_c_2022_n 0.00386309f $X=-0.19 $Y=1.655 $X2=0.615
+ $Y2=0.445
cc_315 VPB N_A_245_409#_c_2023_n 0.0106538f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.11
cc_316 VPB N_A_245_409#_c_2024_n 0.00378074f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=0.855
cc_317 VPB N_A_245_409#_c_2025_n 0.00922767f $X=-0.19 $Y=1.655 $X2=2.655
+ $Y2=2.545
cc_318 VPB N_A_352_409#_c_2090_n 0.0137929f $X=-0.19 $Y=1.655 $X2=2.555
+ $Y2=0.445
cc_319 VPB N_A_352_409#_c_2091_n 0.00245018f $X=-0.19 $Y=1.655 $X2=2.585
+ $Y2=0.88
cc_320 VPB N_A_352_409#_c_2075_n 0.0026312f $X=-0.19 $Y=1.655 $X2=2.655
+ $Y2=2.545
cc_321 VPB N_A_352_409#_c_2093_n 0.00656379f $X=-0.19 $Y=1.655 $X2=2.672
+ $Y2=1.285
cc_322 VPB N_A_352_409#_c_2089_n 0.00619447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_A_352_409#_c_2095_n 0.0157462f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.045
cc_324 VPB N_Q_N_c_2268_n 0.00124977f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.445
cc_325 VPB N_Q_N_c_2273_n 0.00470039f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.855
cc_326 VPB N_Q_N_c_2270_n 0.0029883f $X=-0.19 $Y=1.655 $X2=2.57 $Y2=0.73
cc_327 VPB Q 0.043263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_Q_c_2314_n 0.0284669f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.12
cc_329 VPB N_Q_c_2312_n 0.00986018f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.625
cc_330 N_SCE_c_343_n N_A_27_409#_c_440_n 0.0182902f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_331 N_SCE_M1007_g N_A_27_409#_c_441_n 0.00685901f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_332 N_SCE_M1010_g N_A_27_409#_c_442_n 0.00979362f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_333 N_SCE_c_341_n N_A_27_409#_c_442_n 0.0106932f $X=1.095 $Y=1.02 $X2=0 $Y2=0
cc_334 N_SCE_c_346_n N_A_27_409#_c_442_n 0.0103951f $X=1.565 $Y=1.045 $X2=0
+ $Y2=0
cc_335 N_SCE_c_343_n N_A_27_409#_c_443_n 7.75503e-19 $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_336 N_SCE_M1007_g N_A_27_409#_c_444_n 0.00333275f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_337 N_SCE_c_341_n N_A_27_409#_c_444_n 0.0125709f $X=1.095 $Y=1.02 $X2=0 $Y2=0
cc_338 N_SCE_c_342_n N_A_27_409#_c_444_n 0.00119626f $X=2.04 $Y=1.045 $X2=0
+ $Y2=0
cc_339 N_SCE_c_343_n N_A_27_409#_c_444_n 0.00893034f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_340 N_SCE_M1010_g N_A_27_409#_c_445_n 0.0181295f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_341 N_SCE_M1023_g N_A_27_409#_c_445_n 0.0213242f $X=0.615 $Y=0.445 $X2=0
+ $Y2=0
cc_342 N_SCE_M1007_g N_A_27_409#_c_445_n 0.00204936f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_343 N_SCE_c_335_n N_A_27_409#_c_445_n 0.0113095f $X=0.555 $Y=1.11 $X2=0 $Y2=0
cc_344 N_SCE_c_346_n N_A_27_409#_c_445_n 0.0144418f $X=1.565 $Y=1.045 $X2=0
+ $Y2=0
cc_345 N_SCE_M1010_g N_A_27_409#_c_451_n 0.0366051f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_346 N_SCE_M1010_g N_A_27_409#_c_446_n 0.0173611f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_347 N_SCE_c_335_n N_A_27_409#_c_446_n 0.0134343f $X=0.555 $Y=1.11 $X2=0 $Y2=0
cc_348 N_SCE_c_341_n N_A_27_409#_c_446_n 7.69499e-19 $X=1.095 $Y=1.02 $X2=0
+ $Y2=0
cc_349 N_SCE_c_346_n N_A_27_409#_c_446_n 0.0269786f $X=1.565 $Y=1.045 $X2=0
+ $Y2=0
cc_350 N_SCE_M1010_g N_A_27_409#_c_447_n 0.0173508f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_351 N_SCE_M1046_g N_D_M1031_g 0.0765858f $X=2.655 $Y=2.545 $X2=0 $Y2=0
cc_352 N_SCE_c_336_n N_D_M1016_g 0.0174476f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_353 N_SCE_c_338_n N_D_M1016_g 0.0228082f $X=2.675 $Y=1.12 $X2=0 $Y2=0
cc_354 N_SCE_c_351_n N_D_M1016_g 0.00109329f $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_355 N_SCE_c_347_n N_D_M1016_g 0.0222793f $X=2.275 $Y=1.045 $X2=0 $Y2=0
cc_356 N_SCE_c_339_n D 0.00113718f $X=2.675 $Y=1.625 $X2=0 $Y2=0
cc_357 N_SCE_c_343_n D 0.0566403f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_358 N_SCE_c_351_n D 0.0220339f $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_359 N_SCE_c_339_n N_D_c_509_n 0.0207503f $X=2.675 $Y=1.625 $X2=0 $Y2=0
cc_360 N_SCE_c_342_n N_D_c_509_n 0.00186599f $X=2.04 $Y=1.045 $X2=0 $Y2=0
cc_361 N_SCE_c_351_n N_D_c_509_n 4.1374e-19 $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_362 N_SCE_c_347_n N_D_c_509_n 0.00262094f $X=2.275 $Y=1.045 $X2=0 $Y2=0
cc_363 N_SCE_c_336_n N_SCD_c_550_n 0.032078f $X=2.57 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_364 N_SCE_M1046_g N_SCD_M1024_g 0.0469913f $X=2.655 $Y=2.545 $X2=0 $Y2=0
cc_365 N_SCE_c_339_n N_SCD_M1024_g 0.0197752f $X=2.675 $Y=1.625 $X2=0 $Y2=0
cc_366 N_SCE_c_337_n N_SCD_c_551_n 0.00972694f $X=2.57 $Y=0.88 $X2=0 $Y2=0
cc_367 N_SCE_c_338_n N_SCD_c_553_n 2.64808e-19 $X=2.675 $Y=1.12 $X2=0 $Y2=0
cc_368 N_SCE_c_344_n N_SCD_c_553_n 2.1929e-19 $X=2.51 $Y=1.195 $X2=0 $Y2=0
cc_369 N_SCE_c_351_n N_SCD_c_553_n 5.76172e-19 $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_370 N_SCE_c_345_n N_SCD_c_553_n 0.0197752f $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_371 N_SCE_c_338_n N_SCD_c_554_n 0.00556564f $X=2.675 $Y=1.12 $X2=0 $Y2=0
cc_372 N_SCE_M1010_g N_VPWR_c_1854_n 0.0250662f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_373 N_SCE_M1046_g N_VPWR_c_1855_n 0.011031f $X=2.655 $Y=2.545 $X2=0 $Y2=0
cc_374 N_SCE_M1046_g N_VPWR_c_1863_n 0.0073986f $X=2.655 $Y=2.545 $X2=0 $Y2=0
cc_375 N_SCE_M1010_g N_VPWR_c_1853_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_376 N_SCE_M1046_g N_VPWR_c_1853_n 0.00723273f $X=2.655 $Y=2.545 $X2=0 $Y2=0
cc_377 N_SCE_M1010_g N_VPWR_c_1872_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_378 N_SCE_M1010_g N_A_245_409#_c_2022_n 3.95513e-19 $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_379 N_SCE_M1010_g N_A_245_409#_c_2023_n 0.00155163f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_380 N_SCE_M1046_g N_A_245_409#_c_2024_n 0.00522741f $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_381 N_SCE_M1046_g N_A_245_409#_c_2029_n 0.00993317f $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_382 N_SCE_M1046_g N_A_245_409#_c_2030_n 0.0127459f $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_383 N_SCE_M1046_g N_A_245_409#_c_2031_n 0.00238028f $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_384 N_SCE_M1046_g N_A_245_409#_c_2025_n 8.77766e-19 $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_385 N_SCE_M1046_g N_A_352_409#_c_2096_n 0.00108911f $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_386 N_SCE_M1046_g N_A_352_409#_c_2090_n 0.0146911f $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_387 N_SCE_c_340_n N_A_352_409#_c_2090_n 7.46077e-19 $X=2.675 $Y=1.79 $X2=0
+ $Y2=0
cc_388 N_SCE_c_351_n N_A_352_409#_c_2090_n 0.0237712f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_389 N_SCE_c_337_n N_A_352_409#_c_2074_n 0.00196542f $X=2.57 $Y=0.88 $X2=0
+ $Y2=0
cc_390 N_SCE_c_338_n N_A_352_409#_c_2074_n 0.00139015f $X=2.675 $Y=1.12 $X2=0
+ $Y2=0
cc_391 N_SCE_c_344_n N_A_352_409#_c_2074_n 0.0167042f $X=2.51 $Y=1.195 $X2=0
+ $Y2=0
cc_392 N_SCE_c_345_n N_A_352_409#_c_2074_n 0.00137074f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_393 N_SCE_M1046_g N_A_352_409#_c_2075_n 0.00348712f $X=2.655 $Y=2.545 $X2=0
+ $Y2=0
cc_394 N_SCE_c_338_n N_A_352_409#_c_2075_n 0.00318194f $X=2.675 $Y=1.12 $X2=0
+ $Y2=0
cc_395 N_SCE_c_344_n N_A_352_409#_c_2075_n 0.0130532f $X=2.51 $Y=1.195 $X2=0
+ $Y2=0
cc_396 N_SCE_c_351_n N_A_352_409#_c_2075_n 0.0365638f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_397 N_SCE_c_345_n N_A_352_409#_c_2075_n 0.00365786f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_398 N_SCE_c_336_n N_A_352_409#_c_2087_n 0.0125964f $X=2.57 $Y=0.73 $X2=0
+ $Y2=0
cc_399 N_SCE_c_337_n N_A_352_409#_c_2087_n 0.00343365f $X=2.57 $Y=0.88 $X2=0
+ $Y2=0
cc_400 N_SCE_c_338_n N_A_352_409#_c_2087_n 0.00250647f $X=2.675 $Y=1.12 $X2=0
+ $Y2=0
cc_401 N_SCE_c_344_n N_A_352_409#_c_2087_n 0.0197901f $X=2.51 $Y=1.195 $X2=0
+ $Y2=0
cc_402 N_SCE_c_347_n N_A_352_409#_c_2087_n 0.0161592f $X=2.275 $Y=1.045 $X2=0
+ $Y2=0
cc_403 N_SCE_M1023_g N_VGND_c_2335_n 0.00239701f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_404 N_SCE_M1007_g N_VGND_c_2335_n 0.0137855f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_405 N_SCE_c_341_n N_VGND_c_2335_n 0.00417255f $X=1.095 $Y=1.02 $X2=0 $Y2=0
cc_406 N_SCE_c_346_n N_VGND_c_2335_n 0.0262295f $X=1.565 $Y=1.045 $X2=0 $Y2=0
cc_407 N_SCE_c_336_n N_VGND_c_2336_n 0.00207237f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_408 N_SCE_M1023_g N_VGND_c_2345_n 0.00549284f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_409 N_SCE_M1007_g N_VGND_c_2345_n 0.00486043f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_410 N_SCE_c_336_n N_VGND_c_2346_n 0.00362516f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_411 N_SCE_c_337_n N_VGND_c_2346_n 4.97855e-19 $X=2.57 $Y=0.88 $X2=0 $Y2=0
cc_412 N_SCE_M1023_g N_VGND_c_2353_n 0.0110955f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_413 N_SCE_M1007_g N_VGND_c_2353_n 0.0045337f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_414 N_SCE_c_336_n N_VGND_c_2353_n 0.00539979f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_415 N_SCE_c_337_n N_VGND_c_2353_n 8.18184e-19 $X=2.57 $Y=0.88 $X2=0 $Y2=0
cc_416 N_SCE_c_343_n N_VGND_c_2353_n 0.0215311f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_417 N_SCE_c_346_n N_VGND_c_2353_n 0.0112235f $X=1.565 $Y=1.045 $X2=0 $Y2=0
cc_418 N_A_27_409#_M1045_g N_D_M1031_g 0.0336853f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_419 N_A_27_409#_c_440_n N_D_M1016_g 0.0216441f $X=1.655 $Y=1.425 $X2=0 $Y2=0
cc_420 N_A_27_409#_c_441_n N_D_M1016_g 0.0419662f $X=1.735 $Y=0.73 $X2=0 $Y2=0
cc_421 N_A_27_409#_c_443_n N_D_M1016_g 0.00182095f $X=1.635 $Y=1.59 $X2=0 $Y2=0
cc_422 N_A_27_409#_M1045_g D 0.0108293f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_423 N_A_27_409#_c_443_n D 0.0149066f $X=1.635 $Y=1.59 $X2=0 $Y2=0
cc_424 N_A_27_409#_c_446_n D 0.0236784f $X=1.22 $Y=1.59 $X2=0 $Y2=0
cc_425 N_A_27_409#_c_443_n N_D_c_509_n 0.0214736f $X=1.635 $Y=1.59 $X2=0 $Y2=0
cc_426 N_A_27_409#_M1045_g N_VPWR_c_1854_n 0.00380434f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_427 N_A_27_409#_c_451_n N_VPWR_c_1854_n 0.0685263f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_428 N_A_27_409#_c_446_n N_VPWR_c_1854_n 0.0207871f $X=1.22 $Y=1.59 $X2=0
+ $Y2=0
cc_429 N_A_27_409#_M1045_g N_VPWR_c_1863_n 0.00546179f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_430 N_A_27_409#_M1045_g N_VPWR_c_1853_n 0.00832053f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_431 N_A_27_409#_c_451_n N_VPWR_c_1853_n 0.0125808f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_432 N_A_27_409#_c_451_n N_VPWR_c_1872_n 0.0220321f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_433 N_A_27_409#_M1045_g N_A_245_409#_c_2022_n 9.65935e-19 $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_434 N_A_27_409#_M1045_g N_A_245_409#_c_2023_n 0.0167532f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_435 N_A_27_409#_c_442_n N_A_245_409#_c_2023_n 0.00891589f $X=1.51 $Y=1.59
+ $X2=0 $Y2=0
cc_436 N_A_27_409#_c_446_n N_A_245_409#_c_2023_n 0.0106951f $X=1.22 $Y=1.59
+ $X2=0 $Y2=0
cc_437 N_A_27_409#_M1045_g N_A_245_409#_c_2024_n 0.0164696f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_438 N_A_27_409#_M1045_g N_A_352_409#_c_2096_n 0.0103858f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_439 N_A_27_409#_M1045_g N_A_352_409#_c_2091_n 0.00598618f $X=1.635 $Y=2.545
+ $X2=0 $Y2=0
cc_440 N_A_27_409#_c_441_n N_A_352_409#_c_2087_n 0.00180434f $X=1.735 $Y=0.73
+ $X2=0 $Y2=0
cc_441 N_A_27_409#_c_441_n N_VGND_c_2335_n 0.0122158f $X=1.735 $Y=0.73 $X2=0
+ $Y2=0
cc_442 N_A_27_409#_c_445_n N_VGND_c_2335_n 0.0133046f $X=0.4 $Y=0.47 $X2=0 $Y2=0
cc_443 N_A_27_409#_c_445_n N_VGND_c_2345_n 0.0278794f $X=0.4 $Y=0.47 $X2=0 $Y2=0
cc_444 N_A_27_409#_c_441_n N_VGND_c_2346_n 0.00585385f $X=1.735 $Y=0.73 $X2=0
+ $Y2=0
cc_445 N_A_27_409#_c_444_n N_VGND_c_2346_n 0.0016562f $X=1.735 $Y=0.805 $X2=0
+ $Y2=0
cc_446 N_A_27_409#_M1023_s N_VGND_c_2353_n 0.00232985f $X=0.255 $Y=0.235 $X2=0
+ $Y2=0
cc_447 N_A_27_409#_c_441_n N_VGND_c_2353_n 0.0070095f $X=1.735 $Y=0.73 $X2=0
+ $Y2=0
cc_448 N_A_27_409#_c_444_n N_VGND_c_2353_n 0.00218182f $X=1.735 $Y=0.805 $X2=0
+ $Y2=0
cc_449 N_A_27_409#_c_445_n N_VGND_c_2353_n 0.017224f $X=0.4 $Y=0.47 $X2=0 $Y2=0
cc_450 N_D_M1031_g N_VPWR_c_1855_n 8.56804e-19 $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_451 N_D_M1031_g N_VPWR_c_1863_n 0.00546209f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_452 N_D_M1031_g N_VPWR_c_1853_n 0.00735468f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_453 N_D_M1031_g N_A_245_409#_c_2023_n 8.93568e-19 $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_454 N_D_M1031_g N_A_245_409#_c_2024_n 0.0199598f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_455 N_D_M1031_g N_A_245_409#_c_2029_n 0.00579089f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_456 N_D_M1031_g N_A_245_409#_c_2031_n 0.00169926f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_457 N_D_M1031_g N_A_352_409#_c_2096_n 0.0102338f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_458 N_D_M1031_g N_A_352_409#_c_2090_n 0.0183326f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_459 D N_A_352_409#_c_2090_n 0.0160355f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_460 N_D_c_509_n N_A_352_409#_c_2090_n 2.22766e-19 $X=2.135 $Y=1.625 $X2=0
+ $Y2=0
cc_461 N_D_M1031_g N_A_352_409#_c_2091_n 0.00163487f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_462 D N_A_352_409#_c_2091_n 0.027305f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_463 N_D_c_509_n N_A_352_409#_c_2091_n 0.00162266f $X=2.135 $Y=1.625 $X2=0
+ $Y2=0
cc_464 N_D_M1016_g N_A_352_409#_c_2087_n 0.0109415f $X=2.125 $Y=0.445 $X2=0
+ $Y2=0
cc_465 N_D_M1016_g N_VGND_c_2346_n 0.0054778f $X=2.125 $Y=0.445 $X2=0 $Y2=0
cc_466 N_D_M1016_g N_VGND_c_2353_n 0.00623217f $X=2.125 $Y=0.445 $X2=0 $Y2=0
cc_467 N_SCD_c_553_n N_CLK_M1042_g 0.0167961f $X=3.525 $Y=1.275 $X2=0 $Y2=0
cc_468 N_SCD_M1024_g N_A_761_113#_c_1305_n 0.00597732f $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_469 N_SCD_M1024_g N_A_761_113#_c_1292_n 0.00435208f $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_470 SCD N_A_761_113#_c_1292_n 0.048119f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_471 N_SCD_c_553_n N_A_761_113#_c_1292_n 0.00573299f $X=3.525 $Y=1.275 $X2=0
+ $Y2=0
cc_472 N_SCD_M1024_g N_A_761_113#_c_1310_n 0.00308709f $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_473 N_SCD_c_551_n N_A_761_113#_c_1295_n 5.47566e-19 $X=3.155 $Y=0.805 $X2=0
+ $Y2=0
cc_474 N_SCD_c_554_n N_A_761_113#_c_1295_n 0.00387488f $X=3.375 $Y=1.11 $X2=0
+ $Y2=0
cc_475 N_SCD_M1024_g N_VPWR_c_1855_n 0.0122002f $X=3.185 $Y=2.545 $X2=0 $Y2=0
cc_476 N_SCD_M1024_g N_VPWR_c_1865_n 0.00769046f $X=3.185 $Y=2.545 $X2=0 $Y2=0
cc_477 N_SCD_M1024_g N_VPWR_c_1853_n 0.00833754f $X=3.185 $Y=2.545 $X2=0 $Y2=0
cc_478 N_SCD_M1024_g N_A_245_409#_c_2029_n 8.04314e-19 $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_479 N_SCD_M1024_g N_A_245_409#_c_2030_n 0.0167894f $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_480 N_SCD_M1024_g N_A_245_409#_c_2025_n 0.012954f $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_481 SCD N_A_245_409#_c_2025_n 0.00879654f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_482 N_SCD_c_553_n N_A_245_409#_c_2025_n 0.00161435f $X=3.525 $Y=1.275 $X2=0
+ $Y2=0
cc_483 N_SCD_M1024_g N_A_352_409#_c_2090_n 0.00925578f $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_484 N_SCD_c_551_n N_A_352_409#_c_2074_n 0.00838022f $X=3.155 $Y=0.805 $X2=0
+ $Y2=0
cc_485 N_SCD_M1024_g N_A_352_409#_c_2075_n 0.010005f $X=3.185 $Y=2.545 $X2=0
+ $Y2=0
cc_486 SCD N_A_352_409#_c_2075_n 0.0455899f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_487 N_SCD_c_553_n N_A_352_409#_c_2075_n 0.0194436f $X=3.525 $Y=1.275 $X2=0
+ $Y2=0
cc_488 N_SCD_c_554_n N_A_352_409#_c_2075_n 0.0097416f $X=3.375 $Y=1.11 $X2=0
+ $Y2=0
cc_489 N_SCD_c_551_n N_A_352_409#_c_2076_n 0.00337262f $X=3.155 $Y=0.805 $X2=0
+ $Y2=0
cc_490 SCD N_A_352_409#_c_2076_n 0.0250574f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_491 N_SCD_c_553_n N_A_352_409#_c_2076_n 0.00782825f $X=3.525 $Y=1.275 $X2=0
+ $Y2=0
cc_492 N_SCD_c_554_n N_A_352_409#_c_2076_n 0.00320065f $X=3.375 $Y=1.11 $X2=0
+ $Y2=0
cc_493 N_SCD_c_550_n N_A_352_409#_c_2077_n 0.00355564f $X=2.945 $Y=0.73 $X2=0
+ $Y2=0
cc_494 N_SCD_c_551_n N_A_352_409#_c_2077_n 0.00100252f $X=3.155 $Y=0.805 $X2=0
+ $Y2=0
cc_495 SCD N_A_352_409#_c_2078_n 2.33898e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_496 N_SCD_c_550_n N_A_352_409#_c_2087_n 0.00224553f $X=2.945 $Y=0.73 $X2=0
+ $Y2=0
cc_497 N_SCD_c_551_n N_A_352_409#_c_2139_n 0.00425826f $X=3.155 $Y=0.805 $X2=0
+ $Y2=0
cc_498 N_SCD_c_554_n N_A_352_409#_c_2139_n 0.00125883f $X=3.375 $Y=1.11 $X2=0
+ $Y2=0
cc_499 N_SCD_c_550_n N_VGND_c_2336_n 0.0112135f $X=2.945 $Y=0.73 $X2=0 $Y2=0
cc_500 N_SCD_c_551_n N_VGND_c_2336_n 0.0052461f $X=3.155 $Y=0.805 $X2=0 $Y2=0
cc_501 N_SCD_c_550_n N_VGND_c_2346_n 0.00367954f $X=2.945 $Y=0.73 $X2=0 $Y2=0
cc_502 N_SCD_c_550_n N_VGND_c_2353_n 0.0043701f $X=2.945 $Y=0.73 $X2=0 $Y2=0
cc_503 N_CLK_M1006_g N_A_761_113#_c_1276_n 0.0108964f $X=4.525 $Y=0.775 $X2=0
+ $Y2=0
cc_504 N_CLK_c_604_n N_A_761_113#_c_1277_n 0.00762099f $X=4.282 $Y=1.588 $X2=0
+ $Y2=0
cc_505 CLK N_A_761_113#_c_1277_n 0.00124206f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_506 N_CLK_c_606_n N_A_761_113#_c_1290_n 0.0108964f $X=4.345 $Y=1.315 $X2=0
+ $Y2=0
cc_507 N_CLK_M1047_g N_A_761_113#_c_1305_n 0.0168451f $X=4.28 $Y=2.545 $X2=0
+ $Y2=0
cc_508 N_CLK_M1042_g N_A_761_113#_c_1292_n 0.0123407f $X=4.165 $Y=0.775 $X2=0
+ $Y2=0
cc_509 N_CLK_M1047_g N_A_761_113#_c_1292_n 0.00686465f $X=4.28 $Y=2.545 $X2=0
+ $Y2=0
cc_510 CLK N_A_761_113#_c_1292_n 0.0241667f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_511 N_CLK_M1047_g N_A_761_113#_c_1307_n 0.0188849f $X=4.28 $Y=2.545 $X2=0
+ $Y2=0
cc_512 CLK N_A_761_113#_c_1307_n 0.030946f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_513 N_CLK_c_608_n N_A_761_113#_c_1307_n 0.00183219f $X=4.31 $Y=1.615 $X2=0
+ $Y2=0
cc_514 N_CLK_M1047_g N_A_761_113#_c_1293_n 8.93373e-19 $X=4.28 $Y=2.545 $X2=0
+ $Y2=0
cc_515 CLK N_A_761_113#_c_1293_n 0.0173664f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_516 N_CLK_c_604_n N_A_761_113#_c_1294_n 0.0142084f $X=4.282 $Y=1.588 $X2=0
+ $Y2=0
cc_517 N_CLK_M1047_g N_A_761_113#_c_1294_n 0.0312092f $X=4.28 $Y=2.545 $X2=0
+ $Y2=0
cc_518 CLK N_A_761_113#_c_1294_n 0.00180942f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_519 N_CLK_M1047_g N_A_761_113#_c_1310_n 0.00338717f $X=4.28 $Y=2.545 $X2=0
+ $Y2=0
cc_520 N_CLK_c_608_n N_A_761_113#_c_1310_n 0.00311128f $X=4.31 $Y=1.615 $X2=0
+ $Y2=0
cc_521 N_CLK_M1042_g N_A_761_113#_c_1295_n 0.0057338f $X=4.165 $Y=0.775 $X2=0
+ $Y2=0
cc_522 N_CLK_M1006_g N_A_761_113#_c_1295_n 3.08234e-19 $X=4.525 $Y=0.775 $X2=0
+ $Y2=0
cc_523 N_CLK_M1047_g N_VPWR_c_1856_n 0.0189165f $X=4.28 $Y=2.545 $X2=0 $Y2=0
cc_524 N_CLK_M1047_g N_VPWR_c_1865_n 0.00769046f $X=4.28 $Y=2.545 $X2=0 $Y2=0
cc_525 N_CLK_M1047_g N_VPWR_c_1853_n 0.0143431f $X=4.28 $Y=2.545 $X2=0 $Y2=0
cc_526 N_CLK_M1047_g N_A_245_409#_c_2025_n 0.00105075f $X=4.28 $Y=2.545 $X2=0
+ $Y2=0
cc_527 N_CLK_M1042_g N_A_352_409#_c_2077_n 0.00311563f $X=4.165 $Y=0.775 $X2=0
+ $Y2=0
cc_528 N_CLK_M1042_g N_A_352_409#_c_2078_n 0.00707754f $X=4.165 $Y=0.775 $X2=0
+ $Y2=0
cc_529 N_CLK_M1006_g N_A_352_409#_c_2078_n 2.48962e-19 $X=4.525 $Y=0.775 $X2=0
+ $Y2=0
cc_530 N_CLK_M1042_g N_A_352_409#_c_2080_n 0.00366721f $X=4.165 $Y=0.775 $X2=0
+ $Y2=0
cc_531 N_CLK_M1006_g N_A_352_409#_c_2080_n 0.0117179f $X=4.525 $Y=0.775 $X2=0
+ $Y2=0
cc_532 N_CLK_M1006_g N_A_352_409#_c_2081_n 0.00727325f $X=4.525 $Y=0.775 $X2=0
+ $Y2=0
cc_533 N_CLK_c_606_n N_A_352_409#_c_2081_n 0.00348762f $X=4.345 $Y=1.315 $X2=0
+ $Y2=0
cc_534 CLK N_A_352_409#_c_2081_n 0.0131191f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_535 N_CLK_M1042_g N_A_352_409#_c_2082_n 5.77011e-19 $X=4.165 $Y=0.775 $X2=0
+ $Y2=0
cc_536 N_CLK_M1006_g N_A_352_409#_c_2082_n 4.60164e-19 $X=4.525 $Y=0.775 $X2=0
+ $Y2=0
cc_537 N_CLK_c_606_n N_A_352_409#_c_2082_n 0.00624734f $X=4.345 $Y=1.315 $X2=0
+ $Y2=0
cc_538 CLK N_A_352_409#_c_2082_n 0.0129587f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_539 N_CLK_M1006_g N_A_352_409#_c_2083_n 6.6435e-19 $X=4.525 $Y=0.775 $X2=0
+ $Y2=0
cc_540 N_CLK_c_604_n N_A_352_409#_c_2088_n 2.00473e-19 $X=4.282 $Y=1.588 $X2=0
+ $Y2=0
cc_541 N_CLK_c_606_n N_A_352_409#_c_2088_n 2.455e-19 $X=4.345 $Y=1.315 $X2=0
+ $Y2=0
cc_542 CLK N_A_352_409#_c_2089_n 0.00317994f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_543 N_CLK_M1006_g N_VGND_c_2337_n 9.43806e-19 $X=4.525 $Y=0.775 $X2=0 $Y2=0
cc_544 N_CLK_M1006_g N_VGND_c_2343_n 0.00409299f $X=4.525 $Y=0.775 $X2=0 $Y2=0
cc_545 N_CLK_M1006_g N_VGND_c_2353_n 0.00437698f $X=4.525 $Y=0.775 $X2=0 $Y2=0
cc_546 N_A_987_409#_c_681_p N_A_1423_99#_M1026_d 0.00473561f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_547 N_A_987_409#_M1018_g N_A_1423_99#_M1011_g 0.03516f $X=6.83 $Y=0.835 $X2=0
+ $Y2=0
cc_548 N_A_987_409#_c_658_n N_A_1423_99#_M1011_g 3.85439e-19 $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_549 N_A_987_409#_c_684_p N_A_1423_99#_M1004_g 0.0195517f $X=7.39 $Y=2.98
+ $X2=0 $Y2=0
cc_550 N_A_987_409#_c_685_p N_A_1423_99#_M1004_g 0.00652195f $X=7.475 $Y=2.895
+ $X2=0 $Y2=0
cc_551 N_A_987_409#_c_686_p N_A_1423_99#_M1004_g 0.0071872f $X=7.56 $Y=2.6 $X2=0
+ $Y2=0
cc_552 N_A_987_409#_c_659_n N_A_1423_99#_c_870_n 0.03516f $X=6.74 $Y=1.465 $X2=0
+ $Y2=0
cc_553 N_A_987_409#_c_681_p N_A_1423_99#_c_870_n 5.40025e-19 $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_554 N_A_987_409#_c_686_p N_A_1423_99#_c_870_n 3.45105e-19 $X=7.56 $Y=2.6
+ $X2=0 $Y2=0
cc_555 N_A_987_409#_c_681_p N_A_1423_99#_c_888_n 0.0159455f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_556 N_A_987_409#_c_686_p N_A_1423_99#_c_888_n 0.009183f $X=7.56 $Y=2.6 $X2=0
+ $Y2=0
cc_557 N_A_987_409#_c_681_p N_A_1423_99#_c_878_n 0.0461265f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_558 N_A_987_409#_c_674_n N_A_1201_419#_M1008_d 0.0086935f $X=6.045 $Y=2.895
+ $X2=0 $Y2=0
cc_559 N_A_987_409#_c_684_p N_A_1201_419#_M1008_d 0.0159428f $X=7.39 $Y=2.98
+ $X2=0 $Y2=0
cc_560 N_A_987_409#_c_695_p N_A_1201_419#_M1008_d 6.69812e-19 $X=6.045 $Y=2.98
+ $X2=0 $Y2=0
cc_561 N_A_987_409#_c_685_p N_A_1201_419#_M1026_g 0.00253853f $X=7.475 $Y=2.895
+ $X2=0 $Y2=0
cc_562 N_A_987_409#_c_681_p N_A_1201_419#_M1026_g 0.0183911f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_563 N_A_987_409#_c_681_p N_A_1201_419#_M1025_g 0.0215879f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_564 N_A_987_409#_c_660_n N_A_1201_419#_M1002_g 2.89045e-19 $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_565 N_A_987_409#_c_661_n N_A_1201_419#_M1002_g 0.00249151f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_566 N_A_987_409#_c_668_n N_A_1201_419#_M1002_g 0.0223907f $X=9.98 $Y=1.155
+ $X2=0 $Y2=0
cc_567 N_A_987_409#_c_660_n N_A_1201_419#_c_953_n 0.00300375f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_568 N_A_987_409#_c_666_n N_A_1201_419#_c_953_n 0.00222853f $X=9.98 $Y=1.69
+ $X2=0 $Y2=0
cc_569 N_A_987_409#_c_681_p N_A_1201_419#_c_972_n 2.07832e-19 $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_570 N_A_987_409#_c_675_n N_A_1201_419#_c_972_n 0.00620283f $X=9.9 $Y=2.515
+ $X2=0 $Y2=0
cc_571 N_A_987_409#_M1008_g N_A_1201_419#_c_992_n 0.00152258f $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_572 N_A_987_409#_c_674_n N_A_1201_419#_c_992_n 0.0343853f $X=6.045 $Y=2.895
+ $X2=0 $Y2=0
cc_573 N_A_987_409#_c_684_p N_A_1201_419#_c_992_n 0.0194739f $X=7.39 $Y=2.98
+ $X2=0 $Y2=0
cc_574 N_A_987_409#_c_658_n N_A_1201_419#_c_973_n 0.00881594f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_575 N_A_987_409#_c_659_n N_A_1201_419#_c_973_n 0.00150336f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_576 N_A_987_409#_c_684_p N_A_1201_419#_c_973_n 0.0120907f $X=7.39 $Y=2.98
+ $X2=0 $Y2=0
cc_577 N_A_987_409#_M1008_g N_A_1201_419#_c_974_n 6.20042e-19 $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_578 N_A_987_409#_c_674_n N_A_1201_419#_c_974_n 0.0133149f $X=6.045 $Y=2.895
+ $X2=0 $Y2=0
cc_579 N_A_987_409#_c_658_n N_A_1201_419#_c_974_n 0.0142118f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_580 N_A_987_409#_M1018_g N_A_1201_419#_c_1001_n 0.00850648f $X=6.83 $Y=0.835
+ $X2=0 $Y2=0
cc_581 N_A_987_409#_c_658_n N_A_1201_419#_c_1001_n 0.00645661f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_582 N_A_987_409#_M1018_g N_A_1201_419#_c_954_n 0.00476116f $X=6.83 $Y=0.835
+ $X2=0 $Y2=0
cc_583 N_A_987_409#_c_658_n N_A_1201_419#_c_954_n 0.0250969f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_584 N_A_987_409#_c_659_n N_A_1201_419#_c_954_n 9.7274e-19 $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_585 N_A_987_409#_c_681_p N_A_1201_419#_c_959_n 3.87968e-19 $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_586 N_A_987_409#_M1018_g N_A_1201_419#_c_965_n 0.00738595f $X=6.83 $Y=0.835
+ $X2=0 $Y2=0
cc_587 N_A_987_409#_c_657_n N_A_1201_419#_c_965_n 0.00191579f $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_588 N_A_987_409#_c_658_n N_A_1201_419#_c_965_n 0.0214455f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_589 N_A_987_409#_c_659_n N_A_1201_419#_c_965_n 0.00398645f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_590 N_A_987_409#_c_663_n N_A_1201_419#_c_965_n 0.00519813f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_591 N_A_987_409#_c_681_p N_A_1201_419#_c_966_n 0.00760442f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_592 N_A_987_409#_c_660_n N_A_1201_419#_c_966_n 0.026624f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_593 N_A_987_409#_c_661_n N_A_1201_419#_c_966_n 9.90146e-19 $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_594 N_A_987_409#_c_675_n N_A_1201_419#_c_966_n 0.00606062f $X=9.9 $Y=2.515
+ $X2=0 $Y2=0
cc_595 N_A_987_409#_c_666_n N_A_1201_419#_c_966_n 0.0101635f $X=9.98 $Y=1.69
+ $X2=0 $Y2=0
cc_596 N_A_987_409#_c_660_n N_A_1201_419#_c_967_n 2.14095e-19 $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_597 N_A_987_409#_c_661_n N_A_1201_419#_c_967_n 0.0176692f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_598 N_A_987_409#_c_681_p N_SET_B_M1005_g 0.0241312f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_599 N_A_987_409#_c_660_n N_SET_B_c_1151_n 0.00847092f $X=9.98 $Y=1.32 $X2=0
+ $Y2=0
cc_600 N_A_987_409#_c_662_n N_SET_B_c_1151_n 0.0350015f $X=10.715 $Y=1.69 $X2=0
+ $Y2=0
cc_601 N_A_987_409#_c_666_n N_SET_B_c_1151_n 0.0223376f $X=9.98 $Y=1.69 $X2=0
+ $Y2=0
cc_602 N_A_987_409#_c_667_n N_SET_B_c_1151_n 0.00277703f $X=10.88 $Y=1.77 $X2=0
+ $Y2=0
cc_603 N_A_987_409#_c_681_p N_SET_B_c_1153_n 0.00616039f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_604 N_A_987_409#_c_681_p N_SET_B_c_1155_n 9.98371e-19 $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_605 N_A_987_409#_c_671_n N_A_761_113#_M1034_g 0.0108317f $X=5.075 $Y=2.475
+ $X2=0 $Y2=0
cc_606 N_A_987_409#_c_673_n N_A_761_113#_M1034_g 0.00359736f $X=5.24 $Y=2.98
+ $X2=0 $Y2=0
cc_607 N_A_987_409#_c_663_n N_A_761_113#_c_1276_n 3.04539e-19 $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_608 N_A_987_409#_c_657_n N_A_761_113#_c_1277_n 2.53501e-19 $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_609 N_A_987_409#_c_664_n N_A_761_113#_c_1277_n 0.00117f $X=5.84 $Y=1.615
+ $X2=0 $Y2=0
cc_610 N_A_987_409#_c_657_n N_A_761_113#_c_1279_n 0.00105896f $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_611 N_A_987_409#_c_663_n N_A_761_113#_c_1279_n 0.00497645f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_612 N_A_987_409#_c_657_n N_A_761_113#_c_1280_n 0.0153148f $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_613 N_A_987_409#_c_663_n N_A_761_113#_c_1280_n 0.0115092f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_614 N_A_987_409#_c_664_n N_A_761_113#_c_1280_n 0.0172301f $X=5.84 $Y=1.615
+ $X2=0 $Y2=0
cc_615 N_A_987_409#_c_665_n N_A_761_113#_c_1280_n 0.00816481f $X=6.13 $Y=1.54
+ $X2=0 $Y2=0
cc_616 N_A_987_409#_M1018_g N_A_761_113#_c_1281_n 0.00967771f $X=6.83 $Y=0.835
+ $X2=0 $Y2=0
cc_617 N_A_987_409#_c_657_n N_A_761_113#_c_1281_n 0.00103285f $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_618 N_A_987_409#_c_658_n N_A_761_113#_c_1281_n 0.00123456f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_619 N_A_987_409#_c_663_n N_A_761_113#_c_1281_n 0.00188274f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_620 N_A_987_409#_c_657_n N_A_761_113#_c_1282_n 0.00246531f $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_621 N_A_987_409#_c_674_n N_A_761_113#_c_1282_n 0.00547693f $X=6.045 $Y=2.895
+ $X2=0 $Y2=0
cc_622 N_A_987_409#_c_658_n N_A_761_113#_c_1282_n 0.0236476f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_623 N_A_987_409#_c_659_n N_A_761_113#_c_1282_n 0.021337f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_624 N_A_987_409#_c_664_n N_A_761_113#_c_1282_n 0.0176878f $X=5.84 $Y=1.615
+ $X2=0 $Y2=0
cc_625 N_A_987_409#_c_665_n N_A_761_113#_c_1282_n 0.00402605f $X=6.13 $Y=1.54
+ $X2=0 $Y2=0
cc_626 N_A_987_409#_M1018_g N_A_761_113#_M1043_g 0.0104517f $X=6.83 $Y=0.835
+ $X2=0 $Y2=0
cc_627 N_A_987_409#_c_663_n N_A_761_113#_M1043_g 0.00156348f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_628 N_A_987_409#_c_658_n N_A_761_113#_c_1298_n 0.0057037f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_629 N_A_987_409#_c_659_n N_A_761_113#_c_1298_n 0.0167375f $X=6.74 $Y=1.465
+ $X2=0 $Y2=0
cc_630 N_A_987_409#_M1008_g N_A_761_113#_c_1299_n 0.0176878f $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_631 N_A_987_409#_M1018_g N_A_761_113#_c_1284_n 0.00860793f $X=6.83 $Y=0.835
+ $X2=0 $Y2=0
cc_632 N_A_987_409#_c_668_n N_A_761_113#_c_1284_n 0.00907339f $X=9.98 $Y=1.155
+ $X2=0 $Y2=0
cc_633 N_A_987_409#_M1008_g N_A_761_113#_c_1300_n 0.0145942f $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_634 N_A_987_409#_c_674_n N_A_761_113#_c_1300_n 0.00490093f $X=6.045 $Y=2.895
+ $X2=0 $Y2=0
cc_635 N_A_987_409#_c_684_p N_A_761_113#_c_1300_n 0.0182317f $X=7.39 $Y=2.98
+ $X2=0 $Y2=0
cc_636 N_A_987_409#_c_685_p N_A_761_113#_c_1300_n 8.76528e-19 $X=7.475 $Y=2.895
+ $X2=0 $Y2=0
cc_637 N_A_987_409#_c_686_p N_A_761_113#_c_1300_n 7.00849e-19 $X=7.56 $Y=2.6
+ $X2=0 $Y2=0
cc_638 N_A_987_409#_c_681_p N_A_761_113#_M1000_g 0.00878814f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_639 N_A_987_409#_c_675_n N_A_761_113#_M1000_g 0.0218613f $X=9.9 $Y=2.515
+ $X2=0 $Y2=0
cc_640 N_A_987_409#_c_662_n N_A_761_113#_M1000_g 3.1459e-19 $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_641 N_A_987_409#_c_667_n N_A_761_113#_M1000_g 0.019313f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_642 N_A_987_409#_c_662_n N_A_761_113#_c_1302_n 0.0119165f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_643 N_A_987_409#_c_666_n N_A_761_113#_c_1302_n 0.00284081f $X=9.98 $Y=1.69
+ $X2=0 $Y2=0
cc_644 N_A_987_409#_c_661_n N_A_761_113#_c_1303_n 0.0165547f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_645 N_A_987_409#_c_675_n N_A_761_113#_c_1303_n 0.00573205f $X=9.9 $Y=2.515
+ $X2=0 $Y2=0
cc_646 N_A_987_409#_c_666_n N_A_761_113#_c_1303_n 0.00958194f $X=9.98 $Y=1.69
+ $X2=0 $Y2=0
cc_647 N_A_987_409#_c_660_n N_A_761_113#_c_1286_n 0.00415815f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_648 N_A_987_409#_c_662_n N_A_761_113#_c_1286_n 0.00779306f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_649 N_A_987_409#_c_667_n N_A_761_113#_c_1286_n 0.0180907f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_650 N_A_987_409#_c_662_n N_A_761_113#_c_1287_n 0.00494977f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_651 N_A_987_409#_c_667_n N_A_761_113#_c_1287_n 0.00825615f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_652 N_A_987_409#_c_660_n N_A_761_113#_c_1288_n 0.0019115f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_653 N_A_987_409#_c_661_n N_A_761_113#_c_1288_n 0.018124f $X=9.98 $Y=1.32
+ $X2=0 $Y2=0
cc_654 N_A_987_409#_c_668_n N_A_761_113#_M1028_g 0.00735708f $X=9.98 $Y=1.155
+ $X2=0 $Y2=0
cc_655 N_A_987_409#_M1034_d N_A_761_113#_c_1307_n 0.00263338f $X=4.935 $Y=2.045
+ $X2=0 $Y2=0
cc_656 N_A_987_409#_M1008_g N_A_761_113#_c_1307_n 5.67789e-19 $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_657 N_A_987_409#_c_671_n N_A_761_113#_c_1307_n 0.0145008f $X=5.075 $Y=2.475
+ $X2=0 $Y2=0
cc_658 N_A_987_409#_M1008_g N_A_761_113#_c_1294_n 0.00131971f $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_659 N_A_987_409#_c_671_n N_A_761_113#_c_1294_n 0.00100762f $X=5.075 $Y=2.475
+ $X2=0 $Y2=0
cc_660 N_A_987_409#_c_664_n N_A_761_113#_c_1294_n 0.00379283f $X=5.84 $Y=1.615
+ $X2=0 $Y2=0
cc_661 N_A_987_409#_c_662_n N_A_2220_40#_c_1488_n 3.28355e-19 $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_662 N_A_987_409#_c_667_n N_A_2220_40#_c_1488_n 0.0181784f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_663 N_A_987_409#_M1035_g N_A_2220_40#_M1021_g 0.0549773f $X=10.84 $Y=2.595
+ $X2=0 $Y2=0
cc_664 N_A_987_409#_c_667_n N_A_2220_40#_M1021_g 0.00258148f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_665 N_A_987_409#_c_668_n N_A_2019_419#_c_1592_n 0.0114537f $X=9.98 $Y=1.155
+ $X2=0 $Y2=0
cc_666 N_A_987_409#_M1035_g N_A_2019_419#_c_1609_n 0.023789f $X=10.84 $Y=2.595
+ $X2=0 $Y2=0
cc_667 N_A_987_409#_c_662_n N_A_2019_419#_c_1609_n 0.0225963f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_668 N_A_987_409#_c_667_n N_A_2019_419#_c_1609_n 0.00171515f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_669 N_A_987_409#_c_662_n N_A_2019_419#_c_1593_n 0.00602547f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_670 N_A_987_409#_c_667_n N_A_2019_419#_c_1593_n 0.00216442f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_671 N_A_987_409#_c_662_n N_A_2019_419#_c_1594_n 0.00772114f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_672 N_A_987_409#_c_668_n N_A_2019_419#_c_1594_n 0.0049388f $X=9.98 $Y=1.155
+ $X2=0 $Y2=0
cc_673 N_A_987_409#_M1035_g N_A_2019_419#_c_1595_n 0.00333471f $X=10.84 $Y=2.595
+ $X2=0 $Y2=0
cc_674 N_A_987_409#_c_662_n N_A_2019_419#_c_1595_n 0.0224635f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_675 N_A_987_409#_c_667_n N_A_2019_419#_c_1595_n 0.00184117f $X=10.88 $Y=1.77
+ $X2=0 $Y2=0
cc_676 N_A_987_409#_M1035_g N_A_2019_419#_c_1606_n 0.0217744f $X=10.84 $Y=2.595
+ $X2=0 $Y2=0
cc_677 N_A_987_409#_c_681_p N_A_2019_419#_c_1606_n 0.0114736f $X=9.815 $Y=2.6
+ $X2=0 $Y2=0
cc_678 N_A_987_409#_c_675_n N_A_2019_419#_c_1606_n 0.0273782f $X=9.9 $Y=2.515
+ $X2=0 $Y2=0
cc_679 N_A_987_409#_c_662_n N_A_2019_419#_c_1606_n 0.0144528f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_680 N_A_987_409#_c_684_p N_VPWR_M1004_d 0.00277849f $X=7.39 $Y=2.98 $X2=0
+ $Y2=0
cc_681 N_A_987_409#_c_685_p N_VPWR_M1004_d 0.00300067f $X=7.475 $Y=2.895 $X2=0
+ $Y2=0
cc_682 N_A_987_409#_c_681_p N_VPWR_M1004_d 0.0129248f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_683 N_A_987_409#_c_686_p N_VPWR_M1004_d 0.00113058f $X=7.56 $Y=2.6 $X2=0
+ $Y2=0
cc_684 N_A_987_409#_c_681_p N_VPWR_M1005_d 0.0188519f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_685 N_A_987_409#_c_671_n N_VPWR_c_1856_n 0.0385131f $X=5.075 $Y=2.475 $X2=0
+ $Y2=0
cc_686 N_A_987_409#_c_673_n N_VPWR_c_1856_n 0.0119061f $X=5.24 $Y=2.98 $X2=0
+ $Y2=0
cc_687 N_A_987_409#_c_684_p N_VPWR_c_1857_n 0.0138719f $X=7.39 $Y=2.98 $X2=0
+ $Y2=0
cc_688 N_A_987_409#_c_685_p N_VPWR_c_1857_n 0.00216246f $X=7.475 $Y=2.895 $X2=0
+ $Y2=0
cc_689 N_A_987_409#_c_681_p N_VPWR_c_1857_n 0.019543f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_690 N_A_987_409#_c_681_p N_VPWR_c_1858_n 0.0110845f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_691 N_A_987_409#_c_681_p N_VPWR_c_1859_n 0.019543f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_692 N_A_987_409#_M1035_g N_VPWR_c_1860_n 0.00350452f $X=10.84 $Y=2.595 $X2=0
+ $Y2=0
cc_693 N_A_987_409#_M1008_g N_VPWR_c_1866_n 0.00599878f $X=5.88 $Y=2.595 $X2=0
+ $Y2=0
cc_694 N_A_987_409#_c_672_n N_VPWR_c_1866_n 0.0412372f $X=5.96 $Y=2.98 $X2=0
+ $Y2=0
cc_695 N_A_987_409#_c_673_n N_VPWR_c_1866_n 0.0221635f $X=5.24 $Y=2.98 $X2=0
+ $Y2=0
cc_696 N_A_987_409#_c_684_p N_VPWR_c_1866_n 0.078901f $X=7.39 $Y=2.98 $X2=0
+ $Y2=0
cc_697 N_A_987_409#_c_681_p N_VPWR_c_1866_n 0.00305828f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_698 N_A_987_409#_c_695_p N_VPWR_c_1866_n 0.00921724f $X=6.045 $Y=2.98 $X2=0
+ $Y2=0
cc_699 N_A_987_409#_M1035_g N_VPWR_c_1867_n 0.00975641f $X=10.84 $Y=2.595 $X2=0
+ $Y2=0
cc_700 N_A_987_409#_c_681_p N_VPWR_c_1867_n 0.0130784f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_701 N_A_987_409#_M1008_g N_VPWR_c_1853_n 0.0100086f $X=5.88 $Y=2.595 $X2=0
+ $Y2=0
cc_702 N_A_987_409#_M1035_g N_VPWR_c_1853_n 0.0179933f $X=10.84 $Y=2.595 $X2=0
+ $Y2=0
cc_703 N_A_987_409#_c_672_n N_VPWR_c_1853_n 0.0259624f $X=5.96 $Y=2.98 $X2=0
+ $Y2=0
cc_704 N_A_987_409#_c_673_n N_VPWR_c_1853_n 0.0126536f $X=5.24 $Y=2.98 $X2=0
+ $Y2=0
cc_705 N_A_987_409#_c_684_p N_VPWR_c_1853_n 0.0513336f $X=7.39 $Y=2.98 $X2=0
+ $Y2=0
cc_706 N_A_987_409#_c_681_p N_VPWR_c_1853_n 0.0491788f $X=9.815 $Y=2.6 $X2=0
+ $Y2=0
cc_707 N_A_987_409#_c_695_p N_VPWR_c_1853_n 0.00636028f $X=6.045 $Y=2.98 $X2=0
+ $Y2=0
cc_708 N_A_987_409#_c_672_n N_A_352_409#_M1008_s 0.00534965f $X=5.96 $Y=2.98
+ $X2=0 $Y2=0
cc_709 N_A_987_409#_c_657_n N_A_352_409#_c_2083_n 0.00313309f $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_710 N_A_987_409#_c_663_n N_A_352_409#_c_2083_n 0.0154314f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_711 N_A_987_409#_c_663_n N_A_352_409#_c_2084_n 0.0317334f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_712 N_A_987_409#_M1008_g N_A_352_409#_c_2093_n 0.0140272f $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_713 N_A_987_409#_c_671_n N_A_352_409#_c_2093_n 0.0290823f $X=5.075 $Y=2.475
+ $X2=0 $Y2=0
cc_714 N_A_987_409#_c_672_n N_A_352_409#_c_2093_n 0.0196499f $X=5.96 $Y=2.98
+ $X2=0 $Y2=0
cc_715 N_A_987_409#_M1018_g N_A_352_409#_c_2086_n 5.96497e-19 $X=6.83 $Y=0.835
+ $X2=0 $Y2=0
cc_716 N_A_987_409#_c_663_n N_A_352_409#_c_2086_n 0.0190233f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_717 N_A_987_409#_c_665_n N_A_352_409#_c_2086_n 0.0108641f $X=6.13 $Y=1.54
+ $X2=0 $Y2=0
cc_718 N_A_987_409#_c_657_n N_A_352_409#_c_2088_n 0.0117982f $X=5.755 $Y=1.3
+ $X2=0 $Y2=0
cc_719 N_A_987_409#_c_663_n N_A_352_409#_c_2088_n 0.0100256f $X=5.755 $Y=0.81
+ $X2=0 $Y2=0
cc_720 N_A_987_409#_c_665_n N_A_352_409#_c_2088_n 0.00472989f $X=6.13 $Y=1.54
+ $X2=0 $Y2=0
cc_721 N_A_987_409#_M1008_g N_A_352_409#_c_2089_n 0.00272709f $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_722 N_A_987_409#_c_674_n N_A_352_409#_c_2089_n 0.00597942f $X=6.045 $Y=2.895
+ $X2=0 $Y2=0
cc_723 N_A_987_409#_c_664_n N_A_352_409#_c_2089_n 0.00127551f $X=5.84 $Y=1.615
+ $X2=0 $Y2=0
cc_724 N_A_987_409#_c_665_n N_A_352_409#_c_2089_n 0.0339659f $X=6.13 $Y=1.54
+ $X2=0 $Y2=0
cc_725 N_A_987_409#_M1008_g N_A_352_409#_c_2095_n 0.00691144f $X=5.88 $Y=2.595
+ $X2=0 $Y2=0
cc_726 N_A_987_409#_c_674_n N_A_352_409#_c_2095_n 0.0517827f $X=6.045 $Y=2.895
+ $X2=0 $Y2=0
cc_727 N_A_987_409#_c_664_n N_A_352_409#_c_2095_n 0.00185447f $X=5.84 $Y=1.615
+ $X2=0 $Y2=0
cc_728 N_A_987_409#_c_665_n N_A_352_409#_c_2095_n 0.00894917f $X=6.13 $Y=1.54
+ $X2=0 $Y2=0
cc_729 N_A_987_409#_c_684_p A_1373_419# 0.00497901f $X=7.39 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_730 N_A_987_409#_c_681_p A_1921_419# 0.00702693f $X=9.815 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_731 N_A_987_409#_M1018_g N_VGND_c_2353_n 9.49986e-19 $X=6.83 $Y=0.835 $X2=0
+ $Y2=0
cc_732 N_A_987_409#_c_668_n N_VGND_c_2353_n 9.49986e-19 $X=9.98 $Y=1.155 $X2=0
+ $Y2=0
cc_733 N_A_1423_99#_M1004_g N_A_1201_419#_M1026_g 0.0158161f $X=7.27 $Y=2.595
+ $X2=0 $Y2=0
cc_734 N_A_1423_99#_c_869_n N_A_1201_419#_M1026_g 0.00433088f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_735 N_A_1423_99#_c_878_n N_A_1201_419#_M1026_g 0.0179387f $X=8.435 $Y=2.25
+ $X2=0 $Y2=0
cc_736 N_A_1423_99#_c_871_n N_A_1201_419#_c_950_n 0.00397756f $X=8.095 $Y=1.31
+ $X2=0 $Y2=0
cc_737 N_A_1423_99#_c_873_n N_A_1201_419#_c_950_n 0.00391855f $X=8.18 $Y=1.225
+ $X2=0 $Y2=0
cc_738 N_A_1423_99#_c_874_n N_A_1201_419#_c_950_n 0.00633505f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_739 N_A_1423_99#_c_873_n N_A_1201_419#_c_951_n 0.00283292f $X=8.18 $Y=1.225
+ $X2=0 $Y2=0
cc_740 N_A_1423_99#_c_874_n N_A_1201_419#_c_951_n 0.00508231f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_741 N_A_1423_99#_M1004_g N_A_1201_419#_c_992_n 0.00201989f $X=7.27 $Y=2.595
+ $X2=0 $Y2=0
cc_742 N_A_1423_99#_M1004_g N_A_1201_419#_c_973_n 0.00860303f $X=7.27 $Y=2.595
+ $X2=0 $Y2=0
cc_743 N_A_1423_99#_c_869_n N_A_1201_419#_c_973_n 7.633e-19 $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_744 N_A_1423_99#_c_888_n N_A_1201_419#_c_973_n 0.00686956f $X=7.765 $Y=2.21
+ $X2=0 $Y2=0
cc_745 N_A_1423_99#_M1011_g N_A_1201_419#_c_954_n 0.0151046f $X=7.19 $Y=0.835
+ $X2=0 $Y2=0
cc_746 N_A_1423_99#_M1004_g N_A_1201_419#_c_954_n 0.00595154f $X=7.27 $Y=2.595
+ $X2=0 $Y2=0
cc_747 N_A_1423_99#_c_869_n N_A_1201_419#_c_954_n 0.0476903f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_748 N_A_1423_99#_c_870_n N_A_1201_419#_c_954_n 0.0129121f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_749 N_A_1423_99#_c_872_n N_A_1201_419#_c_954_n 0.01314f $X=7.765 $Y=1.31
+ $X2=0 $Y2=0
cc_750 N_A_1423_99#_M1011_g N_A_1201_419#_c_955_n 0.0046703f $X=7.19 $Y=0.835
+ $X2=0 $Y2=0
cc_751 N_A_1423_99#_c_870_n N_A_1201_419#_c_955_n 0.00558962f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_752 N_A_1423_99#_c_871_n N_A_1201_419#_c_955_n 0.0121295f $X=8.095 $Y=1.31
+ $X2=0 $Y2=0
cc_753 N_A_1423_99#_c_872_n N_A_1201_419#_c_955_n 0.0266476f $X=7.765 $Y=1.31
+ $X2=0 $Y2=0
cc_754 N_A_1423_99#_c_873_n N_A_1201_419#_c_955_n 0.00202762f $X=8.18 $Y=1.225
+ $X2=0 $Y2=0
cc_755 N_A_1423_99#_c_874_n N_A_1201_419#_c_955_n 0.0125113f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_756 N_A_1423_99#_M1011_g N_A_1201_419#_c_956_n 0.00469758f $X=7.19 $Y=0.835
+ $X2=0 $Y2=0
cc_757 N_A_1423_99#_c_874_n N_A_1201_419#_c_956_n 0.0201782f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_758 N_A_1423_99#_c_874_n N_A_1201_419#_c_957_n 0.0306148f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_759 N_A_1423_99#_c_869_n N_A_1201_419#_c_959_n 0.0199475f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_760 N_A_1423_99#_c_870_n N_A_1201_419#_c_959_n 0.00110518f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_761 N_A_1423_99#_c_871_n N_A_1201_419#_c_959_n 0.0191949f $X=8.095 $Y=1.31
+ $X2=0 $Y2=0
cc_762 N_A_1423_99#_c_878_n N_A_1201_419#_c_959_n 0.0445136f $X=8.435 $Y=2.25
+ $X2=0 $Y2=0
cc_763 N_A_1423_99#_c_874_n N_A_1201_419#_c_959_n 0.00596349f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_764 N_A_1423_99#_M1004_g N_A_1201_419#_c_960_n 7.90626e-19 $X=7.27 $Y=2.595
+ $X2=0 $Y2=0
cc_765 N_A_1423_99#_c_869_n N_A_1201_419#_c_960_n 6.23797e-19 $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_766 N_A_1423_99#_c_870_n N_A_1201_419#_c_960_n 0.0148975f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_767 N_A_1423_99#_c_871_n N_A_1201_419#_c_960_n 0.00459618f $X=8.095 $Y=1.31
+ $X2=0 $Y2=0
cc_768 N_A_1423_99#_c_878_n N_A_1201_419#_c_960_n 0.00195488f $X=8.435 $Y=2.25
+ $X2=0 $Y2=0
cc_769 N_A_1423_99#_c_871_n N_A_1201_419#_c_961_n 0.00191269f $X=8.095 $Y=1.31
+ $X2=0 $Y2=0
cc_770 N_A_1423_99#_c_873_n N_A_1201_419#_c_962_n 0.00634916f $X=8.18 $Y=1.225
+ $X2=0 $Y2=0
cc_771 N_A_1423_99#_c_874_n N_A_1201_419#_c_962_n 0.0153823f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_772 N_A_1423_99#_c_871_n N_A_1201_419#_c_964_n 0.0118646f $X=8.095 $Y=1.31
+ $X2=0 $Y2=0
cc_773 N_A_1423_99#_c_873_n N_A_1201_419#_c_964_n 0.0017133f $X=8.18 $Y=1.225
+ $X2=0 $Y2=0
cc_774 N_A_1423_99#_c_874_n N_A_1201_419#_c_964_n 0.00332007f $X=8.355 $Y=0.815
+ $X2=0 $Y2=0
cc_775 N_A_1423_99#_M1011_g N_A_1201_419#_c_965_n 0.00125843f $X=7.19 $Y=0.835
+ $X2=0 $Y2=0
cc_776 N_A_1423_99#_M1011_g N_A_1201_419#_c_1062_n 0.00690009f $X=7.19 $Y=0.835
+ $X2=0 $Y2=0
cc_777 N_A_1423_99#_c_869_n N_A_1201_419#_c_968_n 0.00362518f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_778 N_A_1423_99#_c_870_n N_A_1201_419#_c_968_n 0.00183234f $X=7.6 $Y=1.675
+ $X2=0 $Y2=0
cc_779 N_A_1423_99#_c_871_n N_A_1201_419#_c_968_n 0.00438268f $X=8.095 $Y=1.31
+ $X2=0 $Y2=0
cc_780 N_A_1423_99#_c_878_n N_SET_B_M1005_g 0.0127902f $X=8.435 $Y=2.25 $X2=0
+ $Y2=0
cc_781 N_A_1423_99#_M1004_g N_A_761_113#_c_1298_n 0.0643022f $X=7.27 $Y=2.595
+ $X2=0 $Y2=0
cc_782 N_A_1423_99#_M1011_g N_A_761_113#_c_1284_n 0.00866183f $X=7.19 $Y=0.835
+ $X2=0 $Y2=0
cc_783 N_A_1423_99#_c_888_n N_VPWR_M1004_d 0.00771208f $X=7.765 $Y=2.21 $X2=0
+ $Y2=0
cc_784 N_A_1423_99#_c_878_n N_VPWR_M1004_d 0.00376162f $X=8.435 $Y=2.25 $X2=0
+ $Y2=0
cc_785 N_A_1423_99#_M1004_g N_VPWR_c_1857_n 0.00309907f $X=7.27 $Y=2.595 $X2=0
+ $Y2=0
cc_786 N_A_1423_99#_M1004_g N_VPWR_c_1866_n 0.00599934f $X=7.27 $Y=2.595 $X2=0
+ $Y2=0
cc_787 N_A_1423_99#_M1026_d N_VPWR_c_1853_n 0.00329651f $X=8.295 $Y=2.095 $X2=0
+ $Y2=0
cc_788 N_A_1423_99#_M1004_g N_VPWR_c_1853_n 0.0086712f $X=7.27 $Y=2.595 $X2=0
+ $Y2=0
cc_789 N_A_1423_99#_M1011_g N_VGND_c_2338_n 0.0063844f $X=7.19 $Y=0.835 $X2=0
+ $Y2=0
cc_790 N_A_1423_99#_M1011_g N_VGND_c_2353_n 9.49986e-19 $X=7.19 $Y=0.835 $X2=0
+ $Y2=0
cc_791 N_A_1201_419#_M1026_g N_SET_B_M1005_g 0.0489488f $X=8.17 $Y=2.595 $X2=0
+ $Y2=0
cc_792 N_A_1201_419#_M1025_g N_SET_B_M1005_g 0.0307071f $X=9.48 $Y=2.595 $X2=0
+ $Y2=0
cc_793 N_A_1201_419#_c_959_n N_SET_B_M1005_g 0.00215524f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_794 N_A_1201_419#_c_960_n N_SET_B_M1005_g 0.0096933f $X=8.17 $Y=1.74 $X2=0
+ $Y2=0
cc_795 N_A_1201_419#_c_951_n N_SET_B_M1037_g 0.0367242f $X=8.57 $Y=1.16 $X2=0
+ $Y2=0
cc_796 N_A_1201_419#_M1002_g N_SET_B_M1037_g 0.0130154f $X=9.5 $Y=0.835 $X2=0
+ $Y2=0
cc_797 N_A_1201_419#_c_961_n N_SET_B_M1037_g 0.00194401f $X=8.53 $Y=1.575 $X2=0
+ $Y2=0
cc_798 N_A_1201_419#_c_962_n N_SET_B_M1037_g 0.00639012f $X=8.785 $Y=1.2 $X2=0
+ $Y2=0
cc_799 N_A_1201_419#_c_963_n N_SET_B_M1037_g 0.0148626f $X=9.275 $Y=1.285 $X2=0
+ $Y2=0
cc_800 N_A_1201_419#_c_966_n N_SET_B_M1037_g 7.2647e-19 $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_801 N_A_1201_419#_c_967_n N_SET_B_M1037_g 0.018824f $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_802 N_A_1201_419#_c_968_n N_SET_B_M1037_g 0.00320945f $X=8.17 $Y=1.575 $X2=0
+ $Y2=0
cc_803 N_A_1201_419#_c_953_n N_SET_B_c_1151_n 0.00232868f $X=9.44 $Y=1.705 $X2=0
+ $Y2=0
cc_804 N_A_1201_419#_c_972_n N_SET_B_c_1151_n 5.32754e-19 $X=9.44 $Y=1.87 $X2=0
+ $Y2=0
cc_805 N_A_1201_419#_c_963_n N_SET_B_c_1151_n 0.00928499f $X=9.275 $Y=1.285
+ $X2=0 $Y2=0
cc_806 N_A_1201_419#_c_966_n N_SET_B_c_1151_n 0.0355884f $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_807 N_A_1201_419#_c_959_n N_SET_B_c_1152_n 0.00618466f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_808 N_A_1201_419#_c_961_n N_SET_B_c_1152_n 6.47208e-19 $X=8.53 $Y=1.575 $X2=0
+ $Y2=0
cc_809 N_A_1201_419#_c_964_n N_SET_B_c_1152_n 0.004311f $X=8.87 $Y=1.285 $X2=0
+ $Y2=0
cc_810 N_A_1201_419#_c_966_n N_SET_B_c_1152_n 5.88013e-19 $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_811 N_A_1201_419#_c_953_n N_SET_B_c_1153_n 0.00109422f $X=9.44 $Y=1.705 $X2=0
+ $Y2=0
cc_812 N_A_1201_419#_c_959_n N_SET_B_c_1153_n 0.0200517f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_813 N_A_1201_419#_c_960_n N_SET_B_c_1153_n 2.64093e-19 $X=8.17 $Y=1.74 $X2=0
+ $Y2=0
cc_814 N_A_1201_419#_c_961_n N_SET_B_c_1153_n 0.00136625f $X=8.53 $Y=1.575 $X2=0
+ $Y2=0
cc_815 N_A_1201_419#_c_964_n N_SET_B_c_1153_n 0.0157687f $X=8.87 $Y=1.285 $X2=0
+ $Y2=0
cc_816 N_A_1201_419#_c_966_n N_SET_B_c_1153_n 0.0178208f $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_817 N_A_1201_419#_c_949_n N_SET_B_c_1155_n 0.00390359f $X=8.495 $Y=1.235
+ $X2=0 $Y2=0
cc_818 N_A_1201_419#_M1025_g N_SET_B_c_1155_n 4.71348e-19 $X=9.48 $Y=2.595 $X2=0
+ $Y2=0
cc_819 N_A_1201_419#_c_953_n N_SET_B_c_1155_n 0.0212605f $X=9.44 $Y=1.705 $X2=0
+ $Y2=0
cc_820 N_A_1201_419#_c_959_n N_SET_B_c_1155_n 0.00857431f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_821 N_A_1201_419#_c_961_n N_SET_B_c_1155_n 8.22677e-19 $X=8.53 $Y=1.575 $X2=0
+ $Y2=0
cc_822 N_A_1201_419#_c_963_n N_SET_B_c_1155_n 2.01906e-19 $X=9.275 $Y=1.285
+ $X2=0 $Y2=0
cc_823 N_A_1201_419#_c_964_n N_SET_B_c_1155_n 0.00702384f $X=8.87 $Y=1.285 $X2=0
+ $Y2=0
cc_824 N_A_1201_419#_c_966_n N_SET_B_c_1155_n 0.00116218f $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_825 N_A_1201_419#_c_968_n N_SET_B_c_1155_n 0.0096933f $X=8.17 $Y=1.575 $X2=0
+ $Y2=0
cc_826 N_A_1201_419#_c_965_n N_A_761_113#_M1043_g 0.00444953f $X=6.615 $Y=0.835
+ $X2=0 $Y2=0
cc_827 N_A_1201_419#_c_954_n N_A_761_113#_c_1298_n 0.00417154f $X=7.17 $Y=2.075
+ $X2=0 $Y2=0
cc_828 N_A_1201_419#_c_974_n N_A_761_113#_c_1299_n 0.00892503f $X=6.64 $Y=2.16
+ $X2=0 $Y2=0
cc_829 N_A_1201_419#_c_951_n N_A_761_113#_c_1284_n 0.00737233f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_830 N_A_1201_419#_M1002_g N_A_761_113#_c_1284_n 0.00907339f $X=9.5 $Y=0.835
+ $X2=0 $Y2=0
cc_831 N_A_1201_419#_c_1001_n N_A_761_113#_c_1284_n 0.0033529f $X=7.085 $Y=0.96
+ $X2=0 $Y2=0
cc_832 N_A_1201_419#_c_955_n N_A_761_113#_c_1284_n 0.00462744f $X=7.745 $Y=0.96
+ $X2=0 $Y2=0
cc_833 N_A_1201_419#_c_957_n N_A_761_113#_c_1284_n 0.0201004f $X=8.7 $Y=0.35
+ $X2=0 $Y2=0
cc_834 N_A_1201_419#_c_958_n N_A_761_113#_c_1284_n 0.00418768f $X=7.915 $Y=0.35
+ $X2=0 $Y2=0
cc_835 N_A_1201_419#_c_965_n N_A_761_113#_c_1284_n 0.00527611f $X=6.615 $Y=0.835
+ $X2=0 $Y2=0
cc_836 N_A_1201_419#_c_1062_n N_A_761_113#_c_1284_n 4.39455e-19 $X=7.17 $Y=0.96
+ $X2=0 $Y2=0
cc_837 N_A_1201_419#_c_992_n N_A_761_113#_c_1300_n 0.011874f $X=6.475 $Y=2.395
+ $X2=0 $Y2=0
cc_838 N_A_1201_419#_c_973_n N_A_761_113#_c_1300_n 0.0153824f $X=7.085 $Y=2.16
+ $X2=0 $Y2=0
cc_839 N_A_1201_419#_c_974_n N_A_761_113#_c_1300_n 0.00277341f $X=6.64 $Y=2.16
+ $X2=0 $Y2=0
cc_840 N_A_1201_419#_M1025_g N_A_761_113#_M1000_g 0.0415468f $X=9.48 $Y=2.595
+ $X2=0 $Y2=0
cc_841 N_A_1201_419#_c_972_n N_A_761_113#_c_1303_n 0.0415468f $X=9.44 $Y=1.87
+ $X2=0 $Y2=0
cc_842 N_A_1201_419#_M1026_g N_VPWR_c_1857_n 0.0105816f $X=8.17 $Y=2.595 $X2=0
+ $Y2=0
cc_843 N_A_1201_419#_M1026_g N_VPWR_c_1858_n 0.00639129f $X=8.17 $Y=2.595 $X2=0
+ $Y2=0
cc_844 N_A_1201_419#_M1026_g N_VPWR_c_1859_n 0.00184932f $X=8.17 $Y=2.595 $X2=0
+ $Y2=0
cc_845 N_A_1201_419#_M1025_g N_VPWR_c_1859_n 0.00795191f $X=9.48 $Y=2.595 $X2=0
+ $Y2=0
cc_846 N_A_1201_419#_M1025_g N_VPWR_c_1867_n 0.00710941f $X=9.48 $Y=2.595 $X2=0
+ $Y2=0
cc_847 N_A_1201_419#_M1008_d N_VPWR_c_1853_n 0.00499582f $X=6.005 $Y=2.095 $X2=0
+ $Y2=0
cc_848 N_A_1201_419#_M1026_g N_VPWR_c_1853_n 0.00713465f $X=8.17 $Y=2.595 $X2=0
+ $Y2=0
cc_849 N_A_1201_419#_M1025_g N_VPWR_c_1853_n 0.0094236f $X=9.48 $Y=2.595 $X2=0
+ $Y2=0
cc_850 N_A_1201_419#_c_965_n N_A_352_409#_c_2086_n 0.00934633f $X=6.615 $Y=0.835
+ $X2=0 $Y2=0
cc_851 N_A_1201_419#_c_973_n A_1373_419# 0.00336478f $X=7.085 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_852 N_A_1201_419#_c_955_n N_VGND_M1011_d 0.00862469f $X=7.745 $Y=0.96 $X2=0
+ $Y2=0
cc_853 N_A_1201_419#_c_955_n N_VGND_c_2338_n 0.0188647f $X=7.745 $Y=0.96 $X2=0
+ $Y2=0
cc_854 N_A_1201_419#_c_956_n N_VGND_c_2338_n 0.0189539f $X=7.83 $Y=0.875 $X2=0
+ $Y2=0
cc_855 N_A_1201_419#_c_958_n N_VGND_c_2338_n 0.0140867f $X=7.915 $Y=0.35 $X2=0
+ $Y2=0
cc_856 N_A_1201_419#_c_965_n N_VGND_c_2338_n 0.00165761f $X=6.615 $Y=0.835 $X2=0
+ $Y2=0
cc_857 N_A_1201_419#_M1002_g N_VGND_c_2339_n 0.00598495f $X=9.5 $Y=0.835 $X2=0
+ $Y2=0
cc_858 N_A_1201_419#_c_957_n N_VGND_c_2339_n 0.0144411f $X=8.7 $Y=0.35 $X2=0
+ $Y2=0
cc_859 N_A_1201_419#_c_962_n N_VGND_c_2339_n 0.0143489f $X=8.785 $Y=1.2 $X2=0
+ $Y2=0
cc_860 N_A_1201_419#_c_963_n N_VGND_c_2339_n 0.0154758f $X=9.275 $Y=1.285 $X2=0
+ $Y2=0
cc_861 N_A_1201_419#_c_966_n N_VGND_c_2339_n 0.00796253f $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_862 N_A_1201_419#_c_967_n N_VGND_c_2339_n 7.7371e-19 $X=9.44 $Y=1.365 $X2=0
+ $Y2=0
cc_863 N_A_1201_419#_c_965_n N_VGND_c_2347_n 0.00662562f $X=6.615 $Y=0.835 $X2=0
+ $Y2=0
cc_864 N_A_1201_419#_c_957_n N_VGND_c_2348_n 0.0589829f $X=8.7 $Y=0.35 $X2=0
+ $Y2=0
cc_865 N_A_1201_419#_c_958_n N_VGND_c_2348_n 0.0114574f $X=7.915 $Y=0.35 $X2=0
+ $Y2=0
cc_866 N_A_1201_419#_M1002_g N_VGND_c_2353_n 9.49986e-19 $X=9.5 $Y=0.835 $X2=0
+ $Y2=0
cc_867 N_A_1201_419#_c_957_n N_VGND_c_2353_n 0.032098f $X=8.7 $Y=0.35 $X2=0
+ $Y2=0
cc_868 N_A_1201_419#_c_958_n N_VGND_c_2353_n 0.00589978f $X=7.915 $Y=0.35 $X2=0
+ $Y2=0
cc_869 N_A_1201_419#_c_965_n N_VGND_c_2353_n 0.00866864f $X=6.615 $Y=0.835 $X2=0
+ $Y2=0
cc_870 N_A_1201_419#_c_1001_n A_1381_125# 0.00529857f $X=7.085 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_871 N_A_1201_419#_c_962_n A_1729_125# 0.00276176f $X=8.785 $Y=1.2 $X2=-0.19
+ $Y2=-0.245
cc_872 N_SET_B_M1037_g N_A_761_113#_c_1284_n 0.00907339f $X=8.96 $Y=0.835 $X2=0
+ $Y2=0
cc_873 N_SET_B_c_1151_n N_A_761_113#_c_1286_n 0.00205714f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_874 N_SET_B_c_1151_n N_A_761_113#_c_1287_n 0.00616986f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_875 N_SET_B_c_1148_n N_A_2220_40#_M1029_g 0.0486362f $X=11.54 $Y=0.825 $X2=0
+ $Y2=0
cc_876 N_SET_B_c_1150_n N_A_2220_40#_c_1488_n 0.0172822f $X=11.615 $Y=0.9 $X2=0
+ $Y2=0
cc_877 N_SET_B_c_1151_n N_A_2220_40#_c_1488_n 0.0102798f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_878 N_SET_B_c_1157_n N_A_2220_40#_c_1488_n 0.00122707f $X=12.15 $Y=1.725
+ $X2=0 $Y2=0
cc_879 N_SET_B_c_1158_n N_A_2220_40#_c_1488_n 0.0443147f $X=12.15 $Y=1.56 $X2=0
+ $Y2=0
cc_880 N_SET_B_c_1156_n N_A_2220_40#_M1021_g 0.0254547f $X=12.15 $Y=1.725 $X2=0
+ $Y2=0
cc_881 N_SET_B_c_1151_n N_A_2220_40#_c_1496_n 0.0178437f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_882 SET_B N_A_2220_40#_c_1496_n 4.85279e-19 $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_883 N_SET_B_c_1157_n N_A_2220_40#_c_1496_n 0.0189633f $X=12.15 $Y=1.725 $X2=0
+ $Y2=0
cc_884 N_SET_B_c_1158_n N_A_2220_40#_c_1496_n 0.00172347f $X=12.15 $Y=1.56 $X2=0
+ $Y2=0
cc_885 N_SET_B_c_1149_n N_A_2220_40#_c_1489_n 0.00505022f $X=11.985 $Y=0.9 $X2=0
+ $Y2=0
cc_886 N_SET_B_c_1151_n N_A_2220_40#_c_1489_n 0.00970372f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_887 SET_B N_A_2220_40#_c_1489_n 0.00834942f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_888 N_SET_B_c_1156_n N_A_2220_40#_c_1489_n 0.0012094f $X=12.15 $Y=1.725 $X2=0
+ $Y2=0
cc_889 N_SET_B_c_1157_n N_A_2220_40#_c_1489_n 0.0229166f $X=12.15 $Y=1.725 $X2=0
+ $Y2=0
cc_890 N_SET_B_c_1158_n N_A_2220_40#_c_1489_n 0.014828f $X=12.15 $Y=1.56 $X2=0
+ $Y2=0
cc_891 N_SET_B_c_1150_n N_A_2220_40#_c_1490_n 0.00377533f $X=11.615 $Y=0.9 $X2=0
+ $Y2=0
cc_892 N_SET_B_c_1148_n N_A_2220_40#_c_1491_n 0.00251281f $X=11.54 $Y=0.825
+ $X2=0 $Y2=0
cc_893 N_SET_B_c_1149_n N_A_2220_40#_c_1491_n 0.0110799f $X=11.985 $Y=0.9 $X2=0
+ $Y2=0
cc_894 N_SET_B_M1027_g N_A_2220_40#_c_1497_n 0.00192995f $X=12.11 $Y=2.595 $X2=0
+ $Y2=0
cc_895 N_SET_B_M1027_g N_A_2220_40#_c_1493_n 0.00536067f $X=12.11 $Y=2.595 $X2=0
+ $Y2=0
cc_896 SET_B N_A_2220_40#_c_1493_n 0.00696049f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_897 N_SET_B_c_1156_n N_A_2220_40#_c_1493_n 0.00128137f $X=12.15 $Y=1.725
+ $X2=0 $Y2=0
cc_898 N_SET_B_c_1157_n N_A_2220_40#_c_1493_n 0.0151755f $X=12.15 $Y=1.725 $X2=0
+ $Y2=0
cc_899 N_SET_B_c_1158_n N_A_2220_40#_c_1493_n 0.00295925f $X=12.15 $Y=1.56 $X2=0
+ $Y2=0
cc_900 N_SET_B_c_1149_n N_A_2019_419#_M1013_g 0.0082552f $X=11.985 $Y=0.9 $X2=0
+ $Y2=0
cc_901 N_SET_B_c_1158_n N_A_2019_419#_c_1576_n 0.0082552f $X=12.15 $Y=1.56 $X2=0
+ $Y2=0
cc_902 N_SET_B_c_1151_n N_A_2019_419#_c_1609_n 0.00881833f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_903 N_SET_B_c_1150_n N_A_2019_419#_c_1593_n 7.27547e-19 $X=11.615 $Y=0.9
+ $X2=0 $Y2=0
cc_904 N_SET_B_c_1151_n N_A_2019_419#_c_1593_n 0.0125971f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_905 N_SET_B_c_1158_n N_A_2019_419#_c_1593_n 0.00360267f $X=12.15 $Y=1.56
+ $X2=0 $Y2=0
cc_906 N_SET_B_c_1151_n N_A_2019_419#_c_1594_n 0.00688932f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_907 N_SET_B_c_1151_n N_A_2019_419#_c_1595_n 0.0204771f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_908 N_SET_B_c_1156_n N_A_2019_419#_c_1595_n 0.00104215f $X=12.15 $Y=1.725
+ $X2=0 $Y2=0
cc_909 N_SET_B_c_1158_n N_A_2019_419#_c_1595_n 0.00178611f $X=12.15 $Y=1.56
+ $X2=0 $Y2=0
cc_910 N_SET_B_M1027_g N_A_2019_419#_c_1633_n 0.0197366f $X=12.11 $Y=2.595 $X2=0
+ $Y2=0
cc_911 N_SET_B_c_1151_n N_A_2019_419#_c_1633_n 0.015145f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_912 SET_B N_A_2019_419#_c_1633_n 6.03144e-19 $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_913 N_SET_B_c_1157_n N_A_2019_419#_c_1633_n 0.0116644f $X=12.15 $Y=1.725
+ $X2=0 $Y2=0
cc_914 N_SET_B_M1027_g N_A_2019_419#_c_1603_n 0.0020085f $X=12.11 $Y=2.595 $X2=0
+ $Y2=0
cc_915 SET_B N_A_2019_419#_c_1603_n 0.00239488f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_916 N_SET_B_c_1156_n N_A_2019_419#_c_1603_n 0.00184978f $X=12.15 $Y=1.725
+ $X2=0 $Y2=0
cc_917 N_SET_B_c_1157_n N_A_2019_419#_c_1603_n 0.0105389f $X=12.15 $Y=1.725
+ $X2=0 $Y2=0
cc_918 N_SET_B_M1027_g N_A_2019_419#_c_1641_n 0.0165497f $X=12.11 $Y=2.595 $X2=0
+ $Y2=0
cc_919 N_SET_B_M1027_g N_A_2019_419#_c_1642_n 0.00317906f $X=12.11 $Y=2.595
+ $X2=0 $Y2=0
cc_920 N_SET_B_c_1156_n N_A_2019_419#_c_1597_n 0.00484093f $X=12.15 $Y=1.725
+ $X2=0 $Y2=0
cc_921 N_SET_B_c_1158_n N_A_2019_419#_c_1597_n 0.00247486f $X=12.15 $Y=1.56
+ $X2=0 $Y2=0
cc_922 N_SET_B_c_1151_n N_A_2019_419#_c_1606_n 0.00256847f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_923 N_SET_B_M1005_g N_VPWR_c_1857_n 0.00184932f $X=8.7 $Y=2.595 $X2=0 $Y2=0
cc_924 N_SET_B_M1005_g N_VPWR_c_1858_n 0.00639129f $X=8.7 $Y=2.595 $X2=0 $Y2=0
cc_925 N_SET_B_M1005_g N_VPWR_c_1859_n 0.0103951f $X=8.7 $Y=2.595 $X2=0 $Y2=0
cc_926 N_SET_B_M1027_g N_VPWR_c_1860_n 0.0101241f $X=12.11 $Y=2.595 $X2=0 $Y2=0
cc_927 N_SET_B_M1027_g N_VPWR_c_1868_n 0.00938036f $X=12.11 $Y=2.595 $X2=0 $Y2=0
cc_928 N_SET_B_M1005_g N_VPWR_c_1853_n 0.00713465f $X=8.7 $Y=2.595 $X2=0 $Y2=0
cc_929 N_SET_B_M1027_g N_VPWR_c_1853_n 0.0179032f $X=12.11 $Y=2.595 $X2=0 $Y2=0
cc_930 N_SET_B_M1037_g N_VGND_c_2339_n 0.00135982f $X=8.96 $Y=0.835 $X2=0 $Y2=0
cc_931 N_SET_B_c_1151_n N_VGND_c_2339_n 4.14819e-19 $X=12.095 $Y=1.665 $X2=0
+ $Y2=0
cc_932 N_SET_B_c_1148_n N_VGND_c_2340_n 0.0145721f $X=11.54 $Y=0.825 $X2=0 $Y2=0
cc_933 N_SET_B_c_1149_n N_VGND_c_2340_n 0.00845669f $X=11.985 $Y=0.9 $X2=0 $Y2=0
cc_934 N_SET_B_c_1148_n N_VGND_c_2349_n 0.00411131f $X=11.54 $Y=0.825 $X2=0
+ $Y2=0
cc_935 N_SET_B_M1037_g N_VGND_c_2353_n 9.49986e-19 $X=8.96 $Y=0.835 $X2=0 $Y2=0
cc_936 N_SET_B_c_1148_n N_VGND_c_2353_n 0.00779341f $X=11.54 $Y=0.825 $X2=0
+ $Y2=0
cc_937 N_SET_B_c_1149_n N_VGND_c_2353_n 0.00521992f $X=11.985 $Y=0.9 $X2=0 $Y2=0
cc_938 N_A_761_113#_c_1284_n N_A_2220_40#_M1029_g 0.0332721f $X=10.71 $Y=0.18
+ $X2=0 $Y2=0
cc_939 N_A_761_113#_M1028_g N_A_2220_40#_c_1488_n 0.0332721f $X=10.785 $Y=0.54
+ $X2=0 $Y2=0
cc_940 N_A_761_113#_c_1284_n N_A_2019_419#_c_1592_n 0.00710251f $X=10.71 $Y=0.18
+ $X2=0 $Y2=0
cc_941 N_A_761_113#_M1028_g N_A_2019_419#_c_1592_n 0.0109782f $X=10.785 $Y=0.54
+ $X2=0 $Y2=0
cc_942 N_A_761_113#_c_1287_n N_A_2019_419#_c_1593_n 0.00133388f $X=10.71 $Y=1.29
+ $X2=0 $Y2=0
cc_943 N_A_761_113#_M1028_g N_A_2019_419#_c_1593_n 0.0160735f $X=10.785 $Y=0.54
+ $X2=0 $Y2=0
cc_944 N_A_761_113#_c_1288_n N_A_2019_419#_c_1594_n 0.00925811f $X=10.505
+ $Y=1.29 $X2=0 $Y2=0
cc_945 N_A_761_113#_c_1286_n N_A_2019_419#_c_1595_n 0.00487906f $X=10.43
+ $Y=1.725 $X2=0 $Y2=0
cc_946 N_A_761_113#_M1028_g N_A_2019_419#_c_1595_n 0.00158722f $X=10.785 $Y=0.54
+ $X2=0 $Y2=0
cc_947 N_A_761_113#_M1000_g N_A_2019_419#_c_1606_n 0.018646f $X=9.97 $Y=2.595
+ $X2=0 $Y2=0
cc_948 N_A_761_113#_c_1302_n N_A_2019_419#_c_1606_n 0.0073295f $X=10.355 $Y=1.8
+ $X2=0 $Y2=0
cc_949 N_A_761_113#_c_1307_n N_VPWR_M1047_d 0.00180746f $X=4.825 $Y=2.045 $X2=0
+ $Y2=0
cc_950 N_A_761_113#_M1034_g N_VPWR_c_1856_n 0.0189096f $X=4.81 $Y=2.545 $X2=0
+ $Y2=0
cc_951 N_A_761_113#_c_1305_n N_VPWR_c_1856_n 0.0497475f $X=4.015 $Y=2.19 $X2=0
+ $Y2=0
cc_952 N_A_761_113#_c_1307_n N_VPWR_c_1856_n 0.0163515f $X=4.825 $Y=2.045 $X2=0
+ $Y2=0
cc_953 N_A_761_113#_c_1305_n N_VPWR_c_1865_n 0.0220321f $X=4.015 $Y=2.19 $X2=0
+ $Y2=0
cc_954 N_A_761_113#_M1034_g N_VPWR_c_1866_n 0.00767656f $X=4.81 $Y=2.545 $X2=0
+ $Y2=0
cc_955 N_A_761_113#_c_1300_n N_VPWR_c_1866_n 0.00599941f $X=6.74 $Y=2.02 $X2=0
+ $Y2=0
cc_956 N_A_761_113#_M1000_g N_VPWR_c_1867_n 0.00827272f $X=9.97 $Y=2.595 $X2=0
+ $Y2=0
cc_957 N_A_761_113#_M1034_g N_VPWR_c_1853_n 0.014306f $X=4.81 $Y=2.545 $X2=0
+ $Y2=0
cc_958 N_A_761_113#_c_1300_n N_VPWR_c_1853_n 0.00861537f $X=6.74 $Y=2.02 $X2=0
+ $Y2=0
cc_959 N_A_761_113#_M1000_g N_VPWR_c_1853_n 0.0131771f $X=9.97 $Y=2.595 $X2=0
+ $Y2=0
cc_960 N_A_761_113#_c_1305_n N_VPWR_c_1853_n 0.0125808f $X=4.015 $Y=2.19 $X2=0
+ $Y2=0
cc_961 N_A_761_113#_c_1305_n N_A_245_409#_c_2025_n 0.0501419f $X=4.015 $Y=2.19
+ $X2=0 $Y2=0
cc_962 N_A_761_113#_c_1305_n N_A_352_409#_c_2090_n 2.78788e-19 $X=4.015 $Y=2.19
+ $X2=0 $Y2=0
cc_963 N_A_761_113#_c_1310_n N_A_352_409#_c_2090_n 0.0050211f $X=4.015 $Y=2.045
+ $X2=0 $Y2=0
cc_964 N_A_761_113#_c_1310_n N_A_352_409#_c_2075_n 2.76809e-19 $X=4.015 $Y=2.045
+ $X2=0 $Y2=0
cc_965 N_A_761_113#_c_1295_n N_A_352_409#_c_2076_n 0.0133765f $X=3.95 $Y=0.81
+ $X2=0 $Y2=0
cc_966 N_A_761_113#_c_1295_n N_A_352_409#_c_2077_n 0.0101504f $X=3.95 $Y=0.81
+ $X2=0 $Y2=0
cc_967 N_A_761_113#_c_1295_n N_A_352_409#_c_2078_n 0.0160399f $X=3.95 $Y=0.81
+ $X2=0 $Y2=0
cc_968 N_A_761_113#_c_1276_n N_A_352_409#_c_2080_n 6.99561e-19 $X=4.955 $Y=1.06
+ $X2=0 $Y2=0
cc_969 N_A_761_113#_c_1292_n N_A_352_409#_c_2080_n 0.00525652f $X=3.95 $Y=1.96
+ $X2=0 $Y2=0
cc_970 N_A_761_113#_c_1295_n N_A_352_409#_c_2080_n 0.0140824f $X=3.95 $Y=0.81
+ $X2=0 $Y2=0
cc_971 N_A_761_113#_c_1277_n N_A_352_409#_c_2081_n 0.0038277f $X=4.955 $Y=1.555
+ $X2=0 $Y2=0
cc_972 N_A_761_113#_c_1290_n N_A_352_409#_c_2081_n 0.00842211f $X=4.955 $Y=1.135
+ $X2=0 $Y2=0
cc_973 N_A_761_113#_c_1293_n N_A_352_409#_c_2081_n 0.00956149f $X=4.98 $Y=1.72
+ $X2=0 $Y2=0
cc_974 N_A_761_113#_c_1294_n N_A_352_409#_c_2081_n 0.00551261f $X=4.98 $Y=1.72
+ $X2=0 $Y2=0
cc_975 N_A_761_113#_c_1292_n N_A_352_409#_c_2082_n 0.0101592f $X=3.95 $Y=1.96
+ $X2=0 $Y2=0
cc_976 N_A_761_113#_c_1276_n N_A_352_409#_c_2083_n 0.0107945f $X=4.955 $Y=1.06
+ $X2=0 $Y2=0
cc_977 N_A_761_113#_c_1278_n N_A_352_409#_c_2083_n 0.00223445f $X=5.24 $Y=1.135
+ $X2=0 $Y2=0
cc_978 N_A_761_113#_c_1279_n N_A_352_409#_c_2083_n 0.00499645f $X=5.315 $Y=1.06
+ $X2=0 $Y2=0
cc_979 N_A_761_113#_c_1290_n N_A_352_409#_c_2083_n 6.70354e-19 $X=4.955 $Y=1.135
+ $X2=0 $Y2=0
cc_980 N_A_761_113#_c_1279_n N_A_352_409#_c_2084_n 0.00706035f $X=5.315 $Y=1.06
+ $X2=0 $Y2=0
cc_981 N_A_761_113#_c_1280_n N_A_352_409#_c_2084_n 0.00384822f $X=6.215 $Y=1.135
+ $X2=0 $Y2=0
cc_982 N_A_761_113#_M1043_g N_A_352_409#_c_2084_n 0.0122097f $X=6.32 $Y=0.625
+ $X2=0 $Y2=0
cc_983 N_A_761_113#_c_1276_n N_A_352_409#_c_2085_n 2.48962e-19 $X=4.955 $Y=1.06
+ $X2=0 $Y2=0
cc_984 N_A_761_113#_M1034_g N_A_352_409#_c_2093_n 0.0052504f $X=4.81 $Y=2.545
+ $X2=0 $Y2=0
cc_985 N_A_761_113#_c_1279_n N_A_352_409#_c_2086_n 0.00399822f $X=5.315 $Y=1.06
+ $X2=0 $Y2=0
cc_986 N_A_761_113#_c_1280_n N_A_352_409#_c_2086_n 0.00501084f $X=6.215 $Y=1.135
+ $X2=0 $Y2=0
cc_987 N_A_761_113#_c_1281_n N_A_352_409#_c_2086_n 0.00107968f $X=6.29 $Y=1.21
+ $X2=0 $Y2=0
cc_988 N_A_761_113#_M1043_g N_A_352_409#_c_2086_n 0.00842726f $X=6.32 $Y=0.625
+ $X2=0 $Y2=0
cc_989 N_A_761_113#_c_1277_n N_A_352_409#_c_2088_n 0.00512935f $X=4.955 $Y=1.555
+ $X2=0 $Y2=0
cc_990 N_A_761_113#_c_1278_n N_A_352_409#_c_2088_n 0.00815679f $X=5.24 $Y=1.135
+ $X2=0 $Y2=0
cc_991 N_A_761_113#_c_1280_n N_A_352_409#_c_2088_n 0.00385197f $X=6.215 $Y=1.135
+ $X2=0 $Y2=0
cc_992 N_A_761_113#_c_1291_n N_A_352_409#_c_2088_n 0.00974583f $X=5.315 $Y=1.135
+ $X2=0 $Y2=0
cc_993 N_A_761_113#_c_1293_n N_A_352_409#_c_2088_n 0.00958947f $X=4.98 $Y=1.72
+ $X2=0 $Y2=0
cc_994 N_A_761_113#_c_1294_n N_A_352_409#_c_2088_n 9.48313e-19 $X=4.98 $Y=1.72
+ $X2=0 $Y2=0
cc_995 N_A_761_113#_M1034_g N_A_352_409#_c_2089_n 0.00114776f $X=4.81 $Y=2.545
+ $X2=0 $Y2=0
cc_996 N_A_761_113#_c_1277_n N_A_352_409#_c_2089_n 0.00402544f $X=4.955 $Y=1.555
+ $X2=0 $Y2=0
cc_997 N_A_761_113#_c_1293_n N_A_352_409#_c_2089_n 0.0292866f $X=4.98 $Y=1.72
+ $X2=0 $Y2=0
cc_998 N_A_761_113#_c_1294_n N_A_352_409#_c_2089_n 0.00327845f $X=4.98 $Y=1.72
+ $X2=0 $Y2=0
cc_999 N_A_761_113#_c_1307_n N_A_352_409#_c_2095_n 0.0146392f $X=4.825 $Y=2.045
+ $X2=0 $Y2=0
cc_1000 N_A_761_113#_c_1276_n N_VGND_c_2337_n 9.43806e-19 $X=4.955 $Y=1.06 $X2=0
+ $Y2=0
cc_1001 N_A_761_113#_c_1284_n N_VGND_c_2338_n 0.0210961f $X=10.71 $Y=0.18 $X2=0
+ $Y2=0
cc_1002 N_A_761_113#_c_1284_n N_VGND_c_2339_n 0.0261591f $X=10.71 $Y=0.18 $X2=0
+ $Y2=0
cc_1003 N_A_761_113#_c_1276_n N_VGND_c_2347_n 0.00409299f $X=4.955 $Y=1.06 $X2=0
+ $Y2=0
cc_1004 N_A_761_113#_c_1285_n N_VGND_c_2347_n 0.0346424f $X=6.395 $Y=0.18 $X2=0
+ $Y2=0
cc_1005 N_A_761_113#_c_1284_n N_VGND_c_2348_n 0.0354719f $X=10.71 $Y=0.18 $X2=0
+ $Y2=0
cc_1006 N_A_761_113#_c_1284_n N_VGND_c_2349_n 0.0483643f $X=10.71 $Y=0.18 $X2=0
+ $Y2=0
cc_1007 N_A_761_113#_c_1276_n N_VGND_c_2353_n 0.00437698f $X=4.955 $Y=1.06 $X2=0
+ $Y2=0
cc_1008 N_A_761_113#_c_1284_n N_VGND_c_2353_n 0.144365f $X=10.71 $Y=0.18 $X2=0
+ $Y2=0
cc_1009 N_A_761_113#_c_1285_n N_VGND_c_2353_n 0.0106778f $X=6.395 $Y=0.18 $X2=0
+ $Y2=0
cc_1010 N_A_2220_40#_c_1491_n N_A_2019_419#_M1013_g 0.0226906f $X=12.33 $Y=0.495
+ $X2=0 $Y2=0
cc_1011 N_A_2220_40#_c_1492_n N_A_2019_419#_c_1575_n 0.0148533f $X=12.725
+ $Y=1.285 $X2=0 $Y2=0
cc_1012 N_A_2220_40#_c_1497_n N_A_2019_419#_c_1575_n 5.4511e-19 $X=12.93
+ $Y=2.185 $X2=0 $Y2=0
cc_1013 N_A_2220_40#_c_1493_n N_A_2019_419#_c_1575_n 0.00153997f $X=12.827
+ $Y=2.02 $X2=0 $Y2=0
cc_1014 N_A_2220_40#_c_1491_n N_A_2019_419#_c_1576_n 0.00125587f $X=12.33
+ $Y=0.495 $X2=0 $Y2=0
cc_1015 N_A_2220_40#_c_1492_n N_A_2019_419#_c_1576_n 0.0112235f $X=12.725
+ $Y=1.285 $X2=0 $Y2=0
cc_1016 N_A_2220_40#_c_1491_n N_A_2019_419#_M1014_g 0.00347898f $X=12.33
+ $Y=0.495 $X2=0 $Y2=0
cc_1017 N_A_2220_40#_c_1493_n N_A_2019_419#_M1012_g 0.00342875f $X=12.827
+ $Y=2.02 $X2=0 $Y2=0
cc_1018 N_A_2220_40#_c_1497_n N_A_2019_419#_c_1590_n 0.00785035f $X=12.93
+ $Y=2.185 $X2=0 $Y2=0
cc_1019 N_A_2220_40#_M1029_g N_A_2019_419#_c_1592_n 0.00140589f $X=11.175
+ $Y=0.54 $X2=0 $Y2=0
cc_1020 N_A_2220_40#_M1029_g N_A_2019_419#_c_1593_n 0.0148867f $X=11.175 $Y=0.54
+ $X2=0 $Y2=0
cc_1021 N_A_2220_40#_M1029_g N_A_2019_419#_c_1595_n 0.0034779f $X=11.175 $Y=0.54
+ $X2=0 $Y2=0
cc_1022 N_A_2220_40#_c_1488_n N_A_2019_419#_c_1595_n 0.0259362f $X=11.41
+ $Y=1.885 $X2=0 $Y2=0
cc_1023 N_A_2220_40#_M1021_g N_A_2019_419#_c_1595_n 0.00683409f $X=11.41
+ $Y=2.595 $X2=0 $Y2=0
cc_1024 N_A_2220_40#_c_1496_n N_A_2019_419#_c_1595_n 0.0336422f $X=11.61 $Y=1.38
+ $X2=0 $Y2=0
cc_1025 N_A_2220_40#_c_1490_n N_A_2019_419#_c_1595_n 0.0124915f $X=11.775
+ $Y=1.285 $X2=0 $Y2=0
cc_1026 N_A_2220_40#_c_1488_n N_A_2019_419#_c_1633_n 0.00141747f $X=11.41
+ $Y=1.885 $X2=0 $Y2=0
cc_1027 N_A_2220_40#_M1021_g N_A_2019_419#_c_1633_n 0.0182238f $X=11.41 $Y=2.595
+ $X2=0 $Y2=0
cc_1028 N_A_2220_40#_c_1496_n N_A_2019_419#_c_1633_n 0.0135177f $X=11.61 $Y=1.38
+ $X2=0 $Y2=0
cc_1029 N_A_2220_40#_c_1497_n N_A_2019_419#_c_1603_n 0.0173771f $X=12.93
+ $Y=2.185 $X2=0 $Y2=0
cc_1030 N_A_2220_40#_M1021_g N_A_2019_419#_c_1641_n 6.66307e-19 $X=11.41
+ $Y=2.595 $X2=0 $Y2=0
cc_1031 N_A_2220_40#_c_1497_n N_A_2019_419#_c_1641_n 0.0333503f $X=12.93
+ $Y=2.185 $X2=0 $Y2=0
cc_1032 N_A_2220_40#_M1012_s N_A_2019_419#_c_1604_n 0.00300374f $X=12.79 $Y=2
+ $X2=0 $Y2=0
cc_1033 N_A_2220_40#_c_1497_n N_A_2019_419#_c_1604_n 0.0274783f $X=12.93
+ $Y=2.185 $X2=0 $Y2=0
cc_1034 N_A_2220_40#_c_1491_n N_A_2019_419#_c_1596_n 9.51712e-19 $X=12.33
+ $Y=0.495 $X2=0 $Y2=0
cc_1035 N_A_2220_40#_c_1492_n N_A_2019_419#_c_1596_n 0.0131113f $X=12.725
+ $Y=1.285 $X2=0 $Y2=0
cc_1036 N_A_2220_40#_c_1493_n N_A_2019_419#_c_1596_n 0.0336164f $X=12.827
+ $Y=2.02 $X2=0 $Y2=0
cc_1037 N_A_2220_40#_c_1492_n N_A_2019_419#_c_1597_n 8.08074e-19 $X=12.725
+ $Y=1.285 $X2=0 $Y2=0
cc_1038 N_A_2220_40#_c_1493_n N_A_2019_419#_c_1597_n 0.00657618f $X=12.827
+ $Y=2.02 $X2=0 $Y2=0
cc_1039 N_A_2220_40#_c_1493_n N_A_2019_419#_c_1605_n 0.00693763f $X=12.827
+ $Y=2.02 $X2=0 $Y2=0
cc_1040 N_A_2220_40#_M1021_g N_A_2019_419#_c_1685_n 0.00523371f $X=11.41
+ $Y=2.595 $X2=0 $Y2=0
cc_1041 N_A_2220_40#_c_1497_n N_A_2019_419#_c_1607_n 0.00188032f $X=12.93
+ $Y=2.185 $X2=0 $Y2=0
cc_1042 N_A_2220_40#_M1021_g N_VPWR_c_1860_n 0.0187395f $X=11.41 $Y=2.595 $X2=0
+ $Y2=0
cc_1043 N_A_2220_40#_M1021_g N_VPWR_c_1867_n 0.008763f $X=11.41 $Y=2.595 $X2=0
+ $Y2=0
cc_1044 N_A_2220_40#_M1021_g N_VPWR_c_1853_n 0.0146671f $X=11.41 $Y=2.595 $X2=0
+ $Y2=0
cc_1045 N_A_2220_40#_M1029_g N_VGND_c_2340_n 0.00300553f $X=11.175 $Y=0.54 $X2=0
+ $Y2=0
cc_1046 N_A_2220_40#_c_1489_n N_VGND_c_2340_n 0.00633469f $X=12.165 $Y=1.285
+ $X2=0 $Y2=0
cc_1047 N_A_2220_40#_c_1490_n N_VGND_c_2340_n 0.00888302f $X=11.775 $Y=1.285
+ $X2=0 $Y2=0
cc_1048 N_A_2220_40#_c_1491_n N_VGND_c_2340_n 0.0325934f $X=12.33 $Y=0.495 $X2=0
+ $Y2=0
cc_1049 N_A_2220_40#_c_1491_n N_VGND_c_2341_n 0.0153904f $X=12.33 $Y=0.495 $X2=0
+ $Y2=0
cc_1050 N_A_2220_40#_M1029_g N_VGND_c_2349_n 0.00495161f $X=11.175 $Y=0.54 $X2=0
+ $Y2=0
cc_1051 N_A_2220_40#_c_1491_n N_VGND_c_2350_n 0.0220321f $X=12.33 $Y=0.495 $X2=0
+ $Y2=0
cc_1052 N_A_2220_40#_M1029_g N_VGND_c_2353_n 0.00974028f $X=11.175 $Y=0.54 $X2=0
+ $Y2=0
cc_1053 N_A_2220_40#_c_1491_n N_VGND_c_2353_n 0.0125808f $X=12.33 $Y=0.495 $X2=0
+ $Y2=0
cc_1054 N_A_2019_419#_c_1588_n N_A_2865_74#_M1003_g 0.00970668f $X=15.04
+ $Y=0.865 $X2=0 $Y2=0
cc_1055 N_A_2019_419#_M1009_g N_A_2865_74#_c_1786_n 0.0163172f $X=14.985 $Y=2.37
+ $X2=0 $Y2=0
cc_1056 N_A_2019_419#_M1009_g N_A_2865_74#_c_1787_n 0.0306346f $X=14.985 $Y=2.37
+ $X2=0 $Y2=0
cc_1057 N_A_2019_419#_c_1591_n N_A_2865_74#_c_1787_n 0.00970668f $X=15.04
+ $Y=0.94 $X2=0 $Y2=0
cc_1058 N_A_2019_419#_c_1583_n N_A_2865_74#_c_1788_n 0.0101733f $X=13.895
+ $Y=1.32 $X2=0 $Y2=0
cc_1059 N_A_2019_419#_c_1585_n N_A_2865_74#_c_1788_n 0.0110965f $X=14.605
+ $Y=0.94 $X2=0 $Y2=0
cc_1060 N_A_2019_419#_c_1586_n N_A_2865_74#_c_1788_n 0.00177493f $X=14.68
+ $Y=0.865 $X2=0 $Y2=0
cc_1061 N_A_2019_419#_M1009_g N_A_2865_74#_c_1788_n 0.0161425f $X=14.985 $Y=2.37
+ $X2=0 $Y2=0
cc_1062 N_A_2019_419#_c_1591_n N_A_2865_74#_c_1788_n 0.00719114f $X=15.04
+ $Y=0.94 $X2=0 $Y2=0
cc_1063 N_A_2019_419#_M1017_g N_A_2865_74#_c_1796_n 0.00337976f $X=13.895 $Y=2.5
+ $X2=0 $Y2=0
cc_1064 N_A_2019_419#_M1009_g N_A_2865_74#_c_1796_n 0.0267026f $X=14.985 $Y=2.37
+ $X2=0 $Y2=0
cc_1065 N_A_2019_419#_M1009_g N_A_2865_74#_c_1789_n 0.0246017f $X=14.985 $Y=2.37
+ $X2=0 $Y2=0
cc_1066 N_A_2019_419#_M1009_g N_A_2865_74#_c_1790_n 0.00311526f $X=14.985
+ $Y=2.37 $X2=0 $Y2=0
cc_1067 N_A_2019_419#_c_1582_n N_A_2865_74#_c_1792_n 0.00121425f $X=13.695
+ $Y=0.78 $X2=0 $Y2=0
cc_1068 N_A_2019_419#_c_1585_n N_A_2865_74#_c_1792_n 0.0069861f $X=14.605
+ $Y=0.94 $X2=0 $Y2=0
cc_1069 N_A_2019_419#_c_1586_n N_A_2865_74#_c_1792_n 0.00897908f $X=14.68
+ $Y=0.865 $X2=0 $Y2=0
cc_1070 N_A_2019_419#_c_1588_n N_A_2865_74#_c_1792_n 0.00152256f $X=15.04
+ $Y=0.865 $X2=0 $Y2=0
cc_1071 N_A_2019_419#_M1017_g N_A_2865_74#_c_1793_n 0.00269891f $X=13.895 $Y=2.5
+ $X2=0 $Y2=0
cc_1072 N_A_2019_419#_M1009_g N_A_2865_74#_c_1793_n 0.00531849f $X=14.985
+ $Y=2.37 $X2=0 $Y2=0
cc_1073 N_A_2019_419#_c_1591_n N_A_2865_74#_c_1793_n 0.00491571f $X=15.04
+ $Y=0.94 $X2=0 $Y2=0
cc_1074 N_A_2019_419#_c_1633_n N_VPWR_M1021_d 0.0111002f $X=12.21 $Y=2.2 $X2=0
+ $Y2=0
cc_1075 N_A_2019_419#_c_1633_n N_VPWR_c_1860_n 0.0209601f $X=12.21 $Y=2.2 $X2=0
+ $Y2=0
cc_1076 N_A_2019_419#_c_1641_n N_VPWR_c_1860_n 0.0179821f $X=12.335 $Y=2.895
+ $X2=0 $Y2=0
cc_1077 N_A_2019_419#_c_1642_n N_VPWR_c_1860_n 0.00767604f $X=12.46 $Y=2.98
+ $X2=0 $Y2=0
cc_1078 N_A_2019_419#_M1012_g N_VPWR_c_1861_n 0.00495448f $X=13.195 $Y=2.5 $X2=0
+ $Y2=0
cc_1079 N_A_2019_419#_c_1579_n N_VPWR_c_1861_n 9.33255e-19 $X=13.62 $Y=1.245
+ $X2=0 $Y2=0
cc_1080 N_A_2019_419#_M1017_g N_VPWR_c_1861_n 0.0245573f $X=13.895 $Y=2.5 $X2=0
+ $Y2=0
cc_1081 N_A_2019_419#_c_1604_n N_VPWR_c_1861_n 0.0092562f $X=13.195 $Y=2.98
+ $X2=0 $Y2=0
cc_1082 N_A_2019_419#_c_1605_n N_VPWR_c_1861_n 0.0344562f $X=13.28 $Y=2.895
+ $X2=0 $Y2=0
cc_1083 N_A_2019_419#_M1009_g N_VPWR_c_1862_n 0.0257488f $X=14.985 $Y=2.37 $X2=0
+ $Y2=0
cc_1084 N_A_2019_419#_c_1606_n N_VPWR_c_1867_n 0.0216692f $X=10.37 $Y=2.24 $X2=0
+ $Y2=0
cc_1085 N_A_2019_419#_M1012_g N_VPWR_c_1868_n 0.00502067f $X=13.195 $Y=2.5 $X2=0
+ $Y2=0
cc_1086 N_A_2019_419#_c_1604_n N_VPWR_c_1868_n 0.0550914f $X=13.195 $Y=2.98
+ $X2=0 $Y2=0
cc_1087 N_A_2019_419#_c_1642_n N_VPWR_c_1868_n 0.014577f $X=12.46 $Y=2.98 $X2=0
+ $Y2=0
cc_1088 N_A_2019_419#_M1017_g N_VPWR_c_1869_n 0.00711337f $X=13.895 $Y=2.5 $X2=0
+ $Y2=0
cc_1089 N_A_2019_419#_M1009_g N_VPWR_c_1869_n 0.00747382f $X=14.985 $Y=2.37
+ $X2=0 $Y2=0
cc_1090 N_A_2019_419#_M1000_d N_VPWR_c_1853_n 0.0152343f $X=10.095 $Y=2.095
+ $X2=0 $Y2=0
cc_1091 N_A_2019_419#_M1027_d N_VPWR_c_1853_n 0.00232188f $X=12.235 $Y=2.095
+ $X2=0 $Y2=0
cc_1092 N_A_2019_419#_M1012_g N_VPWR_c_1853_n 0.00731936f $X=13.195 $Y=2.5 $X2=0
+ $Y2=0
cc_1093 N_A_2019_419#_M1017_g N_VPWR_c_1853_n 0.0135914f $X=13.895 $Y=2.5 $X2=0
+ $Y2=0
cc_1094 N_A_2019_419#_M1009_g N_VPWR_c_1853_n 0.00779694f $X=14.985 $Y=2.37
+ $X2=0 $Y2=0
cc_1095 N_A_2019_419#_c_1604_n N_VPWR_c_1853_n 0.0328859f $X=13.195 $Y=2.98
+ $X2=0 $Y2=0
cc_1096 N_A_2019_419#_c_1642_n N_VPWR_c_1853_n 0.00948536f $X=12.46 $Y=2.98
+ $X2=0 $Y2=0
cc_1097 N_A_2019_419#_c_1606_n N_VPWR_c_1853_n 0.0126914f $X=10.37 $Y=2.24 $X2=0
+ $Y2=0
cc_1098 N_A_2019_419#_c_1609_n A_2193_419# 0.00719976f $X=11.16 $Y=2.2 $X2=-0.19
+ $Y2=-0.245
cc_1099 N_A_2019_419#_c_1595_n A_2193_419# 2.60378e-19 $X=11.245 $Y=2.115
+ $X2=-0.19 $Y2=-0.245
cc_1100 N_A_2019_419#_c_1685_n A_2193_419# 0.0030224f $X=11.245 $Y=2.2 $X2=-0.19
+ $Y2=-0.245
cc_1101 N_A_2019_419#_M1017_g N_Q_N_c_2268_n 0.0255508f $X=13.895 $Y=2.5 $X2=0
+ $Y2=0
cc_1102 N_A_2019_419#_c_1585_n N_Q_N_c_2268_n 0.00356886f $X=14.605 $Y=0.94
+ $X2=0 $Y2=0
cc_1103 N_A_2019_419#_M1009_g N_Q_N_c_2268_n 6.18397e-19 $X=14.985 $Y=2.37 $X2=0
+ $Y2=0
cc_1104 N_A_2019_419#_M1017_g N_Q_N_c_2273_n 0.0267255f $X=13.895 $Y=2.5 $X2=0
+ $Y2=0
cc_1105 N_A_2019_419#_M1009_g N_Q_N_c_2273_n 0.00432563f $X=14.985 $Y=2.37 $X2=0
+ $Y2=0
cc_1106 N_A_2019_419#_c_1590_n N_Q_N_c_2273_n 3.50661e-19 $X=13.075 $Y=1.84
+ $X2=0 $Y2=0
cc_1107 N_A_2019_419#_c_1607_n N_Q_N_c_2273_n 0.00552042f $X=13.177 $Y=1.84
+ $X2=0 $Y2=0
cc_1108 N_A_2019_419#_M1014_g Q_N 0.00559888f $X=12.905 $Y=0.495 $X2=0 $Y2=0
cc_1109 N_A_2019_419#_c_1579_n Q_N 0.00418706f $X=13.62 $Y=1.245 $X2=0 $Y2=0
cc_1110 N_A_2019_419#_c_1580_n Q_N 0.00492302f $X=13.62 $Y=0.855 $X2=0 $Y2=0
cc_1111 N_A_2019_419#_c_1582_n Q_N 0.00166615f $X=13.695 $Y=0.78 $X2=0 $Y2=0
cc_1112 N_A_2019_419#_c_1583_n Q_N 0.0229876f $X=13.895 $Y=1.32 $X2=0 $Y2=0
cc_1113 N_A_2019_419#_M1017_g Q_N 0.0104873f $X=13.895 $Y=2.5 $X2=0 $Y2=0
cc_1114 N_A_2019_419#_c_1596_n Q_N 0.0308571f $X=13.155 $Y=1.335 $X2=0 $Y2=0
cc_1115 N_A_2019_419#_c_1597_n Q_N 9.93497e-19 $X=13.155 $Y=1.335 $X2=0 $Y2=0
cc_1116 N_A_2019_419#_M1017_g N_Q_N_c_2270_n 0.00282089f $X=13.895 $Y=2.5 $X2=0
+ $Y2=0
cc_1117 N_A_2019_419#_c_1590_n N_Q_N_c_2270_n 7.02529e-19 $X=13.075 $Y=1.84
+ $X2=0 $Y2=0
cc_1118 N_A_2019_419#_c_1596_n N_Q_N_c_2270_n 0.0134146f $X=13.155 $Y=1.335
+ $X2=0 $Y2=0
cc_1119 N_A_2019_419#_c_1578_n N_Q_N_c_2271_n 0.00255628f $X=13.335 $Y=0.78
+ $X2=0 $Y2=0
cc_1120 N_A_2019_419#_c_1582_n N_Q_N_c_2271_n 0.0104082f $X=13.695 $Y=0.78 $X2=0
+ $Y2=0
cc_1121 N_A_2019_419#_c_1583_n N_Q_N_c_2271_n 0.010152f $X=13.895 $Y=1.32 $X2=0
+ $Y2=0
cc_1122 N_A_2019_419#_c_1586_n N_Q_N_c_2271_n 0.00307579f $X=14.68 $Y=0.865
+ $X2=0 $Y2=0
cc_1123 N_A_2019_419#_M1009_g N_Q_c_2314_n 2.74822e-19 $X=14.985 $Y=2.37 $X2=0
+ $Y2=0
cc_1124 N_A_2019_419#_M1013_g N_VGND_c_2340_n 0.00295332f $X=12.545 $Y=0.495
+ $X2=0 $Y2=0
cc_1125 N_A_2019_419#_M1013_g N_VGND_c_2341_n 0.002112f $X=12.545 $Y=0.495 $X2=0
+ $Y2=0
cc_1126 N_A_2019_419#_M1014_g N_VGND_c_2341_n 0.0134712f $X=12.905 $Y=0.495
+ $X2=0 $Y2=0
cc_1127 N_A_2019_419#_c_1578_n N_VGND_c_2341_n 0.0109841f $X=13.335 $Y=0.78
+ $X2=0 $Y2=0
cc_1128 N_A_2019_419#_c_1582_n N_VGND_c_2341_n 0.00130587f $X=13.695 $Y=0.78
+ $X2=0 $Y2=0
cc_1129 N_A_2019_419#_c_1589_n N_VGND_c_2341_n 0.00132199f $X=13.075 $Y=1.245
+ $X2=0 $Y2=0
cc_1130 N_A_2019_419#_c_1596_n N_VGND_c_2341_n 0.0125555f $X=13.155 $Y=1.335
+ $X2=0 $Y2=0
cc_1131 N_A_2019_419#_c_1586_n N_VGND_c_2342_n 0.00182089f $X=14.68 $Y=0.865
+ $X2=0 $Y2=0
cc_1132 N_A_2019_419#_c_1588_n N_VGND_c_2342_n 0.0130702f $X=15.04 $Y=0.865
+ $X2=0 $Y2=0
cc_1133 N_A_2019_419#_c_1592_n N_VGND_c_2349_n 0.0174108f $X=10.49 $Y=0.475
+ $X2=0 $Y2=0
cc_1134 N_A_2019_419#_M1013_g N_VGND_c_2350_n 0.00502664f $X=12.545 $Y=0.495
+ $X2=0 $Y2=0
cc_1135 N_A_2019_419#_M1014_g N_VGND_c_2350_n 0.00445056f $X=12.905 $Y=0.495
+ $X2=0 $Y2=0
cc_1136 N_A_2019_419#_c_1578_n N_VGND_c_2351_n 0.00445056f $X=13.335 $Y=0.78
+ $X2=0 $Y2=0
cc_1137 N_A_2019_419#_c_1580_n N_VGND_c_2351_n 4.57848e-19 $X=13.62 $Y=0.855
+ $X2=0 $Y2=0
cc_1138 N_A_2019_419#_c_1582_n N_VGND_c_2351_n 0.00327544f $X=13.695 $Y=0.78
+ $X2=0 $Y2=0
cc_1139 N_A_2019_419#_c_1586_n N_VGND_c_2351_n 0.00434272f $X=14.68 $Y=0.865
+ $X2=0 $Y2=0
cc_1140 N_A_2019_419#_c_1588_n N_VGND_c_2351_n 0.00383152f $X=15.04 $Y=0.865
+ $X2=0 $Y2=0
cc_1141 N_A_2019_419#_M1013_g N_VGND_c_2353_n 0.010303f $X=12.545 $Y=0.495 $X2=0
+ $Y2=0
cc_1142 N_A_2019_419#_M1014_g N_VGND_c_2353_n 0.00796275f $X=12.905 $Y=0.495
+ $X2=0 $Y2=0
cc_1143 N_A_2019_419#_c_1578_n N_VGND_c_2353_n 0.00796275f $X=13.335 $Y=0.78
+ $X2=0 $Y2=0
cc_1144 N_A_2019_419#_c_1580_n N_VGND_c_2353_n 6.33118e-19 $X=13.62 $Y=0.855
+ $X2=0 $Y2=0
cc_1145 N_A_2019_419#_c_1582_n N_VGND_c_2353_n 0.00563474f $X=13.695 $Y=0.78
+ $X2=0 $Y2=0
cc_1146 N_A_2019_419#_c_1585_n N_VGND_c_2353_n 0.00475329f $X=14.605 $Y=0.94
+ $X2=0 $Y2=0
cc_1147 N_A_2019_419#_c_1586_n N_VGND_c_2353_n 0.00825516f $X=14.68 $Y=0.865
+ $X2=0 $Y2=0
cc_1148 N_A_2019_419#_c_1588_n N_VGND_c_2353_n 0.00756787f $X=15.04 $Y=0.865
+ $X2=0 $Y2=0
cc_1149 N_A_2019_419#_c_1591_n N_VGND_c_2353_n 7.5656e-19 $X=15.04 $Y=0.94 $X2=0
+ $Y2=0
cc_1150 N_A_2019_419#_c_1592_n N_VGND_c_2353_n 0.0110845f $X=10.49 $Y=0.475
+ $X2=0 $Y2=0
cc_1151 N_A_2865_74#_c_1794_n N_VPWR_c_1862_n 0.0257237f $X=15.515 $Y=1.785
+ $X2=0 $Y2=0
cc_1152 N_A_2865_74#_c_1796_n N_VPWR_c_1862_n 0.0698785f $X=14.72 $Y=2.015 $X2=0
+ $Y2=0
cc_1153 N_A_2865_74#_c_1789_n N_VPWR_c_1862_n 0.025331f $X=15.395 $Y=1.575 $X2=0
+ $Y2=0
cc_1154 N_A_2865_74#_c_1796_n N_VPWR_c_1869_n 0.0137683f $X=14.72 $Y=2.015 $X2=0
+ $Y2=0
cc_1155 N_A_2865_74#_c_1794_n N_VPWR_c_1870_n 0.00747382f $X=15.515 $Y=1.785
+ $X2=0 $Y2=0
cc_1156 N_A_2865_74#_c_1794_n N_VPWR_c_1853_n 0.00779694f $X=15.515 $Y=1.785
+ $X2=0 $Y2=0
cc_1157 N_A_2865_74#_c_1796_n N_VPWR_c_1853_n 0.0147251f $X=14.72 $Y=2.015 $X2=0
+ $Y2=0
cc_1158 N_A_2865_74#_c_1796_n N_Q_N_c_2268_n 0.00912624f $X=14.72 $Y=2.015 $X2=0
+ $Y2=0
cc_1159 N_A_2865_74#_c_1793_n N_Q_N_c_2268_n 0.00396702f $X=14.672 $Y=1.575
+ $X2=0 $Y2=0
cc_1160 N_A_2865_74#_c_1796_n N_Q_N_c_2273_n 0.0769354f $X=14.72 $Y=2.015 $X2=0
+ $Y2=0
cc_1161 N_A_2865_74#_c_1788_n Q_N 0.0171935f $X=14.545 $Y=1.49 $X2=0 $Y2=0
cc_1162 N_A_2865_74#_c_1792_n Q_N 0.00322358f $X=14.465 $Y=0.58 $X2=0 $Y2=0
cc_1163 N_A_2865_74#_c_1793_n Q_N 0.00349829f $X=14.672 $Y=1.575 $X2=0 $Y2=0
cc_1164 N_A_2865_74#_c_1792_n N_Q_N_c_2271_n 0.0265419f $X=14.465 $Y=0.58 $X2=0
+ $Y2=0
cc_1165 N_A_2865_74#_M1003_g N_Q_c_2311_n 0.00125204f $X=15.47 $Y=0.58 $X2=0
+ $Y2=0
cc_1166 N_A_2865_74#_M1041_g N_Q_c_2311_n 0.0100639f $X=15.83 $Y=0.58 $X2=0
+ $Y2=0
cc_1167 N_A_2865_74#_c_1794_n Q 0.0134352f $X=15.515 $Y=1.785 $X2=0 $Y2=0
cc_1168 N_A_2865_74#_c_1794_n N_Q_c_2314_n 0.00589385f $X=15.515 $Y=1.785 $X2=0
+ $Y2=0
cc_1169 N_A_2865_74#_c_1786_n N_Q_c_2314_n 6.55907e-19 $X=15.56 $Y=1.495 $X2=0
+ $Y2=0
cc_1170 N_A_2865_74#_c_1789_n N_Q_c_2314_n 0.00881185f $X=15.395 $Y=1.575 $X2=0
+ $Y2=0
cc_1171 N_A_2865_74#_M1041_g N_Q_c_2312_n 0.00870018f $X=15.83 $Y=0.58 $X2=0
+ $Y2=0
cc_1172 N_A_2865_74#_c_1786_n N_Q_c_2312_n 0.00397155f $X=15.56 $Y=1.495 $X2=0
+ $Y2=0
cc_1173 N_A_2865_74#_c_1789_n N_Q_c_2312_n 0.00851731f $X=15.395 $Y=1.575 $X2=0
+ $Y2=0
cc_1174 N_A_2865_74#_c_1790_n N_Q_c_2312_n 0.0236709f $X=15.56 $Y=1.155 $X2=0
+ $Y2=0
cc_1175 N_A_2865_74#_c_1791_n N_Q_c_2312_n 0.00811515f $X=15.56 $Y=1.155 $X2=0
+ $Y2=0
cc_1176 N_A_2865_74#_M1003_g N_VGND_c_2342_n 0.012197f $X=15.47 $Y=0.58 $X2=0
+ $Y2=0
cc_1177 N_A_2865_74#_M1041_g N_VGND_c_2342_n 0.00182089f $X=15.83 $Y=0.58 $X2=0
+ $Y2=0
cc_1178 N_A_2865_74#_c_1790_n N_VGND_c_2342_n 0.00185662f $X=15.56 $Y=1.155
+ $X2=0 $Y2=0
cc_1179 N_A_2865_74#_c_1792_n N_VGND_c_2342_n 0.0153904f $X=14.465 $Y=0.58 $X2=0
+ $Y2=0
cc_1180 N_A_2865_74#_c_1792_n N_VGND_c_2351_n 0.014367f $X=14.465 $Y=0.58 $X2=0
+ $Y2=0
cc_1181 N_A_2865_74#_M1003_g N_VGND_c_2352_n 0.00383152f $X=15.47 $Y=0.58 $X2=0
+ $Y2=0
cc_1182 N_A_2865_74#_M1041_g N_VGND_c_2352_n 0.00434272f $X=15.83 $Y=0.58 $X2=0
+ $Y2=0
cc_1183 N_A_2865_74#_M1003_g N_VGND_c_2353_n 0.00756787f $X=15.47 $Y=0.58 $X2=0
+ $Y2=0
cc_1184 N_A_2865_74#_M1041_g N_VGND_c_2353_n 0.00824158f $X=15.83 $Y=0.58 $X2=0
+ $Y2=0
cc_1185 N_A_2865_74#_c_1792_n N_VGND_c_2353_n 0.0119227f $X=14.465 $Y=0.58 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1854_n N_A_245_409#_c_2022_n 0.0121616f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1863_n N_A_245_409#_c_2022_n 0.0221635f $X=2.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1853_n N_A_245_409#_c_2022_n 0.0126536f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1854_n N_A_245_409#_c_2023_n 0.0586203f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1855_n N_A_245_409#_c_2024_n 0.0129587f $X=2.92 $Y=2.865 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1863_n N_A_245_409#_c_2024_n 0.0626461f $X=2.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1853_n N_A_245_409#_c_2024_n 0.0367028f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1855_n N_A_245_409#_c_2029_n 0.0153156f $X=2.92 $Y=2.865 $X2=0
+ $Y2=0
cc_1194 N_VPWR_M1046_d N_A_245_409#_c_2030_n 0.00356107f $X=2.78 $Y=2.045 $X2=0
+ $Y2=0
cc_1195 N_VPWR_c_1855_n N_A_245_409#_c_2030_n 0.0159264f $X=2.92 $Y=2.865 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1853_n N_A_245_409#_c_2030_n 0.0115006f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1855_n N_A_245_409#_c_2025_n 0.0260268f $X=2.92 $Y=2.865 $X2=0
+ $Y2=0
cc_1198 N_VPWR_c_1865_n N_A_245_409#_c_2025_n 0.0220321f $X=4.38 $Y=3.33 $X2=0
+ $Y2=0
cc_1199 N_VPWR_c_1853_n N_A_245_409#_c_2025_n 0.0125808f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1200 N_VPWR_c_1853_n N_A_352_409#_M1008_s 0.00224633f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1201 N_VPWR_M1046_d N_A_352_409#_c_2090_n 0.00181172f $X=2.78 $Y=2.045 $X2=0
+ $Y2=0
cc_1202 N_VPWR_c_1853_n A_1373_419# 0.00225465f $X=16.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1203 N_VPWR_c_1853_n A_1921_419# 0.00282515f $X=16.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1204 N_VPWR_c_1853_n A_2193_419# 0.0137053f $X=16.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1205 N_VPWR_c_1861_n N_Q_N_c_2273_n 0.065672f $X=13.63 $Y=2.145 $X2=0 $Y2=0
cc_1206 N_VPWR_c_1869_n N_Q_N_c_2273_n 0.0130952f $X=15.085 $Y=3.33 $X2=0 $Y2=0
cc_1207 N_VPWR_c_1853_n N_Q_N_c_2273_n 0.00926016f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1208 N_VPWR_c_1861_n N_Q_N_c_2270_n 0.0188952f $X=13.63 $Y=2.145 $X2=0 $Y2=0
cc_1209 N_VPWR_c_1870_n Q 0.0193272f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1210 N_VPWR_c_1853_n Q 0.0206525f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1211 N_VPWR_c_1862_n N_Q_c_2314_n 0.0717213f $X=15.25 $Y=2.015 $X2=0 $Y2=0
cc_1212 N_A_245_409#_c_2024_n N_A_352_409#_M1045_d 0.00180746f $X=2.405 $Y=2.98
+ $X2=0 $Y2=0
cc_1213 N_A_245_409#_c_2023_n N_A_352_409#_c_2096_n 0.0378542f $X=1.37 $Y=2.19
+ $X2=0 $Y2=0
cc_1214 N_A_245_409#_c_2024_n N_A_352_409#_c_2096_n 0.015238f $X=2.405 $Y=2.98
+ $X2=0 $Y2=0
cc_1215 N_A_245_409#_c_2029_n N_A_352_409#_c_2096_n 0.00972699f $X=2.49 $Y=2.895
+ $X2=0 $Y2=0
cc_1216 N_A_245_409#_c_2031_n N_A_352_409#_c_2096_n 0.00823843f $X=2.575
+ $Y=2.405 $X2=0 $Y2=0
cc_1217 N_A_245_409#_c_2030_n N_A_352_409#_c_2090_n 0.0338482f $X=3.285 $Y=2.405
+ $X2=0 $Y2=0
cc_1218 N_A_245_409#_c_2031_n N_A_352_409#_c_2090_n 0.00857425f $X=2.575
+ $Y=2.405 $X2=0 $Y2=0
cc_1219 N_A_245_409#_c_2023_n N_A_352_409#_c_2091_n 0.00805415f $X=1.37 $Y=2.19
+ $X2=0 $Y2=0
cc_1220 N_A_245_409#_c_2024_n A_458_409# 0.00217487f $X=2.405 $Y=2.98 $X2=-0.19
+ $Y2=1.655
cc_1221 N_A_245_409#_c_2029_n A_458_409# 0.00445973f $X=2.49 $Y=2.895 $X2=-0.19
+ $Y2=1.655
cc_1222 N_A_245_409#_c_2031_n A_458_409# 0.00271405f $X=2.575 $Y=2.405 $X2=-0.19
+ $Y2=1.655
cc_1223 N_A_352_409#_c_2090_n A_458_409# 0.00295343f $X=3.015 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_1224 N_A_352_409#_c_2074_n N_VGND_c_2336_n 0.00130213f $X=3.015 $Y=0.845
+ $X2=0 $Y2=0
cc_1225 N_A_352_409#_c_2076_n N_VGND_c_2336_n 0.0104637f $X=3.505 $Y=0.845 $X2=0
+ $Y2=0
cc_1226 N_A_352_409#_c_2077_n N_VGND_c_2336_n 0.0110062f $X=3.59 $Y=0.76 $X2=0
+ $Y2=0
cc_1227 N_A_352_409#_c_2079_n N_VGND_c_2336_n 0.0144409f $X=3.675 $Y=0.35 $X2=0
+ $Y2=0
cc_1228 N_A_352_409#_c_2087_n N_VGND_c_2336_n 0.0129945f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_1229 N_A_352_409#_c_2139_n N_VGND_c_2336_n 0.0111573f $X=3.1 $Y=0.845 $X2=0
+ $Y2=0
cc_1230 N_A_352_409#_c_2078_n N_VGND_c_2337_n 0.0132716f $X=4.295 $Y=0.35 $X2=0
+ $Y2=0
cc_1231 N_A_352_409#_c_2080_n N_VGND_c_2337_n 0.0194919f $X=4.38 $Y=1.1 $X2=0
+ $Y2=0
cc_1232 N_A_352_409#_c_2081_n N_VGND_c_2337_n 0.013238f $X=5.015 $Y=1.185 $X2=0
+ $Y2=0
cc_1233 N_A_352_409#_c_2083_n N_VGND_c_2337_n 0.0194919f $X=5.1 $Y=1.1 $X2=0
+ $Y2=0
cc_1234 N_A_352_409#_c_2085_n N_VGND_c_2337_n 0.0132716f $X=5.185 $Y=0.35 $X2=0
+ $Y2=0
cc_1235 N_A_352_409#_c_2076_n N_VGND_c_2343_n 0.00254764f $X=3.505 $Y=0.845
+ $X2=0 $Y2=0
cc_1236 N_A_352_409#_c_2078_n N_VGND_c_2343_n 0.049001f $X=4.295 $Y=0.35 $X2=0
+ $Y2=0
cc_1237 N_A_352_409#_c_2079_n N_VGND_c_2343_n 0.0114429f $X=3.675 $Y=0.35 $X2=0
+ $Y2=0
cc_1238 N_A_352_409#_c_2074_n N_VGND_c_2346_n 0.00496182f $X=3.015 $Y=0.845
+ $X2=0 $Y2=0
cc_1239 N_A_352_409#_c_2087_n N_VGND_c_2346_n 0.0250411f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_1240 N_A_352_409#_c_2084_n N_VGND_c_2347_n 0.0671687f $X=6.02 $Y=0.35 $X2=0
+ $Y2=0
cc_1241 N_A_352_409#_c_2085_n N_VGND_c_2347_n 0.0114622f $X=5.185 $Y=0.35 $X2=0
+ $Y2=0
cc_1242 N_A_352_409#_M1016_d N_VGND_c_2353_n 0.0022543f $X=2.2 $Y=0.235 $X2=0
+ $Y2=0
cc_1243 N_A_352_409#_c_2074_n N_VGND_c_2353_n 0.0090016f $X=3.015 $Y=0.845 $X2=0
+ $Y2=0
cc_1244 N_A_352_409#_c_2076_n N_VGND_c_2353_n 0.00519846f $X=3.505 $Y=0.845
+ $X2=0 $Y2=0
cc_1245 N_A_352_409#_c_2078_n N_VGND_c_2353_n 0.0297409f $X=4.295 $Y=0.35 $X2=0
+ $Y2=0
cc_1246 N_A_352_409#_c_2079_n N_VGND_c_2353_n 0.00657383f $X=3.675 $Y=0.35 $X2=0
+ $Y2=0
cc_1247 N_A_352_409#_c_2084_n N_VGND_c_2353_n 0.0407196f $X=6.02 $Y=0.35 $X2=0
+ $Y2=0
cc_1248 N_A_352_409#_c_2085_n N_VGND_c_2353_n 0.00657784f $X=5.185 $Y=0.35 $X2=0
+ $Y2=0
cc_1249 N_A_352_409#_c_2087_n N_VGND_c_2353_n 0.016432f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_1250 N_A_352_409#_c_2139_n N_VGND_c_2353_n 6.51182e-19 $X=3.1 $Y=0.845 $X2=0
+ $Y2=0
cc_1251 N_Q_N_c_2271_n N_VGND_c_2341_n 0.0127769f $X=13.91 $Y=0.495 $X2=0 $Y2=0
cc_1252 N_Q_N_c_2271_n N_VGND_c_2351_n 0.033192f $X=13.91 $Y=0.495 $X2=0 $Y2=0
cc_1253 N_Q_N_c_2271_n N_VGND_c_2353_n 0.0188539f $X=13.91 $Y=0.495 $X2=0 $Y2=0
cc_1254 N_Q_c_2311_n N_VGND_c_2342_n 0.0153904f $X=16.045 $Y=0.58 $X2=0 $Y2=0
cc_1255 N_Q_c_2311_n N_VGND_c_2352_n 0.0143708f $X=16.045 $Y=0.58 $X2=0 $Y2=0
cc_1256 N_Q_c_2311_n N_VGND_c_2353_n 0.011923f $X=16.045 $Y=0.58 $X2=0 $Y2=0
cc_1257 A_138_47# N_VGND_c_2353_n 0.010279f $X=0.69 $Y=0.235 $X2=16.08 $Y2=0
cc_1258 N_VGND_c_2353_n A_362_47# 0.0034141f $X=16.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1259 N_VGND_c_2353_n A_526_47# 0.00323414f $X=16.08 $Y=0 $X2=-0.19 $Y2=-0.245
