* File: sky130_fd_sc_lp__o2111a_4.spice
* Created: Wed Sep  2 10:12:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111a_4.pex.spice"
.subckt sky130_fd_sc_lp__o2111a_4  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1018 N_A_32_65#_M1018_d N_D1_M1018_g N_A_32_367#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.231 AS=0.1176 PD=2.23 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1021 N_A_32_65#_M1021_d N_D1_M1021_g N_A_32_367#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1007 N_A_289_65#_M1007_d N_C1_M1007_g N_A_32_65#_M1021_d VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1005 N_A_389_65#_M1005_d N_B1_M1005_g N_A_289_65#_M1007_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_A_389_65#_M1005_d N_B1_M1015_g N_A_289_65#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1027 N_A_289_65#_M1015_s N_C1_M1027_g N_A_32_65#_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.3066 PD=1.12 PS=2.41 NRD=0 NRS=9.996 M=1 R=5.6
+ SA=75002.4 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1019 N_A_389_65#_M1019_d N_A2_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_389_65#_M1019_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1000_d N_A1_M1008_g N_A_389_65#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1023 N_A_389_65#_M1008_s N_A2_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75001.5
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1023_s N_A_32_367#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A_32_367#_M1010_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1010_d N_A_32_367#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1020 N_VGND_M1020_d N_A_32_367#_M1020_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_D1_M1013_g N_A_32_367#_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.6 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1013_d N_D1_M1026_g N_A_32_367#_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.2 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_C1_M1016_g N_A_32_367#_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1016_d N_B1_M1004_g N_A_32_367#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=7.0329 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_B1_M1017_g N_A_32_367#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75002.8
+ A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1017_d N_C1_M1022_g N_A_32_367#_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4725 PD=1.54 PS=2.01 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1006 N_A_741_367#_M1006_d N_A2_M1006_g N_A_32_367#_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4725 PD=1.54 PS=2.01 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1001 N_A_741_367#_M1006_d N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_A_741_367#_M1011_d N_A1_M1011_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1024 N_A_741_367#_M1011_d N_A2_M1024_g N_A_32_367#_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_32_367#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_32_367#_M1009_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1009_d N_A_32_367#_M1014_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_A_32_367#_M1025_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.0319 P=19.85
c_81 VNB 0 1.86413e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o2111a_4.pxi.spice"
*
.ends
*
*
