* File: sky130_fd_sc_lp__nor4_0.pxi.spice
* Created: Fri Aug 28 10:57:08 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4_0%A N_A_M1006_g N_A_c_65_n N_A_M1003_g N_A_c_62_n
+ N_A_c_68_n N_A_c_69_n A A N_A_c_64_n PM_SKY130_FD_SC_LP__NOR4_0%A
x_PM_SKY130_FD_SC_LP__NOR4_0%B N_B_M1007_g N_B_M1005_g N_B_c_101_n N_B_c_106_n B
+ B N_B_c_103_n PM_SKY130_FD_SC_LP__NOR4_0%B
x_PM_SKY130_FD_SC_LP__NOR4_0%C N_C_c_138_n N_C_M1000_g N_C_M1004_g N_C_c_144_n C
+ C N_C_c_141_n PM_SKY130_FD_SC_LP__NOR4_0%C
x_PM_SKY130_FD_SC_LP__NOR4_0%D N_D_M1002_g N_D_c_175_n N_D_M1001_g D D D D
+ N_D_c_176_n N_D_c_177_n N_D_c_178_n D PM_SKY130_FD_SC_LP__NOR4_0%D
x_PM_SKY130_FD_SC_LP__NOR4_0%VPWR N_VPWR_M1003_s N_VPWR_c_214_n VPWR
+ N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_213_n N_VPWR_c_218_n
+ PM_SKY130_FD_SC_LP__NOR4_0%VPWR
x_PM_SKY130_FD_SC_LP__NOR4_0%Y N_Y_M1006_d N_Y_M1004_d N_Y_M1002_d N_Y_c_235_n
+ N_Y_c_243_n N_Y_c_244_n N_Y_c_236_n N_Y_c_245_n N_Y_c_237_n N_Y_c_238_n Y Y Y
+ N_Y_c_240_n N_Y_c_241_n PM_SKY130_FD_SC_LP__NOR4_0%Y
x_PM_SKY130_FD_SC_LP__NOR4_0%VGND N_VGND_M1006_s N_VGND_M1007_d N_VGND_M1001_d
+ N_VGND_c_298_n N_VGND_c_299_n N_VGND_c_300_n N_VGND_c_301_n N_VGND_c_302_n
+ N_VGND_c_303_n VGND N_VGND_c_304_n N_VGND_c_305_n
+ PM_SKY130_FD_SC_LP__NOR4_0%VGND
cc_1 VNB N_A_M1006_g 0.0390532f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.56
cc_2 VNB N_A_c_62_n 0.0209276f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.695
cc_3 VNB A 0.00517371f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_c_64_n 0.0165043f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_5 VNB N_B_M1007_g 0.0370158f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.56
cc_6 VNB N_B_c_101_n 0.0192457f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_7 VNB B 0.00545467f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.695
cc_8 VNB N_B_c_103_n 0.0157577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_c_138_n 0.0207164f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.56
cc_10 VNB N_C_M1004_g 0.0361447f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.735
cc_11 VNB C 0.00153965f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.19
cc_12 VNB N_C_c_141_n 0.0181673f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.175
cc_13 VNB N_D_c_175_n 0.00602066f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.1
cc_14 VNB N_D_c_176_n 0.0977548f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_15 VNB N_D_c_177_n 0.0399158f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_16 VNB N_D_c_178_n 0.0219673f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.295
cc_17 VNB D 0.00199964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_213_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_235_n 0.0301657f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_20 VNB N_Y_c_236_n 0.00124925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_237_n 0.011329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_238_n 0.0269801f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_23 VNB Y 0.00295071f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_24 VNB N_Y_c_240_n 0.00798359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_241_n 0.00124584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_298_n 0.0144275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_299_n 0.0207953f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.19
cc_28 VNB N_VGND_c_300_n 0.0224213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_301_n 0.0115308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_302_n 0.0149083f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_31 VNB N_VGND_c_303_n 0.00600627f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB N_VGND_c_304_n 0.0317808f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_33 VNB N_VGND_c_305_n 0.180499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A_c_65_n 0.0151477f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.1
cc_35 VPB N_A_M1003_g 0.0254466f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.735
cc_36 VPB N_A_c_62_n 0.00272969f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.695
cc_37 VPB N_A_c_68_n 0.0165321f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.86
cc_38 VPB N_A_c_69_n 0.0217259f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.175
cc_39 VPB A 0.0032759f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_40 VPB N_B_M1005_g 0.0385196f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.25
cc_41 VPB N_B_c_101_n 0.00251031f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_42 VPB N_B_c_106_n 0.0155978f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.19
cc_43 VPB B 0.00322855f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.695
cc_44 VPB N_C_c_138_n 0.00207881f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.56
cc_45 VPB N_C_M1000_g 0.0384151f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.86
cc_46 VPB N_C_c_144_n 0.0182114f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_47 VPB C 0.00176287f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.19
cc_48 VPB N_D_M1002_g 0.0236552f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.56
cc_49 VPB N_D_c_175_n 0.0505403f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.1
cc_50 VPB D 0.0454572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB D 0.0180805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_214_n 0.0320463f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.1
cc_53 VPB N_VPWR_c_215_n 0.0153494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_216_n 0.0652498f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.175
cc_55 VPB N_VPWR_c_213_n 0.0983778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_218_n 0.00541171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_235_n 0.0194346f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_58 VPB N_Y_c_243_n 0.0600903f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.19
cc_59 VPB N_Y_c_244_n 0.0150699f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.695
cc_60 VPB N_Y_c_245_n 0.024005f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_61 N_A_M1006_g N_B_M1007_g 0.0252673f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_62 N_A_c_65_n N_B_M1005_g 0.00797626f $X=0.615 $Y=2.1 $X2=0 $Y2=0
cc_63 N_A_c_69_n N_B_M1005_g 0.0597303f $X=0.795 $Y=2.175 $X2=0 $Y2=0
cc_64 N_A_c_62_n N_B_c_101_n 0.0116022f $X=0.525 $Y=1.695 $X2=0 $Y2=0
cc_65 N_A_c_68_n N_B_c_106_n 0.0116022f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_66 A B 0.0541544f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_c_64_n B 5.69245e-19 $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_68 A N_B_c_103_n 0.00484707f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_64_n N_B_c_103_n 0.0116022f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_VPWR_c_214_n 0.0177941f $X=0.795 $Y=2.735 $X2=0 $Y2=0
cc_71 N_A_c_69_n N_VPWR_c_214_n 0.00479998f $X=0.795 $Y=2.175 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_VPWR_c_216_n 0.00452967f $X=0.795 $Y=2.735 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_VPWR_c_213_n 0.00809218f $X=0.795 $Y=2.735 $X2=0 $Y2=0
cc_74 N_A_M1006_g N_Y_c_235_n 0.00538517f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_75 N_A_c_65_n N_Y_c_235_n 0.00592428f $X=0.615 $Y=2.1 $X2=0 $Y2=0
cc_76 A N_Y_c_235_n 0.0512332f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_64_n N_Y_c_235_n 0.016285f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_78 N_A_c_65_n N_Y_c_243_n 0.00443615f $X=0.615 $Y=2.1 $X2=0 $Y2=0
cc_79 N_A_c_68_n N_Y_c_243_n 0.00357851f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_80 N_A_c_69_n N_Y_c_243_n 0.0175089f $X=0.795 $Y=2.175 $X2=0 $Y2=0
cc_81 A N_Y_c_243_n 0.0294637f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 A Y 0.013393f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_Y_c_240_n 0.0137646f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_84 A N_Y_c_240_n 0.020579f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_c_64_n N_Y_c_240_n 0.00369723f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_86 N_A_M1006_g N_Y_c_241_n 0.00174332f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_87 N_A_M1006_g N_VGND_c_299_n 0.00946566f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_88 N_A_M1006_g N_VGND_c_304_n 0.00450927f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_89 N_A_M1006_g N_VGND_c_305_n 0.00398153f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_90 N_B_c_101_n N_C_c_138_n 0.0279903f $X=1.095 $Y=1.695 $X2=0 $Y2=0
cc_91 N_B_M1005_g N_C_M1000_g 0.0279903f $X=1.185 $Y=2.735 $X2=0 $Y2=0
cc_92 N_B_M1007_g N_C_M1004_g 0.0103405f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_93 N_B_c_106_n N_C_c_144_n 0.0279903f $X=1.095 $Y=1.86 $X2=0 $Y2=0
cc_94 B C 0.0528286f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B_c_103_n C 6.57212e-19 $X=1.095 $Y=1.355 $X2=0 $Y2=0
cc_96 B N_C_c_141_n 0.00439319f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B_c_103_n N_C_c_141_n 0.0279903f $X=1.095 $Y=1.355 $X2=0 $Y2=0
cc_98 N_B_M1005_g N_VPWR_c_214_n 0.0041831f $X=1.185 $Y=2.735 $X2=0 $Y2=0
cc_99 N_B_M1005_g N_VPWR_c_216_n 0.00545548f $X=1.185 $Y=2.735 $X2=0 $Y2=0
cc_100 N_B_M1005_g N_VPWR_c_213_n 0.0104231f $X=1.185 $Y=2.735 $X2=0 $Y2=0
cc_101 N_B_M1005_g N_Y_c_243_n 0.0148742f $X=1.185 $Y=2.735 $X2=0 $Y2=0
cc_102 N_B_c_106_n N_Y_c_243_n 0.00394184f $X=1.095 $Y=1.86 $X2=0 $Y2=0
cc_103 B N_Y_c_243_n 0.0253015f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_Y_c_238_n 0.0158491f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_105 B N_Y_c_238_n 0.0285049f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B_c_103_n N_Y_c_238_n 0.00125743f $X=1.095 $Y=1.355 $X2=0 $Y2=0
cc_107 N_B_M1007_g N_Y_c_241_n 0.00173197f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_VGND_c_299_n 5.3482e-19 $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_109 N_B_M1007_g N_VGND_c_304_n 0.0135334f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_110 N_B_M1007_g N_VGND_c_305_n 0.00382481f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_111 N_C_c_138_n N_D_c_175_n 0.0321832f $X=1.675 $Y=1.685 $X2=0 $Y2=0
cc_112 N_C_M1000_g N_D_c_175_n 0.067245f $X=1.575 $Y=2.735 $X2=0 $Y2=0
cc_113 N_C_M1004_g N_D_c_176_n 0.0321832f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_114 C N_D_c_176_n 0.00275859f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_C_M1004_g N_D_c_177_n 0.00158289f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_116 C N_D_c_177_n 0.0219398f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_C_M1004_g N_D_c_178_n 0.0106599f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_118 N_C_M1000_g N_VPWR_c_216_n 0.00545548f $X=1.575 $Y=2.735 $X2=0 $Y2=0
cc_119 N_C_M1000_g N_VPWR_c_213_n 0.0104231f $X=1.575 $Y=2.735 $X2=0 $Y2=0
cc_120 N_C_M1000_g N_Y_c_243_n 0.0159278f $X=1.575 $Y=2.735 $X2=0 $Y2=0
cc_121 N_C_c_144_n N_Y_c_243_n 0.00205848f $X=1.675 $Y=1.86 $X2=0 $Y2=0
cc_122 C N_Y_c_243_n 0.0206412f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_123 N_C_M1004_g N_Y_c_236_n 0.00175182f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_124 N_C_M1000_g N_Y_c_245_n 0.00415793f $X=1.575 $Y=2.735 $X2=0 $Y2=0
cc_125 N_C_M1004_g N_Y_c_238_n 0.0135767f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_126 C N_Y_c_238_n 0.022998f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_C_c_141_n N_Y_c_238_n 0.00264837f $X=1.665 $Y=1.355 $X2=0 $Y2=0
cc_128 N_C_M1004_g N_VGND_c_300_n 5.47421e-19 $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_129 N_C_M1004_g N_VGND_c_302_n 0.00398346f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_130 N_C_M1004_g N_VGND_c_304_n 0.00939667f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_131 N_C_M1004_g N_VGND_c_305_n 0.00398153f $X=1.775 $Y=0.56 $X2=0 $Y2=0
cc_132 N_D_M1002_g N_VPWR_c_216_n 0.00511657f $X=1.965 $Y=2.735 $X2=0 $Y2=0
cc_133 D N_VPWR_c_216_n 0.00467679f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_134 N_D_M1002_g N_VPWR_c_213_n 0.0105917f $X=1.965 $Y=2.735 $X2=0 $Y2=0
cc_135 D N_VPWR_c_213_n 0.00786317f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_136 N_D_c_175_n N_Y_c_243_n 0.0272366f $X=2.152 $Y=2.1 $X2=0 $Y2=0
cc_137 D N_Y_c_243_n 0.0148625f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_138 N_D_c_176_n N_Y_c_243_n 0.00297382f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_139 D N_Y_c_243_n 0.00112929f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_140 N_D_c_178_n N_Y_c_236_n 0.00175182f $X=2.36 $Y=0.88 $X2=0 $Y2=0
cc_141 N_D_M1002_g N_Y_c_245_n 0.0180914f $X=1.965 $Y=2.735 $X2=0 $Y2=0
cc_142 N_D_c_175_n N_Y_c_245_n 0.00641191f $X=2.152 $Y=2.1 $X2=0 $Y2=0
cc_143 D N_Y_c_245_n 0.0308006f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_144 N_D_c_176_n N_Y_c_238_n 0.00585157f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_145 N_D_c_177_n N_Y_c_238_n 0.00854528f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_146 N_D_c_178_n N_Y_c_238_n 0.00127713f $X=2.36 $Y=0.88 $X2=0 $Y2=0
cc_147 N_D_c_176_n N_VGND_c_300_n 0.00196253f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_148 N_D_c_177_n N_VGND_c_300_n 0.0219111f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_149 N_D_c_178_n N_VGND_c_300_n 0.0107449f $X=2.36 $Y=0.88 $X2=0 $Y2=0
cc_150 N_D_c_178_n N_VGND_c_302_n 0.00396895f $X=2.36 $Y=0.88 $X2=0 $Y2=0
cc_151 N_D_c_178_n N_VGND_c_304_n 5.35708e-19 $X=2.36 $Y=0.88 $X2=0 $Y2=0
cc_152 N_D_c_176_n N_VGND_c_305_n 0.00113681f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_153 N_D_c_178_n N_VGND_c_305_n 0.00771726f $X=2.36 $Y=0.88 $X2=0 $Y2=0
cc_154 N_VPWR_c_214_n N_Y_c_243_n 0.0257154f $X=0.58 $Y=2.57 $X2=0 $Y2=0
cc_155 N_VPWR_c_216_n N_Y_c_245_n 0.0220321f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_156 N_VPWR_c_213_n N_Y_c_245_n 0.0125808f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_157 N_Y_c_237_n N_VGND_c_299_n 0.00579027f $X=0.26 $Y=0.93 $X2=0 $Y2=0
cc_158 N_Y_c_240_n N_VGND_c_299_n 0.0186359f $X=0.695 $Y=0.93 $X2=0 $Y2=0
cc_159 N_Y_c_236_n N_VGND_c_302_n 0.0064776f $X=1.99 $Y=0.56 $X2=0 $Y2=0
cc_160 N_Y_c_238_n N_VGND_c_304_n 0.0490802f $X=1.895 $Y=0.93 $X2=0 $Y2=0
cc_161 N_Y_c_241_n N_VGND_c_304_n 0.00637979f $X=0.79 $Y=0.56 $X2=0 $Y2=0
cc_162 N_Y_c_236_n N_VGND_c_305_n 0.00673089f $X=1.99 $Y=0.56 $X2=0 $Y2=0
cc_163 N_Y_c_237_n N_VGND_c_305_n 0.00460967f $X=0.26 $Y=0.93 $X2=0 $Y2=0
cc_164 N_Y_c_238_n N_VGND_c_305_n 0.0122233f $X=1.895 $Y=0.93 $X2=0 $Y2=0
cc_165 N_Y_c_240_n N_VGND_c_305_n 0.00585948f $X=0.695 $Y=0.93 $X2=0 $Y2=0
cc_166 N_Y_c_241_n N_VGND_c_305_n 0.00655188f $X=0.79 $Y=0.56 $X2=0 $Y2=0
