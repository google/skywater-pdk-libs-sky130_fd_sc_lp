* File: sky130_fd_sc_lp__and4bb_2.spice
* Created: Fri Aug 28 10:09:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4bb_2.pex.spice"
.subckt sky130_fd_sc_lp__and4bb_2  VNB VPB A_N C D B_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B_N	B_N
* D	D
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_27_133#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_185_23#_M1006_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_X_M1006_d N_A_185_23#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 A_516_125# N_A_27_133#_M1015_g N_A_185_23#_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1011 A_588_125# N_A_558_99#_M1011_g A_516_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 A_696_125# N_C_M1001_g A_588_125# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g A_696_125# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_558_99#_M1005_d N_B_N_M1005_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0819 PD=1.41 PS=0.81 NRD=0 NRS=31.428 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_N_M1009_g N_A_27_133#_M1009_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=80.3169 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_185_23#_M1003_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.285075 PD=1.54 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1012 N_X_M1003_d N_A_185_23#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.43785 PD=1.54 PS=3.18 NRD=0 NRS=29.6879 M=1 R=8.4 SA=75000.8
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_A_185_23#_M1008_d N_A_27_133#_M1008_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.14595 PD=0.7 PS=1.06 NRD=0 NRS=93.7917 M=1 R=2.8
+ SA=75001.9 SB=75002 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_558_99#_M1004_g N_A_185_23#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_185_23#_M1002_d N_C_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06615 AS=0.0672 PD=0.735 PS=0.74 NRD=0 NRS=18.7544 M=1 R=2.8 SA=75002.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_185_23#_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.05985 AS=0.06615 PD=0.705 PS=0.735 NRD=0 NRS=16.4101 M=1 R=2.8 SA=75003.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_558_99#_M1007_d N_B_N_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.05985 PD=1.37 PS=0.705 NRD=0 NRS=2.3443 M=1 R=2.8
+ SA=75003.7 SB=75000.2 A=0.063 P=1.14 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
c_53 VNB 0 4.80826e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__and4bb_2.pxi.spice"
*
.ends
*
*
