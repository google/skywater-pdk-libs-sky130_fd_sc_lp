# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfstp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.915000 2.340000 2.245000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.800000 0.255000 11.025000 1.075000 ;
        RECT 10.800000 1.075000 12.390000 1.245000 ;
        RECT 10.800000 1.765000 12.390000 1.935000 ;
        RECT 10.800000 1.935000 11.025000 3.075000 ;
        RECT 11.695000 0.255000 11.885000 1.075000 ;
        RECT 11.695000 1.935000 11.885000 3.075000 ;
        RECT 12.145000 1.245000 12.390000 1.765000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645000 0.780000 5.110000 1.765000 ;
        RECT 4.645000 1.765000 8.485000 1.835000 ;
        RECT 4.645000 1.835000 6.350000 1.935000 ;
        RECT 4.645000 1.935000 4.845000 2.155000 ;
        RECT 6.180000 1.325000 8.485000 1.765000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.380000 0.815000 2.130000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.480000 0.085000 ;
        RECT  0.985000  0.085000  1.205000 0.870000 ;
        RECT  1.985000  0.085000  2.225000 0.970000 ;
        RECT  3.575000  0.085000  3.905000 0.815000 ;
        RECT  4.905000  0.085000  5.750000 0.610000 ;
        RECT  5.420000  0.610000  5.750000 0.885000 ;
        RECT  7.475000  0.085000  8.145000 0.785000 ;
        RECT 10.370000  0.085000 10.630000 1.105000 ;
        RECT 11.195000  0.085000 11.525000 0.905000 ;
        RECT 12.055000  0.085000 12.385000 0.905000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.480000 3.415000 ;
        RECT  0.695000 2.640000  1.025000 3.245000 ;
        RECT  2.135000 2.415000  2.465000 3.245000 ;
        RECT  3.805000 2.360000  4.135000 3.245000 ;
        RECT  5.015000 2.105000  5.275000 3.245000 ;
        RECT  7.995000 2.355000  8.325000 3.245000 ;
        RECT  9.005000 1.720000  9.265000 3.245000 ;
        RECT 10.375000 1.795000 10.630000 3.245000 ;
        RECT 11.195000 2.105000 11.525000 3.245000 ;
        RECT 12.055000 2.105000 12.385000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.170000 0.540000  0.360000 2.300000 ;
      RECT 0.170000 2.300000  1.260000 2.470000 ;
      RECT 0.170000 2.470000  0.525000 2.975000 ;
      RECT 1.000000 1.495000  1.260000 2.300000 ;
      RECT 1.195000 2.640000  1.600000 2.970000 ;
      RECT 1.375000 0.540000  1.815000 0.935000 ;
      RECT 1.430000 0.935000  1.815000 1.485000 ;
      RECT 1.430000 1.485000  2.600000 1.745000 ;
      RECT 1.430000 1.745000  1.600000 2.640000 ;
      RECT 2.395000 0.640000  2.650000 1.085000 ;
      RECT 2.395000 1.085000  2.950000 1.255000 ;
      RECT 2.635000 1.915000  2.950000 2.085000 ;
      RECT 2.635000 2.085000  2.865000 2.690000 ;
      RECT 2.780000 1.255000  2.950000 1.915000 ;
      RECT 2.820000 0.585000  3.300000 0.915000 ;
      RECT 3.035000 2.295000  3.300000 2.690000 ;
      RECT 3.130000 0.915000  3.300000 1.555000 ;
      RECT 3.130000 1.555000  4.465000 1.725000 ;
      RECT 3.130000 1.725000  3.300000 2.295000 ;
      RECT 3.480000 0.985000  4.445000 1.155000 ;
      RECT 3.480000 1.155000  3.810000 1.385000 ;
      RECT 3.660000 1.895000  4.475000 2.155000 ;
      RECT 4.115000 0.285000  4.445000 0.985000 ;
      RECT 4.135000 1.325000  4.465000 1.555000 ;
      RECT 4.305000 2.155000  4.475000 2.325000 ;
      RECT 4.305000 2.325000  4.660000 2.690000 ;
      RECT 5.370000 1.150000  6.010000 1.595000 ;
      RECT 5.445000 2.105000  5.775000 2.865000 ;
      RECT 5.445000 2.865000  7.345000 3.065000 ;
      RECT 5.965000 2.105000  6.295000 2.525000 ;
      RECT 5.965000 2.525000  7.825000 2.695000 ;
      RECT 6.210000 0.255000  6.705000 0.955000 ;
      RECT 6.210000 0.955000  9.265000 1.125000 ;
      RECT 6.520000 2.015000  8.835000 2.185000 ;
      RECT 6.520000 2.185000  6.795000 2.355000 ;
      RECT 7.565000 2.355000  7.825000 2.525000 ;
      RECT 8.315000 0.265000  9.775000 0.435000 ;
      RECT 8.315000 0.435000  8.575000 0.785000 ;
      RECT 8.495000 2.185000  8.835000 2.660000 ;
      RECT 8.655000 1.125000  9.265000 1.205000 ;
      RECT 8.655000 1.205000  8.835000 2.015000 ;
      RECT 8.935000 0.605000  9.265000 0.955000 ;
      RECT 9.435000 0.435000  9.775000 3.075000 ;
      RECT 9.945000 0.255000 10.200000 1.425000 ;
      RECT 9.945000 1.425000 11.975000 1.595000 ;
      RECT 9.945000 1.595000 10.205000 3.075000 ;
    LAYER mcon ;
      RECT 1.595000 1.210000 1.765000 1.380000 ;
      RECT 5.435000 1.210000 5.605000 1.380000 ;
    LAYER met1 ;
      RECT 1.535000 1.180000 1.825000 1.225000 ;
      RECT 1.535000 1.225000 5.665000 1.365000 ;
      RECT 1.535000 1.365000 1.825000 1.410000 ;
      RECT 5.375000 1.180000 5.665000 1.225000 ;
      RECT 5.375000 1.365000 5.665000 1.410000 ;
  END
END sky130_fd_sc_lp__dfstp_4
