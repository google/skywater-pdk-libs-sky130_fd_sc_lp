* NGSPICE file created from sky130_fd_sc_lp__nand4_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand4_2 A B C D VGND VNB VPB VPWR Y
M1000 VPWR D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=2.5704e+12p pd=1.668e+07u as=1.4112e+12p ps=1.232e+07u
M1001 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_69_47# D VGND VNB nshort w=840000u l=150000u
+  ad=7.056e+11p pd=6.72e+06u as=2.352e+11p ps=2.24e+06u
M1005 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_523_67# A Y VNB nshort w=840000u l=150000u
+  ad=6.972e+11p pd=6.7e+06u as=2.352e+11p ps=2.24e+06u
M1007 a_523_67# B a_330_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1008 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_330_47# C a_69_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND D a_69_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A a_523_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_330_47# B a_523_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_69_47# C a_330_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

