* File: sky130_fd_sc_lp__a21boi_4.pex.spice
* Created: Wed Sep  2 09:19:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BOI_4%B1_N 3 5 7 8 10 21
c34 3 0 7.98929e-20 $X=0.505 $Y=2.465
r35 19 21 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.595 $Y=1.35
+ $X2=0.705 $Y2=1.35
r36 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.35 $X2=0.595 $Y2=1.35
r37 16 19 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.35
+ $X2=0.595 $Y2=1.35
r38 10 20 2.7687 $w=5.38e-07 $l=1.25e-07 $layer=LI1_cond $X=0.72 $Y=1.48
+ $X2=0.595 $Y2=1.48
r39 8 20 7.86311 $w=5.38e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.595 $Y2=1.48
r40 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.185
+ $X2=0.705 $Y2=1.35
r41 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.705 $Y=1.185
+ $X2=0.705 $Y2=0.655
r42 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.505 $Y2=1.35
r43 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.505 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%A_33_367# 1 2 9 13 17 21 25 29 33 37 39 41
+ 45 47 49 50 52 54 57 63 73
c129 73 0 6.85997e-20 $X=2.445 $Y=1.45
c130 63 0 7.98929e-20 $X=1.19 $Y=1.46
c131 37 0 1.75263e-19 $X=2.745 $Y=2.465
r132 72 73 19.6426 $w=3.19e-07 $l=1.3e-07 $layer=POLY_cond $X=2.315 $Y=1.45
+ $X2=2.445 $Y2=1.45
r133 69 70 19.6426 $w=3.19e-07 $l=1.3e-07 $layer=POLY_cond $X=1.885 $Y=1.45
+ $X2=2.015 $Y2=1.45
r134 68 69 45.3292 $w=3.19e-07 $l=3e-07 $layer=POLY_cond $X=1.585 $Y=1.45
+ $X2=1.885 $Y2=1.45
r135 67 68 19.6426 $w=3.19e-07 $l=1.3e-07 $layer=POLY_cond $X=1.455 $Y=1.45
+ $X2=1.585 $Y2=1.45
r136 64 67 40.0408 $w=3.19e-07 $l=2.65e-07 $layer=POLY_cond $X=1.19 $Y=1.45
+ $X2=1.455 $Y2=1.45
r137 64 65 5.2884 $w=3.19e-07 $l=3.5e-08 $layer=POLY_cond $X=1.19 $Y=1.45
+ $X2=1.155 $Y2=1.45
r138 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.19
+ $Y=1.46 $X2=1.19 $Y2=1.46
r139 58 72 15.8652 $w=3.19e-07 $l=1.05e-07 $layer=POLY_cond $X=2.21 $Y=1.45
+ $X2=2.315 $Y2=1.45
r140 58 70 29.4639 $w=3.19e-07 $l=1.95e-07 $layer=POLY_cond $X=2.21 $Y=1.45
+ $X2=2.015 $Y2=1.45
r141 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.21
+ $Y=1.46 $X2=2.21 $Y2=1.46
r142 55 63 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.195 $Y=1.46
+ $X2=1.085 $Y2=1.46
r143 55 57 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=1.195 $Y=1.46
+ $X2=2.21 $Y2=1.46
r144 53 63 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=1.545
+ $X2=1.085 $Y2=1.46
r145 53 54 19.6439 $w=2.18e-07 $l=3.75e-07 $layer=LI1_cond $X=1.085 $Y=1.545
+ $X2=1.085 $Y2=1.92
r146 52 63 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=1.06 $Y=1.375
+ $X2=1.085 $Y2=1.46
r147 51 52 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.06 $Y=1.04
+ $X2=1.06 $Y2=1.375
r148 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=0.955
+ $X2=1.06 $Y2=1.04
r149 49 50 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.975 $Y=0.955
+ $X2=0.605 $Y2=0.955
r150 48 61 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.385 $Y=2.005
+ $X2=0.255 $Y2=2.005
r151 47 54 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.975 $Y=2.005
+ $X2=1.085 $Y2=1.92
r152 47 48 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.975 $Y=2.005
+ $X2=0.385 $Y2=2.005
r153 43 50 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.465 $Y=0.87
+ $X2=0.605 $Y2=0.955
r154 43 45 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=0.465 $Y=0.87
+ $X2=0.465 $Y2=0.42
r155 39 61 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=2.09
+ $X2=0.255 $Y2=2.005
r156 39 41 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=0.255 $Y=2.09
+ $X2=0.255 $Y2=2.455
r157 35 73 45.3292 $w=3.19e-07 $l=3.77492e-07 $layer=POLY_cond $X=2.745 $Y=1.625
+ $X2=2.445 $Y2=1.45
r158 35 37 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.745 $Y=1.625
+ $X2=2.745 $Y2=2.465
r159 31 73 20.418 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.445 $Y=1.275
+ $X2=2.445 $Y2=1.45
r160 31 33 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.445 $Y=1.275
+ $X2=2.445 $Y2=0.655
r161 27 72 20.418 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.315 $Y=1.625
+ $X2=2.315 $Y2=1.45
r162 27 29 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.315 $Y=1.625
+ $X2=2.315 $Y2=2.465
r163 23 70 20.418 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.015 $Y=1.275
+ $X2=2.015 $Y2=1.45
r164 23 25 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.015 $Y=1.275
+ $X2=2.015 $Y2=0.655
r165 19 69 20.418 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.885 $Y=1.625
+ $X2=1.885 $Y2=1.45
r166 19 21 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.885 $Y=1.625
+ $X2=1.885 $Y2=2.465
r167 15 68 20.418 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.585 $Y=1.275
+ $X2=1.585 $Y2=1.45
r168 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.585 $Y=1.275
+ $X2=1.585 $Y2=0.655
r169 11 67 20.418 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.455 $Y=1.625
+ $X2=1.455 $Y2=1.45
r170 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.455 $Y=1.625
+ $X2=1.455 $Y2=2.465
r171 7 65 20.418 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.155 $Y=1.275
+ $X2=1.155 $Y2=1.45
r172 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.155 $Y=1.275
+ $X2=1.155 $Y2=0.655
r173 2 61 600 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.005
r174 2 41 300 $w=1.7e-07 $l=6.79632e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.455
r175 1 45 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.365
+ $Y=0.235 $X2=0.49 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%A2 3 7 8 10 13 15 17 20 22 24 27 31 35 37
+ 38 39 45 55 67
c112 37 0 8.76637e-20 $X=5.52 $Y=1.295
c113 35 0 1.85116e-19 $X=3.195 $Y=1.35
c114 31 0 1.64578e-19 $X=3.172 $Y=1.16
c115 13 0 1.20647e-19 $X=5.365 $Y=2.465
r116 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.28
+ $Y=1.35 $X2=6.28 $Y2=1.35
r117 53 55 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.225 $Y=1.35
+ $X2=6.28 $Y2=1.35
r118 52 53 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.795 $Y=1.35
+ $X2=6.225 $Y2=1.35
r119 50 52 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.6 $Y=1.35
+ $X2=5.795 $Y2=1.35
r120 47 50 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=5.365 $Y=1.35
+ $X2=5.6 $Y2=1.35
r121 39 56 7.557 $w=3.03e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.362 $X2=6.28
+ $Y2=1.362
r122 38 56 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=6 $Y=1.362 $X2=6.28
+ $Y2=1.362
r123 37 67 9.35915 $w=4.38e-07 $l=1.85e-07 $layer=LI1_cond $X=5.52 $Y=1.295
+ $X2=5.335 $Y2=1.295
r124 37 38 11.474 $w=4.73e-07 $l=3.95e-07 $layer=LI1_cond $X=5.605 $Y=1.362
+ $X2=6 $Y2=1.362
r125 37 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=1.35 $X2=5.6 $Y2=1.35
r126 35 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.35
+ $X2=3.195 $Y2=1.515
r127 35 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.35
+ $X2=3.195 $Y2=1.185
r128 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=1.35 $X2=3.195 $Y2=1.35
r129 31 34 7.68295 $w=2.83e-07 $l=1.9e-07 $layer=LI1_cond $X=3.172 $Y=1.16
+ $X2=3.172 $Y2=1.35
r130 30 31 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.315 $Y=1.16
+ $X2=3.172 $Y2=1.16
r131 30 67 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=3.315 $Y=1.16
+ $X2=5.335 $Y2=1.16
r132 25 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.515
+ $X2=6.225 $Y2=1.35
r133 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.225 $Y=1.515
+ $X2=6.225 $Y2=2.465
r134 22 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.185
+ $X2=6.225 $Y2=1.35
r135 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.225 $Y=1.185
+ $X2=6.225 $Y2=0.655
r136 18 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=1.515
+ $X2=5.795 $Y2=1.35
r137 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.795 $Y=1.515
+ $X2=5.795 $Y2=2.465
r138 15 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=1.185
+ $X2=5.795 $Y2=1.35
r139 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.795 $Y=1.185
+ $X2=5.795 $Y2=0.655
r140 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.365 $Y=1.515
+ $X2=5.365 $Y2=1.35
r141 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.365 $Y=1.515
+ $X2=5.365 $Y2=2.465
r142 8 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.365 $Y=1.185
+ $X2=5.365 $Y2=1.35
r143 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.365 $Y=1.185
+ $X2=5.365 $Y2=0.655
r144 7 45 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.215 $Y=0.655
+ $X2=3.215 $Y2=1.185
r145 3 46 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.205 $Y=2.465
+ $X2=3.205 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 53
c78 53 0 1.83642e-19 $X=4.935 $Y=1.51
r79 51 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.845 $Y=1.51
+ $X2=4.935 $Y2=1.51
r80 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.845
+ $Y=1.51 $X2=4.845 $Y2=1.51
r81 48 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.505 $Y=1.51
+ $X2=4.845 $Y2=1.51
r82 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.505
+ $Y=1.51 $X2=4.505 $Y2=1.51
r83 46 48 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.075 $Y=1.51
+ $X2=4.505 $Y2=1.51
r84 44 46 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.825 $Y=1.51
+ $X2=4.075 $Y2=1.51
r85 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.51 $X2=3.825 $Y2=1.51
r86 41 44 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.645 $Y=1.51
+ $X2=3.825 $Y2=1.51
r87 36 52 6.70825 $w=3.33e-07 $l=1.95e-07 $layer=LI1_cond $X=5.04 $Y=1.582
+ $X2=4.845 $Y2=1.582
r88 35 52 9.80437 $w=3.33e-07 $l=2.85e-07 $layer=LI1_cond $X=4.56 $Y=1.582
+ $X2=4.845 $Y2=1.582
r89 35 49 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=4.56 $Y=1.582
+ $X2=4.505 $Y2=1.582
r90 34 49 14.6205 $w=3.33e-07 $l=4.25e-07 $layer=LI1_cond $X=4.08 $Y=1.582
+ $X2=4.505 $Y2=1.582
r91 34 45 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=4.08 $Y=1.582
+ $X2=3.825 $Y2=1.582
r92 33 45 7.74029 $w=3.33e-07 $l=2.25e-07 $layer=LI1_cond $X=3.6 $Y=1.582
+ $X2=3.825 $Y2=1.582
r93 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.675
+ $X2=4.935 $Y2=1.51
r94 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.935 $Y=1.675
+ $X2=4.935 $Y2=2.465
r95 25 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.345
+ $X2=4.935 $Y2=1.51
r96 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.935 $Y=1.345
+ $X2=4.935 $Y2=0.655
r97 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.675
+ $X2=4.505 $Y2=1.51
r98 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.505 $Y=1.675
+ $X2=4.505 $Y2=2.465
r99 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.345
+ $X2=4.505 $Y2=1.51
r100 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.505 $Y=1.345
+ $X2=4.505 $Y2=0.655
r101 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.675
+ $X2=4.075 $Y2=1.51
r102 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.075 $Y=1.675
+ $X2=4.075 $Y2=2.465
r103 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.345
+ $X2=4.075 $Y2=1.51
r104 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.075 $Y=1.345
+ $X2=4.075 $Y2=0.655
r105 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.675
+ $X2=3.645 $Y2=1.51
r106 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.645 $Y=1.675
+ $X2=3.645 $Y2=2.465
r107 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.345
+ $X2=3.645 $Y2=1.51
r108 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.645 $Y=1.345
+ $X2=3.645 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%VPWR 1 2 3 4 5 18 20 21 24 28 32 39 40 41
+ 43 55 59 66 67 70 73 76
r104 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r105 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 67 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r108 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r109 64 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.01 $Y2=3.33
r110 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r112 63 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 60 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.15 $Y2=3.33
r115 60 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.52 $Y2=3.33
r116 59 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6.01 $Y2=3.33
r117 59 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.52 $Y2=3.33
r118 58 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=5.15 $Y2=3.33
r121 55 57 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r122 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r123 51 54 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r124 51 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 50 53 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 48 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 46 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 43 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 41 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 41 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r135 39 53 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.43 $Y2=3.33
r137 38 57 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.6 $Y2=3.33
r138 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.43 $Y2=3.33
r139 32 35 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.01 $Y=2.19
+ $X2=6.01 $Y2=2.95
r140 30 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r141 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.95
r142 26 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=3.33
r143 26 28 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=2.375
r144 22 37 4.12218 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=2.377
+ $X2=3.43 $Y2=2.377
r145 22 24 34.0829 $w=2.33e-07 $l=6.95e-07 $layer=LI1_cond $X=3.595 $Y=2.377
+ $X2=4.29 $Y2=2.377
r146 21 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r147 20 37 2.94799 $w=3.3e-07 $l=1.18e-07 $layer=LI1_cond $X=3.43 $Y=2.495
+ $X2=3.43 $Y2=2.377
r148 20 21 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.43 $Y=2.495
+ $X2=3.43 $Y2=3.245
r149 16 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r150 16 18 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.345
r151 5 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=1.835 $X2=6.01 $Y2=2.95
r152 5 32 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=1.835 $X2=6.01 $Y2=2.19
r153 4 28 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=5.01
+ $Y=1.835 $X2=5.15 $Y2=2.375
r154 3 24 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=4.15
+ $Y=1.835 $X2=4.29 $Y2=2.375
r155 2 37 300 $w=1.7e-07 $l=6.1041e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=1.835 $X2=3.43 $Y2=2.375
r156 1 18 300 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%A_223_367# 1 2 3 4 5 6 7 22 24 26 30 32 35
+ 37 38 39 40 45 46 50 52 56 63 67 70
c99 52 0 1.20647e-19 $X=6.345 $Y=1.805
c100 30 0 1.75263e-19 $X=2.1 $Y=2.29
r101 74 75 5.33268 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=2.005
+ $X2=5.5 $Y2=2.09
r102 73 74 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.5 $Y=1.98
+ $X2=5.5 $Y2=2.005
r103 70 73 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.5 $Y=1.805
+ $X2=5.5 $Y2=1.98
r104 56 58 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=6.475 $Y=1.98
+ $X2=6.475 $Y2=2.91
r105 54 56 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=6.475 $Y=1.925
+ $X2=6.475 $Y2=1.98
r106 53 70 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=1.805
+ $X2=5.5 $Y2=1.805
r107 52 54 6.83069 $w=2.4e-07 $l=1.80278e-07 $layer=LI1_cond $X=6.345 $Y=1.805
+ $X2=6.475 $Y2=1.925
r108 52 53 32.6526 $w=2.38e-07 $l=6.8e-07 $layer=LI1_cond $X=6.345 $Y=1.805
+ $X2=5.665 $Y2=1.805
r109 50 75 21.8737 $w=1.78e-07 $l=3.55e-07 $layer=LI1_cond $X=5.575 $Y=2.445
+ $X2=5.575 $Y2=2.09
r110 47 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.815 $Y=2.005
+ $X2=4.72 $Y2=2.005
r111 46 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.005
+ $X2=5.5 $Y2=2.005
r112 46 47 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.335 $Y=2.005
+ $X2=4.815 $Y2=2.005
r113 45 69 5.42706 $w=1.9e-07 $l=2e-07 $layer=LI1_cond $X=4.72 $Y=2.665 $X2=4.72
+ $Y2=2.865
r114 44 67 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.72 $Y=2.09
+ $X2=4.72 $Y2=2.005
r115 44 45 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=4.72 $Y=2.09
+ $X2=4.72 $Y2=2.665
r116 40 69 2.57785 $w=4e-07 $l=9.5e-08 $layer=LI1_cond $X=4.625 $Y=2.865
+ $X2=4.72 $Y2=2.865
r117 40 42 22.0405 $w=3.98e-07 $l=7.65e-07 $layer=LI1_cond $X=4.625 $Y=2.865
+ $X2=3.86 $Y2=2.865
r118 38 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.625 $Y=2.005
+ $X2=4.72 $Y2=2.005
r119 38 39 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=4.625 $Y=2.005
+ $X2=3.095 $Y2=2.005
r120 35 65 3.75819 $w=2e-07 $l=1.2e-07 $layer=LI1_cond $X=2.995 $Y=2.835
+ $X2=2.995 $Y2=2.955
r121 35 37 37.4318 $w=1.98e-07 $l=6.75e-07 $layer=LI1_cond $X=2.995 $Y=2.835
+ $X2=2.995 $Y2=2.16
r122 34 39 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.995 $Y=2.09
+ $X2=3.095 $Y2=2.005
r123 34 37 3.88182 $w=1.98e-07 $l=7e-08 $layer=LI1_cond $X=2.995 $Y=2.09
+ $X2=2.995 $Y2=2.16
r124 33 63 5.23199 $w=3.25e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.265 $Y=2.955
+ $X2=2.1 $Y2=2.87
r125 32 65 3.13183 $w=2.4e-07 $l=1e-07 $layer=LI1_cond $X=2.895 $Y=2.955
+ $X2=2.995 $Y2=2.955
r126 32 33 30.2516 $w=2.38e-07 $l=6.3e-07 $layer=LI1_cond $X=2.895 $Y=2.955
+ $X2=2.265 $Y2=2.955
r127 28 63 1.28764 $w=3.3e-07 $l=2.05e-07 $layer=LI1_cond $X=2.1 $Y=2.665
+ $X2=2.1 $Y2=2.87
r128 28 30 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.1 $Y=2.665
+ $X2=2.1 $Y2=2.29
r129 27 61 2.82139 $w=4.1e-07 $l=1.3e-07 $layer=LI1_cond $X=1.335 $Y=2.87
+ $X2=1.205 $Y2=2.87
r130 26 63 5.23199 $w=3.25e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=2.87
+ $X2=2.1 $Y2=2.87
r131 26 27 16.865 $w=4.08e-07 $l=6e-07 $layer=LI1_cond $X=1.935 $Y=2.87
+ $X2=1.335 $Y2=2.87
r132 22 61 4.44912 $w=2.6e-07 $l=2.05e-07 $layer=LI1_cond $X=1.205 $Y=2.665
+ $X2=1.205 $Y2=2.87
r133 22 24 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=1.205 $Y=2.665
+ $X2=1.205 $Y2=2.425
r134 7 58 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.835 $X2=6.44 $Y2=2.91
r135 7 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.835 $X2=6.44 $Y2=1.98
r136 6 73 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.44
+ $Y=1.835 $X2=5.58 $Y2=1.98
r137 6 50 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.835 $X2=5.58 $Y2=2.445
r138 5 69 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=4.58
+ $Y=1.835 $X2=4.72 $Y2=2.9
r139 5 67 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=4.58
+ $Y=1.835 $X2=4.72 $Y2=2.085
r140 4 42 600 $w=1.7e-07 $l=1.0627e-06 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.835 $X2=3.86 $Y2=2.83
r141 3 65 400 $w=1.7e-07 $l=1.15688e-06 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.835 $X2=2.99 $Y2=2.91
r142 3 37 400 $w=1.7e-07 $l=4.01092e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.835 $X2=2.99 $Y2=2.16
r143 2 63 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=2.97
r144 2 30 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=2.29
r145 1 61 600 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.835 $X2=1.24 $Y2=2.91
r146 1 24 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.835 $X2=1.24 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%Y 1 2 3 4 5 6 20 22 25 29 35 38 42 43 44 45
+ 59 67 72
c87 72 0 1.85116e-19 $X=2.86 $Y=0.95
r88 71 72 8.28855 $w=5.08e-07 $l=1.58e-07 $layer=LI1_cond $X=2.702 $Y=0.95
+ $X2=2.86 $Y2=0.95
r89 66 68 0.46905 $w=5.08e-07 $l=2e-08 $layer=LI1_cond $X=2.23 $Y=0.95 $X2=2.25
+ $Y2=0.95
r90 66 67 7.93717 $w=5.08e-07 $l=9.5e-08 $layer=LI1_cond $X=2.23 $Y=0.95
+ $X2=2.135 $Y2=0.95
r91 54 59 1.82927 $w=3.13e-07 $l=5e-08 $layer=LI1_cond $X=2.702 $Y=1.715
+ $X2=2.702 $Y2=1.665
r92 53 71 3.56815 $w=3.15e-07 $l=2.55e-07 $layer=LI1_cond $X=2.702 $Y=1.205
+ $X2=2.702 $Y2=0.95
r93 45 54 5.41218 $w=3.02e-07 $l=2.67e-07 $layer=LI1_cond $X=2.435 $Y=1.715
+ $X2=2.702 $Y2=1.715
r94 45 59 0.658539 $w=3.13e-07 $l=1.8e-08 $layer=LI1_cond $X=2.702 $Y=1.647
+ $X2=2.702 $Y2=1.665
r95 44 45 12.8781 $w=3.13e-07 $l=3.52e-07 $layer=LI1_cond $X=2.702 $Y=1.295
+ $X2=2.702 $Y2=1.647
r96 44 53 3.29269 $w=3.13e-07 $l=9e-08 $layer=LI1_cond $X=2.702 $Y=1.295
+ $X2=2.702 $Y2=1.205
r97 43 71 1.45406 $w=5.08e-07 $l=6.2e-08 $layer=LI1_cond $X=2.64 $Y=0.95
+ $X2=2.702 $Y2=0.95
r98 43 68 9.14648 $w=5.08e-07 $l=3.9e-07 $layer=LI1_cond $X=2.64 $Y=0.95
+ $X2=2.25 $Y2=0.95
r99 38 40 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=0.535
+ $X2=1.38 $Y2=0.7
r100 33 35 47.6909 $w=1.98e-07 $l=8.6e-07 $layer=LI1_cond $X=3.86 $Y=0.795
+ $X2=4.72 $Y2=0.795
r101 33 72 55.4545 $w=1.98e-07 $l=1e-06 $layer=LI1_cond $X=3.86 $Y=0.795
+ $X2=2.86 $Y2=0.795
r102 27 68 5.41923 $w=2.3e-07 $l=2.55e-07 $layer=LI1_cond $X=2.25 $Y=0.695
+ $X2=2.25 $Y2=0.95
r103 27 29 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.25 $Y=0.695
+ $X2=2.25 $Y2=0.42
r104 26 42 3.09839 $w=3.2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.765 $Y=1.875
+ $X2=1.635 $Y2=1.875
r105 25 45 1.14084 $w=3.2e-07 $l=1.6e-07 $layer=LI1_cond $X=2.435 $Y=1.875
+ $X2=2.435 $Y2=1.715
r106 25 26 24.1293 $w=3.18e-07 $l=6.7e-07 $layer=LI1_cond $X=2.435 $Y=1.875
+ $X2=1.765 $Y2=1.875
r107 22 67 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.485 $Y=1.12
+ $X2=2.135 $Y2=1.12
r108 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.4 $Y=1.035
+ $X2=1.485 $Y2=1.12
r109 20 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.4 $Y=1.035
+ $X2=1.4 $Y2=0.7
r110 6 45 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.39
+ $Y=1.835 $X2=2.53 $Y2=1.98
r111 5 42 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.835 $X2=1.67 $Y2=1.98
r112 4 35 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=4.58
+ $Y=0.235 $X2=4.72 $Y2=0.79
r113 3 33 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.235 $X2=3.86 $Y2=0.79
r114 2 66 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.23 $Y2=0.93
r115 2 29 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.23 $Y2=0.42
r116 1 38 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=1.23
+ $Y=0.235 $X2=1.37 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%VGND 1 2 3 4 5 18 20 24 28 30 32 34 35 36
+ 47 52 58 63 66 68 72
r94 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r95 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r96 65 66 8.84873 $w=6.08e-07 $l=9.5e-08 $layer=LI1_cond $X=3 $Y=0.22 $X2=3.095
+ $Y2=0.22
r97 61 65 7.05882 $w=6.08e-07 $l=3.6e-07 $layer=LI1_cond $X=2.64 $Y=0.22 $X2=3
+ $Y2=0.22
r98 61 63 9.0448 $w=6.08e-07 $l=1.05e-07 $layer=LI1_cond $X=2.64 $Y=0.22
+ $X2=2.535 $Y2=0.22
r99 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r100 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r101 56 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r102 56 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r103 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r104 53 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.6
+ $Y2=0
r105 53 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=6
+ $Y2=0
r106 52 71 4.45891 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.305 $Y=0
+ $X2=6.512 $Y2=0
r107 52 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6
+ $Y2=0
r108 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r109 50 66 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.12 $Y=0 $X2=3.095
+ $Y2=0
r110 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r111 47 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.6
+ $Y2=0
r112 47 50 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=5.485 $Y=0
+ $X2=3.12 $Y2=0
r113 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r114 46 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r115 45 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.16 $Y=0
+ $X2=2.535 $Y2=0
r116 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r117 43 58 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=1.81
+ $Y2=0
r118 43 45 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.965 $Y=0
+ $X2=2.16 $Y2=0
r119 40 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r120 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 36 69 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=5.52 $Y2=0
r122 36 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r123 34 39 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.72
+ $Y2=0
r124 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.94
+ $Y2=0
r125 30 71 3.05877 $w=3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.455 $Y=0.085
+ $X2=6.512 $Y2=0
r126 30 32 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=6.455 $Y=0.085
+ $X2=6.455 $Y2=0.38
r127 26 68 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=0.085
+ $X2=5.6 $Y2=0
r128 26 28 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.6 $Y=0.085
+ $X2=5.6 $Y2=0.4
r129 22 58 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0
r130 22 24 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.36
r131 21 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=0.94
+ $Y2=0
r132 20 58 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.81
+ $Y2=0
r133 20 21 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.655 $Y=0
+ $X2=1.105 $Y2=0
r134 16 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=0.085
+ $X2=0.94 $Y2=0
r135 16 18 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.94 $Y=0.085
+ $X2=0.94 $Y2=0.56
r136 5 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.235 $X2=6.44 $Y2=0.38
r137 4 28 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.44
+ $Y=0.235 $X2=5.58 $Y2=0.4
r138 3 65 91 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=0.235 $X2=3 $Y2=0.36
r139 2 24 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.66
+ $Y=0.235 $X2=1.8 $Y2=0.36
r140 1 18 182 $w=1.7e-07 $l=3.9702e-07 $layer=licon1_NDIFF $count=1 $X=0.78
+ $Y=0.235 $X2=0.94 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_4%A_658_47# 1 2 3 4 13 19 20 21 23 25
r38 23 32 3.15628 $w=2.5e-07 $l=1.52e-07 $layer=LI1_cond $X=6.01 $Y=0.735
+ $X2=6.01 $Y2=0.887
r39 23 25 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=6.01 $Y=0.735
+ $X2=6.01 $Y2=0.42
r40 22 30 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.315 $Y=0.82
+ $X2=5.185 $Y2=0.82
r41 21 32 3.98688 $w=1.7e-07 $l=1.54919e-07 $layer=LI1_cond $X=5.885 $Y=0.82
+ $X2=6.01 $Y2=0.887
r42 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.885 $Y=0.82
+ $X2=5.315 $Y2=0.82
r43 20 30 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.185 $Y=0.735
+ $X2=5.185 $Y2=0.82
r44 19 28 3.47416 $w=2.6e-07 $l=1.35e-07 $layer=LI1_cond $X=5.185 $Y=0.525
+ $X2=5.185 $Y2=0.39
r45 19 20 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=5.185 $Y=0.525
+ $X2=5.185 $Y2=0.735
r46 15 18 36.7074 $w=2.68e-07 $l=8.6e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=4.29 $Y2=0.39
r47 13 28 3.34549 $w=2.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.055 $Y=0.39
+ $X2=5.185 $Y2=0.39
r48 13 18 32.6526 $w=2.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.055 $Y=0.39
+ $X2=4.29 $Y2=0.39
r49 4 32 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=0.235 $X2=6.01 $Y2=0.875
r50 4 25 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=0.235 $X2=6.01 $Y2=0.42
r51 3 30 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.235 $X2=5.15 $Y2=0.74
r52 3 28 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.235 $X2=5.15 $Y2=0.4
r53 2 18 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.15
+ $Y=0.235 $X2=4.29 $Y2=0.42
r54 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.235 $X2=3.43 $Y2=0.42
.ends

