# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfstp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfstp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.110000 0.550000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.805000 1.850000 13.325000 2.890000 ;
        RECT 12.995000 0.350000 13.325000 0.810000 ;
        RECT 13.085000 0.810000 13.325000 1.850000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.335000 1.550000 6.625000 1.595000 ;
        RECT 6.335000 1.595000 9.985000 1.735000 ;
        RECT 6.335000 1.735000 6.625000 1.780000 ;
        RECT 9.695000 1.550000 9.985000 1.595000 ;
        RECT 9.695000 1.735000 9.985000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.510000 1.450000 1.840000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.095000  0.085000  0.425000 0.725000 ;
      RECT  0.120000  2.025000  0.450000 3.245000 ;
      RECT  0.650000  2.025000  0.980000 3.065000 ;
      RECT  0.810000  0.265000  2.100000 0.435000 ;
      RECT  0.810000  0.435000  1.215000 0.725000 ;
      RECT  0.810000  0.725000  0.980000 2.025000 ;
      RECT  1.160000  1.100000  1.740000 1.270000 ;
      RECT  1.160000  1.270000  1.330000 1.960000 ;
      RECT  1.160000  1.960000  2.190000 2.130000 ;
      RECT  1.160000  2.130000  1.640000 3.065000 ;
      RECT  1.410000  0.615000  1.740000 1.100000 ;
      RECT  1.840000  2.310000  2.170000 3.245000 ;
      RECT  1.930000  0.435000  2.100000 1.100000 ;
      RECT  1.930000  1.100000  2.800000 1.165000 ;
      RECT  1.930000  1.165000  2.970000 1.270000 ;
      RECT  2.020000  1.515000  2.475000 1.845000 ;
      RECT  2.020000  1.845000  2.190000 1.960000 ;
      RECT  2.100000  1.270000  2.970000 1.335000 ;
      RECT  2.280000  0.085000  2.450000 0.920000 ;
      RECT  2.370000  2.025000  2.620000 2.895000 ;
      RECT  2.370000  2.895000  4.760000 3.065000 ;
      RECT  2.630000  0.265000  3.840000 0.435000 ;
      RECT  2.630000  0.435000  2.800000 1.100000 ;
      RECT  2.800000  1.335000  2.970000 2.075000 ;
      RECT  2.800000  2.075000  3.320000 2.715000 ;
      RECT  2.990000  0.615000  3.320000 0.985000 ;
      RECT  3.150000  0.985000  3.320000 1.245000 ;
      RECT  3.150000  1.245000  4.505000 1.575000 ;
      RECT  3.150000  1.575000  3.670000 1.840000 ;
      RECT  3.500000  1.840000  3.670000 2.895000 ;
      RECT  3.510000  0.435000  3.840000 1.065000 ;
      RECT  3.850000  2.075000  4.855000 2.245000 ;
      RECT  3.850000  2.245000  4.180000 2.715000 ;
      RECT  4.085000  0.605000  4.335000 0.875000 ;
      RECT  4.085000  0.875000  5.515000 1.045000 ;
      RECT  4.085000  1.045000  4.855000 1.065000 ;
      RECT  4.590000  2.435000  5.620000 2.605000 ;
      RECT  4.590000  2.605000  4.760000 2.895000 ;
      RECT  4.685000  1.065000  4.855000 2.075000 ;
      RECT  4.915000  0.085000  5.165000 0.695000 ;
      RECT  4.940000  2.785000  5.270000 3.245000 ;
      RECT  5.035000  1.225000  5.865000 1.395000 ;
      RECT  5.035000  1.395000  5.365000 2.085000 ;
      RECT  5.035000  2.085000  6.155000 2.255000 ;
      RECT  5.345000  0.265000  6.505000 0.435000 ;
      RECT  5.345000  0.435000  5.515000 0.875000 ;
      RECT  5.450000  2.605000  5.620000 2.895000 ;
      RECT  5.450000  2.895000  6.505000 3.065000 ;
      RECT  5.575000  1.575000  6.215000 1.745000 ;
      RECT  5.575000  1.745000  5.905000 1.905000 ;
      RECT  5.695000  0.615000  6.155000 1.020000 ;
      RECT  5.695000  1.020000  5.865000 1.225000 ;
      RECT  5.825000  2.255000  6.155000 2.715000 ;
      RECT  6.045000  1.200000  7.240000 1.370000 ;
      RECT  6.045000  1.370000  6.215000 1.575000 ;
      RECT  6.335000  0.435000  6.505000 1.200000 ;
      RECT  6.335000  2.060000  7.780000 2.230000 ;
      RECT  6.335000  2.230000  6.505000 2.895000 ;
      RECT  6.395000  1.550000  6.700000 1.880000 ;
      RECT  6.685000  0.085000  7.015000 1.020000 ;
      RECT  6.685000  2.410000  7.015000 3.245000 ;
      RECT  6.910000  1.370000  7.240000 1.870000 ;
      RECT  7.450000  1.300000  7.780000 1.510000 ;
      RECT  7.450000  1.510000  8.655000 1.840000 ;
      RECT  7.450000  1.840000  7.780000 2.060000 ;
      RECT  7.960000  0.605000  8.290000 0.895000 ;
      RECT  7.960000  0.895000  9.005000 1.065000 ;
      RECT  8.045000  2.020000 10.255000 2.190000 ;
      RECT  8.045000  2.190000  8.375000 3.065000 ;
      RECT  8.835000  1.065000  9.005000 2.020000 ;
      RECT  9.145000  2.370000  9.475000 3.245000 ;
      RECT  9.185000  1.160000 10.655000 1.330000 ;
      RECT  9.185000  1.330000  9.490000 1.840000 ;
      RECT  9.435000  0.085000  9.765000 0.980000 ;
      RECT  9.700000  1.510000 10.030000 1.840000 ;
      RECT  9.925000  2.190000 10.255000 2.895000 ;
      RECT  9.925000  2.895000 11.085000 3.065000 ;
      RECT 10.065000  0.265000 10.395000 1.160000 ;
      RECT 10.485000  1.330000 10.655000 1.675000 ;
      RECT 10.485000  1.675000 10.735000 2.715000 ;
      RECT 10.835000  0.825000 11.165000 1.495000 ;
      RECT 10.855000  0.085000 11.185000 0.645000 ;
      RECT 10.915000  1.495000 11.085000 2.895000 ;
      RECT 11.265000  1.675000 11.515000 3.245000 ;
      RECT 11.415000  0.350000 11.865000 0.810000 ;
      RECT 11.695000  0.810000 11.865000 1.490000 ;
      RECT 11.695000  1.490000 12.840000 1.660000 ;
      RECT 11.695000  1.660000 12.075000 2.890000 ;
      RECT 12.205000  0.085000 12.535000 0.810000 ;
      RECT 12.275000  1.850000 12.605000 3.245000 ;
      RECT 12.510000  0.990000 12.840000 1.490000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.580000  6.565000 1.750000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.580000  9.925000 1.750000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
  END
END sky130_fd_sc_lp__dfstp_lp
END LIBRARY
