# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a21o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.265000 1.210000 4.645000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.700000 1.295000 4.085000 1.625000 ;
        RECT 3.915000 1.625000 4.085000 1.950000 ;
        RECT 3.915000 1.950000 5.125000 2.120000 ;
        RECT 4.955000 1.345000 5.430000 1.645000 ;
        RECT 4.955000 1.645000 5.125000 1.950000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.210000 2.935000 1.760000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.075000 2.035000 1.245000 ;
        RECT 0.155000 1.245000 0.805000 1.780000 ;
        RECT 0.155000 1.780000 1.915000 1.985000 ;
        RECT 0.865000 1.985000 1.055000 3.075000 ;
        RECT 0.985000 0.255000 1.175000 1.075000 ;
        RECT 1.725000 1.985000 1.915000 3.075000 ;
        RECT 1.845000 0.255000 2.035000 1.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.365000  2.155000 0.695000 3.245000 ;
      RECT 0.485000  0.085000 0.815000 0.905000 ;
      RECT 0.985000  1.415000 2.375000 1.610000 ;
      RECT 1.225000  2.155000 1.555000 3.245000 ;
      RECT 1.345000  0.085000 1.675000 0.905000 ;
      RECT 2.085000  1.815000 2.385000 3.245000 ;
      RECT 2.205000  0.870000 4.625000 1.030000 ;
      RECT 2.205000  1.030000 3.365000 1.040000 ;
      RECT 2.205000  1.040000 2.375000 1.415000 ;
      RECT 2.240000  0.085000 2.895000 0.700000 ;
      RECT 2.605000  1.930000 2.865000 2.905000 ;
      RECT 2.605000  2.905000 3.735000 3.075000 ;
      RECT 3.035000  1.910000 3.365000 2.735000 ;
      RECT 3.065000  0.255000 3.305000 0.860000 ;
      RECT 3.065000  0.860000 4.625000 0.870000 ;
      RECT 3.105000  1.040000 3.365000 1.910000 ;
      RECT 3.475000  0.085000 3.815000 0.690000 ;
      RECT 3.535000  1.815000 3.745000 2.300000 ;
      RECT 3.535000  2.300000 5.495000 2.470000 ;
      RECT 3.535000  2.470000 3.735000 2.905000 ;
      RECT 3.915000  2.640000 4.245000 3.245000 ;
      RECT 3.985000  0.255000 5.090000 0.435000 ;
      RECT 3.985000  0.435000 4.235000 0.690000 ;
      RECT 4.405000  0.605000 4.625000 0.860000 ;
      RECT 4.415000  2.470000 4.625000 3.075000 ;
      RECT 4.795000  0.435000 5.090000 1.105000 ;
      RECT 4.795000  2.640000 5.125000 3.245000 ;
      RECT 5.260000  0.085000 5.555000 1.105000 ;
      RECT 5.295000  1.815000 5.495000 2.300000 ;
      RECT 5.295000  2.470000 5.495000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__a21o_4
