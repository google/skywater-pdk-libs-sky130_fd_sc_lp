# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__srsdfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  20.64000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.840000 2.135000 2.170000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.590100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.995000 1.815000 20.535000 2.150000 ;
        RECT 19.995000 2.150000 20.325000 3.075000 ;
        RECT 20.205000 0.265000 20.535000 1.815000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.598000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.920000 1.550000 4.250000 1.880000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 1.550000 3.715000 1.880000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.500000 0.935000 2.170000 ;
    END
  END SCE
  PIN SLEEP_B
    ANTENNAGATEAREA  0.598000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.235000 1.120000 18.565000 1.450000 ;
    END
  END SLEEP_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 16.590000 1.460000 17.155000 1.790000 ;
    END
  END CLK
  PIN KAPWR
    ANTENNADIFFAREA  1.236750 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 20.570000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 20.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 20.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 20.640000 0.085000 ;
      RECT  0.000000  3.245000 20.640000 3.415000 ;
      RECT  0.105000  0.530000  0.355000 1.160000 ;
      RECT  0.105000  1.160000  1.660000 1.330000 ;
      RECT  0.105000  1.330000  0.435000 2.990000 ;
      RECT  0.535000  0.085000  0.865000 0.990000 ;
      RECT  0.620000  2.340000  0.950000 3.245000 ;
      RECT  1.070000  0.255000  3.405000 0.425000 ;
      RECT  1.070000  0.425000  1.320000 0.990000 ;
      RECT  1.225000  1.500000  2.080000 1.670000 ;
      RECT  1.225000  1.670000  1.395000 2.340000 ;
      RECT  1.225000  2.340000  2.635000 2.510000 ;
      RECT  1.490000  0.595000  2.475000 0.765000 ;
      RECT  1.490000  0.765000  1.660000 1.160000 ;
      RECT  1.830000  0.935000  2.080000 1.500000 ;
      RECT  2.305000  0.765000  2.475000 1.600000 ;
      RECT  2.305000  1.600000  2.880000 1.930000 ;
      RECT  2.305000  2.100000  4.755000 2.270000 ;
      RECT  2.305000  2.270000  2.635000 2.340000 ;
      RECT  2.305000  2.510000  2.635000 2.990000 ;
      RECT  2.645000  0.740000  2.975000 1.210000 ;
      RECT  2.645000  1.210000  4.375000 1.380000 ;
      RECT  3.155000  0.425000  3.405000 1.040000 ;
      RECT  3.245000  2.440000  3.575000 3.245000 ;
      RECT  3.615000  0.085000  3.865000 1.040000 ;
      RECT  4.045000  0.580000  4.375000 1.210000 ;
      RECT  4.425000  2.270000  4.755000 2.990000 ;
      RECT  4.545000  1.250000  5.205000 1.420000 ;
      RECT  4.545000  1.420000  4.715000 2.100000 ;
      RECT  4.615000  0.255000  6.590000 0.425000 ;
      RECT  4.615000  0.425000  4.865000 1.080000 ;
      RECT  4.885000  1.590000  5.215000 1.920000 ;
      RECT  4.925000  1.920000  5.095000 2.600000 ;
      RECT  4.925000  2.600000  5.950000 2.770000 ;
      RECT  5.035000  0.595000  6.055000 0.765000 ;
      RECT  5.035000  0.765000  5.205000 1.250000 ;
      RECT  5.265000  2.090000  7.110000 2.260000 ;
      RECT  5.265000  2.260000  5.555000 2.430000 ;
      RECT  5.375000  0.935000  5.555000 1.265000 ;
      RECT  5.385000  1.265000  5.555000 2.090000 ;
      RECT  5.725000  0.765000  6.055000 1.265000 ;
      RECT  5.780000  2.430000  8.725000 2.435000 ;
      RECT  5.780000  2.435000  7.680000 2.600000 ;
      RECT  5.960000  1.435000  6.610000 1.605000 ;
      RECT  5.960000  1.605000  6.290000 1.825000 ;
      RECT  6.120000  2.770000  6.450000 3.245000 ;
      RECT  6.260000  0.425000  6.590000 0.835000 ;
      RECT  6.280000  1.005000  9.530000 1.165000 ;
      RECT  6.280000  1.165000  8.135000 1.175000 ;
      RECT  6.280000  1.175000  6.610000 1.435000 ;
      RECT  6.780000  1.345000  7.795000 1.675000 ;
      RECT  6.780000  1.675000  7.110000 2.090000 ;
      RECT  7.050000  0.085000  7.380000 0.835000 ;
      RECT  7.340000  1.845000  8.135000 2.095000 ;
      RECT  7.510000  2.265000  8.725000 2.430000 ;
      RECT  7.590000  0.575000  7.840000 0.995000 ;
      RECT  7.590000  0.995000  9.530000 1.005000 ;
      RECT  7.850000  2.605000  8.180000 3.245000 ;
      RECT  7.965000  1.175000  8.135000 1.845000 ;
      RECT  8.020000  0.085000  8.350000 0.825000 ;
      RECT  8.395000  1.335000  8.990000 1.495000 ;
      RECT  8.395000  1.495000  9.540000 1.665000 ;
      RECT  8.395000  1.665000  8.725000 2.265000 ;
      RECT  8.395000  2.435000  8.725000 2.825000 ;
      RECT  8.555000  2.825000  8.725000 2.905000 ;
      RECT  8.555000  2.905000 13.455000 3.075000 ;
      RECT  9.200000  0.265000 10.930000 0.435000 ;
      RECT  9.200000  0.435000  9.530000 0.995000 ;
      RECT  9.200000  1.165000  9.530000 1.285000 ;
      RECT  9.210000  1.665000  9.540000 1.825000 ;
      RECT  9.890000  2.040000 10.500000 2.565000 ;
      RECT  9.890000  2.565000 12.540000 2.735000 ;
      RECT 10.190000  0.605000 10.500000 2.040000 ;
      RECT 10.680000  0.435000 10.930000 2.395000 ;
      RECT 11.100000  1.155000 12.235000 1.325000 ;
      RECT 11.100000  1.325000 11.430000 2.010000 ;
      RECT 11.100000  2.010000 14.955000 2.180000 ;
      RECT 11.365000  0.085000 11.695000 0.985000 ;
      RECT 11.640000  1.510000 11.970000 1.670000 ;
      RECT 11.640000  1.670000 14.525000 1.840000 ;
      RECT 11.905000  0.575000 12.235000 1.155000 ;
      RECT 12.210000  2.350000 19.325000 2.520000 ;
      RECT 12.210000  2.520000 12.540000 2.565000 ;
      RECT 12.695000  0.575000 12.945000 0.980000 ;
      RECT 12.695000  0.980000 13.845000 1.150000 ;
      RECT 12.930000  1.320000 14.185000 1.500000 ;
      RECT 13.125000  0.085000 13.455000 0.810000 ;
      RECT 13.125000  2.745000 13.455000 2.905000 ;
      RECT 13.625000  2.520000 13.955000 2.970000 ;
      RECT 13.675000  0.575000 13.845000 0.980000 ;
      RECT 14.015000  0.600000 15.315000 0.770000 ;
      RECT 14.015000  0.770000 14.185000 1.320000 ;
      RECT 14.355000  0.940000 16.435000 0.950000 ;
      RECT 14.355000  0.950000 16.760000 1.110000 ;
      RECT 14.355000  1.110000 14.525000 1.670000 ;
      RECT 14.525000  2.690000 14.975000 2.970000 ;
      RECT 14.695000  1.280000 14.955000 1.440000 ;
      RECT 14.695000  1.440000 15.815000 1.610000 ;
      RECT 14.695000  1.610000 14.955000 2.010000 ;
      RECT 14.985000  0.255000 17.100000 0.425000 ;
      RECT 14.985000  0.425000 15.315000 0.600000 ;
      RECT 15.645000  1.610000 15.815000 1.930000 ;
      RECT 15.645000  1.930000 16.080000 2.180000 ;
      RECT 15.985000  1.410000 16.420000 1.740000 ;
      RECT 16.105000  0.595000 16.435000 0.940000 ;
      RECT 16.105000  1.110000 16.760000 1.120000 ;
      RECT 16.250000  1.740000 16.420000 2.350000 ;
      RECT 16.280000  2.690000 16.675000 2.970000 ;
      RECT 16.590000  1.120000 17.495000 1.290000 ;
      RECT 16.855000  2.010000 17.495000 2.180000 ;
      RECT 16.925000  2.690000 17.730000 3.025000 ;
      RECT 16.930000  0.425000 17.100000 0.780000 ;
      RECT 16.930000  0.780000 18.345000 0.950000 ;
      RECT 17.325000  1.290000 17.495000 2.010000 ;
      RECT 17.475000  0.085000 17.805000 0.610000 ;
      RECT 17.895000  0.950000 18.065000 1.850000 ;
      RECT 17.895000  1.850000 18.490000 2.180000 ;
      RECT 18.015000  0.345000 18.345000 0.780000 ;
      RECT 18.735000  0.975000 19.685000 1.145000 ;
      RECT 18.735000  1.145000 18.905000 1.815000 ;
      RECT 18.735000  1.815000 18.985000 2.180000 ;
      RECT 18.805000  0.085000 19.055000 0.805000 ;
      RECT 19.075000  1.315000 19.345000 1.645000 ;
      RECT 19.155000  1.645000 19.325000 2.350000 ;
      RECT 19.235000  0.345000 19.685000 0.975000 ;
      RECT 19.495000  1.815000 19.825000 3.245000 ;
      RECT 19.515000  1.145000 19.685000 1.315000 ;
      RECT 19.515000  1.315000 20.020000 1.645000 ;
      RECT 19.855000  0.085000 20.025000 1.145000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  2.735000 14.725000 2.905000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  2.735000 16.645000 2.905000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  2.735000 17.125000 2.905000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.245000 18.565000 3.415000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.245000 19.045000 3.415000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.245000 19.525000 3.415000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.245000 20.005000 3.415000 ;
      RECT 20.315000 -0.085000 20.485000 0.085000 ;
      RECT 20.315000  3.245000 20.485000 3.415000 ;
  END
END sky130_fd_sc_lp__srsdfrtp_1
