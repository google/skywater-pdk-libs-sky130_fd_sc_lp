* File: sky130_fd_sc_lp__a21o_1.spice
* Created: Fri Aug 28 09:50:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21o_1.pex.spice"
.subckt sky130_fd_sc_lp__a21o_1  VNB VPB B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_80_237#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2688 AS=0.2226 PD=1.48 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1003 N_A_80_237#_M1003_d N_B1_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1659 AS=0.2688 PD=1.235 PS=1.48 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1002 A_378_47# N_A1_M1002_g N_A_80_237#_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.1659 PD=1.26 PS=1.235 NRD=22.14 NRS=6.42 M=1 R=5.6 SA=75001.5
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_378_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1764 PD=2.21 PS=1.26 NRD=0 NRS=22.14 M=1 R=5.6 SA=75002.1 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_80_237#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_A_300_367#_M1001_d N_B1_M1001_g N_A_80_237#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_300_367#_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2394 AS=0.1764 PD=1.64 PS=1.54 NRD=8.5892 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1004 N_A_300_367#_M1004_d N_A2_M1004_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2394 PD=3.05 PS=1.64 NRD=0 NRS=7.0329 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__a21o_1.pxi.spice"
*
.ends
*
*
