* NGSPICE file created from sky130_fd_sc_lp__clkinvlp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__clkinvlp_4 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.6e+11p pd=5.12e+06u as=8.1e+11p ps=7.62e+06u
M1001 a_268_67# A Y VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=1.54e+11p ps=1.66e+06u
M1002 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A a_110_67# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.52e+06u
M1004 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_110_67# A VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=2.915e+11p ps=3.26e+06u
M1007 VGND A a_268_67# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

