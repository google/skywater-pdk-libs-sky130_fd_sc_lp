* File: sky130_fd_sc_lp__fahcon_1.pex.spice
* Created: Fri Aug 28 10:35:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A 3 7 8 11 13
r40 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.51
+ $X2=0.55 $Y2=1.675
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.51
+ $X2=0.55 $Y2=1.345
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.55
+ $Y=1.51 $X2=0.55 $Y2=1.51
r43 8 12 4.5038 $w=4.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=1.562 $X2=0.55
+ $Y2=1.562
r44 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.54 $Y=0.815
+ $X2=0.54 $Y2=1.345
r45 3 14 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.525 $Y=2.465
+ $X2=0.525 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_33_367# 1 2 3 4 15 17 19 22 28 30 33 36
+ 37 41 42 44 45 47 49 51 53 59
c116 53 0 5.11154e-20 $X=2.585 $Y=1.93
r117 58 59 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.16 $Y=1.51
+ $X2=1.33 $Y2=1.51
r118 53 54 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=1.93
+ $X2=2.585 $Y2=1.765
r119 48 58 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.09 $Y=1.51 $X2=1.16
+ $Y2=1.51
r120 47 49 9.2829 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.087 $Y=1.51
+ $X2=1.087 $Y2=1.345
r121 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.51 $X2=1.09 $Y2=1.51
r122 44 45 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.282 $Y=2.125
+ $X2=0.282 $Y2=1.96
r123 41 54 45.4063 $w=2.48e-07 $l=9.85e-07 $layer=LI1_cond $X=2.58 $Y=0.78
+ $X2=2.58 $Y2=1.765
r124 38 41 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.58 $Y=0.435
+ $X2=2.58 $Y2=0.78
r125 36 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.455 $Y=0.35
+ $X2=2.58 $Y2=0.435
r126 36 37 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=2.455 $Y=0.35
+ $X2=1.19 $Y2=0.35
r127 34 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=1.165
+ $X2=1.105 $Y2=1.08
r128 34 49 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.105 $Y=1.165
+ $X2=1.105 $Y2=1.345
r129 33 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=0.995
+ $X2=1.105 $Y2=1.08
r130 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=0.435
+ $X2=1.19 $Y2=0.35
r131 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.105 $Y=0.435
+ $X2=1.105 $Y2=0.995
r132 31 42 3.25423 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.49 $Y=1.08 $X2=0.29
+ $Y2=1.08
r133 30 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.02 $Y=1.08
+ $X2=1.105 $Y2=1.08
r134 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.02 $Y=1.08
+ $X2=0.49 $Y2=1.08
r135 26 44 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=0.282 $Y=2.152
+ $X2=0.282 $Y2=2.125
r136 26 28 22.3903 $w=3.83e-07 $l=7.48e-07 $layer=LI1_cond $X=0.282 $Y=2.152
+ $X2=0.282 $Y2=2.9
r137 24 42 3.29812 $w=2.85e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.175 $Y=1.165
+ $X2=0.29 $Y2=1.08
r138 24 45 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.175 $Y=1.165
+ $X2=0.175 $Y2=1.96
r139 20 42 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=0.995
+ $X2=0.29 $Y2=1.08
r140 20 22 13.109 $w=3.98e-07 $l=4.55e-07 $layer=LI1_cond $X=0.29 $Y=0.995
+ $X2=0.29 $Y2=0.54
r141 17 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.345
+ $X2=1.33 $Y2=1.51
r142 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.33 $Y=1.345
+ $X2=1.33 $Y2=0.915
r143 13 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.675
+ $X2=1.16 $Y2=1.51
r144 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.16 $Y=1.675
+ $X2=1.16 $Y2=2.335
r145 4 53 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.795 $X2=2.585 $Y2=1.93
r146 3 44 400 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.31 $Y2=2.125
r147 3 28 400 $w=1.7e-07 $l=1.13519e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.31 $Y2=2.9
r148 2 41 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=2.38
+ $Y=0.635 $X2=2.54 $Y2=0.78
r149 1 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.18
+ $Y=0.395 $X2=0.325 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_329_269# 1 2 9 14 16 20 23 26 28 29 33 35
+ 41 43 44 45 51
c111 44 0 1.06147e-19 $X=4.22 $Y=1.775
c112 43 0 1.23395e-19 $X=3.215 $Y=0.395
c113 33 0 1.89636e-19 $X=4.22 $Y=1.94
c114 9 0 5.11154e-20 $X=1.72 $Y=2.255
r115 50 51 33.6995 $w=4.1e-07 $l=7.5e-08 $layer=POLY_cond $X=2.76 $Y=0.32
+ $X2=2.685 $Y2=0.32
r116 48 49 18.4595 $w=5.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.38 $Y=0.43
+ $X2=4.38 $Y2=1
r117 45 48 1.67871 $w=5.68e-07 $l=8e-08 $layer=LI1_cond $X=4.38 $Y=0.35 $X2=4.38
+ $Y2=0.43
r118 44 49 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=4.18 $Y=1.775
+ $X2=4.18 $Y2=1
r119 41 50 39.3377 $w=4.1e-07 $l=2.9e-07 $layer=POLY_cond $X=3.05 $Y=0.32
+ $X2=2.76 $Y2=0.32
r120 40 43 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0.395
+ $X2=3.215 $Y2=0.395
r121 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.05
+ $Y=0.36 $X2=3.05 $Y2=0.36
r122 33 44 7.56219 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.22 $Y=1.94
+ $X2=4.22 $Y2=1.775
r123 33 35 33.5256 $w=3.28e-07 $l=9.6e-07 $layer=LI1_cond $X=4.22 $Y=1.94
+ $X2=4.22 $Y2=2.9
r124 29 45 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=4.095 $Y=0.35
+ $X2=4.38 $Y2=0.35
r125 29 43 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=4.095 $Y=0.35
+ $X2=3.215 $Y2=0.35
r126 27 28 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=2.78 $Y=1.385
+ $X2=2.78 $Y2=1.535
r127 25 26 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.74 $Y=1.345
+ $X2=1.74 $Y2=1.495
r128 23 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.8 $Y=2.215
+ $X2=2.8 $Y2=1.535
r129 20 27 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.76 $Y=0.955
+ $X2=2.76 $Y2=1.385
r130 17 50 26.4667 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.76 $Y=0.525
+ $X2=2.76 $Y2=0.32
r131 17 20 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.76 $Y=0.525
+ $X2=2.76 $Y2=0.955
r132 16 51 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.835 $Y=0.19
+ $X2=2.685 $Y2=0.19
r133 14 25 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.76 $Y=0.915
+ $X2=1.76 $Y2=1.345
r134 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.76 $Y=0.265
+ $X2=1.835 $Y2=0.19
r135 11 14 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.76 $Y=0.265
+ $X2=1.76 $Y2=0.915
r136 9 26 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.72 $Y=2.255
+ $X2=1.72 $Y2=1.495
r137 2 35 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=4.08
+ $Y=1.795 $X2=4.22 $Y2=2.9
r138 2 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.08
+ $Y=1.795 $X2=4.22 $Y2=1.94
r139 1 48 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.25 $X2=4.5 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%B 3 8 9 10 14 17 19 22 23 24 27 29 31 33 36
+ 38 39 42 45 48 50 51 52 57
c144 42 0 2.38886e-20 $X=5.745 $Y=0.57
c145 38 0 1.23209e-19 $X=5.67 $Y=1.095
c146 27 0 2.02469e-20 $X=4.435 $Y=2.425
c147 23 0 1.89636e-19 $X=4.36 $Y=1.455
c148 17 0 2.29542e-19 $X=3.53 $Y=0.955
c149 3 0 1.47047e-19 $X=2.305 $Y=0.955
r150 56 58 32.3387 $w=3.13e-07 $l=2.1e-07 $layer=POLY_cond $X=4.885 $Y=1.275
+ $X2=5.095 $Y2=1.275
r151 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.365 $X2=4.885 $Y2=1.365
r152 52 57 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=4.56 $Y=1.355
+ $X2=4.885 $Y2=1.355
r153 46 48 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=3.425 $Y=1.61
+ $X2=3.53 $Y2=1.61
r154 44 45 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=2.337 $Y=1.535
+ $X2=2.337 $Y2=1.685
r155 40 42 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.745 $Y=1.02
+ $X2=5.745 $Y2=0.57
r156 39 58 57.0126 $w=3.13e-07 $l=3.6404e-07 $layer=POLY_cond $X=5.38 $Y=1.095
+ $X2=5.095 $Y2=1.275
r157 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.67 $Y=1.095
+ $X2=5.745 $Y2=1.02
r158 38 39 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.67 $Y=1.095
+ $X2=5.38 $Y2=1.095
r159 34 58 19.9686 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.095 $Y=1.53
+ $X2=5.095 $Y2=1.275
r160 34 36 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.095 $Y=1.53
+ $X2=5.095 $Y2=2.4
r161 31 56 13.8594 $w=3.13e-07 $l=9e-08 $layer=POLY_cond $X=4.795 $Y=1.275
+ $X2=4.885 $Y2=1.275
r162 31 33 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.795 $Y=1.2
+ $X2=4.795 $Y2=0.67
r163 30 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.51 $Y=1.455
+ $X2=4.435 $Y2=1.455
r164 29 31 24.674 $w=3.13e-07 $l=2.14243e-07 $layer=POLY_cond $X=4.72 $Y=1.455
+ $X2=4.795 $Y2=1.275
r165 29 30 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.72 $Y=1.455
+ $X2=4.51 $Y2=1.455
r166 25 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.435 $Y=1.53
+ $X2=4.435 $Y2=1.455
r167 25 27 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.435 $Y=1.53
+ $X2=4.435 $Y2=2.425
r168 23 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.36 $Y=1.455
+ $X2=4.435 $Y2=1.455
r169 23 24 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=4.36 $Y=1.455
+ $X2=4.005 $Y2=1.455
r170 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.93 $Y=1.53
+ $X2=4.005 $Y2=1.455
r171 21 22 756.33 $w=1.5e-07 $l=1.475e-06 $layer=POLY_cond $X=3.93 $Y=1.53
+ $X2=3.93 $Y2=3.005
r172 20 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.5 $Y=3.08
+ $X2=3.425 $Y2=3.08
r173 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.855 $Y=3.08
+ $X2=3.93 $Y2=3.005
r174 19 20 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=3.855 $Y=3.08
+ $X2=3.5 $Y2=3.08
r175 15 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.53 $Y=1.535
+ $X2=3.53 $Y2=1.61
r176 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.53 $Y=1.535
+ $X2=3.53 $Y2=0.955
r177 12 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.425 $Y=3.005
+ $X2=3.425 $Y2=3.08
r178 12 14 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.425 $Y=3.005
+ $X2=3.425 $Y2=2.215
r179 11 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.425 $Y=1.685
+ $X2=3.425 $Y2=1.61
r180 11 14 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.425 $Y=1.685
+ $X2=3.425 $Y2=2.215
r181 9 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.35 $Y=3.08
+ $X2=3.425 $Y2=3.08
r182 9 10 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=3.35 $Y=3.08
+ $X2=2.445 $Y2=3.08
r183 8 45 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.37 $Y=2.215
+ $X2=2.37 $Y2=1.685
r184 6 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.37 $Y=3.005
+ $X2=2.445 $Y2=3.08
r185 6 8 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.37 $Y=3.005
+ $X2=2.37 $Y2=2.215
r186 3 44 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.305 $Y=0.955
+ $X2=2.305 $Y2=1.535
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_367_119# 1 2 9 13 16 19 22 23 25 27 28 30
+ 34 35 39 40 44 45 46 47 48 49 50 57 60 62 70 72 75 87
c248 87 0 1.7833e-19 $X=9.585 $Y=0.925
c249 72 0 6.03739e-20 $X=6.82 $Y=1
c250 70 0 1.0543e-19 $X=6.82 $Y=1.165
c251 60 0 1.24317e-19 $X=6.96 $Y=0.925
c252 47 0 1.33605e-19 $X=6.815 $Y=0.925
c253 40 0 1.37952e-19 $X=9.585 $Y=1.35
c254 39 0 8.37252e-20 $X=9.585 $Y=1.35
r255 70 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.82 $Y=1.165
+ $X2=6.82 $Y2=1
r256 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.82
+ $Y=1.165 $X2=6.82 $Y2=1.165
r257 63 87 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=9.36 $Y=0.925
+ $X2=9.585 $Y2=0.925
r258 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0.925
+ $X2=9.36 $Y2=0.925
r259 60 71 7.09196 $w=3.88e-07 $l=2.4e-07 $layer=LI1_cond $X=6.85 $Y=0.925
+ $X2=6.85 $Y2=1.165
r260 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0.925
+ $X2=6.96 $Y2=0.925
r261 57 81 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6 $Y=0.925
+ $X2=5.755 $Y2=0.925
r262 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0.925 $X2=6
+ $Y2=0.925
r263 52 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.925
r264 50 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=0.925
+ $X2=6.96 $Y2=0.925
r265 49 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=9.36 $Y2=0.925
r266 49 50 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=7.105 $Y2=0.925
r267 48 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=0.925
+ $X2=6 $Y2=0.925
r268 47 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=0.925
+ $X2=6.96 $Y2=0.925
r269 47 48 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=6.815 $Y=0.925
+ $X2=6.145 $Y2=0.925
r270 46 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=0.925
+ $X2=2.16 $Y2=0.925
r271 45 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=6 $Y2=0.925
r272 45 46 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=2.305 $Y2=0.925
r273 43 75 19.0078 $w=3.83e-07 $l=6.35e-07 $layer=LI1_cond $X=2.082 $Y=1.415
+ $X2=2.082 $Y2=0.78
r274 43 44 8.7386 $w=3.83e-07 $l=1.7e-07 $layer=LI1_cond $X=1.997 $Y=1.415
+ $X2=1.997 $Y2=1.585
r275 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.585
+ $Y=1.35 $X2=9.585 $Y2=1.35
r276 37 87 2.17527 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=9.585 $Y=1.04
+ $X2=9.585 $Y2=0.925
r277 37 39 19.101 $w=1.78e-07 $l=3.1e-07 $layer=LI1_cond $X=9.585 $Y=1.04
+ $X2=9.585 $Y2=1.35
r278 35 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.755 $Y=1.575
+ $X2=5.755 $Y2=1.74
r279 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.755
+ $Y=1.575 $X2=5.755 $Y2=1.575
r280 32 81 1.55539 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=5.755 $Y=1.04
+ $X2=5.755 $Y2=0.925
r281 32 34 29.6682 $w=1.98e-07 $l=5.35e-07 $layer=LI1_cond $X=5.755 $Y=1.04
+ $X2=5.755 $Y2=1.575
r282 28 30 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=1.89 $Y=2.63
+ $X2=3.095 $Y2=2.63
r283 27 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.805 $Y=2.545
+ $X2=1.89 $Y2=2.63
r284 27 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.805 $Y=2.545
+ $X2=1.805 $Y2=1.585
r285 24 40 46.1022 $w=3.8e-07 $l=3.15e-07 $layer=POLY_cond $X=9.56 $Y=1.665
+ $X2=9.56 $Y2=1.35
r286 24 25 48.9106 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=9.56 $Y=1.665
+ $X2=9.56 $Y2=1.855
r287 23 40 2.19534 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=9.56 $Y=1.335
+ $X2=9.56 $Y2=1.35
r288 22 23 43.0563 $w=3.8e-07 $l=1.5e-07 $layer=POLY_cond $X=9.54 $Y=1.185
+ $X2=9.54 $Y2=1.335
r289 19 25 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=9.445 $Y=2.475
+ $X2=9.445 $Y2=1.855
r290 16 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.405 $Y=0.755
+ $X2=9.405 $Y2=1.185
r291 13 72 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.88 $Y=0.57
+ $X2=6.88 $Y2=1
r292 9 68 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.665 $Y=2.48
+ $X2=5.665 $Y2=1.74
r293 2 30 600 $w=1.7e-07 $l=9.38576e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.795 $X2=3.095 $Y2=2.63
r294 1 75 91 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=2 $X=1.835
+ $Y=0.595 $X2=2.09 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_359_367# 1 2 7 9 11 14 18 22 26 31 33 37
+ 39 40 41 43 44 47 48 49 50 59 67 68 71
c195 68 0 1.33605e-19 $X=6.625 $Y=1.735
c196 49 0 1.0543e-19 $X=8.735 $Y=2.035
c197 44 0 8.37252e-20 $X=8.655 $Y=1.39
c198 43 0 1.37952e-19 $X=8.655 $Y=1.39
c199 26 0 3.15466e-20 $X=6.34 $Y=1.075
c200 18 0 1.7833e-19 $X=8.715 $Y=0.755
c201 11 0 1.24317e-19 $X=6.34 $Y=1.57
r202 66 68 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=6.485 $Y=1.735
+ $X2=6.625 $Y2=1.735
r203 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.485
+ $Y=1.735 $X2=6.485 $Y2=1.735
r204 63 66 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=6.34 $Y=1.735
+ $X2=6.485 $Y2=1.735
r205 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r206 57 67 13.0465 $w=2.63e-07 $l=3e-07 $layer=LI1_cond $X=6.517 $Y=2.035
+ $X2=6.517 $Y2=1.735
r207 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=2.035
+ $X2=6.48 $Y2=2.035
r208 53 71 36.1448 $w=3.28e-07 $l=1.035e-06 $layer=LI1_cond $X=3.095 $Y=2.035
+ $X2=3.095 $Y2=1
r209 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=2.035
+ $X2=3.12 $Y2=2.035
r210 50 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=2.035
+ $X2=6.48 $Y2=2.035
r211 49 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r212 49 50 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=6.625 $Y2=2.035
r213 48 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=2.035
+ $X2=3.12 $Y2=2.035
r214 47 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=2.035
+ $X2=6.48 $Y2=2.035
r215 47 48 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.335 $Y=2.035
+ $X2=3.265 $Y2=2.035
r216 46 53 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.095 $Y=2.195
+ $X2=3.095 $Y2=2.035
r217 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.655
+ $Y=1.39 $X2=8.655 $Y2=1.39
r218 41 60 9.24242 $w=2.97e-07 $l=3.13568e-07 $layer=LI1_cond $X=8.655 $Y=1.725
+ $X2=8.88 $Y2=1.937
r219 41 43 20.6414 $w=1.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.655 $Y=1.725
+ $X2=8.655 $Y2=1.39
r220 39 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.93 $Y=2.28
+ $X2=3.095 $Y2=2.195
r221 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.93 $Y=2.28
+ $X2=2.24 $Y2=2.28
r222 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.155 $Y=2.195
+ $X2=2.24 $Y2=2.28
r223 35 37 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.155 $Y=2.195
+ $X2=2.155 $Y2=2.07
r224 31 44 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.655 $Y=1.745
+ $X2=8.655 $Y2=1.39
r225 31 33 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=8.655 $Y=1.82
+ $X2=9.015 $Y2=1.82
r226 29 44 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=1.225
+ $X2=8.655 $Y2=1.39
r227 24 26 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.175 $Y=1.075
+ $X2=6.34 $Y2=1.075
r228 20 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.015 $Y=1.895
+ $X2=9.015 $Y2=1.82
r229 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.015 $Y=1.895
+ $X2=9.015 $Y2=2.475
r230 18 29 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=8.715 $Y=0.755
+ $X2=8.715 $Y2=1.225
r231 12 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.625 $Y=1.9
+ $X2=6.625 $Y2=1.735
r232 12 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.625 $Y=1.9
+ $X2=6.625 $Y2=2.48
r233 11 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.34 $Y=1.57
+ $X2=6.34 $Y2=1.735
r234 10 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.34 $Y=1.15
+ $X2=6.34 $Y2=1.075
r235 10 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=6.34 $Y=1.15
+ $X2=6.34 $Y2=1.57
r236 7 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.175 $Y=1 $X2=6.175
+ $Y2=1.075
r237 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.175 $Y=1 $X2=6.175
+ $Y2=0.57
r238 2 37 600 $w=1.7e-07 $l=4.62817e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.835 $X2=2.155 $Y2=2.07
r239 1 71 182 $w=1.7e-07 $l=4.77624e-07 $layer=licon1_NDIFF $count=1 $X=2.835
+ $Y=0.635 $X2=3.095 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%CI 3 6 7 9 12 14 16 17 20 25
c65 25 0 1.35641e-20 $X=8.17 $Y=1.35
c66 3 0 1.20808e-19 $X=7.27 $Y=2.335
r67 23 25 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=7.87 $Y=1.35 $X2=8.17
+ $Y2=1.35
r68 21 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.78 $Y=1.35 $X2=7.87
+ $Y2=1.35
r69 19 21 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.63 $Y=1.35
+ $X2=7.78 $Y2=1.35
r70 19 20 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.63 $Y=1.35
+ $X2=7.555 $Y2=1.35
r71 17 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.87
+ $Y=1.35 $X2=7.87 $Y2=1.35
r72 14 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.17 $Y=1.185
+ $X2=8.17 $Y2=1.35
r73 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.17 $Y=1.185
+ $X2=8.17 $Y2=0.655
r74 10 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.78 $Y=1.515
+ $X2=7.78 $Y2=1.35
r75 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.78 $Y=1.515
+ $X2=7.78 $Y2=2.465
r76 7 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.63 $Y=1.185
+ $X2=7.63 $Y2=1.35
r77 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.63 $Y=1.185 $X2=7.63
+ $Y2=0.755
r78 6 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.345 $Y=1.44
+ $X2=7.555 $Y2=1.44
r79 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.27 $Y=1.515
+ $X2=7.345 $Y2=1.44
r80 1 3 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.27 $Y=1.515 $X2=7.27
+ $Y2=2.335
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_1571_367# 1 2 3 12 14 16 18 21 25 29 34
+ 35 36 38 41 42 48 52
c122 35 0 1.44079e-19 $X=8.107 $Y=1.815
c123 21 0 1.20808e-19 $X=7.995 $Y=2.9
r124 49 52 4.44923 $w=3.25e-07 $l=3e-08 $layer=POLY_cond $X=10.125 $Y=1.665
+ $X2=10.155 $Y2=1.665
r125 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.125
+ $Y=1.59 $X2=10.125 $Y2=1.59
r126 45 48 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=9.94 $Y=1.59
+ $X2=10.125 $Y2=1.59
r127 41 43 9.70403 $w=5.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.76 $Y=2.2
+ $X2=9.76 $Y2=2.63
r128 41 42 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.76 $Y=2.2
+ $X2=9.76 $Y2=2.035
r129 38 39 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=8.382 $Y=0.88
+ $X2=8.382 $Y2=1.045
r130 35 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.3 $Y=1.815
+ $X2=8.3 $Y2=1.045
r131 34 35 9.86413 $w=5.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.107 $Y=1.98
+ $X2=8.107 $Y2=1.815
r132 31 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.94 $Y=1.755
+ $X2=9.94 $Y2=1.59
r133 31 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=9.94 $Y=1.755
+ $X2=9.94 $Y2=2.035
r134 30 36 4.93025 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=8.385 $Y=2.63
+ $X2=8.107 $Y2=2.63
r135 29 43 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=9.495 $Y=2.63
+ $X2=9.76 $Y2=2.63
r136 29 30 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=9.495 $Y=2.63
+ $X2=8.385 $Y2=2.63
r137 23 38 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=8.382 $Y=0.878
+ $X2=8.382 $Y2=0.88
r138 23 25 15.4118 $w=3.33e-07 $l=4.48e-07 $layer=LI1_cond $X=8.382 $Y=0.878
+ $X2=8.382 $Y2=0.43
r139 19 36 2.20108 $w=4.42e-07 $l=1.4854e-07 $layer=LI1_cond $X=7.995 $Y=2.715
+ $X2=8.107 $Y2=2.63
r140 19 21 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.995 $Y=2.715
+ $X2=7.995 $Y2=2.9
r141 18 36 2.20108 $w=4.42e-07 $l=8.5e-08 $layer=LI1_cond $X=8.107 $Y=2.545
+ $X2=8.107 $Y2=2.63
r142 17 34 2.41371 $w=5.53e-07 $l=1.12e-07 $layer=LI1_cond $X=8.107 $Y=2.092
+ $X2=8.107 $Y2=1.98
r143 17 18 9.76259 $w=5.53e-07 $l=4.53e-07 $layer=LI1_cond $X=8.107 $Y=2.092
+ $X2=8.107 $Y2=2.545
r144 14 52 51.9077 $w=3.25e-07 $l=4.54423e-07 $layer=POLY_cond $X=10.505
+ $Y=1.905 $X2=10.155 $Y2=1.665
r145 14 16 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.505 $Y=1.905
+ $X2=10.505 $Y2=2.515
r146 10 52 20.86 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.155 $Y=1.425
+ $X2=10.155 $Y2=1.665
r147 10 12 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=10.155 $Y=1.425
+ $X2=10.155 $Y2=0.755
r148 3 41 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.52
+ $Y=2.055 $X2=9.66 $Y2=2.2
r149 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.855
+ $Y=1.835 $X2=7.995 $Y2=1.98
r150 2 21 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=7.855
+ $Y=1.835 $X2=7.995 $Y2=2.9
r151 1 38 182 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_NDIFF $count=1 $X=8.245
+ $Y=0.235 $X2=8.385 $Y2=0.88
r152 1 25 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=8.245
+ $Y=0.235 $X2=8.385 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_1758_87# 1 2 7 9 12 17 19 20 21 24 27 28
+ 29 32 35 38 43
c102 38 0 1.57643e-19 $X=9.23 $Y=1.305
r103 42 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=11.025 $Y=1.35
+ $X2=11.04 $Y2=1.35
r104 36 38 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.01 $Y=1.305
+ $X2=9.23 $Y2=1.305
r105 33 42 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=10.865 $Y=1.35
+ $X2=11.025 $Y2=1.35
r106 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.865
+ $Y=1.35 $X2=10.865 $Y2=1.35
r107 30 32 24.3889 $w=2.13e-07 $l=4.55e-07 $layer=LI1_cond $X=10.867 $Y=0.895
+ $X2=10.867 $Y2=1.35
r108 28 30 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=10.76 $Y=0.81
+ $X2=10.867 $Y2=0.895
r109 28 29 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.76 $Y=0.81
+ $X2=10.375 $Y2=0.81
r110 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.29 $Y=0.725
+ $X2=10.375 $Y2=0.81
r111 26 27 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.29 $Y=0.435
+ $X2=10.29 $Y2=0.725
r112 22 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.23 $Y=1.39
+ $X2=9.23 $Y2=1.305
r113 22 24 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=9.23 $Y=1.39
+ $X2=9.23 $Y2=2.2
r114 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.205 $Y=0.35
+ $X2=10.29 $Y2=0.435
r115 20 21 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=10.205 $Y=0.35
+ $X2=9.095 $Y2=0.35
r116 19 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=1.22
+ $X2=9.01 $Y2=1.305
r117 19 35 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.01 $Y=1.22
+ $X2=9.01 $Y2=1.045
r118 15 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.93 $Y=0.88
+ $X2=8.93 $Y2=1.045
r119 15 17 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=8.93 $Y=0.88
+ $X2=8.93 $Y2=0.73
r120 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.93 $Y=0.435
+ $X2=9.095 $Y2=0.35
r121 14 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.93 $Y=0.435
+ $X2=8.93 $Y2=0.73
r122 10 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.04 $Y=1.515
+ $X2=11.04 $Y2=1.35
r123 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=11.04 $Y=1.515
+ $X2=11.04 $Y2=2.465
r124 7 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.025 $Y=1.185
+ $X2=11.025 $Y2=1.35
r125 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.025 $Y=1.185
+ $X2=11.025 $Y2=0.655
r126 2 24 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.055 $X2=9.23 $Y2=2.2
r127 1 17 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=8.79
+ $Y=0.435 $X2=8.93 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%VPWR 1 2 3 4 17 23 31 35 38 39 40 49 56 66
+ 67 70 73 76
r98 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r99 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r100 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 67 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r102 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r103 64 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.91 $Y=3.33
+ $X2=10.785 $Y2=3.33
r104 64 66 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.91 $Y=3.33
+ $X2=11.28 $Y2=3.33
r105 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r106 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r107 60 63 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r108 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r109 59 62 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r110 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=3.33
+ $X2=7.485 $Y2=3.33
r112 57 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.65 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 56 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.66 $Y=3.33
+ $X2=10.785 $Y2=3.33
r114 56 62 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.66 $Y=3.33
+ $X2=10.32 $Y2=3.33
r115 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=7.485 $Y2=3.33
r120 49 54 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 47 48 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r123 45 48 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r124 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 44 47 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 44 45 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 42 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r128 42 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 40 55 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6.96 $Y2=3.33
r130 40 52 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 38 47 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.565 $Y=3.33
+ $X2=4.56 $Y2=3.33
r132 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=3.33
+ $X2=4.73 $Y2=3.33
r133 37 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=5.04 $Y2=3.33
r134 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=4.73 $Y2=3.33
r135 33 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.785 $Y=3.245
+ $X2=10.785 $Y2=3.33
r136 33 35 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=10.785 $Y=3.245
+ $X2=10.785 $Y2=2.45
r137 29 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=3.245
+ $X2=7.485 $Y2=3.33
r138 29 31 42.6055 $w=3.28e-07 $l=1.22e-06 $layer=LI1_cond $X=7.485 $Y=3.245
+ $X2=7.485 $Y2=2.025
r139 26 28 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=4.73 $Y=2.425
+ $X2=4.73 $Y2=2.91
r140 23 26 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=4.73 $Y=1.94
+ $X2=4.73 $Y2=2.425
r141 21 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=3.245
+ $X2=4.73 $Y2=3.33
r142 21 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.73 $Y=3.245
+ $X2=4.73 $Y2=2.91
r143 17 20 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=0.82 $Y=2.125
+ $X2=0.82 $Y2=2.95
r144 15 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r145 15 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.95
r146 4 35 300 $w=1.7e-07 $l=5.43875e-07 $layer=licon1_PDIFF $count=2 $X=10.58
+ $Y=2.015 $X2=10.825 $Y2=2.45
r147 3 31 300 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=1.835 $X2=7.485 $Y2=2.025
r148 2 28 600 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.795 $X2=4.73 $Y2=2.91
r149 2 26 600 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.795 $X2=4.73 $Y2=2.425
r150 2 23 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.795 $X2=4.73 $Y2=1.94
r151 1 20 600 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.82 $Y2=2.95
r152 1 17 300 $w=1.7e-07 $l=3.84578e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.835 $X2=0.82 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_247_367# 1 2 3 4 16 18 21 25 26 29 34 35
+ 36 37
c74 25 0 2.02469e-20 $X=3.475 $Y=2.98
c75 21 0 1.47047e-19 $X=1.545 $Y=0.925
r76 35 36 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.455 $Y=1.855
+ $X2=1.455 $Y2=1.235
r77 34 37 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=3.64 $Y=1.94
+ $X2=3.64 $Y2=1.295
r78 32 34 33.351 $w=3.28e-07 $l=9.55e-07 $layer=LI1_cond $X=3.64 $Y=2.895
+ $X2=3.64 $Y2=1.94
r79 27 37 6.44801 $w=4.33e-07 $l=2.17e-07 $layer=LI1_cond $X=3.692 $Y=1.078
+ $X2=3.692 $Y2=1.295
r80 27 29 7.8949 $w=4.33e-07 $l=2.98e-07 $layer=LI1_cond $X=3.692 $Y=1.078
+ $X2=3.692 $Y2=0.78
r81 25 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.475 $Y=2.98
+ $X2=3.64 $Y2=2.895
r82 25 26 126.241 $w=1.68e-07 $l=1.935e-06 $layer=LI1_cond $X=3.475 $Y=2.98
+ $X2=1.54 $Y2=2.98
r83 19 36 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.54 $Y=1.065
+ $X2=1.54 $Y2=1.235
r84 19 21 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.54 $Y=1.065
+ $X2=1.54 $Y2=0.925
r85 16 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=2.02
+ $X2=1.375 $Y2=1.855
r86 16 18 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.375 $Y=2.02
+ $X2=1.375 $Y2=2.69
r87 14 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.375 $Y=2.895
+ $X2=1.54 $Y2=2.98
r88 14 18 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.375 $Y=2.895
+ $X2=1.375 $Y2=2.69
r89 4 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.5
+ $Y=1.795 $X2=3.64 $Y2=1.94
r90 3 18 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.835 $X2=1.375 $Y2=2.69
r91 3 16 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.835 $X2=1.375 $Y2=2.02
r92 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.605
+ $Y=0.635 $X2=3.745 $Y2=0.78
r93 1 21 182 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.595 $X2=1.545 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_1034_380# 1 2 9 11 15 16 17 19
c51 19 0 1.62544e-19 $X=5.96 $Y=0.445
c52 17 0 3.15466e-20 $X=5.31 $Y=1.88
r53 19 21 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=5.96 $Y=0.445 $X2=5.96
+ $Y2=0.545
r54 15 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=0.545
+ $X2=5.96 $Y2=0.545
r55 15 16 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.795 $Y=0.545
+ $X2=5.475 $Y2=0.545
r56 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.39 $Y=0.63
+ $X2=5.475 $Y2=0.545
r57 13 17 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=5.39 $Y=0.63
+ $X2=5.39 $Y2=1.88
r58 9 17 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.31 $Y=2.045
+ $X2=5.31 $Y2=1.88
r59 9 11 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.31 $Y=2.045
+ $X2=5.31 $Y2=2.4
r60 2 11 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=5.17
+ $Y=1.9 $X2=5.31 $Y2=2.4
r61 2 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.9 $X2=5.31 $Y2=2.045
r62 1 19 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=5.82
+ $Y=0.25 $X2=5.96 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%COUT_N 1 2 9 14 15 18 20
c59 18 0 1.0217e-19 $X=6.39 $Y=1.305
c60 14 0 1.47098e-19 $X=6.39 $Y=1.22
r61 22 25 2.39469 $w=3.83e-07 $l=8e-08 $layer=LI1_cond $X=6.39 $Y=0.457 $X2=6.47
+ $Y2=0.457
r62 20 25 0.299336 $w=3.83e-07 $l=1e-08 $layer=LI1_cond $X=6.48 $Y=0.457
+ $X2=6.47 $Y2=0.457
r63 16 18 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.12 $Y=1.305
+ $X2=6.39 $Y2=1.305
r64 14 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.22
+ $X2=6.39 $Y2=1.305
r65 13 22 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=6.39 $Y=0.65
+ $X2=6.39 $Y2=0.457
r66 13 14 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.39 $Y=0.65
+ $X2=6.39 $Y2=1.22
r67 11 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=1.39
+ $X2=6.12 $Y2=1.305
r68 11 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.12 $Y=1.39
+ $X2=6.12 $Y2=2.04
r69 9 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.04 $Y=2.205
+ $X2=6.04 $Y2=2.04
r70 2 9 300 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=2 $X=5.74
+ $Y=2.06 $X2=6.04 $Y2=2.205
r71 1 25 182 $w=1.7e-07 $l=3.05778e-07 $layer=licon1_NDIFF $count=1 $X=6.25
+ $Y=0.25 $X2=6.47 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_1340_412# 1 2 9 13 15
r45 15 18 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=7.35 $Y=0.43 $X2=7.35
+ $Y2=0.93
r46 13 18 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=7.35 $Y=1.51
+ $X2=7.35 $Y2=0.93
r47 9 11 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=6.985 $Y=1.98
+ $X2=6.985 $Y2=2.755
r48 7 13 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.985 $Y=1.595
+ $X2=7.35 $Y2=1.595
r49 7 9 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=6.985 $Y=1.68 $X2=6.985
+ $Y2=1.98
r50 2 11 400 $w=1.7e-07 $l=8.0827e-07 $layer=licon1_PDIFF $count=1 $X=6.7
+ $Y=2.06 $X2=6.945 $Y2=2.755
r51 2 9 400 $w=1.7e-07 $l=2.82179e-07 $layer=licon1_PDIFF $count=1 $X=6.7
+ $Y=2.06 $X2=6.945 $Y2=1.98
r52 1 18 182 $w=1.7e-07 $l=8.38928e-07 $layer=licon1_NDIFF $count=1 $X=6.955
+ $Y=0.25 $X2=7.31 $Y2=0.93
r53 1 15 182 $w=1.7e-07 $l=4.35804e-07 $layer=licon1_NDIFF $count=1 $X=6.955
+ $Y=0.25 $X2=7.31 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%A_1708_411# 1 2 3 10 16 18 19 23 28 29
r60 28 29 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=10.392 $Y=1.935
+ $X2=10.392 $Y2=2.105
r61 26 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.495 $Y=1.245
+ $X2=10.495 $Y2=1.935
r62 23 25 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=10.33 $Y=2.16
+ $X2=10.33 $Y2=2.87
r63 23 29 2.53537 $w=2.48e-07 $l=5.5e-08 $layer=LI1_cond $X=10.33 $Y=2.16
+ $X2=10.33 $Y2=2.105
r64 21 25 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=10.33 $Y=2.895
+ $X2=10.33 $Y2=2.87
r65 18 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.41 $Y=1.16
+ $X2=10.495 $Y2=1.245
r66 18 19 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.41 $Y=1.16
+ $X2=10.025 $Y2=1.16
r67 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.94 $Y=1.075
+ $X2=10.025 $Y2=1.16
r68 14 16 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.94 $Y=1.075
+ $X2=9.94 $Y2=0.855
r69 10 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.205 $Y=2.98
+ $X2=10.33 $Y2=2.895
r70 10 12 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=10.205 $Y=2.98
+ $X2=8.685 $Y2=2.98
r71 3 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.145
+ $Y=2.015 $X2=10.29 $Y2=2.87
r72 3 23 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.145
+ $Y=2.015 $X2=10.29 $Y2=2.16
r73 2 12 600 $w=1.7e-07 $l=9.94862e-07 $layer=licon1_PDIFF $count=1 $X=8.54
+ $Y=2.055 $X2=8.685 $Y2=2.98
r74 1 16 182 $w=1.7e-07 $l=6.36239e-07 $layer=licon1_NDIFF $count=1 $X=9.48
+ $Y=0.435 $X2=9.94 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%SUM 1 2 7 8 9 10 11 12 13 22
r12 13 40 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=11.287 $Y=2.775
+ $X2=11.287 $Y2=2.9
r13 12 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.287 $Y=2.405
+ $X2=11.287 $Y2=2.775
r14 11 12 18.4826 $w=2.63e-07 $l=4.25e-07 $layer=LI1_cond $X=11.287 $Y=1.98
+ $X2=11.287 $Y2=2.405
r15 10 11 13.6989 $w=2.63e-07 $l=3.15e-07 $layer=LI1_cond $X=11.287 $Y=1.665
+ $X2=11.287 $Y2=1.98
r16 9 10 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.287 $Y=1.295
+ $X2=11.287 $Y2=1.665
r17 8 9 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.287 $Y=0.925
+ $X2=11.287 $Y2=1.295
r18 7 8 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.287 $Y=0.555
+ $X2=11.287 $Y2=0.925
r19 7 22 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=11.287 $Y=0.555
+ $X2=11.287 $Y2=0.43
r20 2 40 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=11.115
+ $Y=1.835 $X2=11.255 $Y2=2.9
r21 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.115
+ $Y=1.835 $X2=11.255 $Y2=1.98
r22 1 22 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=11.1
+ $Y=0.235 $X2=11.24 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__FAHCON_1%VGND 1 2 3 4 17 21 25 31 34 35 36 38 46 59
+ 60 63 66 69
r112 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r113 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r114 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r115 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r116 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r117 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r118 54 57 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r119 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r120 53 56 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.32
+ $Y2=0
r121 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r122 51 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.035 $Y=0 $X2=7.91
+ $Y2=0
r123 51 53 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.035 $Y=0 $X2=8.4
+ $Y2=0
r124 50 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r125 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r126 47 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=4.97
+ $Y2=0
r127 47 49 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=5.095 $Y=0
+ $X2=7.44 $Y2=0
r128 46 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.785 $Y=0 $X2=7.91
+ $Y2=0
r129 46 49 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.785 $Y=0 $X2=7.44
+ $Y2=0
r130 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r131 44 45 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r132 42 45 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r133 42 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r134 41 44 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r135 41 42 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r136 39 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0 $X2=0.755
+ $Y2=0
r137 39 41 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=1.2
+ $Y2=0
r138 38 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.845 $Y=0 $X2=4.97
+ $Y2=0
r139 38 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.845 $Y=0
+ $X2=4.56 $Y2=0
r140 36 50 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r141 36 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=0 $X2=5.04
+ $Y2=0
r142 34 56 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.61 $Y=0
+ $X2=10.32 $Y2=0
r143 34 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.61 $Y=0
+ $X2=10.735 $Y2=0
r144 33 59 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=0
+ $X2=11.28 $Y2=0
r145 33 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.86 $Y=0
+ $X2=10.735 $Y2=0
r146 29 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.735 $Y=0.085
+ $X2=10.735 $Y2=0
r147 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=10.735 $Y=0.085
+ $X2=10.735 $Y2=0.38
r148 25 27 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=7.91 $Y=0.38
+ $X2=7.91 $Y2=0.835
r149 23 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r150 23 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.38
r151 19 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=0.085
+ $X2=4.97 $Y2=0
r152 19 21 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=4.97 $Y=0.085
+ $X2=4.97 $Y2=0.395
r153 15 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r154 15 17 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.595
r155 4 31 182 $w=1.7e-07 $l=4.91732e-07 $layer=licon1_NDIFF $count=1 $X=10.23
+ $Y=0.435 $X2=10.695 $Y2=0.38
r156 3 27 182 $w=1.7e-07 $l=5.07937e-07 $layer=licon1_NDIFF $count=1 $X=7.705
+ $Y=0.435 $X2=7.95 $Y2=0.835
r157 3 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.705
+ $Y=0.435 $X2=7.95 $Y2=0.38
r158 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.87
+ $Y=0.25 $X2=5.01 $Y2=0.395
r159 1 17 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.395 $X2=0.755 $Y2=0.595
.ends

