* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxtp_lp D GATE VGND VNB VPB VPWR Q
X0 a_824_491# a_463_491# a_933_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_114_102# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_463_491# a_27_102# a_550_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VPWR a_350_102# a_746_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_746_491# a_27_102# a_824_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_27_102# GATE a_114_102# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR D a_278_470# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_1198_47# a_824_491# a_1027_407# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_114_470# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VGND D a_278_102# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_1027_407# a_1474_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_1474_367# a_1027_407# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_463_491# a_27_102# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_278_470# D a_350_102# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_790_47# a_463_491# a_824_491# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_824_491# a_1198_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_824_491# a_27_102# a_982_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1474_53# a_1027_407# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_278_102# D a_350_102# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_350_102# a_790_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_933_535# a_1027_407# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_27_102# GATE a_114_470# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_982_47# a_1027_407# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR a_824_491# a_1204_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_1204_367# a_824_491# a_1027_407# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_550_491# a_27_102# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VGND a_1027_407# a_1474_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_584_47# a_27_102# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
