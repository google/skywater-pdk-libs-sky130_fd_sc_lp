* File: sky130_fd_sc_lp__a21boi_2.spice
* Created: Fri Aug 28 09:50:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21boi_2.pex.spice"
.subckt sky130_fd_sc_lp__a21boi_2  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_B1_N_M1012_g N_A_119_500#_M1012_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_119_500#_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=3.564 M=1 R=5.6 SA=75000.5
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1002_d N_A_119_500#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9 SB=75002.1
+ A=0.126 P=1.98 MULT=1
MM1009 N_A_502_65#_M1009_d N_A2_M1009_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.4
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g N_A_502_65#_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75001.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1003_d N_A1_M1005_g N_A_502_65#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1013 N_A_502_65#_M1005_s N_A2_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_A_119_500#_M1011_d N_B1_N_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_231_367#_M1004_d N_A_119_500#_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1010 N_A_231_367#_M1010_d N_A_119_500#_M1010_g N_Y_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_231_367#_M1010_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1001_d N_A1_M1000_g N_A_231_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75001.6 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_231_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1006_d N_A2_M1008_g N_A_231_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
c_49 VNB 0 1.37558e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a21boi_2.pxi.spice"
*
.ends
*
*
