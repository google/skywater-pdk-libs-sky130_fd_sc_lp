* File: sky130_fd_sc_lp__invlp_4.pex.spice
* Created: Wed Sep  2 09:57:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVLP_4%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 70 71 73 74 75 108 109 119
c169 63 0 1.66076e-19 $X=3.785 $Y=0.685
c170 35 0 6.94355e-20 $X=2.305 $Y=2.465
c171 15 0 5.41714e-20 $X=0.945 $Y=2.465
r172 104 105 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.735 $Y=1.51
+ $X2=3.785 $Y2=1.51
r173 103 104 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.305 $Y=1.51
+ $X2=3.735 $Y2=1.51
r174 102 103 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.285 $Y=1.51
+ $X2=3.305 $Y2=1.51
r175 99 100 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.785 $Y=1.51
+ $X2=2.805 $Y2=1.51
r176 98 108 0.847774 $w=4.33e-07 $l=3.2e-08 $layer=LI1_cond $X=2.57 $Y=1.562
+ $X2=2.538 $Y2=1.562
r177 97 99 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.57 $Y=1.51
+ $X2=2.785 $Y2=1.51
r178 97 98 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.51 $X2=2.57 $Y2=1.51
r179 95 97 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.355 $Y=1.51
+ $X2=2.57 $Y2=1.51
r180 94 95 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.305 $Y=1.51
+ $X2=2.355 $Y2=1.51
r181 93 108 8.15983 $w=4.33e-07 $l=3.08e-07 $layer=LI1_cond $X=2.23 $Y=1.562
+ $X2=2.538 $Y2=1.562
r182 92 94 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.305 $Y2=1.51
r183 92 93 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.51 $X2=2.23 $Y2=1.51
r184 90 92 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.925 $Y=1.51
+ $X2=2.23 $Y2=1.51
r185 89 90 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.805 $Y=1.51
+ $X2=1.925 $Y2=1.51
r186 87 89 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.55 $Y=1.51
+ $X2=1.805 $Y2=1.51
r187 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.51 $X2=1.55 $Y2=1.51
r188 85 87 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.495 $Y=1.51
+ $X2=1.55 $Y2=1.51
r189 84 85 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.375 $Y=1.51
+ $X2=1.495 $Y2=1.51
r190 83 84 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.945 $Y=1.51
+ $X2=1.375 $Y2=1.51
r191 82 83 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.945 $Y2=1.51
r192 81 82 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.515 $Y=1.51
+ $X2=0.925 $Y2=1.51
r193 79 81 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.515 $Y2=1.51
r194 75 119 3.74573 $w=4.33e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=2.755 $Y2=1.562
r195 75 98 1.85451 $w=4.33e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=2.57 $Y2=1.562
r196 74 93 1.85451 $w=4.33e-07 $l=7e-08 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=2.23 $Y2=1.562
r197 74 109 4.23887 $w=4.33e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=2 $Y2=1.562
r198 73 109 9.05536 $w=4.35e-07 $l=3.2e-07 $layer=LI1_cond $X=1.68 $Y=1.562
+ $X2=2 $Y2=1.562
r199 73 88 3.92574 $w=4.04e-07 $l=1.3e-07 $layer=LI1_cond $X=1.68 $Y=1.562
+ $X2=1.55 $Y2=1.562
r200 71 105 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.93 $Y=1.51
+ $X2=3.785 $Y2=1.51
r201 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.93
+ $Y=1.51 $X2=3.93 $Y2=1.51
r202 68 102 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.91 $Y=1.51
+ $X2=3.285 $Y2=1.51
r203 68 100 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=2.91 $Y=1.51
+ $X2=2.805 $Y2=1.51
r204 67 70 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=2.91 $Y=1.51
+ $X2=3.93 $Y2=1.51
r205 67 119 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.91 $Y=1.51
+ $X2=2.755 $Y2=1.51
r206 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.91
+ $Y=1.51 $X2=2.91 $Y2=1.51
r207 61 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.345
+ $X2=3.785 $Y2=1.51
r208 61 63 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.785 $Y=1.345
+ $X2=3.785 $Y2=0.685
r209 57 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.735 $Y=1.675
+ $X2=3.735 $Y2=1.51
r210 57 59 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.735 $Y=1.675
+ $X2=3.735 $Y2=2.465
r211 53 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.675
+ $X2=3.305 $Y2=1.51
r212 53 55 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.305 $Y=1.675
+ $X2=3.305 $Y2=2.465
r213 49 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.345
+ $X2=3.285 $Y2=1.51
r214 49 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.285 $Y=1.345
+ $X2=3.285 $Y2=0.685
r215 45 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.675
+ $X2=2.805 $Y2=1.51
r216 45 47 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.805 $Y=1.675
+ $X2=2.805 $Y2=2.465
r217 41 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.345
+ $X2=2.785 $Y2=1.51
r218 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.785 $Y=1.345
+ $X2=2.785 $Y2=0.685
r219 37 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.345
+ $X2=2.355 $Y2=1.51
r220 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.355 $Y=1.345
+ $X2=2.355 $Y2=0.685
r221 33 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.675
+ $X2=2.305 $Y2=1.51
r222 33 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.305 $Y=1.675
+ $X2=2.305 $Y2=2.465
r223 29 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.345
+ $X2=1.925 $Y2=1.51
r224 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.925 $Y=1.345
+ $X2=1.925 $Y2=0.685
r225 25 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.675
+ $X2=1.805 $Y2=1.51
r226 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.805 $Y=1.675
+ $X2=1.805 $Y2=2.465
r227 21 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.345
+ $X2=1.495 $Y2=1.51
r228 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.495 $Y=1.345
+ $X2=1.495 $Y2=0.685
r229 17 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=1.51
r230 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=2.465
r231 13 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.675
+ $X2=0.945 $Y2=1.51
r232 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.945 $Y=1.675
+ $X2=0.945 $Y2=2.465
r233 9 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=1.51
r234 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=0.685
r235 5 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.675
+ $X2=0.515 $Y2=1.51
r236 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.515 $Y=1.675
+ $X2=0.515 $Y2=2.465
r237 1 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=1.51
r238 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_4%VPWR 1 2 3 10 12 18 20 22 26 28 33 42 46
r57 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 37 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 34 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.12 $Y2=3.33
r63 34 36 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 33 45 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.087 $Y2=3.33
r65 33 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 32 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 29 39 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.192 $Y2=3.33
r70 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 28 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.12 $Y2=3.33
r72 28 31 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 26 37 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r74 26 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 22 25 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=4.02 $Y=2.01
+ $X2=4.02 $Y2=2.95
r76 20 45 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.087 $Y2=3.33
r77 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=2.95
r78 16 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=3.33
r79 16 18 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=2.87
r80 12 15 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=0.26 $Y=1.98
+ $X2=0.26 $Y2=2.95
r81 10 39 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.192 $Y2=3.33
r82 10 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r83 3 25 400 $w=1.7e-07 $l=1.21547e-06 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.835 $X2=4.02 $Y2=2.95
r84 3 22 400 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.835 $X2=4.02 $Y2=2.01
r85 2 18 600 $w=1.7e-07 $l=1.10278e-06 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.835 $X2=1.16 $Y2=2.87
r86 1 15 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.3 $Y2=2.95
r87 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.3 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_4%A_118_367# 1 2 3 4 15 19 21 22 23 24 27 29
+ 31 33 36 39
c58 24 0 5.41714e-20 $X=1.755 $Y=2.99
c59 21 0 6.94355e-20 $X=1.59 $Y=2.46
r60 31 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=2.905
+ $X2=3.56 $Y2=2.99
r61 31 33 41.2575 $w=2.48e-07 $l=8.95e-07 $layer=LI1_cond $X=3.56 $Y=2.905
+ $X2=3.56 $Y2=2.01
r62 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=2.99
+ $X2=2.59 $Y2=2.99
r63 29 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.435 $Y=2.99
+ $X2=3.56 $Y2=2.99
r64 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.435 $Y=2.99
+ $X2=2.755 $Y2=2.99
r65 25 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.905
+ $X2=2.59 $Y2=2.99
r66 25 27 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.59 $Y=2.905
+ $X2=2.59 $Y2=2.455
r67 23 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=2.99
+ $X2=2.59 $Y2=2.99
r68 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.425 $Y=2.99
+ $X2=1.755 $Y2=2.99
r69 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.755 $Y2=2.99
r70 21 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.46 $X2=1.59
+ $Y2=2.375
r71 21 22 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.59 $Y=2.46
+ $X2=1.59 $Y2=2.905
r72 20 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=2.375
+ $X2=0.69 $Y2=2.375
r73 19 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=2.375
+ $X2=1.59 $Y2=2.375
r74 19 20 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.425 $Y=2.375
+ $X2=0.815 $Y2=2.375
r75 13 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.29 $X2=0.69
+ $Y2=2.375
r76 13 15 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.69 $Y=2.29
+ $X2=0.69 $Y2=1.98
r77 4 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.835 $X2=3.52 $Y2=2.91
r78 4 33 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.835 $X2=3.52 $Y2=2.01
r79 3 27 300 $w=1.7e-07 $l=7.17356e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=1.835 $X2=2.59 $Y2=2.455
r80 2 38 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=2.455
r81 1 36 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.835 $X2=0.73 $Y2=2.445
r82 1 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.835 $X2=0.73 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_4%Y 1 2 3 4 14 15 17 18 23 25 27 31 33 35 37
+ 40 42 43 46
c85 31 0 1.66076e-19 $X=3.07 $Y=0.86
r86 40 46 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=1.295
+ $X2=0.72 $Y2=1.295
r87 37 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.13 $Y=1.09
+ $X2=1.13 $Y2=1.295
r88 33 45 3.01048 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=3.09 $Y=2.12
+ $X2=3.09 $Y2=1.982
r89 33 35 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.09 $Y=2.12
+ $X2=3.09 $Y2=2.57
r90 29 31 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=3.07 $Y=1.005
+ $X2=3.07 $Y2=0.86
r91 28 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=2.09 $Y2=2.035
r92 27 45 4.75569 $w=1.7e-07 $l=1.89658e-07 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=3.09 $Y2=1.982
r93 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=2.255 $Y2=2.035
r94 26 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=1.09
+ $X2=2.14 $Y2=1.09
r95 25 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.905 $Y=1.09
+ $X2=3.07 $Y2=1.005
r96 25 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.905 $Y=1.09
+ $X2=2.225 $Y2=1.09
r97 21 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.005
+ $X2=2.14 $Y2=1.09
r98 21 23 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.14 $Y=1.005
+ $X2=2.14 $Y2=0.86
r99 17 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=2.035
+ $X2=2.09 $Y2=2.035
r100 17 18 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.925 $Y=2.035
+ $X2=1.215 $Y2=2.035
r101 16 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=1.09
+ $X2=1.13 $Y2=1.09
r102 15 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.09
+ $X2=2.14 $Y2=1.09
r103 15 16 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.055 $Y=1.09
+ $X2=1.215 $Y2=1.09
r104 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.13 $Y=1.95
+ $X2=1.215 $Y2=2.035
r105 13 40 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.13 $Y=1.41
+ $X2=1.13 $Y2=1.295
r106 13 14 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.13 $Y=1.41
+ $X2=1.13 $Y2=1.95
r107 4 45 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.835 $X2=3.09 $Y2=2.01
r108 4 35 600 $w=1.7e-07 $l=8.33412e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.835 $X2=3.09 $Y2=2.57
r109 3 42 300 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_PDIFF $count=2 $X=1.88
+ $Y=1.835 $X2=2.09 $Y2=2.115
r110 2 31 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.265 $X2=3.07 $Y2=0.86
r111 1 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.265 $X2=2.14 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_4%VGND 1 2 3 10 12 16 18 20 22 24 29 41 45
r54 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r55 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 36 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r58 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r59 33 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r60 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r61 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r62 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r63 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r64 29 44 3.96406 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=4.117
+ $Y2=0
r65 29 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=3.6
+ $Y2=0
r66 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r67 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r68 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 25 38 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r70 25 27 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r71 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r72 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r73 22 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r74 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r75 18 44 3.1791 $w=2.5e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.117 $Y2=0
r76 18 20 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.41
r77 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r78 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.41
r79 10 38 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r80 10 12 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.41
r81 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.265 $X2=4 $Y2=0.41
r82 2 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.265 $X2=1.21 $Y2=0.41
r83 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.265 $X2=0.28 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_4%A_114_53# 1 2 3 4 15 17 18 22 23 24 27 32 34
r71 28 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0.34
+ $X2=2.57 $Y2=0.34
r72 27 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0.34
+ $X2=3.57 $Y2=0.34
r73 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.405 $Y=0.34
+ $X2=2.735 $Y2=0.34
r74 23 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=0.34
+ $X2=2.57 $Y2=0.34
r75 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.405 $Y=0.34
+ $X2=1.875 $Y2=0.34
r76 20 22 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.71 $Y=0.665
+ $X2=1.71 $Y2=0.545
r77 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.71 $Y=0.425
+ $X2=1.875 $Y2=0.34
r78 19 22 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.71 $Y=0.425
+ $X2=1.71 $Y2=0.545
r79 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.545 $Y=0.75
+ $X2=1.71 $Y2=0.665
r80 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=0.75
+ $X2=0.875 $Y2=0.75
r81 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=0.665
+ $X2=0.875 $Y2=0.75
r82 13 15 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.71 $Y=0.665
+ $X2=0.71 $Y2=0.42
r83 4 34 91 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=2 $X=3.36
+ $Y=0.265 $X2=3.57 $Y2=0.42
r84 3 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.265 $X2=2.57 $Y2=0.41
r85 2 22 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.265 $X2=1.71 $Y2=0.545
r86 1 15 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.265 $X2=0.71 $Y2=0.42
.ends

