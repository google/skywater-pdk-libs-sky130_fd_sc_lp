* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__busdriver2_20 A TE_B VGND VNB VPB VPWR Z
X0 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X1 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 VPWR a_114_47# a_286_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X3 VPWR a_114_47# a_286_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X4 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X5 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X7 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X8 VGND TE_B a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X14 VGND A a_1909_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X16 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X20 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X21 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X24 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X25 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X26 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 a_114_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X28 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X29 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 a_286_367# a_114_47# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X31 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X32 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X33 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X34 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 a_286_367# a_114_47# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X36 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X37 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X39 a_286_367# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X40 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X41 VGND A a_1909_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X42 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X43 a_114_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X44 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X45 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X46 a_1909_21# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X47 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X48 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X49 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X50 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X51 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X52 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X53 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X54 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X55 a_1909_21# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X56 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X57 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X58 VGND a_114_47# a_286_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X59 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X60 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X61 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X62 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X63 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X64 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X65 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X66 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X67 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X68 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X69 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X70 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X71 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X72 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X73 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X74 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X75 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X76 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X77 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X78 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X79 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X80 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X81 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X82 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X83 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X84 VPWR TE_B a_114_47# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X85 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X86 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X87 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X88 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X89 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
