* File: sky130_fd_sc_lp__mux2i_4.spice
* Created: Wed Sep  2 10:01:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2i_4.pex.spice"
.subckt sky130_fd_sc_lp__mux2i_4  VNB VPB A0 A1 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1005 N_A_110_69#_M1005_d N_A0_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1020 N_A_110_69#_M1005_d N_A0_M1020_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.6
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1024 N_A_110_69#_M1024_d N_A0_M1024_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75002.7
+ A=0.126 P=1.98 MULT=1
MM1029 N_A_110_69#_M1024_d N_A0_M1029_g N_Y_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1029_s N_A1_M1002_g N_A_470_69#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6 SA=75002
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1018 N_Y_M1018_d N_A1_M1018_g N_A_470_69#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6 SA=75002.6
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1019 N_Y_M1018_d N_A1_M1019_g N_A_470_69#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6 SA=75003
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1030 N_Y_M1030_d N_A1_M1030_g N_A_470_69#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.20075 PD=2.25 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6 SA=75003.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_S_M1010_g N_A_470_69#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_S_M1012_g N_A_470_69#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1012_d N_S_M1031_g N_A_470_69#_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1033 N_VGND_M1033_d N_S_M1033_g N_A_470_69#_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1033_d N_A_1418_21#_M1006_g N_A_110_69#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_1418_21#_M1009_g N_A_110_69#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1027 N_VGND_M1009_d N_A_1418_21#_M1027_g N_A_110_69#_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1028 N_VGND_M1028_d N_A_1418_21#_M1028_g N_A_110_69#_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_A_1418_21#_M1003_d N_S_M1003_g N_VGND_M1028_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_A0_M1001_g N_A_126_367#_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1014_d N_A0_M1014_g N_A_126_367#_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1014_d N_A0_M1016_g N_A_126_367#_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1025 N_Y_M1025_d N_A0_M1025_g N_A_126_367#_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1025_d N_A1_M1007_g N_A_470_367#_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1013 N_Y_M1013_d N_A1_M1013_g N_A_470_367#_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1023 N_Y_M1013_d N_A1_M1023_g N_A_470_367#_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1032 N_Y_M1032_d N_A1_M1032_g N_A_470_367#_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_S_M1000_g N_A_126_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.53155 AS=0.1764 PD=3.51 PS=1.54 NRD=18.7544 NRS=0 M=1 R=8.4 SA=75000.3
+ SB=75003.8 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_S_M1004_g N_A_126_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1004_d N_S_M1017_g N_A_126_367#_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.189 PD=1.54 PS=1.56 NRD=0 NRS=0 M=1 R=8.4 SA=75001.2 SB=75003
+ A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_S_M1026_g N_A_126_367#_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.189 PD=1.54 PS=1.56 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75001.6
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1026_d N_A_1418_21#_M1008_g N_A_470_367#_M1008_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.1 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_1418_21#_M1011_g N_A_470_367#_M1008_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75002.5 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1011_d N_A_1418_21#_M1021_g N_A_470_367#_M1021_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75003.1 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_1418_21#_M1022_g N_A_470_367#_M1021_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.189 AS=0.1764 PD=1.56 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75003.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_1418_21#_M1015_d N_S_M1015_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.189 PD=3.05 PS=1.56 NRD=0 NRS=0 M=1 R=8.4 SA=75004 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=18.6127 P=23.69
*
.include "sky130_fd_sc_lp__mux2i_4.pxi.spice"
*
.ends
*
*
