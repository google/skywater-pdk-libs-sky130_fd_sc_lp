* File: sky130_fd_sc_lp__dlxbn_2.pex.spice
* Created: Fri Aug 28 10:27:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXBN_2%D 3 6 9 10 11 12 13 17
c33 17 0 9.39864e-20 $X=0.545 $Y=1.375
r34 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.545
+ $Y=1.375 $X2=0.545 $Y2=1.375
r35 13 18 7.54049 $w=4.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.375
r36 12 18 2.08014 $w=4.58e-07 $l=8e-08 $layer=LI1_cond $X=0.68 $Y=1.295 $X2=0.68
+ $Y2=1.375
r37 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.545 $Y=1.715
+ $X2=0.545 $Y2=1.375
r38 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.715
+ $X2=0.545 $Y2=1.88
r39 9 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.21
+ $X2=0.545 $Y2=1.375
r40 6 11 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.635 $Y=2.395
+ $X2=0.635 $Y2=1.88
r41 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.565 $Y=0.89
+ $X2=0.565 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%GATE_N 1 3 6 8 11 12 13 16 17
c41 17 0 9.21549e-20 $X=1.445 $Y=0.405
r42 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=0.405
+ $X2=1.445 $Y2=0.57
r43 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=0.405 $X2=1.445 $Y2=0.405
r44 13 17 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.2 $Y=0.485
+ $X2=1.445 $Y2=0.485
r45 11 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.535 $Y=1.21
+ $X2=1.535 $Y2=0.57
r46 9 12 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.14 $Y=1.285
+ $X2=1.03 $Y2=1.285
r47 8 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.46 $Y=1.285
+ $X2=1.535 $Y2=1.21
r48 8 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.46 $Y=1.285 $X2=1.14
+ $Y2=1.285
r49 4 12 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.065 $Y=1.36
+ $X2=1.03 $Y2=1.285
r50 4 6 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=1.065 $Y=1.36
+ $X2=1.065 $Y2=2.395
r51 1 12 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=0.995 $Y=1.21
+ $X2=1.03 $Y2=1.285
r52 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.995 $Y=1.21
+ $X2=0.995 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%A_214_136# 1 2 9 11 14 18 20 24 27 28 29 30
+ 31 40 44 45
c112 44 0 1.53527e-19 $X=2.995 $Y=1.25
c113 40 0 9.39864e-20 $X=1.615 $Y=1.17
c114 31 0 1.53889e-19 $X=2.935 $Y=1.17
c115 30 0 6.46996e-20 $X=2.112 $Y=2.295
c116 9 0 9.21549e-20 $X=2.11 $Y=0.73
r117 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.995
+ $Y=1.25 $X2=2.995 $Y2=1.25
r118 40 42 9.93665 $w=8.84e-07 $l=7.2e-07 $layer=LI1_cond $X=1.615 $Y=1.17
+ $X2=1.615 $Y2=1.89
r119 38 40 0.552036 $w=8.84e-07 $l=4e-08 $layer=LI1_cond $X=1.615 $Y=1.13
+ $X2=1.615 $Y2=1.17
r120 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.985
+ $Y=1.13 $X2=1.985 $Y2=1.13
r121 36 38 2.82919 $w=8.84e-07 $l=4.97041e-07 $layer=LI1_cond $X=1.21 $Y=0.925
+ $X2=1.615 $Y2=1.13
r122 32 40 5.25053 $w=4.1e-07 $l=5.7e-07 $layer=LI1_cond $X=2.185 $Y=1.17
+ $X2=1.615 $Y2=1.17
r123 31 44 2.87083 $w=4.1e-07 $l=1.37e-07 $layer=LI1_cond $X=2.935 $Y=1.17
+ $X2=3.072 $Y2=1.17
r124 31 32 21.0813 $w=4.08e-07 $l=7.5e-07 $layer=LI1_cond $X=2.935 $Y=1.17
+ $X2=2.185 $Y2=1.17
r125 29 30 42.7811 $w=2.25e-07 $l=1.5e-07 $layer=POLY_cond $X=2.112 $Y=2.145
+ $X2=2.112 $Y2=2.295
r126 28 29 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.075 $Y=1.635
+ $X2=2.075 $Y2=2.145
r127 27 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.985 $Y=1.47
+ $X2=1.985 $Y2=1.13
r128 27 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.47
+ $X2=1.985 $Y2=1.635
r129 22 24 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.77 $Y=1.755
+ $X2=3.77 $Y2=2.665
r130 21 45 59.3768 $w=2.76e-07 $l=3.4e-07 $layer=POLY_cond $X=2.995 $Y=1.59
+ $X2=2.995 $Y2=1.25
r131 20 22 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.695 $Y=1.59
+ $X2=3.77 $Y2=1.755
r132 20 21 93.5508 $w=3.3e-07 $l=5.35e-07 $layer=POLY_cond $X=3.695 $Y=1.59
+ $X2=3.16 $Y2=1.59
r133 16 45 38.7914 $w=2.76e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.02 $Y=1.085
+ $X2=2.995 $Y2=1.25
r134 16 18 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.02 $Y=1.085
+ $X2=3.02 $Y2=0.445
r135 14 30 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.15 $Y=2.775
+ $X2=2.15 $Y2=2.295
r136 9 39 81.3502 $w=2.37e-07 $l=4.58258e-07 $layer=POLY_cond $X=2.11 $Y=0.73
+ $X2=1.985 $Y2=1.13
r137 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.11 $Y=0.73 $X2=2.11
+ $Y2=0.445
r138 2 42 600 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=2.075 $X2=1.395 $Y2=1.89
r139 1 36 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.68 $X2=1.21 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%A_45_136# 1 2 8 9 11 12 14 18 21 22 26 35 39
c84 26 0 2.32782e-19 $X=2.525 $Y=1.79
c85 22 0 6.42183e-20 $X=2.435 $Y=2.24
c86 18 0 1.12376e-19 $X=2.66 $Y=0.805
c87 14 0 1.34222e-19 $X=2.87 $Y=2.775
c88 12 0 1.53527e-19 $X=2.87 $Y=2.295
r89 39 41 9.67073 $w=4.1e-07 $l=3.25e-07 $layer=LI1_cond $X=0.32 $Y=2.24
+ $X2=0.32 $Y2=2.565
r90 38 39 0.446341 $w=4.1e-07 $l=1.5e-08 $layer=LI1_cond $X=0.32 $Y=2.225
+ $X2=0.32 $Y2=2.24
r91 32 35 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=0.195 $Y=0.87
+ $X2=0.35 $Y2=0.87
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=2.13 $X2=2.6 $Y2=2.13
r93 27 31 44.4119 $w=3.69e-07 $l=3.4e-07 $layer=POLY_cond $X=2.652 $Y=1.79
+ $X2=2.652 $Y2=2.13
r94 26 30 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=2.597 $Y=1.79
+ $X2=2.597 $Y2=2.13
r95 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.525
+ $Y=1.79 $X2=2.525 $Y2=1.79
r96 24 30 0.886495 $w=3.23e-07 $l=2.5e-08 $layer=LI1_cond $X=2.597 $Y=2.155
+ $X2=2.597 $Y2=2.13
r97 23 39 5.92876 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.53 $Y=2.24 $X2=0.32
+ $Y2=2.24
r98 22 24 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=2.435 $Y=2.24
+ $X2=2.597 $Y2=2.155
r99 22 23 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=2.435 $Y=2.24
+ $X2=0.53 $Y2=2.24
r100 21 38 9.20018 $w=4.1e-07 $l=2.18746e-07 $layer=LI1_cond $X=0.195 $Y=2.06
+ $X2=0.32 $Y2=2.225
r101 20 32 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.195 $Y=1.04
+ $X2=0.195 $Y2=0.87
r102 20 21 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.195 $Y=1.04
+ $X2=0.195 $Y2=2.06
r103 16 18 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.515 $Y=0.805
+ $X2=2.66 $Y2=0.805
r104 12 31 39.0404 $w=3.69e-07 $l=2.88953e-07 $layer=POLY_cond $X=2.87 $Y=2.295
+ $X2=2.652 $Y2=2.13
r105 12 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.87 $Y=2.295
+ $X2=2.87 $Y2=2.775
r106 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.66 $Y=0.73
+ $X2=2.66 $Y2=0.805
r107 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.66 $Y=0.73 $X2=2.66
+ $Y2=0.445
r108 8 27 39.0404 $w=3.69e-07 $l=2.23226e-07 $layer=POLY_cond $X=2.515 $Y=1.625
+ $X2=2.652 $Y2=1.79
r109 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.515 $Y=0.88
+ $X2=2.515 $Y2=0.805
r110 7 8 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.515 $Y=0.88
+ $X2=2.515 $Y2=1.625
r111 2 41 600 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=2.075 $X2=0.365 $Y2=2.565
r112 2 38 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=2.075 $X2=0.365 $Y2=2.225
r113 1 35 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.68 $X2=0.35 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%A_354_47# 1 2 9 13 19 21 22 23 26 27 28 31
+ 35 36 38
c115 31 0 2.323e-19 $X=3.32 $Y=2.13
c116 28 0 1.53889e-19 $X=3.1 $Y=2.092
r117 36 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.02
+ $X2=3.535 $Y2=0.855
r118 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.535
+ $Y=1.02 $X2=3.535 $Y2=1.02
r119 33 35 45.3774 $w=2.38e-07 $l=9.45e-07 $layer=LI1_cond $X=3.5 $Y=1.965
+ $X2=3.5 $Y2=1.02
r120 32 35 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=3.5 $Y=0.795
+ $X2=3.5 $Y2=1.02
r121 31 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.32 $Y=2.13
+ $X2=3.32 $Y2=2.295
r122 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=2.13 $X2=3.32 $Y2=2.13
r123 28 30 9.94265 $w=2.53e-07 $l=2.2e-07 $layer=LI1_cond $X=3.1 $Y=2.092
+ $X2=3.32 $Y2=2.092
r124 27 33 6.82464 $w=2.55e-07 $l=1.77113e-07 $layer=LI1_cond $X=3.38 $Y=2.092
+ $X2=3.5 $Y2=1.965
r125 27 30 2.71163 $w=2.53e-07 $l=6e-08 $layer=LI1_cond $X=3.38 $Y=2.092
+ $X2=3.32 $Y2=2.092
r126 25 28 7.17723 $w=2.55e-07 $l=1.65118e-07 $layer=LI1_cond $X=3.015 $Y=2.22
+ $X2=3.1 $Y2=2.092
r127 25 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.015 $Y=2.22
+ $X2=3.015 $Y2=2.495
r128 24 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=2.58
+ $X2=1.935 $Y2=2.58
r129 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.93 $Y=2.58
+ $X2=3.015 $Y2=2.495
r130 23 24 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.93 $Y=2.58
+ $X2=2.1 $Y2=2.58
r131 21 32 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.38 $Y=0.71
+ $X2=3.5 $Y2=0.795
r132 21 22 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.38 $Y=0.71
+ $X2=2.05 $Y2=0.71
r133 17 22 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.915 $Y=0.625
+ $X2=2.05 $Y2=0.71
r134 17 19 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.915 $Y=0.625
+ $X2=1.915 $Y2=0.445
r135 13 43 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.61 $Y=0.445
+ $X2=3.61 $Y2=0.855
r136 9 41 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.23 $Y=2.775
+ $X2=3.23 $Y2=2.295
r137 2 38 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=1.81
+ $Y=2.455 $X2=1.935 $Y2=2.61
r138 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.235 $X2=1.895 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%A_805_21# 1 2 9 14 18 20 24 26 28 33 35 37
+ 38 39 41 42 43 45 46 48 53 56 59 60 61 62 63 64 65 67 68 69 72 73 77 78 80 87
+ 90 93
r186 92 94 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=8.085 $Y=1.46
+ $X2=8.165 $Y2=1.46
r187 92 93 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.085 $Y=1.46
+ $X2=8.01 $Y2=1.46
r188 83 90 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.875 $Y=0.36
+ $X2=6.05 $Y2=0.36
r189 82 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.875
+ $Y=0.36 $X2=5.875 $Y2=0.36
r190 77 87 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.22 $Y=1.9
+ $X2=4.22 $Y2=2.065
r191 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=1.9 $X2=4.22 $Y2=1.9
r192 73 94 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=8.32 $Y=1.46
+ $X2=8.165 $Y2=1.46
r193 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.32
+ $Y=1.46 $X2=8.32 $Y2=1.46
r194 70 72 36.7477 $w=2.63e-07 $l=8.45e-07 $layer=LI1_cond $X=8.357 $Y=2.305
+ $X2=8.357 $Y2=1.46
r195 68 70 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=8.225 $Y=2.39
+ $X2=8.357 $Y2=2.305
r196 68 69 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=8.225 $Y=2.39
+ $X2=7.445 $Y2=2.39
r197 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.36 $Y=2.305
+ $X2=7.445 $Y2=2.39
r198 66 67 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=7.36 $Y=0.795
+ $X2=7.36 $Y2=2.305
r199 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.275 $Y=0.71
+ $X2=7.36 $Y2=0.795
r200 64 65 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=7.275 $Y=0.71
+ $X2=6.04 $Y2=0.71
r201 63 65 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.875 $Y=0.625
+ $X2=6.04 $Y2=0.71
r202 62 82 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=5.875 $Y=0.455
+ $X2=5.875 $Y2=0.355
r203 62 63 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.875 $Y=0.455
+ $X2=5.875 $Y2=0.625
r204 60 82 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=0.355
+ $X2=5.875 $Y2=0.355
r205 60 61 24.6773 $w=1.98e-07 $l=4.45e-07 $layer=LI1_cond $X=5.71 $Y=0.355
+ $X2=5.265 $Y2=0.355
r206 59 80 6.10429 $w=2.2e-07 $l=1.53704e-07 $layer=LI1_cond $X=5.175 $Y=1.795
+ $X2=5.135 $Y2=1.93
r207 59 78 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=5.175 $Y=1.795
+ $X2=5.175 $Y2=1.125
r208 54 80 6.10429 $w=2.2e-07 $l=1.35e-07 $layer=LI1_cond $X=5.135 $Y=2.065
+ $X2=5.135 $Y2=1.93
r209 54 56 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=5.135 $Y=2.065
+ $X2=5.135 $Y2=2.425
r210 51 78 9.60236 $w=4.18e-07 $l=2.1e-07 $layer=LI1_cond $X=5.055 $Y=0.915
+ $X2=5.055 $Y2=1.125
r211 51 53 12.2104 $w=4.18e-07 $l=4.45e-07 $layer=LI1_cond $X=5.055 $Y=0.915
+ $X2=5.055 $Y2=0.47
r212 50 61 7.99718 $w=2e-07 $l=2.55147e-07 $layer=LI1_cond $X=5.055 $Y=0.455
+ $X2=5.265 $Y2=0.355
r213 50 53 0.411587 $w=4.18e-07 $l=1.5e-08 $layer=LI1_cond $X=5.055 $Y=0.455
+ $X2=5.055 $Y2=0.47
r214 49 76 3.02242 $w=2.7e-07 $l=1.03e-07 $layer=LI1_cond $X=4.335 $Y=1.93
+ $X2=4.232 $Y2=1.93
r215 48 80 0.616579 $w=2.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.005 $Y=1.93
+ $X2=5.135 $Y2=1.93
r216 48 49 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.005 $Y=1.93
+ $X2=4.335 $Y2=1.93
r217 46 77 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.22 $Y=1.56
+ $X2=4.22 $Y2=1.9
r218 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=1.56 $X2=4.22 $Y2=1.56
r219 43 76 3.96142 $w=2.05e-07 $l=1.35e-07 $layer=LI1_cond $X=4.232 $Y=1.795
+ $X2=4.232 $Y2=1.93
r220 43 45 12.714 $w=2.03e-07 $l=2.35e-07 $layer=LI1_cond $X=4.232 $Y=1.795
+ $X2=4.232 $Y2=1.56
r221 41 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.22 $Y=1.395
+ $X2=4.22 $Y2=1.56
r222 39 41 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.13 $Y=0.915
+ $X2=4.13 $Y2=1.395
r223 38 39 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.115 $Y=0.765
+ $X2=4.115 $Y2=0.915
r224 35 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.165 $Y=1.295
+ $X2=8.165 $Y2=1.46
r225 35 37 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.165 $Y=1.295
+ $X2=8.165 $Y2=0.765
r226 31 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.085 $Y=1.625
+ $X2=8.085 $Y2=1.46
r227 31 33 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.085 $Y=1.625
+ $X2=8.085 $Y2=2.465
r228 30 42 5.30422 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=7.81 $Y=1.37
+ $X2=7.695 $Y2=1.37
r229 30 93 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.81 $Y=1.37 $X2=8.01
+ $Y2=1.37
r230 26 42 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=7.735 $Y=1.295
+ $X2=7.695 $Y2=1.37
r231 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.735 $Y=1.295
+ $X2=7.735 $Y2=0.765
r232 22 42 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=7.655 $Y=1.445
+ $X2=7.695 $Y2=1.37
r233 22 24 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=7.655 $Y=1.445
+ $X2=7.655 $Y2=2.465
r234 18 20 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=6.05 $Y=0.975
+ $X2=6.05 $Y2=2.155
r235 16 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=0.525
+ $X2=6.05 $Y2=0.36
r236 16 18 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.05 $Y=0.525
+ $X2=6.05 $Y2=0.975
r237 14 87 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.13 $Y=2.665 $X2=4.13
+ $Y2=2.065
r238 9 38 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.1 $Y=0.445 $X2=4.1
+ $Y2=0.765
r239 2 80 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=1.785 $X2=5.1 $Y2=1.93
r240 2 56 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=4.96
+ $Y=1.785 $X2=5.1 $Y2=2.425
r241 1 53 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.835
+ $Y=0.345 $X2=4.975 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%A_619_47# 1 2 9 12 14 20 24 25 27 29 30 32
+ 36 38
c93 25 0 1.34222e-19 $X=3.61 $Y=2.475
r94 36 39 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.777 $Y=1.46
+ $X2=4.777 $Y2=1.625
r95 36 38 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.777 $Y=1.46
+ $X2=4.777 $Y2=1.295
r96 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.76
+ $Y=1.46 $X2=4.76 $Y2=1.46
r97 31 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=1.14
+ $X2=3.875 $Y2=1.14
r98 30 35 12.6753 $w=3.08e-07 $l=4.09878e-07 $layer=LI1_cond $X=4.505 $Y=1.14
+ $X2=4.71 $Y2=1.46
r99 30 31 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.505 $Y=1.14
+ $X2=3.96 $Y2=1.14
r100 28 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=1.225
+ $X2=3.875 $Y2=1.14
r101 28 29 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=3.875 $Y=1.225
+ $X2=3.875 $Y2=2.39
r102 27 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=1.055
+ $X2=3.875 $Y2=1.14
r103 26 27 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.875 $Y=0.455
+ $X2=3.875 $Y2=1.055
r104 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.79 $Y=2.475
+ $X2=3.875 $Y2=2.39
r105 24 25 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.79 $Y=2.475
+ $X2=3.61 $Y2=2.475
r106 20 22 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.445 $Y=2.6
+ $X2=3.445 $Y2=2.94
r107 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.445 $Y=2.56
+ $X2=3.61 $Y2=2.475
r108 18 20 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=3.445 $Y=2.56
+ $X2=3.445 $Y2=2.6
r109 14 26 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.79 $Y=0.355
+ $X2=3.875 $Y2=0.455
r110 14 16 26.3409 $w=1.98e-07 $l=4.75e-07 $layer=LI1_cond $X=3.79 $Y=0.355
+ $X2=3.315 $Y2=0.355
r111 12 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.885 $Y=2.415
+ $X2=4.885 $Y2=1.625
r112 9 38 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.76 $Y=0.765
+ $X2=4.76 $Y2=1.295
r113 2 22 600 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=2.455 $X2=3.445 $Y2=2.94
r114 2 20 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=2.455 $X2=3.445 $Y2=2.6
r115 1 16 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.235 $X2=3.315 $Y2=0.35
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%A_1138_153# 1 2 7 9 12 14 16 18 21 23 26 30
+ 34 41
r64 40 41 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.715 $Y=1.46
+ $X2=6.79 $Y2=1.46
r65 36 37 5.91831 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=1.46
+ $X2=5.835 $Y2=1.625
r66 34 36 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.835 $Y=1.06 $X2=5.835
+ $Y2=1.46
r67 31 40 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.5 $Y=1.46
+ $X2=6.715 $Y2=1.46
r68 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.5
+ $Y=1.46 $X2=6.5 $Y2=1.46
r69 28 36 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=1.46 $X2=5.835
+ $Y2=1.46
r70 28 30 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6 $Y=1.46 $X2=6.5
+ $Y2=1.46
r71 26 37 13.8684 $w=2.93e-07 $l=3.55e-07 $layer=LI1_cond $X=5.817 $Y=1.98
+ $X2=5.817 $Y2=1.625
r72 19 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.145 $Y=1.445
+ $X2=7.145 $Y2=1.37
r73 19 21 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=7.145 $Y=1.445
+ $X2=7.145 $Y2=2.465
r74 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.145 $Y=1.295
+ $X2=7.145 $Y2=1.37
r75 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.145 $Y=1.295
+ $X2=7.145 $Y2=0.765
r76 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.07 $Y=1.37
+ $X2=7.145 $Y2=1.37
r77 14 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.07 $Y=1.37
+ $X2=6.79 $Y2=1.37
r78 10 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.625
+ $X2=6.715 $Y2=1.46
r79 10 12 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.715 $Y=1.625
+ $X2=6.715 $Y2=2.465
r80 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.295
+ $X2=6.715 $Y2=1.46
r81 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.715 $Y=1.295
+ $X2=6.715 $Y2=0.765
r82 2 26 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.71
+ $Y=1.835 $X2=5.835 $Y2=1.98
r83 1 34 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=5.69
+ $Y=0.765 $X2=5.835 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%VPWR 1 2 3 4 5 6 23 27 31 37 43 45 47 49 51
+ 59 64 72 77 83 86 89 92 95 99
r107 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r108 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r109 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r111 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 81 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r114 81 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r116 78 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.43 $Y2=3.33
r117 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 77 98 4.61575 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=8.135 $Y=3.33
+ $X2=8.387 $Y2=3.33
r119 77 80 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.135 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 76 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r121 76 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 73 92 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.36 $Y2=3.33
r124 73 75 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 72 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.43 $Y2=3.33
r126 72 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=6.96 $Y2=3.33
r127 71 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r128 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r129 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r130 68 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 67 70 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r132 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 65 89 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.835 $Y=3.33
+ $X2=4.54 $Y2=3.33
r134 65 67 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.835 $Y=3.33
+ $X2=5.04 $Y2=3.33
r135 64 92 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.36 $Y2=3.33
r136 64 70 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6 $Y2=3.33
r137 63 87 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r139 60 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.505 $Y2=3.33
r140 60 62 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=4.08 $Y2=3.33
r141 59 89 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.54 $Y2=3.33
r142 59 62 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 58 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r144 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r146 55 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 54 57 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r148 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r149 52 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.85 $Y2=3.33
r150 52 54 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.2 $Y2=3.33
r151 51 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.505 $Y2=3.33
r152 51 57 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.16 $Y2=3.33
r153 49 90 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 49 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r155 45 98 3.15043 $w=3.3e-07 $l=1.22327e-07 $layer=LI1_cond $X=8.3 $Y=3.245
+ $X2=8.387 $Y2=3.33
r156 45 47 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=8.3 $Y=3.245
+ $X2=8.3 $Y2=2.77
r157 41 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=3.245
+ $X2=7.43 $Y2=3.33
r158 41 43 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=7.43 $Y=3.245
+ $X2=7.43 $Y2=2.77
r159 37 40 17.8083 $w=4.48e-07 $l=6.7e-07 $layer=LI1_cond $X=6.36 $Y=1.96
+ $X2=6.36 $Y2=2.63
r160 35 92 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.36 $Y=3.245
+ $X2=6.36 $Y2=3.33
r161 35 40 16.3464 $w=4.48e-07 $l=6.15e-07 $layer=LI1_cond $X=6.36 $Y=3.245
+ $X2=6.36 $Y2=2.63
r162 31 34 12.1635 $w=5.88e-07 $l=6e-07 $layer=LI1_cond $X=4.54 $Y=2.32 $X2=4.54
+ $Y2=2.92
r163 29 89 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=3.245
+ $X2=4.54 $Y2=3.33
r164 29 34 6.58857 $w=5.88e-07 $l=3.25e-07 $layer=LI1_cond $X=4.54 $Y=3.245
+ $X2=4.54 $Y2=2.92
r165 25 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=3.245
+ $X2=2.505 $Y2=3.33
r166 25 27 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.505 $Y=3.245
+ $X2=2.505 $Y2=2.945
r167 21 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=3.33
r168 21 23 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=2.59
r169 6 47 600 $w=1.7e-07 $l=1.00256e-06 $layer=licon1_PDIFF $count=1 $X=8.16
+ $Y=1.835 $X2=8.3 $Y2=2.77
r170 5 43 600 $w=1.7e-07 $l=1.03469e-06 $layer=licon1_PDIFF $count=1 $X=7.22
+ $Y=1.835 $X2=7.43 $Y2=2.77
r171 4 40 300 $w=1.7e-07 $l=9.64443e-07 $layer=licon1_PDIFF $count=2 $X=6.125
+ $Y=1.835 $X2=6.5 $Y2=2.63
r172 4 37 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.125
+ $Y=1.835 $X2=6.265 $Y2=1.96
r173 3 34 400 $w=1.7e-07 $l=6.57609e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=2.455 $X2=4.67 $Y2=2.92
r174 3 31 400 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=2.455 $X2=4.67 $Y2=2.32
r175 2 27 600 $w=1.7e-07 $l=6.14247e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=2.455 $X2=2.505 $Y2=2.945
r176 1 23 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=2.075 $X2=0.85 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%Q_N 1 2 7 8 9 10 11 18
r17 11 32 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.93 $Y=2.775
+ $X2=6.93 $Y2=2.91
r18 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.93 $Y=2.405
+ $X2=6.93 $Y2=2.775
r19 9 10 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.93 $Y=2.015
+ $X2=6.93 $Y2=2.405
r20 8 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.93 $Y=1.665 $X2=6.93
+ $Y2=2.015
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.93 $Y=1.295 $X2=6.93
+ $Y2=1.665
r22 7 18 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=6.93 $Y=1.295
+ $X2=6.93 $Y2=1.06
r23 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.79
+ $Y=1.835 $X2=6.93 $Y2=2.91
r24 2 9 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=6.79 $Y=1.835
+ $X2=6.93 $Y2=2.015
r25 1 18 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=6.79
+ $Y=0.345 $X2=6.93 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%Q 1 2 8 10 11 12 13 14
r26 13 14 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=7.875 $Y=1.665
+ $X2=7.875 $Y2=2.01
r27 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=7.875 $Y=1.295
+ $X2=7.875 $Y2=1.665
r28 11 12 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=7.875 $Y=0.925
+ $X2=7.875 $Y2=1.295
r29 9 10 6.82929 $w=2.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.91 $Y=0.655
+ $X2=7.91 $Y2=0.495
r30 8 11 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=7.875 $Y=0.825
+ $X2=7.875 $Y2=0.925
r31 8 9 6.28338 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=7.875 $Y=0.825
+ $X2=7.875 $Y2=0.655
r32 2 14 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.835 $X2=7.87 $Y2=2.01
r33 1 10 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=7.81
+ $Y=0.345 $X2=7.95 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_2%VGND 1 2 3 4 5 6 23 27 31 35 39 41 43 46 47
+ 49 50 51 60 71 75 81 84 87 91
c112 60 0 1.12376e-19 $X=4.265 $Y=0
r113 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r114 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r115 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r116 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 79 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r118 79 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r119 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r120 76 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=0 $X2=7.44
+ $Y2=0
r121 76 78 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.605 $Y=0
+ $X2=7.92 $Y2=0
r122 75 90 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=8.215 $Y=0
+ $X2=8.427 $Y2=0
r123 75 78 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.215 $Y=0 $X2=7.92
+ $Y2=0
r124 74 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r125 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r126 71 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.275 $Y=0 $X2=7.44
+ $Y2=0
r127 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=6.96 $Y2=0
r128 70 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r129 70 85 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.56
+ $Y2=0
r130 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r131 67 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.43
+ $Y2=0
r132 67 69 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=4.595 $Y=0 $X2=6
+ $Y2=0
r133 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r134 63 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.08 $Y2=0
r135 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r136 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r137 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.43
+ $Y2=0
r138 60 65 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.265 $Y=0
+ $X2=4.08 $Y2=0
r139 59 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r140 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r141 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r142 56 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r143 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r144 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r145 53 81 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.765
+ $Y2=0
r146 53 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r147 51 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r148 51 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r149 49 69 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.22 $Y=0 $X2=6
+ $Y2=0
r150 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.22 $Y=0 $X2=6.385
+ $Y2=0
r151 48 73 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.96
+ $Y2=0
r152 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.385
+ $Y2=0
r153 46 58 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.16
+ $Y2=0
r154 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.385
+ $Y2=0
r155 45 62 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.64
+ $Y2=0
r156 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.385
+ $Y2=0
r157 41 90 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=8.38 $Y=0.085
+ $X2=8.427 $Y2=0
r158 41 43 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=8.38 $Y=0.085
+ $X2=8.38 $Y2=0.49
r159 37 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0
r160 37 39 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0.36
r161 33 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=0.085
+ $X2=6.385 $Y2=0
r162 33 35 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.385 $Y=0.085
+ $X2=6.385 $Y2=0.36
r163 29 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.43 $Y=0.085
+ $X2=4.43 $Y2=0
r164 29 31 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.43 $Y=0.085
+ $X2=4.43 $Y2=0.36
r165 25 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0
r166 25 27 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0.35
r167 21 81 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0
r168 21 23 41.3832 $w=2.18e-07 $l=7.9e-07 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0.875
r169 6 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.24
+ $Y=0.345 $X2=8.38 $Y2=0.49
r170 5 39 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=7.22
+ $Y=0.345 $X2=7.44 $Y2=0.36
r171 4 35 182 $w=1.7e-07 $l=5.18965e-07 $layer=licon1_NDIFF $count=1 $X=6.125
+ $Y=0.765 $X2=6.385 $Y2=0.36
r172 3 31 91 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=2 $X=4.175
+ $Y=0.235 $X2=4.43 $Y2=0.36
r173 2 27 182 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_NDIFF $count=1 $X=2.185
+ $Y=0.235 $X2=2.385 $Y2=0.35
r174 1 23 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.68 $X2=0.78 $Y2=0.875
.ends

