* File: sky130_fd_sc_lp__nor3b_lp.spice
* Created: Wed Sep  2 10:09:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor3b_lp.pex.spice"
.subckt sky130_fd_sc_lp__nor3b_lp  VNB VPB A B C_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C_N	C_N
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_136_57# N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.9
+ A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g A_136_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1002 A_294_57# N_B_M1002_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75002.1 A=0.063
+ P=1.14 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g A_294_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1007 A_452_57# N_A_350_269#_M1007_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_350_269#_M1005_g A_452_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_610_57# N_C_N_M1008_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_350_269#_M1009_d N_C_N_M1009_g A_610_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 A_188_409# N_A_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1003 A_286_409# N_B_M1003_g A_188_409# VPB PHIGHVT L=0.25 W=1 AD=0.16 AS=0.12
+ PD=1.32 PS=1.24 NRD=20.6653 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1000 N_Y_M1000_d N_A_350_269#_M1000_g A_286_409# VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=20.6653 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1006 N_A_350_269#_M1006_d N_C_N_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__nor3b_lp.pxi.spice"
*
.ends
*
*
