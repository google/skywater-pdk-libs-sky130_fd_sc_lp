* NGSPICE file created from sky130_fd_sc_lp__o22ai_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o22ai_m A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A2 a_85_82# VNB nshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=4.074e+11p ps=4.46e+06u
M1001 a_198_535# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.226e+11p ps=2.74e+06u
M1002 Y B2 a_198_535# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1003 a_85_82# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 a_85_82# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1005 VPWR A1 a_356_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_85_82# B2 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_356_535# A2 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

