* File: sky130_fd_sc_lp__nor2b_4.pxi.spice
* Created: Fri Aug 28 10:54:42 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2B_4%B_N N_B_N_M1012_g N_B_N_M1013_g N_B_N_c_85_n
+ N_B_N_c_86_n B_N N_B_N_c_87_n PM_SKY130_FD_SC_LP__NOR2B_4%B_N
x_PM_SKY130_FD_SC_LP__NOR2B_4%A N_A_M1001_g N_A_M1000_g N_A_M1002_g N_A_M1005_g
+ N_A_M1009_g N_A_M1014_g N_A_M1016_g N_A_M1015_g N_A_c_115_n N_A_c_116_n
+ N_A_c_128_n N_A_c_117_n N_A_c_130_n A A A N_A_c_119_n N_A_c_120_n N_A_c_121_n
+ N_A_c_133_n PM_SKY130_FD_SC_LP__NOR2B_4%A
x_PM_SKY130_FD_SC_LP__NOR2B_4%A_60_47# N_A_60_47#_M1012_s N_A_60_47#_M1013_s
+ N_A_60_47#_c_269_n N_A_60_47#_M1004_g N_A_60_47#_M1003_g N_A_60_47#_c_271_n
+ N_A_60_47#_M1006_g N_A_60_47#_M1007_g N_A_60_47#_c_273_n N_A_60_47#_M1010_g
+ N_A_60_47#_M1008_g N_A_60_47#_c_275_n N_A_60_47#_M1017_g N_A_60_47#_M1011_g
+ N_A_60_47#_c_277_n N_A_60_47#_c_290_n N_A_60_47#_c_278_n N_A_60_47#_c_279_n
+ N_A_60_47#_c_280_n N_A_60_47#_c_281_n N_A_60_47#_c_292_n N_A_60_47#_c_282_n
+ N_A_60_47#_c_283_n N_A_60_47#_c_284_n N_A_60_47#_c_285_n
+ PM_SKY130_FD_SC_LP__NOR2B_4%A_60_47#
x_PM_SKY130_FD_SC_LP__NOR2B_4%VPWR N_VPWR_M1013_d N_VPWR_M1005_s N_VPWR_M1015_s
+ N_VPWR_c_430_n N_VPWR_c_444_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_450_n
+ N_VPWR_c_433_n N_VPWR_c_434_n VPWR N_VPWR_c_435_n N_VPWR_c_429_n
+ PM_SKY130_FD_SC_LP__NOR2B_4%VPWR
x_PM_SKY130_FD_SC_LP__NOR2B_4%A_245_367# N_A_245_367#_M1000_d
+ N_A_245_367#_M1007_d N_A_245_367#_M1014_d N_A_245_367#_M1011_d
+ N_A_245_367#_c_508_n N_A_245_367#_c_534_p N_A_245_367#_c_513_n
+ N_A_245_367#_c_537_p N_A_245_367#_c_527_n
+ PM_SKY130_FD_SC_LP__NOR2B_4%A_245_367#
x_PM_SKY130_FD_SC_LP__NOR2B_4%Y N_Y_M1001_s N_Y_M1006_d N_Y_M1009_s N_Y_M1017_d
+ N_Y_M1003_s N_Y_M1008_s N_Y_c_545_n N_Y_c_578_n N_Y_c_546_n N_Y_c_547_n
+ N_Y_c_551_n N_Y_c_553_n N_Y_c_555_n N_Y_c_593_n N_Y_c_622_n N_Y_c_642_p
+ N_Y_c_538_n N_Y_c_561_n N_Y_c_564_n N_Y_c_565_n N_Y_c_566_n N_Y_c_539_n Y Y Y
+ PM_SKY130_FD_SC_LP__NOR2B_4%Y
x_PM_SKY130_FD_SC_LP__NOR2B_4%VGND N_VGND_M1012_d N_VGND_M1004_s N_VGND_M1002_d
+ N_VGND_M1010_s N_VGND_M1016_d N_VGND_c_655_n N_VGND_c_656_n N_VGND_c_657_n
+ N_VGND_c_658_n N_VGND_c_659_n N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n
+ N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n VGND N_VGND_c_666_n
+ N_VGND_c_667_n N_VGND_c_668_n N_VGND_c_669_n PM_SKY130_FD_SC_LP__NOR2B_4%VGND
cc_1 VNB N_B_N_M1012_g 0.0289544f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_2 VNB N_B_N_M1013_g 0.00144514f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_3 VNB N_B_N_c_85_n 0.0618704f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.46
cc_4 VNB N_B_N_c_86_n 0.0094345f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.46
cc_5 VNB N_B_N_c_87_n 0.0013005f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_6 VNB N_A_M1001_g 0.0245055f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_7 VNB N_A_M1002_g 0.0231699f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_M1009_g 0.0231684f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_9 VNB N_A_M1016_g 0.028067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_c_115_n 0.00100953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_116_n 0.0284749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_c_117_n 0.0258606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A 0.00429219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_c_119_n 0.0307246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_120_n 0.00110194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_c_121_n 0.0018677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_60_47#_c_269_n 0.0154474f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_18 VNB N_A_60_47#_M1003_g 0.00688781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_60_47#_c_271_n 0.0154648f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_20 VNB N_A_60_47#_M1007_g 0.00649604f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_21 VNB N_A_60_47#_c_273_n 0.015451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_60_47#_M1008_g 0.00725423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_60_47#_c_275_n 0.0161411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_60_47#_M1011_g 0.00705913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_60_47#_c_277_n 0.0284746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_60_47#_c_278_n 0.00312582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_60_47#_c_279_n 0.0169982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_60_47#_c_280_n 0.00987776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_60_47#_c_281_n 0.0159407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_60_47#_c_282_n 0.00336158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_60_47#_c_283_n 0.0041807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_60_47#_c_284_n 0.0371712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_60_47#_c_285_n 0.0383868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_429_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_538_n 0.0204402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_539_n 0.00384819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB Y 0.0244346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_655_n 0.002833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_656_n 0.00422004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_657_n 0.0167176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_658_n 0.003699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_659_n 0.00178362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_660_n 0.0156289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_661_n 0.0261041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_662_n 0.0176482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_663_n 0.00362148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_664_n 0.0167176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_665_n 0.00375786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_666_n 0.0124089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_667_n 0.0257608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_668_n 0.00362148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_669_n 0.261468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_B_N_M1013_g 0.0252636f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.465
cc_54 VPB N_B_N_c_87_n 0.0120687f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_55 VPB N_A_M1000_g 0.0183582f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.465
cc_56 VPB N_A_M1005_g 0.0174407f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_57 VPB N_A_M1014_g 0.0174407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_M1015_g 0.0216056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_c_115_n 3.78445e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_c_116_n 0.00657527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_c_128_n 0.00152935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_c_117_n 0.00648788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_c_130_n 0.00860397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB A 4.27982e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_c_119_n 0.00462236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_c_133_n 0.00557666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_60_47#_M1003_g 0.0186604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_60_47#_M1007_g 0.0185055f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.665
cc_69 VPB N_A_60_47#_M1008_g 0.0186928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_60_47#_M1011_g 0.018667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_60_47#_c_290_n 0.0372327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_60_47#_c_278_n 0.00116368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_60_47#_c_292_n 0.00724748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_430_n 0.00528682f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_75 VPB N_VPWR_c_431_n 0.015603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_432_n 0.0308394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_433_n 0.0234885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_434_n 0.00535984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_435_n 0.0731845f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_429_n 0.0580147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB Y 0.0174827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB Y 0.0150631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 N_B_N_M1012_g N_A_M1001_g 0.026222f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_84 N_B_N_M1013_g N_A_M1000_g 0.035239f $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_85 N_B_N_M1013_g N_A_c_128_n 6.09633e-19 $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_N_c_86_n N_A_c_128_n 2.77268e-19 $X=0.64 $Y=1.46 $X2=0 $Y2=0
cc_87 N_B_N_c_86_n N_A_c_117_n 0.0165311f $X=0.64 $Y=1.46 $X2=0 $Y2=0
cc_88 N_B_N_M1012_g N_A_60_47#_c_278_n 0.0020275f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_89 N_B_N_M1013_g N_A_60_47#_c_278_n 0.0123206f $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_90 N_B_N_c_86_n N_A_60_47#_c_278_n 0.0107096f $X=0.64 $Y=1.46 $X2=0 $Y2=0
cc_91 N_B_N_c_87_n N_A_60_47#_c_278_n 0.028833f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_92 N_B_N_M1012_g N_A_60_47#_c_280_n 0.0202943f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_93 N_B_N_c_85_n N_A_60_47#_c_280_n 0.0101056f $X=0.565 $Y=1.46 $X2=0 $Y2=0
cc_94 N_B_N_c_87_n N_A_60_47#_c_280_n 0.0149787f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_95 N_B_N_M1013_g N_A_60_47#_c_292_n 0.0126358f $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_96 N_B_N_c_85_n N_A_60_47#_c_292_n 0.00426347f $X=0.565 $Y=1.46 $X2=0 $Y2=0
cc_97 N_B_N_c_87_n N_A_60_47#_c_292_n 0.0139366f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_98 N_B_N_M1013_g N_VPWR_c_430_n 0.00758344f $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_99 N_B_N_M1013_g N_VPWR_c_433_n 0.00585385f $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B_N_M1013_g N_VPWR_c_429_n 0.0119758f $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B_N_M1012_g N_VGND_c_655_n 0.0119707f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_102 N_B_N_M1012_g N_VGND_c_667_n 0.00486043f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_103 N_B_N_M1012_g N_VGND_c_669_n 0.00930295f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_104 N_A_M1001_g N_A_60_47#_c_269_n 0.0228177f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_105 N_A_M1000_g N_A_60_47#_M1003_g 0.0565185f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_c_128_n N_A_60_47#_M1003_g 6.13968e-19 $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_107 N_A_c_121_n N_A_60_47#_M1003_g 8.56965e-19 $X=2.285 $Y=1.645 $X2=0 $Y2=0
cc_108 N_A_c_133_n N_A_60_47#_M1003_g 0.0121214f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_109 N_A_M1002_g N_A_60_47#_c_271_n 0.0321878f $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_110 N_A_M1005_g N_A_60_47#_M1007_g 0.0321878f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_c_121_n N_A_60_47#_M1007_g 0.00815428f $X=2.285 $Y=1.645 $X2=0 $Y2=0
cc_112 N_A_c_133_n N_A_60_47#_M1007_g 0.00874416f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_113 N_A_M1009_g N_A_60_47#_c_273_n 0.0255219f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_114 N_A_M1014_g N_A_60_47#_M1008_g 0.0255219f $X=2.87 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_c_130_n N_A_60_47#_M1008_g 0.0118551f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_116 N_A_M1016_g N_A_60_47#_c_275_n 0.0228151f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_117 N_A_M1015_g N_A_60_47#_M1011_g 0.0372564f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_c_115_n N_A_60_47#_M1011_g 3.95394e-19 $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_119 N_A_c_130_n N_A_60_47#_M1011_g 0.0150272f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_120 N_A_M1001_g N_A_60_47#_c_278_n 0.00165347f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A_M1000_g N_A_60_47#_c_278_n 0.00170593f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_c_128_n N_A_60_47#_c_278_n 0.0323762f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_123 N_A_c_117_n N_A_60_47#_c_278_n 0.00310735f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_124 N_A_M1001_g N_A_60_47#_c_279_n 0.0146378f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_125 N_A_c_128_n N_A_60_47#_c_279_n 0.0247643f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_126 N_A_c_117_n N_A_60_47#_c_279_n 0.00446668f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_127 N_A_c_133_n N_A_60_47#_c_279_n 0.0100815f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_128 N_A_M1001_g N_A_60_47#_c_280_n 0.0018506f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_129 N_A_M1002_g N_A_60_47#_c_281_n 0.010445f $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A_M1009_g N_A_60_47#_c_281_n 0.010445f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_131 N_A_c_130_n N_A_60_47#_c_281_n 0.00547072f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_132 N_A_c_119_n N_A_60_47#_c_281_n 0.00246472f $X=2.87 $Y=1.51 $X2=0 $Y2=0
cc_133 N_A_c_121_n N_A_60_47#_c_281_n 0.0886373f $X=2.285 $Y=1.645 $X2=0 $Y2=0
cc_134 N_A_c_133_n N_A_60_47#_c_281_n 0.00547454f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_135 N_A_M1000_g N_A_60_47#_c_292_n 0.00388625f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_M1001_g N_A_60_47#_c_282_n 5.92537e-19 $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_137 N_A_M1002_g N_A_60_47#_c_282_n 8.26584e-19 $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_138 N_A_c_128_n N_A_60_47#_c_282_n 0.00466679f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_139 N_A_c_117_n N_A_60_47#_c_282_n 7.81434e-19 $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_140 N_A_c_121_n N_A_60_47#_c_282_n 0.0071044f $X=2.285 $Y=1.645 $X2=0 $Y2=0
cc_141 N_A_c_133_n N_A_60_47#_c_282_n 0.0238747f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_142 N_A_M1009_g N_A_60_47#_c_283_n 8.91486e-19 $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_143 N_A_M1016_g N_A_60_47#_c_283_n 7.18948e-19 $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_144 N_A_c_115_n N_A_60_47#_c_283_n 0.00604552f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A_c_116_n N_A_60_47#_c_283_n 4.84402e-19 $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_146 N_A_c_130_n N_A_60_47#_c_283_n 0.0190444f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_147 A N_A_60_47#_c_283_n 0.00738405f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A_c_128_n N_A_60_47#_c_284_n 0.00142755f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A_c_117_n N_A_60_47#_c_284_n 0.0217612f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A_c_119_n N_A_60_47#_c_284_n 0.0321878f $X=2.87 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A_c_121_n N_A_60_47#_c_284_n 0.00280374f $X=2.285 $Y=1.645 $X2=0 $Y2=0
cc_152 N_A_c_133_n N_A_60_47#_c_284_n 6.96228e-19 $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_153 N_A_c_115_n N_A_60_47#_c_285_n 0.00180178f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A_c_116_n N_A_60_47#_c_285_n 0.0184358f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A_c_130_n N_A_60_47#_c_285_n 6.96228e-19 $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_156 A N_A_60_47#_c_285_n 0.00686345f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_c_119_n N_A_60_47#_c_285_n 0.0255219f $X=2.87 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A_c_128_n N_VPWR_M1013_d 0.00113435f $X=1.13 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_c_120_n N_VPWR_M1005_s 0.00182141f $X=2.985 $Y=1.645 $X2=0 $Y2=0
cc_160 N_A_c_130_n N_VPWR_M1015_s 4.64841e-19 $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_161 N_A_M1000_g N_VPWR_c_430_n 0.00356843f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_M1000_g N_VPWR_c_444_n 0.0135463f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_M1005_g N_VPWR_c_444_n 0.0102746f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A_M1014_g N_VPWR_c_444_n 0.00302552f $X=2.87 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_c_128_n N_VPWR_c_444_n 0.00446839f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A_c_133_n N_VPWR_c_444_n 0.00793549f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_167 N_A_M1015_g N_VPWR_c_432_n 0.0154314f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_M1000_g N_VPWR_c_450_n 0.00438118f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_c_128_n N_VPWR_c_450_n 0.00252065f $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A_c_117_n N_VPWR_c_450_n 3.75316e-19 $X=1.13 $Y=1.51 $X2=0 $Y2=0
cc_171 N_A_M1000_g N_VPWR_c_435_n 0.004201f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_M1005_g N_VPWR_c_435_n 0.00359964f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A_M1014_g N_VPWR_c_435_n 0.00359964f $X=2.87 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_M1015_g N_VPWR_c_435_n 0.00486043f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_M1000_g N_VPWR_c_429_n 0.00588888f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_M1005_g N_VPWR_c_429_n 0.00537821f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A_M1014_g N_VPWR_c_429_n 0.00537821f $X=2.87 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_M1015_g N_VPWR_c_429_n 0.0082726f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A_c_128_n N_A_245_367#_M1000_d 3.08849e-19 $X=1.13 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_c_133_n N_A_245_367#_M1000_d 0.00300445f $X=2.065 $Y=1.645 $X2=-0.19
+ $Y2=-0.245
cc_181 N_A_c_120_n N_A_245_367#_M1007_d 2.41392e-19 $X=2.985 $Y=1.645 $X2=0
+ $Y2=0
cc_182 N_A_c_121_n N_A_245_367#_M1007_d 0.00156905f $X=2.285 $Y=1.645 $X2=0
+ $Y2=0
cc_183 A N_A_245_367#_M1014_d 0.00182141f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A_c_130_n N_A_245_367#_M1011_d 0.00176891f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_185 N_A_M1000_g N_A_245_367#_c_508_n 0.00299722f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_M1005_g N_A_245_367#_c_508_n 0.00958686f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_M1014_g N_A_245_367#_c_508_n 0.0113783f $X=2.87 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_c_133_n N_Y_M1003_s 0.00176891f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_189 N_A_c_130_n N_Y_M1008_s 0.00176461f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_190 N_A_M1001_g N_Y_c_545_n 0.00531616f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A_M1001_g N_Y_c_546_n 0.00296375f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_M1005_g N_Y_c_547_n 0.010745f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_M1014_g N_Y_c_547_n 0.0122549f $X=2.87 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_c_119_n N_Y_c_547_n 4.50113e-19 $X=2.87 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A_c_120_n N_Y_c_547_n 0.0475739f $X=2.985 $Y=1.645 $X2=0 $Y2=0
cc_196 N_A_M1002_g N_Y_c_551_n 0.00637926f $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_197 N_A_M1009_g N_Y_c_551_n 5.25381e-19 $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_198 N_A_M1002_g N_Y_c_553_n 0.00886808f $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_199 N_A_M1009_g N_Y_c_553_n 0.00886808f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A_M1002_g N_Y_c_555_n 5.25381e-19 $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_M1009_g N_Y_c_555_n 0.00637926f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_202 N_A_M1016_g N_Y_c_538_n 0.0144627f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_203 N_A_c_115_n N_Y_c_538_n 0.0196225f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_204 N_A_c_116_n N_Y_c_538_n 0.00342855f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_205 N_A_c_130_n N_Y_c_538_n 5.03485e-19 $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_206 N_A_M1000_g N_Y_c_561_n 0.00105603f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_M1005_g N_Y_c_561_n 2.39364e-19 $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_c_133_n N_Y_c_561_n 0.0475739f $X=2.065 $Y=1.645 $X2=0 $Y2=0
cc_209 N_A_M1002_g N_Y_c_564_n 7.17169e-19 $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A_M1009_g N_Y_c_565_n 7.17169e-19 $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_211 N_A_c_130_n N_Y_c_566_n 0.0135055f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_212 N_A_c_130_n N_Y_c_539_n 0.00728863f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_213 N_A_M1016_g Y 0.00554833f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A_M1015_g Y 0.00672111f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_c_115_n Y 0.026444f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A_c_116_n Y 0.00809258f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_217 N_A_c_130_n Y 0.014541f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_218 N_A_M1015_g Y 0.0160093f $X=4.16 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A_c_116_n Y 0.00239032f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_220 N_A_c_130_n Y 0.0344005f $X=4.045 $Y=1.78 $X2=0 $Y2=0
cc_221 N_A_M1001_g N_VGND_c_655_n 0.00615664f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A_M1002_g N_VGND_c_657_n 0.00428252f $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_223 N_A_M1002_g N_VGND_c_658_n 0.00153274f $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_224 N_A_M1009_g N_VGND_c_658_n 0.00153274f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_225 N_A_M1016_g N_VGND_c_659_n 5.35628e-19 $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_226 N_A_M1016_g N_VGND_c_661_n 0.0113738f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_227 N_A_M1001_g N_VGND_c_662_n 0.0054895f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_228 N_A_M1009_g N_VGND_c_664_n 0.00428252f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_229 N_A_M1016_g N_VGND_c_666_n 0.00486043f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_230 N_A_M1001_g N_VGND_c_669_n 0.0101477f $X=1.15 $Y=0.655 $X2=0 $Y2=0
cc_231 N_A_M1002_g N_VGND_c_669_n 0.00587209f $X=2.44 $Y=0.655 $X2=0 $Y2=0
cc_232 N_A_M1009_g N_VGND_c_669_n 0.00587209f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_233 N_A_M1016_g N_VGND_c_669_n 0.0082726f $X=4.16 $Y=0.655 $X2=0 $Y2=0
cc_234 N_A_60_47#_c_278_n N_VPWR_M1013_d 0.00112373f $X=0.7 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_60_47#_c_292_n N_VPWR_M1013_d 0.00261557f $X=0.7 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_60_47#_M1003_g N_VPWR_c_444_n 0.0143483f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_60_47#_M1007_g N_VPWR_c_444_n 0.0129984f $X=2.01 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_60_47#_M1011_g N_VPWR_c_432_n 0.00111968f $X=3.73 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A_60_47#_M1003_g N_VPWR_c_450_n 8.31629e-19 $X=1.58 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A_60_47#_c_292_n N_VPWR_c_450_n 0.00102118f $X=0.7 $Y=2.015 $X2=0 $Y2=0
cc_241 N_A_60_47#_c_290_n N_VPWR_c_433_n 0.0181659f $X=0.425 $Y=2.91 $X2=0 $Y2=0
cc_242 N_A_60_47#_M1003_g N_VPWR_c_435_n 0.00359964f $X=1.58 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_A_60_47#_M1007_g N_VPWR_c_435_n 0.00359964f $X=2.01 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_A_60_47#_M1008_g N_VPWR_c_435_n 0.00359964f $X=3.3 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A_60_47#_M1011_g N_VPWR_c_435_n 0.00359964f $X=3.73 $Y=2.465 $X2=0
+ $Y2=0
cc_246 N_A_60_47#_M1013_s N_VPWR_c_429_n 0.00336915f $X=0.3 $Y=1.835 $X2=0 $Y2=0
cc_247 N_A_60_47#_M1003_g N_VPWR_c_429_n 0.00537821f $X=1.58 $Y=2.465 $X2=0
+ $Y2=0
cc_248 N_A_60_47#_M1007_g N_VPWR_c_429_n 0.00537821f $X=2.01 $Y=2.465 $X2=0
+ $Y2=0
cc_249 N_A_60_47#_M1008_g N_VPWR_c_429_n 0.00537821f $X=3.3 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A_60_47#_M1011_g N_VPWR_c_429_n 0.00537821f $X=3.73 $Y=2.465 $X2=0
+ $Y2=0
cc_251 N_A_60_47#_c_290_n N_VPWR_c_429_n 0.0104192f $X=0.425 $Y=2.91 $X2=0 $Y2=0
cc_252 N_A_60_47#_M1003_g N_A_245_367#_c_508_n 0.00960322f $X=1.58 $Y=2.465
+ $X2=0 $Y2=0
cc_253 N_A_60_47#_M1007_g N_A_245_367#_c_508_n 0.00960322f $X=2.01 $Y=2.465
+ $X2=0 $Y2=0
cc_254 N_A_60_47#_M1008_g N_A_245_367#_c_513_n 0.012559f $X=3.3 $Y=2.465 $X2=0
+ $Y2=0
cc_255 N_A_60_47#_M1011_g N_A_245_367#_c_513_n 0.0126083f $X=3.73 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_A_60_47#_c_269_n N_Y_c_545_n 0.00637926f $X=1.58 $Y=1.185 $X2=0 $Y2=0
cc_257 N_A_60_47#_c_271_n N_Y_c_545_n 5.25381e-19 $X=2.01 $Y=1.185 $X2=0 $Y2=0
cc_258 N_A_60_47#_c_269_n N_Y_c_578_n 0.00885073f $X=1.58 $Y=1.185 $X2=0 $Y2=0
cc_259 N_A_60_47#_c_271_n N_Y_c_578_n 0.00886808f $X=2.01 $Y=1.185 $X2=0 $Y2=0
cc_260 N_A_60_47#_c_279_n N_Y_c_578_n 0.00233842f $X=1.565 $Y=1.17 $X2=0 $Y2=0
cc_261 N_A_60_47#_c_281_n N_Y_c_578_n 0.00994467f $X=3.375 $Y=1.17 $X2=0 $Y2=0
cc_262 N_A_60_47#_c_282_n N_Y_c_578_n 0.0229896f $X=1.73 $Y=1.17 $X2=0 $Y2=0
cc_263 N_A_60_47#_c_284_n N_Y_c_578_n 5.4431e-19 $X=2.01 $Y=1.35 $X2=0 $Y2=0
cc_264 N_A_60_47#_c_269_n N_Y_c_546_n 7.17169e-19 $X=1.58 $Y=1.185 $X2=0 $Y2=0
cc_265 N_A_60_47#_c_279_n N_Y_c_546_n 0.0217194f $X=1.565 $Y=1.17 $X2=0 $Y2=0
cc_266 N_A_60_47#_M1007_g N_Y_c_547_n 0.00756348f $X=2.01 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A_60_47#_M1008_g N_Y_c_547_n 0.0129469f $X=3.3 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A_60_47#_c_269_n N_Y_c_551_n 5.25381e-19 $X=1.58 $Y=1.185 $X2=0 $Y2=0
cc_269 N_A_60_47#_c_271_n N_Y_c_551_n 0.00637926f $X=2.01 $Y=1.185 $X2=0 $Y2=0
cc_270 N_A_60_47#_c_281_n N_Y_c_553_n 0.033448f $X=3.375 $Y=1.17 $X2=0 $Y2=0
cc_271 N_A_60_47#_c_273_n N_Y_c_555_n 0.00656525f $X=3.3 $Y=1.185 $X2=0 $Y2=0
cc_272 N_A_60_47#_c_275_n N_Y_c_555_n 4.4915e-19 $X=3.73 $Y=1.185 $X2=0 $Y2=0
cc_273 N_A_60_47#_c_273_n N_Y_c_593_n 0.00882151f $X=3.3 $Y=1.185 $X2=0 $Y2=0
cc_274 N_A_60_47#_c_275_n N_Y_c_593_n 0.0144821f $X=3.73 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A_60_47#_c_281_n N_Y_c_593_n 0.00843866f $X=3.375 $Y=1.17 $X2=0 $Y2=0
cc_276 N_A_60_47#_c_283_n N_Y_c_593_n 0.01729f $X=3.505 $Y=1.17 $X2=0 $Y2=0
cc_277 N_A_60_47#_c_285_n N_Y_c_593_n 5.4431e-19 $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_278 N_A_60_47#_M1003_g N_Y_c_561_n 0.00490528f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A_60_47#_M1007_g N_Y_c_561_n 0.0019458f $X=2.01 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A_60_47#_c_271_n N_Y_c_564_n 6.5926e-19 $X=2.01 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A_60_47#_c_281_n N_Y_c_564_n 0.0217194f $X=3.375 $Y=1.17 $X2=0 $Y2=0
cc_282 N_A_60_47#_c_273_n N_Y_c_565_n 7.17169e-19 $X=3.3 $Y=1.185 $X2=0 $Y2=0
cc_283 N_A_60_47#_c_281_n N_Y_c_565_n 0.0217194f $X=3.375 $Y=1.17 $X2=0 $Y2=0
cc_284 N_A_60_47#_c_275_n N_Y_c_539_n 9.41618e-19 $X=3.73 $Y=1.185 $X2=0 $Y2=0
cc_285 N_A_60_47#_c_283_n N_Y_c_539_n 0.00618498f $X=3.505 $Y=1.17 $X2=0 $Y2=0
cc_286 N_A_60_47#_M1011_g Y 0.0129469f $X=3.73 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A_60_47#_c_280_n N_VGND_M1012_d 0.00116574f $X=0.785 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_60_47#_c_279_n N_VGND_c_655_n 0.0145829f $X=1.565 $Y=1.17 $X2=0 $Y2=0
cc_289 N_A_60_47#_c_280_n N_VGND_c_655_n 0.0031614f $X=0.785 $Y=1.17 $X2=0 $Y2=0
cc_290 N_A_60_47#_c_269_n N_VGND_c_656_n 0.00280293f $X=1.58 $Y=1.185 $X2=0
+ $Y2=0
cc_291 N_A_60_47#_c_271_n N_VGND_c_656_n 0.00153274f $X=2.01 $Y=1.185 $X2=0
+ $Y2=0
cc_292 N_A_60_47#_c_271_n N_VGND_c_657_n 0.00428252f $X=2.01 $Y=1.185 $X2=0
+ $Y2=0
cc_293 N_A_60_47#_c_273_n N_VGND_c_659_n 0.00157435f $X=3.3 $Y=1.185 $X2=0 $Y2=0
cc_294 N_A_60_47#_c_275_n N_VGND_c_659_n 0.00720164f $X=3.73 $Y=1.185 $X2=0
+ $Y2=0
cc_295 N_A_60_47#_c_275_n N_VGND_c_661_n 5.96445e-19 $X=3.73 $Y=1.185 $X2=0
+ $Y2=0
cc_296 N_A_60_47#_c_269_n N_VGND_c_662_n 0.00428252f $X=1.58 $Y=1.185 $X2=0
+ $Y2=0
cc_297 N_A_60_47#_c_273_n N_VGND_c_664_n 0.00428252f $X=3.3 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A_60_47#_c_275_n N_VGND_c_666_n 0.00366311f $X=3.73 $Y=1.185 $X2=0
+ $Y2=0
cc_299 N_A_60_47#_c_277_n N_VGND_c_667_n 0.0178111f $X=0.425 $Y=0.42 $X2=0 $Y2=0
cc_300 N_A_60_47#_M1012_s N_VGND_c_669_n 0.00371702f $X=0.3 $Y=0.235 $X2=0 $Y2=0
cc_301 N_A_60_47#_c_269_n N_VGND_c_669_n 0.00587209f $X=1.58 $Y=1.185 $X2=0
+ $Y2=0
cc_302 N_A_60_47#_c_271_n N_VGND_c_669_n 0.00587209f $X=2.01 $Y=1.185 $X2=0
+ $Y2=0
cc_303 N_A_60_47#_c_273_n N_VGND_c_669_n 0.00587209f $X=3.3 $Y=1.185 $X2=0 $Y2=0
cc_304 N_A_60_47#_c_275_n N_VGND_c_669_n 0.00436859f $X=3.73 $Y=1.185 $X2=0
+ $Y2=0
cc_305 N_A_60_47#_c_277_n N_VGND_c_669_n 0.0100304f $X=0.425 $Y=0.42 $X2=0 $Y2=0
cc_306 N_VPWR_c_444_n N_A_245_367#_M1000_d 0.00491738f $X=2.655 $Y=2.55
+ $X2=-0.19 $Y2=-0.245
cc_307 N_VPWR_c_429_n N_A_245_367#_M1000_d 0.00223855f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_308 N_VPWR_c_444_n N_A_245_367#_M1007_d 0.00372618f $X=2.655 $Y=2.55 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_429_n N_A_245_367#_M1007_d 0.00223855f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_429_n N_A_245_367#_M1014_d 0.00223829f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_429_n N_A_245_367#_M1011_d 0.00376848f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_M1005_s N_A_245_367#_c_508_n 0.00339837f $X=2.515 $Y=1.835 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_444_n N_A_245_367#_c_508_n 0.0820672f $X=2.655 $Y=2.55 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_435_n N_A_245_367#_c_508_n 0.0939794f $X=4.21 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_429_n N_A_245_367#_c_508_n 0.0641898f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_435_n N_A_245_367#_c_513_n 0.0455271f $X=4.21 $Y=3.33 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_429_n N_A_245_367#_c_513_n 0.0305365f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_435_n N_A_245_367#_c_527_n 0.0121175f $X=4.21 $Y=3.33 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_429_n N_A_245_367#_c_527_n 0.0077417f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_444_n N_Y_M1003_s 0.00351361f $X=2.655 $Y=2.55 $X2=0 $Y2=0
cc_321 N_VPWR_c_429_n N_Y_M1003_s 0.00225465f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_322 N_VPWR_c_429_n N_Y_M1008_s 0.00225465f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_323 N_VPWR_M1005_s N_Y_c_547_n 0.00358342f $X=2.515 $Y=1.835 $X2=0 $Y2=0
cc_324 N_VPWR_c_444_n N_Y_c_547_n 0.0372465f $X=2.655 $Y=2.55 $X2=0 $Y2=0
cc_325 N_VPWR_c_444_n N_Y_c_561_n 0.0160416f $X=2.655 $Y=2.55 $X2=0 $Y2=0
cc_326 N_VPWR_M1015_s Y 0.00264236f $X=4.235 $Y=1.835 $X2=0 $Y2=0
cc_327 N_VPWR_M1015_s Y 0.00781961f $X=4.235 $Y=1.835 $X2=0 $Y2=0
cc_328 N_VPWR_c_432_n Y 0.0225014f $X=4.375 $Y=2.475 $X2=0 $Y2=0
cc_329 N_A_245_367#_c_508_n N_Y_M1003_s 0.00339837f $X=2.99 $Y=2.945 $X2=1.15
+ $Y2=1.675
cc_330 N_A_245_367#_c_513_n N_Y_M1008_s 0.00336401f $X=3.84 $Y=2.975 $X2=1.15
+ $Y2=2.465
cc_331 N_A_245_367#_M1007_d N_Y_c_547_n 0.00374812f $X=2.085 $Y=1.835 $X2=4.16
+ $Y2=1.345
cc_332 N_A_245_367#_M1014_d N_Y_c_547_n 0.00353353f $X=2.945 $Y=1.835 $X2=4.16
+ $Y2=1.345
cc_333 N_A_245_367#_c_508_n N_Y_c_547_n 0.00296302f $X=2.99 $Y=2.945 $X2=4.16
+ $Y2=1.345
cc_334 N_A_245_367#_c_534_p N_Y_c_547_n 0.0135217f $X=3.085 $Y=2.54 $X2=4.16
+ $Y2=1.345
cc_335 N_A_245_367#_c_513_n N_Y_c_622_n 0.0127409f $X=3.84 $Y=2.975 $X2=1.13
+ $Y2=1.51
cc_336 N_A_245_367#_M1011_d Y 0.00353353f $X=3.805 $Y=1.835 $X2=4.21 $Y2=1.675
cc_337 N_A_245_367#_c_537_p Y 0.0135217f $X=3.945 $Y=2.54 $X2=4.21 $Y2=1.675
cc_338 N_Y_c_578_n N_VGND_M1004_s 0.00329366f $X=2.06 $Y=0.83 $X2=0 $Y2=0
cc_339 N_Y_c_553_n N_VGND_M1002_d 0.00335318f $X=2.92 $Y=0.83 $X2=0 $Y2=0
cc_340 N_Y_c_593_n N_VGND_M1010_s 0.00329366f $X=3.84 $Y=0.83 $X2=0 $Y2=0
cc_341 N_Y_c_538_n N_VGND_M1016_d 0.00253355f $X=4.475 $Y=1.09 $X2=0 $Y2=0
cc_342 N_Y_c_578_n N_VGND_c_656_n 0.0130506f $X=2.06 $Y=0.83 $X2=0 $Y2=0
cc_343 N_Y_c_578_n N_VGND_c_657_n 0.00191958f $X=2.06 $Y=0.83 $X2=0 $Y2=0
cc_344 N_Y_c_551_n N_VGND_c_657_n 0.0188913f $X=2.225 $Y=0.42 $X2=0 $Y2=0
cc_345 N_Y_c_553_n N_VGND_c_657_n 0.00191958f $X=2.92 $Y=0.83 $X2=0 $Y2=0
cc_346 N_Y_c_553_n N_VGND_c_658_n 0.0130506f $X=2.92 $Y=0.83 $X2=0 $Y2=0
cc_347 N_Y_c_593_n N_VGND_c_659_n 0.0147753f $X=3.84 $Y=0.83 $X2=0 $Y2=0
cc_348 N_Y_c_538_n N_VGND_c_661_n 0.0225465f $X=4.475 $Y=1.09 $X2=0 $Y2=0
cc_349 N_Y_c_545_n N_VGND_c_662_n 0.0188913f $X=1.365 $Y=0.42 $X2=0 $Y2=0
cc_350 N_Y_c_578_n N_VGND_c_662_n 0.00191958f $X=2.06 $Y=0.83 $X2=0 $Y2=0
cc_351 N_Y_c_553_n N_VGND_c_664_n 0.00191958f $X=2.92 $Y=0.83 $X2=0 $Y2=0
cc_352 N_Y_c_555_n N_VGND_c_664_n 0.0188913f $X=3.085 $Y=0.42 $X2=0 $Y2=0
cc_353 N_Y_c_593_n N_VGND_c_664_n 0.00191958f $X=3.84 $Y=0.83 $X2=0 $Y2=0
cc_354 N_Y_c_593_n N_VGND_c_666_n 0.00184586f $X=3.84 $Y=0.83 $X2=0 $Y2=0
cc_355 N_Y_c_642_p N_VGND_c_666_n 0.0120977f $X=3.945 $Y=0.42 $X2=0 $Y2=0
cc_356 N_Y_M1001_s N_VGND_c_669_n 0.00223559f $X=1.225 $Y=0.235 $X2=0 $Y2=0
cc_357 N_Y_M1006_d N_VGND_c_669_n 0.00223559f $X=2.085 $Y=0.235 $X2=0 $Y2=0
cc_358 N_Y_M1009_s N_VGND_c_669_n 0.00223559f $X=2.945 $Y=0.235 $X2=0 $Y2=0
cc_359 N_Y_M1017_d N_VGND_c_669_n 0.00435668f $X=3.805 $Y=0.235 $X2=0 $Y2=0
cc_360 N_Y_c_545_n N_VGND_c_669_n 0.012376f $X=1.365 $Y=0.42 $X2=0 $Y2=0
cc_361 N_Y_c_578_n N_VGND_c_669_n 0.00827851f $X=2.06 $Y=0.83 $X2=0 $Y2=0
cc_362 N_Y_c_551_n N_VGND_c_669_n 0.012376f $X=2.225 $Y=0.42 $X2=0 $Y2=0
cc_363 N_Y_c_553_n N_VGND_c_669_n 0.00827851f $X=2.92 $Y=0.83 $X2=0 $Y2=0
cc_364 N_Y_c_555_n N_VGND_c_669_n 0.012376f $X=3.085 $Y=0.42 $X2=0 $Y2=0
cc_365 N_Y_c_593_n N_VGND_c_669_n 0.00829644f $X=3.84 $Y=0.83 $X2=0 $Y2=0
cc_366 N_Y_c_642_p N_VGND_c_669_n 0.00691495f $X=3.945 $Y=0.42 $X2=0 $Y2=0
cc_367 N_Y_c_539_n N_VGND_c_669_n 2.3963e-19 $X=3.935 $Y=0.83 $X2=0 $Y2=0
