# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.190000 1.815000 1.800000 2.075000 ;
        RECT 1.515000 0.385000 1.800000 1.815000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.898800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.110000 0.255000 14.775000 1.095000 ;
        RECT 14.525000 1.095000 14.775000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.155000 0.265000 12.460000 1.815000 ;
        RECT 12.155000 1.815000 12.585000 2.120000 ;
        RECT 12.290000 2.120000 12.585000 3.075000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.510000 1.535000 2.890000 2.250000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 1.155000 0.885000 2.245000 ;
        RECT 0.555000 2.245000 2.340000 2.415000 ;
        RECT 0.555000 2.415000 0.985000 2.490000 ;
        RECT 2.090000 1.165000 2.340000 2.245000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.295000 1.920000  7.585000 1.965000 ;
        RECT  7.295000 1.965000 10.945000 2.105000 ;
        RECT  7.295000 2.105000  7.585000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.995000 0.775000 3.380000 1.025000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.245000 15.360000 3.415000 ;
      RECT  0.095000  0.275000  0.660000 0.815000 ;
      RECT  0.095000  0.815000  1.345000 0.985000 ;
      RECT  0.095000  0.985000  0.355000 2.985000 ;
      RECT  0.525000  2.660000  0.855000 3.245000 ;
      RECT  0.830000  0.085000  1.160000 0.605000 ;
      RECT  1.055000  0.985000  1.345000 1.485000 ;
      RECT  1.425000  2.585000  3.230000 2.805000 ;
      RECT  1.970000  0.280000  2.220000 0.705000 ;
      RECT  1.970000  0.705000  2.690000 0.875000 ;
      RECT  2.445000  2.975000  2.775000 3.245000 ;
      RECT  2.520000  0.875000  2.690000 1.195000 ;
      RECT  2.520000  1.195000  3.230000 1.365000 ;
      RECT  2.690000  0.085000  3.020000 0.535000 ;
      RECT  3.060000  1.365000  3.230000 2.585000 ;
      RECT  3.060000  2.805000  3.930000 2.995000 ;
      RECT  3.190000  0.275000  3.940000 0.605000 ;
      RECT  3.400000  1.195000  4.405000 1.565000 ;
      RECT  3.400000  1.565000  3.590000 2.635000 ;
      RECT  3.550000  0.605000  3.940000 0.895000 ;
      RECT  3.550000  0.895000  4.405000 1.195000 ;
      RECT  3.760000  2.335000  5.655000 2.360000 ;
      RECT  3.760000  2.360000  5.780000 2.505000 ;
      RECT  3.760000  2.505000  3.930000 2.805000 ;
      RECT  4.100000  2.675000  4.360000 3.245000 ;
      RECT  4.145000  0.085000  4.405000 0.725000 ;
      RECT  4.575000  0.410000  4.905000 1.485000 ;
      RECT  4.575000  1.485000  5.295000 2.165000 ;
      RECT  5.360000  0.640000  5.655000 1.235000 ;
      RECT  5.475000  1.235000  5.655000 2.335000 ;
      RECT  5.475000  2.505000  5.780000 2.705000 ;
      RECT  5.825000  0.640000  6.120000 1.140000 ;
      RECT  5.825000  1.140000  7.505000 1.205000 ;
      RECT  5.825000  1.205000  8.575000 1.345000 ;
      RECT  5.825000  1.345000  5.995000 2.020000 ;
      RECT  5.825000  2.020000  6.250000 2.190000 ;
      RECT  5.950000  2.190000  6.250000 2.690000 ;
      RECT  6.165000  1.515000  6.430000 1.545000 ;
      RECT  6.165000  1.545000  8.215000 1.725000 ;
      RECT  6.165000  1.725000  6.425000 1.845000 ;
      RECT  6.580000  0.085000  6.910000 0.970000 ;
      RECT  6.635000  1.905000  6.965000 2.300000 ;
      RECT  6.635000  2.300000  9.485000 2.375000 ;
      RECT  6.635000  2.375000  8.215000 2.470000 ;
      RECT  6.790000  2.640000  7.120000 3.245000 ;
      RECT  7.175000  1.345000  8.575000 1.375000 ;
      RECT  7.255000  0.640000  7.960000 0.865000 ;
      RECT  7.255000  0.865000  8.915000 0.970000 ;
      RECT  7.265000  1.895000  7.865000 2.130000 ;
      RECT  7.300000  2.470000  7.630000 2.690000 ;
      RECT  7.790000  0.970000  8.915000 1.030000 ;
      RECT  7.790000  1.030000  9.485000 1.035000 ;
      RECT  7.950000  2.640000  8.280000 3.245000 ;
      RECT  8.045000  1.725000  8.215000 1.855000 ;
      RECT  8.045000  1.855000  9.145000 2.025000 ;
      RECT  8.045000  2.205000  9.485000 2.300000 ;
      RECT  8.140000  0.085000  8.470000 0.695000 ;
      RECT  8.385000  1.375000  8.575000 1.675000 ;
      RECT  8.745000  1.035000  9.485000 1.200000 ;
      RECT  8.885000  1.370000  9.145000 1.855000 ;
      RECT  8.970000  2.555000  9.835000 2.885000 ;
      RECT  9.135000  0.590000  9.835000 0.860000 ;
      RECT  9.315000  1.200000  9.485000 2.205000 ;
      RECT  9.665000  0.860000  9.835000 2.155000 ;
      RECT  9.665000  2.155000 10.535000 2.335000 ;
      RECT  9.665000  2.335000  9.835000 2.555000 ;
      RECT 10.005000  2.505000 10.195000 3.245000 ;
      RECT 10.015000  1.085000 11.925000 1.255000 ;
      RECT 10.015000  1.255000 10.345000 1.845000 ;
      RECT 10.340000  0.085000 10.670000 0.915000 ;
      RECT 10.365000  2.335000 10.535000 2.505000 ;
      RECT 10.365000  2.505000 11.235000 2.835000 ;
      RECT 10.705000  1.630000 10.895000 2.300000 ;
      RECT 11.065000  1.425000 11.575000 1.645000 ;
      RECT 11.065000  1.645000 11.235000 2.505000 ;
      RECT 11.120000  0.710000 11.380000 1.085000 ;
      RECT 11.415000  1.815000 11.925000 2.145000 ;
      RECT 11.550000  0.085000 11.985000 0.915000 ;
      RECT 11.755000  1.255000 11.925000 1.815000 ;
      RECT 11.860000  2.315000 12.120000 3.245000 ;
      RECT 12.630000  0.085000 12.965000 1.105000 ;
      RECT 12.755000  1.815000 13.095000 3.245000 ;
      RECT 13.135000  0.290000 13.475000 0.620000 ;
      RECT 13.265000  0.620000 13.475000 1.275000 ;
      RECT 13.265000  1.275000 14.355000 1.605000 ;
      RECT 13.265000  1.605000 13.575000 2.495000 ;
      RECT 13.655000  0.085000 13.940000 1.095000 ;
      RECT 14.025000  1.820000 14.355000 3.245000 ;
      RECT 14.945000  0.085000 15.215000 1.095000 ;
      RECT 14.945000  1.820000 15.215000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.950000  7.525000 2.120000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfsbp_2
