# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxbn_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.450000 1.210000 0.910000 1.880000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 0.655000 8.045000 2.135000 ;
        RECT 7.775000 0.330000 8.045000 0.655000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765000 0.965000 7.095000 3.075000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.320000 1.610000 0.650000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.640000 0.085000 ;
        RECT 0.655000  0.085000 0.875000 1.040000 ;
        RECT 2.220000  0.085000 2.550000 0.455000 ;
        RECT 4.265000  0.085000 4.595000 0.885000 ;
        RECT 6.220000  0.085000 6.550000 0.455000 ;
        RECT 7.275000  0.085000 7.605000 0.455000 ;
        RECT 8.215000  0.085000 8.545000 1.125000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.640000 3.415000 ;
        RECT 0.685000 2.495000 1.015000 3.245000 ;
        RECT 2.340000 2.835000 2.670000 3.245000 ;
        RECT 4.245000 2.235000 4.835000 3.245000 ;
        RECT 6.135000 1.795000 6.585000 3.245000 ;
        RECT 7.265000 2.645000 7.595000 3.245000 ;
        RECT 8.135000 2.645000 8.465000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 0.700000 0.485000 1.040000 ;
      RECT 0.110000 1.040000 0.280000 2.060000 ;
      RECT 0.110000 2.060000 0.530000 2.155000 ;
      RECT 0.110000 2.155000 2.760000 2.325000 ;
      RECT 0.110000 2.325000 0.515000 2.730000 ;
      RECT 1.045000 0.820000 1.400000 0.965000 ;
      RECT 1.045000 0.965000 3.210000 1.090000 ;
      RECT 1.230000 1.090000 3.210000 1.375000 ;
      RECT 1.230000 1.375000 2.185000 1.955000 ;
      RECT 1.230000 1.955000 1.560000 1.985000 ;
      RECT 1.770000 2.495000 3.100000 2.665000 ;
      RECT 1.770000 2.665000 2.100000 3.075000 ;
      RECT 1.780000 0.280000 2.050000 0.625000 ;
      RECT 1.780000 0.625000 3.620000 0.795000 ;
      RECT 2.435000 1.625000 2.760000 2.155000 ;
      RECT 2.930000 1.965000 3.620000 2.220000 ;
      RECT 2.930000 2.220000 3.100000 2.495000 ;
      RECT 2.935000 1.375000 3.210000 1.755000 ;
      RECT 3.150000 0.255000 3.960000 0.455000 ;
      RECT 3.280000 2.390000 3.960000 2.560000 ;
      RECT 3.280000 2.560000 3.610000 3.075000 ;
      RECT 3.380000 0.795000 3.620000 1.965000 ;
      RECT 3.790000 0.455000 3.960000 1.055000 ;
      RECT 3.790000 1.055000 4.675000 1.225000 ;
      RECT 3.790000 1.225000 3.960000 2.390000 ;
      RECT 4.130000 1.395000 4.335000 1.795000 ;
      RECT 4.130000 1.795000 5.265000 2.065000 ;
      RECT 4.505000 1.225000 4.675000 1.295000 ;
      RECT 4.505000 1.295000 4.915000 1.625000 ;
      RECT 4.845000 0.255000 6.040000 0.455000 ;
      RECT 4.845000 0.455000 5.265000 1.125000 ;
      RECT 5.005000 2.065000 5.265000 3.075000 ;
      RECT 5.085000 1.125000 5.265000 1.795000 ;
      RECT 5.670000 0.965000 6.000000 1.295000 ;
      RECT 5.670000 1.295000 6.585000 1.625000 ;
      RECT 5.670000 1.625000 5.965000 2.485000 ;
      RECT 5.710000 0.455000 6.040000 0.625000 ;
      RECT 5.710000 0.625000 7.445000 0.795000 ;
      RECT 7.275000 0.795000 7.445000 2.305000 ;
      RECT 7.275000 2.305000 8.490000 2.475000 ;
      RECT 8.225000 1.295000 8.490000 2.305000 ;
  END
END sky130_fd_sc_lp__dlxbn_2
