* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_823_367# B2 a_547_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 X a_547_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND A2 a_44_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR B1 a_823_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_547_367# B2 a_44_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_823_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_112_367# A2 a_195_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 X a_547_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR a_547_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_112_367# A3 a_547_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_195_367# A2 a_112_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND a_547_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR A1 a_195_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 X a_547_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_195_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_547_367# B1 a_44_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND a_547_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_44_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VGND A3 a_44_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_547_367# A3 a_112_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VGND A1 a_44_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_44_65# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_44_65# B1 a_547_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 X a_547_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_547_367# B2 a_823_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VPWR a_547_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_44_65# B2 a_547_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_44_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
