* File: sky130_fd_sc_lp__dlrbn_lp.spice
* Created: Fri Aug 28 10:25:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrbn_lp.pex.spice"
.subckt sky130_fd_sc_lp__dlrbn_lp  VNB VPB D GATE_N RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1015 A_114_68# N_D_M1015_g N_A_27_68#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_D_M1002_g A_114_68# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1018 A_272_68# N_GATE_N_M1018_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_A_252_396#_M1019_d N_GATE_N_M1019_g A_272_68# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 A_542_47# N_A_252_396#_M1021_g N_A_451_419#_M1021_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_252_396#_M1007_g A_542_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=0.99 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1011 A_758_47# N_A_27_68#_M1011_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=0.99 NRD=18.564 NRS=82.848 M=1 R=2.8 SA=75001.3
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1012 N_A_796_419#_M1012_d N_A_252_396#_M1012_g A_758_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8
+ SA=75001.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1022 A_950_47# N_A_451_419#_M1022_g N_A_796_419#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0882 PD=0.81 PS=0.84 NRD=39.996 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_952_305#_M1029_g A_950_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1626 AS=0.0819 PD=1.64 PS=0.81 NRD=22.848 NRS=39.996 M=1 R=2.8 SA=75002.8
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1024 A_1277_153# N_A_796_419#_M1024_g N_A_952_305#_M1024_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_RESET_B_M1010_g A_1277_153# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1014 A_1435_153# N_A_952_305#_M1014_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_Q_M1008_d N_A_952_305#_M1008_g A_1435_153# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_1703_76# N_A_952_305#_M1004_g N_A_1617_76#_M1004_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_952_305#_M1006_g A_1703_76# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1023 A_1861_76# N_A_1617_76#_M1023_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_Q_N_M1025_d N_A_1617_76#_M1025_g A_1861_76# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_D_M1013_g N_A_27_68#_M1013_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_252_396#_M1003_d N_GATE_N_M1003_g N_VPWR_M1013_d VPB PHIGHVT L=0.25
+ W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1017 N_VPWR_M1017_d N_A_252_396#_M1017_g N_A_451_419#_M1017_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.225 AS=0.285 PD=1.45 PS=2.57 NRD=33.4703 NRS=0 M=1 R=4
+ SA=125000 SB=125005 A=0.25 P=2.5 MULT=1
MM1020 A_698_419# N_A_27_68#_M1020_g N_VPWR_M1017_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.225 PD=1.24 PS=1.45 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_796_419#_M1000_d N_A_451_419#_M1000_g A_698_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.145 AS=0.12 PD=1.29 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1009 A_904_419# N_A_252_396#_M1009_g N_A_796_419#_M1000_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.145 PD=1.24 PS=1.29 NRD=12.7853 NRS=0 M=1 R=4 SA=125002
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1026 N_VPWR_M1026_d N_A_952_305#_M1026_g A_904_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.295 AS=0.12 PD=1.59 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1005 N_A_952_305#_M1005_d N_A_796_419#_M1005_g N_VPWR_M1026_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.295 PD=1.28 PS=1.59 NRD=0 NRS=61.0503 M=1 R=4
+ SA=125003 SB=125002 A=0.25 P=2.5 MULT=1
MM1028 N_VPWR_M1028_d N_RESET_B_M1028_g N_A_952_305#_M1005_d VPB PHIGHVT L=0.25
+ W=1 AD=0.56 AS=0.14 PD=2.12 PS=1.28 NRD=165.48 NRS=0 M=1 R=4 SA=125004
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1001 N_Q_M1001_d N_A_952_305#_M1001_g N_VPWR_M1028_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.56 PD=2.57 PS=2.12 NRD=0 NRS=0 M=1 R=4 SA=125005 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1027 N_VPWR_M1027_d N_A_952_305#_M1027_g N_A_1617_76#_M1027_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1016 N_Q_N_M1016_d N_A_1617_76#_M1016_g N_VPWR_M1027_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX30_noxref VNB VPB NWDIODE A=19.5079 P=24.65
*
.include "sky130_fd_sc_lp__dlrbn_lp.pxi.spice"
*
.ends
*
*
