* File: sky130_fd_sc_lp__a2bb2o_0.pxi.spice
* Created: Wed Sep  2 09:23:36 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2O_0%A_59_194# N_A_59_194#_M1006_d N_A_59_194#_M1011_s
+ N_A_59_194#_c_95_n N_A_59_194#_M1003_g N_A_59_194#_c_96_n N_A_59_194#_c_97_n
+ N_A_59_194#_M1000_g N_A_59_194#_c_102_n N_A_59_194#_c_103_n
+ N_A_59_194#_c_104_n N_A_59_194#_c_105_n N_A_59_194#_c_106_n
+ N_A_59_194#_c_135_p N_A_59_194#_c_99_n N_A_59_194#_c_108_n N_A_59_194#_c_109_n
+ PM_SKY130_FD_SC_LP__A2BB2O_0%A_59_194#
x_PM_SKY130_FD_SC_LP__A2BB2O_0%A1_N N_A1_N_c_196_n N_A1_N_M1004_g N_A1_N_M1009_g
+ N_A1_N_c_197_n N_A1_N_c_198_n A1_N A1_N A1_N N_A1_N_c_200_n
+ PM_SKY130_FD_SC_LP__A2BB2O_0%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2O_0%A2_N N_A2_N_M1010_g N_A2_N_M1001_g N_A2_N_c_255_n
+ N_A2_N_c_259_n A2_N A2_N N_A2_N_c_257_n PM_SKY130_FD_SC_LP__A2BB2O_0%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2O_0%A_237_47# N_A_237_47#_M1009_d N_A_237_47#_M1010_d
+ N_A_237_47#_M1006_g N_A_237_47#_c_315_n N_A_237_47#_c_316_n
+ N_A_237_47#_c_317_n N_A_237_47#_M1011_g N_A_237_47#_c_307_n
+ N_A_237_47#_c_320_n N_A_237_47#_c_308_n N_A_237_47#_c_309_n
+ N_A_237_47#_c_310_n N_A_237_47#_c_321_n N_A_237_47#_c_311_n
+ N_A_237_47#_c_312_n N_A_237_47#_c_313_n N_A_237_47#_c_323_n
+ N_A_237_47#_c_314_n N_A_237_47#_c_324_n PM_SKY130_FD_SC_LP__A2BB2O_0%A_237_47#
x_PM_SKY130_FD_SC_LP__A2BB2O_0%B2 N_B2_M1007_g N_B2_M1005_g B2 B2 B2 B2
+ N_B2_c_392_n PM_SKY130_FD_SC_LP__A2BB2O_0%B2
x_PM_SKY130_FD_SC_LP__A2BB2O_0%B1 N_B1_c_432_n N_B1_M1008_g N_B1_c_433_n
+ N_B1_c_434_n N_B1_M1002_g N_B1_c_436_n B1 B1 B1 B1 B1 N_B1_c_438_n
+ PM_SKY130_FD_SC_LP__A2BB2O_0%B1
x_PM_SKY130_FD_SC_LP__A2BB2O_0%X N_X_M1000_s N_X_M1003_s N_X_c_468_n X X X X X X
+ X PM_SKY130_FD_SC_LP__A2BB2O_0%X
x_PM_SKY130_FD_SC_LP__A2BB2O_0%VPWR N_VPWR_M1003_d N_VPWR_M1005_d N_VPWR_c_496_n
+ N_VPWR_c_497_n VPWR N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_495_n N_VPWR_c_502_n N_VPWR_c_503_n PM_SKY130_FD_SC_LP__A2BB2O_0%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2O_0%A_516_535# N_A_516_535#_M1011_d
+ N_A_516_535#_M1002_d N_A_516_535#_c_546_n N_A_516_535#_c_547_n
+ N_A_516_535#_c_548_n N_A_516_535#_c_549_n
+ PM_SKY130_FD_SC_LP__A2BB2O_0%A_516_535#
x_PM_SKY130_FD_SC_LP__A2BB2O_0%VGND N_VGND_M1000_d N_VGND_M1001_d N_VGND_M1008_d
+ N_VGND_c_572_n N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n N_VGND_c_576_n
+ N_VGND_c_577_n VGND N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n
+ N_VGND_c_581_n N_VGND_c_582_n PM_SKY130_FD_SC_LP__A2BB2O_0%VGND
cc_1 VNB N_A_59_194#_c_95_n 0.0327876f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.93
cc_2 VNB N_A_59_194#_c_96_n 0.0198695f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.045
cc_3 VNB N_A_59_194#_c_97_n 0.0111043f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.045
cc_4 VNB N_A_59_194#_M1000_g 0.031025f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.445
cc_5 VNB N_A_59_194#_c_99_n 0.00697405f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.075
cc_6 VNB N_A1_N_c_196_n 0.0233696f $X=-0.19 $Y=-0.245 $X2=2.165 $Y2=2.675
cc_7 VNB N_A1_N_c_197_n 0.0167333f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.77
cc_8 VNB N_A1_N_c_198_n 0.0126653f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.77
cc_9 VNB A1_N 0.0121937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_N_c_200_n 0.0273921f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.095
cc_11 VNB N_A2_N_M1001_g 0.0390271f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.12
cc_12 VNB N_A2_N_c_255_n 0.0210424f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.77
cc_13 VNB A2_N 0.0041829f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.045
cc_14 VNB N_A2_N_c_257_n 0.0159034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_237_47#_M1006_g 0.0448374f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.26
cc_16 VNB N_A_237_47#_c_307_n 0.0163505f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.095
cc_17 VNB N_A_237_47#_c_308_n 0.00280087f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.88
cc_18 VNB N_A_237_47#_c_309_n 0.0132721f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.965
cc_19 VNB N_A_237_47#_c_310_n 0.00407421f $X=-0.19 $Y=-0.245 $X2=2.302 $Y2=2.245
cc_20 VNB N_A_237_47#_c_311_n 0.00221284f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.445
cc_21 VNB N_A_237_47#_c_312_n 0.00160777f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.245
cc_22 VNB N_A_237_47#_c_313_n 0.0159705f $X=-0.19 $Y=-0.245 $X2=2.302 $Y2=2.965
cc_23 VNB N_A_237_47#_c_314_n 0.00454865f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.095
cc_24 VNB N_B2_M1007_g 0.0366674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB B2 0.00985248f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.26
cc_26 VNB N_B2_c_392_n 0.0539929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_c_432_n 0.0188191f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=0.235
cc_28 VNB N_B1_c_433_n 0.0425904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_c_434_n 0.00596089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_M1002_g 0.00183788f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.93
cc_31 VNB N_B1_c_436_n 0.0242645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB B1 0.0557f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.045
cc_33 VNB N_B1_c_438_n 0.0483171f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.26
cc_34 VNB N_X_c_468_n 0.0179499f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.77
cc_35 VNB X 0.043387f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.045
cc_36 VNB N_VPWR_c_495_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=0.445
cc_37 VNB N_VGND_c_572_n 0.00465702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_573_n 0.0177423f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.045
cc_39 VNB N_VGND_c_574_n 0.00500436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_575_n 0.00251179f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.095
cc_41 VNB N_VGND_c_576_n 0.021923f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.26
cc_42 VNB N_VGND_c_577_n 0.00497572f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.88
cc_43 VNB N_VGND_c_578_n 0.027394f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=0.445
cc_44 VNB N_VGND_c_579_n 0.01856f $X=-0.19 $Y=-0.245 $X2=2.302 $Y2=2.965
cc_45 VNB N_VGND_c_580_n 0.214536f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=2.885
cc_46 VNB N_VGND_c_581_n 0.00632231f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.095
cc_47 VNB N_VGND_c_582_n 0.00395493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_A_59_194#_c_95_n 0.016784f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.93
cc_49 VPB N_A_59_194#_M1003_g 0.0275018f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.77
cc_50 VPB N_A_59_194#_c_102_n 0.00927654f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=2.095
cc_51 VPB N_A_59_194#_c_103_n 0.00341265f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.88
cc_52 VPB N_A_59_194#_c_104_n 0.019158f $X=-0.19 $Y=1.655 $X2=2.185 $Y2=2.965
cc_53 VPB N_A_59_194#_c_105_n 0.00254213f $X=-0.19 $Y=1.655 $X2=1.31 $Y2=2.965
cc_54 VPB N_A_59_194#_c_106_n 0.00868471f $X=-0.19 $Y=1.655 $X2=2.302 $Y2=2.88
cc_55 VPB N_A_59_194#_c_99_n 0.00447633f $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.075
cc_56 VPB N_A_59_194#_c_108_n 6.4611e-19 $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.245
cc_57 VPB N_A_59_194#_c_109_n 0.0446692f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.095
cc_58 VPB N_A1_N_M1004_g 0.047763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB A1_N 0.00415569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A1_N_c_200_n 0.00907134f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.095
cc_61 VPB N_A2_N_M1010_g 0.0486712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A2_N_c_259_n 0.0178564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB A2_N 0.00246263f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.045
cc_64 VPB N_A_237_47#_c_315_n 0.0112533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_237_47#_c_316_n 0.0249515f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.045
cc_66 VPB N_A_237_47#_c_317_n 0.0117573f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.045
cc_67 VPB N_A_237_47#_M1011_g 0.0392998f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.445
cc_68 VPB N_A_237_47#_c_307_n 0.00540727f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.095
cc_69 VPB N_A_237_47#_c_320_n 0.0170565f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.095
cc_70 VPB N_A_237_47#_c_321_n 0.0151865f $X=-0.19 $Y=1.655 $X2=2.302 $Y2=2.88
cc_71 VPB N_A_237_47#_c_312_n 5.52478e-19 $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.245
cc_72 VPB N_A_237_47#_c_323_n 0.0108712f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.93
cc_73 VPB N_A_237_47#_c_324_n 0.00460777f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.095
cc_74 VPB N_B2_M1005_g 0.0527667f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.12
cc_75 VPB B2 0.010674f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.26
cc_76 VPB N_B2_c_392_n 0.0253405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_B1_M1002_g 0.0805493f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.93
cc_78 VPB B1 0.0255992f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.045
cc_79 VPB X 0.0321746f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.045
cc_80 VPB X 0.00841927f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.445
cc_81 VPB X 0.0191643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_496_n 0.0101534f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.26
cc_83 VPB N_VPWR_c_497_n 0.00524934f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.045
cc_84 VPB N_VPWR_c_498_n 0.0182217f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.445
cc_85 VPB N_VPWR_c_499_n 0.0509229f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.095
cc_86 VPB N_VPWR_c_500_n 0.0165716f $X=-0.19 $Y=1.655 $X2=2.325 $Y2=0.445
cc_87 VPB N_VPWR_c_495_n 0.0569166f $X=-0.19 $Y=1.655 $X2=2.325 $Y2=0.445
cc_88 VPB N_VPWR_c_502_n 0.00679912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_503_n 0.00507051f $X=-0.19 $Y=1.655 $X2=2.302 $Y2=2.965
cc_90 VPB N_A_516_535#_c_546_n 0.00153267f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.26
cc_91 VPB N_A_516_535#_c_547_n 0.0180563f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.77
cc_92 VPB N_A_516_535#_c_548_n 0.00483007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_516_535#_c_549_n 0.0189967f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.97
cc_94 N_A_59_194#_c_95_n N_A1_N_c_196_n 0.00201508f $X=0.37 $Y=1.93 $X2=0 $Y2=0
cc_95 N_A_59_194#_c_96_n N_A1_N_c_196_n 0.0104484f $X=0.605 $Y=1.045 $X2=0 $Y2=0
cc_96 N_A_59_194#_c_95_n N_A1_N_M1004_g 0.00286399f $X=0.37 $Y=1.93 $X2=0 $Y2=0
cc_97 N_A_59_194#_M1003_g N_A1_N_M1004_g 0.0113426f $X=0.495 $Y=2.77 $X2=0 $Y2=0
cc_98 N_A_59_194#_c_102_n N_A1_N_M1004_g 0.0238583f $X=1.14 $Y=2.095 $X2=0 $Y2=0
cc_99 N_A_59_194#_c_103_n N_A1_N_M1004_g 0.00593714f $X=1.225 $Y=2.88 $X2=0
+ $Y2=0
cc_100 N_A_59_194#_c_105_n N_A1_N_M1004_g 9.63942e-19 $X=1.31 $Y=2.965 $X2=0
+ $Y2=0
cc_101 N_A_59_194#_c_109_n N_A1_N_M1004_g 0.0213522f $X=0.495 $Y=2.095 $X2=0
+ $Y2=0
cc_102 N_A_59_194#_M1000_g N_A1_N_c_197_n 0.0129369f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_103 N_A_59_194#_M1000_g N_A1_N_c_198_n 0.0104484f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_104 N_A_59_194#_c_95_n A1_N 0.00459074f $X=0.37 $Y=1.93 $X2=0 $Y2=0
cc_105 N_A_59_194#_c_96_n A1_N 0.0120439f $X=0.605 $Y=1.045 $X2=0 $Y2=0
cc_106 N_A_59_194#_M1000_g A1_N 0.010689f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_59_194#_c_102_n A1_N 0.0347234f $X=1.14 $Y=2.095 $X2=0 $Y2=0
cc_108 N_A_59_194#_c_109_n A1_N 0.00419868f $X=0.495 $Y=2.095 $X2=0 $Y2=0
cc_109 N_A_59_194#_c_95_n N_A1_N_c_200_n 0.0162994f $X=0.37 $Y=1.93 $X2=0 $Y2=0
cc_110 N_A_59_194#_c_96_n N_A1_N_c_200_n 0.00386578f $X=0.605 $Y=1.045 $X2=0
+ $Y2=0
cc_111 N_A_59_194#_c_102_n N_A1_N_c_200_n 0.0023418f $X=1.14 $Y=2.095 $X2=0
+ $Y2=0
cc_112 N_A_59_194#_c_109_n N_A1_N_c_200_n 0.00368758f $X=0.495 $Y=2.095 $X2=0
+ $Y2=0
cc_113 N_A_59_194#_c_102_n N_A2_N_M1010_g 0.00468085f $X=1.14 $Y=2.095 $X2=0
+ $Y2=0
cc_114 N_A_59_194#_c_103_n N_A2_N_M1010_g 0.0038169f $X=1.225 $Y=2.88 $X2=0
+ $Y2=0
cc_115 N_A_59_194#_c_104_n N_A2_N_M1010_g 0.0136076f $X=2.185 $Y=2.965 $X2=0
+ $Y2=0
cc_116 N_A_59_194#_c_106_n N_A2_N_M1010_g 0.00297994f $X=2.302 $Y=2.88 $X2=0
+ $Y2=0
cc_117 N_A_59_194#_c_108_n N_A2_N_M1010_g 2.28469e-19 $X=2.34 $Y=2.245 $X2=0
+ $Y2=0
cc_118 N_A_59_194#_c_102_n A2_N 0.0179025f $X=1.14 $Y=2.095 $X2=0 $Y2=0
cc_119 N_A_59_194#_c_135_p N_A_237_47#_M1006_g 0.00477325f $X=2.41 $Y=0.445
+ $X2=0 $Y2=0
cc_120 N_A_59_194#_c_99_n N_A_237_47#_M1006_g 0.00701897f $X=2.34 $Y=2.075 $X2=0
+ $Y2=0
cc_121 N_A_59_194#_c_99_n N_A_237_47#_c_316_n 0.00402232f $X=2.34 $Y=2.075 $X2=0
+ $Y2=0
cc_122 N_A_59_194#_c_108_n N_A_237_47#_c_316_n 0.0139788f $X=2.34 $Y=2.245 $X2=0
+ $Y2=0
cc_123 N_A_59_194#_c_104_n N_A_237_47#_c_317_n 0.00273032f $X=2.185 $Y=2.965
+ $X2=0 $Y2=0
cc_124 N_A_59_194#_c_108_n N_A_237_47#_c_317_n 0.00466008f $X=2.34 $Y=2.245
+ $X2=0 $Y2=0
cc_125 N_A_59_194#_c_106_n N_A_237_47#_M1011_g 0.013571f $X=2.302 $Y=2.88 $X2=0
+ $Y2=0
cc_126 N_A_59_194#_c_108_n N_A_237_47#_M1011_g 0.00449554f $X=2.34 $Y=2.245
+ $X2=0 $Y2=0
cc_127 N_A_59_194#_c_99_n N_A_237_47#_c_309_n 0.0105757f $X=2.34 $Y=2.075 $X2=0
+ $Y2=0
cc_128 N_A_59_194#_c_103_n N_A_237_47#_c_321_n 0.0119385f $X=1.225 $Y=2.88 $X2=0
+ $Y2=0
cc_129 N_A_59_194#_c_104_n N_A_237_47#_c_321_n 0.0370849f $X=2.185 $Y=2.965
+ $X2=0 $Y2=0
cc_130 N_A_59_194#_c_106_n N_A_237_47#_c_321_n 0.0226955f $X=2.302 $Y=2.88 $X2=0
+ $Y2=0
cc_131 N_A_59_194#_c_99_n N_A_237_47#_c_311_n 0.0500828f $X=2.34 $Y=2.075 $X2=0
+ $Y2=0
cc_132 N_A_59_194#_c_99_n N_A_237_47#_c_313_n 0.00668054f $X=2.34 $Y=2.075 $X2=0
+ $Y2=0
cc_133 N_A_59_194#_c_102_n N_A_237_47#_c_323_n 0.0126249f $X=1.14 $Y=2.095 $X2=0
+ $Y2=0
cc_134 N_A_59_194#_c_103_n N_A_237_47#_c_323_n 0.0057828f $X=1.225 $Y=2.88 $X2=0
+ $Y2=0
cc_135 N_A_59_194#_c_99_n N_A_237_47#_c_323_n 0.00815338f $X=2.34 $Y=2.075 $X2=0
+ $Y2=0
cc_136 N_A_59_194#_c_108_n N_A_237_47#_c_323_n 0.0259457f $X=2.34 $Y=2.245 $X2=0
+ $Y2=0
cc_137 N_A_59_194#_c_99_n N_A_237_47#_c_314_n 0.012549f $X=2.34 $Y=2.075 $X2=0
+ $Y2=0
cc_138 N_A_59_194#_c_135_p N_B2_M1007_g 0.00590825f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_59_194#_c_99_n N_B2_M1007_g 0.0116798f $X=2.34 $Y=2.075 $X2=0 $Y2=0
cc_140 N_A_59_194#_c_99_n N_B2_M1005_g 9.20219e-19 $X=2.34 $Y=2.075 $X2=0 $Y2=0
cc_141 N_A_59_194#_c_108_n N_B2_M1005_g 2.60415e-19 $X=2.34 $Y=2.245 $X2=0 $Y2=0
cc_142 N_A_59_194#_c_99_n B2 0.0776817f $X=2.34 $Y=2.075 $X2=0 $Y2=0
cc_143 N_A_59_194#_c_99_n N_B2_c_392_n 0.0179832f $X=2.34 $Y=2.075 $X2=0 $Y2=0
cc_144 N_A_59_194#_c_135_p N_B1_c_432_n 9.37141e-19 $X=2.41 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_59_194#_c_99_n N_B1_c_432_n 8.70625e-19 $X=2.34 $Y=2.075 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_59_194#_c_96_n N_X_c_468_n 2.24176e-19 $X=0.605 $Y=1.045 $X2=0 $Y2=0
cc_147 N_A_59_194#_c_97_n N_X_c_468_n 0.00673155f $X=0.445 $Y=1.045 $X2=0 $Y2=0
cc_148 N_A_59_194#_c_95_n X 0.0272167f $X=0.37 $Y=1.93 $X2=0 $Y2=0
cc_149 N_A_59_194#_c_97_n X 0.0063258f $X=0.445 $Y=1.045 $X2=0 $Y2=0
cc_150 N_A_59_194#_M1000_g X 0.00614841f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_151 N_A_59_194#_c_102_n X 0.0263713f $X=1.14 $Y=2.095 $X2=0 $Y2=0
cc_152 N_A_59_194#_c_109_n X 0.0175036f $X=0.495 $Y=2.095 $X2=0 $Y2=0
cc_153 N_A_59_194#_M1003_g X 0.00348303f $X=0.495 $Y=2.77 $X2=0 $Y2=0
cc_154 N_A_59_194#_c_109_n X 0.00335397f $X=0.495 $Y=2.095 $X2=0 $Y2=0
cc_155 N_A_59_194#_M1003_g X 0.00499291f $X=0.495 $Y=2.77 $X2=0 $Y2=0
cc_156 N_A_59_194#_M1003_g N_VPWR_c_496_n 0.00655064f $X=0.495 $Y=2.77 $X2=0
+ $Y2=0
cc_157 N_A_59_194#_c_102_n N_VPWR_c_496_n 0.0306186f $X=1.14 $Y=2.095 $X2=0
+ $Y2=0
cc_158 N_A_59_194#_c_103_n N_VPWR_c_496_n 0.0180907f $X=1.225 $Y=2.88 $X2=0
+ $Y2=0
cc_159 N_A_59_194#_c_105_n N_VPWR_c_496_n 0.0146155f $X=1.31 $Y=2.965 $X2=0
+ $Y2=0
cc_160 N_A_59_194#_c_109_n N_VPWR_c_496_n 0.0032381f $X=0.495 $Y=2.095 $X2=0
+ $Y2=0
cc_161 N_A_59_194#_M1003_g N_VPWR_c_498_n 0.00544103f $X=0.495 $Y=2.77 $X2=0
+ $Y2=0
cc_162 N_A_59_194#_c_104_n N_VPWR_c_499_n 0.0486835f $X=2.185 $Y=2.965 $X2=0
+ $Y2=0
cc_163 N_A_59_194#_c_105_n N_VPWR_c_499_n 0.0105206f $X=1.31 $Y=2.965 $X2=0
+ $Y2=0
cc_164 N_A_59_194#_c_106_n N_VPWR_c_499_n 0.0128088f $X=2.302 $Y=2.88 $X2=0
+ $Y2=0
cc_165 N_A_59_194#_M1011_s N_VPWR_c_495_n 0.00251649f $X=2.165 $Y=2.675 $X2=0
+ $Y2=0
cc_166 N_A_59_194#_M1003_g N_VPWR_c_495_n 0.0120229f $X=0.495 $Y=2.77 $X2=0
+ $Y2=0
cc_167 N_A_59_194#_c_104_n N_VPWR_c_495_n 0.0323925f $X=2.185 $Y=2.965 $X2=0
+ $Y2=0
cc_168 N_A_59_194#_c_105_n N_VPWR_c_495_n 0.00652894f $X=1.31 $Y=2.965 $X2=0
+ $Y2=0
cc_169 N_A_59_194#_c_106_n N_VPWR_c_495_n 0.00901394f $X=2.302 $Y=2.88 $X2=0
+ $Y2=0
cc_170 N_A_59_194#_c_103_n A_223_490# 0.00177857f $X=1.225 $Y=2.88 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_59_194#_c_106_n N_A_516_535#_c_546_n 0.00699485f $X=2.302 $Y=2.88
+ $X2=0 $Y2=0
cc_172 N_A_59_194#_c_106_n N_A_516_535#_c_548_n 0.0146715f $X=2.302 $Y=2.88
+ $X2=0 $Y2=0
cc_173 N_A_59_194#_M1000_g N_VGND_c_572_n 0.00316145f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_174 N_A_59_194#_c_135_p N_VGND_c_575_n 0.0103611f $X=2.41 $Y=0.445 $X2=0
+ $Y2=0
cc_175 N_A_59_194#_M1000_g N_VGND_c_576_n 0.00585385f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_A_59_194#_c_135_p N_VGND_c_578_n 0.0159982f $X=2.41 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_59_194#_M1006_d N_VGND_c_580_n 0.00226211f $X=2.185 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_A_59_194#_M1000_g N_VGND_c_580_n 0.00732527f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_59_194#_c_135_p N_VGND_c_580_n 0.0123335f $X=2.41 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A1_N_M1004_g N_A2_N_M1010_g 0.0549786f $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_181 N_A1_N_c_196_n N_A2_N_M1001_g 0.00805717f $X=1.04 $Y=1.36 $X2=0 $Y2=0
cc_182 N_A1_N_c_197_n N_A2_N_M1001_g 0.0168818f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_183 A1_N N_A2_N_c_255_n 2.13715e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_184 N_A1_N_c_200_n N_A2_N_c_255_n 0.0145504f $X=1.04 $Y=1.525 $X2=0 $Y2=0
cc_185 N_A1_N_M1004_g N_A2_N_c_259_n 0.0145504f $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_186 N_A1_N_c_196_n A2_N 0.00447435f $X=1.04 $Y=1.36 $X2=0 $Y2=0
cc_187 N_A1_N_M1004_g A2_N 0.00122159f $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_188 N_A1_N_c_198_n A2_N 0.00311359f $X=1.075 $Y=0.915 $X2=0 $Y2=0
cc_189 A1_N A2_N 0.0490416f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_190 N_A1_N_c_200_n A2_N 0.00791503f $X=1.04 $Y=1.525 $X2=0 $Y2=0
cc_191 N_A1_N_c_196_n N_A2_N_c_257_n 0.0145504f $X=1.04 $Y=1.36 $X2=0 $Y2=0
cc_192 N_A1_N_c_197_n N_A_237_47#_c_308_n 0.003496f $X=1.075 $Y=0.765 $X2=0
+ $Y2=0
cc_193 N_A1_N_c_196_n N_A_237_47#_c_310_n 6.16991e-19 $X=1.04 $Y=1.36 $X2=0
+ $Y2=0
cc_194 N_A1_N_c_198_n N_A_237_47#_c_310_n 0.00154531f $X=1.075 $Y=0.915 $X2=0
+ $Y2=0
cc_195 A1_N N_A_237_47#_c_310_n 0.0129805f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_196 A1_N N_X_c_468_n 0.00348693f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_197 N_A1_N_M1004_g X 0.00153476f $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_198 A1_N X 0.0698584f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_199 N_A1_N_c_200_n X 2.72214e-19 $X=1.04 $Y=1.525 $X2=0 $Y2=0
cc_200 N_A1_N_M1004_g X 2.26563e-19 $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_201 N_A1_N_M1004_g N_VPWR_c_496_n 0.00803424f $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_202 N_A1_N_M1004_g N_VPWR_c_499_n 0.00495467f $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_203 N_A1_N_M1004_g N_VPWR_c_495_n 0.00503696f $X=1.04 $Y=2.66 $X2=0 $Y2=0
cc_204 N_A1_N_c_197_n N_VGND_c_572_n 0.00174527f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_205 N_A1_N_c_198_n N_VGND_c_572_n 0.00176781f $X=1.075 $Y=0.915 $X2=0 $Y2=0
cc_206 A1_N N_VGND_c_572_n 0.0129121f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_207 N_A1_N_c_197_n N_VGND_c_573_n 0.00585385f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_208 N_A1_N_c_197_n N_VGND_c_580_n 0.010818f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_209 N_A1_N_c_198_n N_VGND_c_580_n 2.68819e-19 $X=1.075 $Y=0.915 $X2=0 $Y2=0
cc_210 A1_N N_VGND_c_580_n 0.0067001f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_211 N_A2_N_M1001_g N_A_237_47#_M1006_g 0.0252209f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_212 N_A2_N_c_257_n N_A_237_47#_M1006_g 0.00192071f $X=1.49 $Y=1.32 $X2=0
+ $Y2=0
cc_213 N_A2_N_M1010_g N_A_237_47#_c_315_n 0.00405672f $X=1.43 $Y=2.66 $X2=0
+ $Y2=0
cc_214 N_A2_N_c_255_n N_A_237_47#_c_307_n 0.0103437f $X=1.49 $Y=1.66 $X2=0 $Y2=0
cc_215 N_A2_N_M1010_g N_A_237_47#_c_320_n 0.00212294f $X=1.43 $Y=2.66 $X2=0
+ $Y2=0
cc_216 N_A2_N_c_259_n N_A_237_47#_c_320_n 0.0103437f $X=1.49 $Y=1.825 $X2=0
+ $Y2=0
cc_217 N_A2_N_M1001_g N_A_237_47#_c_308_n 0.00349423f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A2_N_M1001_g N_A_237_47#_c_309_n 0.0129839f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_219 A2_N N_A_237_47#_c_309_n 0.014678f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A2_N_c_257_n N_A_237_47#_c_309_n 2.64151e-19 $X=1.49 $Y=1.32 $X2=0
+ $Y2=0
cc_221 A2_N N_A_237_47#_c_310_n 0.0251167f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_222 N_A2_N_c_257_n N_A_237_47#_c_310_n 0.00106118f $X=1.49 $Y=1.32 $X2=0
+ $Y2=0
cc_223 N_A2_N_M1010_g N_A_237_47#_c_321_n 0.00471181f $X=1.43 $Y=2.66 $X2=0
+ $Y2=0
cc_224 N_A2_N_c_259_n N_A_237_47#_c_321_n 0.00415876f $X=1.49 $Y=1.825 $X2=0
+ $Y2=0
cc_225 N_A2_N_c_255_n N_A_237_47#_c_311_n 0.0018095f $X=1.49 $Y=1.66 $X2=0 $Y2=0
cc_226 N_A2_N_c_259_n N_A_237_47#_c_312_n 0.0018095f $X=1.49 $Y=1.825 $X2=0
+ $Y2=0
cc_227 A2_N N_A_237_47#_c_313_n 5.82486e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A2_N_c_257_n N_A_237_47#_c_313_n 0.0103437f $X=1.49 $Y=1.32 $X2=0 $Y2=0
cc_229 N_A2_N_M1001_g N_A_237_47#_c_314_n 0.00357277f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_230 A2_N N_A_237_47#_c_314_n 0.0470402f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_231 N_A2_N_c_257_n N_A_237_47#_c_314_n 0.0018095f $X=1.49 $Y=1.32 $X2=0 $Y2=0
cc_232 N_A2_N_M1010_g N_A_237_47#_c_324_n 0.00864466f $X=1.43 $Y=2.66 $X2=0
+ $Y2=0
cc_233 N_A2_N_M1010_g N_VPWR_c_496_n 2.21287e-19 $X=1.43 $Y=2.66 $X2=0 $Y2=0
cc_234 N_A2_N_M1010_g N_VPWR_c_499_n 8.13067e-19 $X=1.43 $Y=2.66 $X2=0 $Y2=0
cc_235 N_A2_N_M1001_g N_VGND_c_573_n 0.00585385f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A2_N_M1001_g N_VGND_c_574_n 0.00406743f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A2_N_M1001_g N_VGND_c_580_n 0.00659198f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_238 N_A_237_47#_M1006_g N_B2_M1007_g 0.0312845f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A_237_47#_c_316_n N_B2_M1005_g 0.0336228f $X=2.43 $Y=2.14 $X2=0 $Y2=0
cc_240 N_A_237_47#_c_320_n N_B2_M1005_g 0.0026426f $X=2.06 $Y=1.905 $X2=0 $Y2=0
cc_241 N_A_237_47#_c_316_n B2 0.00109563f $X=2.43 $Y=2.14 $X2=0 $Y2=0
cc_242 N_A_237_47#_c_316_n N_B2_c_392_n 0.00797592f $X=2.43 $Y=2.14 $X2=0 $Y2=0
cc_243 N_A_237_47#_c_311_n N_B2_c_392_n 5.1372e-19 $X=1.995 $Y=1.395 $X2=0 $Y2=0
cc_244 N_A_237_47#_c_313_n N_B2_c_392_n 0.0308103f $X=2.06 $Y=1.4 $X2=0 $Y2=0
cc_245 N_A_237_47#_M1011_g N_VPWR_c_499_n 0.00585385f $X=2.505 $Y=2.885 $X2=0
+ $Y2=0
cc_246 N_A_237_47#_M1011_g N_VPWR_c_495_n 0.0124078f $X=2.505 $Y=2.885 $X2=0
+ $Y2=0
cc_247 N_A_237_47#_M1011_g N_A_516_535#_c_546_n 7.75802e-19 $X=2.505 $Y=2.885
+ $X2=0 $Y2=0
cc_248 N_A_237_47#_M1011_g N_A_516_535#_c_548_n 0.00151072f $X=2.505 $Y=2.885
+ $X2=0 $Y2=0
cc_249 N_A_237_47#_c_308_n N_VGND_c_573_n 0.0135213f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_250 N_A_237_47#_M1006_g N_VGND_c_574_n 0.00537835f $X=2.11 $Y=0.445 $X2=0
+ $Y2=0
cc_251 N_A_237_47#_c_309_n N_VGND_c_574_n 0.0264043f $X=1.835 $Y=0.877 $X2=0
+ $Y2=0
cc_252 N_A_237_47#_c_313_n N_VGND_c_574_n 2.81358e-19 $X=2.06 $Y=1.4 $X2=0 $Y2=0
cc_253 N_A_237_47#_M1006_g N_VGND_c_578_n 0.0054833f $X=2.11 $Y=0.445 $X2=0
+ $Y2=0
cc_254 N_A_237_47#_M1009_d N_VGND_c_580_n 0.00277345f $X=1.185 $Y=0.235 $X2=0
+ $Y2=0
cc_255 N_A_237_47#_M1006_g N_VGND_c_580_n 0.0102652f $X=2.11 $Y=0.445 $X2=0
+ $Y2=0
cc_256 N_A_237_47#_c_308_n N_VGND_c_580_n 0.0102992f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_257 N_A_237_47#_c_309_n N_VGND_c_580_n 0.0079296f $X=1.835 $Y=0.877 $X2=0
+ $Y2=0
cc_258 N_B2_M1007_g N_B1_c_432_n 0.0420827f $X=2.54 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_259 B2 N_B1_c_433_n 0.012037f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_260 B2 N_B1_c_434_n 0.00773704f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_261 N_B2_c_392_n N_B1_c_434_n 0.00856468f $X=2.845 $Y=1.32 $X2=0 $Y2=0
cc_262 N_B2_M1005_g N_B1_c_436_n 0.0370686f $X=2.935 $Y=2.885 $X2=0 $Y2=0
cc_263 B2 B1 0.115017f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_264 N_B2_c_392_n B1 7.45613e-19 $X=2.845 $Y=1.32 $X2=0 $Y2=0
cc_265 N_B2_M1007_g N_B1_c_438_n 0.00225316f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_266 B2 N_B1_c_438_n 0.0123233f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_267 N_B2_c_392_n N_B1_c_438_n 0.0370686f $X=2.845 $Y=1.32 $X2=0 $Y2=0
cc_268 N_B2_M1005_g N_VPWR_c_497_n 0.0031034f $X=2.935 $Y=2.885 $X2=0 $Y2=0
cc_269 N_B2_M1005_g N_VPWR_c_499_n 0.00440547f $X=2.935 $Y=2.885 $X2=0 $Y2=0
cc_270 N_B2_M1005_g N_VPWR_c_495_n 0.00602924f $X=2.935 $Y=2.885 $X2=0 $Y2=0
cc_271 N_B2_M1005_g N_A_516_535#_c_546_n 0.0012913f $X=2.935 $Y=2.885 $X2=0
+ $Y2=0
cc_272 N_B2_M1005_g N_A_516_535#_c_547_n 0.0122172f $X=2.935 $Y=2.885 $X2=0
+ $Y2=0
cc_273 B2 N_A_516_535#_c_547_n 0.0285595f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_274 B2 N_A_516_535#_c_548_n 0.00497163f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_275 N_B2_c_392_n N_A_516_535#_c_548_n 0.00547084f $X=2.845 $Y=1.32 $X2=0
+ $Y2=0
cc_276 N_B2_M1007_g N_VGND_c_575_n 0.00223131f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_277 B2 N_VGND_c_575_n 0.020051f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_278 N_B2_M1007_g N_VGND_c_578_n 0.00540919f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_279 N_B2_M1007_g N_VGND_c_580_n 0.00980721f $X=2.54 $Y=0.445 $X2=0 $Y2=0
cc_280 B2 N_VGND_c_580_n 0.00913252f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_281 N_B1_M1002_g N_VPWR_c_497_n 0.0031336f $X=3.365 $Y=2.885 $X2=0 $Y2=0
cc_282 N_B1_M1002_g N_VPWR_c_500_n 0.00440547f $X=3.365 $Y=2.885 $X2=0 $Y2=0
cc_283 N_B1_M1002_g N_VPWR_c_495_n 0.00699263f $X=3.365 $Y=2.885 $X2=0 $Y2=0
cc_284 N_B1_M1002_g N_A_516_535#_c_547_n 0.0176924f $X=3.365 $Y=2.885 $X2=0
+ $Y2=0
cc_285 B1 N_A_516_535#_c_547_n 0.0247285f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_286 N_B1_M1002_g N_A_516_535#_c_549_n 0.00300843f $X=3.365 $Y=2.885 $X2=0
+ $Y2=0
cc_287 N_B1_c_432_n N_VGND_c_575_n 0.0125866f $X=2.93 $Y=0.765 $X2=0 $Y2=0
cc_288 N_B1_c_433_n N_VGND_c_575_n 0.00475697f $X=3.29 $Y=0.84 $X2=0 $Y2=0
cc_289 B1 N_VGND_c_575_n 0.0169364f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_290 N_B1_c_432_n N_VGND_c_578_n 0.00486043f $X=2.93 $Y=0.765 $X2=0 $Y2=0
cc_291 N_B1_c_433_n N_VGND_c_579_n 0.00385916f $X=3.29 $Y=0.84 $X2=0 $Y2=0
cc_292 B1 N_VGND_c_579_n 0.0123662f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_293 N_B1_c_432_n N_VGND_c_580_n 0.00441005f $X=2.93 $Y=0.765 $X2=0 $Y2=0
cc_294 N_B1_c_433_n N_VGND_c_580_n 0.00436486f $X=3.29 $Y=0.84 $X2=0 $Y2=0
cc_295 B1 N_VGND_c_580_n 0.011921f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_296 X N_VPWR_c_496_n 0.0252877f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_297 X N_VPWR_c_498_n 0.0231836f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_298 N_X_M1003_s N_VPWR_c_495_n 0.00213729f $X=0.155 $Y=2.45 $X2=0 $Y2=0
cc_299 X N_VPWR_c_495_n 0.0137294f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_300 N_X_c_468_n N_VGND_c_576_n 0.0281909f $X=0.465 $Y=0.445 $X2=0 $Y2=0
cc_301 N_X_M1000_s N_VGND_c_580_n 0.00247877f $X=0.31 $Y=0.235 $X2=0 $Y2=0
cc_302 N_X_c_468_n N_VGND_c_580_n 0.0191928f $X=0.465 $Y=0.445 $X2=0 $Y2=0
cc_303 N_VPWR_c_495_n N_A_516_535#_M1011_d 0.00281679f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_304 N_VPWR_c_495_n N_A_516_535#_M1002_d 0.00223845f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_499_n N_A_516_535#_c_546_n 0.0120755f $X=3.02 $Y=3.33 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_495_n N_A_516_535#_c_546_n 0.00893098f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_497_n N_A_516_535#_c_547_n 0.0166679f $X=3.15 $Y=2.92 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_499_n N_A_516_535#_c_547_n 0.00256486f $X=3.02 $Y=3.33 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_500_n N_A_516_535#_c_547_n 0.00219893f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_495_n N_A_516_535#_c_547_n 0.00896087f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_500_n N_A_516_535#_c_549_n 0.0162027f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_312 N_VPWR_c_495_n N_A_516_535#_c_549_n 0.0110391f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VGND_c_580_n A_523_47# 0.00754654f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
