* File: sky130_fd_sc_lp__dlrtn_2.pxi.spice
* Created: Wed Sep  2 09:46:57 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTN_2%D N_D_M1013_g N_D_M1003_g N_D_c_150_n N_D_c_151_n
+ N_D_c_152_n D D D N_D_c_154_n PM_SKY130_FD_SC_LP__DLRTN_2%D
x_PM_SKY130_FD_SC_LP__DLRTN_2%GATE_N N_GATE_N_M1004_g N_GATE_N_M1005_g
+ N_GATE_N_c_190_n N_GATE_N_c_191_n N_GATE_N_c_192_n GATE_N GATE_N GATE_N
+ N_GATE_N_c_194_n PM_SKY130_FD_SC_LP__DLRTN_2%GATE_N
x_PM_SKY130_FD_SC_LP__DLRTN_2%A_31_464# N_A_31_464#_M1003_s N_A_31_464#_M1013_s
+ N_A_31_464#_M1019_g N_A_31_464#_M1007_g N_A_31_464#_c_244_n
+ N_A_31_464#_c_245_n N_A_31_464#_c_239_n N_A_31_464#_c_247_n
+ N_A_31_464#_c_248_n N_A_31_464#_c_249_n N_A_31_464#_c_250_n
+ N_A_31_464#_c_251_n N_A_31_464#_c_252_n N_A_31_464#_c_279_p
+ N_A_31_464#_c_253_n N_A_31_464#_c_240_n N_A_31_464#_c_241_n
+ N_A_31_464#_c_242_n N_A_31_464#_c_256_n PM_SKY130_FD_SC_LP__DLRTN_2%A_31_464#
x_PM_SKY130_FD_SC_LP__DLRTN_2%A_372_397# N_A_372_397#_M1018_s
+ N_A_372_397#_M1000_s N_A_372_397#_M1009_g N_A_372_397#_M1016_g
+ N_A_372_397#_c_352_n N_A_372_397#_c_353_n N_A_372_397#_c_354_n
+ N_A_372_397#_c_355_n N_A_372_397#_c_356_n N_A_372_397#_c_357_n
+ N_A_372_397#_c_358_n N_A_372_397#_c_359_n N_A_372_397#_c_364_n
+ N_A_372_397#_c_365_n N_A_372_397#_c_360_n N_A_372_397#_c_361_n
+ PM_SKY130_FD_SC_LP__DLRTN_2%A_372_397#
x_PM_SKY130_FD_SC_LP__DLRTN_2%A_221_70# N_A_221_70#_M1004_d N_A_221_70#_M1005_d
+ N_A_221_70#_c_459_n N_A_221_70#_c_460_n N_A_221_70#_c_461_n
+ N_A_221_70#_c_462_n N_A_221_70#_c_473_n N_A_221_70#_c_474_n
+ N_A_221_70#_c_463_n N_A_221_70#_M1018_g N_A_221_70#_M1000_g
+ N_A_221_70#_c_464_n N_A_221_70#_M1015_g N_A_221_70#_c_466_n
+ N_A_221_70#_M1012_g N_A_221_70#_c_467_n N_A_221_70#_c_468_n
+ N_A_221_70#_c_469_n N_A_221_70#_c_470_n N_A_221_70#_c_471_n
+ N_A_221_70#_c_480_n N_A_221_70#_c_481_n N_A_221_70#_c_472_n
+ N_A_221_70#_c_482_n PM_SKY130_FD_SC_LP__DLRTN_2%A_221_70#
x_PM_SKY130_FD_SC_LP__DLRTN_2%A_776_99# N_A_776_99#_M1017_s N_A_776_99#_M1002_d
+ N_A_776_99#_c_589_n N_A_776_99#_M1021_g N_A_776_99#_M1014_g
+ N_A_776_99#_M1001_g N_A_776_99#_M1008_g N_A_776_99#_M1006_g
+ N_A_776_99#_M1020_g N_A_776_99#_c_594_n N_A_776_99#_c_604_n
+ N_A_776_99#_c_595_n N_A_776_99#_c_596_n N_A_776_99#_c_647_p
+ N_A_776_99#_c_686_p N_A_776_99#_c_606_n N_A_776_99#_c_597_n
+ N_A_776_99#_c_598_n N_A_776_99#_c_608_n N_A_776_99#_c_609_n
+ N_A_776_99#_c_599_n N_A_776_99#_c_610_n N_A_776_99#_c_650_p
+ N_A_776_99#_c_600_n PM_SKY130_FD_SC_LP__DLRTN_2%A_776_99#
x_PM_SKY130_FD_SC_LP__DLRTN_2%A_626_125# N_A_626_125#_M1015_d
+ N_A_626_125#_M1009_d N_A_626_125#_M1017_g N_A_626_125#_M1002_g
+ N_A_626_125#_c_725_n N_A_626_125#_c_726_n N_A_626_125#_c_738_n
+ N_A_626_125#_c_727_n N_A_626_125#_c_728_n N_A_626_125#_c_731_n
+ N_A_626_125#_c_732_n N_A_626_125#_c_729_n
+ PM_SKY130_FD_SC_LP__DLRTN_2%A_626_125#
x_PM_SKY130_FD_SC_LP__DLRTN_2%RESET_B N_RESET_B_M1011_g N_RESET_B_M1010_g
+ N_RESET_B_c_826_n N_RESET_B_c_817_n N_RESET_B_c_818_n RESET_B
+ N_RESET_B_c_819_n PM_SKY130_FD_SC_LP__DLRTN_2%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTN_2%VPWR N_VPWR_M1013_d N_VPWR_M1000_d N_VPWR_M1014_d
+ N_VPWR_M1010_d N_VPWR_M1020_s N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_865_n
+ N_VPWR_c_866_n N_VPWR_c_867_n N_VPWR_c_868_n N_VPWR_c_869_n N_VPWR_c_911_n
+ VPWR N_VPWR_c_870_n N_VPWR_c_871_n N_VPWR_c_872_n N_VPWR_c_873_n
+ N_VPWR_c_874_n N_VPWR_c_875_n N_VPWR_c_876_n N_VPWR_c_877_n N_VPWR_c_878_n
+ N_VPWR_c_862_n PM_SKY130_FD_SC_LP__DLRTN_2%VPWR
x_PM_SKY130_FD_SC_LP__DLRTN_2%Q N_Q_M1001_d N_Q_M1008_d Q Q Q Q Q N_Q_c_965_n
+ PM_SKY130_FD_SC_LP__DLRTN_2%Q
x_PM_SKY130_FD_SC_LP__DLRTN_2%VGND N_VGND_M1003_d N_VGND_M1018_d N_VGND_M1021_d
+ N_VGND_M1011_d N_VGND_M1006_s N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n
+ N_VGND_c_987_n N_VGND_c_988_n N_VGND_c_989_n N_VGND_c_990_n VGND
+ N_VGND_c_991_n N_VGND_c_992_n N_VGND_c_993_n N_VGND_c_994_n N_VGND_c_995_n
+ N_VGND_c_996_n N_VGND_c_997_n N_VGND_c_998_n PM_SKY130_FD_SC_LP__DLRTN_2%VGND
cc_1 VNB N_D_M1013_g 0.00611532f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_2 VNB N_D_c_150_n 0.0216291f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.88
cc_3 VNB N_D_c_151_n 0.023176f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_4 VNB N_D_c_152_n 0.01653f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.55
cc_5 VNB D 0.00749522f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_D_c_154_n 0.0163048f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_7 VNB N_GATE_N_M1005_g 0.00504793f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.56
cc_8 VNB N_GATE_N_c_190_n 0.0196332f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.88
cc_9 VNB N_GATE_N_c_191_n 0.02206f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_10 VNB N_GATE_N_c_192_n 0.0157532f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.55
cc_11 VNB GATE_N 0.0076926f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_12 VNB N_GATE_N_c_194_n 0.0168341f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_13 VNB N_A_31_464#_M1019_g 0.0333397f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.88
cc_14 VNB N_A_31_464#_c_239_n 0.0457063f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_15 VNB N_A_31_464#_c_240_n 0.00183416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_31_464#_c_241_n 0.0164908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_31_464#_c_242_n 0.013225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_372_397#_c_352_n 0.00590329f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_19 VNB N_A_372_397#_c_353_n 0.0135649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_372_397#_c_354_n 0.00179308f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_21 VNB N_A_372_397#_c_355_n 0.00228326f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_22 VNB N_A_372_397#_c_356_n 0.00638651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_372_397#_c_357_n 0.0400066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_372_397#_c_358_n 0.00738366f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.295
cc_25 VNB N_A_372_397#_c_359_n 0.00258241f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.665
cc_26 VNB N_A_372_397#_c_360_n 0.00651305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_372_397#_c_361_n 0.0151577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_221_70#_c_459_n 0.053657f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_29 VNB N_A_221_70#_c_460_n 0.0918944f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.88
cc_30 VNB N_A_221_70#_c_461_n 0.0122674f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_31 VNB N_A_221_70#_c_462_n 0.0252395f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.55
cc_32 VNB N_A_221_70#_c_463_n 0.0148465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_221_70#_c_464_n 0.0408489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_221_70#_M1015_g 0.0241772f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.295
cc_35 VNB N_A_221_70#_c_466_n 0.0229519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_221_70#_c_467_n 0.0120692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_221_70#_c_468_n 0.0146449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_221_70#_c_469_n 0.00252237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_221_70#_c_470_n 0.00218799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_221_70#_c_471_n 0.0207071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_221_70#_c_472_n 0.00894616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_776_99#_c_589_n 0.0193714f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.56
cc_43 VNB N_A_776_99#_M1001_g 0.0227123f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_44 VNB N_A_776_99#_M1008_g 0.00155732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_776_99#_M1006_g 0.0295969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_776_99#_M1020_g 0.00157373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_776_99#_c_594_n 0.0205769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_776_99#_c_595_n 0.0078774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_776_99#_c_596_n 0.00352708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_776_99#_c_597_n 0.00394259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_776_99#_c_598_n 0.0784787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_776_99#_c_599_n 0.00605682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_776_99#_c_600_n 0.0187537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_626_125#_M1017_g 0.0245906f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.88
cc_55 VNB N_A_626_125#_M1002_g 0.00203294f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_56 VNB N_A_626_125#_c_725_n 0.0421004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_626_125#_c_726_n 0.00893659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_626_125#_c_727_n 0.00430502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_626_125#_c_728_n 0.0203943f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.665
cc_60 VNB N_A_626_125#_c_729_n 9.63934e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_M1010_g 0.00770343f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.56
cc_62 VNB N_RESET_B_c_817_n 0.00199476f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_63 VNB N_RESET_B_c_818_n 0.0326051f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.55
cc_64 VNB N_RESET_B_c_819_n 0.0162494f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.925
cc_65 VNB N_VPWR_c_862_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_965_n 0.00441612f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_67 VNB N_VGND_c_984_n 0.0082898f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.045
cc_68 VNB N_VGND_c_985_n 0.00749495f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.045
cc_69 VNB N_VGND_c_986_n 0.0336253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_987_n 0.0171797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_988_n 0.00500655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_989_n 0.0106846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_990_n 0.0380491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_991_n 0.0373883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_992_n 0.0275949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_993_n 0.016026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_994_n 0.0260672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_995_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_996_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_997_n 0.00631736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_998_n 0.357085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VPB N_D_M1013_g 0.0586192f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.64
cc_83 VPB D 0.00353065f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_84 VPB N_GATE_N_M1005_g 0.0551932f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=0.56
cc_85 VPB GATE_N 0.00429085f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_86 VPB N_A_31_464#_M1007_g 0.0205247f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_87 VPB N_A_31_464#_c_244_n 0.0246762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_31_464#_c_245_n 0.0163815f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.045
cc_89 VPB N_A_31_464#_c_239_n 0.0144429f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.045
cc_90 VPB N_A_31_464#_c_247_n 0.0368503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_31_464#_c_248_n 0.0166753f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.295
cc_92 VPB N_A_31_464#_c_249_n 0.00173063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_31_464#_c_250_n 0.0142295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_31_464#_c_251_n 0.00125455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_31_464#_c_252_n 0.00262807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_31_464#_c_253_n 0.00197871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_31_464#_c_240_n 0.0017827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_31_464#_c_241_n 0.00209066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_31_464#_c_256_n 0.012132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_372_397#_M1009_g 0.0230157f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.88
cc_101 VPB N_A_372_397#_c_359_n 0.00382031f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.665
cc_102 VPB N_A_372_397#_c_364_n 0.0313281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_372_397#_c_365_n 0.00590201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_372_397#_c_360_n 0.00321103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_221_70#_c_473_n 0.0325233f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_106 VPB N_A_221_70#_c_474_n 0.0178793f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_107 VPB N_A_221_70#_M1000_g 0.0462109f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.045
cc_108 VPB N_A_221_70#_c_464_n 0.00179984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_221_70#_c_466_n 0.0106645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_221_70#_M1012_g 0.0454682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_221_70#_c_471_n 8.85307e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_221_70#_c_480_n 0.0103426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_221_70#_c_481_n 0.0113823f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_221_70#_c_482_n 0.00588699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_776_99#_M1014_g 0.0222674f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_116 VPB N_A_776_99#_M1008_g 0.0203026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_776_99#_M1020_g 0.0222114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_776_99#_c_604_n 0.00676278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_776_99#_c_596_n 6.14258e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_776_99#_c_606_n 0.00752299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_776_99#_c_597_n 0.0260969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_776_99#_c_608_n 0.00381421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_776_99#_c_609_n 0.0356509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_776_99#_c_610_n 0.00739675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_776_99#_c_600_n 0.011748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_626_125#_M1002_g 0.0223538f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_127 VPB N_A_626_125#_c_731_n 0.00501268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_626_125#_c_732_n 0.00518895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_RESET_B_M1010_g 0.0193656f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=0.56
cc_130 VPB N_VPWR_c_863_n 0.0112691f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.045
cc_131 VPB N_VPWR_c_864_n 0.00853103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_865_n 0.0116242f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.665
cc_133 VPB N_VPWR_c_866_n 0.00353629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_867_n 3.16188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_868_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_869_n 0.0199138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_870_n 0.0183556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_871_n 0.0413059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_872_n 0.0406504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_873_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_874_n 0.0153449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_875_n 0.00430193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_876_n 0.00632006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_877_n 0.0123215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_878_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_862_n 0.0905415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_Q_c_965_n 0.00283085f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.045
cc_148 N_D_M1013_g N_GATE_N_M1005_g 0.0221151f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_149 D N_GATE_N_M1005_g 8.01422e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_150 N_D_c_150_n N_GATE_N_c_190_n 0.0131786f $X=0.55 $Y=0.88 $X2=0 $Y2=0
cc_151 D N_GATE_N_c_190_n 2.59881e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_152 N_D_c_151_n N_GATE_N_c_191_n 0.0137828f $X=0.55 $Y=1.385 $X2=0 $Y2=0
cc_153 N_D_c_152_n N_GATE_N_c_192_n 0.0137828f $X=0.55 $Y=1.55 $X2=0 $Y2=0
cc_154 N_D_M1013_g GATE_N 5.40026e-19 $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_155 D GATE_N 0.0760295f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_156 N_D_c_154_n GATE_N 5.8438e-19 $X=0.55 $Y=1.045 $X2=0 $Y2=0
cc_157 D N_GATE_N_c_194_n 0.00448642f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_158 N_D_c_154_n N_GATE_N_c_194_n 0.0137828f $X=0.55 $Y=1.045 $X2=0 $Y2=0
cc_159 N_D_M1013_g N_A_31_464#_c_239_n 0.0108171f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_160 N_D_c_150_n N_A_31_464#_c_239_n 0.00430388f $X=0.55 $Y=0.88 $X2=0 $Y2=0
cc_161 D N_A_31_464#_c_239_n 0.069043f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_162 N_D_c_154_n N_A_31_464#_c_239_n 0.0163648f $X=0.55 $Y=1.045 $X2=0 $Y2=0
cc_163 N_D_M1013_g N_A_31_464#_c_247_n 0.00575074f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_164 N_D_M1013_g N_A_31_464#_c_248_n 0.0189186f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_165 N_D_c_152_n N_A_31_464#_c_248_n 8.89382e-19 $X=0.55 $Y=1.55 $X2=0 $Y2=0
cc_166 D N_A_31_464#_c_248_n 0.0302195f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_167 N_D_M1013_g N_A_31_464#_c_249_n 0.00206124f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_168 N_D_c_150_n N_A_31_464#_c_242_n 0.00239439f $X=0.55 $Y=0.88 $X2=0 $Y2=0
cc_169 D N_A_31_464#_c_242_n 0.00304282f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_170 N_D_c_154_n N_A_31_464#_c_242_n 0.00361721f $X=0.55 $Y=1.045 $X2=0 $Y2=0
cc_171 N_D_c_152_n N_A_31_464#_c_256_n 9.30767e-19 $X=0.55 $Y=1.55 $X2=0 $Y2=0
cc_172 N_D_M1013_g N_VPWR_c_863_n 0.00390064f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_173 N_D_M1013_g N_VPWR_c_870_n 0.00461464f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_174 N_D_M1013_g N_VPWR_c_862_n 0.00912986f $X=0.495 $Y=2.64 $X2=0 $Y2=0
cc_175 N_D_c_150_n N_VGND_c_984_n 0.00331625f $X=0.55 $Y=0.88 $X2=0 $Y2=0
cc_176 D N_VGND_c_984_n 0.0105289f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_177 N_D_c_150_n N_VGND_c_994_n 0.00472388f $X=0.55 $Y=0.88 $X2=0 $Y2=0
cc_178 N_D_c_150_n N_VGND_c_998_n 0.00509226f $X=0.55 $Y=0.88 $X2=0 $Y2=0
cc_179 D N_VGND_c_998_n 0.00622581f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_180 N_GATE_N_M1005_g N_A_31_464#_c_248_n 0.0063468f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_181 N_GATE_N_c_192_n N_A_31_464#_c_248_n 0.00320349f $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_182 GATE_N N_A_31_464#_c_248_n 0.0126619f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_183 N_GATE_N_M1005_g N_A_31_464#_c_249_n 0.0186388f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_184 N_GATE_N_M1005_g N_A_31_464#_c_250_n 0.0116719f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_185 N_GATE_N_M1005_g N_A_31_464#_c_251_n 0.00300044f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_186 N_GATE_N_M1005_g N_A_31_464#_c_252_n 0.00238622f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_187 N_GATE_N_c_194_n N_A_221_70#_c_459_n 0.00635393f $X=1.09 $Y=1.045 $X2=0
+ $Y2=0
cc_188 N_GATE_N_c_190_n N_A_221_70#_c_461_n 0.00780985f $X=1.09 $Y=0.88 $X2=0
+ $Y2=0
cc_189 N_GATE_N_M1005_g N_A_221_70#_c_474_n 0.0122097f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_190 N_GATE_N_c_191_n N_A_221_70#_c_467_n 0.0122097f $X=1.09 $Y=1.385 $X2=0
+ $Y2=0
cc_191 GATE_N N_A_221_70#_c_467_n 0.00195322f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_192 GATE_N N_A_221_70#_c_468_n 0.0134801f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_193 N_GATE_N_c_194_n N_A_221_70#_c_468_n 8.28126e-19 $X=1.09 $Y=1.045 $X2=0
+ $Y2=0
cc_194 N_GATE_N_c_191_n N_A_221_70#_c_469_n 6.95221e-19 $X=1.09 $Y=1.385 $X2=0
+ $Y2=0
cc_195 N_GATE_N_c_192_n N_A_221_70#_c_470_n 6.95221e-19 $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_196 N_GATE_N_c_192_n N_A_221_70#_c_471_n 0.0122097f $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_197 N_GATE_N_M1005_g N_A_221_70#_c_481_n 0.00142509f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_198 N_GATE_N_c_190_n N_A_221_70#_c_472_n 0.0031016f $X=1.09 $Y=0.88 $X2=0
+ $Y2=0
cc_199 GATE_N N_A_221_70#_c_472_n 0.0764322f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_200 N_GATE_N_c_194_n N_A_221_70#_c_472_n 6.95221e-19 $X=1.09 $Y=1.045 $X2=0
+ $Y2=0
cc_201 N_GATE_N_M1005_g N_A_221_70#_c_482_n 0.0125797f $X=1.18 $Y=2.64 $X2=0
+ $Y2=0
cc_202 N_GATE_N_M1005_g N_VPWR_c_863_n 0.00421734f $X=1.18 $Y=2.64 $X2=0 $Y2=0
cc_203 N_GATE_N_M1005_g N_VPWR_c_871_n 0.00291612f $X=1.18 $Y=2.64 $X2=0 $Y2=0
cc_204 N_GATE_N_M1005_g N_VPWR_c_862_n 0.00366095f $X=1.18 $Y=2.64 $X2=0 $Y2=0
cc_205 N_GATE_N_c_190_n N_VGND_c_984_n 0.00321079f $X=1.09 $Y=0.88 $X2=0 $Y2=0
cc_206 N_GATE_N_c_190_n N_VGND_c_991_n 0.00478016f $X=1.09 $Y=0.88 $X2=0 $Y2=0
cc_207 N_GATE_N_c_190_n N_VGND_c_998_n 0.00653901f $X=1.09 $Y=0.88 $X2=0 $Y2=0
cc_208 GATE_N N_VGND_c_998_n 0.00367754f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_209 N_GATE_N_c_194_n N_VGND_c_998_n 3.9536e-19 $X=1.09 $Y=1.045 $X2=0 $Y2=0
cc_210 N_A_31_464#_c_250_n N_A_372_397#_M1000_s 0.00486566f $X=1.815 $Y=2.895
+ $X2=0 $Y2=0
cc_211 N_A_31_464#_c_252_n N_A_372_397#_M1000_s 0.00406698f $X=1.9 $Y=2.81 $X2=0
+ $Y2=0
cc_212 N_A_31_464#_c_279_p N_A_372_397#_M1000_s 0.00574821f $X=2.58 $Y=2.51
+ $X2=0 $Y2=0
cc_213 N_A_31_464#_c_253_n N_A_372_397#_M1000_s 0.00243323f $X=1.985 $Y=2.51
+ $X2=0 $Y2=0
cc_214 N_A_31_464#_c_245_n N_A_372_397#_M1009_g 0.0376202f $X=2.745 $Y=2.185
+ $X2=0 $Y2=0
cc_215 N_A_31_464#_c_279_p N_A_372_397#_M1009_g 5.74605e-19 $X=2.58 $Y=2.51
+ $X2=0 $Y2=0
cc_216 N_A_31_464#_M1019_g N_A_372_397#_c_353_n 0.0138859f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_217 N_A_31_464#_c_240_n N_A_372_397#_c_353_n 0.0209609f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_218 N_A_31_464#_c_241_n N_A_372_397#_c_353_n 0.00117149f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_219 N_A_31_464#_M1019_g N_A_372_397#_c_354_n 0.00313447f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_220 N_A_31_464#_M1019_g N_A_372_397#_c_359_n 0.00129909f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_221 N_A_31_464#_c_244_n N_A_372_397#_c_359_n 0.00113602f $X=2.745 $Y=2.02
+ $X2=0 $Y2=0
cc_222 N_A_31_464#_c_240_n N_A_372_397#_c_359_n 0.0441079f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_223 N_A_31_464#_c_241_n N_A_372_397#_c_359_n 0.00538706f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_224 N_A_31_464#_c_244_n N_A_372_397#_c_364_n 0.0376202f $X=2.745 $Y=2.02
+ $X2=0 $Y2=0
cc_225 N_A_31_464#_c_240_n N_A_372_397#_c_364_n 0.00199931f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_226 N_A_31_464#_c_279_p N_A_372_397#_c_365_n 0.0133754f $X=2.58 $Y=2.51 $X2=0
+ $Y2=0
cc_227 N_A_31_464#_c_253_n N_A_372_397#_c_365_n 0.0140669f $X=1.985 $Y=2.51
+ $X2=0 $Y2=0
cc_228 N_A_31_464#_M1019_g N_A_372_397#_c_360_n 0.00545049f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_229 N_A_31_464#_c_240_n N_A_372_397#_c_360_n 0.028313f $X=2.745 $Y=1.68 $X2=0
+ $Y2=0
cc_230 N_A_31_464#_c_241_n N_A_372_397#_c_360_n 0.00336889f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_231 N_A_31_464#_c_250_n N_A_221_70#_M1005_d 0.00361268f $X=1.815 $Y=2.895
+ $X2=0 $Y2=0
cc_232 N_A_31_464#_M1019_g N_A_221_70#_c_460_n 0.00894529f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_233 N_A_31_464#_c_279_p N_A_221_70#_c_473_n 0.00139819f $X=2.58 $Y=2.51 $X2=0
+ $Y2=0
cc_234 N_A_31_464#_c_240_n N_A_221_70#_c_473_n 0.00197171f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_235 N_A_31_464#_c_241_n N_A_221_70#_c_473_n 0.015797f $X=2.745 $Y=1.68 $X2=0
+ $Y2=0
cc_236 N_A_31_464#_c_253_n N_A_221_70#_c_474_n 3.28957e-19 $X=1.985 $Y=2.51
+ $X2=0 $Y2=0
cc_237 N_A_31_464#_M1019_g N_A_221_70#_c_463_n 0.0187215f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_238 N_A_31_464#_M1007_g N_A_221_70#_M1000_g 0.0178656f $X=2.835 $Y=2.685
+ $X2=0 $Y2=0
cc_239 N_A_31_464#_c_244_n N_A_221_70#_M1000_g 0.015797f $X=2.745 $Y=2.02 $X2=0
+ $Y2=0
cc_240 N_A_31_464#_c_250_n N_A_221_70#_M1000_g 0.00369802f $X=1.815 $Y=2.895
+ $X2=0 $Y2=0
cc_241 N_A_31_464#_c_252_n N_A_221_70#_M1000_g 0.00630929f $X=1.9 $Y=2.81 $X2=0
+ $Y2=0
cc_242 N_A_31_464#_c_279_p N_A_221_70#_M1000_g 0.0189f $X=2.58 $Y=2.51 $X2=0
+ $Y2=0
cc_243 N_A_31_464#_c_240_n N_A_221_70#_M1000_g 0.00464023f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_244 N_A_31_464#_M1019_g N_A_221_70#_c_464_n 0.00744075f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_245 N_A_31_464#_c_240_n N_A_221_70#_c_464_n 3.20169e-19 $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_246 N_A_31_464#_c_241_n N_A_221_70#_c_464_n 0.00855568f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_247 N_A_31_464#_M1019_g N_A_221_70#_M1015_g 0.0482266f $X=2.695 $Y=0.835
+ $X2=0 $Y2=0
cc_248 N_A_31_464#_c_248_n N_A_221_70#_c_480_n 0.00843867f $X=0.975 $Y=2.045
+ $X2=0 $Y2=0
cc_249 N_A_31_464#_c_249_n N_A_221_70#_c_480_n 0.00757517f $X=1.06 $Y=2.81 $X2=0
+ $Y2=0
cc_250 N_A_31_464#_c_249_n N_A_221_70#_c_481_n 0.0232469f $X=1.06 $Y=2.81 $X2=0
+ $Y2=0
cc_251 N_A_31_464#_c_250_n N_A_221_70#_c_481_n 0.0218465f $X=1.815 $Y=2.895
+ $X2=0 $Y2=0
cc_252 N_A_31_464#_c_252_n N_A_221_70#_c_481_n 0.00255157f $X=1.9 $Y=2.81 $X2=0
+ $Y2=0
cc_253 N_A_31_464#_c_253_n N_A_221_70#_c_481_n 0.0144401f $X=1.985 $Y=2.51 $X2=0
+ $Y2=0
cc_254 N_A_31_464#_M1007_g N_A_626_125#_c_731_n 0.00178891f $X=2.835 $Y=2.685
+ $X2=0 $Y2=0
cc_255 N_A_31_464#_c_279_p N_A_626_125#_c_731_n 0.00767514f $X=2.58 $Y=2.51
+ $X2=0 $Y2=0
cc_256 N_A_31_464#_c_240_n N_A_626_125#_c_731_n 0.00210951f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_257 N_A_31_464#_M1007_g N_A_626_125#_c_732_n 3.87407e-19 $X=2.835 $Y=2.685
+ $X2=0 $Y2=0
cc_258 N_A_31_464#_c_240_n N_A_626_125#_c_732_n 0.00459713f $X=2.745 $Y=1.68
+ $X2=0 $Y2=0
cc_259 N_A_31_464#_c_249_n N_VPWR_M1013_d 0.00448184f $X=1.06 $Y=2.81 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_31_464#_c_251_n N_VPWR_M1013_d 0.00143095f $X=1.145 $Y=2.895
+ $X2=-0.19 $Y2=-0.245
cc_261 N_A_31_464#_c_279_p N_VPWR_M1000_d 0.00896492f $X=2.58 $Y=2.51 $X2=0
+ $Y2=0
cc_262 N_A_31_464#_c_240_n N_VPWR_M1000_d 7.62831e-19 $X=2.745 $Y=1.68 $X2=0
+ $Y2=0
cc_263 N_A_31_464#_c_247_n N_VPWR_c_863_n 0.00224457f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_31_464#_c_248_n N_VPWR_c_863_n 0.0188347f $X=0.975 $Y=2.045 $X2=0
+ $Y2=0
cc_265 N_A_31_464#_c_249_n N_VPWR_c_863_n 0.0378558f $X=1.06 $Y=2.81 $X2=0 $Y2=0
cc_266 N_A_31_464#_c_251_n N_VPWR_c_863_n 0.0141604f $X=1.145 $Y=2.895 $X2=0
+ $Y2=0
cc_267 N_A_31_464#_M1007_g N_VPWR_c_864_n 0.00340614f $X=2.835 $Y=2.685 $X2=0
+ $Y2=0
cc_268 N_A_31_464#_c_245_n N_VPWR_c_864_n 4.61086e-19 $X=2.745 $Y=2.185 $X2=0
+ $Y2=0
cc_269 N_A_31_464#_c_279_p N_VPWR_c_864_n 0.0225799f $X=2.58 $Y=2.51 $X2=0 $Y2=0
cc_270 N_A_31_464#_c_247_n N_VPWR_c_870_n 0.0125692f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_31_464#_c_250_n N_VPWR_c_871_n 0.0340589f $X=1.815 $Y=2.895 $X2=0
+ $Y2=0
cc_272 N_A_31_464#_c_251_n N_VPWR_c_871_n 0.00746599f $X=1.145 $Y=2.895 $X2=0
+ $Y2=0
cc_273 N_A_31_464#_c_279_p N_VPWR_c_871_n 0.00512613f $X=2.58 $Y=2.51 $X2=0
+ $Y2=0
cc_274 N_A_31_464#_M1007_g N_VPWR_c_872_n 0.00367486f $X=2.835 $Y=2.685 $X2=0
+ $Y2=0
cc_275 N_A_31_464#_c_279_p N_VPWR_c_872_n 0.00237568f $X=2.58 $Y=2.51 $X2=0
+ $Y2=0
cc_276 N_A_31_464#_M1007_g N_VPWR_c_862_n 0.00508165f $X=2.835 $Y=2.685 $X2=0
+ $Y2=0
cc_277 N_A_31_464#_c_247_n N_VPWR_c_862_n 0.0107561f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_A_31_464#_c_250_n N_VPWR_c_862_n 0.0293944f $X=1.815 $Y=2.895 $X2=0
+ $Y2=0
cc_279 N_A_31_464#_c_251_n N_VPWR_c_862_n 0.00608573f $X=1.145 $Y=2.895 $X2=0
+ $Y2=0
cc_280 N_A_31_464#_c_279_p N_VPWR_c_862_n 0.0159015f $X=2.58 $Y=2.51 $X2=0 $Y2=0
cc_281 N_A_31_464#_M1019_g N_VGND_c_985_n 0.00683104f $X=2.695 $Y=0.835 $X2=0
+ $Y2=0
cc_282 N_A_31_464#_c_242_n N_VGND_c_994_n 0.0135109f $X=0.365 $Y=0.56 $X2=0
+ $Y2=0
cc_283 N_A_31_464#_M1019_g N_VGND_c_998_n 7.97988e-19 $X=2.695 $Y=0.835 $X2=0
+ $Y2=0
cc_284 N_A_31_464#_c_242_n N_VGND_c_998_n 0.0143973f $X=0.365 $Y=0.56 $X2=0
+ $Y2=0
cc_285 N_A_372_397#_c_352_n N_A_221_70#_c_459_n 0.00374508f $X=2.037 $Y=1.295
+ $X2=0 $Y2=0
cc_286 N_A_372_397#_c_352_n N_A_221_70#_c_460_n 0.00425784f $X=2.037 $Y=1.295
+ $X2=0 $Y2=0
cc_287 N_A_372_397#_c_355_n N_A_221_70#_c_460_n 0.0032544f $X=2.985 $Y=0.377
+ $X2=0 $Y2=0
cc_288 N_A_372_397#_c_357_n N_A_221_70#_c_460_n 0.0218618f $X=3.505 $Y=0.35
+ $X2=0 $Y2=0
cc_289 N_A_372_397#_c_352_n N_A_221_70#_c_462_n 0.00923756f $X=2.037 $Y=1.295
+ $X2=0 $Y2=0
cc_290 N_A_372_397#_c_353_n N_A_221_70#_c_462_n 0.00675243f $X=2.815 $Y=1.21
+ $X2=0 $Y2=0
cc_291 N_A_372_397#_c_360_n N_A_221_70#_c_462_n 0.00377784f $X=1.985 $Y=1.995
+ $X2=0 $Y2=0
cc_292 N_A_372_397#_c_352_n N_A_221_70#_c_473_n 4.28753e-19 $X=2.037 $Y=1.295
+ $X2=0 $Y2=0
cc_293 N_A_372_397#_c_353_n N_A_221_70#_c_473_n 0.0022402f $X=2.815 $Y=1.21
+ $X2=0 $Y2=0
cc_294 N_A_372_397#_c_360_n N_A_221_70#_c_473_n 0.0156912f $X=1.985 $Y=1.995
+ $X2=0 $Y2=0
cc_295 N_A_372_397#_c_365_n N_A_221_70#_c_474_n 0.00376577f $X=1.985 $Y=2.15
+ $X2=0 $Y2=0
cc_296 N_A_372_397#_c_352_n N_A_221_70#_c_463_n 0.00210862f $X=2.037 $Y=1.295
+ $X2=0 $Y2=0
cc_297 N_A_372_397#_c_353_n N_A_221_70#_c_463_n 0.00697157f $X=2.815 $Y=1.21
+ $X2=0 $Y2=0
cc_298 N_A_372_397#_c_360_n N_A_221_70#_M1000_g 0.0110144f $X=1.985 $Y=1.995
+ $X2=0 $Y2=0
cc_299 N_A_372_397#_c_356_n N_A_221_70#_c_464_n 3.20457e-19 $X=3.505 $Y=0.35
+ $X2=0 $Y2=0
cc_300 N_A_372_397#_c_358_n N_A_221_70#_c_464_n 0.0143646f $X=3.25 $Y=1.295
+ $X2=0 $Y2=0
cc_301 N_A_372_397#_c_359_n N_A_221_70#_c_464_n 0.0155314f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_302 N_A_372_397#_c_364_n N_A_221_70#_c_464_n 0.0210518f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_303 N_A_372_397#_c_361_n N_A_221_70#_c_464_n 0.00117185f $X=3.505 $Y=0.515
+ $X2=0 $Y2=0
cc_304 N_A_372_397#_c_354_n N_A_221_70#_M1015_g 0.0120989f $X=2.9 $Y=1.125 $X2=0
+ $Y2=0
cc_305 N_A_372_397#_c_355_n N_A_221_70#_M1015_g 0.00437034f $X=2.985 $Y=0.377
+ $X2=0 $Y2=0
cc_306 N_A_372_397#_c_356_n N_A_221_70#_M1015_g 0.0106486f $X=3.505 $Y=0.35
+ $X2=0 $Y2=0
cc_307 N_A_372_397#_c_358_n N_A_221_70#_M1015_g 0.00492083f $X=3.25 $Y=1.295
+ $X2=0 $Y2=0
cc_308 N_A_372_397#_c_361_n N_A_221_70#_M1015_g 0.0136875f $X=3.505 $Y=0.515
+ $X2=0 $Y2=0
cc_309 N_A_372_397#_c_358_n N_A_221_70#_c_466_n 3.32335e-19 $X=3.25 $Y=1.295
+ $X2=0 $Y2=0
cc_310 N_A_372_397#_c_359_n N_A_221_70#_c_466_n 0.00528327f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_311 N_A_372_397#_c_361_n N_A_221_70#_c_466_n 0.0058952f $X=3.505 $Y=0.515
+ $X2=0 $Y2=0
cc_312 N_A_372_397#_M1009_g N_A_221_70#_M1012_g 0.0118555f $X=3.195 $Y=2.685
+ $X2=0 $Y2=0
cc_313 N_A_372_397#_c_359_n N_A_221_70#_M1012_g 0.00145648f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_314 N_A_372_397#_c_364_n N_A_221_70#_M1012_g 0.0197546f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_315 N_A_372_397#_c_352_n N_A_221_70#_c_469_n 0.011072f $X=2.037 $Y=1.295
+ $X2=0 $Y2=0
cc_316 N_A_372_397#_c_360_n N_A_221_70#_c_469_n 0.0395079f $X=1.985 $Y=1.995
+ $X2=0 $Y2=0
cc_317 N_A_372_397#_c_360_n N_A_221_70#_c_471_n 0.00465937f $X=1.985 $Y=1.995
+ $X2=0 $Y2=0
cc_318 N_A_372_397#_c_365_n N_A_221_70#_c_480_n 0.0194227f $X=1.985 $Y=2.15
+ $X2=0 $Y2=0
cc_319 N_A_372_397#_c_360_n N_A_221_70#_c_480_n 0.00896202f $X=1.985 $Y=1.995
+ $X2=0 $Y2=0
cc_320 N_A_372_397#_c_352_n N_A_221_70#_c_472_n 0.0278769f $X=2.037 $Y=1.295
+ $X2=0 $Y2=0
cc_321 N_A_372_397#_c_357_n N_A_776_99#_c_589_n 0.00129958f $X=3.505 $Y=0.35
+ $X2=0 $Y2=0
cc_322 N_A_372_397#_c_361_n N_A_776_99#_c_589_n 0.0316785f $X=3.505 $Y=0.515
+ $X2=0 $Y2=0
cc_323 N_A_372_397#_c_359_n N_A_776_99#_c_600_n 5.30945e-19 $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_324 N_A_372_397#_c_356_n N_A_626_125#_c_738_n 0.0321506f $X=3.505 $Y=0.35
+ $X2=0 $Y2=0
cc_325 N_A_372_397#_c_357_n N_A_626_125#_c_738_n 0.00308941f $X=3.505 $Y=0.35
+ $X2=0 $Y2=0
cc_326 N_A_372_397#_c_358_n N_A_626_125#_c_738_n 0.015291f $X=3.25 $Y=1.295
+ $X2=0 $Y2=0
cc_327 N_A_372_397#_c_361_n N_A_626_125#_c_738_n 0.00876809f $X=3.505 $Y=0.515
+ $X2=0 $Y2=0
cc_328 N_A_372_397#_c_354_n N_A_626_125#_c_727_n 0.004275f $X=2.9 $Y=1.125 $X2=0
+ $Y2=0
cc_329 N_A_372_397#_c_358_n N_A_626_125#_c_727_n 0.014003f $X=3.25 $Y=1.295
+ $X2=0 $Y2=0
cc_330 N_A_372_397#_c_359_n N_A_626_125#_c_727_n 0.00540853f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_331 N_A_372_397#_c_361_n N_A_626_125#_c_727_n 0.00663848f $X=3.505 $Y=0.515
+ $X2=0 $Y2=0
cc_332 N_A_372_397#_M1009_g N_A_626_125#_c_731_n 0.00969667f $X=3.195 $Y=2.685
+ $X2=0 $Y2=0
cc_333 N_A_372_397#_c_359_n N_A_626_125#_c_731_n 0.00723171f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_334 N_A_372_397#_c_364_n N_A_626_125#_c_731_n 0.00379559f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_335 N_A_372_397#_M1009_g N_A_626_125#_c_732_n 0.00153789f $X=3.195 $Y=2.685
+ $X2=0 $Y2=0
cc_336 N_A_372_397#_c_359_n N_A_626_125#_c_732_n 0.0487175f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_337 N_A_372_397#_c_364_n N_A_626_125#_c_732_n 0.00203002f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_338 N_A_372_397#_c_359_n N_A_626_125#_c_729_n 0.0157919f $X=3.285 $Y=2.04
+ $X2=0 $Y2=0
cc_339 N_A_372_397#_M1009_g N_VPWR_c_872_n 0.00494541f $X=3.195 $Y=2.685 $X2=0
+ $Y2=0
cc_340 N_A_372_397#_M1009_g N_VPWR_c_862_n 0.0101609f $X=3.195 $Y=2.685 $X2=0
+ $Y2=0
cc_341 N_A_372_397#_c_353_n N_VGND_c_985_n 0.0216087f $X=2.815 $Y=1.21 $X2=0
+ $Y2=0
cc_342 N_A_372_397#_c_354_n N_VGND_c_985_n 0.0217004f $X=2.9 $Y=1.125 $X2=0
+ $Y2=0
cc_343 N_A_372_397#_c_355_n N_VGND_c_985_n 0.0216513f $X=2.985 $Y=0.377 $X2=0
+ $Y2=0
cc_344 N_A_372_397#_c_357_n N_VGND_c_985_n 2.91442e-19 $X=3.505 $Y=0.35 $X2=0
+ $Y2=0
cc_345 N_A_372_397#_c_355_n N_VGND_c_986_n 0.0115566f $X=2.985 $Y=0.377 $X2=0
+ $Y2=0
cc_346 N_A_372_397#_c_356_n N_VGND_c_986_n 0.0437853f $X=3.505 $Y=0.35 $X2=0
+ $Y2=0
cc_347 N_A_372_397#_c_357_n N_VGND_c_986_n 0.00647615f $X=3.505 $Y=0.35 $X2=0
+ $Y2=0
cc_348 N_A_372_397#_c_356_n N_VGND_c_987_n 0.0122488f $X=3.505 $Y=0.35 $X2=0
+ $Y2=0
cc_349 N_A_372_397#_c_357_n N_VGND_c_987_n 0.0033626f $X=3.505 $Y=0.35 $X2=0
+ $Y2=0
cc_350 N_A_372_397#_c_361_n N_VGND_c_987_n 0.00107406f $X=3.505 $Y=0.515 $X2=0
+ $Y2=0
cc_351 N_A_372_397#_c_352_n N_VGND_c_991_n 0.00454067f $X=2.037 $Y=1.295 $X2=0
+ $Y2=0
cc_352 N_A_372_397#_c_352_n N_VGND_c_998_n 0.00663239f $X=2.037 $Y=1.295 $X2=0
+ $Y2=0
cc_353 N_A_372_397#_c_355_n N_VGND_c_998_n 0.00579705f $X=2.985 $Y=0.377 $X2=0
+ $Y2=0
cc_354 N_A_372_397#_c_356_n N_VGND_c_998_n 0.0237901f $X=3.505 $Y=0.35 $X2=0
+ $Y2=0
cc_355 N_A_372_397#_c_357_n N_VGND_c_998_n 0.00941423f $X=3.505 $Y=0.35 $X2=0
+ $Y2=0
cc_356 N_A_221_70#_c_464_n N_A_776_99#_c_594_n 0.00163639f $X=3.055 $Y=1.155
+ $X2=0 $Y2=0
cc_357 N_A_221_70#_M1012_g N_A_776_99#_c_608_n 0.0015349f $X=3.74 $Y=2.575 $X2=0
+ $Y2=0
cc_358 N_A_221_70#_M1012_g N_A_776_99#_c_609_n 0.0412023f $X=3.74 $Y=2.575 $X2=0
+ $Y2=0
cc_359 N_A_221_70#_c_466_n N_A_776_99#_c_600_n 0.0412023f $X=3.665 $Y=1.59 $X2=0
+ $Y2=0
cc_360 N_A_221_70#_c_464_n N_A_626_125#_c_738_n 6.08449e-19 $X=3.055 $Y=1.155
+ $X2=0 $Y2=0
cc_361 N_A_221_70#_c_466_n N_A_626_125#_c_738_n 0.0019762f $X=3.665 $Y=1.59
+ $X2=0 $Y2=0
cc_362 N_A_221_70#_c_464_n N_A_626_125#_c_727_n 7.29842e-19 $X=3.055 $Y=1.155
+ $X2=0 $Y2=0
cc_363 N_A_221_70#_M1015_g N_A_626_125#_c_727_n 6.02455e-19 $X=3.055 $Y=0.835
+ $X2=0 $Y2=0
cc_364 N_A_221_70#_c_466_n N_A_626_125#_c_728_n 0.00644146f $X=3.665 $Y=1.59
+ $X2=0 $Y2=0
cc_365 N_A_221_70#_M1012_g N_A_626_125#_c_731_n 0.0186172f $X=3.74 $Y=2.575
+ $X2=0 $Y2=0
cc_366 N_A_221_70#_c_466_n N_A_626_125#_c_732_n 0.00757007f $X=3.665 $Y=1.59
+ $X2=0 $Y2=0
cc_367 N_A_221_70#_M1012_g N_A_626_125#_c_732_n 0.0180612f $X=3.74 $Y=2.575
+ $X2=0 $Y2=0
cc_368 N_A_221_70#_c_464_n N_A_626_125#_c_729_n 9.56206e-19 $X=3.055 $Y=1.155
+ $X2=0 $Y2=0
cc_369 N_A_221_70#_c_466_n N_A_626_125#_c_729_n 0.00434185f $X=3.665 $Y=1.59
+ $X2=0 $Y2=0
cc_370 N_A_221_70#_M1000_g N_VPWR_c_864_n 0.00353601f $X=2.295 $Y=2.685 $X2=0
+ $Y2=0
cc_371 N_A_221_70#_M1012_g N_VPWR_c_911_n 0.00134237f $X=3.74 $Y=2.575 $X2=0
+ $Y2=0
cc_372 N_A_221_70#_M1000_g N_VPWR_c_871_n 0.00367597f $X=2.295 $Y=2.685 $X2=0
+ $Y2=0
cc_373 N_A_221_70#_M1012_g N_VPWR_c_872_n 0.00319315f $X=3.74 $Y=2.575 $X2=0
+ $Y2=0
cc_374 N_A_221_70#_M1000_g N_VPWR_c_862_n 0.00564401f $X=2.295 $Y=2.685 $X2=0
+ $Y2=0
cc_375 N_A_221_70#_M1012_g N_VPWR_c_862_n 0.0031495f $X=3.74 $Y=2.575 $X2=0
+ $Y2=0
cc_376 N_A_221_70#_c_468_n N_VGND_c_984_n 6.7721e-19 $X=1.465 $Y=0.505 $X2=0
+ $Y2=0
cc_377 N_A_221_70#_c_459_n N_VGND_c_985_n 0.0048624f $X=1.75 $Y=1.155 $X2=0
+ $Y2=0
cc_378 N_A_221_70#_c_460_n N_VGND_c_985_n 0.0249217f $X=2.98 $Y=0.18 $X2=0 $Y2=0
cc_379 N_A_221_70#_c_463_n N_VGND_c_985_n 0.00861793f $X=2.265 $Y=1.155 $X2=0
+ $Y2=0
cc_380 N_A_221_70#_M1015_g N_VGND_c_985_n 0.00156431f $X=3.055 $Y=0.835 $X2=0
+ $Y2=0
cc_381 N_A_221_70#_c_460_n N_VGND_c_986_n 0.0131953f $X=2.98 $Y=0.18 $X2=0 $Y2=0
cc_382 N_A_221_70#_c_461_n N_VGND_c_991_n 0.020754f $X=1.825 $Y=0.18 $X2=0 $Y2=0
cc_383 N_A_221_70#_c_468_n N_VGND_c_991_n 0.0234831f $X=1.465 $Y=0.505 $X2=0
+ $Y2=0
cc_384 N_A_221_70#_c_460_n N_VGND_c_998_n 0.0326784f $X=2.98 $Y=0.18 $X2=0 $Y2=0
cc_385 N_A_221_70#_c_461_n N_VGND_c_998_n 0.011455f $X=1.825 $Y=0.18 $X2=0 $Y2=0
cc_386 N_A_221_70#_c_463_n N_VGND_c_998_n 7.97988e-19 $X=2.265 $Y=1.155 $X2=0
+ $Y2=0
cc_387 N_A_221_70#_c_468_n N_VGND_c_998_n 0.0191913f $X=1.465 $Y=0.505 $X2=0
+ $Y2=0
cc_388 N_A_776_99#_c_594_n N_A_626_125#_M1017_g 0.00278593f $X=4.1 $Y=1.23 $X2=0
+ $Y2=0
cc_389 N_A_776_99#_c_596_n N_A_626_125#_M1017_g 0.00467715f $X=5.005 $Y=1.72
+ $X2=0 $Y2=0
cc_390 N_A_776_99#_c_599_n N_A_626_125#_M1017_g 0.0133001f $X=5.005 $Y=1.11
+ $X2=0 $Y2=0
cc_391 N_A_776_99#_M1014_g N_A_626_125#_M1002_g 0.00204187f $X=4.1 $Y=2.575
+ $X2=0 $Y2=0
cc_392 N_A_776_99#_c_604_n N_A_626_125#_M1002_g 0.00988784f $X=4.92 $Y=1.805
+ $X2=0 $Y2=0
cc_393 N_A_776_99#_c_596_n N_A_626_125#_M1002_g 0.00485775f $X=5.005 $Y=1.72
+ $X2=0 $Y2=0
cc_394 N_A_776_99#_c_608_n N_A_626_125#_M1002_g 4.54438e-19 $X=4.19 $Y=1.805
+ $X2=0 $Y2=0
cc_395 N_A_776_99#_c_609_n N_A_626_125#_M1002_g 0.00459209f $X=4.19 $Y=2.025
+ $X2=0 $Y2=0
cc_396 N_A_776_99#_c_610_n N_A_626_125#_M1002_g 0.00530394f $X=5.23 $Y=1.805
+ $X2=0 $Y2=0
cc_397 N_A_776_99#_c_600_n N_A_626_125#_M1002_g 0.0038763f $X=4.19 $Y=1.86 $X2=0
+ $Y2=0
cc_398 N_A_776_99#_c_594_n N_A_626_125#_c_725_n 0.0196771f $X=4.1 $Y=1.23 $X2=0
+ $Y2=0
cc_399 N_A_776_99#_c_604_n N_A_626_125#_c_725_n 0.0105422f $X=4.92 $Y=1.805
+ $X2=0 $Y2=0
cc_400 N_A_776_99#_c_599_n N_A_626_125#_c_725_n 0.00778893f $X=5.005 $Y=1.11
+ $X2=0 $Y2=0
cc_401 N_A_776_99#_c_596_n N_A_626_125#_c_726_n 0.0121833f $X=5.005 $Y=1.72
+ $X2=0 $Y2=0
cc_402 N_A_776_99#_c_589_n N_A_626_125#_c_738_n 0.00220931f $X=3.955 $Y=1.155
+ $X2=0 $Y2=0
cc_403 N_A_776_99#_c_589_n N_A_626_125#_c_727_n 0.00718209f $X=3.955 $Y=1.155
+ $X2=0 $Y2=0
cc_404 N_A_776_99#_c_600_n N_A_626_125#_c_727_n 0.00174876f $X=4.19 $Y=1.86
+ $X2=0 $Y2=0
cc_405 N_A_776_99#_c_594_n N_A_626_125#_c_728_n 0.00656673f $X=4.1 $Y=1.23 $X2=0
+ $Y2=0
cc_406 N_A_776_99#_c_604_n N_A_626_125#_c_728_n 0.0286353f $X=4.92 $Y=1.805
+ $X2=0 $Y2=0
cc_407 N_A_776_99#_c_596_n N_A_626_125#_c_728_n 0.0139401f $X=5.005 $Y=1.72
+ $X2=0 $Y2=0
cc_408 N_A_776_99#_c_608_n N_A_626_125#_c_728_n 0.0258275f $X=4.19 $Y=1.805
+ $X2=0 $Y2=0
cc_409 N_A_776_99#_c_609_n N_A_626_125#_c_728_n 8.97603e-19 $X=4.19 $Y=2.025
+ $X2=0 $Y2=0
cc_410 N_A_776_99#_c_599_n N_A_626_125#_c_728_n 0.0161913f $X=5.005 $Y=1.11
+ $X2=0 $Y2=0
cc_411 N_A_776_99#_c_600_n N_A_626_125#_c_728_n 0.0124158f $X=4.19 $Y=1.86 $X2=0
+ $Y2=0
cc_412 N_A_776_99#_c_609_n N_A_626_125#_c_731_n 0.00244846f $X=4.19 $Y=2.025
+ $X2=0 $Y2=0
cc_413 N_A_776_99#_c_608_n N_A_626_125#_c_732_n 0.0210045f $X=4.19 $Y=1.805
+ $X2=0 $Y2=0
cc_414 N_A_776_99#_c_600_n N_A_626_125#_c_732_n 0.00244846f $X=4.19 $Y=1.86
+ $X2=0 $Y2=0
cc_415 N_A_776_99#_c_596_n N_RESET_B_M1010_g 0.00421859f $X=5.005 $Y=1.72 $X2=0
+ $Y2=0
cc_416 N_A_776_99#_c_647_p N_RESET_B_M1010_g 0.00997615f $X=5.12 $Y=1.98 $X2=0
+ $Y2=0
cc_417 N_A_776_99#_c_598_n N_RESET_B_M1010_g 0.0481778f $X=6.45 $Y=1.46 $X2=0
+ $Y2=0
cc_418 N_A_776_99#_c_610_n N_RESET_B_M1010_g 0.00743185f $X=5.23 $Y=1.805 $X2=0
+ $Y2=0
cc_419 N_A_776_99#_c_650_p N_RESET_B_M1010_g 0.00870484f $X=5.282 $Y=2.4 $X2=0
+ $Y2=0
cc_420 N_A_776_99#_M1001_g N_RESET_B_c_826_n 0.00163405f $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_421 N_A_776_99#_c_599_n N_RESET_B_c_826_n 0.00622188f $X=5.005 $Y=1.11 $X2=0
+ $Y2=0
cc_422 N_A_776_99#_M1001_g N_RESET_B_c_817_n 0.00426907f $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_423 N_A_776_99#_c_596_n N_RESET_B_c_817_n 0.0236172f $X=5.005 $Y=1.72 $X2=0
+ $Y2=0
cc_424 N_A_776_99#_c_599_n N_RESET_B_c_817_n 0.0136055f $X=5.005 $Y=1.11 $X2=0
+ $Y2=0
cc_425 N_A_776_99#_c_610_n N_RESET_B_c_817_n 0.0192315f $X=5.23 $Y=1.805 $X2=0
+ $Y2=0
cc_426 N_A_776_99#_M1001_g N_RESET_B_c_818_n 0.0212037f $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_427 N_A_776_99#_c_596_n N_RESET_B_c_818_n 0.00194387f $X=5.005 $Y=1.72 $X2=0
+ $Y2=0
cc_428 N_A_776_99#_c_610_n N_RESET_B_c_818_n 0.0041043f $X=5.23 $Y=1.805 $X2=0
+ $Y2=0
cc_429 N_A_776_99#_M1001_g N_RESET_B_c_819_n 0.0242997f $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_430 N_A_776_99#_c_599_n N_RESET_B_c_819_n 0.00105933f $X=5.005 $Y=1.11 $X2=0
+ $Y2=0
cc_431 N_A_776_99#_c_604_n N_VPWR_M1014_d 0.00246514f $X=4.92 $Y=1.805 $X2=0
+ $Y2=0
cc_432 N_A_776_99#_c_647_p N_VPWR_M1010_d 0.00531774f $X=5.12 $Y=1.98 $X2=0
+ $Y2=0
cc_433 N_A_776_99#_c_606_n N_VPWR_M1010_d 0.00642121f $X=6.345 $Y=2.4 $X2=0
+ $Y2=0
cc_434 N_A_776_99#_c_610_n N_VPWR_M1010_d 6.64614e-19 $X=5.23 $Y=1.805 $X2=0
+ $Y2=0
cc_435 N_A_776_99#_c_650_p N_VPWR_M1010_d 7.9716e-19 $X=5.282 $Y=2.4 $X2=0 $Y2=0
cc_436 N_A_776_99#_c_606_n N_VPWR_M1020_s 0.00307117f $X=6.345 $Y=2.4 $X2=0
+ $Y2=0
cc_437 N_A_776_99#_c_597_n N_VPWR_M1020_s 0.00430282f $X=6.45 $Y=1.46 $X2=0
+ $Y2=0
cc_438 N_A_776_99#_M1014_g N_VPWR_c_865_n 0.00580703f $X=4.1 $Y=2.575 $X2=0
+ $Y2=0
cc_439 N_A_776_99#_M1014_g N_VPWR_c_866_n 0.00458822f $X=4.1 $Y=2.575 $X2=0
+ $Y2=0
cc_440 N_A_776_99#_c_604_n N_VPWR_c_866_n 0.0220025f $X=4.92 $Y=1.805 $X2=0
+ $Y2=0
cc_441 N_A_776_99#_c_608_n N_VPWR_c_866_n 0.0102881f $X=4.19 $Y=1.805 $X2=0
+ $Y2=0
cc_442 N_A_776_99#_c_609_n N_VPWR_c_866_n 0.00115192f $X=4.19 $Y=2.025 $X2=0
+ $Y2=0
cc_443 N_A_776_99#_M1008_g N_VPWR_c_867_n 0.0119953f $X=5.805 $Y=2.465 $X2=0
+ $Y2=0
cc_444 N_A_776_99#_M1020_g N_VPWR_c_867_n 0.00166911f $X=6.235 $Y=2.465 $X2=0
+ $Y2=0
cc_445 N_A_776_99#_c_606_n N_VPWR_c_867_n 0.0108094f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_446 N_A_776_99#_c_650_p N_VPWR_c_867_n 0.0067145f $X=5.282 $Y=2.4 $X2=0 $Y2=0
cc_447 N_A_776_99#_M1008_g N_VPWR_c_869_n 0.001741f $X=5.805 $Y=2.465 $X2=0
+ $Y2=0
cc_448 N_A_776_99#_M1020_g N_VPWR_c_869_n 0.0153451f $X=6.235 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A_776_99#_c_606_n N_VPWR_c_869_n 0.0236251f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_450 N_A_776_99#_M1014_g N_VPWR_c_911_n 0.00579726f $X=4.1 $Y=2.575 $X2=0
+ $Y2=0
cc_451 N_A_776_99#_c_604_n N_VPWR_c_911_n 0.00627492f $X=4.92 $Y=1.805 $X2=0
+ $Y2=0
cc_452 N_A_776_99#_c_608_n N_VPWR_c_911_n 0.0119208f $X=4.19 $Y=1.805 $X2=0
+ $Y2=0
cc_453 N_A_776_99#_c_609_n N_VPWR_c_911_n 0.00117341f $X=4.19 $Y=2.025 $X2=0
+ $Y2=0
cc_454 N_A_776_99#_M1014_g N_VPWR_c_872_n 0.00382362f $X=4.1 $Y=2.575 $X2=0
+ $Y2=0
cc_455 N_A_776_99#_c_686_p N_VPWR_c_873_n 0.0131621f $X=5.12 $Y=2.91 $X2=0 $Y2=0
cc_456 N_A_776_99#_M1008_g N_VPWR_c_874_n 0.00564095f $X=5.805 $Y=2.465 $X2=0
+ $Y2=0
cc_457 N_A_776_99#_M1020_g N_VPWR_c_874_n 0.00486043f $X=6.235 $Y=2.465 $X2=0
+ $Y2=0
cc_458 N_A_776_99#_M1002_d N_VPWR_c_862_n 0.00395361f $X=4.98 $Y=1.835 $X2=0
+ $Y2=0
cc_459 N_A_776_99#_M1014_g N_VPWR_c_862_n 0.00413371f $X=4.1 $Y=2.575 $X2=0
+ $Y2=0
cc_460 N_A_776_99#_M1008_g N_VPWR_c_862_n 0.00527412f $X=5.805 $Y=2.465 $X2=0
+ $Y2=0
cc_461 N_A_776_99#_M1020_g N_VPWR_c_862_n 0.00462979f $X=6.235 $Y=2.465 $X2=0
+ $Y2=0
cc_462 N_A_776_99#_c_686_p N_VPWR_c_862_n 0.00808656f $X=5.12 $Y=2.91 $X2=0
+ $Y2=0
cc_463 N_A_776_99#_c_606_n N_VPWR_c_862_n 0.0188091f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_464 N_A_776_99#_c_650_p N_VPWR_c_862_n 0.00600135f $X=5.282 $Y=2.4 $X2=0
+ $Y2=0
cc_465 N_A_776_99#_c_606_n N_Q_M1008_d 0.00504536f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_466 N_A_776_99#_M1001_g N_Q_c_965_n 0.00291372f $X=5.805 $Y=0.655 $X2=0 $Y2=0
cc_467 N_A_776_99#_M1008_g N_Q_c_965_n 0.00365595f $X=5.805 $Y=2.465 $X2=0 $Y2=0
cc_468 N_A_776_99#_M1006_g N_Q_c_965_n 0.00568661f $X=6.235 $Y=0.655 $X2=0 $Y2=0
cc_469 N_A_776_99#_M1020_g N_Q_c_965_n 0.00171653f $X=6.235 $Y=2.465 $X2=0 $Y2=0
cc_470 N_A_776_99#_c_606_n N_Q_c_965_n 0.0135055f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_471 N_A_776_99#_c_597_n N_Q_c_965_n 0.0318985f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_472 N_A_776_99#_c_598_n N_Q_c_965_n 0.0213915f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_473 N_A_776_99#_c_610_n N_Q_c_965_n 0.0071569f $X=5.23 $Y=1.805 $X2=0 $Y2=0
cc_474 N_A_776_99#_c_589_n N_VGND_c_986_n 0.00345209f $X=3.955 $Y=1.155 $X2=0
+ $Y2=0
cc_475 N_A_776_99#_c_589_n N_VGND_c_987_n 0.0110351f $X=3.955 $Y=1.155 $X2=0
+ $Y2=0
cc_476 N_A_776_99#_c_594_n N_VGND_c_987_n 0.00411397f $X=4.1 $Y=1.23 $X2=0 $Y2=0
cc_477 N_A_776_99#_c_595_n N_VGND_c_987_n 0.0561862f $X=4.69 $Y=0.42 $X2=0 $Y2=0
cc_478 N_A_776_99#_M1001_g N_VGND_c_988_n 0.0032697f $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_479 N_A_776_99#_M1001_g N_VGND_c_990_n 7.15687e-19 $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_480 N_A_776_99#_M1006_g N_VGND_c_990_n 0.0185691f $X=6.235 $Y=0.655 $X2=0
+ $Y2=0
cc_481 N_A_776_99#_c_597_n N_VGND_c_990_n 0.0211258f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_482 N_A_776_99#_c_598_n N_VGND_c_990_n 0.00362701f $X=6.45 $Y=1.46 $X2=0
+ $Y2=0
cc_483 N_A_776_99#_c_595_n N_VGND_c_992_n 0.0174563f $X=4.69 $Y=0.42 $X2=0 $Y2=0
cc_484 N_A_776_99#_M1001_g N_VGND_c_993_n 0.00585385f $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_485 N_A_776_99#_M1006_g N_VGND_c_993_n 0.00486043f $X=6.235 $Y=0.655 $X2=0
+ $Y2=0
cc_486 N_A_776_99#_M1017_s N_VGND_c_998_n 0.0040649f $X=4.565 $Y=0.235 $X2=0
+ $Y2=0
cc_487 N_A_776_99#_c_589_n N_VGND_c_998_n 0.00394323f $X=3.955 $Y=1.155 $X2=0
+ $Y2=0
cc_488 N_A_776_99#_M1001_g N_VGND_c_998_n 0.0110135f $X=5.805 $Y=0.655 $X2=0
+ $Y2=0
cc_489 N_A_776_99#_M1006_g N_VGND_c_998_n 0.00824727f $X=6.235 $Y=0.655 $X2=0
+ $Y2=0
cc_490 N_A_776_99#_c_595_n N_VGND_c_998_n 0.00963639f $X=4.69 $Y=0.42 $X2=0
+ $Y2=0
cc_491 N_A_776_99#_c_599_n A_996_47# 9.80878e-19 $X=5.005 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_492 N_A_626_125#_c_726_n N_RESET_B_M1010_g 0.0256704f $X=4.905 $Y=1.455 $X2=0
+ $Y2=0
cc_493 N_A_626_125#_M1017_g N_RESET_B_c_826_n 0.00410868f $X=4.905 $Y=0.655
+ $X2=0 $Y2=0
cc_494 N_A_626_125#_M1017_g N_RESET_B_c_817_n 9.78614e-19 $X=4.905 $Y=0.655
+ $X2=0 $Y2=0
cc_495 N_A_626_125#_c_726_n N_RESET_B_c_818_n 0.0428038f $X=4.905 $Y=1.455 $X2=0
+ $Y2=0
cc_496 N_A_626_125#_M1017_g RESET_B 0.00624655f $X=4.905 $Y=0.655 $X2=0 $Y2=0
cc_497 N_A_626_125#_M1017_g N_RESET_B_c_819_n 0.0428038f $X=4.905 $Y=0.655 $X2=0
+ $Y2=0
cc_498 N_A_626_125#_c_731_n N_VPWR_c_864_n 0.00401629f $X=3.43 $Y=2.51 $X2=0
+ $Y2=0
cc_499 N_A_626_125#_M1002_g N_VPWR_c_865_n 0.00869849f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_500 N_A_626_125#_M1002_g N_VPWR_c_866_n 0.00443908f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_501 N_A_626_125#_M1002_g N_VPWR_c_867_n 5.48646e-19 $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_502 N_A_626_125#_M1002_g N_VPWR_c_911_n 0.00355517f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_503 N_A_626_125#_c_731_n N_VPWR_c_911_n 0.024188f $X=3.43 $Y=2.51 $X2=0 $Y2=0
cc_504 N_A_626_125#_c_731_n N_VPWR_c_872_n 0.0234244f $X=3.43 $Y=2.51 $X2=0
+ $Y2=0
cc_505 N_A_626_125#_M1002_g N_VPWR_c_873_n 0.00486043f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_A_626_125#_M1002_g N_VPWR_c_862_n 0.0082726f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_507 N_A_626_125#_c_731_n N_VPWR_c_862_n 0.0170351f $X=3.43 $Y=2.51 $X2=0
+ $Y2=0
cc_508 N_A_626_125#_c_738_n N_VGND_c_986_n 7.42881e-19 $X=3.55 $Y=0.812 $X2=0
+ $Y2=0
cc_509 N_A_626_125#_M1017_g N_VGND_c_987_n 0.00345876f $X=4.905 $Y=0.655 $X2=0
+ $Y2=0
cc_510 N_A_626_125#_c_738_n N_VGND_c_987_n 0.0155438f $X=3.55 $Y=0.812 $X2=0
+ $Y2=0
cc_511 N_A_626_125#_c_727_n N_VGND_c_987_n 0.00220954f $X=3.635 $Y=1.365 $X2=0
+ $Y2=0
cc_512 N_A_626_125#_c_728_n N_VGND_c_987_n 0.0137053f $X=4.575 $Y=1.455 $X2=0
+ $Y2=0
cc_513 N_A_626_125#_M1017_g N_VGND_c_992_n 0.00538152f $X=4.905 $Y=0.655 $X2=0
+ $Y2=0
cc_514 N_A_626_125#_M1017_g N_VGND_c_998_n 0.0107178f $X=4.905 $Y=0.655 $X2=0
+ $Y2=0
cc_515 N_A_626_125#_c_738_n N_VGND_c_998_n 0.00173642f $X=3.55 $Y=0.812 $X2=0
+ $Y2=0
cc_516 N_A_626_125#_c_738_n A_726_125# 0.00363995f $X=3.55 $Y=0.812 $X2=-0.19
+ $Y2=-0.245
cc_517 N_A_626_125#_c_727_n A_726_125# 9.70695e-19 $X=3.635 $Y=1.365 $X2=-0.19
+ $Y2=-0.245
cc_518 N_RESET_B_M1010_g N_VPWR_c_867_n 0.00876677f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_519 N_RESET_B_M1010_g N_VPWR_c_911_n 6.40375e-19 $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_520 N_RESET_B_M1010_g N_VPWR_c_873_n 0.00564095f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_521 N_RESET_B_M1010_g N_VPWR_c_862_n 0.00521882f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_522 N_RESET_B_M1010_g N_Q_c_965_n 4.83547e-19 $X=5.335 $Y=2.465 $X2=0 $Y2=0
cc_523 N_RESET_B_c_817_n N_Q_c_965_n 0.0221528f $X=5.355 $Y=1.35 $X2=0 $Y2=0
cc_524 N_RESET_B_c_818_n N_Q_c_965_n 5.91817e-19 $X=5.355 $Y=1.35 $X2=0 $Y2=0
cc_525 N_RESET_B_c_826_n N_VGND_M1011_d 0.00366335f $X=5.39 $Y=0.855 $X2=0 $Y2=0
cc_526 N_RESET_B_c_817_n N_VGND_M1011_d 0.00302103f $X=5.355 $Y=1.35 $X2=0 $Y2=0
cc_527 N_RESET_B_c_826_n N_VGND_c_988_n 0.0095183f $X=5.39 $Y=0.855 $X2=0 $Y2=0
cc_528 N_RESET_B_c_819_n N_VGND_c_988_n 0.00331551f $X=5.355 $Y=1.185 $X2=0
+ $Y2=0
cc_529 N_RESET_B_c_826_n N_VGND_c_992_n 0.00237326f $X=5.39 $Y=0.855 $X2=0 $Y2=0
cc_530 RESET_B N_VGND_c_992_n 0.00706477f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_531 N_RESET_B_c_819_n N_VGND_c_992_n 0.00432313f $X=5.355 $Y=1.185 $X2=0
+ $Y2=0
cc_532 N_RESET_B_c_826_n N_VGND_c_998_n 0.00460257f $X=5.39 $Y=0.855 $X2=0 $Y2=0
cc_533 RESET_B N_VGND_c_998_n 0.00826571f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_534 N_RESET_B_c_819_n N_VGND_c_998_n 0.00594161f $X=5.355 $Y=1.185 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_826_n A_996_47# 0.00247373f $X=5.39 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_536 RESET_B A_996_47# 0.00144399f $X=4.955 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_537 N_VPWR_c_862_n N_Q_M1008_d 0.00412982f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_538 N_Q_c_965_n N_VGND_c_990_n 0.032257f $X=6.02 $Y=0.42 $X2=0 $Y2=0
cc_539 N_Q_c_965_n N_VGND_c_993_n 0.0131621f $X=6.02 $Y=0.42 $X2=0 $Y2=0
cc_540 N_Q_M1001_d N_VGND_c_998_n 0.00467071f $X=5.88 $Y=0.235 $X2=0 $Y2=0
cc_541 N_Q_c_965_n N_VGND_c_998_n 0.00808656f $X=6.02 $Y=0.42 $X2=0 $Y2=0
cc_542 N_VGND_c_998_n A_996_47# 0.00181742f $X=6.48 $Y=0 $X2=-0.19 $Y2=-0.245
