* File: sky130_fd_sc_lp__nor4_lp.pex.spice
* Created: Fri Aug 28 10:57:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4_LP%C 3 7 9 13 16 18 19 21 28
c41 28 0 1.68228e-19 $X=0.525 $Y=1.275
c42 9 0 1.55496e-19 $X=0.9 $Y=1.185
r43 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.275 $X2=0.525 $Y2=1.275
r44 21 29 3.48112 $w=6.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.72 $Y=1.445
+ $X2=0.525 $Y2=1.445
r45 19 29 5.0878 $w=6.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=1.445
+ $X2=0.525 $Y2=1.445
r46 17 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=1.615
+ $X2=0.525 $Y2=1.275
r47 17 18 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.615
+ $X2=0.525 $Y2=1.78
r48 15 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.525 $Y=1.26
+ $X2=0.525 $Y2=1.275
r49 15 16 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=0.525 $Y=1.26
+ $X2=0.525 $Y2=1.185
r50 11 13 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.975 $Y=1.11
+ $X2=0.975 $Y2=0.495
r51 10 16 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.69 $Y=1.185
+ $X2=0.525 $Y2=1.185
r52 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.9 $Y=1.185
+ $X2=0.975 $Y2=1.11
r53 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.9 $Y=1.185 $X2=0.69
+ $Y2=1.185
r54 5 16 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.615 $Y=1.11
+ $X2=0.525 $Y2=1.185
r55 5 7 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.615 $Y=1.11
+ $X2=0.615 $Y2=0.495
r56 3 18 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.545 $Y=2.545
+ $X2=0.545 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%D 3 7 11 13 14 20
c43 20 0 3.67825e-19 $X=1.675 $Y=1.29
c44 14 0 8.73928e-20 $X=2.16 $Y=1.295
r45 20 22 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=1.675 $Y=1.29
+ $X2=1.765 $Y2=1.29
r46 18 20 7.24812 $w=2.66e-07 $l=4e-08 $layer=POLY_cond $X=1.635 $Y=1.29
+ $X2=1.675 $Y2=1.29
r47 13 14 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.675 $Y=1.29
+ $X2=2.16 $Y2=1.29
r48 13 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.29 $X2=1.675 $Y2=1.29
r49 9 22 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.125
+ $X2=1.765 $Y2=1.29
r50 9 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.765 $Y=1.125
+ $X2=1.765 $Y2=0.495
r51 5 18 4.31405 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.455
+ $X2=1.635 $Y2=1.29
r52 5 7 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.635 $Y=1.455 $X2=1.635
+ $Y2=2.155
r53 1 18 41.6767 $w=2.66e-07 $l=3.01413e-07 $layer=POLY_cond $X=1.405 $Y=1.125
+ $X2=1.635 $Y2=1.29
r54 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.405 $Y=1.125
+ $X2=1.405 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%B 1 3 4 5 6 8 12 15 17 18 19 20 24 26
c57 19 0 1.99597e-19 $X=2.64 $Y=1.295
c58 17 0 2.52295e-20 $X=2.555 $Y=0.855
c59 12 0 1.57071e-19 $X=2.665 $Y=1.66
r60 24 26 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.34
+ $X2=2.665 $Y2=1.175
r61 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=1.295
+ $X2=2.645 $Y2=1.665
r62 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.645
+ $Y=1.34 $X2=2.645 $Y2=1.34
r63 15 18 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.725 $Y=2.545
+ $X2=2.725 $Y2=1.845
r64 12 18 34.9505 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.665 $Y=1.66
+ $X2=2.665 $Y2=1.845
r65 11 24 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=2.665 $Y=1.36
+ $X2=2.665 $Y2=1.34
r66 11 12 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=2.665 $Y=1.36
+ $X2=2.665 $Y2=1.66
r67 9 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.555 $Y=0.93
+ $X2=2.555 $Y2=0.855
r68 9 26 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=2.555 $Y=0.93
+ $X2=2.555 $Y2=1.175
r69 6 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.555 $Y=0.78
+ $X2=2.555 $Y2=0.855
r70 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.555 $Y=0.78 $X2=2.555
+ $Y2=0.495
r71 4 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.48 $Y=0.855
+ $X2=2.555 $Y2=0.855
r72 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.48 $Y=0.855 $X2=2.27
+ $Y2=0.855
r73 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.195 $Y=0.78
+ $X2=2.27 $Y2=0.855
r74 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.195 $Y=0.78 $X2=2.195
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%A 1 3 6 8 10 15 17 18 19 23 24
c41 24 0 2.52295e-20 $X=3.355 $Y=1.07
c42 23 0 9.31175e-20 $X=3.355 $Y=1.07
c43 8 0 4.46818e-20 $X=3.345 $Y=0.785
r44 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.355
+ $Y=1.07 $X2=3.355 $Y2=1.07
r45 18 19 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=3.452 $Y=1.295
+ $X2=3.452 $Y2=1.665
r46 18 24 5.12605 $w=5.23e-07 $l=2.25e-07 $layer=LI1_cond $X=3.452 $Y=1.295
+ $X2=3.452 $Y2=1.07
r47 17 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.355 $Y=1.41
+ $X2=3.355 $Y2=1.07
r48 15 23 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.355 $Y=0.935
+ $X2=3.355 $Y2=1.07
r49 13 15 5.12766 $w=1.5e-07 $l=1e-08 $layer=POLY_cond $X=3.345 $Y=0.86
+ $X2=3.355 $Y2=0.86
r50 11 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.985 $Y=0.86
+ $X2=3.345 $Y2=0.86
r51 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.345 $Y=0.785
+ $X2=3.345 $Y2=0.86
r52 8 10 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.345 $Y=0.785
+ $X2=3.345 $Y2=0.495
r53 4 17 47.383 $w=2.95e-07 $l=3.53129e-07 $layer=POLY_cond $X=3.215 $Y=1.7
+ $X2=3.355 $Y2=1.41
r54 4 6 209.943 $w=2.5e-07 $l=8.45e-07 $layer=POLY_cond $X=3.215 $Y=1.7
+ $X2=3.215 $Y2=2.545
r55 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.985 $Y=0.785
+ $X2=2.985 $Y2=0.86
r56 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.985 $Y=0.785
+ $X2=2.985 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%A_27_409# 1 2 7 9 11 15 19 23
r35 17 23 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.9 $Y=2.315 $X2=1.9
+ $Y2=2.23
r36 17 19 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.9 $Y=2.315
+ $X2=1.9 $Y2=2.51
r37 13 23 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.9 $Y=2.145 $X2=1.9
+ $Y2=2.23
r38 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.9 $Y=2.145
+ $X2=1.9 $Y2=1.8
r39 12 22 4.72267 $w=1.7e-07 $l=1.92678e-07 $layer=LI1_cond $X=0.445 $Y=2.23
+ $X2=0.28 $Y2=2.17
r40 11 23 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=2.23
+ $X2=1.9 $Y2=2.23
r41 11 12 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=1.735 $Y=2.23
+ $X2=0.445 $Y2=2.23
r42 7 22 3.0435 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=0.28 $Y=2.315 $X2=0.28
+ $Y2=2.17
r43 7 9 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=0.28 $Y=2.315
+ $X2=0.28 $Y2=2.9
r44 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=1.655 $X2=1.9 $Y2=2.51
r45 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=1.655 $X2=1.9 $Y2=1.8
r46 1 22 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r47 1 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%A_134_409# 1 2 9 11 12 13 15
r31 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.895 $X2=2.46
+ $Y2=2.98
r32 13 15 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=2.46 $Y=2.895
+ $X2=2.46 $Y2=2.19
r33 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=2.98
+ $X2=2.46 $Y2=2.98
r34 11 12 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=2.295 $Y=2.98
+ $X2=0.975 $Y2=2.98
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.81 $Y=2.895
+ $X2=0.975 $Y2=2.98
r36 7 9 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.81 $Y=2.895
+ $X2=0.81 $Y2=2.78
r37 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.045 $X2=2.46 $Y2=2.9
r38 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.045 $X2=2.46 $Y2=2.19
r39 1 9 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%Y 1 2 3 12 14 18 20 21 22 41
c56 41 0 2.54009e-19 $X=1.37 $Y=1.8
c57 14 0 1.37799e-19 $X=2.605 $Y=0.86
r58 29 36 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=1.635
+ $X2=1.17 $Y2=1.8
r59 22 41 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.2 $Y=1.8 $X2=1.37
+ $Y2=1.8
r60 22 36 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.2 $Y=1.8 $X2=1.17
+ $Y2=1.8
r61 22 29 1.1127 $w=2.88e-07 $l=2.8e-08 $layer=LI1_cond $X=1.17 $Y=1.607
+ $X2=1.17 $Y2=1.635
r62 21 22 12.3987 $w=2.88e-07 $l=3.12e-07 $layer=LI1_cond $X=1.17 $Y=1.295
+ $X2=1.17 $Y2=1.607
r63 20 28 3.05675 $w=3.1e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.19 $Y=0.86
+ $X2=1.17 $Y2=0.945
r64 20 21 12.6371 $w=2.88e-07 $l=3.18e-07 $layer=LI1_cond $X=1.17 $Y=0.977
+ $X2=1.17 $Y2=1.295
r65 20 28 1.27166 $w=2.88e-07 $l=3.2e-08 $layer=LI1_cond $X=1.17 $Y=0.977
+ $X2=1.17 $Y2=0.945
r66 16 18 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.77 $Y=0.775
+ $X2=2.77 $Y2=0.495
r67 15 20 3.57226 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0.86
+ $X2=1.19 $Y2=0.86
r68 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.605 $Y=0.86
+ $X2=2.77 $Y2=0.775
r69 14 15 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.605 $Y=0.86
+ $X2=1.355 $Y2=0.86
r70 10 20 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=0.775
+ $X2=1.19 $Y2=0.86
r71 10 12 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.19 $Y=0.775
+ $X2=1.19 $Y2=0.495
r72 3 41 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=1.655 $X2=1.37 $Y2=1.8
r73 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.63
+ $Y=0.285 $X2=2.77 $Y2=0.495
r74 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.285 $X2=1.19 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%VPWR 1 4 6 10 12 22
r23 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r24 19 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r25 18 19 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r26 14 18 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.12 $Y2=3.33
r27 14 15 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 12 21 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.577 $Y2=3.33
r29 12 18 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.12 $Y2=3.33
r30 10 19 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r31 10 15 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 6 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.48 $Y=2.19 $X2=3.48
+ $Y2=2.9
r33 4 21 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.577 $Y2=3.33
r34 4 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.48 $Y2=2.9
r35 1 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.045 $X2=3.48 $Y2=2.9
r36 1 6 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.045 $X2=3.48 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_LP%VGND 1 2 3 10 12 16 18 20 23 24 25 34 46
r49 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 40 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r52 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r54 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r55 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 34 45 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.617
+ $Y2=0
r57 34 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.12
+ $Y2=0
r58 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r60 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r61 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r62 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r63 27 42 4.52228 $w=1.7e-07 $l=2.83e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.282
+ $Y2=0
r64 27 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.72
+ $Y2=0
r65 25 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r66 25 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r67 23 32 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.68
+ $Y2=0
r68 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r69 22 36 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.16
+ $Y2=0
r70 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r71 18 45 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.617 $Y2=0
r72 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0.495
r73 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r74 14 16 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.43
r75 10 42 3.2439 $w=3.3e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.4 $Y=0.085
+ $X2=0.282 $Y2=0
r76 10 12 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.4 $Y=0.085 $X2=0.4
+ $Y2=0.495
r77 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.285 $X2=3.56 $Y2=0.495
r78 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.285 $X2=1.98 $Y2=0.43
r79 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.285 $X2=0.4 $Y2=0.495
.ends

