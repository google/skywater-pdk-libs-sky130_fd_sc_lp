* File: sky130_fd_sc_lp__a2bb2oi_4.spice
* Created: Fri Aug 28 09:56:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2oi_4.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2oi_4  VNB VPB B1 B2 A1_N A2_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2_N	A2_N
* A1_N	A1_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_B1_M1003_g N_A_157_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75009
+ A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_B1_M1013_g N_A_157_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75008.5 A=0.126 P=1.98 MULT=1
MM1025 N_VGND_M1013_d N_B1_M1025_g N_A_157_47#_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75008.1 A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_B2_M1004_g N_A_157_47#_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75007.7 A=0.126 P=1.98 MULT=1
MM1010 N_Y_M1004_d N_B2_M1010_g N_A_157_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75007.2 A=0.126 P=1.98 MULT=1
MM1020 N_Y_M1020_d N_B2_M1020_g N_A_157_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75006.8 A=0.126 P=1.98 MULT=1
MM1023 N_Y_M1020_d N_B2_M1023_g N_A_157_47#_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75006.4 A=0.126 P=1.98 MULT=1
MM1035 N_VGND_M1035_d N_B1_M1035_g N_A_157_47#_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1533 AS=0.1176 PD=1.205 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75006 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1035_d N_A_832_21#_M1017_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1533 AS=0.1176 PD=1.205 PS=1.12 NRD=6.42 NRS=0 M=1 R=5.6 SA=75003.7
+ SB=75005.4 A=0.126 P=1.98 MULT=1
MM1030 N_VGND_M1030_d N_A_832_21#_M1030_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1 SB=75005
+ A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1030_d N_A_832_21#_M1031_g N_Y_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.6
+ SB=75004.6 A=0.126 P=1.98 MULT=1
MM1037 N_VGND_M1037_d N_A_832_21#_M1037_g N_Y_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005 SB=75004.1
+ A=0.126 P=1.98 MULT=1
MM1006 N_A_832_21#_M1006_d N_A1_N_M1006_g N_VGND_M1037_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.4
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1011 N_A_832_21#_M1006_d N_A1_N_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.9
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1022 N_A_832_21#_M1022_d N_A1_N_M1022_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.3
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1026 N_A_832_21#_M1022_d N_A1_N_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.336 PD=1.12 PS=1.64 NRD=0 NRS=24.756 M=1 R=5.6
+ SA=75006.7 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1007 N_A_832_21#_M1007_d N_A2_N_M1007_g N_VGND_M1026_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.336 PD=1.12 PS=1.64 NRD=0 NRS=49.512 M=1 R=5.6
+ SA=75007.7 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1024 N_A_832_21#_M1007_d N_A2_N_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1027 N_A_832_21#_M1027_d N_A2_N_M1027_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1039 N_A_832_21#_M1027_d N_A2_N_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75009
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_73_367#_M1002_d N_B1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1005 N_A_73_367#_M1005_d N_B1_M1005_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_73_367#_M1005_d N_B1_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_73_367#_M1000_d N_B2_M1000_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.8 A=0.189 P=2.82 MULT=1
MM1012 N_A_73_367#_M1000_d N_B2_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1021 N_A_73_367#_M1021_d N_B2_M1021_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1034 N_A_73_367#_M1021_d N_B2_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.283 PD=1.54 PS=1.74 NRD=0 NRS=12.8838 M=1 R=8.4 SA=75002.8
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1018 N_A_73_367#_M1018_d N_B1_M1018_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.283 PD=1.54 PS=1.74 NRD=0 NRS=12.8838 M=1 R=8.4 SA=75003.4
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_832_21#_M1001_g N_A_73_367#_M1018_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1001_d N_A_832_21#_M1016_g N_A_73_367#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1028 N_Y_M1028_d N_A_832_21#_M1028_g N_A_73_367#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1036 N_Y_M1028_d N_A_832_21#_M1036_g N_A_73_367#_M1036_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1008 N_A_1241_367#_M1008_d N_A1_N_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1019 N_A_1241_367#_M1019_d N_A1_N_M1019_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1029 N_A_1241_367#_M1019_d N_A1_N_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1038 N_A_1241_367#_M1038_d N_A1_N_M1038_g N_VPWR_M1029_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_A_832_21#_M1009_d N_A2_N_M1009_g N_A_1241_367#_M1038_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1015 N_A_832_21#_M1009_d N_A2_N_M1015_g N_A_1241_367#_M1015_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1032 N_A_832_21#_M1032_d N_A2_N_M1032_g N_A_1241_367#_M1015_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1033 N_A_832_21#_M1032_d N_A2_N_M1033_g N_A_1241_367#_M1033_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.5079 P=24.65
c_156 VPB 0 9.18783e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a2bb2oi_4.pxi.spice"
*
.ends
*
*
