* File: sky130_fd_sc_lp__nor4bb_1.pxi.spice
* Created: Fri Aug 28 10:58:54 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4BB_1%D_N N_D_N_M1002_g N_D_N_M1006_g D_N D_N D_N
+ N_D_N_c_75_n PM_SKY130_FD_SC_LP__NOR4BB_1%D_N
x_PM_SKY130_FD_SC_LP__NOR4BB_1%A_27_508# N_A_27_508#_M1006_s N_A_27_508#_M1002_s
+ N_A_27_508#_c_106_n N_A_27_508#_M1009_g N_A_27_508#_c_107_n
+ N_A_27_508#_M1004_g N_A_27_508#_c_113_n N_A_27_508#_c_114_n
+ N_A_27_508#_c_115_n N_A_27_508#_c_108_n N_A_27_508#_c_109_n
+ N_A_27_508#_c_110_n N_A_27_508#_c_111_n PM_SKY130_FD_SC_LP__NOR4BB_1%A_27_508#
x_PM_SKY130_FD_SC_LP__NOR4BB_1%A_375_269# N_A_375_269#_M1010_d
+ N_A_375_269#_M1003_d N_A_375_269#_M1011_g N_A_375_269#_M1001_g
+ N_A_375_269#_c_174_n N_A_375_269#_c_168_n N_A_375_269#_c_184_p
+ N_A_375_269#_c_181_n N_A_375_269#_c_169_n N_A_375_269#_c_170_n
+ N_A_375_269#_c_171_n N_A_375_269#_c_177_n N_A_375_269#_c_172_n
+ N_A_375_269#_c_203_p PM_SKY130_FD_SC_LP__NOR4BB_1%A_375_269#
x_PM_SKY130_FD_SC_LP__NOR4BB_1%B N_B_M1005_g N_B_M1007_g B N_B_c_245_n
+ N_B_c_248_n PM_SKY130_FD_SC_LP__NOR4BB_1%B
x_PM_SKY130_FD_SC_LP__NOR4BB_1%A N_A_M1000_g N_A_M1008_g A A N_A_c_280_n
+ N_A_c_281_n PM_SKY130_FD_SC_LP__NOR4BB_1%A
x_PM_SKY130_FD_SC_LP__NOR4BB_1%C_N N_C_N_M1003_g N_C_N_M1010_g C_N N_C_N_c_319_n
+ PM_SKY130_FD_SC_LP__NOR4BB_1%C_N
x_PM_SKY130_FD_SC_LP__NOR4BB_1%VPWR N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_c_346_n
+ N_VPWR_c_347_n VPWR N_VPWR_c_348_n N_VPWR_c_349_n N_VPWR_c_350_n
+ N_VPWR_c_345_n N_VPWR_c_352_n N_VPWR_c_353_n PM_SKY130_FD_SC_LP__NOR4BB_1%VPWR
x_PM_SKY130_FD_SC_LP__NOR4BB_1%Y N_Y_M1009_d N_Y_M1007_d N_Y_M1004_s N_Y_c_387_n
+ N_Y_c_429_p N_Y_c_384_n N_Y_c_388_n N_Y_c_385_n N_Y_c_386_n Y Y N_Y_c_416_n
+ PM_SKY130_FD_SC_LP__NOR4BB_1%Y
x_PM_SKY130_FD_SC_LP__NOR4BB_1%VGND N_VGND_M1006_d N_VGND_M1001_d N_VGND_M1000_d
+ N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n
+ VGND N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n
+ N_VGND_c_454_n N_VGND_c_455_n PM_SKY130_FD_SC_LP__NOR4BB_1%VGND
cc_1 VNB N_D_N_M1006_g 0.0276641f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_2 VNB D_N 0.0362377f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_D_N_c_75_n 0.0504562f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.375
cc_4 VNB N_A_27_508#_c_106_n 0.0188815f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_5 VNB N_A_27_508#_c_107_n 0.0581885f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_508#_c_108_n 0.0143362f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.88
cc_7 VNB N_A_27_508#_c_109_n 0.00152445f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=1.665
cc_8 VNB N_A_27_508#_c_110_n 0.00170072f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=2.035
cc_9 VNB N_A_27_508#_c_111_n 0.00711827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_375_269#_M1001_g 0.0247792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_375_269#_c_168_n 0.0254562f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.21
cc_12 VNB N_A_375_269#_c_169_n 0.00513817f $X=-0.19 $Y=-0.245 $X2=0.367
+ $Y2=1.375
cc_13 VNB N_A_375_269#_c_170_n 0.0142114f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=1.665
cc_14 VNB N_A_375_269#_c_171_n 0.00367898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_375_269#_c_172_n 0.0145889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1007_g 0.0254607f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_17 VNB N_B_c_245_n 0.0254884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_M1008_g 0.0069202f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_19 VNB A 0.00253756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_280_n 0.0359503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_281_n 0.0193341f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.375
cc_22 VNB N_C_N_M1010_g 0.0352907f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_23 VNB C_N 0.0126655f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_C_N_c_319_n 0.0422892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_345_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_384_n 0.015057f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=1.295
cc_27 VNB N_Y_c_385_n 0.00318663f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=1.665
cc_28 VNB N_Y_c_386_n 0.00678913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_445_n 0.0166662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_446_n 0.0149824f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.375
cc_31 VNB N_VGND_c_447_n 0.00461085f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=1.295
cc_32 VNB N_VGND_c_448_n 0.0180616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_449_n 0.0197888f $X=-0.19 $Y=-0.245 $X2=0.367 $Y2=2.035
cc_34 VNB N_VGND_c_450_n 0.0368914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_451_n 0.0193417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_452_n 0.26509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_453_n 0.00609605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_454_n 0.00519006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_455_n 0.0116741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_D_N_M1002_g 0.066891f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.75
cc_41 VPB D_N 0.0272189f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_42 VPB N_D_N_c_75_n 0.0326751f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.375
cc_43 VPB N_A_27_508#_c_107_n 0.0299584f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_44 VPB N_A_27_508#_c_113_n 0.0186382f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.375
cc_45 VPB N_A_27_508#_c_114_n 0.0176419f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.375
cc_46 VPB N_A_27_508#_c_115_n 0.0101244f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.21
cc_47 VPB N_A_27_508#_c_110_n 0.0101313f $X=-0.19 $Y=1.655 $X2=0.367 $Y2=2.035
cc_48 VPB N_A_375_269#_M1011_g 0.0187018f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_49 VPB N_A_375_269#_c_174_n 0.0013665f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.375
cc_50 VPB N_A_375_269#_c_168_n 0.00647803f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.21
cc_51 VPB N_A_375_269#_c_169_n 0.00145323f $X=-0.19 $Y=1.655 $X2=0.367 $Y2=1.375
cc_52 VPB N_A_375_269#_c_177_n 0.0106564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B_M1005_g 0.0211083f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.75
cc_54 VPB N_B_c_245_n 0.00647941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B_c_248_n 0.00228237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_M1008_g 0.0233589f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.865
cc_57 VPB A 0.00168545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_C_N_M1003_g 0.0300554f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.75
cc_59 VPB C_N 0.0172265f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_60 VPB N_C_N_c_319_n 0.0137141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_346_n 0.0108563f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_62 VPB N_VPWR_c_347_n 0.0312261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_348_n 0.0169002f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.375
cc_64 VPB N_VPWR_c_349_n 0.0649802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_350_n 0.0311013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_345_n 0.0969339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_352_n 0.00613202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_353_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_Y_c_387_n 0.0123337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_Y_c_388_n 0.00521053f $X=-0.19 $Y=1.655 $X2=0.367 $Y2=1.375
cc_71 VPB N_Y_c_385_n 9.76208e-19 $X=-0.19 $Y=1.655 $X2=0.367 $Y2=1.665
cc_72 N_D_N_M1006_g N_A_27_508#_c_106_n 0.00536942f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_73 N_D_N_M1006_g N_A_27_508#_c_107_n 0.0214965f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_74 N_D_N_c_75_n N_A_27_508#_c_107_n 0.00752086f $X=0.565 $Y=1.375 $X2=0 $Y2=0
cc_75 N_D_N_M1002_g N_A_27_508#_c_113_n 0.0036463f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_76 N_D_N_M1002_g N_A_27_508#_c_114_n 0.0172689f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_77 D_N N_A_27_508#_c_114_n 0.0235506f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_D_N_c_75_n N_A_27_508#_c_114_n 0.00586566f $X=0.565 $Y=1.375 $X2=0 $Y2=0
cc_79 D_N N_A_27_508#_c_115_n 0.0242234f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_D_N_M1006_g N_A_27_508#_c_108_n 0.0154328f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_81 D_N N_A_27_508#_c_108_n 0.0190988f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_D_N_c_75_n N_A_27_508#_c_108_n 0.00419582f $X=0.565 $Y=1.375 $X2=0 $Y2=0
cc_83 N_D_N_M1006_g N_A_27_508#_c_109_n 0.00850397f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_84 N_D_N_M1002_g N_A_27_508#_c_110_n 0.00668891f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_85 D_N N_A_27_508#_c_110_n 0.0478149f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_D_N_c_75_n N_A_27_508#_c_110_n 0.0129697f $X=0.565 $Y=1.375 $X2=0 $Y2=0
cc_87 N_D_N_M1006_g N_A_27_508#_c_111_n 0.00154751f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_88 D_N N_A_27_508#_c_111_n 0.0251789f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_D_N_c_75_n N_A_27_508#_c_111_n 0.00918793f $X=0.565 $Y=1.375 $X2=0 $Y2=0
cc_90 N_D_N_M1002_g N_VPWR_c_346_n 0.0140126f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_91 N_D_N_M1002_g N_VPWR_c_348_n 0.00383152f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_92 N_D_N_M1002_g N_VPWR_c_345_n 0.00761127f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_93 N_D_N_M1002_g N_Y_c_387_n 0.00526703f $X=0.475 $Y=2.75 $X2=0 $Y2=0
cc_94 N_D_N_c_75_n N_Y_c_388_n 2.14269e-19 $X=0.565 $Y=1.375 $X2=0 $Y2=0
cc_95 N_D_N_c_75_n N_Y_c_385_n 3.38322e-19 $X=0.565 $Y=1.375 $X2=0 $Y2=0
cc_96 N_D_N_M1006_g N_VGND_c_445_n 0.00499928f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_97 N_D_N_M1006_g N_VGND_c_450_n 0.00313467f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_98 N_D_N_M1006_g N_VGND_c_452_n 0.0046122f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_99 N_A_27_508#_c_106_n N_A_375_269#_M1001_g 0.0225548f $X=1.59 $Y=1.185 $X2=0
+ $Y2=0
cc_100 N_A_27_508#_c_107_n N_A_375_269#_c_174_n 5.98135e-19 $X=1.59 $Y=1.725
+ $X2=0 $Y2=0
cc_101 N_A_27_508#_c_107_n N_A_375_269#_c_168_n 0.114699f $X=1.59 $Y=1.725 $X2=0
+ $Y2=0
cc_102 N_A_27_508#_c_107_n N_A_375_269#_c_181_n 2.56625e-19 $X=1.59 $Y=1.725
+ $X2=0 $Y2=0
cc_103 N_A_27_508#_c_107_n N_VPWR_c_346_n 0.00281504f $X=1.59 $Y=1.725 $X2=0
+ $Y2=0
cc_104 N_A_27_508#_c_114_n N_VPWR_c_346_n 0.0247108f $X=0.82 $Y=2.375 $X2=0
+ $Y2=0
cc_105 N_A_27_508#_c_113_n N_VPWR_c_348_n 0.00880077f $X=0.26 $Y=2.755 $X2=0
+ $Y2=0
cc_106 N_A_27_508#_c_107_n N_VPWR_c_349_n 0.00357668f $X=1.59 $Y=1.725 $X2=0
+ $Y2=0
cc_107 N_A_27_508#_c_107_n N_VPWR_c_345_n 0.00648284f $X=1.59 $Y=1.725 $X2=0
+ $Y2=0
cc_108 N_A_27_508#_c_113_n N_VPWR_c_345_n 0.00914991f $X=0.26 $Y=2.755 $X2=0
+ $Y2=0
cc_109 N_A_27_508#_c_107_n N_Y_c_387_n 0.0207279f $X=1.59 $Y=1.725 $X2=0 $Y2=0
cc_110 N_A_27_508#_c_114_n N_Y_c_387_n 0.0148498f $X=0.82 $Y=2.375 $X2=0 $Y2=0
cc_111 N_A_27_508#_c_107_n N_Y_c_388_n 0.0167529f $X=1.59 $Y=1.725 $X2=0 $Y2=0
cc_112 N_A_27_508#_c_110_n N_Y_c_388_n 0.0377917f $X=0.925 $Y=2.29 $X2=0 $Y2=0
cc_113 N_A_27_508#_c_111_n N_Y_c_388_n 0.0079548f $X=1.26 $Y=1.35 $X2=0 $Y2=0
cc_114 N_A_27_508#_c_107_n N_Y_c_385_n 0.0174164f $X=1.59 $Y=1.725 $X2=0 $Y2=0
cc_115 N_A_27_508#_c_110_n N_Y_c_385_n 0.00977417f $X=0.925 $Y=2.29 $X2=0 $Y2=0
cc_116 N_A_27_508#_c_111_n N_Y_c_385_n 0.0193384f $X=1.26 $Y=1.35 $X2=0 $Y2=0
cc_117 N_A_27_508#_c_106_n N_Y_c_386_n 0.0101766f $X=1.59 $Y=1.185 $X2=0 $Y2=0
cc_118 N_A_27_508#_c_107_n N_Y_c_386_n 0.00312522f $X=1.59 $Y=1.725 $X2=0 $Y2=0
cc_119 N_A_27_508#_c_109_n N_Y_c_386_n 0.0039268f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_120 N_A_27_508#_c_111_n N_Y_c_386_n 0.00565311f $X=1.26 $Y=1.35 $X2=0 $Y2=0
cc_121 N_A_27_508#_c_108_n N_VGND_M1006_d 0.00530753f $X=0.82 $Y=0.87 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_27_508#_c_109_n N_VGND_M1006_d 6.14954e-19 $X=0.905 $Y=1.185
+ $X2=-0.19 $Y2=-0.245
cc_123 N_A_27_508#_c_106_n N_VGND_c_445_n 0.0130474f $X=1.59 $Y=1.185 $X2=0
+ $Y2=0
cc_124 N_A_27_508#_c_107_n N_VGND_c_445_n 0.00976971f $X=1.59 $Y=1.725 $X2=0
+ $Y2=0
cc_125 N_A_27_508#_c_108_n N_VGND_c_445_n 0.016103f $X=0.82 $Y=0.87 $X2=0 $Y2=0
cc_126 N_A_27_508#_c_111_n N_VGND_c_445_n 0.01063f $X=1.26 $Y=1.35 $X2=0 $Y2=0
cc_127 N_A_27_508#_c_106_n N_VGND_c_446_n 0.00486043f $X=1.59 $Y=1.185 $X2=0
+ $Y2=0
cc_128 N_A_27_508#_c_108_n N_VGND_c_450_n 0.00785591f $X=0.82 $Y=0.87 $X2=0
+ $Y2=0
cc_129 N_A_27_508#_c_106_n N_VGND_c_452_n 0.0082726f $X=1.59 $Y=1.185 $X2=0
+ $Y2=0
cc_130 N_A_27_508#_c_108_n N_VGND_c_452_n 0.0154756f $X=0.82 $Y=0.87 $X2=0 $Y2=0
cc_131 N_A_375_269#_M1011_g N_B_M1005_g 0.0529322f $X=1.95 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_375_269#_c_174_n N_B_M1005_g 0.00456423f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_133 N_A_375_269#_c_184_p N_B_M1005_g 0.0182416f $X=3.385 $Y=2.037 $X2=0 $Y2=0
cc_134 N_A_375_269#_M1001_g N_B_M1007_g 0.024764f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_135 N_A_375_269#_c_174_n N_B_c_245_n 8.70727e-19 $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_136 N_A_375_269#_c_168_n N_B_c_245_n 0.0211796f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A_375_269#_c_184_p N_B_c_245_n 9.11359e-19 $X=3.385 $Y=2.037 $X2=0
+ $Y2=0
cc_138 N_A_375_269#_c_174_n N_B_c_248_n 0.0215553f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_139 N_A_375_269#_c_168_n N_B_c_248_n 8.70727e-19 $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_140 N_A_375_269#_c_184_p N_B_c_248_n 0.0230127f $X=3.385 $Y=2.037 $X2=0 $Y2=0
cc_141 N_A_375_269#_c_184_p N_A_M1008_g 0.019789f $X=3.385 $Y=2.037 $X2=0 $Y2=0
cc_142 N_A_375_269#_c_169_n N_A_M1008_g 0.00387478f $X=3.47 $Y=1.93 $X2=0 $Y2=0
cc_143 N_A_375_269#_c_184_p A 0.0131192f $X=3.385 $Y=2.037 $X2=0 $Y2=0
cc_144 N_A_375_269#_c_169_n A 0.0373118f $X=3.47 $Y=1.93 $X2=0 $Y2=0
cc_145 N_A_375_269#_c_171_n A 0.0124961f $X=3.555 $Y=1.17 $X2=0 $Y2=0
cc_146 N_A_375_269#_c_184_p N_A_c_280_n 0.00247727f $X=3.385 $Y=2.037 $X2=0
+ $Y2=0
cc_147 N_A_375_269#_c_169_n N_A_c_280_n 0.00241564f $X=3.47 $Y=1.93 $X2=0 $Y2=0
cc_148 N_A_375_269#_c_171_n N_A_c_280_n 7.20846e-19 $X=3.555 $Y=1.17 $X2=0 $Y2=0
cc_149 N_A_375_269#_c_171_n N_A_c_281_n 5.41505e-19 $X=3.555 $Y=1.17 $X2=0 $Y2=0
cc_150 N_A_375_269#_c_169_n N_C_N_M1003_g 0.0106432f $X=3.47 $Y=1.93 $X2=0 $Y2=0
cc_151 N_A_375_269#_c_177_n N_C_N_M1003_g 0.0075316f $X=3.785 $Y=2.035 $X2=0
+ $Y2=0
cc_152 N_A_375_269#_c_203_p N_C_N_M1003_g 0.00717876f $X=3.47 $Y=2.037 $X2=0
+ $Y2=0
cc_153 N_A_375_269#_c_169_n N_C_N_M1010_g 0.00470672f $X=3.47 $Y=1.93 $X2=0
+ $Y2=0
cc_154 N_A_375_269#_c_170_n N_C_N_M1010_g 0.0161569f $X=3.92 $Y=1.17 $X2=0 $Y2=0
cc_155 N_A_375_269#_c_172_n N_C_N_M1010_g 7.53159e-19 $X=4.015 $Y=0.86 $X2=0
+ $Y2=0
cc_156 N_A_375_269#_c_169_n C_N 0.0243178f $X=3.47 $Y=1.93 $X2=0 $Y2=0
cc_157 N_A_375_269#_c_170_n C_N 0.033691f $X=3.92 $Y=1.17 $X2=0 $Y2=0
cc_158 N_A_375_269#_c_177_n C_N 0.0171153f $X=3.785 $Y=2.035 $X2=0 $Y2=0
cc_159 N_A_375_269#_c_169_n N_C_N_c_319_n 0.00553422f $X=3.47 $Y=1.93 $X2=0
+ $Y2=0
cc_160 N_A_375_269#_c_170_n N_C_N_c_319_n 0.00898108f $X=3.92 $Y=1.17 $X2=0
+ $Y2=0
cc_161 N_A_375_269#_c_177_n N_C_N_c_319_n 0.00289471f $X=3.785 $Y=2.035 $X2=0
+ $Y2=0
cc_162 N_A_375_269#_c_184_p N_VPWR_M1008_d 0.00814043f $X=3.385 $Y=2.037 $X2=0
+ $Y2=0
cc_163 N_A_375_269#_c_169_n N_VPWR_M1008_d 0.00118786f $X=3.47 $Y=1.93 $X2=0
+ $Y2=0
cc_164 N_A_375_269#_c_203_p N_VPWR_M1008_d 0.00156273f $X=3.47 $Y=2.037 $X2=0
+ $Y2=0
cc_165 N_A_375_269#_c_184_p N_VPWR_c_347_n 0.0202393f $X=3.385 $Y=2.037 $X2=0
+ $Y2=0
cc_166 N_A_375_269#_c_203_p N_VPWR_c_347_n 0.00216123f $X=3.47 $Y=2.037 $X2=0
+ $Y2=0
cc_167 N_A_375_269#_M1011_g N_VPWR_c_349_n 0.00585385f $X=1.95 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_375_269#_M1011_g N_VPWR_c_345_n 0.011101f $X=1.95 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_375_269#_M1001_g N_Y_c_384_n 0.013485f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A_375_269#_c_168_n N_Y_c_384_n 0.00272601f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_171 N_A_375_269#_c_184_p N_Y_c_384_n 0.00850133f $X=3.385 $Y=2.037 $X2=0
+ $Y2=0
cc_172 N_A_375_269#_c_171_n N_Y_c_384_n 8.40809e-19 $X=3.555 $Y=1.17 $X2=0 $Y2=0
cc_173 N_A_375_269#_M1011_g N_Y_c_388_n 0.00197296f $X=1.95 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_375_269#_M1001_g N_Y_c_385_n 0.00168714f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_175 N_A_375_269#_c_174_n N_Y_c_385_n 0.0328943f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A_375_269#_c_168_n N_Y_c_385_n 0.00197296f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A_375_269#_M1001_g N_Y_c_386_n 0.00225377f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A_375_269#_c_174_n N_Y_c_386_n 0.0257811f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A_375_269#_c_168_n N_Y_c_386_n 0.00204664f $X=2.04 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_375_269#_M1001_g N_Y_c_416_n 6.59762e-19 $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_181 N_A_375_269#_c_174_n A_405_367# 0.00121536f $X=2.04 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_375_269#_c_184_p A_405_367# 0.00955666f $X=3.385 $Y=2.037 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_375_269#_c_181_n A_405_367# 0.00554129f $X=2.205 $Y=2.037 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_375_269#_c_184_p A_513_367# 0.0163054f $X=3.385 $Y=2.037 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_375_269#_M1001_g N_VGND_c_445_n 6.52048e-19 $X=2.02 $Y=0.655 $X2=0
+ $Y2=0
cc_186 N_A_375_269#_M1001_g N_VGND_c_446_n 0.00585385f $X=2.02 $Y=0.655 $X2=0
+ $Y2=0
cc_187 N_A_375_269#_M1001_g N_VGND_c_447_n 0.00172463f $X=2.02 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A_375_269#_c_170_n N_VGND_c_449_n 0.0132473f $X=3.92 $Y=1.17 $X2=0
+ $Y2=0
cc_189 N_A_375_269#_c_171_n N_VGND_c_449_n 0.015628f $X=3.555 $Y=1.17 $X2=0
+ $Y2=0
cc_190 N_A_375_269#_c_172_n N_VGND_c_451_n 0.00391489f $X=4.015 $Y=0.86 $X2=0
+ $Y2=0
cc_191 N_A_375_269#_M1001_g N_VGND_c_452_n 0.0108326f $X=2.02 $Y=0.655 $X2=0
+ $Y2=0
cc_192 N_A_375_269#_c_172_n N_VGND_c_452_n 0.00684471f $X=4.015 $Y=0.86 $X2=0
+ $Y2=0
cc_193 N_B_M1005_g N_A_M1008_g 0.051009f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_194 N_B_c_248_n N_A_M1008_g 6.67716e-19 $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_195 N_B_M1007_g A 6.00536e-19 $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_196 N_B_c_245_n A 0.0012738f $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_197 N_B_c_248_n A 0.0165228f $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_198 N_B_c_245_n N_A_c_280_n 0.0203278f $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_199 N_B_c_248_n N_A_c_280_n 8.4048e-19 $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_200 N_B_M1007_g N_A_c_281_n 0.0192029f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_201 N_B_M1005_g N_VPWR_c_347_n 0.00449866f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B_M1005_g N_VPWR_c_349_n 0.00585385f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B_M1005_g N_VPWR_c_345_n 0.011557f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B_M1007_g N_Y_c_384_n 0.0119565f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_205 N_B_c_245_n N_Y_c_384_n 0.00484477f $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_206 N_B_c_248_n N_Y_c_384_n 0.0258896f $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_207 N_B_M1007_g N_Y_c_416_n 0.0147175f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_208 N_B_M1007_g N_VGND_c_447_n 0.00841701f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_209 N_B_M1007_g N_VGND_c_448_n 0.00473044f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_210 N_B_M1007_g N_VGND_c_449_n 0.0013481f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_211 N_B_M1007_g N_VGND_c_452_n 0.00856428f $X=2.555 $Y=0.655 $X2=0 $Y2=0
cc_212 A N_C_N_M1010_g 2.62766e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_213 N_A_c_280_n N_C_N_M1010_g 0.00674763f $X=3.12 $Y=1.35 $X2=0 $Y2=0
cc_214 N_A_c_281_n N_C_N_M1010_g 0.0039192f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_215 N_A_M1008_g N_C_N_c_319_n 0.0229798f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_216 A N_C_N_c_319_n 6.28413e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_217 N_A_M1008_g N_VPWR_c_347_n 0.0245543f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_M1008_g N_VPWR_c_349_n 0.00486043f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A_M1008_g N_VPWR_c_345_n 0.00864313f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_220 A N_Y_c_384_n 0.0121549f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A_c_281_n N_Y_c_384_n 0.00151672f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_222 N_A_c_281_n N_Y_c_416_n 0.00662676f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_223 N_A_c_281_n N_VGND_c_448_n 0.00486043f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_224 A N_VGND_c_449_n 0.00866012f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_225 N_A_c_280_n N_VGND_c_449_n 0.00337719f $X=3.12 $Y=1.35 $X2=0 $Y2=0
cc_226 N_A_c_281_n N_VGND_c_449_n 0.0157935f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_227 N_A_c_281_n N_VGND_c_452_n 0.00837755f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_228 N_C_N_M1003_g N_VPWR_c_347_n 0.00191978f $X=3.57 $Y=2.045 $X2=0 $Y2=0
cc_229 N_C_N_M1010_g N_VGND_c_449_n 0.0137526f $X=3.8 $Y=0.865 $X2=0 $Y2=0
cc_230 N_C_N_c_319_n N_VGND_c_449_n 3.63003e-19 $X=3.8 $Y=1.51 $X2=0 $Y2=0
cc_231 N_C_N_M1010_g N_VGND_c_451_n 0.00332367f $X=3.8 $Y=0.865 $X2=0 $Y2=0
cc_232 N_C_N_M1010_g N_VGND_c_452_n 0.00387424f $X=3.8 $Y=0.865 $X2=0 $Y2=0
cc_233 N_VPWR_c_345_n N_Y_M1004_s 0.00215158f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_234 N_VPWR_c_346_n N_Y_c_387_n 0.0229383f $X=0.69 $Y=2.755 $X2=0 $Y2=0
cc_235 N_VPWR_c_349_n N_Y_c_387_n 0.0306326f $X=3.08 $Y=3.33 $X2=0 $Y2=0
cc_236 N_VPWR_c_345_n N_Y_c_387_n 0.0180137f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_237 N_VPWR_c_345_n A_333_367# 0.00798529f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_238 N_VPWR_c_345_n A_405_367# 0.0167135f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_239 N_VPWR_c_345_n A_513_367# 0.0167135f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_240 N_Y_c_386_n N_VGND_c_445_n 0.00107468f $X=1.945 $Y=1.16 $X2=0 $Y2=0
cc_241 N_Y_c_429_p N_VGND_c_446_n 0.0140491f $X=1.805 $Y=0.42 $X2=0 $Y2=0
cc_242 N_Y_c_384_n N_VGND_c_447_n 0.0205451f $X=2.555 $Y=1.17 $X2=0 $Y2=0
cc_243 N_Y_c_416_n N_VGND_c_447_n 0.0500922f $X=2.77 $Y=0.42 $X2=0 $Y2=0
cc_244 N_Y_c_416_n N_VGND_c_448_n 0.0187767f $X=2.77 $Y=0.42 $X2=0 $Y2=0
cc_245 N_Y_c_416_n N_VGND_c_449_n 0.0432671f $X=2.77 $Y=0.42 $X2=0 $Y2=0
cc_246 N_Y_M1009_d N_VGND_c_452_n 0.00380103f $X=1.665 $Y=0.235 $X2=0 $Y2=0
cc_247 N_Y_M1007_d N_VGND_c_452_n 0.00607622f $X=2.63 $Y=0.235 $X2=0 $Y2=0
cc_248 N_Y_c_429_p N_VGND_c_452_n 0.0090585f $X=1.805 $Y=0.42 $X2=0 $Y2=0
cc_249 N_Y_c_416_n N_VGND_c_452_n 0.0111738f $X=2.77 $Y=0.42 $X2=0 $Y2=0
