* File: sky130_fd_sc_lp__inv_4.pex.spice
* Created: Wed Sep  2 09:55:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31 32
+ 47
r66 45 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.68 $Y=1.35 $X2=1.77
+ $Y2=1.35
r67 43 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.34 $Y=1.35
+ $X2=1.68 $Y2=1.35
r68 42 43 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.91 $Y=1.35
+ $X2=1.34 $Y2=1.35
r69 41 42 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.48 $Y=1.35
+ $X2=0.91 $Y2=1.35
r70 38 41 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.32 $Y=1.35
+ $X2=0.48 $Y2=1.35
r71 32 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.35 $X2=1.68 $Y2=1.35
r72 31 32 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.362
+ $X2=1.68 $Y2=1.362
r73 30 31 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.362
+ $X2=1.2 $Y2=1.362
r74 29 30 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.362
+ $X2=0.72 $Y2=1.362
r75 29 38 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.35 $X2=0.32 $Y2=1.35
r76 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.515
+ $X2=1.77 $Y2=1.35
r77 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.77 $Y=1.515
+ $X2=1.77 $Y2=2.465
r78 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.185
+ $X2=1.77 $Y2=1.35
r79 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.77 $Y=1.185
+ $X2=1.77 $Y2=0.655
r80 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.515
+ $X2=1.34 $Y2=1.35
r81 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.34 $Y=1.515
+ $X2=1.34 $Y2=2.465
r82 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.185
+ $X2=1.34 $Y2=1.35
r83 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.34 $Y=1.185
+ $X2=1.34 $Y2=0.655
r84 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.515
+ $X2=0.91 $Y2=1.35
r85 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.91 $Y=1.515
+ $X2=0.91 $Y2=2.465
r86 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.185
+ $X2=0.91 $Y2=1.35
r87 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.91 $Y=1.185
+ $X2=0.91 $Y2=0.655
r88 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.515
+ $X2=0.48 $Y2=1.35
r89 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.48 $Y=1.515 $X2=0.48
+ $Y2=2.465
r90 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.185
+ $X2=0.48 $Y2=1.35
r91 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.48 $Y=1.185 $X2=0.48
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__INV_4%VPWR 1 2 3 10 12 18 22 24 29 30 31 37 46
r35 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 40 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 37 45 4.21968 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=2.127 $Y2=3.33
r40 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 36 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 33 42 4.39509 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r44 33 35 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 31 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 31 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 29 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 29 30 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.122 $Y2=3.33
r49 28 39 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 28 30 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.122 $Y2=3.33
r51 24 27 26.9554 $w=2.93e-07 $l=6.9e-07 $layer=LI1_cond $X=2.002 $Y=2.26
+ $X2=2.002 $Y2=2.95
r52 22 45 3.25784 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.002 $Y=3.245
+ $X2=2.127 $Y2=3.33
r53 22 27 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=2.002 $Y=3.245
+ $X2=2.002 $Y2=2.95
r54 18 21 31.1838 $w=2.53e-07 $l=6.9e-07 $layer=LI1_cond $X=1.122 $Y=2.26
+ $X2=1.122 $Y2=2.95
r55 16 30 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.122 $Y=3.245
+ $X2=1.122 $Y2=3.33
r56 16 21 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.122 $Y=3.245
+ $X2=1.122 $Y2=2.95
r57 12 15 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=0.245 $Y=1.98
+ $X2=0.245 $Y2=2.95
r58 10 42 3.04275 $w=2.9e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.195 $Y2=3.33
r59 10 15 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.245 $Y2=2.95
r60 3 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.835 $X2=1.985 $Y2=2.95
r61 3 24 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.835 $X2=1.985 $Y2=2.26
r62 2 21 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.95
r63 2 18 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.26
r64 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.95
r65 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__INV_4%Y 1 2 3 4 15 21 23 24 25 26 29 35 37 39 41 42
+ 44 45 46 50
r57 45 46 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.162 $Y=1.295
+ $X2=2.162 $Y2=1.665
r58 45 50 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=2.162 $Y=1.295
+ $X2=2.162 $Y2=1.04
r59 44 50 2.97041 $w=2.75e-07 $l=1e-07 $layer=LI1_cond $X=2.162 $Y=0.94
+ $X2=2.162 $Y2=1.04
r60 43 46 3.77163 $w=2.73e-07 $l=9e-08 $layer=LI1_cond $X=2.162 $Y=1.755
+ $X2=2.162 $Y2=1.665
r61 40 41 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.685 $Y=1.84
+ $X2=1.552 $Y2=1.84
r62 39 43 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=2.025 $Y=1.84
+ $X2=2.162 $Y2=1.755
r63 39 40 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.025 $Y=1.84
+ $X2=1.685 $Y2=1.84
r64 38 42 6.78838 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=1.685 $Y=0.94
+ $X2=1.555 $Y2=0.94
r65 37 44 4.06946 $w=2e-07 $l=1.37e-07 $layer=LI1_cond $X=2.025 $Y=0.94
+ $X2=2.162 $Y2=0.94
r66 37 38 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.025 $Y=0.94
+ $X2=1.685 $Y2=0.94
r67 33 42 0.150961 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=1.555 $Y=0.84
+ $X2=1.555 $Y2=0.94
r68 33 35 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.555 $Y=0.84
+ $X2=1.555 $Y2=0.42
r69 29 31 40.4442 $w=2.63e-07 $l=9.3e-07 $layer=LI1_cond $X=1.552 $Y=1.98
+ $X2=1.552 $Y2=2.91
r70 27 41 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.552 $Y=1.925
+ $X2=1.552 $Y2=1.84
r71 27 29 2.39186 $w=2.63e-07 $l=5.5e-08 $layer=LI1_cond $X=1.552 $Y=1.925
+ $X2=1.552 $Y2=1.98
r72 25 41 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.42 $Y=1.84
+ $X2=1.552 $Y2=1.84
r73 25 26 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.42 $Y=1.84
+ $X2=0.825 $Y2=1.84
r74 23 42 6.78838 $w=1.85e-07 $l=1.37295e-07 $layer=LI1_cond $X=1.425 $Y=0.955
+ $X2=1.555 $Y2=0.94
r75 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.425 $Y=0.955
+ $X2=0.825 $Y2=0.955
r76 19 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.695 $Y=0.87
+ $X2=0.825 $Y2=0.955
r77 19 21 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=0.695 $Y=0.87
+ $X2=0.695 $Y2=0.42
r78 15 17 40.4442 $w=2.63e-07 $l=9.3e-07 $layer=LI1_cond $X=0.692 $Y=1.98
+ $X2=0.692 $Y2=2.91
r79 13 26 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.692 $Y=1.925
+ $X2=0.825 $Y2=1.84
r80 13 15 2.39186 $w=2.63e-07 $l=5.5e-08 $layer=LI1_cond $X=0.692 $Y=1.925
+ $X2=0.692 $Y2=1.98
r81 4 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.415
+ $Y=1.835 $X2=1.555 $Y2=2.91
r82 4 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.415
+ $Y=1.835 $X2=1.555 $Y2=1.98
r83 3 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.91
r84 3 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=1.98
r85 2 35 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.42
r86 1 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=0.695 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__INV_4%VGND 1 2 3 10 12 16 18 20 23 24 25 31 40
r38 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 34 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r41 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r42 31 39 4.21968 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.127
+ $Y2=0
r43 31 33 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.68
+ $Y2=0
r44 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r45 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 27 36 4.4461 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r47 27 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.72
+ $Y2=0
r48 25 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r49 25 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r50 23 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.72
+ $Y2=0
r51 23 24 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.125
+ $Y2=0
r52 22 33 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.68
+ $Y2=0
r53 22 24 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.125
+ $Y2=0
r54 18 39 3.25784 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.002 $Y=0.085
+ $X2=2.127 $Y2=0
r55 18 20 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=2.002 $Y=0.085
+ $X2=2.002 $Y2=0.505
r56 14 24 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0
r57 14 16 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0.535
r58 10 36 3.03143 $w=2.95e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.247 $Y=0.085
+ $X2=0.197 $Y2=0
r59 10 12 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.247 $Y=0.085
+ $X2=0.247 $Y2=0.38
r60 3 20 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=1.985 $Y2=0.505
r61 2 16 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.125 $Y2=0.535
r62 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.38
.ends

