* File: sky130_fd_sc_lp__and3_4.pex.spice
* Created: Wed Sep  2 09:31:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3_4%A 3 6 8 9 13 15
r27 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=1.35
+ $X2=0.635 $Y2=1.515
r28 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=1.35
+ $X2=0.635 $Y2=1.185
r29 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=1.35 $X2=0.635 $Y2=1.35
r30 8 9 14.9251 $w=3.03e-07 $l=3.95e-07 $layer=LI1_cond $X=0.24 $Y=1.362
+ $X2=0.635 $Y2=1.362
r31 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.725 $Y=2.465
+ $X2=0.725 $Y2=1.515
r32 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.725 $Y=0.655
+ $X2=0.725 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_4%B 3 7 9 12
c29 7 0 4.04067e-20 $X=1.235 $Y=2.465
r30 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.375
+ $X2=1.175 $Y2=1.54
r31 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.375
+ $X2=1.175 $Y2=1.21
r32 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=1.375 $X2=1.175 $Y2=1.375
r33 7 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.235 $Y=2.465
+ $X2=1.235 $Y2=1.54
r34 3 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.085 $Y=0.655
+ $X2=1.085 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_4%C 3 7 9 12
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.375
+ $X2=1.715 $Y2=1.54
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.375
+ $X2=1.715 $Y2=1.21
r36 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.715
+ $Y=1.375 $X2=1.715 $Y2=1.375
r37 7 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.665 $Y=2.465
+ $X2=1.665 $Y2=1.54
r38 3 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.625 $Y=0.655
+ $X2=1.625 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_4%A_77_47# 1 2 3 12 16 20 24 28 32 36 40 44 48
+ 52 53 54 55 58 62 65 71 72 74 75
c137 75 0 4.04067e-20 $X=2.065 $Y=1.5
r138 82 83 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.06 $Y=1.5
+ $X2=3.49 $Y2=1.5
r139 81 82 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.63 $Y=1.5
+ $X2=3.06 $Y2=1.5
r140 75 76 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.065 $Y=1.5
+ $X2=2.065 $Y2=1.795
r141 72 83 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.65 $Y=1.5
+ $X2=3.49 $Y2=1.5
r142 71 72 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.65
+ $Y=1.5 $X2=3.65 $Y2=1.5
r143 69 81 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.29 $Y=1.5
+ $X2=2.63 $Y2=1.5
r144 69 78 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.29 $Y=1.5 $X2=2.2
+ $Y2=1.5
r145 68 71 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.29 $Y=1.5
+ $X2=3.65 $Y2=1.5
r146 68 69 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.5 $X2=2.29 $Y2=1.5
r147 66 75 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=1.5
+ $X2=2.065 $Y2=1.5
r148 66 68 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.15 $Y=1.5
+ $X2=2.29 $Y2=1.5
r149 65 75 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=1.415
+ $X2=2.065 $Y2=1.5
r150 64 65 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.065 $Y=1.04
+ $X2=2.065 $Y2=1.415
r151 63 74 6.28297 $w=1.92e-07 $l=1.33548e-07 $layer=LI1_cond $X=1.595 $Y=1.795
+ $X2=1.472 $Y2=1.817
r152 62 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.795
+ $X2=2.065 $Y2=1.795
r153 62 63 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.98 $Y=1.795
+ $X2=1.595 $Y2=1.795
r154 58 60 43.7458 $w=2.43e-07 $l=9.3e-07 $layer=LI1_cond $X=1.472 $Y=1.98
+ $X2=1.472 $Y2=2.91
r155 56 74 0.490351 $w=2.45e-07 $l=1.08e-07 $layer=LI1_cond $X=1.472 $Y=1.925
+ $X2=1.472 $Y2=1.817
r156 56 58 2.58712 $w=2.43e-07 $l=5.5e-08 $layer=LI1_cond $X=1.472 $Y=1.925
+ $X2=1.472 $Y2=1.98
r157 54 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.98 $Y=0.955
+ $X2=2.065 $Y2=1.04
r158 54 55 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=1.98 $Y=0.955
+ $X2=0.675 $Y2=0.955
r159 52 74 6.28297 $w=1.92e-07 $l=1.22e-07 $layer=LI1_cond $X=1.35 $Y=1.817
+ $X2=1.472 $Y2=1.817
r160 52 53 39.3975 $w=2.13e-07 $l=7.35e-07 $layer=LI1_cond $X=1.35 $Y=1.817
+ $X2=0.615 $Y2=1.817
r161 48 50 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.48 $Y=1.98
+ $X2=0.48 $Y2=2.91
r162 46 53 6.93113 $w=2.15e-07 $l=1.81122e-07 $layer=LI1_cond $X=0.48 $Y=1.925
+ $X2=0.615 $Y2=1.817
r163 46 48 2.34757 $w=2.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.48 $Y=1.925
+ $X2=0.48 $Y2=1.98
r164 42 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.51 $Y=0.87
+ $X2=0.675 $Y2=0.955
r165 42 44 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.51 $Y=0.87
+ $X2=0.51 $Y2=0.38
r166 38 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.665
+ $X2=3.49 $Y2=1.5
r167 38 40 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.49 $Y=1.665
+ $X2=3.49 $Y2=2.465
r168 34 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.335
+ $X2=3.49 $Y2=1.5
r169 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.49 $Y=1.335
+ $X2=3.49 $Y2=0.655
r170 30 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.665
+ $X2=3.06 $Y2=1.5
r171 30 32 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.06 $Y=1.665
+ $X2=3.06 $Y2=2.465
r172 26 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.335
+ $X2=3.06 $Y2=1.5
r173 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.06 $Y=1.335
+ $X2=3.06 $Y2=0.655
r174 22 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.665
+ $X2=2.63 $Y2=1.5
r175 22 24 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.63 $Y=1.665
+ $X2=2.63 $Y2=2.465
r176 18 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.335
+ $X2=2.63 $Y2=1.5
r177 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.63 $Y=1.335
+ $X2=2.63 $Y2=0.655
r178 14 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.665
+ $X2=2.2 $Y2=1.5
r179 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=2.465
r180 10 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.335
+ $X2=2.2 $Y2=1.5
r181 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.2 $Y=1.335
+ $X2=2.2 $Y2=0.655
r182 3 60 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.835 $X2=1.45 $Y2=2.91
r183 3 58 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.835 $X2=1.45 $Y2=1.98
r184 2 50 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.835 $X2=0.51 $Y2=2.91
r185 2 48 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.835 $X2=0.51 $Y2=1.98
r186 1 44 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.385
+ $Y=0.235 $X2=0.51 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_4%VPWR 1 2 3 4 15 21 27 31 35 40 41 43 44 45 46
+ 47 61 62 65
r61 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 59 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=3.705 $Y2=3.33
r65 59 61 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 58 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 47 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 47 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 45 57 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r74 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=2.845 $Y2=3.33
r75 43 54 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.93 $Y2=3.33
r77 42 57 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.93 $Y2=3.33
r79 40 50 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.98 $Y2=3.33
r81 39 54 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=0.98 $Y2=3.33
r83 35 38 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.705 $Y=2.18
+ $X2=3.705 $Y2=2.95
r84 33 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=3.245
+ $X2=3.705 $Y2=3.33
r85 33 38 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.705 $Y=3.245
+ $X2=3.705 $Y2=2.95
r86 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=2.845 $Y2=3.33
r87 31 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=3.705 $Y2=3.33
r88 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=3.01 $Y2=3.33
r89 27 30 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.845 $Y=2.18
+ $X2=2.845 $Y2=2.97
r90 25 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=3.245
+ $X2=2.845 $Y2=3.33
r91 25 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.845 $Y=3.245
+ $X2=2.845 $Y2=2.97
r92 21 24 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=1.93 $Y=2.135
+ $X2=1.93 $Y2=2.95
r93 19 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r94 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.95
r95 15 18 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.98 $Y=2.19
+ $X2=0.98 $Y2=2.95
r96 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.98 $Y=3.245
+ $X2=0.98 $Y2=3.33
r97 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.98 $Y=3.245
+ $X2=0.98 $Y2=2.95
r98 4 38 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.835 $X2=3.705 $Y2=2.95
r99 4 35 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.835 $X2=3.705 $Y2=2.18
r100 3 30 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.845 $Y2=2.97
r101 3 27 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.845 $Y2=2.18
r102 2 24 400 $w=1.7e-07 $l=1.20626e-06 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.835 $X2=1.93 $Y2=2.95
r103 2 21 400 $w=1.7e-07 $l=3.83406e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.835 $X2=1.93 $Y2=2.135
r104 1 18 400 $w=1.7e-07 $l=1.20163e-06 $layer=licon1_PDIFF $count=1 $X=0.8
+ $Y=1.835 $X2=0.98 $Y2=2.95
r105 1 15 400 $w=1.7e-07 $l=4.35804e-07 $layer=licon1_PDIFF $count=1 $X=0.8
+ $Y=1.835 $X2=0.98 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 40 41 43
+ 44 45 46 61
r65 59 61 3.00637 $w=2.28e-07 $l=6e-08 $layer=LI1_cond $X=4.11 $Y=1.235 $X2=4.11
+ $Y2=1.295
r66 45 53 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=1.15 $X2=4.11
+ $Y2=1.065
r67 45 59 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=1.15 $X2=4.11
+ $Y2=1.235
r68 45 46 17.938 $w=2.28e-07 $l=3.58e-07 $layer=LI1_cond $X=4.11 $Y=1.307
+ $X2=4.11 $Y2=1.665
r69 45 61 0.601275 $w=2.28e-07 $l=1.2e-08 $layer=LI1_cond $X=4.11 $Y=1.307
+ $X2=4.11 $Y2=1.295
r70 44 53 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.11 $Y=0.925
+ $X2=4.11 $Y2=1.065
r71 43 44 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.11 $Y=0.555
+ $X2=4.11 $Y2=0.925
r72 42 46 4.50956 $w=2.28e-07 $l=9e-08 $layer=LI1_cond $X=4.11 $Y=1.755 $X2=4.11
+ $Y2=1.665
r73 39 45 35.7594 $w=1.93e-07 $l=6.25e-07 $layer=LI1_cond $X=3.37 $Y=1.15
+ $X2=3.995 $Y2=1.15
r74 39 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.37 $Y=1.15
+ $X2=3.275 $Y2=1.15
r75 38 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.37 $Y=1.84
+ $X2=3.275 $Y2=1.84
r76 37 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.995 $Y=1.84
+ $X2=4.11 $Y2=1.755
r77 37 38 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.995 $Y=1.84
+ $X2=3.37 $Y2=1.84
r78 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.275 $Y=1.98
+ $X2=3.275 $Y2=2.91
r79 31 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=1.925
+ $X2=3.275 $Y2=1.84
r80 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=3.275 $Y=1.925
+ $X2=3.275 $Y2=1.98
r81 27 40 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=1.065
+ $X2=3.275 $Y2=1.15
r82 27 29 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=3.275 $Y=1.065
+ $X2=3.275 $Y2=0.42
r83 25 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.18 $Y=1.84
+ $X2=3.275 $Y2=1.84
r84 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.18 $Y=1.84
+ $X2=2.51 $Y2=1.84
r85 23 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.18 $Y=1.15
+ $X2=3.275 $Y2=1.15
r86 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.18 $Y=1.15
+ $X2=2.51 $Y2=1.15
r87 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.415 $Y=1.98
+ $X2=2.415 $Y2=2.91
r88 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.415 $Y=1.925
+ $X2=2.51 $Y2=1.84
r89 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=2.415 $Y=1.925
+ $X2=2.415 $Y2=1.98
r90 13 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.415 $Y=1.065
+ $X2=2.51 $Y2=1.15
r91 13 15 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=2.415 $Y=1.065
+ $X2=2.415 $Y2=0.42
r92 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.135
+ $Y=1.835 $X2=3.275 $Y2=2.91
r93 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.135
+ $Y=1.835 $X2=3.275 $Y2=1.98
r94 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=2.91
r95 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=1.98
r96 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.135
+ $Y=0.235 $X2=3.275 $Y2=0.42
r97 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.275
+ $Y=0.235 $X2=2.415 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_4%VGND 1 2 3 12 16 18 22 25 26 27 28 29 43 44
+ 47
r54 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 44 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r56 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 41 47 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.682
+ $Y2=0
r58 41 43 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=4.08
+ $Y2=0
r59 40 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r60 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r61 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r62 33 37 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r63 32 36 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r64 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r66 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r67 27 39 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.64
+ $Y2=0
r68 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.845
+ $Y2=0
r69 25 36 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.68
+ $Y2=0
r70 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.91
+ $Y2=0
r71 24 39 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.64
+ $Y2=0
r72 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=1.91
+ $Y2=0
r73 20 47 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.682 $Y=0.085
+ $X2=3.682 $Y2=0
r74 20 22 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=3.682 $Y=0.085
+ $X2=3.682 $Y2=0.38
r75 19 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.845
+ $Y2=0
r76 18 47 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.682
+ $Y2=0
r77 18 19 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.01
+ $Y2=0
r78 14 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0
r79 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0.38
r80 10 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=0.085
+ $X2=1.91 $Y2=0
r81 10 12 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.91 $Y=0.085
+ $X2=1.91 $Y2=0.56
r82 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.565
+ $Y=0.235 $X2=3.705 $Y2=0.38
r83 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.705
+ $Y=0.235 $X2=2.845 $Y2=0.38
r84 1 12 182 $w=1.7e-07 $l=4.16983e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=1.91 $Y2=0.56
.ends

