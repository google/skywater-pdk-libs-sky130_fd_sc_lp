* File: sky130_fd_sc_lp__bufinv_16.pex.spice
* Created: Fri Aug 28 10:11:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFINV_16%A 3 7 11 15 19 23 25 26 27 31 43 44
c60 43 0 9.89959e-20 $X=1.405 $Y=1.51
r61 42 44 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.405 $Y=1.51
+ $X2=1.515 $Y2=1.51
r62 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=1.51 $X2=1.405 $Y2=1.51
r63 40 42 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.085 $Y=1.51
+ $X2=1.405 $Y2=1.51
r64 38 40 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.065 $Y=1.51
+ $X2=1.085 $Y2=1.51
r65 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=1.51 $X2=1.065 $Y2=1.51
r66 36 38 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.655 $Y=1.51
+ $X2=1.065 $Y2=1.51
r67 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.51 $X2=0.385 $Y2=1.51
r68 31 36 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.58 $Y=1.51
+ $X2=0.655 $Y2=1.51
r69 31 33 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.58 $Y=1.51
+ $X2=0.385 $Y2=1.51
r70 27 43 6.84785 $w=3.43e-07 $l=2.05e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.405 $Y2=1.587
r71 27 39 4.50956 $w=3.43e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.065 $Y2=1.587
r72 26 39 11.5244 $w=3.43e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=1.065 $Y2=1.587
r73 26 34 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=0.385 $Y2=1.587
r74 25 34 4.8436 $w=3.43e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.587
+ $X2=0.385 $Y2=1.587
r75 21 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.675
+ $X2=1.515 $Y2=1.51
r76 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.515 $Y=1.675
+ $X2=1.515 $Y2=2.465
r77 17 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.345
+ $X2=1.515 $Y2=1.51
r78 17 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.515 $Y=1.345
+ $X2=1.515 $Y2=0.665
r79 13 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.675
+ $X2=1.085 $Y2=1.51
r80 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.085 $Y=1.675
+ $X2=1.085 $Y2=2.465
r81 9 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.345
+ $X2=1.085 $Y2=1.51
r82 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.085 $Y=1.345
+ $X2=1.085 $Y2=0.665
r83 5 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.675
+ $X2=0.655 $Y2=1.51
r84 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.655 $Y=1.675
+ $X2=0.655 $Y2=2.465
r85 1 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.345
+ $X2=0.655 $Y2=1.51
r86 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.655 $Y=1.345
+ $X2=0.655 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_16%A_63_49# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 65 67 69 70 71 75 79 81 83 86 88 94 99 101 102 111
c158 94 0 1.68532e-19 $X=4.005 $Y=1.49
c159 19 0 9.89959e-20 $X=1.99 $Y=2.465
r160 108 109 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.28 $Y=1.49
+ $X2=3.71 $Y2=1.49
r161 107 108 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.85 $Y=1.49
+ $X2=3.28 $Y2=1.49
r162 106 107 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.42 $Y=1.49
+ $X2=2.85 $Y2=1.49
r163 105 106 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.99 $Y=1.49
+ $X2=2.42 $Y2=1.49
r164 95 111 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.005 $Y=1.49
+ $X2=4.14 $Y2=1.49
r165 95 109 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=4.005 $Y=1.49
+ $X2=3.71 $Y2=1.49
r166 94 95 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=4.005
+ $Y=1.49 $X2=4.005 $Y2=1.49
r167 92 105 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.965 $Y=1.49
+ $X2=1.99 $Y2=1.49
r168 91 94 119.081 $w=1.88e-07 $l=2.04e-06 $layer=LI1_cond $X=1.965 $Y=1.49
+ $X2=4.005 $Y2=1.49
r169 91 92 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=1.965
+ $Y=1.49 $X2=1.965 $Y2=1.49
r170 89 102 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=1.49
+ $X2=1.835 $Y2=1.49
r171 89 91 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=1.92 $Y=1.49
+ $X2=1.965 $Y2=1.49
r172 87 102 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.835 $Y=1.585
+ $X2=1.835 $Y2=1.49
r173 87 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.835 $Y=1.585
+ $X2=1.835 $Y2=1.93
r174 86 102 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.835 $Y=1.395
+ $X2=1.835 $Y2=1.49
r175 85 86 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.835 $Y=1.245
+ $X2=1.835 $Y2=1.395
r176 84 101 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.43 $Y=2.015
+ $X2=1.3 $Y2=2.015
r177 83 88 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.75 $Y=2.015
+ $X2=1.835 $Y2=1.93
r178 83 84 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.75 $Y=2.015
+ $X2=1.43 $Y2=2.015
r179 82 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.43 $Y=1.16 $X2=1.3
+ $Y2=1.16
r180 81 85 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.75 $Y=1.16
+ $X2=1.835 $Y2=1.245
r181 81 82 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.75 $Y=1.16
+ $X2=1.43 $Y2=1.16
r182 77 101 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.1 $X2=1.3
+ $Y2=2.015
r183 77 79 33.6868 $w=2.58e-07 $l=7.6e-07 $layer=LI1_cond $X=1.3 $Y=2.1 $X2=1.3
+ $Y2=2.86
r184 73 99 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=1.075
+ $X2=1.3 $Y2=1.16
r185 73 75 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=1.3 $Y=1.075
+ $X2=1.3 $Y2=0.48
r186 72 98 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.57 $Y=2.015
+ $X2=0.422 $Y2=2.015
r187 71 101 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.17 $Y=2.015
+ $X2=1.3 $Y2=2.015
r188 71 72 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.17 $Y=2.015
+ $X2=0.57 $Y2=2.015
r189 69 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.17 $Y=1.16 $X2=1.3
+ $Y2=1.16
r190 69 70 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.17 $Y=1.16 $X2=0.57
+ $Y2=1.16
r191 65 98 2.72785 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.422 $Y=2.1
+ $X2=0.422 $Y2=2.015
r192 65 67 29.6901 $w=2.93e-07 $l=7.6e-07 $layer=LI1_cond $X=0.422 $Y=2.1
+ $X2=0.422 $Y2=2.86
r193 61 70 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.422 $Y=1.075
+ $X2=0.57 $Y2=1.16
r194 61 63 23.2442 $w=2.93e-07 $l=5.95e-07 $layer=LI1_cond $X=0.422 $Y=1.075
+ $X2=0.422 $Y2=0.48
r195 57 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.655
+ $X2=4.14 $Y2=1.49
r196 57 59 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.14 $Y=1.655
+ $X2=4.14 $Y2=2.465
r197 53 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.325
+ $X2=4.14 $Y2=1.49
r198 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.14 $Y=1.325
+ $X2=4.14 $Y2=0.665
r199 49 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.655
+ $X2=3.71 $Y2=1.49
r200 49 51 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.71 $Y=1.655
+ $X2=3.71 $Y2=2.465
r201 45 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.325
+ $X2=3.71 $Y2=1.49
r202 45 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.71 $Y=1.325
+ $X2=3.71 $Y2=0.665
r203 41 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.28 $Y=1.655
+ $X2=3.28 $Y2=1.49
r204 41 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.28 $Y=1.655
+ $X2=3.28 $Y2=2.465
r205 37 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.28 $Y=1.325
+ $X2=3.28 $Y2=1.49
r206 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.28 $Y=1.325
+ $X2=3.28 $Y2=0.665
r207 33 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.655
+ $X2=2.85 $Y2=1.49
r208 33 35 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.85 $Y=1.655
+ $X2=2.85 $Y2=2.465
r209 29 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.325
+ $X2=2.85 $Y2=1.49
r210 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.85 $Y=1.325
+ $X2=2.85 $Y2=0.665
r211 25 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.655
+ $X2=2.42 $Y2=1.49
r212 25 27 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.42 $Y=1.655
+ $X2=2.42 $Y2=2.465
r213 21 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.325
+ $X2=2.42 $Y2=1.49
r214 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.42 $Y=1.325
+ $X2=2.42 $Y2=0.665
r215 17 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.655
+ $X2=1.99 $Y2=1.49
r216 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.99 $Y=1.655
+ $X2=1.99 $Y2=2.465
r217 13 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.325
+ $X2=1.99 $Y2=1.49
r218 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.99 $Y=1.325
+ $X2=1.99 $Y2=0.665
r219 4 101 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.835 $X2=1.3 $Y2=2.095
r220 4 79 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.835 $X2=1.3 $Y2=2.86
r221 3 98 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=1.835 $X2=0.44 $Y2=2.095
r222 3 67 400 $w=1.7e-07 $l=1.0857e-06 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=1.835 $X2=0.44 $Y2=2.86
r223 2 75 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=1.16
+ $Y=0.245 $X2=1.3 $Y2=0.48
r224 1 63 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=0.315
+ $Y=0.245 $X2=0.44 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_16%A_413_49# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 153 157 158 159 160 163 167 171 173 177 181 185 187 189 190 191
+ 192 197 218 226 231 236 241 246 251 256 258
c366 258 0 1.68532e-19 $X=11.02 $Y=1.51
c367 187 0 1.57775e-19 $X=4.34 $Y=1.84
r368 257 258 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=10.59 $Y=1.51
+ $X2=11.02 $Y2=1.51
r369 255 257 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=10.375 $Y=1.51
+ $X2=10.59 $Y2=1.51
r370 255 256 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.375
+ $Y=1.51 $X2=10.375 $Y2=1.51
r371 253 255 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=10.16 $Y=1.51
+ $X2=10.375 $Y2=1.51
r372 252 253 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=9.73 $Y=1.51
+ $X2=10.16 $Y2=1.51
r373 250 252 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=9.515 $Y=1.51
+ $X2=9.73 $Y2=1.51
r374 250 251 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.515
+ $Y=1.51 $X2=9.515 $Y2=1.51
r375 248 250 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=9.3 $Y=1.51
+ $X2=9.515 $Y2=1.51
r376 247 248 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.87 $Y=1.51
+ $X2=9.3 $Y2=1.51
r377 245 247 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.655 $Y=1.51
+ $X2=8.87 $Y2=1.51
r378 245 246 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.655
+ $Y=1.51 $X2=8.655 $Y2=1.51
r379 243 245 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.44 $Y=1.51
+ $X2=8.655 $Y2=1.51
r380 242 243 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.01 $Y=1.51
+ $X2=8.44 $Y2=1.51
r381 240 242 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.795 $Y=1.51
+ $X2=8.01 $Y2=1.51
r382 240 241 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.795
+ $Y=1.51 $X2=7.795 $Y2=1.51
r383 238 240 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.58 $Y=1.51
+ $X2=7.795 $Y2=1.51
r384 237 238 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.15 $Y=1.51
+ $X2=7.58 $Y2=1.51
r385 235 237 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.935 $Y=1.51
+ $X2=7.15 $Y2=1.51
r386 235 236 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.935
+ $Y=1.51 $X2=6.935 $Y2=1.51
r387 233 235 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.72 $Y=1.51
+ $X2=6.935 $Y2=1.51
r388 232 233 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.29 $Y=1.51
+ $X2=6.72 $Y2=1.51
r389 230 232 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.075 $Y=1.51
+ $X2=6.29 $Y2=1.51
r390 230 231 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.075
+ $Y=1.51 $X2=6.075 $Y2=1.51
r391 228 230 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.86 $Y=1.51
+ $X2=6.075 $Y2=1.51
r392 227 228 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.43 $Y=1.51
+ $X2=5.86 $Y2=1.51
r393 225 227 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.215 $Y=1.51
+ $X2=5.43 $Y2=1.51
r394 225 226 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.215
+ $Y=1.51 $X2=5.215 $Y2=1.51
r395 223 225 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5 $Y=1.51
+ $X2=5.215 $Y2=1.51
r396 221 223 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.57 $Y=1.51
+ $X2=5 $Y2=1.51
r397 218 256 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.375 $Y=1.665
+ $X2=10.375 $Y2=1.665
r398 215 218 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.515 $Y=1.665
+ $X2=10.375 $Y2=1.665
r399 215 251 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.515 $Y=1.665
+ $X2=9.515 $Y2=1.665
r400 212 215 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=8.655 $Y=1.665
+ $X2=9.515 $Y2=1.665
r401 212 246 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.655 $Y=1.665
+ $X2=8.655 $Y2=1.665
r402 209 212 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.795 $Y=1.665
+ $X2=8.655 $Y2=1.665
r403 209 241 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.795 $Y=1.665
+ $X2=7.795 $Y2=1.665
r404 206 209 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.935 $Y=1.665
+ $X2=7.795 $Y2=1.665
r405 206 236 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.935 $Y=1.665
+ $X2=6.935 $Y2=1.665
r406 203 206 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.075 $Y=1.665
+ $X2=6.935 $Y2=1.665
r407 203 231 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.075 $Y=1.665
+ $X2=6.075 $Y2=1.665
r408 200 203 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.215 $Y=1.665
+ $X2=6.075 $Y2=1.665
r409 200 226 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.215 $Y=1.665
+ $X2=5.215 $Y2=1.665
r410 196 200 0.500451 $w=2.3e-07 $l=7.8e-07 $layer=MET1_cond $X=4.435 $Y=1.665
+ $X2=5.215 $Y2=1.665
r411 196 197 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.435 $Y=1.665
+ $X2=4.435 $Y2=1.665
r412 194 197 5.54545 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=4.43 $Y=1.755
+ $X2=4.43 $Y2=1.665
r413 193 197 27.1111 $w=1.78e-07 $l=4.4e-07 $layer=LI1_cond $X=4.43 $Y=1.225
+ $X2=4.43 $Y2=1.665
r414 188 192 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.055 $Y=1.84
+ $X2=3.925 $Y2=1.84
r415 187 194 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.34 $Y=1.84
+ $X2=4.43 $Y2=1.755
r416 187 188 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.34 $Y=1.84
+ $X2=4.055 $Y2=1.84
r417 186 191 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.055 $Y=1.14
+ $X2=3.925 $Y2=1.14
r418 185 193 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.34 $Y=1.14
+ $X2=4.43 $Y2=1.225
r419 185 186 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.34 $Y=1.14
+ $X2=4.055 $Y2=1.14
r420 181 183 33.9084 $w=2.58e-07 $l=7.65e-07 $layer=LI1_cond $X=3.925 $Y=2.095
+ $X2=3.925 $Y2=2.86
r421 179 192 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=1.925
+ $X2=3.925 $Y2=1.84
r422 179 181 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=3.925 $Y=1.925
+ $X2=3.925 $Y2=2.095
r423 175 191 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=1.055
+ $X2=3.925 $Y2=1.14
r424 175 177 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.925 $Y=1.055
+ $X2=3.925 $Y2=0.48
r425 174 190 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.195 $Y=1.84
+ $X2=3.065 $Y2=1.84
r426 173 192 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.795 $Y=1.84
+ $X2=3.925 $Y2=1.84
r427 173 174 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.795 $Y=1.84
+ $X2=3.195 $Y2=1.84
r428 172 189 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.195 $Y=1.14
+ $X2=3.065 $Y2=1.14
r429 171 191 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.795 $Y=1.14
+ $X2=3.925 $Y2=1.14
r430 171 172 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.795 $Y=1.14
+ $X2=3.195 $Y2=1.14
r431 167 169 33.9084 $w=2.58e-07 $l=7.65e-07 $layer=LI1_cond $X=3.065 $Y=2.095
+ $X2=3.065 $Y2=2.86
r432 165 190 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=1.925
+ $X2=3.065 $Y2=1.84
r433 165 167 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=3.065 $Y=1.925
+ $X2=3.065 $Y2=2.095
r434 161 189 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=1.055
+ $X2=3.065 $Y2=1.14
r435 161 163 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.065 $Y=1.055
+ $X2=3.065 $Y2=0.48
r436 159 190 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.935 $Y=1.84
+ $X2=3.065 $Y2=1.84
r437 159 160 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.935 $Y=1.84
+ $X2=2.335 $Y2=1.84
r438 157 189 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.935 $Y=1.14
+ $X2=3.065 $Y2=1.14
r439 157 158 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.935 $Y=1.14
+ $X2=2.335 $Y2=1.14
r440 153 155 35.9844 $w=2.43e-07 $l=7.65e-07 $layer=LI1_cond $X=2.212 $Y=2.095
+ $X2=2.212 $Y2=2.86
r441 151 160 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=2.212 $Y=1.925
+ $X2=2.335 $Y2=1.84
r442 151 153 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=2.212 $Y=1.925
+ $X2=2.212 $Y2=2.095
r443 147 158 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=2.212 $Y=1.055
+ $X2=2.335 $Y2=1.14
r444 147 149 27.0471 $w=2.43e-07 $l=5.75e-07 $layer=LI1_cond $X=2.212 $Y=1.055
+ $X2=2.212 $Y2=0.48
r445 143 258 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.02 $Y=1.675
+ $X2=11.02 $Y2=1.51
r446 143 145 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.02 $Y=1.675
+ $X2=11.02 $Y2=2.465
r447 139 258 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.02 $Y=1.345
+ $X2=11.02 $Y2=1.51
r448 139 141 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=11.02 $Y=1.345
+ $X2=11.02 $Y2=0.665
r449 135 257 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.59 $Y=1.675
+ $X2=10.59 $Y2=1.51
r450 135 137 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.59 $Y=1.675
+ $X2=10.59 $Y2=2.465
r451 131 257 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.59 $Y=1.345
+ $X2=10.59 $Y2=1.51
r452 131 133 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.59 $Y=1.345
+ $X2=10.59 $Y2=0.665
r453 127 253 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.16 $Y=1.675
+ $X2=10.16 $Y2=1.51
r454 127 129 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.16 $Y=1.675
+ $X2=10.16 $Y2=2.465
r455 123 253 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.16 $Y=1.345
+ $X2=10.16 $Y2=1.51
r456 123 125 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.16 $Y=1.345
+ $X2=10.16 $Y2=0.665
r457 119 252 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.73 $Y=1.675
+ $X2=9.73 $Y2=1.51
r458 119 121 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.73 $Y=1.675
+ $X2=9.73 $Y2=2.465
r459 115 252 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.73 $Y=1.345
+ $X2=9.73 $Y2=1.51
r460 115 117 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.73 $Y=1.345
+ $X2=9.73 $Y2=0.665
r461 111 248 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.3 $Y=1.675
+ $X2=9.3 $Y2=1.51
r462 111 113 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.3 $Y=1.675
+ $X2=9.3 $Y2=2.465
r463 107 248 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.3 $Y=1.345
+ $X2=9.3 $Y2=1.51
r464 107 109 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.3 $Y=1.345
+ $X2=9.3 $Y2=0.665
r465 103 247 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.87 $Y=1.675
+ $X2=8.87 $Y2=1.51
r466 103 105 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.87 $Y=1.675
+ $X2=8.87 $Y2=2.465
r467 99 247 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.87 $Y=1.345
+ $X2=8.87 $Y2=1.51
r468 99 101 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.87 $Y=1.345
+ $X2=8.87 $Y2=0.665
r469 95 243 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.44 $Y=1.675
+ $X2=8.44 $Y2=1.51
r470 95 97 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.44 $Y=1.675
+ $X2=8.44 $Y2=2.465
r471 91 243 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.44 $Y=1.345
+ $X2=8.44 $Y2=1.51
r472 91 93 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.44 $Y=1.345
+ $X2=8.44 $Y2=0.665
r473 87 242 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.01 $Y=1.675
+ $X2=8.01 $Y2=1.51
r474 87 89 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.01 $Y=1.675
+ $X2=8.01 $Y2=2.465
r475 83 242 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.01 $Y=1.345
+ $X2=8.01 $Y2=1.51
r476 83 85 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.01 $Y=1.345
+ $X2=8.01 $Y2=0.665
r477 79 238 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.58 $Y=1.675
+ $X2=7.58 $Y2=1.51
r478 79 81 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.58 $Y=1.675
+ $X2=7.58 $Y2=2.465
r479 75 238 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.58 $Y=1.345
+ $X2=7.58 $Y2=1.51
r480 75 77 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.58 $Y=1.345
+ $X2=7.58 $Y2=0.665
r481 71 237 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.15 $Y=1.675
+ $X2=7.15 $Y2=1.51
r482 71 73 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.15 $Y=1.675
+ $X2=7.15 $Y2=2.465
r483 67 237 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.15 $Y=1.345
+ $X2=7.15 $Y2=1.51
r484 67 69 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.15 $Y=1.345
+ $X2=7.15 $Y2=0.665
r485 63 233 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.72 $Y=1.675
+ $X2=6.72 $Y2=1.51
r486 63 65 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.72 $Y=1.675
+ $X2=6.72 $Y2=2.465
r487 59 233 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.72 $Y=1.345
+ $X2=6.72 $Y2=1.51
r488 59 61 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.72 $Y=1.345
+ $X2=6.72 $Y2=0.665
r489 55 232 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.29 $Y=1.675
+ $X2=6.29 $Y2=1.51
r490 55 57 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.29 $Y=1.675
+ $X2=6.29 $Y2=2.465
r491 51 232 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.29 $Y=1.345
+ $X2=6.29 $Y2=1.51
r492 51 53 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.29 $Y=1.345
+ $X2=6.29 $Y2=0.665
r493 47 228 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.86 $Y=1.675
+ $X2=5.86 $Y2=1.51
r494 47 49 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.86 $Y=1.675
+ $X2=5.86 $Y2=2.465
r495 43 228 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.86 $Y=1.345
+ $X2=5.86 $Y2=1.51
r496 43 45 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.86 $Y=1.345
+ $X2=5.86 $Y2=0.665
r497 39 227 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.43 $Y=1.675
+ $X2=5.43 $Y2=1.51
r498 39 41 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.43 $Y=1.675
+ $X2=5.43 $Y2=2.465
r499 35 227 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.43 $Y=1.345
+ $X2=5.43 $Y2=1.51
r500 35 37 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.43 $Y=1.345
+ $X2=5.43 $Y2=0.665
r501 31 223 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5 $Y=1.675 $X2=5
+ $Y2=1.51
r502 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5 $Y=1.675 $X2=5
+ $Y2=2.465
r503 27 223 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5 $Y=1.345 $X2=5
+ $Y2=1.51
r504 27 29 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5 $Y=1.345 $X2=5
+ $Y2=0.665
r505 23 221 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.675
+ $X2=4.57 $Y2=1.51
r506 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.57 $Y=1.675
+ $X2=4.57 $Y2=2.465
r507 19 221 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.345
+ $X2=4.57 $Y2=1.51
r508 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.57 $Y=1.345
+ $X2=4.57 $Y2=0.665
r509 6 183 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.835 $X2=3.925 $Y2=2.86
r510 6 181 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.835 $X2=3.925 $Y2=2.095
r511 5 169 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=2.86
r512 5 167 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=2.095
r513 4 155 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.835 $X2=2.205 $Y2=2.86
r514 4 153 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.835 $X2=2.205 $Y2=2.095
r515 3 177 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.785
+ $Y=0.245 $X2=3.925 $Y2=0.48
r516 2 163 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.925
+ $Y=0.245 $X2=3.065 $Y2=0.48
r517 1 149 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.065
+ $Y=0.245 $X2=2.205 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 42 44
+ 48 52 58 64 70 74 78 84 90 96 102 106 110 114 116 120 121 123 124 126 127 128
+ 129 131 132 134 135 136 137 138 144 159 174 180 183 186 189 192 196
r219 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r220 192 193 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r221 189 190 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r222 186 187 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r223 183 184 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r224 180 181 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 178 196 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r226 178 193 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r227 177 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r228 175 192 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.505 $Y=3.33
+ $X2=10.375 $Y2=3.33
r229 175 177 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.505 $Y=3.33
+ $X2=10.8 $Y2=3.33
r230 174 195 4.39729 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=11.105 $Y=3.33
+ $X2=11.312 $Y2=3.33
r231 174 177 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.105 $Y=3.33
+ $X2=10.8 $Y2=3.33
r232 173 193 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r233 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r234 170 173 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r235 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r236 167 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r237 167 190 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r238 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r239 164 189 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.065 $Y=3.33
+ $X2=6.935 $Y2=3.33
r240 164 166 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.065 $Y=3.33
+ $X2=7.44 $Y2=3.33
r241 163 190 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r242 163 187 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r243 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r244 160 186 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.205 $Y=3.33
+ $X2=6.075 $Y2=3.33
r245 160 162 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.205 $Y=3.33
+ $X2=6.48 $Y2=3.33
r246 159 189 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.935 $Y2=3.33
r247 159 162 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.48 $Y2=3.33
r248 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r249 155 158 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r250 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r251 152 155 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r252 152 184 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r253 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r254 149 183 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.635 $Y2=3.33
r255 149 151 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=3.12 $Y2=3.33
r256 148 184 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r257 148 181 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r258 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r259 145 180 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.752 $Y2=3.33
r260 145 147 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r261 144 183 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.635 $Y2=3.33
r262 144 147 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r263 142 181 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r264 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r265 138 187 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r266 138 158 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.04 $Y2=3.33
r267 136 172 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=9.385 $Y=3.33
+ $X2=9.36 $Y2=3.33
r268 136 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.385 $Y=3.33
+ $X2=9.515 $Y2=3.33
r269 134 169 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.525 $Y=3.33
+ $X2=8.4 $Y2=3.33
r270 134 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.525 $Y=3.33
+ $X2=8.655 $Y2=3.33
r271 133 172 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=8.785 $Y=3.33
+ $X2=9.36 $Y2=3.33
r272 133 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.785 $Y=3.33
+ $X2=8.655 $Y2=3.33
r273 131 166 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.44 $Y2=3.33
r274 131 132 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.795 $Y2=3.33
r275 130 169 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=8.4 $Y2=3.33
r276 130 132 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=7.795 $Y2=3.33
r277 128 157 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.085 $Y=3.33
+ $X2=5.04 $Y2=3.33
r278 128 129 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.085 $Y=3.33
+ $X2=5.215 $Y2=3.33
r279 126 154 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.08 $Y2=3.33
r280 126 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.355 $Y2=3.33
r281 125 157 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.485 $Y=3.33
+ $X2=5.04 $Y2=3.33
r282 125 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.485 $Y=3.33
+ $X2=4.355 $Y2=3.33
r283 123 151 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.12 $Y2=3.33
r284 123 124 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.495 $Y2=3.33
r285 122 154 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=4.08 $Y2=3.33
r286 122 124 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=3.495 $Y2=3.33
r287 120 141 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.74 $Y=3.33
+ $X2=0.72 $Y2=3.33
r288 120 121 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.74 $Y=3.33
+ $X2=0.87 $Y2=3.33
r289 116 119 30.862 $w=2.93e-07 $l=7.9e-07 $layer=LI1_cond $X=11.252 $Y=2.12
+ $X2=11.252 $Y2=2.91
r290 114 195 3.08023 $w=2.95e-07 $l=1.11018e-07 $layer=LI1_cond $X=11.252
+ $Y=3.245 $X2=11.312 $Y2=3.33
r291 114 119 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=11.252 $Y=3.245
+ $X2=11.252 $Y2=2.91
r292 110 113 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=10.375 $Y=2.12
+ $X2=10.375 $Y2=2.91
r293 108 192 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.375 $Y=3.245
+ $X2=10.375 $Y2=3.33
r294 108 113 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=10.375 $Y=3.245
+ $X2=10.375 $Y2=2.91
r295 107 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.645 $Y=3.33
+ $X2=9.515 $Y2=3.33
r296 106 192 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.245 $Y=3.33
+ $X2=10.375 $Y2=3.33
r297 106 107 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=10.245 $Y=3.33
+ $X2=9.645 $Y2=3.33
r298 102 105 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=9.515 $Y=2.12
+ $X2=9.515 $Y2=2.91
r299 100 137 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=3.245
+ $X2=9.515 $Y2=3.33
r300 100 105 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=9.515 $Y=3.245
+ $X2=9.515 $Y2=2.91
r301 96 99 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=8.655 $Y=2.12
+ $X2=8.655 $Y2=2.91
r302 94 135 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.655 $Y=3.245
+ $X2=8.655 $Y2=3.33
r303 94 99 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=8.655 $Y=3.245
+ $X2=8.655 $Y2=2.91
r304 90 93 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=7.795 $Y=2.12
+ $X2=7.795 $Y2=2.91
r305 88 132 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.795 $Y=3.245
+ $X2=7.795 $Y2=3.33
r306 88 93 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=7.795 $Y=3.245
+ $X2=7.795 $Y2=2.91
r307 84 87 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=6.935 $Y=2.12
+ $X2=6.935 $Y2=2.91
r308 82 189 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.935 $Y=3.245
+ $X2=6.935 $Y2=3.33
r309 82 87 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=6.935 $Y=3.245
+ $X2=6.935 $Y2=2.91
r310 78 81 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=6.075 $Y=2.12
+ $X2=6.075 $Y2=2.91
r311 76 186 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=3.245
+ $X2=6.075 $Y2=3.33
r312 76 81 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=6.075 $Y=3.245
+ $X2=6.075 $Y2=2.91
r313 75 129 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.345 $Y=3.33
+ $X2=5.215 $Y2=3.33
r314 74 186 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=6.075 $Y2=3.33
r315 74 75 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=5.345 $Y2=3.33
r316 70 73 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=5.215 $Y=2.12
+ $X2=5.215 $Y2=2.91
r317 68 129 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=3.245
+ $X2=5.215 $Y2=3.33
r318 68 73 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=5.215 $Y=3.245
+ $X2=5.215 $Y2=2.91
r319 64 67 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=4.355 $Y=2.27
+ $X2=4.355 $Y2=2.95
r320 62 127 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=3.245
+ $X2=4.355 $Y2=3.33
r321 62 67 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=4.355 $Y=3.245
+ $X2=4.355 $Y2=2.95
r322 58 61 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.495 $Y=2.27
+ $X2=3.495 $Y2=2.95
r323 56 124 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=3.33
r324 56 61 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=2.95
r325 52 55 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=2.635 $Y=2.27
+ $X2=2.635 $Y2=2.95
r326 50 183 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=3.33
r327 50 55 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=2.95
r328 46 180 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.752 $Y=3.245
+ $X2=1.752 $Y2=3.33
r329 46 48 30.6059 $w=3.03e-07 $l=8.1e-07 $layer=LI1_cond $X=1.752 $Y=3.245
+ $X2=1.752 $Y2=2.435
r330 45 121 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=0.87
+ $Y2=3.33
r331 44 180 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=1.6 $Y=3.33
+ $X2=1.752 $Y2=3.33
r332 44 45 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.6 $Y=3.33 $X2=1
+ $Y2=3.33
r333 40 121 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=3.33
r334 40 42 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=2.435
r335 13 119 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.095
+ $Y=1.835 $X2=11.235 $Y2=2.91
r336 13 116 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=11.095
+ $Y=1.835 $X2=11.235 $Y2=2.12
r337 12 113 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.235
+ $Y=1.835 $X2=10.375 $Y2=2.91
r338 12 110 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=10.235
+ $Y=1.835 $X2=10.375 $Y2=2.12
r339 11 105 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.375
+ $Y=1.835 $X2=9.515 $Y2=2.91
r340 11 102 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=9.375
+ $Y=1.835 $X2=9.515 $Y2=2.12
r341 10 99 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.515
+ $Y=1.835 $X2=8.655 $Y2=2.91
r342 10 96 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=8.515
+ $Y=1.835 $X2=8.655 $Y2=2.12
r343 9 93 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.655
+ $Y=1.835 $X2=7.795 $Y2=2.91
r344 9 90 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=7.655
+ $Y=1.835 $X2=7.795 $Y2=2.12
r345 8 87 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.835 $X2=6.935 $Y2=2.91
r346 8 84 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.835 $X2=6.935 $Y2=2.12
r347 7 81 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.935
+ $Y=1.835 $X2=6.075 $Y2=2.91
r348 7 78 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=5.935
+ $Y=1.835 $X2=6.075 $Y2=2.12
r349 6 73 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.075
+ $Y=1.835 $X2=5.215 $Y2=2.91
r350 6 70 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=5.075
+ $Y=1.835 $X2=5.215 $Y2=2.12
r351 5 67 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.215
+ $Y=1.835 $X2=4.355 $Y2=2.95
r352 5 64 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=4.215
+ $Y=1.835 $X2=4.355 $Y2=2.27
r353 4 61 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.355
+ $Y=1.835 $X2=3.495 $Y2=2.95
r354 4 58 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=3.355
+ $Y=1.835 $X2=3.495 $Y2=2.27
r355 3 55 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.835 $X2=2.635 $Y2=2.95
r356 3 52 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.835 $X2=2.635 $Y2=2.27
r357 2 48 300 $w=1.7e-07 $l=6.75278e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.835 $X2=1.75 $Y2=2.435
r358 1 42 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.835 $X2=0.87 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 49 52 62 72 82 92 102 112 122 126
c185 126 0 1.57775e-19 $X=10.805 $Y=2.035
r186 125 129 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=10.805 $Y=2.035
+ $X2=10.805 $Y2=2.86
r187 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.805 $Y=2.035
+ $X2=10.805 $Y2=2.035
r188 122 125 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=10.805 $Y=0.48
+ $X2=10.805 $Y2=2.035
r189 116 126 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.945 $Y=2.035
+ $X2=10.805 $Y2=2.035
r190 115 119 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=9.945 $Y=2.035
+ $X2=9.945 $Y2=2.86
r191 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.945 $Y=2.035
+ $X2=9.945 $Y2=2.035
r192 112 115 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=9.945 $Y=0.48
+ $X2=9.945 $Y2=2.035
r193 106 116 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.085 $Y=2.035
+ $X2=9.945 $Y2=2.035
r194 105 109 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=9.085 $Y=2.035
+ $X2=9.085 $Y2=2.86
r195 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.085 $Y=2.035
+ $X2=9.085 $Y2=2.035
r196 102 105 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=9.085 $Y=0.48
+ $X2=9.085 $Y2=2.035
r197 96 106 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=8.225 $Y=2.035
+ $X2=9.085 $Y2=2.035
r198 95 99 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=8.225 $Y=2.035
+ $X2=8.225 $Y2=2.86
r199 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.225 $Y=2.035
+ $X2=8.225 $Y2=2.035
r200 92 95 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=8.225 $Y=0.48
+ $X2=8.225 $Y2=2.035
r201 85 89 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=7.365 $Y=2.035
+ $X2=7.365 $Y2=2.86
r202 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.365 $Y=2.035
+ $X2=7.365 $Y2=2.035
r203 82 85 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=7.365 $Y=0.48
+ $X2=7.365 $Y2=2.035
r204 76 86 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.505 $Y=2.035
+ $X2=7.365 $Y2=2.035
r205 75 79 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=6.505 $Y=2.035
+ $X2=6.505 $Y2=2.86
r206 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.505 $Y=2.035
+ $X2=6.505 $Y2=2.035
r207 72 75 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=6.505 $Y=0.48
+ $X2=6.505 $Y2=2.035
r208 66 76 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=5.645 $Y=2.035
+ $X2=6.505 $Y2=2.035
r209 65 69 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=5.645 $Y=2.035
+ $X2=5.645 $Y2=2.86
r210 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.645 $Y=2.035
+ $X2=5.645 $Y2=2.035
r211 62 65 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=5.645 $Y=0.48
+ $X2=5.645 $Y2=2.035
r212 56 66 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.785 $Y=2.035
+ $X2=5.645 $Y2=2.035
r213 55 59 42.2562 $w=2.23e-07 $l=8.25e-07 $layer=LI1_cond $X=4.802 $Y=2.035
+ $X2=4.802 $Y2=2.86
r214 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.785 $Y=2.035
+ $X2=4.785 $Y2=2.035
r215 52 55 79.6466 $w=2.23e-07 $l=1.555e-06 $layer=LI1_cond $X=4.802 $Y=0.48
+ $X2=4.802 $Y2=2.035
r216 49 96 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=7.795 $Y=2.035
+ $X2=8.225 $Y2=2.035
r217 49 86 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=7.795 $Y=2.035
+ $X2=7.365 $Y2=2.035
r218 16 129 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=10.665
+ $Y=1.835 $X2=10.805 $Y2=2.86
r219 16 125 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=10.665
+ $Y=1.835 $X2=10.805 $Y2=2.07
r220 15 119 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=9.805
+ $Y=1.835 $X2=9.945 $Y2=2.86
r221 15 115 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=9.805
+ $Y=1.835 $X2=9.945 $Y2=2.07
r222 14 109 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=1.835 $X2=9.085 $Y2=2.86
r223 14 105 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=1.835 $X2=9.085 $Y2=2.07
r224 13 99 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=8.085
+ $Y=1.835 $X2=8.225 $Y2=2.86
r225 13 95 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=8.085
+ $Y=1.835 $X2=8.225 $Y2=2.07
r226 12 89 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=1.835 $X2=7.365 $Y2=2.86
r227 12 85 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=1.835 $X2=7.365 $Y2=2.07
r228 11 79 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=1.835 $X2=6.505 $Y2=2.86
r229 11 75 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=1.835 $X2=6.505 $Y2=2.07
r230 10 69 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.835 $X2=5.645 $Y2=2.86
r231 10 65 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.835 $X2=5.645 $Y2=2.07
r232 9 59 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.835 $X2=4.785 $Y2=2.86
r233 9 55 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.835 $X2=4.785 $Y2=2.07
r234 8 122 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=10.665
+ $Y=0.245 $X2=10.805 $Y2=0.48
r235 7 112 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=9.805
+ $Y=0.245 $X2=9.945 $Y2=0.48
r236 6 102 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=8.945
+ $Y=0.245 $X2=9.085 $Y2=0.48
r237 5 92 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=8.085
+ $Y=0.245 $X2=8.225 $Y2=0.48
r238 4 82 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.225
+ $Y=0.245 $X2=7.365 $Y2=0.48
r239 3 72 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=6.365
+ $Y=0.245 $X2=6.505 $Y2=0.48
r240 2 62 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.505
+ $Y=0.245 $X2=5.645 $Y2=0.48
r241 1 52 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.645
+ $Y=0.245 $X2=4.785 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 42 44
+ 48 52 56 60 64 66 70 74 78 82 86 88 92 94 96 98 99 101 102 104 105 106 107 109
+ 110 112 113 114 115 116 122 137 152 158 161 164 167 170 174
r186 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r187 170 171 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r188 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r189 164 165 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r190 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r191 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r192 156 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r193 156 171 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r194 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r195 153 170 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.505 $Y=0
+ $X2=10.375 $Y2=0
r196 153 155 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.505 $Y=0
+ $X2=10.8 $Y2=0
r197 152 173 4.39729 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=11.105 $Y=0
+ $X2=11.312 $Y2=0
r198 152 155 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.105 $Y=0
+ $X2=10.8 $Y2=0
r199 151 171 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r200 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r201 148 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=9.36 $Y2=0
r202 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r203 145 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.4 $Y2=0
r204 145 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r205 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r206 142 167 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.065 $Y=0
+ $X2=6.935 $Y2=0
r207 142 144 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.065 $Y=0
+ $X2=7.44 $Y2=0
r208 141 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r209 141 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r210 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r211 138 164 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=6.075 $Y2=0
r212 138 140 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=6.48 $Y2=0
r213 137 167 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.805 $Y=0
+ $X2=6.935 $Y2=0
r214 137 140 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=0
+ $X2=6.48 $Y2=0
r215 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r216 133 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r217 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r218 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r219 130 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.64 $Y2=0
r220 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r221 127 161 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.765 $Y=0
+ $X2=2.635 $Y2=0
r222 127 129 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.765 $Y=0
+ $X2=3.12 $Y2=0
r223 126 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r224 126 159 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r225 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r226 123 158 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.87 $Y=0
+ $X2=1.735 $Y2=0
r227 123 125 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.87 $Y=0
+ $X2=2.16 $Y2=0
r228 122 161 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=0
+ $X2=2.635 $Y2=0
r229 122 125 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=0
+ $X2=2.16 $Y2=0
r230 120 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r231 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r232 116 165 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0 $X2=6
+ $Y2=0
r233 116 136 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.04 $Y2=0
r234 114 150 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=9.385 $Y=0
+ $X2=9.36 $Y2=0
r235 114 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.385 $Y=0
+ $X2=9.515 $Y2=0
r236 112 147 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.525 $Y=0
+ $X2=8.4 $Y2=0
r237 112 113 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.525 $Y=0
+ $X2=8.655 $Y2=0
r238 111 150 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=8.785 $Y=0
+ $X2=9.36 $Y2=0
r239 111 113 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.785 $Y=0
+ $X2=8.655 $Y2=0
r240 109 144 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.44 $Y2=0
r241 109 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.795 $Y2=0
r242 108 147 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=7.925 $Y=0
+ $X2=8.4 $Y2=0
r243 108 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.925 $Y=0
+ $X2=7.795 $Y2=0
r244 106 135 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.085 $Y=0
+ $X2=5.04 $Y2=0
r245 106 107 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.085 $Y=0
+ $X2=5.215 $Y2=0
r246 104 132 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.08 $Y2=0
r247 104 105 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.355 $Y2=0
r248 103 135 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.485 $Y=0
+ $X2=5.04 $Y2=0
r249 103 105 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.485 $Y=0
+ $X2=4.355 $Y2=0
r250 101 129 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.365 $Y=0
+ $X2=3.12 $Y2=0
r251 101 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.365 $Y=0
+ $X2=3.495 $Y2=0
r252 100 132 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=0
+ $X2=4.08 $Y2=0
r253 100 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.625 $Y=0
+ $X2=3.495 $Y2=0
r254 98 119 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.72
+ $Y2=0
r255 98 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.87
+ $Y2=0
r256 94 173 3.08023 $w=2.95e-07 $l=1.11018e-07 $layer=LI1_cond $X=11.252
+ $Y=0.085 $X2=11.312 $Y2=0
r257 94 96 15.431 $w=2.93e-07 $l=3.95e-07 $layer=LI1_cond $X=11.252 $Y=0.085
+ $X2=11.252 $Y2=0.48
r258 90 170 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.375 $Y=0.085
+ $X2=10.375 $Y2=0
r259 90 92 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=10.375 $Y=0.085
+ $X2=10.375 $Y2=0.48
r260 89 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.645 $Y=0
+ $X2=9.515 $Y2=0
r261 88 170 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.245 $Y=0
+ $X2=10.375 $Y2=0
r262 88 89 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=10.245 $Y=0 $X2=9.645
+ $Y2=0
r263 84 115 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=0.085
+ $X2=9.515 $Y2=0
r264 84 86 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=9.515 $Y=0.085
+ $X2=9.515 $Y2=0.48
r265 80 113 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.655 $Y=0.085
+ $X2=8.655 $Y2=0
r266 80 82 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=8.655 $Y=0.085
+ $X2=8.655 $Y2=0.48
r267 76 110 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.795 $Y=0.085
+ $X2=7.795 $Y2=0
r268 76 78 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=7.795 $Y=0.085
+ $X2=7.795 $Y2=0.48
r269 72 167 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.935 $Y=0.085
+ $X2=6.935 $Y2=0
r270 72 74 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=6.935 $Y=0.085
+ $X2=6.935 $Y2=0.48
r271 68 164 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=0.085
+ $X2=6.075 $Y2=0
r272 68 70 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=6.075 $Y=0.085
+ $X2=6.075 $Y2=0.48
r273 67 107 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.215 $Y2=0
r274 66 164 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=6.075 $Y2=0
r275 66 67 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.945 $Y=0 $X2=5.345
+ $Y2=0
r276 62 107 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=0.085
+ $X2=5.215 $Y2=0
r277 62 64 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=5.215 $Y=0.085
+ $X2=5.215 $Y2=0.48
r278 58 105 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=0.085
+ $X2=4.355 $Y2=0
r279 58 60 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=4.355 $Y=0.085
+ $X2=4.355 $Y2=0.38
r280 54 102 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=0.085
+ $X2=3.495 $Y2=0
r281 54 56 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.495 $Y=0.085
+ $X2=3.495 $Y2=0.38
r282 50 161 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0
r283 50 52 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0.38
r284 46 158 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r285 46 48 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.4
r286 45 99 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.87
+ $Y2=0
r287 44 158 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=1.735
+ $Y2=0
r288 44 45 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=1 $Y2=0
r289 40 99 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=0.085
+ $X2=0.87 $Y2=0
r290 40 42 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.87 $Y=0.085
+ $X2=0.87 $Y2=0.4
r291 13 96 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=11.095
+ $Y=0.245 $X2=11.235 $Y2=0.48
r292 12 92 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=10.235
+ $Y=0.245 $X2=10.375 $Y2=0.48
r293 11 86 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=9.375
+ $Y=0.245 $X2=9.515 $Y2=0.48
r294 10 82 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=8.515
+ $Y=0.245 $X2=8.655 $Y2=0.48
r295 9 78 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.655
+ $Y=0.245 $X2=7.795 $Y2=0.48
r296 8 74 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=6.795
+ $Y=0.245 $X2=6.935 $Y2=0.48
r297 7 70 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.935
+ $Y=0.245 $X2=6.075 $Y2=0.48
r298 6 64 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.075
+ $Y=0.245 $X2=5.215 $Y2=0.48
r299 5 60 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.215
+ $Y=0.245 $X2=4.355 $Y2=0.38
r300 4 56 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.355
+ $Y=0.245 $X2=3.495 $Y2=0.38
r301 3 52 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.495
+ $Y=0.245 $X2=2.635 $Y2=0.38
r302 2 48 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=1.59
+ $Y=0.245 $X2=1.73 $Y2=0.4
r303 1 42 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.73
+ $Y=0.245 $X2=0.87 $Y2=0.4
.ends

