* File: sky130_fd_sc_lp__xnor2_0.pex.spice
* Created: Fri Aug 28 11:34:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR2_0%A 3 7 10 11 12 13 15 18 23 24 25 27 28 30 33
+ 34 38 42
c84 34 0 1.34543e-19 $X=0.24 $Y=2.035
r85 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.74 $X2=0.385 $Y2=1.74
r86 34 39 5.96849 $w=6.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.4 $Y=2.035
+ $X2=0.4 $Y2=1.74
r87 33 39 1.51741 $w=6.03e-07 $l=7.5e-08 $layer=LI1_cond $X=0.4 $Y=1.665 $X2=0.4
+ $Y2=1.74
r88 31 42 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.175 $Y=0.35
+ $X2=1.325 $Y2=0.35
r89 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=0.35 $X2=1.175 $Y2=0.35
r90 28 30 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=0.715 $Y=0.385
+ $X2=1.175 $Y2=0.385
r91 27 33 11.7954 $w=6.03e-07 $l=3.30568e-07 $layer=LI1_cond $X=0.63 $Y=1.43
+ $X2=0.4 $Y2=1.665
r92 26 28 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.63 $Y=0.515
+ $X2=0.715 $Y2=0.385
r93 26 27 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=0.63 $Y=0.515
+ $X2=0.63 $Y2=1.43
r94 23 38 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.385 $Y=2.095
+ $X2=0.385 $Y2=1.74
r95 23 24 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.467 $Y=2.095
+ $X2=0.467 $Y2=2.245
r96 21 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.575
+ $X2=0.385 $Y2=1.74
r97 16 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=0.98
+ $X2=1.84 $Y2=0.905
r98 16 18 910.16 $w=1.5e-07 $l=1.775e-06 $layer=POLY_cond $X=1.84 $Y=0.98
+ $X2=1.84 $Y2=2.755
r99 13 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=0.83
+ $X2=1.84 $Y2=0.905
r100 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.84 $Y=0.83
+ $X2=1.84 $Y2=0.51
r101 11 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=0.905
+ $X2=1.84 $Y2=0.905
r102 11 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.765 $Y=0.905
+ $X2=1.4 $Y2=0.905
r103 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.325 $Y=0.83
+ $X2=1.4 $Y2=0.905
r104 9 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=0.515
+ $X2=1.325 $Y2=0.35
r105 9 10 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.325 $Y=0.515
+ $X2=1.325 $Y2=0.83
r106 7 24 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.64 $Y=2.755
+ $X2=0.64 $Y2=2.245
r107 3 21 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.475 $Y=1.095
+ $X2=0.475 $Y2=1.575
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_0%B 1 3 6 10 14 18 19 20 21 25 28
c75 25 0 1.78581e-19 $X=2.29 $Y=1.385
c76 14 0 4.16037e-20 $X=2.27 $Y=0.51
c77 6 0 1.34543e-19 $X=1.07 $Y=2.755
c78 1 0 5.50351e-20 $X=0.835 $Y=1.425
r79 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.39
+ $Y=1.59 $X2=1.39 $Y2=1.59
r80 28 30 29.8915 $w=5.16e-07 $l=3.2e-07 $layer=POLY_cond $X=1.07 $Y=1.76
+ $X2=1.39 $Y2=1.76
r81 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.385 $X2=2.29 $Y2=1.385
r82 21 26 2.3707 $w=6.69e-07 $l=1.3e-07 $layer=LI1_cond $X=2.16 $Y=1.657
+ $X2=2.29 $Y2=1.657
r83 20 21 8.75336 $w=6.69e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.657
+ $X2=2.16 $Y2=1.657
r84 20 31 5.28849 $w=6.69e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.657
+ $X2=1.39 $Y2=1.657
r85 18 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.29 $Y=1.725
+ $X2=2.29 $Y2=1.385
r86 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.725
+ $X2=2.29 $Y2=1.89
r87 17 25 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.22
+ $X2=2.29 $Y2=1.385
r88 14 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.27 $Y=0.51
+ $X2=2.27 $Y2=1.22
r89 10 19 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=2.2 $Y=2.755
+ $X2=2.2 $Y2=1.89
r90 4 28 32.2057 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.07 $Y=2.095
+ $X2=1.07 $Y2=1.76
r91 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.07 $Y=2.095 $X2=1.07
+ $Y2=2.755
r92 1 28 21.9515 $w=5.16e-07 $l=4.36978e-07 $layer=POLY_cond $X=0.835 $Y=1.425
+ $X2=1.07 $Y2=1.76
r93 1 3 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.835 $Y=1.425
+ $X2=0.835 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_0%A_143_487# 1 2 9 13 16 18 19 22 25 26 28 32
+ 33 35 37 40
r82 40 42 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.015 $Y=2.15
+ $X2=2.015 $Y2=2.35
r83 37 39 6.63994 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.05 $Y=1.095
+ $X2=1.05 $Y2=1.26
r84 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.835
+ $Y=1.73 $X2=2.835 $Y2=1.73
r85 30 32 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.8 $Y=2.065
+ $X2=2.8 $Y2=1.73
r86 29 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=2.15
+ $X2=2.015 $Y2=2.15
r87 28 30 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.67 $Y=2.15
+ $X2=2.8 $Y2=2.065
r88 28 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.67 $Y=2.15 $X2=2.1
+ $Y2=2.15
r89 27 35 2.68609 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.125 $Y=2.35
+ $X2=0.932 $Y2=2.35
r90 26 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=2.35
+ $X2=2.015 $Y2=2.35
r91 26 27 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.93 $Y=2.35
+ $X2=1.125 $Y2=2.35
r92 25 35 3.77418 $w=2.45e-07 $l=1.15888e-07 $layer=LI1_cond $X=1.005 $Y=2.265
+ $X2=0.932 $Y2=2.35
r93 25 39 48.2585 $w=2.38e-07 $l=1.005e-06 $layer=LI1_cond $X=1.005 $Y=2.265
+ $X2=1.005 $Y2=1.26
r94 20 35 3.77418 $w=2.45e-07 $l=1.13666e-07 $layer=LI1_cond $X=0.865 $Y=2.435
+ $X2=0.932 $Y2=2.35
r95 20 22 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.865 $Y=2.435
+ $X2=0.865 $Y2=2.56
r96 19 33 131.146 $w=3.3e-07 $l=7.5e-07 $layer=POLY_cond $X=2.835 $Y=0.98
+ $X2=2.835 $Y2=1.73
r97 18 19 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.812 $Y=0.83
+ $X2=2.812 $Y2=0.98
r98 15 33 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=2.835 $Y=2.13
+ $X2=2.835 $Y2=1.73
r99 15 16 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.787 $Y=2.13
+ $X2=2.787 $Y2=2.28
r100 13 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.7 $Y=0.51 $X2=2.7
+ $Y2=0.83
r101 9 16 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=2.65 $Y=2.755
+ $X2=2.65 $Y2=2.28
r102 2 22 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.715
+ $Y=2.435 $X2=0.855 $Y2=2.56
r103 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.885 $X2=1.05 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_0%VPWR 1 2 3 10 12 14 18 22 24 25 26 27 35 40
r41 40 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 38 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 29 40 12.9051 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=1.79 $Y=3.33
+ $X2=1.475 $Y2=3.33
r48 29 31 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.79 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 27 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 27 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 27 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 25 31 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 25 26 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.915 $Y2=3.33
r54 24 34 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=3.06 $Y=3.33 $X2=3.12
+ $Y2=3.33
r55 24 26 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.06 $Y=3.33
+ $X2=2.915 $Y2=3.33
r56 20 26 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=3.33
r57 20 22 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=2.91
r58 16 40 2.6323 $w=6.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=3.33
r59 16 18 9.01805 $w=6.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=2.77
r60 15 37 4.33154 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.285 $Y2=3.33
r61 14 40 12.9051 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=1.475 $Y2=3.33
r62 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.16 $Y=3.33 $X2=0.57
+ $Y2=3.33
r63 10 37 3.26765 $w=3.1e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.285 $Y2=3.33
r64 10 12 24.7218 $w=3.08e-07 $l=6.65e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.415 $Y2=2.58
r65 3 22 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=2.725
+ $Y=2.435 $X2=2.865 $Y2=2.91
r66 2 18 300 $w=1.7e-07 $l=6.2546e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.435 $X2=1.625 $Y2=2.77
r67 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=2.435 $X2=0.425 $Y2=2.58
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_0%Y 1 2 9 11 12 13 14 15 16 23
c41 16 0 1.78581e-19 $X=3.12 $Y=1.295
r42 16 21 4.02526 $w=5.18e-07 $l=1.75e-07 $layer=LI1_cond $X=3.01 $Y=1.295
+ $X2=3.01 $Y2=1.12
r43 15 21 4.48529 $w=5.18e-07 $l=1.95e-07 $layer=LI1_cond $X=3.01 $Y=0.925
+ $X2=3.01 $Y2=1.12
r44 14 15 8.51056 $w=5.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.01 $Y=0.555
+ $X2=3.01 $Y2=0.925
r45 14 23 1.03507 $w=5.18e-07 $l=4.5e-08 $layer=LI1_cond $X=3.01 $Y=0.555
+ $X2=3.01 $Y2=0.51
r46 13 16 44.1806 $w=2.73e-07 $l=1.025e-06 $layer=LI1_cond $X=3.185 $Y=2.405
+ $X2=3.185 $Y2=1.38
r47 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.49
+ $X2=3.185 $Y2=2.405
r48 11 12 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.1 $Y=2.49 $X2=2.6
+ $Y2=2.49
r49 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.435 $Y=2.575
+ $X2=2.6 $Y2=2.49
r50 7 9 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.435 $Y=2.575
+ $X2=2.435 $Y2=2.58
r51 2 9 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=2.435 $X2=2.435 $Y2=2.58
r52 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.3 $X2=2.915 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_0%VGND 1 2 7 9 13 15 17 27 28 34
r39 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 28 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r42 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 25 34 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.052
+ $Y2=0
r44 25 27 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=3.12
+ $Y2=0
r45 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r46 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r47 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 18 31 4.31056 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=0.187
+ $Y2=0
r49 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=0.72
+ $Y2=0
r50 17 34 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=2.052
+ $Y2=0
r51 17 23 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=1.68
+ $Y2=0
r52 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r53 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r54 15 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 11 34 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.052 $Y=0.085
+ $X2=2.052 $Y2=0
r56 11 13 19.2074 $w=2.53e-07 $l=4.25e-07 $layer=LI1_cond $X=2.052 $Y=0.085
+ $X2=2.052 $Y2=0.51
r57 7 31 3.04949 $w=2.8e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.187 $Y2=0
r58 7 9 41.5703 $w=2.78e-07 $l=1.01e-06 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.235 $Y2=1.095
r59 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.3 $X2=2.055 $Y2=0.51
r60 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.885 $X2=0.26 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_0%A_300_60# 1 2 9 11 12 15
c31 9 0 9.66388e-20 $X=1.625 $Y=0.51
r32 13 15 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.465 $Y=0.845
+ $X2=2.465 $Y2=0.51
r33 11 13 6.89722 $w=1.9e-07 $l=1.55403e-07 $layer=LI1_cond $X=2.35 $Y=0.94
+ $X2=2.465 $Y2=0.845
r34 11 12 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=2.35 $Y=0.94
+ $X2=1.755 $Y2=0.94
r35 7 12 6.95919 $w=1.9e-07 $l=1.6375e-07 $layer=LI1_cond $X=1.632 $Y=0.845
+ $X2=1.755 $Y2=0.94
r36 7 9 15.7579 $w=2.43e-07 $l=3.35e-07 $layer=LI1_cond $X=1.632 $Y=0.845
+ $X2=1.632 $Y2=0.51
r37 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.3 $X2=2.485 $Y2=0.51
r38 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.5 $Y=0.3
+ $X2=1.625 $Y2=0.51
.ends

