* File: sky130_fd_sc_lp__dfstp_4.pxi.spice
* Created: Fri Aug 28 10:23:26 2020
* 
x_PM_SKY130_FD_SC_LP__DFSTP_4%CLK N_CLK_M1013_g N_CLK_c_249_n N_CLK_M1005_g
+ N_CLK_c_250_n CLK CLK CLK CLK CLK N_CLK_c_252_n N_CLK_c_253_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%CLK
x_PM_SKY130_FD_SC_LP__DFSTP_4%D N_D_c_288_n N_D_c_289_n N_D_c_292_n N_D_c_290_n
+ N_D_M1037_g N_D_c_293_n N_D_M1031_g D N_D_c_295_n N_D_c_291_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%D
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_230_465# N_A_230_465#_M1001_d
+ N_A_230_465#_M1025_d N_A_230_465#_c_340_n N_A_230_465#_M1019_g
+ N_A_230_465#_M1027_g N_A_230_465#_M1018_g N_A_230_465#_M1036_g
+ N_A_230_465#_c_345_n N_A_230_465#_c_357_n N_A_230_465#_c_346_n
+ N_A_230_465#_c_359_n N_A_230_465#_c_347_n N_A_230_465#_c_348_n
+ N_A_230_465#_c_349_n N_A_230_465#_c_350_n N_A_230_465#_c_351_n
+ N_A_230_465#_c_399_p N_A_230_465#_c_352_n N_A_230_465#_c_353_n
+ N_A_230_465#_c_354_n PM_SKY130_FD_SC_LP__DFSTP_4%A_230_465#
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_690_93# N_A_690_93#_M1007_s N_A_690_93#_M1016_d
+ N_A_690_93#_c_513_n N_A_690_93#_M1035_g N_A_690_93#_M1006_g
+ N_A_690_93#_c_520_n N_A_690_93#_c_521_n N_A_690_93#_c_514_n
+ N_A_690_93#_c_515_n N_A_690_93#_c_516_n N_A_690_93#_c_532_p
+ N_A_690_93#_c_522_n N_A_690_93#_c_517_n N_A_690_93#_c_518_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%A_690_93#
x_PM_SKY130_FD_SC_LP__DFSTP_4%SET_B N_SET_B_M1003_g N_SET_B_M1009_g
+ N_SET_B_c_597_n N_SET_B_M1034_g N_SET_B_c_598_n N_SET_B_c_599_n
+ N_SET_B_c_600_n N_SET_B_M1032_g N_SET_B_c_601_n N_SET_B_c_602_n
+ N_SET_B_c_610_n N_SET_B_c_611_n N_SET_B_c_612_n N_SET_B_c_603_n SET_B SET_B
+ SET_B SET_B SET_B N_SET_B_c_605_n PM_SKY130_FD_SC_LP__DFSTP_4%SET_B
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_562_119# N_A_562_119#_M1002_d
+ N_A_562_119#_M1019_d N_A_562_119#_M1016_g N_A_562_119#_M1007_g
+ N_A_562_119#_c_715_n N_A_562_119#_c_716_n N_A_562_119#_M1020_g
+ N_A_562_119#_c_718_n N_A_562_119#_c_719_n N_A_562_119#_c_720_n
+ N_A_562_119#_M1015_g N_A_562_119#_c_721_n N_A_562_119#_c_722_n
+ N_A_562_119#_c_723_n N_A_562_119#_c_724_n N_A_562_119#_c_730_n
+ N_A_562_119#_c_731_n N_A_562_119#_c_732_n N_A_562_119#_c_725_n
+ N_A_562_119#_c_726_n PM_SKY130_FD_SC_LP__DFSTP_4%A_562_119#
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_30_99# N_A_30_99#_M1013_s N_A_30_99#_M1005_s
+ N_A_30_99#_c_857_n N_A_30_99#_M1025_g N_A_30_99#_c_859_n N_A_30_99#_c_860_n
+ N_A_30_99#_M1001_g N_A_30_99#_c_850_n N_A_30_99#_c_851_n N_A_30_99#_M1002_g
+ N_A_30_99#_M1000_g N_A_30_99#_c_862_n N_A_30_99#_M1021_g N_A_30_99#_M1026_g
+ N_A_30_99#_c_865_n N_A_30_99#_c_866_n N_A_30_99#_c_867_n N_A_30_99#_c_854_n
+ N_A_30_99#_c_869_n N_A_30_99#_c_870_n N_A_30_99#_c_855_n N_A_30_99#_c_856_n
+ N_A_30_99#_c_873_n PM_SKY130_FD_SC_LP__DFSTP_4%A_30_99#
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_1398_65# N_A_1398_65#_M1028_d
+ N_A_1398_65#_M1024_d N_A_1398_65#_M1008_g N_A_1398_65#_c_988_n
+ N_A_1398_65#_c_989_n N_A_1398_65#_c_990_n N_A_1398_65#_c_996_n
+ N_A_1398_65#_c_997_n N_A_1398_65#_M1014_g N_A_1398_65#_c_999_n
+ N_A_1398_65#_c_1000_n N_A_1398_65#_c_991_n N_A_1398_65#_c_992_n
+ N_A_1398_65#_c_993_n N_A_1398_65#_c_994_n N_A_1398_65#_c_1002_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%A_1398_65#
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_1247_47# N_A_1247_47#_M1018_d
+ N_A_1247_47#_M1036_d N_A_1247_47#_M1032_d N_A_1247_47#_c_1079_n
+ N_A_1247_47#_M1028_g N_A_1247_47#_c_1080_n N_A_1247_47#_c_1081_n
+ N_A_1247_47#_c_1082_n N_A_1247_47#_c_1095_n N_A_1247_47#_M1024_g
+ N_A_1247_47#_c_1083_n N_A_1247_47#_M1012_g N_A_1247_47#_M1011_g
+ N_A_1247_47#_c_1086_n N_A_1247_47#_c_1087_n N_A_1247_47#_c_1088_n
+ N_A_1247_47#_c_1089_n N_A_1247_47#_c_1099_n N_A_1247_47#_c_1100_n
+ N_A_1247_47#_c_1090_n N_A_1247_47#_c_1091_n N_A_1247_47#_c_1147_n
+ N_A_1247_47#_c_1092_n N_A_1247_47#_c_1102_n N_A_1247_47#_c_1103_n
+ N_A_1247_47#_c_1093_n N_A_1247_47#_c_1094_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%A_1247_47#
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_1989_49# N_A_1989_49#_M1012_s
+ N_A_1989_49#_M1011_s N_A_1989_49#_M1010_g N_A_1989_49#_M1004_g
+ N_A_1989_49#_M1023_g N_A_1989_49#_M1017_g N_A_1989_49#_M1029_g
+ N_A_1989_49#_M1022_g N_A_1989_49#_M1030_g N_A_1989_49#_M1033_g
+ N_A_1989_49#_c_1204_n N_A_1989_49#_c_1205_n N_A_1989_49#_c_1206_n
+ N_A_1989_49#_c_1207_n N_A_1989_49#_c_1208_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%A_1989_49#
x_PM_SKY130_FD_SC_LP__DFSTP_4%VPWR N_VPWR_M1005_d N_VPWR_M1031_s N_VPWR_M1006_d
+ N_VPWR_M1003_d N_VPWR_M1014_d N_VPWR_M1024_s N_VPWR_M1011_d N_VPWR_M1017_s
+ N_VPWR_M1033_s N_VPWR_c_1296_n N_VPWR_c_1297_n N_VPWR_c_1298_n N_VPWR_c_1299_n
+ N_VPWR_c_1300_n N_VPWR_c_1301_n N_VPWR_c_1302_n N_VPWR_c_1303_n
+ N_VPWR_c_1304_n N_VPWR_c_1305_n N_VPWR_c_1306_n N_VPWR_c_1307_n
+ N_VPWR_c_1308_n N_VPWR_c_1309_n N_VPWR_c_1310_n N_VPWR_c_1311_n
+ N_VPWR_c_1312_n VPWR N_VPWR_c_1313_n N_VPWR_c_1314_n N_VPWR_c_1315_n
+ N_VPWR_c_1316_n N_VPWR_c_1317_n N_VPWR_c_1318_n N_VPWR_c_1319_n
+ N_VPWR_c_1320_n N_VPWR_c_1321_n N_VPWR_c_1295_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%VPWR
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_476_119# N_A_476_119#_M1037_d
+ N_A_476_119#_M1031_d N_A_476_119#_c_1458_n N_A_476_119#_c_1461_n
+ N_A_476_119#_c_1459_n N_A_476_119#_c_1460_n N_A_476_119#_c_1463_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%A_476_119#
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_1094_379# N_A_1094_379#_M1020_d
+ N_A_1094_379#_M1026_d N_A_1094_379#_c_1506_n N_A_1094_379#_c_1507_n
+ N_A_1094_379#_c_1508_n PM_SKY130_FD_SC_LP__DFSTP_4%A_1094_379#
x_PM_SKY130_FD_SC_LP__DFSTP_4%A_1201_407# N_A_1201_407#_M1036_s
+ N_A_1201_407#_M1014_s N_A_1201_407#_c_1533_n N_A_1201_407#_c_1534_n
+ N_A_1201_407#_c_1535_n N_A_1201_407#_c_1536_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%A_1201_407#
x_PM_SKY130_FD_SC_LP__DFSTP_4%Q N_Q_M1010_s N_Q_M1029_s N_Q_M1004_d N_Q_M1022_d
+ N_Q_c_1616_p N_Q_c_1601_n N_Q_c_1562_n N_Q_c_1563_n N_Q_c_1568_n N_Q_c_1569_n
+ N_Q_c_1617_p N_Q_c_1606_n N_Q_c_1564_n N_Q_c_1570_n N_Q_c_1565_n N_Q_c_1571_n
+ Q N_Q_c_1566_n Q PM_SKY130_FD_SC_LP__DFSTP_4%Q
x_PM_SKY130_FD_SC_LP__DFSTP_4%VGND N_VGND_M1013_d N_VGND_M1037_s N_VGND_M1035_d
+ N_VGND_M1009_d N_VGND_M1034_d N_VGND_M1012_d N_VGND_M1023_d N_VGND_M1030_d
+ N_VGND_c_1622_n N_VGND_c_1623_n N_VGND_c_1624_n N_VGND_c_1625_n
+ N_VGND_c_1626_n N_VGND_c_1627_n N_VGND_c_1628_n N_VGND_c_1629_n
+ N_VGND_c_1630_n N_VGND_c_1631_n N_VGND_c_1632_n N_VGND_c_1633_n
+ N_VGND_c_1634_n VGND N_VGND_c_1635_n N_VGND_c_1636_n N_VGND_c_1637_n
+ N_VGND_c_1638_n N_VGND_c_1639_n N_VGND_c_1640_n N_VGND_c_1641_n
+ N_VGND_c_1642_n N_VGND_c_1643_n N_VGND_c_1644_n N_VGND_c_1645_n
+ PM_SKY130_FD_SC_LP__DFSTP_4%VGND
cc_1 VNB N_CLK_c_249_n 0.0238051f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.508
cc_2 VNB N_CLK_c_250_n 0.0107798f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.695
cc_3 VNB CLK 0.0107565f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_4 VNB N_CLK_c_252_n 0.0216237f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.19
cc_5 VNB N_CLK_c_253_n 0.0220103f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.025
cc_6 VNB N_D_c_288_n 0.023366f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.705
cc_7 VNB N_D_c_289_n 0.0131447f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.212
cc_8 VNB N_D_c_290_n 0.0165279f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.645
cc_9 VNB N_D_c_291_n 0.0221554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_230_465#_c_340_n 0.0178293f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.645
cc_11 VNB N_A_230_465#_M1019_g 0.00108725f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_12 VNB N_A_230_465#_M1027_g 0.035274f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_13 VNB N_A_230_465#_M1018_g 0.0398602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_230_465#_M1036_g 0.00497212f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.19
cc_15 VNB N_A_230_465#_c_345_n 0.0224342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_230_465#_c_346_n 0.00229714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_230_465#_c_347_n 0.0093691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_230_465#_c_348_n 0.00268581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_230_465#_c_349_n 0.0331545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_230_465#_c_350_n 0.00167695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_230_465#_c_351_n 0.0179553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_230_465#_c_352_n 0.0156662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_230_465#_c_353_n 0.0129604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_230_465#_c_354_n 0.0472022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_690_93#_c_513_n 0.0189474f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.645
cc_26 VNB N_A_690_93#_c_514_n 0.0132074f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.19
cc_27 VNB N_A_690_93#_c_515_n 0.00926378f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.555
cc_28 VNB N_A_690_93#_c_516_n 2.63896e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_690_93#_c_517_n 0.035552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_690_93#_c_518_n 0.0111411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_SET_B_c_597_n 0.0175787f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.645
cc_32 VNB N_SET_B_c_598_n 0.0158366f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_33 VNB N_SET_B_c_599_n 0.00677902f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_34 VNB N_SET_B_c_600_n 0.0831283f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_35 VNB N_SET_B_c_601_n 0.010839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_SET_B_c_602_n 0.0325651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_SET_B_c_603_n 0.00225764f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.19
cc_38 VNB SET_B 0.012893f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=2.035
cc_39 VNB N_SET_B_c_605_n 0.0193038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_562_119#_M1016_g 0.00427787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_562_119#_M1007_g 0.0501049f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_42 VNB N_A_562_119#_c_715_n 0.0374332f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_43 VNB N_A_562_119#_c_716_n 0.0188014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_562_119#_M1020_g 0.00375483f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.19
cc_45 VNB N_A_562_119#_c_718_n 0.0220705f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.19
cc_46 VNB N_A_562_119#_c_719_n 0.00947912f $X=-0.19 $Y=-0.245 $X2=0.602
+ $Y2=1.025
cc_47 VNB N_A_562_119#_c_720_n 0.0187524f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.555
cc_48 VNB N_A_562_119#_c_721_n 0.00391059f $X=-0.19 $Y=-0.245 $X2=0.672
+ $Y2=0.925
cc_49 VNB N_A_562_119#_c_722_n 0.00367596f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.19
cc_50 VNB N_A_562_119#_c_723_n 0.00625022f $X=-0.19 $Y=-0.245 $X2=0.672
+ $Y2=1.665
cc_51 VNB N_A_562_119#_c_724_n 0.00419806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_562_119#_c_725_n 8.09904e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_562_119#_c_726_n 0.0445073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_30_99#_M1001_g 0.0547976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_30_99#_c_850_n 0.10775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_30_99#_c_851_n 0.0125015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_30_99#_M1002_g 0.0344914f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.19
cc_58 VNB N_A_30_99#_M1021_g 0.0468852f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.665
cc_59 VNB N_A_30_99#_c_854_n 0.0349844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_30_99#_c_855_n 0.00363788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_30_99#_c_856_n 0.0189896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1398_65#_M1008_g 0.0355071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1398_65#_c_988_n 0.022656f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_64 VNB N_A_1398_65#_c_989_n 0.00819273f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_65 VNB N_A_1398_65#_c_990_n 0.00575531f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_66 VNB N_A_1398_65#_c_991_n 0.00442222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1398_65#_c_992_n 0.0178933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1398_65#_c_993_n 5.317e-19 $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.19
cc_69 VNB N_A_1398_65#_c_994_n 0.0239186f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.665
cc_70 VNB N_A_1247_47#_c_1079_n 0.0178311f $X=-0.19 $Y=-0.245 $X2=0.602
+ $Y2=1.695
cc_71 VNB N_A_1247_47#_c_1080_n 0.059437f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_72 VNB N_A_1247_47#_c_1081_n 0.0114857f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_73 VNB N_A_1247_47#_c_1082_n 0.0132775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1247_47#_c_1083_n 0.0395841f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.19
cc_75 VNB N_A_1247_47#_M1012_g 0.0318087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1247_47#_M1011_g 0.00497788f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.19
cc_77 VNB N_A_1247_47#_c_1086_n 0.00378487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1247_47#_c_1087_n 0.00436351f $X=-0.19 $Y=-0.245 $X2=0.672
+ $Y2=1.665
cc_79 VNB N_A_1247_47#_c_1088_n 0.0043288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1247_47#_c_1089_n 0.003552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1247_47#_c_1090_n 0.0102409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1247_47#_c_1091_n 0.0117868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1247_47#_c_1092_n 0.0895241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1247_47#_c_1093_n 0.038651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1247_47#_c_1094_n 0.0129439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1989_49#_M1010_g 0.0242526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1989_49#_M1023_g 0.0222627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1989_49#_M1029_g 0.0222413f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.555
cc_89 VNB N_A_1989_49#_M1030_g 0.027033f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.665
cc_90 VNB N_A_1989_49#_c_1204_n 0.00682622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1989_49#_c_1205_n 9.93652e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1989_49#_c_1206_n 0.00632282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1989_49#_c_1207_n 2.23393e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1989_49#_c_1208_n 0.0682463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VPWR_c_1295_n 0.521925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_476_119#_c_1458_n 0.00187788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_476_119#_c_1459_n 0.00831614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_476_119#_c_1460_n 0.00677324f $X=-0.19 $Y=-0.245 $X2=0.602
+ $Y2=1.19
cc_99 VNB N_Q_c_1562_n 0.00310505f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.19
cc_100 VNB N_Q_c_1563_n 0.00375808f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.025
cc_101 VNB N_Q_c_1564_n 0.0012391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_Q_c_1565_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_Q_c_1566_n 0.0083195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB Q 0.0205513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1622_n 0.0149278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1623_n 0.0104221f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.295
cc_107 VNB N_VGND_c_1624_n 0.0383277f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.665
cc_108 VNB N_VGND_c_1625_n 0.0211512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1626_n 0.0107141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1627_n 0.00839581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1628_n 4.81113e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1629_n 0.0104415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1630_n 0.0289266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1631_n 0.0303931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1632_n 0.00423165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1633_n 0.0544519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1634_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1635_n 0.0213055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1636_n 0.0277957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1637_n 0.0490112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1638_n 0.0148369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1639_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1640_n 0.00319606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1641_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1642_n 0.0215379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1643_n 0.0123565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1644_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1645_n 0.647038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VPB N_CLK_M1005_g 0.0507229f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.645
cc_130 VPB N_CLK_c_250_n 0.0101651f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.695
cc_131 VPB CLK 0.00825547f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_132 VPB N_D_c_292_n 0.0350806f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.508
cc_133 VPB N_D_c_293_n 0.0185375f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.695
cc_134 VPB D 0.00950335f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_135 VPB N_D_c_295_n 0.0428749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_D_c_291_n 0.0173662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_230_465#_M1019_g 0.0512347f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_138 VPB N_A_230_465#_M1036_g 0.0355337f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.19
cc_139 VPB N_A_230_465#_c_357_n 0.0248042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_230_465#_c_346_n 0.00253593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_230_465#_c_359_n 0.0106447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_230_465#_c_348_n 0.00651127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_230_465#_c_352_n 0.0164856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_230_465#_c_354_n 0.00904803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_690_93#_M1006_g 0.0181012f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_146 VPB N_A_690_93#_c_520_n 0.0107669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_690_93#_c_521_n 0.0321364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_690_93#_c_522_n 0.0014421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_690_93#_c_518_n 0.0107065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_SET_B_M1003_g 0.0203374f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.705
cc_151 VPB N_SET_B_c_600_n 0.043107f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_152 VPB N_SET_B_M1032_g 0.0362486f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_153 VPB N_SET_B_c_601_n 0.00214154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_SET_B_c_610_n 0.00865654f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.19
cc_155 VPB N_SET_B_c_611_n 0.0347557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_SET_B_c_612_n 0.0183394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_SET_B_c_603_n 0.00473642f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=1.19
cc_158 VPB SET_B 0.0135107f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=2.035
cc_159 VPB N_A_562_119#_M1016_g 0.0419977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_562_119#_M1020_g 0.0290611f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.19
cc_161 VPB N_A_562_119#_c_723_n 0.0117158f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=1.665
cc_162 VPB N_A_562_119#_c_730_n 0.00201425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_562_119#_c_731_n 0.0120155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_562_119#_c_732_n 4.27224e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_562_119#_c_725_n 0.00246222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_30_99#_c_857_n 0.0254972f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.645
cc_167 VPB N_A_30_99#_M1025_g 0.011352f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_168 VPB N_A_30_99#_c_859_n 0.165146f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_169 VPB N_A_30_99#_c_860_n 0.0113013f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_170 VPB N_A_30_99#_M1000_g 0.0366071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_30_99#_c_862_n 0.255799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_30_99#_M1021_g 0.00575531f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=1.665
cc_173 VPB N_A_30_99#_M1026_g 0.0193446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_30_99#_c_865_n 0.0206327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_30_99#_c_866_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_30_99#_c_867_n 0.0192814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_30_99#_c_854_n 0.0312541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_30_99#_c_869_n 0.0242427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_30_99#_c_870_n 0.00769821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_30_99#_c_855_n 0.00105281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_30_99#_c_856_n 0.00162808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_30_99#_c_873_n 0.011795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1398_65#_c_990_n 0.0837868f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_184 VPB N_A_1398_65#_c_996_n 0.020976f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_185 VPB N_A_1398_65#_c_997_n 0.0104278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1398_65#_M1014_g 0.0303173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1398_65#_c_999_n 0.125784f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.19
cc_188 VPB N_A_1398_65#_c_1000_n 0.00732516f $X=-0.19 $Y=1.655 $X2=0.625
+ $Y2=1.19
cc_189 VPB N_A_1398_65#_c_994_n 0.0189899f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=1.665
cc_190 VPB N_A_1398_65#_c_1002_n 0.0656568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1247_47#_c_1095_n 0.0235434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_1247_47#_c_1083_n 0.0149597f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.19
cc_193 VPB N_A_1247_47#_M1011_g 0.0215564f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=1.19
cc_194 VPB N_A_1247_47#_c_1086_n 0.00331176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1247_47#_c_1099_n 0.0186175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1247_47#_c_1100_n 0.00844457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_1247_47#_c_1090_n 0.00987268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1247_47#_c_1102_n 0.00230666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_1247_47#_c_1103_n 0.00892077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1989_49#_M1004_g 0.0190266f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_201 VPB N_A_1989_49#_M1017_g 0.0179297f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.19
cc_202 VPB N_A_1989_49#_M1022_g 0.0179086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1989_49#_M1033_g 0.0212797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1989_49#_c_1205_n 0.00353669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1989_49#_c_1208_n 0.0117266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1296_n 0.00216255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1297_n 0.0220996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1298_n 0.0129695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1299_n 0.0242902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1300_n 0.0162292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1301_n 0.00943361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1302_n 0.0271946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1303_n 0.00788231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1304_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1305_n 0.0102373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1306_n 0.0412014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1307_n 0.0647557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1308_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1309_n 0.0180783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1310_n 0.0034365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1311_n 0.0284413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1312_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1313_n 0.0300585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1314_n 0.03832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1315_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1316_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1317_n 0.0263077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1318_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1319_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1320_n 0.0034365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1321_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1295_n 0.0599778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_476_119#_c_1461_n 0.00402093f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.21
cc_234 VPB N_A_476_119#_c_1460_n 0.00463266f $X=-0.19 $Y=1.655 $X2=0.602
+ $Y2=1.19
cc_235 VPB N_A_476_119#_c_1463_n 0.00343104f $X=-0.19 $Y=1.655 $X2=0.625
+ $Y2=1.19
cc_236 VPB N_A_1094_379#_c_1506_n 0.0127277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_1094_379#_c_1507_n 0.00448509f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=0.47
cc_238 VPB N_A_1094_379#_c_1508_n 0.0260455f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.21
cc_239 VPB N_A_1201_407#_c_1533_n 0.00423352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1201_407#_c_1534_n 0.00786899f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=0.47
cc_241 VPB N_A_1201_407#_c_1535_n 0.00408906f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=0.84
cc_242 VPB N_A_1201_407#_c_1536_n 0.00281309f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.58
cc_243 VPB N_Q_c_1568_n 0.00304538f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=0.555
cc_244 VPB N_Q_c_1569_n 0.00248092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_Q_c_1570_n 0.00922706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_Q_c_1571_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB Q 0.00547496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 CLK N_A_230_465#_c_347_n 0.00143727f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_249 CLK N_A_230_465#_c_348_n 3.52783e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_250 CLK N_A_230_465#_c_351_n 0.0184962f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_251 N_CLK_M1005_g N_A_30_99#_c_857_n 0.0447826f $X=0.645 $Y=2.645 $X2=0 $Y2=0
cc_252 N_CLK_c_250_n N_A_30_99#_c_857_n 0.00627853f $X=0.602 $Y=1.695 $X2=0
+ $Y2=0
cc_253 CLK N_A_30_99#_M1001_g 0.00597124f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_254 N_CLK_c_252_n N_A_30_99#_M1001_g 0.0114299f $X=0.625 $Y=1.19 $X2=0 $Y2=0
cc_255 N_CLK_c_253_n N_A_30_99#_M1001_g 0.00522735f $X=0.602 $Y=1.025 $X2=0
+ $Y2=0
cc_256 N_CLK_M1005_g N_A_30_99#_c_854_n 0.00666253f $X=0.645 $Y=2.645 $X2=0
+ $Y2=0
cc_257 CLK N_A_30_99#_c_854_n 0.106441f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_258 N_CLK_c_253_n N_A_30_99#_c_854_n 0.0203662f $X=0.602 $Y=1.025 $X2=0 $Y2=0
cc_259 N_CLK_M1005_g N_A_30_99#_c_869_n 2.23931e-19 $X=0.645 $Y=2.645 $X2=0
+ $Y2=0
cc_260 N_CLK_M1005_g N_A_30_99#_c_870_n 0.0101336f $X=0.645 $Y=2.645 $X2=0 $Y2=0
cc_261 N_CLK_c_250_n N_A_30_99#_c_870_n 4.60615e-19 $X=0.602 $Y=1.695 $X2=0
+ $Y2=0
cc_262 CLK N_A_30_99#_c_870_n 0.0226595f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_263 N_CLK_c_249_n N_A_30_99#_c_855_n 2.38298e-19 $X=0.602 $Y=1.508 $X2=0
+ $Y2=0
cc_264 N_CLK_M1005_g N_A_30_99#_c_855_n 0.00115789f $X=0.645 $Y=2.645 $X2=0
+ $Y2=0
cc_265 CLK N_A_30_99#_c_855_n 0.045751f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_266 N_CLK_c_249_n N_A_30_99#_c_856_n 0.00627853f $X=0.602 $Y=1.508 $X2=0
+ $Y2=0
cc_267 CLK N_A_30_99#_c_856_n 0.00397226f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_268 N_CLK_c_250_n N_A_30_99#_c_873_n 0.00336442f $X=0.602 $Y=1.695 $X2=0
+ $Y2=0
cc_269 N_CLK_M1005_g N_VPWR_c_1296_n 0.010927f $X=0.645 $Y=2.645 $X2=0 $Y2=0
cc_270 N_CLK_M1005_g N_VPWR_c_1317_n 0.00386543f $X=0.645 $Y=2.645 $X2=0 $Y2=0
cc_271 N_CLK_M1005_g N_VPWR_c_1295_n 0.00400158f $X=0.645 $Y=2.645 $X2=0 $Y2=0
cc_272 CLK N_VGND_M1013_d 0.00551703f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_273 CLK N_VGND_c_1622_n 0.0380544f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_274 N_CLK_c_253_n N_VGND_c_1622_n 0.00143165f $X=0.602 $Y=1.025 $X2=0 $Y2=0
cc_275 CLK N_VGND_c_1631_n 0.0111708f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_276 N_CLK_c_253_n N_VGND_c_1631_n 0.00459873f $X=0.602 $Y=1.025 $X2=0 $Y2=0
cc_277 CLK N_VGND_c_1645_n 0.0102313f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_278 N_CLK_c_253_n N_VGND_c_1645_n 0.00506877f $X=0.602 $Y=1.025 $X2=0 $Y2=0
cc_279 N_D_c_292_n N_A_230_465#_M1019_g 0.0170347f $X=2.44 $Y=2.13 $X2=0 $Y2=0
cc_280 D N_A_230_465#_M1019_g 6.7384e-19 $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_281 N_D_c_288_n N_A_230_465#_M1027_g 0.00144221f $X=2.23 $Y=1.2 $X2=0 $Y2=0
cc_282 D N_A_230_465#_c_357_n 0.0258441f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_283 N_D_c_295_n N_A_230_465#_c_357_n 0.00435208f $X=1.865 $Y=2.08 $X2=0 $Y2=0
cc_284 N_D_c_291_n N_A_230_465#_c_357_n 0.00338869f $X=1.865 $Y=1.915 $X2=0
+ $Y2=0
cc_285 N_D_c_288_n N_A_230_465#_c_346_n 0.00580301f $X=2.23 $Y=1.2 $X2=0 $Y2=0
cc_286 N_D_c_292_n N_A_230_465#_c_346_n 0.00258601f $X=2.44 $Y=2.13 $X2=0 $Y2=0
cc_287 D N_A_230_465#_c_346_n 0.0398977f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_288 N_D_c_295_n N_A_230_465#_c_346_n 0.00146958f $X=1.865 $Y=2.08 $X2=0 $Y2=0
cc_289 N_D_c_291_n N_A_230_465#_c_346_n 0.0150553f $X=1.865 $Y=1.915 $X2=0 $Y2=0
cc_290 N_D_c_290_n N_A_230_465#_c_347_n 0.00313795f $X=2.305 $Y=1.125 $X2=0
+ $Y2=0
cc_291 D N_A_230_465#_c_348_n 0.0036789f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_292 N_D_c_295_n N_A_230_465#_c_348_n 0.00415919f $X=1.865 $Y=2.08 $X2=0 $Y2=0
cc_293 N_D_c_288_n N_A_230_465#_c_349_n 0.0114656f $X=2.23 $Y=1.2 $X2=0 $Y2=0
cc_294 N_D_c_289_n N_A_230_465#_c_349_n 0.00473931f $X=2.03 $Y=1.2 $X2=0 $Y2=0
cc_295 N_D_c_291_n N_A_230_465#_c_349_n 0.0023102f $X=1.865 $Y=1.915 $X2=0 $Y2=0
cc_296 N_D_c_289_n N_A_230_465#_c_350_n 9.08494e-19 $X=2.03 $Y=1.2 $X2=0 $Y2=0
cc_297 N_D_c_291_n N_A_230_465#_c_350_n 8.22677e-19 $X=1.865 $Y=1.915 $X2=0
+ $Y2=0
cc_298 N_D_c_289_n N_A_230_465#_c_351_n 0.00834959f $X=2.03 $Y=1.2 $X2=0 $Y2=0
cc_299 N_D_c_288_n N_A_230_465#_c_352_n 0.00790592f $X=2.23 $Y=1.2 $X2=0 $Y2=0
cc_300 N_D_c_292_n N_A_230_465#_c_352_n 0.0183022f $X=2.44 $Y=2.13 $X2=0 $Y2=0
cc_301 D N_A_230_465#_c_352_n 4.86409e-19 $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_302 N_D_c_291_n N_A_230_465#_c_352_n 0.0184532f $X=1.865 $Y=1.915 $X2=0 $Y2=0
cc_303 N_D_c_295_n N_A_30_99#_c_857_n 0.00786636f $X=1.865 $Y=2.08 $X2=0 $Y2=0
cc_304 N_D_c_293_n N_A_30_99#_c_859_n 0.0103107f $X=2.515 $Y=2.205 $X2=0 $Y2=0
cc_305 N_D_c_289_n N_A_30_99#_M1001_g 0.00633944f $X=2.03 $Y=1.2 $X2=0 $Y2=0
cc_306 N_D_c_290_n N_A_30_99#_c_850_n 0.0104164f $X=2.305 $Y=1.125 $X2=0 $Y2=0
cc_307 N_D_c_290_n N_A_30_99#_M1002_g 0.0119551f $X=2.305 $Y=1.125 $X2=0 $Y2=0
cc_308 N_D_c_291_n N_A_30_99#_c_856_n 0.00633944f $X=1.865 $Y=1.915 $X2=0 $Y2=0
cc_309 N_D_c_292_n N_VPWR_c_1297_n 0.00347026f $X=2.44 $Y=2.13 $X2=0 $Y2=0
cc_310 N_D_c_293_n N_VPWR_c_1297_n 0.009325f $X=2.515 $Y=2.205 $X2=0 $Y2=0
cc_311 D N_VPWR_c_1297_n 0.0177532f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_312 N_D_c_293_n N_VPWR_c_1295_n 7.88961e-19 $X=2.515 $Y=2.205 $X2=0 $Y2=0
cc_313 N_D_c_290_n N_A_476_119#_c_1458_n 0.00103784f $X=2.305 $Y=1.125 $X2=0
+ $Y2=0
cc_314 N_D_c_293_n N_A_476_119#_c_1461_n 0.00194527f $X=2.515 $Y=2.205 $X2=0
+ $Y2=0
cc_315 N_D_c_290_n N_A_476_119#_c_1459_n 0.00341677f $X=2.305 $Y=1.125 $X2=0
+ $Y2=0
cc_316 N_D_c_288_n N_A_476_119#_c_1460_n 2.5815e-19 $X=2.23 $Y=1.2 $X2=0 $Y2=0
cc_317 N_D_c_292_n N_A_476_119#_c_1463_n 0.00194527f $X=2.44 $Y=2.13 $X2=0 $Y2=0
cc_318 D N_A_476_119#_c_1463_n 0.0184794f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_319 N_D_c_289_n N_VGND_c_1623_n 0.00595345f $X=2.03 $Y=1.2 $X2=0 $Y2=0
cc_320 N_D_c_290_n N_VGND_c_1623_n 0.00573363f $X=2.305 $Y=1.125 $X2=0 $Y2=0
cc_321 N_D_c_290_n N_VGND_c_1645_n 9.39239e-19 $X=2.305 $Y=1.125 $X2=0 $Y2=0
cc_322 N_A_230_465#_M1027_g N_A_690_93#_c_513_n 0.0603908f $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_323 N_A_230_465#_c_349_n N_A_690_93#_c_520_n 0.00163982f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_324 N_A_230_465#_c_349_n N_A_690_93#_c_514_n 0.0195529f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_325 N_A_230_465#_M1027_g N_A_690_93#_c_516_n 5.07813e-19 $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_326 N_A_230_465#_c_349_n N_A_690_93#_c_516_n 0.0213277f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_327 N_A_230_465#_c_349_n N_A_690_93#_c_517_n 0.00333286f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_328 N_A_230_465#_M1019_g N_A_690_93#_c_518_n 0.0059144f $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_329 N_A_230_465#_M1027_g N_A_690_93#_c_518_n 0.00447365f $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_330 N_A_230_465#_c_349_n N_SET_B_c_601_n 0.0387858f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_331 N_A_230_465#_c_399_p N_SET_B_c_601_n 7.06517e-19 $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_332 N_A_230_465#_c_353_n N_SET_B_c_601_n 0.0235549f $X=5.845 $Y=1.51 $X2=0
+ $Y2=0
cc_333 N_A_230_465#_c_349_n N_SET_B_c_611_n 8.15906e-19 $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_334 N_A_230_465#_c_349_n N_SET_B_c_612_n 0.0090884f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_335 N_A_230_465#_c_399_p N_SET_B_c_612_n 0.00139624f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_336 N_A_230_465#_c_353_n N_SET_B_c_612_n 0.0485061f $X=5.845 $Y=1.51 $X2=0
+ $Y2=0
cc_337 N_A_230_465#_c_354_n N_SET_B_c_612_n 0.0142067f $X=6.16 $Y=1.51 $X2=0
+ $Y2=0
cc_338 N_A_230_465#_M1018_g N_SET_B_c_603_n 0.00243307f $X=6.16 $Y=0.555 $X2=0
+ $Y2=0
cc_339 N_A_230_465#_M1036_g N_SET_B_c_603_n 0.0128519f $X=6.345 $Y=2.245 $X2=0
+ $Y2=0
cc_340 N_A_230_465#_c_399_p N_SET_B_c_603_n 3.13728e-19 $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_341 N_A_230_465#_c_353_n N_SET_B_c_603_n 0.0227064f $X=5.845 $Y=1.51 $X2=0
+ $Y2=0
cc_342 N_A_230_465#_c_354_n N_SET_B_c_603_n 0.0118216f $X=6.16 $Y=1.51 $X2=0
+ $Y2=0
cc_343 N_A_230_465#_M1036_g SET_B 0.00822448f $X=6.345 $Y=2.245 $X2=0 $Y2=0
cc_344 N_A_230_465#_c_354_n SET_B 0.00338654f $X=6.16 $Y=1.51 $X2=0 $Y2=0
cc_345 N_A_230_465#_c_349_n N_A_562_119#_M1007_g 0.00612695f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_346 N_A_230_465#_c_349_n N_A_562_119#_c_715_n 0.00271119f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_347 N_A_230_465#_M1018_g N_A_562_119#_c_716_n 0.00261287f $X=6.16 $Y=0.555
+ $X2=0 $Y2=0
cc_348 N_A_230_465#_c_349_n N_A_562_119#_c_716_n 0.00350816f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_349 N_A_230_465#_c_353_n N_A_562_119#_c_716_n 0.0103838f $X=5.845 $Y=1.51
+ $X2=0 $Y2=0
cc_350 N_A_230_465#_c_354_n N_A_562_119#_c_716_n 0.0215981f $X=6.16 $Y=1.51
+ $X2=0 $Y2=0
cc_351 N_A_230_465#_c_353_n N_A_562_119#_M1020_g 0.00164381f $X=5.845 $Y=1.51
+ $X2=0 $Y2=0
cc_352 N_A_230_465#_c_353_n N_A_562_119#_c_718_n 0.0098714f $X=5.845 $Y=1.51
+ $X2=0 $Y2=0
cc_353 N_A_230_465#_c_354_n N_A_562_119#_c_718_n 0.0123946f $X=6.16 $Y=1.51
+ $X2=0 $Y2=0
cc_354 N_A_230_465#_M1018_g N_A_562_119#_c_720_n 0.0622402f $X=6.16 $Y=0.555
+ $X2=0 $Y2=0
cc_355 N_A_230_465#_c_353_n N_A_562_119#_c_721_n 0.00551683f $X=5.845 $Y=1.51
+ $X2=0 $Y2=0
cc_356 N_A_230_465#_M1027_g N_A_562_119#_c_722_n 0.0123374f $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_357 N_A_230_465#_c_345_n N_A_562_119#_c_722_n 0.00219912f $X=3.165 $Y=1.56
+ $X2=0 $Y2=0
cc_358 N_A_230_465#_c_349_n N_A_562_119#_c_722_n 0.0167692f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_359 N_A_230_465#_c_349_n N_A_562_119#_c_723_n 0.019355f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_360 N_A_230_465#_M1027_g N_A_562_119#_c_724_n 0.00919626f $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_361 N_A_230_465#_c_345_n N_A_562_119#_c_724_n 0.00301787f $X=3.165 $Y=1.56
+ $X2=0 $Y2=0
cc_362 N_A_230_465#_c_349_n N_A_562_119#_c_724_n 0.00862887f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_363 N_A_230_465#_M1019_g N_A_562_119#_c_730_n 2.23879e-19 $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_364 N_A_230_465#_c_345_n N_A_562_119#_c_730_n 0.00233075f $X=3.165 $Y=1.56
+ $X2=0 $Y2=0
cc_365 N_A_230_465#_M1019_g N_A_562_119#_c_731_n 0.00556012f $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_366 N_A_230_465#_M1019_g N_A_562_119#_c_732_n 9.92457e-19 $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_367 N_A_230_465#_c_345_n N_A_562_119#_c_732_n 0.00608487f $X=3.165 $Y=1.56
+ $X2=0 $Y2=0
cc_368 N_A_230_465#_c_349_n N_A_562_119#_c_725_n 0.010265f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_369 N_A_230_465#_c_349_n N_A_562_119#_c_726_n 0.00846729f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_370 N_A_230_465#_c_357_n N_A_30_99#_c_857_n 0.00402267f $X=1.515 $Y=2.64
+ $X2=0 $Y2=0
cc_371 N_A_230_465#_c_357_n N_A_30_99#_M1025_g 0.00589423f $X=1.515 $Y=2.64
+ $X2=0 $Y2=0
cc_372 N_A_230_465#_M1019_g N_A_30_99#_c_859_n 0.0104164f $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_373 N_A_230_465#_c_359_n N_A_30_99#_c_859_n 0.00814764f $X=1.515 $Y=2.805
+ $X2=0 $Y2=0
cc_374 N_A_230_465#_c_347_n N_A_30_99#_M1001_g 8.97897e-19 $X=1.5 $Y=0.705 $X2=0
+ $Y2=0
cc_375 N_A_230_465#_c_348_n N_A_30_99#_M1001_g 0.00320088f $X=1.622 $Y=1.615
+ $X2=0 $Y2=0
cc_376 N_A_230_465#_c_351_n N_A_30_99#_M1001_g 0.0113711f $X=1.68 $Y=1.295 $X2=0
+ $Y2=0
cc_377 N_A_230_465#_c_347_n N_A_30_99#_c_850_n 0.00759179f $X=1.5 $Y=0.705 $X2=0
+ $Y2=0
cc_378 N_A_230_465#_c_340_n N_A_30_99#_M1002_g 0.00486943f $X=2.87 $Y=1.56 $X2=0
+ $Y2=0
cc_379 N_A_230_465#_M1027_g N_A_30_99#_M1002_g 0.0145242f $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_380 N_A_230_465#_M1019_g N_A_30_99#_M1000_g 0.0124449f $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_381 N_A_230_465#_M1036_g N_A_30_99#_c_862_n 0.00262437f $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_382 N_A_230_465#_M1018_g N_A_30_99#_M1021_g 0.0221782f $X=6.16 $Y=0.555 $X2=0
+ $Y2=0
cc_383 N_A_230_465#_c_354_n N_A_30_99#_M1021_g 0.0177004f $X=6.16 $Y=1.51 $X2=0
+ $Y2=0
cc_384 N_A_230_465#_M1036_g N_A_30_99#_M1026_g 0.014804f $X=6.345 $Y=2.245 $X2=0
+ $Y2=0
cc_385 N_A_230_465#_c_359_n N_A_30_99#_c_865_n 0.00346325f $X=1.515 $Y=2.805
+ $X2=0 $Y2=0
cc_386 N_A_230_465#_M1036_g N_A_30_99#_c_867_n 0.0177004f $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_387 N_A_230_465#_M1025_d N_A_30_99#_c_870_n 0.00217079f $X=1.15 $Y=2.325
+ $X2=0 $Y2=0
cc_388 N_A_230_465#_c_357_n N_A_30_99#_c_870_n 0.0141004f $X=1.515 $Y=2.64 $X2=0
+ $Y2=0
cc_389 N_A_230_465#_c_359_n N_A_30_99#_c_870_n 0.0044056f $X=1.515 $Y=2.805
+ $X2=0 $Y2=0
cc_390 N_A_230_465#_c_357_n N_A_30_99#_c_855_n 0.0413865f $X=1.515 $Y=2.64 $X2=0
+ $Y2=0
cc_391 N_A_230_465#_c_348_n N_A_30_99#_c_855_n 0.0207061f $X=1.622 $Y=1.615
+ $X2=0 $Y2=0
cc_392 N_A_230_465#_M1018_g N_A_1247_47#_c_1088_n 0.0170917f $X=6.16 $Y=0.555
+ $X2=0 $Y2=0
cc_393 N_A_230_465#_M1018_g N_A_1247_47#_c_1089_n 0.00616991f $X=6.16 $Y=0.555
+ $X2=0 $Y2=0
cc_394 N_A_230_465#_c_354_n N_A_1247_47#_c_1089_n 0.00128241f $X=6.16 $Y=1.51
+ $X2=0 $Y2=0
cc_395 N_A_230_465#_M1036_g N_A_1247_47#_c_1102_n 0.00447464f $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_396 N_A_230_465#_c_359_n N_VPWR_c_1296_n 0.0124952f $X=1.515 $Y=2.805 $X2=0
+ $Y2=0
cc_397 N_A_230_465#_M1019_g N_VPWR_c_1297_n 8.66328e-19 $X=2.945 $Y=2.525 $X2=0
+ $Y2=0
cc_398 N_A_230_465#_c_357_n N_VPWR_c_1297_n 0.0080616f $X=1.515 $Y=2.64 $X2=0
+ $Y2=0
cc_399 N_A_230_465#_c_346_n N_VPWR_c_1297_n 0.00240946f $X=2.435 $Y=1.65 $X2=0
+ $Y2=0
cc_400 N_A_230_465#_c_359_n N_VPWR_c_1297_n 0.0125581f $X=1.515 $Y=2.805 $X2=0
+ $Y2=0
cc_401 N_A_230_465#_c_359_n N_VPWR_c_1313_n 0.0164226f $X=1.515 $Y=2.805 $X2=0
+ $Y2=0
cc_402 N_A_230_465#_M1019_g N_VPWR_c_1295_n 9.39239e-19 $X=2.945 $Y=2.525 $X2=0
+ $Y2=0
cc_403 N_A_230_465#_c_359_n N_VPWR_c_1295_n 0.0128812f $X=1.515 $Y=2.805 $X2=0
+ $Y2=0
cc_404 N_A_230_465#_c_349_n N_A_476_119#_c_1458_n 0.00142378f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_405 N_A_230_465#_c_351_n N_A_476_119#_c_1458_n 0.00324369f $X=1.68 $Y=1.295
+ $X2=0 $Y2=0
cc_406 N_A_230_465#_M1019_g N_A_476_119#_c_1461_n 0.00223916f $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_407 N_A_230_465#_c_340_n N_A_476_119#_c_1459_n 5.85719e-19 $X=2.87 $Y=1.56
+ $X2=0 $Y2=0
cc_408 N_A_230_465#_M1027_g N_A_476_119#_c_1459_n 0.00151488f $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_409 N_A_230_465#_c_346_n N_A_476_119#_c_1459_n 0.00939313f $X=2.435 $Y=1.65
+ $X2=0 $Y2=0
cc_410 N_A_230_465#_c_349_n N_A_476_119#_c_1459_n 0.0158922f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_411 N_A_230_465#_c_350_n N_A_476_119#_c_1459_n 0.00104488f $X=1.825 $Y=1.295
+ $X2=0 $Y2=0
cc_412 N_A_230_465#_c_351_n N_A_476_119#_c_1459_n 0.00492759f $X=1.68 $Y=1.295
+ $X2=0 $Y2=0
cc_413 N_A_230_465#_c_352_n N_A_476_119#_c_1459_n 0.00678853f $X=2.435 $Y=1.56
+ $X2=0 $Y2=0
cc_414 N_A_230_465#_c_340_n N_A_476_119#_c_1460_n 0.00678326f $X=2.87 $Y=1.56
+ $X2=0 $Y2=0
cc_415 N_A_230_465#_M1019_g N_A_476_119#_c_1460_n 0.00665476f $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_416 N_A_230_465#_M1027_g N_A_476_119#_c_1460_n 0.0039897f $X=3.165 $Y=0.805
+ $X2=0 $Y2=0
cc_417 N_A_230_465#_c_345_n N_A_476_119#_c_1460_n 0.00472402f $X=3.165 $Y=1.56
+ $X2=0 $Y2=0
cc_418 N_A_230_465#_c_346_n N_A_476_119#_c_1460_n 0.0191788f $X=2.435 $Y=1.65
+ $X2=0 $Y2=0
cc_419 N_A_230_465#_c_349_n N_A_476_119#_c_1460_n 0.0113446f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_420 N_A_230_465#_c_352_n N_A_476_119#_c_1460_n 0.00183048f $X=2.435 $Y=1.56
+ $X2=0 $Y2=0
cc_421 N_A_230_465#_c_340_n N_A_476_119#_c_1463_n 0.00332614f $X=2.87 $Y=1.56
+ $X2=0 $Y2=0
cc_422 N_A_230_465#_M1019_g N_A_476_119#_c_1463_n 0.00951851f $X=2.945 $Y=2.525
+ $X2=0 $Y2=0
cc_423 N_A_230_465#_c_349_n N_A_476_119#_c_1463_n 0.00320368f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_424 N_A_230_465#_M1036_g N_A_1094_379#_c_1506_n 0.00109574f $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_425 N_A_230_465#_M1036_g N_A_1094_379#_c_1508_n 4.34847e-19 $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_426 N_A_230_465#_M1036_g N_A_1201_407#_c_1533_n 0.00824985f $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_427 N_A_230_465#_c_354_n N_A_1201_407#_c_1533_n 2.24398e-19 $X=6.16 $Y=1.51
+ $X2=0 $Y2=0
cc_428 N_A_230_465#_M1036_g N_A_1201_407#_c_1534_n 0.00739251f $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_429 N_A_230_465#_M1036_g N_A_1201_407#_c_1535_n 0.00161284f $X=6.345 $Y=2.245
+ $X2=0 $Y2=0
cc_430 N_A_230_465#_c_346_n N_VGND_c_1623_n 0.00342779f $X=2.435 $Y=1.65 $X2=0
+ $Y2=0
cc_431 N_A_230_465#_c_347_n N_VGND_c_1623_n 0.0351477f $X=1.5 $Y=0.705 $X2=0
+ $Y2=0
cc_432 N_A_230_465#_c_349_n N_VGND_c_1623_n 0.00608029f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_433 N_A_230_465#_M1027_g N_VGND_c_1624_n 0.00329607f $X=3.165 $Y=0.805 $X2=0
+ $Y2=0
cc_434 N_A_230_465#_M1027_g N_VGND_c_1625_n 8.26459e-19 $X=3.165 $Y=0.805 $X2=0
+ $Y2=0
cc_435 N_A_230_465#_c_349_n N_VGND_c_1625_n 0.00118069f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_436 N_A_230_465#_c_347_n N_VGND_c_1635_n 0.0102224f $X=1.5 $Y=0.705 $X2=0
+ $Y2=0
cc_437 N_A_230_465#_M1018_g N_VGND_c_1637_n 0.0054895f $X=6.16 $Y=0.555 $X2=0
+ $Y2=0
cc_438 N_A_230_465#_M1018_g N_VGND_c_1642_n 0.00301978f $X=6.16 $Y=0.555 $X2=0
+ $Y2=0
cc_439 N_A_230_465#_c_349_n N_VGND_c_1642_n 0.00968962f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_440 N_A_230_465#_c_399_p N_VGND_c_1642_n 0.00225748f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_441 N_A_230_465#_c_353_n N_VGND_c_1642_n 0.0204898f $X=5.845 $Y=1.51 $X2=0
+ $Y2=0
cc_442 N_A_230_465#_M1027_g N_VGND_c_1645_n 0.00477801f $X=3.165 $Y=0.805 $X2=0
+ $Y2=0
cc_443 N_A_230_465#_M1018_g N_VGND_c_1645_n 0.0111524f $X=6.16 $Y=0.555 $X2=0
+ $Y2=0
cc_444 N_A_230_465#_c_347_n N_VGND_c_1645_n 0.012461f $X=1.5 $Y=0.705 $X2=0
+ $Y2=0
cc_445 N_A_690_93#_c_532_p N_SET_B_M1003_g 0.00650213f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_446 N_A_690_93#_c_522_n N_SET_B_M1003_g 0.00160565f $X=4.482 $Y=2.325 $X2=0
+ $Y2=0
cc_447 N_A_690_93#_c_514_n N_SET_B_c_601_n 0.0128863f $X=4.115 $Y=1.07 $X2=0
+ $Y2=0
cc_448 N_A_690_93#_c_515_n N_SET_B_c_601_n 0.0147331f $X=4.28 $Y=0.45 $X2=0
+ $Y2=0
cc_449 N_A_690_93#_c_520_n N_SET_B_c_610_n 0.0215956f $X=4.305 $Y=2.025 $X2=0
+ $Y2=0
cc_450 N_A_690_93#_c_532_p N_SET_B_c_610_n 0.00113158f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_451 N_A_690_93#_c_520_n N_SET_B_c_611_n 0.00187038f $X=4.305 $Y=2.025 $X2=0
+ $Y2=0
cc_452 N_A_690_93#_c_532_p N_SET_B_c_611_n 0.00168675f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_453 N_A_690_93#_c_515_n N_SET_B_c_605_n 0.00173672f $X=4.28 $Y=0.45 $X2=0
+ $Y2=0
cc_454 N_A_690_93#_M1006_g N_A_562_119#_M1016_g 0.0134634f $X=3.735 $Y=2.525
+ $X2=0 $Y2=0
cc_455 N_A_690_93#_c_520_n N_A_562_119#_M1016_g 0.0139557f $X=4.305 $Y=2.025
+ $X2=0 $Y2=0
cc_456 N_A_690_93#_c_521_n N_A_562_119#_M1016_g 0.0209683f $X=3.825 $Y=1.99
+ $X2=0 $Y2=0
cc_457 N_A_690_93#_c_532_p N_A_562_119#_M1016_g 0.0055379f $X=4.495 $Y=2.525
+ $X2=0 $Y2=0
cc_458 N_A_690_93#_c_522_n N_A_562_119#_M1016_g 0.00457654f $X=4.482 $Y=2.325
+ $X2=0 $Y2=0
cc_459 N_A_690_93#_c_518_n N_A_562_119#_M1016_g 0.00763805f $X=3.825 $Y=1.825
+ $X2=0 $Y2=0
cc_460 N_A_690_93#_c_514_n N_A_562_119#_M1007_g 0.00600597f $X=4.115 $Y=1.07
+ $X2=0 $Y2=0
cc_461 N_A_690_93#_c_515_n N_A_562_119#_M1007_g 0.0173835f $X=4.28 $Y=0.45 $X2=0
+ $Y2=0
cc_462 N_A_690_93#_c_516_n N_A_562_119#_M1007_g 8.31653e-19 $X=3.645 $Y=1.07
+ $X2=0 $Y2=0
cc_463 N_A_690_93#_c_517_n N_A_562_119#_M1007_g 0.00247751f $X=3.735 $Y=1.29
+ $X2=0 $Y2=0
cc_464 N_A_690_93#_c_513_n N_A_562_119#_c_722_n 0.00489262f $X=3.525 $Y=1.125
+ $X2=0 $Y2=0
cc_465 N_A_690_93#_c_516_n N_A_562_119#_c_722_n 0.0275907f $X=3.645 $Y=1.07
+ $X2=0 $Y2=0
cc_466 N_A_690_93#_c_518_n N_A_562_119#_c_722_n 0.00173517f $X=3.825 $Y=1.825
+ $X2=0 $Y2=0
cc_467 N_A_690_93#_c_520_n N_A_562_119#_c_723_n 0.0339504f $X=4.305 $Y=2.025
+ $X2=0 $Y2=0
cc_468 N_A_690_93#_c_521_n N_A_562_119#_c_723_n 0.00438376f $X=3.825 $Y=1.99
+ $X2=0 $Y2=0
cc_469 N_A_690_93#_c_514_n N_A_562_119#_c_723_n 0.00678611f $X=4.115 $Y=1.07
+ $X2=0 $Y2=0
cc_470 N_A_690_93#_c_516_n N_A_562_119#_c_723_n 0.0224531f $X=3.645 $Y=1.07
+ $X2=0 $Y2=0
cc_471 N_A_690_93#_c_517_n N_A_562_119#_c_723_n 0.00625126f $X=3.735 $Y=1.29
+ $X2=0 $Y2=0
cc_472 N_A_690_93#_c_518_n N_A_562_119#_c_723_n 0.0114843f $X=3.825 $Y=1.825
+ $X2=0 $Y2=0
cc_473 N_A_690_93#_c_513_n N_A_562_119#_c_724_n 0.00413697f $X=3.525 $Y=1.125
+ $X2=0 $Y2=0
cc_474 N_A_690_93#_c_520_n N_A_562_119#_c_731_n 0.011725f $X=4.305 $Y=2.025
+ $X2=0 $Y2=0
cc_475 N_A_690_93#_c_521_n N_A_562_119#_c_731_n 0.00253402f $X=3.825 $Y=1.99
+ $X2=0 $Y2=0
cc_476 N_A_690_93#_c_518_n N_A_562_119#_c_731_n 0.00328764f $X=3.825 $Y=1.825
+ $X2=0 $Y2=0
cc_477 N_A_690_93#_c_520_n N_A_562_119#_c_725_n 0.0262847f $X=4.305 $Y=2.025
+ $X2=0 $Y2=0
cc_478 N_A_690_93#_c_514_n N_A_562_119#_c_725_n 0.0214981f $X=4.115 $Y=1.07
+ $X2=0 $Y2=0
cc_479 N_A_690_93#_c_516_n N_A_562_119#_c_725_n 0.00211591f $X=3.645 $Y=1.07
+ $X2=0 $Y2=0
cc_480 N_A_690_93#_c_517_n N_A_562_119#_c_725_n 0.00130835f $X=3.735 $Y=1.29
+ $X2=0 $Y2=0
cc_481 N_A_690_93#_c_520_n N_A_562_119#_c_726_n 9.1978e-19 $X=4.305 $Y=2.025
+ $X2=0 $Y2=0
cc_482 N_A_690_93#_c_514_n N_A_562_119#_c_726_n 0.00617004f $X=4.115 $Y=1.07
+ $X2=0 $Y2=0
cc_483 N_A_690_93#_c_516_n N_A_562_119#_c_726_n 9.05892e-19 $X=3.645 $Y=1.07
+ $X2=0 $Y2=0
cc_484 N_A_690_93#_c_517_n N_A_562_119#_c_726_n 0.0142083f $X=3.735 $Y=1.29
+ $X2=0 $Y2=0
cc_485 N_A_690_93#_M1006_g N_A_30_99#_M1000_g 0.0403652f $X=3.735 $Y=2.525 $X2=0
+ $Y2=0
cc_486 N_A_690_93#_M1006_g N_A_30_99#_c_862_n 0.0104018f $X=3.735 $Y=2.525 $X2=0
+ $Y2=0
cc_487 N_A_690_93#_c_532_p N_A_30_99#_c_862_n 0.0048403f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_488 N_A_690_93#_M1006_g N_VPWR_c_1298_n 0.00973884f $X=3.735 $Y=2.525 $X2=0
+ $Y2=0
cc_489 N_A_690_93#_c_520_n N_VPWR_c_1298_n 0.0213738f $X=4.305 $Y=2.025 $X2=0
+ $Y2=0
cc_490 N_A_690_93#_c_521_n N_VPWR_c_1298_n 0.00392572f $X=3.825 $Y=1.99 $X2=0
+ $Y2=0
cc_491 N_A_690_93#_c_532_p N_VPWR_c_1298_n 0.0257553f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_492 N_A_690_93#_c_532_p N_VPWR_c_1299_n 0.00544268f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_493 N_A_690_93#_c_532_p N_VPWR_c_1300_n 0.0158879f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_494 N_A_690_93#_c_522_n N_VPWR_c_1300_n 0.00582606f $X=4.482 $Y=2.325 $X2=0
+ $Y2=0
cc_495 N_A_690_93#_M1006_g N_VPWR_c_1295_n 9.14192e-19 $X=3.735 $Y=2.525 $X2=0
+ $Y2=0
cc_496 N_A_690_93#_c_532_p N_VPWR_c_1295_n 0.00901867f $X=4.495 $Y=2.525 $X2=0
+ $Y2=0
cc_497 N_A_690_93#_c_514_n N_VGND_M1035_d 8.68247e-19 $X=4.115 $Y=1.07 $X2=0
+ $Y2=0
cc_498 N_A_690_93#_c_516_n N_VGND_M1035_d 0.00173531f $X=3.645 $Y=1.07 $X2=0
+ $Y2=0
cc_499 N_A_690_93#_c_513_n N_VGND_c_1624_n 0.0035863f $X=3.525 $Y=1.125 $X2=0
+ $Y2=0
cc_500 N_A_690_93#_c_513_n N_VGND_c_1625_n 0.00840033f $X=3.525 $Y=1.125 $X2=0
+ $Y2=0
cc_501 N_A_690_93#_c_514_n N_VGND_c_1625_n 0.00729832f $X=4.115 $Y=1.07 $X2=0
+ $Y2=0
cc_502 N_A_690_93#_c_515_n N_VGND_c_1625_n 0.0380585f $X=4.28 $Y=0.45 $X2=0
+ $Y2=0
cc_503 N_A_690_93#_c_516_n N_VGND_c_1625_n 0.0143553f $X=3.645 $Y=1.07 $X2=0
+ $Y2=0
cc_504 N_A_690_93#_c_517_n N_VGND_c_1625_n 0.00103664f $X=3.735 $Y=1.29 $X2=0
+ $Y2=0
cc_505 N_A_690_93#_c_515_n N_VGND_c_1636_n 0.0176612f $X=4.28 $Y=0.45 $X2=0
+ $Y2=0
cc_506 N_A_690_93#_c_515_n N_VGND_c_1642_n 0.0115331f $X=4.28 $Y=0.45 $X2=0
+ $Y2=0
cc_507 N_A_690_93#_M1007_s N_VGND_c_1645_n 0.002172f $X=4.155 $Y=0.235 $X2=0
+ $Y2=0
cc_508 N_A_690_93#_c_513_n N_VGND_c_1645_n 0.00401353f $X=3.525 $Y=1.125 $X2=0
+ $Y2=0
cc_509 N_A_690_93#_c_515_n N_VGND_c_1645_n 0.0124419f $X=4.28 $Y=0.45 $X2=0
+ $Y2=0
cc_510 N_SET_B_M1003_g N_A_562_119#_M1016_g 0.013392f $X=4.71 $Y=2.525 $X2=0
+ $Y2=0
cc_511 N_SET_B_c_601_n N_A_562_119#_M1016_g 0.00216007f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_512 N_SET_B_c_610_n N_A_562_119#_M1016_g 0.00278161f $X=5.11 $Y=1.85 $X2=0
+ $Y2=0
cc_513 N_SET_B_c_611_n N_A_562_119#_M1016_g 0.020573f $X=4.73 $Y=1.99 $X2=0
+ $Y2=0
cc_514 N_SET_B_c_601_n N_A_562_119#_M1007_g 0.012725f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_515 N_SET_B_c_605_n N_A_562_119#_M1007_g 0.059964f $X=4.945 $Y=0.775 $X2=0
+ $Y2=0
cc_516 N_SET_B_c_601_n N_A_562_119#_c_715_n 0.0255302f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_517 N_SET_B_c_602_n N_A_562_119#_c_715_n 0.0120691f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_518 N_SET_B_c_612_n N_A_562_119#_c_715_n 0.00404713f $X=6.18 $Y=1.63 $X2=0
+ $Y2=0
cc_519 N_SET_B_M1003_g N_A_562_119#_M1020_g 0.00578083f $X=4.71 $Y=2.525 $X2=0
+ $Y2=0
cc_520 N_SET_B_c_601_n N_A_562_119#_M1020_g 0.0064889f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_521 N_SET_B_c_610_n N_A_562_119#_M1020_g 8.13102e-19 $X=5.11 $Y=1.85 $X2=0
+ $Y2=0
cc_522 N_SET_B_c_611_n N_A_562_119#_M1020_g 0.00830808f $X=4.73 $Y=1.99 $X2=0
+ $Y2=0
cc_523 N_SET_B_c_612_n N_A_562_119#_M1020_g 0.0178021f $X=6.18 $Y=1.63 $X2=0
+ $Y2=0
cc_524 N_SET_B_c_601_n N_A_562_119#_c_719_n 0.00772659f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_525 N_SET_B_c_602_n N_A_562_119#_c_719_n 0.00841384f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_526 N_SET_B_c_601_n N_A_562_119#_c_720_n 5.24671e-19 $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_527 N_SET_B_c_602_n N_A_562_119#_c_720_n 0.0029115f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_528 N_SET_B_c_601_n N_A_562_119#_c_725_n 0.0305912f $X=4.945 $Y=0.94 $X2=0
+ $Y2=0
cc_529 N_SET_B_c_611_n N_A_562_119#_c_726_n 0.0192183f $X=4.73 $Y=1.99 $X2=0
+ $Y2=0
cc_530 N_SET_B_M1003_g N_A_30_99#_c_862_n 0.0103162f $X=4.71 $Y=2.525 $X2=0
+ $Y2=0
cc_531 SET_B N_A_30_99#_M1021_g 0.0194598f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_532 N_SET_B_c_603_n N_A_30_99#_c_867_n 5.37053e-19 $X=6.35 $Y=1.63 $X2=0
+ $Y2=0
cc_533 SET_B N_A_30_99#_c_867_n 0.0103806f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_534 N_SET_B_c_597_n N_A_1398_65#_M1008_g 0.049823f $X=7.425 $Y=0.985 $X2=0
+ $Y2=0
cc_535 N_SET_B_c_600_n N_A_1398_65#_M1008_g 0.00588534f $X=8.375 $Y=1.915 $X2=0
+ $Y2=0
cc_536 SET_B N_A_1398_65#_M1008_g 0.00480385f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_537 N_SET_B_c_599_n N_A_1398_65#_c_988_n 0.00937621f $X=7.5 $Y=1.06 $X2=0
+ $Y2=0
cc_538 N_SET_B_c_600_n N_A_1398_65#_c_988_n 0.0352136f $X=8.375 $Y=1.915 $X2=0
+ $Y2=0
cc_539 SET_B N_A_1398_65#_c_988_n 0.0155671f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_540 SET_B N_A_1398_65#_c_989_n 0.00650599f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_541 SET_B N_A_1398_65#_c_990_n 0.0146667f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_542 N_SET_B_c_600_n N_A_1398_65#_M1014_g 0.00828166f $X=8.375 $Y=1.915 $X2=0
+ $Y2=0
cc_543 N_SET_B_M1032_g N_A_1398_65#_M1014_g 0.0132048f $X=8.375 $Y=2.495 $X2=0
+ $Y2=0
cc_544 N_SET_B_M1032_g N_A_1398_65#_c_999_n 0.00894529f $X=8.375 $Y=2.495 $X2=0
+ $Y2=0
cc_545 N_SET_B_c_600_n N_A_1247_47#_c_1079_n 0.00945476f $X=8.375 $Y=1.915 $X2=0
+ $Y2=0
cc_546 N_SET_B_c_597_n N_A_1247_47#_c_1081_n 0.00465384f $X=7.425 $Y=0.985 $X2=0
+ $Y2=0
cc_547 N_SET_B_c_603_n N_A_1247_47#_c_1089_n 0.0394568f $X=6.35 $Y=1.63 $X2=0
+ $Y2=0
cc_548 N_SET_B_c_600_n N_A_1247_47#_c_1099_n 0.0127721f $X=8.375 $Y=1.915 $X2=0
+ $Y2=0
cc_549 N_SET_B_M1032_g N_A_1247_47#_c_1099_n 0.0174712f $X=8.375 $Y=2.495 $X2=0
+ $Y2=0
cc_550 SET_B N_A_1247_47#_c_1099_n 0.12713f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_551 N_SET_B_M1032_g N_A_1247_47#_c_1100_n 0.00451166f $X=8.375 $Y=2.495 $X2=0
+ $Y2=0
cc_552 N_SET_B_c_600_n N_A_1247_47#_c_1090_n 0.0130019f $X=8.375 $Y=1.915 $X2=0
+ $Y2=0
cc_553 SET_B N_A_1247_47#_c_1090_n 0.0430671f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_554 SET_B N_A_1247_47#_c_1102_n 0.0219994f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_555 N_SET_B_c_597_n N_A_1247_47#_c_1093_n 0.00689717f $X=7.425 $Y=0.985 $X2=0
+ $Y2=0
cc_556 N_SET_B_c_598_n N_A_1247_47#_c_1093_n 0.00794724f $X=7.74 $Y=1.06 $X2=0
+ $Y2=0
cc_557 N_SET_B_c_599_n N_A_1247_47#_c_1093_n 0.00402599f $X=7.5 $Y=1.06 $X2=0
+ $Y2=0
cc_558 N_SET_B_c_600_n N_A_1247_47#_c_1093_n 0.0221466f $X=8.375 $Y=1.915 $X2=0
+ $Y2=0
cc_559 SET_B N_A_1247_47#_c_1093_n 0.12319f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_560 N_SET_B_c_610_n N_VPWR_M1003_d 6.86134e-19 $X=5.11 $Y=1.85 $X2=0 $Y2=0
cc_561 N_SET_B_c_612_n N_VPWR_M1003_d 0.00167839f $X=6.18 $Y=1.63 $X2=0 $Y2=0
cc_562 N_SET_B_M1003_g N_VPWR_c_1300_n 0.00935574f $X=4.71 $Y=2.525 $X2=0 $Y2=0
cc_563 N_SET_B_c_610_n N_VPWR_c_1300_n 0.0123766f $X=5.11 $Y=1.85 $X2=0 $Y2=0
cc_564 N_SET_B_c_611_n N_VPWR_c_1300_n 4.49476e-19 $X=4.73 $Y=1.99 $X2=0 $Y2=0
cc_565 N_SET_B_c_612_n N_VPWR_c_1300_n 0.0124114f $X=6.18 $Y=1.63 $X2=0 $Y2=0
cc_566 N_SET_B_M1032_g N_VPWR_c_1301_n 0.0131227f $X=8.375 $Y=2.495 $X2=0 $Y2=0
cc_567 N_SET_B_M1032_g N_VPWR_c_1302_n 0.00524649f $X=8.375 $Y=2.495 $X2=0 $Y2=0
cc_568 N_SET_B_M1003_g N_VPWR_c_1295_n 9.39239e-19 $X=4.71 $Y=2.525 $X2=0 $Y2=0
cc_569 N_SET_B_M1032_g N_VPWR_c_1295_n 7.97988e-19 $X=8.375 $Y=2.495 $X2=0 $Y2=0
cc_570 N_SET_B_c_612_n N_A_1094_379#_M1020_d 0.00239457f $X=6.18 $Y=1.63
+ $X2=-0.19 $Y2=-0.245
cc_571 N_SET_B_c_612_n N_A_1094_379#_c_1506_n 0.0220025f $X=6.18 $Y=1.63 $X2=0
+ $Y2=0
cc_572 N_SET_B_c_612_n N_A_1201_407#_c_1533_n 0.0250457f $X=6.18 $Y=1.63 $X2=0
+ $Y2=0
cc_573 N_SET_B_c_603_n N_A_1201_407#_c_1534_n 0.00146619f $X=6.35 $Y=1.63 $X2=0
+ $Y2=0
cc_574 N_SET_B_c_597_n N_VGND_c_1626_n 0.0120566f $X=7.425 $Y=0.985 $X2=0 $Y2=0
cc_575 N_SET_B_c_598_n N_VGND_c_1626_n 0.00268383f $X=7.74 $Y=1.06 $X2=0 $Y2=0
cc_576 N_SET_B_c_605_n N_VGND_c_1636_n 0.00486043f $X=4.945 $Y=0.775 $X2=0 $Y2=0
cc_577 N_SET_B_c_597_n N_VGND_c_1637_n 0.00429764f $X=7.425 $Y=0.985 $X2=0 $Y2=0
cc_578 N_SET_B_c_601_n N_VGND_c_1642_n 0.0198211f $X=4.945 $Y=0.94 $X2=0 $Y2=0
cc_579 N_SET_B_c_602_n N_VGND_c_1642_n 0.00516611f $X=4.945 $Y=0.94 $X2=0 $Y2=0
cc_580 N_SET_B_c_605_n N_VGND_c_1642_n 0.0172703f $X=4.945 $Y=0.775 $X2=0 $Y2=0
cc_581 N_SET_B_c_597_n N_VGND_c_1645_n 0.00435987f $X=7.425 $Y=0.985 $X2=0 $Y2=0
cc_582 N_SET_B_c_601_n N_VGND_c_1645_n 0.0105322f $X=4.945 $Y=0.94 $X2=0 $Y2=0
cc_583 N_SET_B_c_605_n N_VGND_c_1645_n 0.00430516f $X=4.945 $Y=0.775 $X2=0 $Y2=0
cc_584 N_A_562_119#_c_730_n N_A_30_99#_c_859_n 0.00308102f $X=3.16 $Y=2.525
+ $X2=0 $Y2=0
cc_585 N_A_562_119#_c_722_n N_A_30_99#_M1002_g 5.72651e-19 $X=3.215 $Y=1.555
+ $X2=0 $Y2=0
cc_586 N_A_562_119#_c_723_n N_A_30_99#_M1000_g 0.00457527f $X=4.135 $Y=1.64
+ $X2=0 $Y2=0
cc_587 N_A_562_119#_c_731_n N_A_30_99#_M1000_g 0.00340148f $X=3.167 $Y=2.295
+ $X2=0 $Y2=0
cc_588 N_A_562_119#_M1016_g N_A_30_99#_c_862_n 0.0102119f $X=4.28 $Y=2.525 $X2=0
+ $Y2=0
cc_589 N_A_562_119#_M1020_g N_A_30_99#_c_862_n 0.0101457f $X=5.395 $Y=2.315
+ $X2=0 $Y2=0
cc_590 N_A_562_119#_c_720_n N_A_1247_47#_c_1088_n 0.00205415f $X=5.8 $Y=0.985
+ $X2=0 $Y2=0
cc_591 N_A_562_119#_c_720_n N_A_1247_47#_c_1089_n 9.33767e-19 $X=5.8 $Y=0.985
+ $X2=0 $Y2=0
cc_592 N_A_562_119#_M1016_g N_VPWR_c_1298_n 0.00774805f $X=4.28 $Y=2.525 $X2=0
+ $Y2=0
cc_593 N_A_562_119#_c_730_n N_VPWR_c_1298_n 0.0112789f $X=3.16 $Y=2.525 $X2=0
+ $Y2=0
cc_594 N_A_562_119#_c_715_n N_VPWR_c_1300_n 5.62536e-19 $X=5.32 $Y=1.51 $X2=0
+ $Y2=0
cc_595 N_A_562_119#_M1020_g N_VPWR_c_1300_n 0.00136252f $X=5.395 $Y=2.315 $X2=0
+ $Y2=0
cc_596 N_A_562_119#_c_730_n N_VPWR_c_1314_n 0.00406468f $X=3.16 $Y=2.525 $X2=0
+ $Y2=0
cc_597 N_A_562_119#_M1016_g N_VPWR_c_1295_n 9.39239e-19 $X=4.28 $Y=2.525 $X2=0
+ $Y2=0
cc_598 N_A_562_119#_M1020_g N_VPWR_c_1295_n 7.82699e-19 $X=5.395 $Y=2.315 $X2=0
+ $Y2=0
cc_599 N_A_562_119#_c_730_n N_VPWR_c_1295_n 0.00684884f $X=3.16 $Y=2.525 $X2=0
+ $Y2=0
cc_600 N_A_562_119#_c_722_n N_A_476_119#_c_1458_n 0.00381069f $X=3.215 $Y=1.555
+ $X2=0 $Y2=0
cc_601 N_A_562_119#_c_730_n N_A_476_119#_c_1461_n 0.00151307f $X=3.16 $Y=2.525
+ $X2=0 $Y2=0
cc_602 N_A_562_119#_c_731_n N_A_476_119#_c_1461_n 0.0118063f $X=3.167 $Y=2.295
+ $X2=0 $Y2=0
cc_603 N_A_562_119#_c_722_n N_A_476_119#_c_1459_n 0.0124531f $X=3.215 $Y=1.555
+ $X2=0 $Y2=0
cc_604 N_A_562_119#_c_724_n N_A_476_119#_c_1459_n 0.00777965f $X=3.215 $Y=0.75
+ $X2=0 $Y2=0
cc_605 N_A_562_119#_c_722_n N_A_476_119#_c_1460_n 0.0197032f $X=3.215 $Y=1.555
+ $X2=0 $Y2=0
cc_606 N_A_562_119#_c_731_n N_A_476_119#_c_1460_n 0.0251422f $X=3.167 $Y=2.295
+ $X2=0 $Y2=0
cc_607 N_A_562_119#_c_732_n N_A_476_119#_c_1460_n 0.0127427f $X=3.215 $Y=1.64
+ $X2=0 $Y2=0
cc_608 N_A_562_119#_M1020_g N_A_1094_379#_c_1506_n 0.0108426f $X=5.395 $Y=2.315
+ $X2=0 $Y2=0
cc_609 N_A_562_119#_c_724_n N_VGND_c_1623_n 2.76242e-19 $X=3.215 $Y=0.75 $X2=0
+ $Y2=0
cc_610 N_A_562_119#_c_724_n N_VGND_c_1624_n 0.00991306f $X=3.215 $Y=0.75 $X2=0
+ $Y2=0
cc_611 N_A_562_119#_M1007_g N_VGND_c_1625_n 0.0040953f $X=4.495 $Y=0.445 $X2=0
+ $Y2=0
cc_612 N_A_562_119#_c_724_n N_VGND_c_1625_n 0.0127203f $X=3.215 $Y=0.75 $X2=0
+ $Y2=0
cc_613 N_A_562_119#_M1007_g N_VGND_c_1636_n 0.00549943f $X=4.495 $Y=0.445 $X2=0
+ $Y2=0
cc_614 N_A_562_119#_c_720_n N_VGND_c_1637_n 0.00486043f $X=5.8 $Y=0.985 $X2=0
+ $Y2=0
cc_615 N_A_562_119#_M1007_g N_VGND_c_1642_n 0.00233777f $X=4.495 $Y=0.445 $X2=0
+ $Y2=0
cc_616 N_A_562_119#_c_719_n N_VGND_c_1642_n 0.0107259f $X=5.47 $Y=1.06 $X2=0
+ $Y2=0
cc_617 N_A_562_119#_c_720_n N_VGND_c_1642_n 0.0173038f $X=5.8 $Y=0.985 $X2=0
+ $Y2=0
cc_618 N_A_562_119#_M1007_g N_VGND_c_1645_n 0.0113244f $X=4.495 $Y=0.445 $X2=0
+ $Y2=0
cc_619 N_A_562_119#_c_720_n N_VGND_c_1645_n 0.00813827f $X=5.8 $Y=0.985 $X2=0
+ $Y2=0
cc_620 N_A_562_119#_c_724_n N_VGND_c_1645_n 0.0144659f $X=3.215 $Y=0.75 $X2=0
+ $Y2=0
cc_621 N_A_562_119#_c_722_n A_648_119# 0.00104803f $X=3.215 $Y=1.555 $X2=-0.19
+ $Y2=-0.245
cc_622 N_A_562_119#_c_724_n A_648_119# 0.00357461f $X=3.215 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_623 N_A_30_99#_M1021_g N_A_1398_65#_M1008_g 0.0751595f $X=6.705 $Y=0.665
+ $X2=0 $Y2=0
cc_624 N_A_30_99#_M1021_g N_A_1398_65#_c_990_n 0.00323922f $X=6.705 $Y=0.665
+ $X2=0 $Y2=0
cc_625 N_A_30_99#_c_867_n N_A_1398_65#_c_990_n 0.0206213f $X=6.87 $Y=1.85 $X2=0
+ $Y2=0
cc_626 N_A_30_99#_M1026_g N_A_1398_65#_c_997_n 0.0206213f $X=6.87 $Y=2.455 $X2=0
+ $Y2=0
cc_627 N_A_30_99#_M1021_g N_A_1247_47#_c_1088_n 0.0192635f $X=6.705 $Y=0.665
+ $X2=0 $Y2=0
cc_628 N_A_30_99#_M1021_g N_A_1247_47#_c_1089_n 0.00494803f $X=6.705 $Y=0.665
+ $X2=0 $Y2=0
cc_629 N_A_30_99#_M1026_g N_A_1247_47#_c_1099_n 0.0101652f $X=6.87 $Y=2.455
+ $X2=0 $Y2=0
cc_630 N_A_30_99#_M1026_g N_A_1247_47#_c_1102_n 3.07718e-19 $X=6.87 $Y=2.455
+ $X2=0 $Y2=0
cc_631 N_A_30_99#_c_867_n N_A_1247_47#_c_1102_n 0.00473964f $X=6.87 $Y=1.85
+ $X2=0 $Y2=0
cc_632 N_A_30_99#_M1021_g N_A_1247_47#_c_1093_n 0.00693431f $X=6.705 $Y=0.665
+ $X2=0 $Y2=0
cc_633 N_A_30_99#_c_867_n N_A_1247_47#_c_1093_n 4.68003e-19 $X=6.87 $Y=1.85
+ $X2=0 $Y2=0
cc_634 N_A_30_99#_c_870_n N_VPWR_M1005_d 0.00174317f $X=1 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_635 N_A_30_99#_M1025_g N_VPWR_c_1296_n 0.0103232f $X=1.075 $Y=2.645 $X2=0
+ $Y2=0
cc_636 N_A_30_99#_c_860_n N_VPWR_c_1296_n 0.00746875f $X=1.15 $Y=3.15 $X2=0
+ $Y2=0
cc_637 N_A_30_99#_c_869_n N_VPWR_c_1296_n 0.0129486f $X=0.41 $Y=2.47 $X2=0 $Y2=0
cc_638 N_A_30_99#_c_870_n N_VPWR_c_1296_n 0.0168841f $X=1 $Y=2.385 $X2=0 $Y2=0
cc_639 N_A_30_99#_c_859_n N_VPWR_c_1297_n 0.0256494f $X=3.3 $Y=3.15 $X2=0 $Y2=0
cc_640 N_A_30_99#_M1000_g N_VPWR_c_1298_n 0.00811041f $X=3.375 $Y=2.525 $X2=0
+ $Y2=0
cc_641 N_A_30_99#_c_862_n N_VPWR_c_1298_n 0.0259148f $X=6.795 $Y=3.15 $X2=0
+ $Y2=0
cc_642 N_A_30_99#_c_862_n N_VPWR_c_1299_n 0.0272691f $X=6.795 $Y=3.15 $X2=0
+ $Y2=0
cc_643 N_A_30_99#_c_862_n N_VPWR_c_1300_n 0.0221956f $X=6.795 $Y=3.15 $X2=0
+ $Y2=0
cc_644 N_A_30_99#_c_862_n N_VPWR_c_1307_n 0.0372577f $X=6.795 $Y=3.15 $X2=0
+ $Y2=0
cc_645 N_A_30_99#_c_860_n N_VPWR_c_1313_n 0.0343499f $X=1.15 $Y=3.15 $X2=0 $Y2=0
cc_646 N_A_30_99#_c_859_n N_VPWR_c_1314_n 0.0432246f $X=3.3 $Y=3.15 $X2=0 $Y2=0
cc_647 N_A_30_99#_c_869_n N_VPWR_c_1317_n 0.0154375f $X=0.41 $Y=2.47 $X2=0 $Y2=0
cc_648 N_A_30_99#_c_859_n N_VPWR_c_1295_n 0.0658176f $X=3.3 $Y=3.15 $X2=0 $Y2=0
cc_649 N_A_30_99#_c_860_n N_VPWR_c_1295_n 0.00380229f $X=1.15 $Y=3.15 $X2=0
+ $Y2=0
cc_650 N_A_30_99#_c_862_n N_VPWR_c_1295_n 0.0921811f $X=6.795 $Y=3.15 $X2=0
+ $Y2=0
cc_651 N_A_30_99#_c_866_n N_VPWR_c_1295_n 0.00926736f $X=3.375 $Y=3.15 $X2=0
+ $Y2=0
cc_652 N_A_30_99#_c_869_n N_VPWR_c_1295_n 0.0129967f $X=0.41 $Y=2.47 $X2=0 $Y2=0
cc_653 N_A_30_99#_c_870_n N_VPWR_c_1295_n 0.0114703f $X=1 $Y=2.385 $X2=0 $Y2=0
cc_654 N_A_30_99#_c_850_n N_A_476_119#_c_1458_n 0.00303985f $X=2.66 $Y=0.18
+ $X2=0 $Y2=0
cc_655 N_A_30_99#_M1002_g N_A_476_119#_c_1458_n 9.59553e-19 $X=2.735 $Y=0.805
+ $X2=0 $Y2=0
cc_656 N_A_30_99#_c_859_n N_A_476_119#_c_1461_n 0.00404078f $X=3.3 $Y=3.15 $X2=0
+ $Y2=0
cc_657 N_A_30_99#_M1002_g N_A_476_119#_c_1459_n 0.00962072f $X=2.735 $Y=0.805
+ $X2=0 $Y2=0
cc_658 N_A_30_99#_c_862_n N_A_1094_379#_c_1507_n 0.00771487f $X=6.795 $Y=3.15
+ $X2=0 $Y2=0
cc_659 N_A_30_99#_c_862_n N_A_1094_379#_c_1508_n 0.0199187f $X=6.795 $Y=3.15
+ $X2=0 $Y2=0
cc_660 N_A_30_99#_M1026_g N_A_1094_379#_c_1508_n 0.0139464f $X=6.87 $Y=2.455
+ $X2=0 $Y2=0
cc_661 N_A_30_99#_M1026_g N_A_1201_407#_c_1533_n 7.68964e-19 $X=6.87 $Y=2.455
+ $X2=0 $Y2=0
cc_662 N_A_30_99#_M1026_g N_A_1201_407#_c_1534_n 0.0136029f $X=6.87 $Y=2.455
+ $X2=0 $Y2=0
cc_663 N_A_30_99#_c_851_n N_VGND_c_1622_n 0.0150103f $X=1.36 $Y=0.18 $X2=0 $Y2=0
cc_664 N_A_30_99#_c_855_n N_VGND_c_1622_n 0.00546224f $X=1.165 $Y=1.66 $X2=0
+ $Y2=0
cc_665 N_A_30_99#_c_856_n N_VGND_c_1622_n 0.00103206f $X=1.165 $Y=1.66 $X2=0
+ $Y2=0
cc_666 N_A_30_99#_M1001_g N_VGND_c_1623_n 0.00647046f $X=1.285 $Y=0.705 $X2=0
+ $Y2=0
cc_667 N_A_30_99#_c_850_n N_VGND_c_1623_n 0.0208866f $X=2.66 $Y=0.18 $X2=0 $Y2=0
cc_668 N_A_30_99#_M1002_g N_VGND_c_1623_n 0.00594808f $X=2.735 $Y=0.805 $X2=0
+ $Y2=0
cc_669 N_A_30_99#_c_850_n N_VGND_c_1624_n 0.0188116f $X=2.66 $Y=0.18 $X2=0 $Y2=0
cc_670 N_A_30_99#_c_854_n N_VGND_c_1631_n 0.0045032f $X=0.275 $Y=0.705 $X2=0
+ $Y2=0
cc_671 N_A_30_99#_c_851_n N_VGND_c_1635_n 0.0230985f $X=1.36 $Y=0.18 $X2=0 $Y2=0
cc_672 N_A_30_99#_M1021_g N_VGND_c_1637_n 0.00301185f $X=6.705 $Y=0.665 $X2=0
+ $Y2=0
cc_673 N_A_30_99#_c_850_n N_VGND_c_1645_n 0.0462811f $X=2.66 $Y=0.18 $X2=0 $Y2=0
cc_674 N_A_30_99#_c_851_n N_VGND_c_1645_n 0.0113471f $X=1.36 $Y=0.18 $X2=0 $Y2=0
cc_675 N_A_30_99#_M1021_g N_VGND_c_1645_n 0.00262976f $X=6.705 $Y=0.665 $X2=0
+ $Y2=0
cc_676 N_A_30_99#_c_854_n N_VGND_c_1645_n 0.00610626f $X=0.275 $Y=0.705 $X2=0
+ $Y2=0
cc_677 N_A_1398_65#_c_991_n N_A_1247_47#_c_1079_n 2.30209e-19 $X=8.41 $Y=0.62
+ $X2=0 $Y2=0
cc_678 N_A_1398_65#_c_993_n N_A_1247_47#_c_1079_n 0.00113006f $X=8.575 $Y=0.35
+ $X2=0 $Y2=0
cc_679 N_A_1398_65#_c_992_n N_A_1247_47#_c_1080_n 0.0134287f $X=9.435 $Y=0.35
+ $X2=0 $Y2=0
cc_680 N_A_1398_65#_c_993_n N_A_1247_47#_c_1080_n 0.00956474f $X=8.575 $Y=0.35
+ $X2=0 $Y2=0
cc_681 N_A_1398_65#_c_994_n N_A_1247_47#_c_1095_n 0.00687566f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_682 N_A_1398_65#_c_994_n N_A_1247_47#_c_1083_n 0.0230587f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_683 N_A_1398_65#_c_994_n N_A_1247_47#_M1011_g 0.00144861f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_684 N_A_1398_65#_c_1002_n N_A_1247_47#_M1011_g 0.0118029f $X=9.61 $Y=2.6
+ $X2=0 $Y2=0
cc_685 N_A_1398_65#_M1008_g N_A_1247_47#_c_1088_n 0.00348789f $X=7.065 $Y=0.665
+ $X2=0 $Y2=0
cc_686 N_A_1398_65#_c_989_n N_A_1247_47#_c_1099_n 0.00142837f $X=7.14 $Y=1.46
+ $X2=0 $Y2=0
cc_687 N_A_1398_65#_c_990_n N_A_1247_47#_c_1099_n 0.0139531f $X=7.455 $Y=3.075
+ $X2=0 $Y2=0
cc_688 N_A_1398_65#_M1014_g N_A_1247_47#_c_1099_n 0.00797958f $X=7.945 $Y=2.495
+ $X2=0 $Y2=0
cc_689 N_A_1398_65#_c_999_n N_A_1247_47#_c_1100_n 0.00628853f $X=9.445 $Y=3.15
+ $X2=0 $Y2=0
cc_690 N_A_1398_65#_c_994_n N_A_1247_47#_c_1090_n 0.0155636f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_691 N_A_1398_65#_c_994_n N_A_1247_47#_c_1091_n 0.0208002f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_692 N_A_1398_65#_c_991_n N_A_1247_47#_c_1147_n 0.00799771f $X=8.41 $Y=0.62
+ $X2=0 $Y2=0
cc_693 N_A_1398_65#_c_992_n N_A_1247_47#_c_1147_n 0.0229117f $X=9.435 $Y=0.35
+ $X2=0 $Y2=0
cc_694 N_A_1398_65#_c_994_n N_A_1247_47#_c_1147_n 0.0277603f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_695 N_A_1398_65#_c_992_n N_A_1247_47#_c_1092_n 0.0115705f $X=9.435 $Y=0.35
+ $X2=0 $Y2=0
cc_696 N_A_1398_65#_c_994_n N_A_1247_47#_c_1092_n 0.0272848f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_697 N_A_1398_65#_M1008_g N_A_1247_47#_c_1093_n 0.0140154f $X=7.065 $Y=0.665
+ $X2=0 $Y2=0
cc_698 N_A_1398_65#_c_988_n N_A_1247_47#_c_1093_n 0.00144817f $X=7.38 $Y=1.46
+ $X2=0 $Y2=0
cc_699 N_A_1398_65#_c_991_n N_A_1247_47#_c_1093_n 0.0204732f $X=8.41 $Y=0.62
+ $X2=0 $Y2=0
cc_700 N_A_1398_65#_c_992_n N_A_1247_47#_c_1093_n 0.0128162f $X=9.435 $Y=0.35
+ $X2=0 $Y2=0
cc_701 N_A_1398_65#_c_991_n N_A_1247_47#_c_1094_n 0.00533039f $X=8.41 $Y=0.62
+ $X2=0 $Y2=0
cc_702 N_A_1398_65#_c_992_n N_A_1247_47#_c_1094_n 0.00711491f $X=9.435 $Y=0.35
+ $X2=0 $Y2=0
cc_703 N_A_1398_65#_c_994_n N_A_1247_47#_c_1094_n 0.00304395f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_704 N_A_1398_65#_c_992_n N_A_1989_49#_c_1204_n 0.0145199f $X=9.435 $Y=0.35
+ $X2=0 $Y2=0
cc_705 N_A_1398_65#_c_994_n N_A_1989_49#_c_1204_n 0.0799423f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_706 N_A_1398_65#_c_994_n N_A_1989_49#_c_1205_n 0.116805f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_707 N_A_1398_65#_c_1002_n N_A_1989_49#_c_1205_n 0.00529322f $X=9.61 $Y=2.6
+ $X2=0 $Y2=0
cc_708 N_A_1398_65#_c_994_n N_A_1989_49#_c_1207_n 0.0138591f $X=9.55 $Y=1.885
+ $X2=0 $Y2=0
cc_709 N_A_1398_65#_c_990_n N_VPWR_c_1301_n 0.00147924f $X=7.455 $Y=3.075 $X2=0
+ $Y2=0
cc_710 N_A_1398_65#_M1014_g N_VPWR_c_1301_n 0.0176784f $X=7.945 $Y=2.495 $X2=0
+ $Y2=0
cc_711 N_A_1398_65#_c_999_n N_VPWR_c_1301_n 0.0184416f $X=9.445 $Y=3.15 $X2=0
+ $Y2=0
cc_712 N_A_1398_65#_c_1000_n N_VPWR_c_1301_n 0.00450684f $X=7.945 $Y=3.15 $X2=0
+ $Y2=0
cc_713 N_A_1398_65#_c_999_n N_VPWR_c_1302_n 0.0218601f $X=9.445 $Y=3.15 $X2=0
+ $Y2=0
cc_714 N_A_1398_65#_c_994_n N_VPWR_c_1302_n 0.093335f $X=9.55 $Y=1.885 $X2=0
+ $Y2=0
cc_715 N_A_1398_65#_c_1002_n N_VPWR_c_1302_n 0.00452559f $X=9.61 $Y=2.6 $X2=0
+ $Y2=0
cc_716 N_A_1398_65#_c_997_n N_VPWR_c_1307_n 0.0186077f $X=7.53 $Y=3.15 $X2=0
+ $Y2=0
cc_717 N_A_1398_65#_c_999_n N_VPWR_c_1309_n 0.0204671f $X=9.445 $Y=3.15 $X2=0
+ $Y2=0
cc_718 N_A_1398_65#_c_999_n N_VPWR_c_1311_n 0.0143974f $X=9.445 $Y=3.15 $X2=0
+ $Y2=0
cc_719 N_A_1398_65#_c_994_n N_VPWR_c_1311_n 0.0230096f $X=9.55 $Y=1.885 $X2=0
+ $Y2=0
cc_720 N_A_1398_65#_c_996_n N_VPWR_c_1295_n 0.0108567f $X=7.87 $Y=3.15 $X2=0
+ $Y2=0
cc_721 N_A_1398_65#_c_997_n N_VPWR_c_1295_n 0.00557134f $X=7.53 $Y=3.15 $X2=0
+ $Y2=0
cc_722 N_A_1398_65#_c_999_n N_VPWR_c_1295_n 0.0439328f $X=9.445 $Y=3.15 $X2=0
+ $Y2=0
cc_723 N_A_1398_65#_c_1000_n N_VPWR_c_1295_n 0.00749832f $X=7.945 $Y=3.15 $X2=0
+ $Y2=0
cc_724 N_A_1398_65#_c_994_n N_VPWR_c_1295_n 0.0115598f $X=9.55 $Y=1.885 $X2=0
+ $Y2=0
cc_725 N_A_1398_65#_c_990_n N_A_1094_379#_c_1508_n 0.00374103f $X=7.455 $Y=3.075
+ $X2=0 $Y2=0
cc_726 N_A_1398_65#_c_990_n N_A_1201_407#_c_1534_n 0.0124185f $X=7.455 $Y=3.075
+ $X2=0 $Y2=0
cc_727 N_A_1398_65#_c_990_n N_A_1201_407#_c_1536_n 0.00517187f $X=7.455 $Y=3.075
+ $X2=0 $Y2=0
cc_728 N_A_1398_65#_c_996_n N_A_1201_407#_c_1536_n 0.00295489f $X=7.87 $Y=3.15
+ $X2=0 $Y2=0
cc_729 N_A_1398_65#_M1008_g N_VGND_c_1626_n 0.00228172f $X=7.065 $Y=0.665 $X2=0
+ $Y2=0
cc_730 N_A_1398_65#_c_991_n N_VGND_c_1626_n 0.0153564f $X=8.41 $Y=0.62 $X2=0
+ $Y2=0
cc_731 N_A_1398_65#_c_993_n N_VGND_c_1626_n 0.0146654f $X=8.575 $Y=0.35 $X2=0
+ $Y2=0
cc_732 N_A_1398_65#_c_992_n N_VGND_c_1633_n 0.073533f $X=9.435 $Y=0.35 $X2=0
+ $Y2=0
cc_733 N_A_1398_65#_c_993_n N_VGND_c_1633_n 0.0163156f $X=8.575 $Y=0.35 $X2=0
+ $Y2=0
cc_734 N_A_1398_65#_M1008_g N_VGND_c_1637_n 0.00517164f $X=7.065 $Y=0.665 $X2=0
+ $Y2=0
cc_735 N_A_1398_65#_M1008_g N_VGND_c_1645_n 0.00519032f $X=7.065 $Y=0.665 $X2=0
+ $Y2=0
cc_736 N_A_1398_65#_c_992_n N_VGND_c_1645_n 0.0429212f $X=9.435 $Y=0.35 $X2=0
+ $Y2=0
cc_737 N_A_1398_65#_c_993_n N_VGND_c_1645_n 0.00879198f $X=8.575 $Y=0.35 $X2=0
+ $Y2=0
cc_738 N_A_1247_47#_M1012_g N_A_1989_49#_M1010_g 0.0231319f $X=10.285 $Y=0.665
+ $X2=0 $Y2=0
cc_739 N_A_1247_47#_M1011_g N_A_1989_49#_M1004_g 0.0205849f $X=10.285 $Y=2.465
+ $X2=0 $Y2=0
cc_740 N_A_1247_47#_c_1083_n N_A_1989_49#_c_1204_n 0.00467621f $X=10.21 $Y=1.49
+ $X2=0 $Y2=0
cc_741 N_A_1247_47#_M1012_g N_A_1989_49#_c_1204_n 0.0145217f $X=10.285 $Y=0.665
+ $X2=0 $Y2=0
cc_742 N_A_1247_47#_M1011_g N_A_1989_49#_c_1205_n 0.0111166f $X=10.285 $Y=2.465
+ $X2=0 $Y2=0
cc_743 N_A_1247_47#_M1011_g N_A_1989_49#_c_1206_n 0.00788918f $X=10.285 $Y=2.465
+ $X2=0 $Y2=0
cc_744 N_A_1247_47#_c_1087_n N_A_1989_49#_c_1206_n 0.010183f $X=10.285 $Y=1.49
+ $X2=0 $Y2=0
cc_745 N_A_1247_47#_c_1083_n N_A_1989_49#_c_1207_n 0.00993236f $X=10.21 $Y=1.49
+ $X2=0 $Y2=0
cc_746 N_A_1247_47#_M1012_g N_A_1989_49#_c_1208_n 0.0170849f $X=10.285 $Y=0.665
+ $X2=0 $Y2=0
cc_747 N_A_1247_47#_c_1099_n N_VPWR_c_1301_n 0.0216087f $X=8.495 $Y=2.1 $X2=0
+ $Y2=0
cc_748 N_A_1247_47#_c_1095_n N_VPWR_c_1302_n 0.00750315f $X=9.335 $Y=1.565 $X2=0
+ $Y2=0
cc_749 N_A_1247_47#_c_1100_n N_VPWR_c_1302_n 0.0388996f $X=8.59 $Y=2.495 $X2=0
+ $Y2=0
cc_750 N_A_1247_47#_c_1090_n N_VPWR_c_1302_n 0.0225827f $X=8.745 $Y=2.015 $X2=0
+ $Y2=0
cc_751 N_A_1247_47#_c_1091_n N_VPWR_c_1302_n 0.00768298f $X=9.1 $Y=0.955 $X2=0
+ $Y2=0
cc_752 N_A_1247_47#_c_1092_n N_VPWR_c_1302_n 0.0051035f $X=9.1 $Y=0.7 $X2=0
+ $Y2=0
cc_753 N_A_1247_47#_c_1103_n N_VPWR_c_1302_n 0.0146699f $X=8.665 $Y=2.1 $X2=0
+ $Y2=0
cc_754 N_A_1247_47#_M1011_g N_VPWR_c_1303_n 0.00433507f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_755 N_A_1247_47#_c_1100_n N_VPWR_c_1309_n 0.00605007f $X=8.59 $Y=2.495 $X2=0
+ $Y2=0
cc_756 N_A_1247_47#_M1011_g N_VPWR_c_1311_n 0.00585385f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_757 N_A_1247_47#_M1011_g N_VPWR_c_1295_n 0.0109148f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_758 N_A_1247_47#_c_1100_n N_VPWR_c_1295_n 0.00866112f $X=8.59 $Y=2.495 $X2=0
+ $Y2=0
cc_759 N_A_1247_47#_c_1099_n N_A_1094_379#_M1026_d 0.00508562f $X=8.495 $Y=2.1
+ $X2=0 $Y2=0
cc_760 N_A_1247_47#_M1036_d N_A_1094_379#_c_1508_n 0.00226996f $X=6.42 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_A_1247_47#_c_1102_n N_A_1201_407#_c_1533_n 0.0154283f $X=6.657 $Y=2.1
+ $X2=0 $Y2=0
cc_762 N_A_1247_47#_M1036_d N_A_1201_407#_c_1534_n 0.00411732f $X=6.42 $Y=2.035
+ $X2=0 $Y2=0
cc_763 N_A_1247_47#_c_1099_n N_A_1201_407#_c_1534_n 0.0299986f $X=8.495 $Y=2.1
+ $X2=0 $Y2=0
cc_764 N_A_1247_47#_c_1102_n N_A_1201_407#_c_1534_n 0.0167153f $X=6.657 $Y=2.1
+ $X2=0 $Y2=0
cc_765 N_A_1247_47#_c_1099_n N_A_1201_407#_c_1536_n 0.0198172f $X=8.495 $Y=2.1
+ $X2=0 $Y2=0
cc_766 N_A_1247_47#_c_1079_n N_VGND_c_1626_n 0.00723629f $X=8.195 $Y=0.345 $X2=0
+ $Y2=0
cc_767 N_A_1247_47#_c_1081_n N_VGND_c_1626_n 0.00766183f $X=8.27 $Y=0.27 $X2=0
+ $Y2=0
cc_768 N_A_1247_47#_c_1093_n N_VGND_c_1626_n 0.0497227f $X=8.655 $Y=1.08 $X2=0
+ $Y2=0
cc_769 N_A_1247_47#_M1012_g N_VGND_c_1627_n 0.00389861f $X=10.285 $Y=0.665 $X2=0
+ $Y2=0
cc_770 N_A_1247_47#_c_1081_n N_VGND_c_1633_n 0.0196773f $X=8.27 $Y=0.27 $X2=0
+ $Y2=0
cc_771 N_A_1247_47#_M1012_g N_VGND_c_1633_n 0.00575161f $X=10.285 $Y=0.665 $X2=0
+ $Y2=0
cc_772 N_A_1247_47#_c_1088_n N_VGND_c_1637_n 0.032875f $X=6.375 $Y=0.39 $X2=0
+ $Y2=0
cc_773 N_A_1247_47#_c_1088_n N_VGND_c_1642_n 0.0224954f $X=6.375 $Y=0.39 $X2=0
+ $Y2=0
cc_774 N_A_1247_47#_M1018_d N_VGND_c_1645_n 0.00215158f $X=6.235 $Y=0.235 $X2=0
+ $Y2=0
cc_775 N_A_1247_47#_c_1080_n N_VGND_c_1645_n 0.0220606f $X=8.935 $Y=0.27 $X2=0
+ $Y2=0
cc_776 N_A_1247_47#_c_1081_n N_VGND_c_1645_n 0.00756907f $X=8.27 $Y=0.27 $X2=0
+ $Y2=0
cc_777 N_A_1247_47#_M1012_g N_VGND_c_1645_n 0.0118604f $X=10.285 $Y=0.665 $X2=0
+ $Y2=0
cc_778 N_A_1247_47#_c_1088_n N_VGND_c_1645_n 0.0189837f $X=6.375 $Y=0.39 $X2=0
+ $Y2=0
cc_779 N_A_1989_49#_M1004_g N_VPWR_c_1303_n 0.0028697f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_780 N_A_1989_49#_c_1205_n N_VPWR_c_1303_n 0.00312548f $X=10.07 $Y=1.98 $X2=0
+ $Y2=0
cc_781 N_A_1989_49#_c_1206_n N_VPWR_c_1303_n 0.0190366f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_782 N_A_1989_49#_M1004_g N_VPWR_c_1304_n 7.38561e-19 $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_783 N_A_1989_49#_M1017_g N_VPWR_c_1304_n 0.0141984f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_784 N_A_1989_49#_M1022_g N_VPWR_c_1304_n 0.0141179f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_785 N_A_1989_49#_M1033_g N_VPWR_c_1304_n 7.24342e-19 $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_786 N_A_1989_49#_M1022_g N_VPWR_c_1306_n 7.24342e-19 $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_787 N_A_1989_49#_M1033_g N_VPWR_c_1306_n 0.0151814f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_788 N_A_1989_49#_c_1205_n N_VPWR_c_1311_n 0.0163642f $X=10.07 $Y=1.98 $X2=0
+ $Y2=0
cc_789 N_A_1989_49#_M1004_g N_VPWR_c_1315_n 0.00585385f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_790 N_A_1989_49#_M1017_g N_VPWR_c_1315_n 0.00486043f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_791 N_A_1989_49#_M1022_g N_VPWR_c_1316_n 0.00486043f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_792 N_A_1989_49#_M1033_g N_VPWR_c_1316_n 0.00486043f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_793 N_A_1989_49#_M1011_s N_VPWR_c_1295_n 0.00231412f $X=9.945 $Y=1.835 $X2=0
+ $Y2=0
cc_794 N_A_1989_49#_M1004_g N_VPWR_c_1295_n 0.0105477f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_795 N_A_1989_49#_M1017_g N_VPWR_c_1295_n 0.00824727f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_796 N_A_1989_49#_M1022_g N_VPWR_c_1295_n 0.00824727f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_797 N_A_1989_49#_M1033_g N_VPWR_c_1295_n 0.00824727f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_798 N_A_1989_49#_c_1205_n N_VPWR_c_1295_n 0.0100304f $X=10.07 $Y=1.98 $X2=0
+ $Y2=0
cc_799 N_A_1989_49#_M1023_g N_Q_c_1562_n 0.0139142f $X=11.145 $Y=0.665 $X2=0
+ $Y2=0
cc_800 N_A_1989_49#_M1029_g N_Q_c_1562_n 0.01419f $X=11.575 $Y=0.665 $X2=0 $Y2=0
cc_801 N_A_1989_49#_c_1206_n N_Q_c_1562_n 0.0447065f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_802 N_A_1989_49#_c_1208_n N_Q_c_1562_n 0.00244902f $X=12.005 $Y=1.51 $X2=0
+ $Y2=0
cc_803 N_A_1989_49#_M1010_g N_Q_c_1563_n 0.00255478f $X=10.715 $Y=0.665 $X2=0
+ $Y2=0
cc_804 N_A_1989_49#_c_1204_n N_Q_c_1563_n 0.00496017f $X=10.07 $Y=0.42 $X2=0
+ $Y2=0
cc_805 N_A_1989_49#_c_1206_n N_Q_c_1563_n 0.017393f $X=11.81 $Y=1.51 $X2=0 $Y2=0
cc_806 N_A_1989_49#_c_1208_n N_Q_c_1563_n 0.00255521f $X=12.005 $Y=1.51 $X2=0
+ $Y2=0
cc_807 N_A_1989_49#_M1017_g N_Q_c_1568_n 0.0129531f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_808 N_A_1989_49#_M1022_g N_Q_c_1568_n 0.0130453f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_809 N_A_1989_49#_c_1206_n N_Q_c_1568_n 0.0467265f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_810 N_A_1989_49#_c_1208_n N_Q_c_1568_n 0.00246472f $X=12.005 $Y=1.51 $X2=0
+ $Y2=0
cc_811 N_A_1989_49#_M1004_g N_Q_c_1569_n 8.59182e-19 $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_812 N_A_1989_49#_c_1205_n N_Q_c_1569_n 0.00107121f $X=10.07 $Y=1.98 $X2=0
+ $Y2=0
cc_813 N_A_1989_49#_c_1206_n N_Q_c_1569_n 0.0181554f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_814 N_A_1989_49#_c_1208_n N_Q_c_1569_n 0.00256759f $X=12.005 $Y=1.51 $X2=0
+ $Y2=0
cc_815 N_A_1989_49#_M1030_g N_Q_c_1564_n 0.0167327f $X=12.005 $Y=0.665 $X2=0
+ $Y2=0
cc_816 N_A_1989_49#_c_1206_n N_Q_c_1564_n 0.00596141f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_817 N_A_1989_49#_M1033_g N_Q_c_1570_n 0.0156308f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_818 N_A_1989_49#_c_1206_n N_Q_c_1570_n 0.0062318f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_819 N_A_1989_49#_c_1206_n N_Q_c_1565_n 0.014687f $X=11.81 $Y=1.51 $X2=0 $Y2=0
cc_820 N_A_1989_49#_c_1208_n N_Q_c_1565_n 0.00255521f $X=12.005 $Y=1.51 $X2=0
+ $Y2=0
cc_821 N_A_1989_49#_c_1206_n N_Q_c_1571_n 0.0153308f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_822 N_A_1989_49#_c_1208_n N_Q_c_1571_n 0.00256759f $X=12.005 $Y=1.51 $X2=0
+ $Y2=0
cc_823 N_A_1989_49#_M1030_g Q 0.0204004f $X=12.005 $Y=0.665 $X2=0 $Y2=0
cc_824 N_A_1989_49#_c_1206_n Q 0.0137865f $X=11.81 $Y=1.51 $X2=0 $Y2=0
cc_825 N_A_1989_49#_M1010_g N_VGND_c_1627_n 0.00244279f $X=10.715 $Y=0.665 $X2=0
+ $Y2=0
cc_826 N_A_1989_49#_c_1204_n N_VGND_c_1627_n 0.00152267f $X=10.07 $Y=0.42 $X2=0
+ $Y2=0
cc_827 N_A_1989_49#_c_1206_n N_VGND_c_1627_n 0.0140185f $X=11.81 $Y=1.51 $X2=0
+ $Y2=0
cc_828 N_A_1989_49#_M1010_g N_VGND_c_1628_n 6.29009e-19 $X=10.715 $Y=0.665 $X2=0
+ $Y2=0
cc_829 N_A_1989_49#_M1023_g N_VGND_c_1628_n 0.0113159f $X=11.145 $Y=0.665 $X2=0
+ $Y2=0
cc_830 N_A_1989_49#_M1029_g N_VGND_c_1628_n 0.0112407f $X=11.575 $Y=0.665 $X2=0
+ $Y2=0
cc_831 N_A_1989_49#_M1030_g N_VGND_c_1628_n 6.15775e-19 $X=12.005 $Y=0.665 $X2=0
+ $Y2=0
cc_832 N_A_1989_49#_M1029_g N_VGND_c_1630_n 6.15775e-19 $X=11.575 $Y=0.665 $X2=0
+ $Y2=0
cc_833 N_A_1989_49#_M1030_g N_VGND_c_1630_n 0.0126339f $X=12.005 $Y=0.665 $X2=0
+ $Y2=0
cc_834 N_A_1989_49#_c_1204_n N_VGND_c_1633_n 0.0161868f $X=10.07 $Y=0.42 $X2=0
+ $Y2=0
cc_835 N_A_1989_49#_M1010_g N_VGND_c_1638_n 0.00575161f $X=10.715 $Y=0.665 $X2=0
+ $Y2=0
cc_836 N_A_1989_49#_M1023_g N_VGND_c_1638_n 0.00477554f $X=11.145 $Y=0.665 $X2=0
+ $Y2=0
cc_837 N_A_1989_49#_M1029_g N_VGND_c_1639_n 0.00477554f $X=11.575 $Y=0.665 $X2=0
+ $Y2=0
cc_838 N_A_1989_49#_M1030_g N_VGND_c_1639_n 0.00477554f $X=12.005 $Y=0.665 $X2=0
+ $Y2=0
cc_839 N_A_1989_49#_M1012_s N_VGND_c_1645_n 0.00246284f $X=9.945 $Y=0.245 $X2=0
+ $Y2=0
cc_840 N_A_1989_49#_M1010_g N_VGND_c_1645_n 0.0105607f $X=10.715 $Y=0.665 $X2=0
+ $Y2=0
cc_841 N_A_1989_49#_M1023_g N_VGND_c_1645_n 0.00825815f $X=11.145 $Y=0.665 $X2=0
+ $Y2=0
cc_842 N_A_1989_49#_M1029_g N_VGND_c_1645_n 0.00825815f $X=11.575 $Y=0.665 $X2=0
+ $Y2=0
cc_843 N_A_1989_49#_M1030_g N_VGND_c_1645_n 0.00825815f $X=12.005 $Y=0.665 $X2=0
+ $Y2=0
cc_844 N_A_1989_49#_c_1204_n N_VGND_c_1645_n 0.00983606f $X=10.07 $Y=0.42 $X2=0
+ $Y2=0
cc_845 N_VPWR_c_1314_n N_A_476_119#_c_1461_n 0.00376384f $X=3.805 $Y=3.33 $X2=0
+ $Y2=0
cc_846 N_VPWR_c_1295_n N_A_476_119#_c_1461_n 0.00599747f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_847 N_VPWR_c_1295_n N_A_1094_379#_M1026_d 0.00206351f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_848 N_VPWR_c_1300_n N_A_1094_379#_c_1506_n 0.0336563f $X=5.18 $Y=2.27 $X2=0
+ $Y2=0
cc_849 N_VPWR_c_1300_n N_A_1094_379#_c_1507_n 0.0173959f $X=5.18 $Y=2.27 $X2=0
+ $Y2=0
cc_850 N_VPWR_c_1307_n N_A_1094_379#_c_1507_n 0.0222408f $X=7.995 $Y=3.33 $X2=0
+ $Y2=0
cc_851 N_VPWR_c_1295_n N_A_1094_379#_c_1507_n 0.0114525f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_852 N_VPWR_c_1301_n N_A_1094_379#_c_1508_n 0.00597165f $X=8.16 $Y=2.495 $X2=0
+ $Y2=0
cc_853 N_VPWR_c_1307_n N_A_1094_379#_c_1508_n 0.0955147f $X=7.995 $Y=3.33 $X2=0
+ $Y2=0
cc_854 N_VPWR_c_1295_n N_A_1094_379#_c_1508_n 0.0540983f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_855 N_VPWR_c_1307_n N_A_1201_407#_c_1534_n 0.00372597f $X=7.995 $Y=3.33 $X2=0
+ $Y2=0
cc_856 N_VPWR_c_1295_n N_A_1201_407#_c_1534_n 0.0073838f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_857 N_VPWR_c_1307_n N_A_1201_407#_c_1536_n 0.00467279f $X=7.995 $Y=3.33 $X2=0
+ $Y2=0
cc_858 N_VPWR_c_1295_n N_A_1201_407#_c_1536_n 0.00657532f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_859 N_VPWR_c_1295_n N_Q_M1004_d 0.0041489f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_860 N_VPWR_c_1295_n N_Q_M1022_d 0.00536646f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_861 N_VPWR_c_1315_n N_Q_c_1601_n 0.0136943f $X=11.195 $Y=3.33 $X2=0 $Y2=0
cc_862 N_VPWR_c_1295_n N_Q_c_1601_n 0.00866972f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_863 N_VPWR_M1017_s N_Q_c_1568_n 0.00176461f $X=11.22 $Y=1.835 $X2=0 $Y2=0
cc_864 N_VPWR_c_1304_n N_Q_c_1568_n 0.0170777f $X=11.36 $Y=2.19 $X2=0 $Y2=0
cc_865 N_VPWR_c_1303_n N_Q_c_1569_n 0.00338509f $X=10.5 $Y=1.96 $X2=0 $Y2=0
cc_866 N_VPWR_c_1316_n N_Q_c_1606_n 0.0124525f $X=12.055 $Y=3.33 $X2=0 $Y2=0
cc_867 N_VPWR_c_1295_n N_Q_c_1606_n 0.00730901f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_868 N_VPWR_M1033_s N_Q_c_1570_n 0.00275814f $X=12.08 $Y=1.835 $X2=0 $Y2=0
cc_869 N_VPWR_c_1306_n N_Q_c_1570_n 0.024087f $X=12.22 $Y=2.19 $X2=0 $Y2=0
cc_870 N_A_476_119#_c_1458_n N_VGND_c_1624_n 0.00391143f $X=2.52 $Y=0.805 $X2=0
+ $Y2=0
cc_871 N_A_476_119#_c_1458_n N_VGND_c_1645_n 0.00650784f $X=2.52 $Y=0.805 $X2=0
+ $Y2=0
cc_872 N_A_1094_379#_c_1506_n N_A_1201_407#_c_1533_n 0.0323025f $X=5.61 $Y=2.25
+ $X2=0 $Y2=0
cc_873 N_A_1094_379#_M1026_d N_A_1201_407#_c_1534_n 0.00826751f $X=6.945
+ $Y=2.035 $X2=0 $Y2=0
cc_874 N_A_1094_379#_c_1508_n N_A_1201_407#_c_1534_n 0.0652754f $X=7.18 $Y=2.96
+ $X2=0 $Y2=0
cc_875 N_A_1094_379#_c_1506_n N_A_1201_407#_c_1535_n 0.0139001f $X=5.61 $Y=2.25
+ $X2=0 $Y2=0
cc_876 N_A_1094_379#_c_1508_n N_A_1201_407#_c_1535_n 0.0263122f $X=7.18 $Y=2.96
+ $X2=0 $Y2=0
cc_877 N_Q_c_1562_n N_VGND_M1023_d 0.00176461f $X=11.695 $Y=1.16 $X2=0 $Y2=0
cc_878 N_Q_c_1566_n N_VGND_M1030_d 0.0022603f $X=12.267 $Y=1.245 $X2=0 $Y2=0
cc_879 N_Q_c_1563_n N_VGND_c_1627_n 0.0016514f $X=11.025 $Y=1.16 $X2=0 $Y2=0
cc_880 N_Q_c_1562_n N_VGND_c_1628_n 0.0170777f $X=11.695 $Y=1.16 $X2=0 $Y2=0
cc_881 N_Q_c_1564_n N_VGND_c_1630_n 0.00240047f $X=12.145 $Y=1.16 $X2=0 $Y2=0
cc_882 N_Q_c_1566_n N_VGND_c_1630_n 0.0216866f $X=12.267 $Y=1.245 $X2=0 $Y2=0
cc_883 N_Q_c_1616_p N_VGND_c_1638_n 0.0136943f $X=10.93 $Y=0.42 $X2=0 $Y2=0
cc_884 N_Q_c_1617_p N_VGND_c_1639_n 0.0124525f $X=11.79 $Y=0.42 $X2=0 $Y2=0
cc_885 N_Q_M1010_s N_VGND_c_1645_n 0.0041489f $X=10.79 $Y=0.245 $X2=0 $Y2=0
cc_886 N_Q_M1029_s N_VGND_c_1645_n 0.00536646f $X=11.65 $Y=0.245 $X2=0 $Y2=0
cc_887 N_Q_c_1616_p N_VGND_c_1645_n 0.00866972f $X=10.93 $Y=0.42 $X2=0 $Y2=0
cc_888 N_Q_c_1617_p N_VGND_c_1645_n 0.00730901f $X=11.79 $Y=0.42 $X2=0 $Y2=0
cc_889 N_VGND_c_1645_n A_914_47# 0.00509892f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_890 N_VGND_c_1645_n A_1175_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
