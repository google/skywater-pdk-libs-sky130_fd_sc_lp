* File: sky130_fd_sc_lp__nand4bb_1.pxi.spice
* Created: Wed Sep  2 10:06:39 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4BB_1%B_N N_B_N_M1007_g N_B_N_M1006_g B_N B_N B_N B_N
+ B_N N_B_N_c_75_n PM_SKY130_FD_SC_LP__NAND4BB_1%B_N
x_PM_SKY130_FD_SC_LP__NAND4BB_1%D N_D_M1002_g N_D_M1011_g D D N_D_c_103_n
+ PM_SKY130_FD_SC_LP__NAND4BB_1%D
x_PM_SKY130_FD_SC_LP__NAND4BB_1%C N_C_M1003_g N_C_M1004_g C N_C_c_135_n
+ N_C_c_136_n N_C_c_137_n PM_SKY130_FD_SC_LP__NAND4BB_1%C
x_PM_SKY130_FD_SC_LP__NAND4BB_1%A_49_367# N_A_49_367#_M1006_s
+ N_A_49_367#_M1007_s N_A_49_367#_M1005_g N_A_49_367#_M1000_g
+ N_A_49_367#_c_173_n N_A_49_367#_c_183_n N_A_49_367#_c_174_n
+ N_A_49_367#_c_175_n N_A_49_367#_c_176_n N_A_49_367#_c_177_n
+ PM_SKY130_FD_SC_LP__NAND4BB_1%A_49_367#
x_PM_SKY130_FD_SC_LP__NAND4BB_1%A_552_21# N_A_552_21#_M1001_d
+ N_A_552_21#_M1010_d N_A_552_21#_M1009_g N_A_552_21#_M1008_g
+ N_A_552_21#_c_233_n N_A_552_21#_c_241_n N_A_552_21#_c_234_n
+ N_A_552_21#_c_235_n N_A_552_21#_c_236_n N_A_552_21#_c_237_n
+ N_A_552_21#_c_238_n PM_SKY130_FD_SC_LP__NAND4BB_1%A_552_21#
x_PM_SKY130_FD_SC_LP__NAND4BB_1%A_N N_A_N_M1010_g N_A_N_M1001_g N_A_N_c_287_n
+ N_A_N_c_288_n N_A_N_c_289_n A_N A_N N_A_N_c_291_n
+ PM_SKY130_FD_SC_LP__NAND4BB_1%A_N
x_PM_SKY130_FD_SC_LP__NAND4BB_1%VPWR N_VPWR_M1007_d N_VPWR_M1004_d
+ N_VPWR_M1008_d N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n VPWR
+ N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_323_n
+ N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n
+ PM_SKY130_FD_SC_LP__NAND4BB_1%VPWR
x_PM_SKY130_FD_SC_LP__NAND4BB_1%Y N_Y_M1009_d N_Y_M1011_d N_Y_M1000_d
+ N_Y_c_376_n N_Y_c_370_n N_Y_c_371_n N_Y_c_383_n N_Y_c_368_n N_Y_c_373_n Y Y
+ N_Y_c_369_n PM_SKY130_FD_SC_LP__NAND4BB_1%Y
x_PM_SKY130_FD_SC_LP__NAND4BB_1%VGND N_VGND_M1006_d N_VGND_M1001_s
+ N_VGND_c_428_n N_VGND_c_429_n VGND N_VGND_c_430_n N_VGND_c_431_n
+ N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n
+ PM_SKY130_FD_SC_LP__NAND4BB_1%VGND
cc_1 VNB N_B_N_M1007_g 0.00685826f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_2 VNB N_B_N_M1006_g 0.024705f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_3 VNB B_N 0.00189554f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_B_N_c_75_n 0.0392273f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.375
cc_5 VNB N_D_M1002_g 0.0197187f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_6 VNB N_D_M1011_g 0.00661249f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_7 VNB D 0.00586103f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_D_c_103_n 0.0348252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_M1004_g 0.00810024f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.865
cc_10 VNB N_C_c_135_n 0.0280764f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_11 VNB N_C_c_136_n 0.00872992f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_12 VNB N_C_c_137_n 0.0169066f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_13 VNB N_A_49_367#_M1000_g 0.00793339f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_14 VNB N_A_49_367#_c_173_n 0.0323768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_49_367#_c_174_n 0.0153693f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.375
cc_16 VNB N_A_49_367#_c_175_n 0.00176067f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.375
cc_17 VNB N_A_49_367#_c_176_n 0.0340026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_49_367#_c_177_n 0.0180644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_552_21#_M1009_g 0.0292346f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A_552_21#_c_233_n 0.00643061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_552_21#_c_234_n 0.0450063f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.375
cc_22 VNB N_A_552_21#_c_235_n 0.00269553f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.375
cc_23 VNB N_A_552_21#_c_236_n 0.0337143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_552_21#_c_237_n 0.0128383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_552_21#_c_238_n 0.0142381f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.775
cc_26 VNB N_A_N_M1010_g 0.0110005f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_27 VNB N_A_N_c_287_n 0.0288562f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_A_N_c_288_n 0.0207414f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_29 VNB N_A_N_c_289_n 0.0231237f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_30 VNB A_N 0.00662401f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_31 VNB N_A_N_c_291_n 0.0184953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_323_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_368_n 0.00369944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_369_n 0.0131208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_428_n 0.0156316f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_36 VNB N_VGND_c_429_n 0.00942251f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_37 VNB N_VGND_c_430_n 0.0344426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_431_n 0.059125f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.375
cc_39 VNB N_VGND_c_432_n 0.0190901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_433_n 0.254892f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.405
cc_41 VNB N_VGND_c_434_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_435_n 0.00526527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_B_N_M1007_g 0.0290576f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.045
cc_44 VPB B_N 0.0312941f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_45 VPB N_D_M1011_g 0.0234684f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.865
cc_46 VPB D 0.00373963f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_47 VPB N_C_M1004_g 0.0204011f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.865
cc_48 VPB N_A_49_367#_M1000_g 0.0203946f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_49 VPB N_A_49_367#_c_173_n 0.0249336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_552_21#_M1008_g 0.0223198f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_51 VPB N_A_552_21#_c_233_n 0.00320746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_552_21#_c_241_n 0.0217732f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.375
cc_53 VPB N_A_552_21#_c_235_n 0.00282314f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.375
cc_54 VPB N_A_552_21#_c_236_n 0.0130195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_552_21#_c_237_n 0.0150972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_N_M1010_g 0.0303596f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.045
cc_57 VPB N_VPWR_c_324_n 0.0160694f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_58 VPB N_VPWR_c_325_n 0.00498127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_326_n 0.0392974f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.375
cc_60 VPB N_VPWR_c_327_n 0.0318701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_328_n 0.0155889f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.775
cc_62 VPB N_VPWR_c_329_n 0.0188793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_330_n 0.0290329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_323_n 0.105931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_332_n 0.00587781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_333_n 0.00631862f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_334_n 0.00929964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_Y_c_370_n 0.00516585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_Y_c_371_n 0.00347486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_Y_c_368_n 3.26324e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_Y_c_373_n 0.00486871f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.295
cc_72 N_B_N_M1006_g N_D_M1002_g 0.0169676f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_73 N_B_N_M1007_g N_D_M1011_g 0.00965338f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_74 B_N N_D_M1011_g 0.00473504f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_B_N_M1007_g D 7.08562e-19 $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_76 B_N D 0.0370116f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_B_N_c_75_n D 0.00223211f $X=0.81 $Y=1.375 $X2=0 $Y2=0
cc_78 B_N N_D_c_103_n 3.11554e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B_N_c_75_n N_D_c_103_n 0.0206138f $X=0.81 $Y=1.375 $X2=0 $Y2=0
cc_80 N_B_N_M1006_g N_A_49_367#_c_173_n 0.00485433f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_81 B_N N_A_49_367#_c_173_n 0.0742288f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B_N_c_75_n N_A_49_367#_c_173_n 0.0164641f $X=0.81 $Y=1.375 $X2=0 $Y2=0
cc_83 N_B_N_M1006_g N_A_49_367#_c_183_n 0.0139525f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_84 B_N N_A_49_367#_c_183_n 0.0114984f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_B_N_c_75_n N_A_49_367#_c_183_n 0.00499948f $X=0.81 $Y=1.375 $X2=0 $Y2=0
cc_86 B_N N_VPWR_M1007_d 0.0045141f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_87 N_B_N_M1007_g N_VPWR_c_324_n 0.00154655f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_88 B_N N_VPWR_c_324_n 0.0834399f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 B_N N_VPWR_c_327_n 0.00734884f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 B_N N_VPWR_c_323_n 0.00618612f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B_N_M1006_g N_VGND_c_428_n 0.00329746f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_92 N_B_N_M1006_g N_VGND_c_430_n 0.00399858f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_93 N_B_N_M1006_g N_VGND_c_433_n 0.0046122f $X=0.81 $Y=0.865 $X2=0 $Y2=0
cc_94 D N_C_M1004_g 8.74892e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_D_c_103_n N_C_M1004_g 0.0263314f $X=1.26 $Y=1.375 $X2=0 $Y2=0
cc_96 D N_C_c_135_n 2.31345e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_D_c_103_n N_C_c_135_n 0.0450231f $X=1.26 $Y=1.375 $X2=0 $Y2=0
cc_98 N_D_M1002_g N_C_c_136_n 0.00264675f $X=1.395 $Y=0.655 $X2=0 $Y2=0
cc_99 D N_C_c_136_n 0.0254367f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_D_M1002_g N_C_c_137_n 0.0450231f $X=1.395 $Y=0.655 $X2=0 $Y2=0
cc_101 N_D_M1002_g N_A_49_367#_c_183_n 0.0175985f $X=1.395 $Y=0.655 $X2=0 $Y2=0
cc_102 D N_A_49_367#_c_183_n 0.0235994f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_D_c_103_n N_A_49_367#_c_183_n 0.00145687f $X=1.26 $Y=1.375 $X2=0 $Y2=0
cc_104 N_D_M1011_g N_VPWR_c_324_n 0.0250788f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_105 D N_VPWR_c_324_n 0.0277917f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_D_c_103_n N_VPWR_c_324_n 9.85169e-19 $X=1.26 $Y=1.375 $X2=0 $Y2=0
cc_107 N_D_M1011_g N_VPWR_c_328_n 0.00486043f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_108 N_D_M1011_g N_VPWR_c_323_n 0.0082726f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_109 N_D_M1011_g N_Y_c_371_n 0.00319024f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_110 D N_Y_c_371_n 0.00506958f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_111 N_D_M1002_g N_VGND_c_428_n 0.0152376f $X=1.395 $Y=0.655 $X2=0 $Y2=0
cc_112 N_D_M1002_g N_VGND_c_431_n 0.00486043f $X=1.395 $Y=0.655 $X2=0 $Y2=0
cc_113 N_D_M1002_g N_VGND_c_433_n 0.00440948f $X=1.395 $Y=0.655 $X2=0 $Y2=0
cc_114 N_C_M1004_g N_A_49_367#_M1000_g 0.0377804f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_115 N_C_c_135_n N_A_49_367#_c_183_n 0.00427262f $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_116 N_C_c_136_n N_A_49_367#_c_183_n 0.0326226f $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_117 N_C_c_137_n N_A_49_367#_c_183_n 0.0136379f $X=1.845 $Y=1.185 $X2=0 $Y2=0
cc_118 N_C_c_135_n N_A_49_367#_c_175_n 5.08076e-19 $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_119 N_C_c_136_n N_A_49_367#_c_175_n 0.0205384f $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_120 N_C_c_137_n N_A_49_367#_c_175_n 8.93209e-19 $X=1.845 $Y=1.185 $X2=0 $Y2=0
cc_121 N_C_M1004_g N_A_49_367#_c_176_n 2.06149e-19 $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_122 N_C_c_136_n N_A_49_367#_c_176_n 0.00109322f $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_123 N_C_c_135_n N_A_49_367#_c_177_n 0.0207797f $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_124 N_C_c_137_n N_A_49_367#_c_177_n 0.0373865f $X=1.845 $Y=1.185 $X2=0 $Y2=0
cc_125 N_C_M1004_g N_VPWR_c_324_n 8.76878e-19 $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_126 N_C_M1004_g N_VPWR_c_325_n 0.00823616f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_127 N_C_M1004_g N_VPWR_c_328_n 0.0054895f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_128 N_C_M1004_g N_VPWR_c_323_n 0.0102827f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_129 N_C_M1004_g N_Y_c_376_n 0.015895f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_130 N_C_M1004_g N_Y_c_370_n 0.0118389f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_131 N_C_c_135_n N_Y_c_370_n 7.65356e-19 $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_132 N_C_c_136_n N_Y_c_370_n 0.017569f $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_133 N_C_M1004_g N_Y_c_371_n 0.00209483f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_134 N_C_c_135_n N_Y_c_371_n 5.40806e-19 $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_135 N_C_c_136_n N_Y_c_371_n 0.0227327f $X=1.845 $Y=1.35 $X2=0 $Y2=0
cc_136 N_C_M1004_g N_Y_c_383_n 9.76808e-19 $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_137 N_C_c_137_n N_VGND_c_428_n 0.00321301f $X=1.845 $Y=1.185 $X2=0 $Y2=0
cc_138 N_C_c_137_n N_VGND_c_431_n 0.00585385f $X=1.845 $Y=1.185 $X2=0 $Y2=0
cc_139 N_C_c_137_n N_VGND_c_433_n 0.00660378f $X=1.845 $Y=1.185 $X2=0 $Y2=0
cc_140 N_A_49_367#_c_183_n N_A_552_21#_M1009_g 7.01805e-19 $X=2.22 $Y=0.925
+ $X2=0 $Y2=0
cc_141 N_A_49_367#_c_175_n N_A_552_21#_M1009_g 7.5268e-19 $X=2.385 $Y=1.355
+ $X2=0 $Y2=0
cc_142 N_A_49_367#_c_176_n N_A_552_21#_M1009_g 0.0203967f $X=2.385 $Y=1.355
+ $X2=0 $Y2=0
cc_143 N_A_49_367#_c_177_n N_A_552_21#_M1009_g 0.0306166f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_144 N_A_49_367#_M1000_g N_A_552_21#_c_236_n 0.0267259f $X=2.405 $Y=2.465
+ $X2=0 $Y2=0
cc_145 N_A_49_367#_M1000_g N_VPWR_c_325_n 0.0096695f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_49_367#_M1000_g N_VPWR_c_329_n 0.0054895f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_49_367#_M1000_g N_VPWR_c_323_n 0.0102827f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_49_367#_M1000_g N_Y_c_376_n 9.81598e-19 $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_49_367#_M1000_g N_Y_c_370_n 0.0118338f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_49_367#_c_183_n N_Y_c_370_n 0.00513449f $X=2.22 $Y=0.925 $X2=0 $Y2=0
cc_151 N_A_49_367#_c_175_n N_Y_c_370_n 0.0182423f $X=2.385 $Y=1.355 $X2=0 $Y2=0
cc_152 N_A_49_367#_c_176_n N_Y_c_370_n 7.58131e-19 $X=2.385 $Y=1.355 $X2=0 $Y2=0
cc_153 N_A_49_367#_M1000_g N_Y_c_383_n 0.0163796f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_49_367#_M1000_g N_Y_c_368_n 0.00349481f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_49_367#_c_176_n N_Y_c_368_n 0.00200461f $X=2.385 $Y=1.355 $X2=0 $Y2=0
cc_156 N_A_49_367#_M1000_g N_Y_c_373_n 0.00242472f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_49_367#_c_175_n N_Y_c_373_n 0.00203611f $X=2.385 $Y=1.355 $X2=0 $Y2=0
cc_158 N_A_49_367#_c_176_n N_Y_c_373_n 0.00311089f $X=2.385 $Y=1.355 $X2=0 $Y2=0
cc_159 N_A_49_367#_c_183_n N_Y_c_369_n 0.0186722f $X=2.22 $Y=0.925 $X2=0 $Y2=0
cc_160 N_A_49_367#_c_175_n N_Y_c_369_n 0.0372169f $X=2.385 $Y=1.355 $X2=0 $Y2=0
cc_161 N_A_49_367#_c_177_n N_Y_c_369_n 0.0148378f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_162 N_A_49_367#_c_183_n N_VGND_M1006_d 0.0098952f $X=2.22 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_49_367#_c_183_n N_VGND_c_428_n 0.0217327f $X=2.22 $Y=0.925 $X2=0
+ $Y2=0
cc_164 N_A_49_367#_c_177_n N_VGND_c_431_n 0.00585385f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_165 N_A_49_367#_c_183_n N_VGND_c_433_n 0.0589428f $X=2.22 $Y=0.925 $X2=0
+ $Y2=0
cc_166 N_A_49_367#_c_174_n N_VGND_c_433_n 0.0104335f $X=0.465 $Y=0.925 $X2=0
+ $Y2=0
cc_167 N_A_49_367#_c_177_n N_VGND_c_433_n 0.00705731f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_168 N_A_49_367#_c_183_n A_294_47# 0.00297589f $X=2.22 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_49_367#_c_183_n A_366_47# 0.0101865f $X=2.22 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_49_367#_c_183_n A_474_47# 0.00312524f $X=2.22 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_49_367#_c_175_n A_474_47# 3.88982e-19 $X=2.385 $Y=1.355 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_552_21#_M1008_g N_A_N_M1010_g 0.0078072f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_552_21#_c_233_n N_A_N_M1010_g 0.016097f $X=3.645 $Y=1.645 $X2=0 $Y2=0
cc_174 N_A_552_21#_c_241_n N_A_N_M1010_g 0.00477255f $X=3.75 $Y=2.05 $X2=0 $Y2=0
cc_175 N_A_552_21#_c_234_n N_A_N_M1010_g 0.00263354f $X=4.12 $Y=1.56 $X2=0 $Y2=0
cc_176 N_A_552_21#_M1009_g N_A_N_c_288_n 5.63752e-19 $X=2.835 $Y=0.655 $X2=0
+ $Y2=0
cc_177 N_A_552_21#_c_233_n N_A_N_c_288_n 0.00711919f $X=3.645 $Y=1.645 $X2=0
+ $Y2=0
cc_178 N_A_552_21#_c_235_n N_A_N_c_288_n 0.00123573f $X=3.085 $Y=1.51 $X2=0
+ $Y2=0
cc_179 N_A_552_21#_c_236_n N_A_N_c_288_n 0.0219266f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_552_21#_c_234_n N_A_N_c_289_n 0.02126f $X=4.12 $Y=1.56 $X2=0 $Y2=0
cc_181 N_A_552_21#_M1009_g A_N 0.00236861f $X=2.835 $Y=0.655 $X2=0 $Y2=0
cc_182 N_A_552_21#_c_233_n A_N 0.0341586f $X=3.645 $Y=1.645 $X2=0 $Y2=0
cc_183 N_A_552_21#_c_234_n A_N 0.0450681f $X=4.12 $Y=1.56 $X2=0 $Y2=0
cc_184 N_A_552_21#_c_235_n A_N 0.00358393f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A_552_21#_c_236_n A_N 2.74493e-19 $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A_552_21#_M1009_g N_A_N_c_291_n 0.0048816f $X=2.835 $Y=0.655 $X2=0
+ $Y2=0
cc_187 N_A_552_21#_M1008_g N_VPWR_c_326_n 0.0129258f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_552_21#_c_233_n N_VPWR_c_326_n 0.0158309f $X=3.645 $Y=1.645 $X2=0
+ $Y2=0
cc_189 N_A_552_21#_c_235_n N_VPWR_c_326_n 0.0227268f $X=3.085 $Y=1.51 $X2=0
+ $Y2=0
cc_190 N_A_552_21#_c_236_n N_VPWR_c_326_n 0.00176416f $X=3.085 $Y=1.51 $X2=0
+ $Y2=0
cc_191 N_A_552_21#_M1008_g N_VPWR_c_329_n 0.00495816f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_A_552_21#_M1008_g N_VPWR_c_323_n 0.00988926f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A_552_21#_M1008_g N_Y_c_383_n 0.0184305f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_552_21#_M1009_g N_Y_c_368_n 0.00681985f $X=2.835 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_552_21#_M1008_g N_Y_c_368_n 2.5027e-19 $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_552_21#_c_235_n N_Y_c_368_n 0.0241645f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A_552_21#_c_236_n N_Y_c_368_n 0.00801317f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_198 N_A_552_21#_M1008_g N_Y_c_373_n 0.00566683f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A_552_21#_c_235_n N_Y_c_373_n 0.00329699f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A_552_21#_M1009_g N_Y_c_369_n 0.0292395f $X=2.835 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_552_21#_c_235_n N_Y_c_369_n 0.017323f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_202 N_A_552_21#_c_236_n N_Y_c_369_n 0.00531956f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_203 N_A_552_21#_M1009_g N_VGND_c_429_n 0.00284525f $X=2.835 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A_552_21#_M1009_g N_VGND_c_431_n 0.00357668f $X=2.835 $Y=0.655 $X2=0
+ $Y2=0
cc_205 N_A_552_21#_c_238_n N_VGND_c_432_n 0.0162405f $X=4.12 $Y=0.47 $X2=0 $Y2=0
cc_206 N_A_552_21#_M1009_g N_VGND_c_433_n 0.00693886f $X=2.835 $Y=0.655 $X2=0
+ $Y2=0
cc_207 N_A_552_21#_c_238_n N_VGND_c_433_n 0.0127937f $X=4.12 $Y=0.47 $X2=0 $Y2=0
cc_208 N_A_N_M1010_g N_VPWR_c_326_n 0.0134839f $X=3.535 $Y=2.045 $X2=0 $Y2=0
cc_209 N_A_N_M1010_g N_Y_c_383_n 2.36149e-19 $X=3.535 $Y=2.045 $X2=0 $Y2=0
cc_210 A_N N_Y_c_368_n 0.00702742f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_211 N_A_N_M1010_g N_Y_c_373_n 5.81082e-19 $X=3.535 $Y=2.045 $X2=0 $Y2=0
cc_212 N_A_N_c_289_n N_Y_c_369_n 0.00483889f $X=3.695 $Y=0.79 $X2=0 $Y2=0
cc_213 A_N N_Y_c_369_n 0.027159f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_214 N_A_N_c_291_n N_Y_c_369_n 0.00151229f $X=3.695 $Y=0.955 $X2=0 $Y2=0
cc_215 N_A_N_c_288_n N_VGND_c_429_n 2.04136e-19 $X=3.66 $Y=1.46 $X2=0 $Y2=0
cc_216 N_A_N_c_289_n N_VGND_c_429_n 0.00514396f $X=3.695 $Y=0.79 $X2=0 $Y2=0
cc_217 A_N N_VGND_c_429_n 0.0217184f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_218 N_A_N_c_291_n N_VGND_c_429_n 0.00438301f $X=3.695 $Y=0.955 $X2=0 $Y2=0
cc_219 N_A_N_c_289_n N_VGND_c_432_n 0.00560159f $X=3.695 $Y=0.79 $X2=0 $Y2=0
cc_220 N_A_N_c_289_n N_VGND_c_433_n 0.00794351f $X=3.695 $Y=0.79 $X2=0 $Y2=0
cc_221 A_N N_VGND_c_433_n 0.00637329f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_222 N_A_N_c_291_n N_VGND_c_433_n 4.16503e-19 $X=3.695 $Y=0.955 $X2=0 $Y2=0
cc_223 N_VPWR_c_323_n N_Y_M1011_d 0.00380103f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_c_323_n N_Y_M1000_d 0.00223559f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_225 N_VPWR_c_328_n N_Y_c_376_n 0.015688f $X=1.95 $Y=3.33 $X2=0 $Y2=0
cc_226 N_VPWR_c_323_n N_Y_c_376_n 0.00984745f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_227 N_VPWR_M1004_d N_Y_c_370_n 0.00345213f $X=1.9 $Y=1.835 $X2=0 $Y2=0
cc_228 N_VPWR_c_325_n N_Y_c_370_n 0.0257093f $X=2.115 $Y=2.115 $X2=0 $Y2=0
cc_229 N_VPWR_c_326_n N_Y_c_383_n 0.0946782f $X=3.31 $Y=2.065 $X2=0 $Y2=0
cc_230 N_VPWR_c_329_n N_Y_c_383_n 0.0213097f $X=2.99 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_323_n N_Y_c_383_n 0.0135865f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_232 N_Y_c_369_n N_VGND_c_429_n 0.0327064f $X=3.05 $Y=0.38 $X2=0 $Y2=0
cc_233 N_Y_c_369_n N_VGND_c_431_n 0.0378241f $X=3.05 $Y=0.38 $X2=0 $Y2=0
cc_234 N_Y_M1009_d N_VGND_c_433_n 0.00215158f $X=2.91 $Y=0.235 $X2=0 $Y2=0
cc_235 N_Y_c_369_n N_VGND_c_433_n 0.0224893f $X=3.05 $Y=0.38 $X2=0 $Y2=0
cc_236 N_Y_c_369_n A_474_47# 0.0111295f $X=3.05 $Y=0.38 $X2=-0.19 $Y2=-0.245
cc_237 N_VGND_c_433_n A_294_47# 0.00301881f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_238 N_VGND_c_433_n A_366_47# 0.00561644f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_239 N_VGND_c_433_n A_474_47# 0.00979005f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
