# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.000000 1.355000 2.425000 2.175000 ;
        RECT 2.000000 2.175000 2.550000 2.505000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.040000 0.470000 11.410000 2.225000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.940000 1.740000 12.395000 3.075000 ;
        RECT 12.125000 0.260000 12.395000 1.740000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.165000 1.945000 5.495000 2.245000 ;
        RECT 5.165000 2.245000 6.500000 2.490000 ;
        RECT 6.330000 2.490000 6.500000 2.845000 ;
        RECT 6.330000 2.845000 7.680000 3.075000 ;
        RECT 7.510000 1.715000 8.365000 2.045000 ;
        RECT 7.510000 2.045000 7.680000 2.845000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.470000 2.090000 ;
        RECT 0.085000 2.090000 0.430000 2.490000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 12.480000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 12.670000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.480000 0.085000 ;
      RECT  0.000000  3.245000 12.480000 3.415000 ;
      RECT  0.100000  0.085000  0.430000 1.040000 ;
      RECT  0.100000  2.660000  0.430000 3.245000 ;
      RECT  0.600000  2.260000  1.315000 2.930000 ;
      RECT  0.640000  0.830000  0.900000 1.285000 ;
      RECT  0.640000  1.285000  1.830000 1.455000 ;
      RECT  0.640000  1.455000  0.840000 2.260000 ;
      RECT  0.805000  0.265000  1.465000 0.515000 ;
      RECT  0.965000  2.930000  1.315000 3.075000 ;
      RECT  1.020000  1.815000  1.765000 2.090000 ;
      RECT  1.205000  0.515000  1.465000 0.945000 ;
      RECT  1.485000  2.090000  1.765000 2.975000 ;
      RECT  1.635000  1.015000  2.315000 1.185000 ;
      RECT  1.635000  1.185000  1.830000 1.285000 ;
      RECT  1.645000  0.085000  1.975000 0.845000 ;
      RECT  2.000000  2.675000  2.330000 3.245000 ;
      RECT  2.145000  0.300000  3.495000 0.470000 ;
      RECT  2.145000  0.470000  2.315000 1.015000 ;
      RECT  2.485000  0.645000  2.775000 0.975000 ;
      RECT  2.550000  2.720000  2.890000 3.050000 ;
      RECT  2.605000  0.975000  2.775000 1.765000 ;
      RECT  2.605000  1.765000  2.890000 1.935000 ;
      RECT  2.720000  1.935000  2.890000 2.720000 ;
      RECT  2.945000  0.645000  3.155000 1.415000 ;
      RECT  2.945000  1.415000  3.230000 1.585000 ;
      RECT  3.060000  1.585000  3.230000 2.485000 ;
      RECT  3.060000  2.485000  3.955000 2.655000 ;
      RECT  3.060000  2.655000  3.310000 3.050000 ;
      RECT  3.325000  0.470000  3.495000 1.075000 ;
      RECT  3.325000  1.075000  4.265000 1.235000 ;
      RECT  3.400000  1.235000  4.265000 1.245000 ;
      RECT  3.400000  1.245000  3.615000 2.165000 ;
      RECT  3.725000  0.085000  3.925000 0.905000 ;
      RECT  3.770000  2.825000  4.100000 3.245000 ;
      RECT  3.785000  1.765000  4.985000 1.935000 ;
      RECT  3.785000  1.935000  3.955000 2.485000 ;
      RECT  3.900000  1.415000  4.635000 1.585000 ;
      RECT  4.095000  0.605000  4.985000 0.775000 ;
      RECT  4.095000  0.775000  4.265000 1.075000 ;
      RECT  4.135000  2.175000  4.450000 2.505000 ;
      RECT  4.280000  2.505000  4.450000 2.685000 ;
      RECT  4.280000  2.685000  5.565000 3.015000 ;
      RECT  4.445000  0.955000  4.635000 1.415000 ;
      RECT  4.675000  1.935000  4.985000 2.505000 ;
      RECT  4.815000  0.775000  4.985000 1.245000 ;
      RECT  4.815000  1.245000  6.530000 1.335000 ;
      RECT  4.815000  1.335000  6.765000 1.415000 ;
      RECT  4.815000  1.595000  5.845000 1.685000 ;
      RECT  4.815000  1.685000  6.215000 1.765000 ;
      RECT  5.250000  0.085000  5.520000 1.075000 ;
      RECT  5.675000  1.765000  6.215000 2.015000 ;
      RECT  5.740000  0.265000  7.620000 0.445000 ;
      RECT  5.740000  0.445000  6.010000 1.075000 ;
      RECT  5.820000  2.660000  6.150000 3.245000 ;
      RECT  6.200000  0.615000  8.100000 0.785000 ;
      RECT  6.200000  0.785000  6.530000 1.075000 ;
      RECT  6.270000  1.415000  6.765000 1.505000 ;
      RECT  6.505000  1.505000  6.765000 2.005000 ;
      RECT  6.700000  0.955000  7.105000 1.165000 ;
      RECT  6.810000  2.285000  7.140000 2.675000 ;
      RECT  6.935000  1.165000  7.105000 1.315000 ;
      RECT  6.935000  1.315000  9.595000 1.325000 ;
      RECT  6.935000  1.325000 10.870000 1.485000 ;
      RECT  6.935000  1.485000  7.140000 2.285000 ;
      RECT  7.805000  0.955000  9.435000 1.145000 ;
      RECT  7.830000  0.400000  8.100000 0.615000 ;
      RECT  7.850000  2.280000  8.090000 3.245000 ;
      RECT  8.290000  2.225000  8.705000 2.555000 ;
      RECT  8.535000  1.485000  8.705000 2.225000 ;
      RECT  8.620000  0.085000  8.950000 0.730000 ;
      RECT  8.875000  2.200000  9.400000 2.530000 ;
      RECT  8.875000  2.530000  9.130000 3.065000 ;
      RECT  9.140000  0.640000  9.435000 0.955000 ;
      RECT  9.265000  1.485000 10.870000 1.495000 ;
      RECT  9.265000  1.495000  9.595000 1.985000 ;
      RECT  9.570000  2.155000  9.885000 3.245000 ;
      RECT  9.605000  0.085000  9.865000 0.970000 ;
      RECT 10.035000  0.640000 10.730000 1.155000 ;
      RECT 10.055000  1.985000 10.530000 2.155000 ;
      RECT 10.055000  2.155000 10.340000 2.805000 ;
      RECT 10.280000  1.665000 10.530000 1.985000 ;
      RECT 10.700000  1.495000 10.870000 2.395000 ;
      RECT 10.700000  2.395000 11.750000 2.565000 ;
      RECT 11.440000  2.735000 11.770000 3.245000 ;
      RECT 11.580000  0.085000 11.910000 1.060000 ;
      RECT 11.580000  1.230000 11.955000 1.560000 ;
      RECT 11.580000  1.560000 11.750000 2.395000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
  END
END sky130_fd_sc_lp__dfsbp_1
END LIBRARY
