* File: sky130_fd_sc_lp__nand2_1.pxi.spice
* Created: Wed Sep  2 10:02:36 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_1%B N_B_M1000_g N_B_M1003_g B B N_B_c_29_n
+ N_B_c_30_n PM_SKY130_FD_SC_LP__NAND2_1%B
x_PM_SKY130_FD_SC_LP__NAND2_1%A N_A_c_49_n N_A_M1002_g N_A_M1001_g A A
+ N_A_c_52_n PM_SKY130_FD_SC_LP__NAND2_1%A
x_PM_SKY130_FD_SC_LP__NAND2_1%VPWR N_VPWR_M1003_s N_VPWR_M1001_d N_VPWR_c_74_n
+ N_VPWR_c_75_n N_VPWR_c_76_n N_VPWR_c_77_n VPWR N_VPWR_c_78_n N_VPWR_c_73_n
+ PM_SKY130_FD_SC_LP__NAND2_1%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_1%Y N_Y_M1002_d N_Y_M1003_d Y Y Y Y Y Y Y N_Y_c_96_n
+ PM_SKY130_FD_SC_LP__NAND2_1%Y
x_PM_SKY130_FD_SC_LP__NAND2_1%VGND N_VGND_M1000_s N_VGND_c_112_n N_VGND_c_113_n
+ VGND N_VGND_c_114_n N_VGND_c_115_n PM_SKY130_FD_SC_LP__NAND2_1%VGND
cc_1 VNB N_B_M1003_g 0.00183793f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_2 VNB B 0.0203343f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_B_c_29_n 0.0434285f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_4 VNB N_B_c_30_n 0.020031f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.295
cc_5 VNB N_A_c_49_n 0.0209591f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.295
cc_6 VNB N_A_M1001_g 0.00183777f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_7 VNB A 0.0237775f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_c_52_n 0.0459604f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_9 VNB N_VPWR_c_73_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB Y 0.00433012f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_Y_c_96_n 0.0291598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_112_n 0.0115187f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.625
cc_13 VNB N_VGND_c_113_n 0.0358916f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_14 VNB N_VGND_c_114_n 0.028838f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.46
cc_15 VNB N_VGND_c_115_n 0.117362f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.46
cc_16 VPB N_B_M1003_g 0.0254723f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_17 VPB B 0.00719599f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_18 VPB N_A_M1001_g 0.0254689f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_19 VPB A 0.00880435f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_20 VPB N_VPWR_c_74_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_75_n 0.0483665f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_22 VPB N_VPWR_c_76_n 0.0116683f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.46
cc_23 VPB N_VPWR_c_77_n 0.0480342f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.295
cc_24 VPB N_VPWR_c_78_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.665
cc_25 VPB N_VPWR_c_73_n 0.0456597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB Y 0.0039378f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_27 N_B_c_30_n N_A_c_49_n 0.0307793f $X=0.362 $Y=1.295 $X2=-0.19 $Y2=-0.245
cc_28 N_B_M1003_g N_A_M1001_g 0.0131621f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_29 N_B_c_29_n N_A_c_52_n 0.0439414f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_30 N_B_M1003_g N_VPWR_c_75_n 0.0204427f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_31 B N_VPWR_c_75_n 0.026915f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_32 N_B_c_29_n N_VPWR_c_75_n 0.00129037f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_33 N_B_M1003_g N_VPWR_c_77_n 7.44844e-19 $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_34 N_B_M1003_g N_VPWR_c_78_n 0.00486043f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_35 N_B_M1003_g N_VPWR_c_73_n 0.0082726f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_36 B Y 0.0413494f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_37 N_B_c_30_n Y 0.0105708f $X=0.362 $Y=1.295 $X2=0 $Y2=0
cc_38 B N_VGND_c_113_n 0.0269149f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_39 N_B_c_29_n N_VGND_c_113_n 0.00141307f $X=0.33 $Y=1.46 $X2=0 $Y2=0
cc_40 N_B_c_30_n N_VGND_c_113_n 0.0144544f $X=0.362 $Y=1.295 $X2=0 $Y2=0
cc_41 N_B_c_30_n N_VGND_c_114_n 0.00400407f $X=0.362 $Y=1.295 $X2=0 $Y2=0
cc_42 N_B_c_30_n N_VGND_c_115_n 0.00772763f $X=0.362 $Y=1.295 $X2=0 $Y2=0
cc_43 N_A_M1001_g N_VPWR_c_75_n 7.84844e-19 $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_44 N_A_M1001_g N_VPWR_c_77_n 0.0162443f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_45 A N_VPWR_c_77_n 0.0252511f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_46 N_A_c_52_n N_VPWR_c_77_n 0.00129037f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_47 N_A_M1001_g N_VPWR_c_78_n 0.00564095f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_48 N_A_M1001_g N_VPWR_c_73_n 0.00950825f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_49 N_A_c_49_n Y 0.00957488f $X=0.875 $Y=1.295 $X2=0 $Y2=0
cc_50 A Y 0.0409759f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A_c_52_n Y 0.00909497f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_52 N_A_c_49_n N_Y_c_96_n 0.0239069f $X=0.875 $Y=1.295 $X2=0 $Y2=0
cc_53 A N_Y_c_96_n 0.0233313f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A_c_52_n N_Y_c_96_n 0.00152306f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_55 N_A_c_49_n N_VGND_c_113_n 0.00132793f $X=0.875 $Y=1.295 $X2=0 $Y2=0
cc_56 N_A_c_49_n N_VGND_c_114_n 0.00307037f $X=0.875 $Y=1.295 $X2=0 $Y2=0
cc_57 N_A_c_49_n N_VGND_c_115_n 0.00426815f $X=0.875 $Y=1.295 $X2=0 $Y2=0
cc_58 N_VPWR_c_73_n N_Y_M1003_d 0.00467071f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_59 N_VPWR_c_78_n Y 0.0131621f $X=0.985 $Y=3.33 $X2=0 $Y2=0
cc_60 N_VPWR_c_73_n Y 0.00808656f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_61 N_Y_c_96_n N_VGND_c_114_n 0.0243428f $X=1.09 $Y=0.525 $X2=0 $Y2=0
cc_62 N_Y_c_96_n N_VGND_c_115_n 0.0230493f $X=1.09 $Y=0.525 $X2=0 $Y2=0
cc_63 N_Y_c_96_n A_112_69# 0.00163585f $X=1.09 $Y=0.525 $X2=-0.19 $Y2=-0.245
