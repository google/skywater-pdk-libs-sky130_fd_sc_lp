* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VPWR A2 a_231_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_231_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_231_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Y a_119_500# a_231_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_119_500# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_119_500# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y a_119_500# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VGND A2 a_502_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 Y A1 a_502_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR B1_N a_119_500# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_502_65# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_502_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR A1 a_231_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_231_367# a_119_500# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
