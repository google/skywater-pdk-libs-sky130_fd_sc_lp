* File: sky130_fd_sc_lp__o21a_lp.spice
* Created: Fri Aug 28 11:04:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o21a_lp  VNB VPB A1 A2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_27_57#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_27_57#_M1003_d N_A2_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0756 PD=0.78 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_244_409#_M1005_d N_B1_M1005_g N_A_27_57#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_516_47# N_A_244_409#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_X_M1008_d N_A_244_409#_M1008_g A_516_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_146_409# N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1002 N_A_244_409#_M1002_d N_A2_M1002_g A_146_409# VPB PHIGHVT L=0.25 W=1
+ AD=0.29 AS=0.12 PD=1.58 PS=1.24 NRD=59.0803 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_A_244_409#_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.29 PD=1.28 PS=1.58 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_X_M1006_d N_A_244_409#_M1006_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX9_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o21a_lp.pxi.spice"
*
.ends
*
*
