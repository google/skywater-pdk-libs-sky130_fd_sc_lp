* File: sky130_fd_sc_lp__or3b_m.pex.spice
* Created: Wed Sep  2 10:31:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3B_M%C_N 2 5 9 13 15 18 20 21 22 23 24 31
r36 23 24 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r37 22 23 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r38 21 22 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r39 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r40 20 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r41 16 18 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.36 $Y=2.215
+ $X2=0.485 $Y2=2.215
r42 14 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r43 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r44 13 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.99
+ $X2=0.27 $Y2=1.005
r45 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.332 $Y=0.84
+ $X2=0.332 $Y2=0.99
r46 7 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.485 $Y=2.29
+ $X2=0.485 $Y2=2.215
r47 7 9 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=0.485 $Y=2.29
+ $X2=0.485 $Y2=2.885
r48 5 12 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.485 $Y=0.485
+ $X2=0.485 $Y2=0.84
r49 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.14 $X2=0.36
+ $Y2=2.215
r50 2 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.14 $X2=0.36
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_M%A_112_55# 1 2 8 9 10 11 15 17 19 21 24 27 29
+ 30 33 36
r58 33 36 48.5887 $w=2.08e-07 $l=9.2e-07 $layer=LI1_cond $X=0.7 $Y=2.82 $X2=0.7
+ $Y2=1.9
r59 29 35 7.28026 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=1.395
+ $X2=0.76 $Y2=1.23
r60 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.395 $X2=0.84 $Y2=1.395
r61 27 36 7.28026 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=1.735
+ $X2=0.76 $Y2=1.9
r62 27 29 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.76 $Y=1.735
+ $X2=0.76 $Y2=1.395
r63 24 35 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.7 $Y=0.55 $X2=0.7
+ $Y2=1.23
r64 20 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.84 $Y=1.38
+ $X2=0.84 $Y2=1.395
r65 20 21 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=0.84 $Y=1.38
+ $X2=0.84 $Y2=1.305
r66 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.46 $Y=0.77
+ $X2=1.46 $Y2=0.45
r67 13 15 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.42 $Y=1.38
+ $X2=1.42 $Y2=2.3
r68 12 21 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.305
+ $X2=0.84 $Y2=1.305
r69 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.345 $Y=1.305
+ $X2=1.42 $Y2=1.38
r70 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.345 $Y=1.305
+ $X2=1.005 $Y2=1.305
r71 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.385 $Y=0.845
+ $X2=1.46 $Y2=0.77
r72 9 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.385 $Y=0.845
+ $X2=1.005 $Y2=0.845
r73 8 21 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.93 $Y=1.23
+ $X2=0.84 $Y2=1.305
r74 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=0.92
+ $X2=1.005 $Y2=0.845
r75 7 8 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.93 $Y=0.92 $X2=0.93
+ $Y2=1.23
r76 2 33 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=2.675 $X2=0.7 $Y2=2.82
r77 1 24 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.275 $X2=0.7 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_M%B 3 7 11 12 13 14 18
c36 3 0 1.37734e-19 $X=1.78 $Y=2.3
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.87
+ $Y=1.325 $X2=1.87 $Y2=1.325
r38 14 19 8.90524 $w=4.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.815 $Y=1.665
+ $X2=1.815 $Y2=1.325
r39 13 19 0.785757 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=1.815 $Y=1.295
+ $X2=1.815 $Y2=1.325
r40 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.87 $Y=1.665
+ $X2=1.87 $Y2=1.325
r41 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.665
+ $X2=1.87 $Y2=1.83
r42 10 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.16
+ $X2=1.87 $Y2=1.325
r43 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.89 $Y=0.45 $X2=1.89
+ $Y2=1.16
r44 3 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.78 $Y=2.3 $X2=1.78
+ $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_M%A 3 6 7 8 9 14 15
r32 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=2.835
+ $X2=2.26 $Y2=2.67
r33 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=2.835 $X2=2.26 $Y2=2.835
r34 9 15 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=2.835 $X2=2.26
+ $Y2=2.835
r35 8 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.835 $X2=2.16
+ $Y2=2.835
r36 7 8 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.835 $X2=1.68
+ $Y2=2.835
r37 6 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.32 $Y=2.3 $X2=2.32
+ $Y2=2.67
r38 3 6 948.617 $w=1.5e-07 $l=1.85e-06 $layer=POLY_cond $X=2.32 $Y=0.45 $X2=2.32
+ $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_M%A_212_418# 1 2 3 12 15 18 19 20 22 23 24 27
+ 29 30 31 32 34 39 44 45
c85 44 0 3.14971e-19 $X=2.77 $Y=0.94
c86 22 0 1.37734e-19 $X=1.265 $Y=2.13
r87 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=0.94 $X2=2.77 $Y2=0.94
r88 39 41 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=0.515
+ $X2=1.245 $Y2=0.68
r89 34 45 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.66 $Y=1.93
+ $X2=2.66 $Y2=1.445
r90 32 45 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.715 $Y=1.305
+ $X2=2.715 $Y2=1.445
r91 31 43 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.945
+ $X2=2.715 $Y2=0.86
r92 31 32 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.715 $Y=0.945
+ $X2=2.715 $Y2=1.305
r93 29 43 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.575 $Y=0.86
+ $X2=2.715 $Y2=0.86
r94 29 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.575 $Y=0.86
+ $X2=2.21 $Y2=0.86
r95 25 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.105 $Y=0.775
+ $X2=2.21 $Y2=0.86
r96 25 27 12.6753 $w=2.08e-07 $l=2.4e-07 $layer=LI1_cond $X=2.105 $Y=0.775
+ $X2=2.105 $Y2=0.535
r97 23 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=2.015
+ $X2=2.66 $Y2=1.93
r98 23 24 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.575 $Y=2.015
+ $X2=1.7 $Y2=2.015
r99 22 24 21.8725 $w=2.6e-07 $l=4.9135e-07 $layer=LI1_cond $X=1.265 $Y=2.135
+ $X2=1.7 $Y2=2.015
r100 22 36 3.75385 $w=2.6e-07 $l=8e-08 $layer=LI1_cond $X=1.265 $Y=2.135
+ $X2=1.185 $Y2=2.135
r101 22 41 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=1.265 $Y=2.13
+ $X2=1.265 $Y2=0.68
r102 19 44 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.77 $Y=1.28
+ $X2=2.77 $Y2=0.94
r103 19 20 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.28
+ $X2=2.77 $Y2=1.445
r104 18 44 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=0.775
+ $X2=2.77 $Y2=0.94
r105 15 20 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.795 $Y=2.3
+ $X2=2.795 $Y2=1.445
r106 12 18 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.75 $Y=0.45
+ $X2=2.75 $Y2=0.775
r107 3 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=2.09 $X2=1.185 $Y2=2.235
r108 2 27 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.24 $X2=2.105 $Y2=0.535
r109 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.24 $X2=1.245 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_M%VPWR 1 2 7 9 12 16 19 20 21 31 32
r34 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 26 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 23 35 3.52085 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r42 23 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 21 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 19 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.53 $Y=3.33 $X2=2.16
+ $Y2=3.33
r46 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=3.33
+ $X2=2.615 $Y2=3.33
r47 18 31 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.7 $Y=3.33 $X2=3.12
+ $Y2=3.33
r48 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=3.33 $X2=2.615
+ $Y2=3.33
r49 14 16 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.535 $Y=2.385
+ $X2=2.615 $Y2=2.385
r50 12 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=3.33
r51 11 16 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.615 $Y=2.49
+ $X2=2.615 $Y2=2.385
r52 11 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.615 $Y=2.49
+ $X2=2.615 $Y2=3.245
r53 7 35 3.32305 $w=1.9e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.177 $Y2=3.33
r54 7 9 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r55 2 14 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=2.09 $X2=2.535 $Y2=2.385
r56 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.675 $X2=0.27 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_M%X 1 2 7 8 9 10 11 12 13 36 38
r18 36 38 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=3.065 $Y=2.365
+ $X2=3.065 $Y2=2.405
r19 34 36 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.065 $Y=2.34
+ $X2=3.065 $Y2=2.365
r20 12 34 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=3.065 $Y=2.33
+ $X2=3.065 $Y2=2.34
r21 12 50 7.11633 $w=2.78e-07 $l=1.3e-07 $layer=LI1_cond $X=3.065 $Y=2.33
+ $X2=3.065 $Y2=2.2
r22 12 13 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.065 $Y=2.415
+ $X2=3.065 $Y2=2.775
r23 12 38 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=3.065 $Y=2.415
+ $X2=3.065 $Y2=2.405
r24 11 50 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=2.035
+ $X2=3.12 $Y2=2.2
r25 10 11 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=2.035
r26 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.295 $X2=3.12
+ $Y2=1.665
r27 8 9 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=0.925 $X2=3.12
+ $Y2=1.295
r28 7 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=0.43 $X2=3.12
+ $Y2=0.595
r29 7 44 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.12 $Y=0.43
+ $X2=2.965 $Y2=0.43
r30 7 8 20.0941 $w=1.68e-07 $l=3.08e-07 $layer=LI1_cond $X=3.12 $Y=0.617
+ $X2=3.12 $Y2=0.925
r31 7 23 1.43529 $w=1.68e-07 $l=2.2e-08 $layer=LI1_cond $X=3.12 $Y=0.617
+ $X2=3.12 $Y2=0.595
r32 2 36 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=2.09 $X2=3.03 $Y2=2.365
r33 1 44 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.24 $X2=2.965 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_M%VGND 1 2 3 10 12 16 20 23 24 25 27 37 38 44
c50 38 0 1.32842e-19 $X=3.12 $Y=0
c51 20 0 1.82128e-19 $X=2.535 $Y=0.385
r52 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r55 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 32 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.675
+ $Y2=0
r57 32 34 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=2.16
+ $Y2=0
r58 31 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r59 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r60 28 41 3.65184 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=0.187
+ $Y2=0
r61 28 30 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=1.2
+ $Y2=0
r62 27 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.675
+ $Y2=0
r63 27 30 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.2
+ $Y2=0
r64 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r65 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r66 25 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 23 34 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.16
+ $Y2=0
r68 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.535
+ $Y2=0
r69 22 37 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r70 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.535
+ $Y2=0
r71 18 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0
r72 18 20 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0.385
r73 14 44 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0
r74 14 16 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0.385
r75 10 41 3.26335 $w=2.1e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.187 $Y2=0
r76 10 12 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.42
r77 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.24 $X2=2.535 $Y2=0.385
r78 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.24 $X2=1.675 $Y2=0.385
r79 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.275 $X2=0.27 $Y2=0.42
.ends

