* File: sky130_fd_sc_lp__nor4_1.spice
* Created: Fri Aug 28 10:57:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4_1.pex.spice"
.subckt sky130_fd_sc_lp__nor4_1  VNB VPB A B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001.7 A=0.126
+ P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.84 AD=0.21
+ AS=0.1176 PD=1.34 PS=1.12 NRD=15.708 NRS=0 M=1 R=5.6 SA=75000.6 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_C_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.21 PD=1.12 PS=1.34 NRD=0 NRS=15.708 M=1 R=5.6 SA=75001.3 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.7 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1007 A_110_367# N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26 AD=0.2079
+ AS=0.3339 PD=1.59 PS=3.05 NRD=17.1981 NRS=0 M=1 R=8.4 SA=75000.2 SB=75001.7
+ A=0.189 P=2.82 MULT=1
MM1003 A_206_367# N_B_M1003_g A_110_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2142
+ AS=0.2079 PD=1.6 PS=1.59 NRD=17.9664 NRS=17.1981 M=1 R=8.4 SA=75000.7
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1006 A_304_367# N_C_M1006_g A_206_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.2142 PD=1.65 PS=1.6 NRD=21.8867 NRS=17.9664 M=1 R=8.4 SA=75001.2
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_D_M1001_g A_304_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.3339
+ AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75001.7 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__nor4_1.pxi.spice"
*
.ends
*
*
