* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4_2 A B C D VGND VNB VPB VPWR Y
X0 Y A a_523_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND D a_69_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_69_47# C a_330_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_523_67# B a_330_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_330_47# B a_523_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_523_67# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_69_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_330_47# C a_69_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
