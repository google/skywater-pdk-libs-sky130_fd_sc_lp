* File: sky130_fd_sc_lp__nand4bb_1.pex.spice
* Created: Fri Aug 28 10:52:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%B_N 3 7 9 10 11 12 13 24
c28 9 0 4.42457e-20 $X=0.72 $Y=1.295
r29 22 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.72 $Y=1.375 $X2=0.81
+ $Y2=1.375
r30 19 22 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=0.605 $Y=1.375
+ $X2=0.72 $Y2=1.375
r31 12 13 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.72 $Y2=2.775
r32 11 12 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.405
r33 10 11 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=2.035
r34 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.295 $X2=0.72
+ $Y2=1.665
r35 9 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.375 $X2=0.72 $Y2=1.375
r36 5 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.81 $Y=1.21
+ $X2=0.81 $Y2=1.375
r37 5 7 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.81 $Y=1.21 $X2=0.81
+ $Y2=0.865
r38 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.54
+ $X2=0.605 $Y2=1.375
r39 1 3 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.605 $Y=1.54
+ $X2=0.605 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%D 3 7 9 10 14
c34 3 0 4.42457e-20 $X=1.395 $Y=0.655
r35 14 17 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.282 $Y=1.375
+ $X2=1.282 $Y2=1.54
r36 14 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.282 $Y=1.375
+ $X2=1.282 $Y2=1.21
r37 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.295
+ $X2=1.175 $Y2=1.665
r38 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=1.375 $X2=1.26 $Y2=1.375
r39 7 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.395 $Y=2.465
+ $X2=1.395 $Y2=1.54
r40 3 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.395 $Y=0.655
+ $X2=1.395 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%C 3 6 8 11 12 13
r38 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.35
+ $X2=1.845 $Y2=1.515
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.35
+ $X2=1.845 $Y2=1.185
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.35 $X2=1.845 $Y2=1.35
r41 8 12 5.94228 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.36
+ $X2=1.845 $Y2=1.36
r42 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.825 $Y=2.465
+ $X2=1.825 $Y2=1.515
r43 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.755 $Y=0.655
+ $X2=1.755 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%A_49_367# 1 2 9 12 16 18 19 24 25 28
r60 25 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.355
+ $X2=2.385 $Y2=1.52
r61 25 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.355
+ $X2=2.385 $Y2=1.19
r62 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.355 $X2=2.385 $Y2=1.355
r63 22 24 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=2.35 $Y=1.03
+ $X2=2.35 $Y2=1.355
r64 19 21 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=0.465 $Y=0.925
+ $X2=0.575 $Y2=0.925
r65 18 22 6.91731 $w=2.1e-07 $l=1.74786e-07 $layer=LI1_cond $X=2.22 $Y=0.925
+ $X2=2.35 $Y2=1.03
r66 18 21 86.8788 $w=2.08e-07 $l=1.645e-06 $layer=LI1_cond $X=2.22 $Y=0.925
+ $X2=0.575 $Y2=0.925
r67 14 19 6.91731 $w=2.1e-07 $l=1.74786e-07 $layer=LI1_cond $X=0.335 $Y=1.03
+ $X2=0.465 $Y2=0.925
r68 14 16 44.9896 $w=2.58e-07 $l=1.015e-06 $layer=LI1_cond $X=0.335 $Y=1.03
+ $X2=0.335 $Y2=2.045
r69 12 29 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=2.405 $Y=2.465
+ $X2=2.405 $Y2=1.52
r70 9 28 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.295 $Y=0.655
+ $X2=2.295 $Y2=1.19
r71 2 16 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.045
r72 1 21 182 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_NDIFF $count=1 $X=0.45
+ $Y=0.655 $X2=0.575 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%A_552_21# 1 2 9 13 15 19 22 24 25 30 35
c54 24 0 1.54797e-19 $X=3.085 $Y=1.51
r55 33 35 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4 $Y=0.47 $X2=4.12
+ $Y2=0.47
r56 25 37 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.085 $Y=1.51
+ $X2=2.835 $Y2=1.51
r57 24 27 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=3.12 $Y=1.51
+ $X2=3.12 $Y2=1.645
r58 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.085
+ $Y=1.51 $X2=3.085 $Y2=1.51
r59 22 30 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=1.56
+ $X2=4.12 $Y2=1.645
r60 21 35 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=0.635
+ $X2=4.12 $Y2=0.47
r61 21 22 56.9949 $w=1.78e-07 $l=9.25e-07 $layer=LI1_cond $X=4.12 $Y=0.635
+ $X2=4.12 $Y2=1.56
r62 17 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.78 $Y=1.645
+ $X2=4.12 $Y2=1.645
r63 17 19 13.6586 $w=2.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.78 $Y=1.73
+ $X2=3.78 $Y2=2.05
r64 16 27 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.25 $Y=1.645
+ $X2=3.12 $Y2=1.645
r65 15 17 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.645 $Y=1.645
+ $X2=3.78 $Y2=1.645
r66 15 16 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.645 $Y=1.645
+ $X2=3.25 $Y2=1.645
r67 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.675
+ $X2=2.835 $Y2=1.51
r68 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.835 $Y=1.675
+ $X2=2.835 $Y2=2.465
r69 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.345
+ $X2=2.835 $Y2=1.51
r70 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.835 $Y=1.345
+ $X2=2.835 $Y2=0.655
r71 2 19 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=1.835 $X2=3.75 $Y2=2.05
r72 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.86
+ $Y=0.26 $X2=4 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%A_N 3 7 9 10 12 13 14 18
c37 10 0 4.08416e-20 $X=3.66 $Y=1.46
c38 3 0 1.54797e-19 $X=3.535 $Y=2.045
r39 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.695
+ $Y=0.955 $X2=3.695 $Y2=0.955
r40 14 19 8.90524 $w=4.38e-07 $l=3.4e-07 $layer=LI1_cond $X=3.64 $Y=1.295
+ $X2=3.64 $Y2=0.955
r41 13 19 0.785757 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=3.64 $Y=0.925
+ $X2=3.64 $Y2=0.955
r42 12 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=0.79
+ $X2=3.695 $Y2=0.955
r43 9 18 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.695 $Y=1.31
+ $X2=3.695 $Y2=0.955
r44 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.66 $Y=1.31 $X2=3.66
+ $Y2=1.46
r45 7 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.785 $Y=0.47
+ $X2=3.785 $Y2=0.79
r46 3 10 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=3.535 $Y=2.045
+ $X2=3.535 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%VPWR 1 2 3 12 18 24 28 30 35 40 47 48 51
+ 54 57
r45 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 48 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 45 57 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=3.475 $Y=3.33
+ $X2=3.232 $Y2=3.33
r50 45 47 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.475 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 44 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 41 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.115 $Y2=3.33
r54 41 43 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 40 57 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=3.232 $Y2=3.33
r56 40 43 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 36 51 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.16 $Y2=3.33
r60 36 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=3.33
+ $X2=2.115 $Y2=3.33
r62 35 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.95 $Y=3.33 $X2=1.68
+ $Y2=3.33
r63 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 30 51 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.16 $Y2=3.33
r66 30 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 28 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 24 27 10.3578 $w=4.83e-07 $l=4.2e-07 $layer=LI1_cond $X=3.232 $Y=2.065
+ $X2=3.232 $Y2=2.485
r71 22 57 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.232 $Y=3.245
+ $X2=3.232 $Y2=3.33
r72 22 27 18.7427 $w=4.83e-07 $l=7.6e-07 $layer=LI1_cond $X=3.232 $Y=3.245
+ $X2=3.232 $Y2=2.485
r73 18 21 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.115 $Y=2.115
+ $X2=2.115 $Y2=2.95
r74 16 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=3.245
+ $X2=2.115 $Y2=3.33
r75 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.115 $Y=3.245
+ $X2=2.115 $Y2=2.95
r76 12 15 13.2375 $w=3.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.16 $Y=2.085
+ $X2=1.16 $Y2=2.51
r77 10 51 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=3.245
+ $X2=1.16 $Y2=3.33
r78 10 15 22.8931 $w=3.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.16 $Y=3.245
+ $X2=1.16 $Y2=2.51
r79 3 27 300 $w=1.7e-07 $l=7.27839e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=1.835 $X2=3.075 $Y2=2.485
r80 3 24 600 $w=1.7e-07 $l=5.01996e-07 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=1.835 $X2=3.31 $Y2=2.065
r81 2 21 400 $w=1.7e-07 $l=1.21776e-06 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.835 $X2=2.115 $Y2=2.95
r82 2 18 400 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.835 $X2=2.115 $Y2=2.115
r83 1 15 300 $w=1.7e-07 $l=8.90576e-07 $layer=licon1_PDIFF $count=2 $X=0.68
+ $Y=1.835 $X2=1.18 $Y2=2.51
r84 1 12 600 $w=1.7e-07 $l=5.09902e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.835 $X2=1.08 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%Y 1 2 3 12 16 17 20 25 26 27 28 32
c60 25 0 4.08416e-20 $X=2.735 $Y=1.69
r61 28 38 10.5548 $w=5.98e-07 $l=1.85e-07 $layer=LI1_cond $X=2.95 $Y=0.925
+ $X2=2.95 $Y2=1.11
r62 27 28 7.37582 $w=5.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.95 $Y=0.555
+ $X2=2.95 $Y2=0.925
r63 27 32 3.48856 $w=5.98e-07 $l=1.75e-07 $layer=LI1_cond $X=2.95 $Y=0.555
+ $X2=2.95 $Y2=0.38
r64 25 26 3.49088 $w=2.67e-07 $l=1.33918e-07 $layer=LI1_cond $X=2.735 $Y=1.69
+ $X2=2.637 $Y2=1.775
r65 25 38 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.735 $Y=1.69
+ $X2=2.735 $Y2=1.11
r66 20 22 29.3636 $w=3.63e-07 $l=9.3e-07 $layer=LI1_cond $X=2.637 $Y=1.98
+ $X2=2.637 $Y2=2.91
r67 18 26 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=2.637 $Y=1.86
+ $X2=2.637 $Y2=1.775
r68 18 20 3.78885 $w=3.63e-07 $l=1.2e-07 $layer=LI1_cond $X=2.637 $Y=1.86
+ $X2=2.637 $Y2=1.98
r69 16 26 3.01551 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.455 $Y=1.775
+ $X2=2.637 $Y2=1.775
r70 16 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.455 $Y=1.775
+ $X2=1.775 $Y2=1.775
r71 12 14 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=1.645 $Y=1.98
+ $X2=1.645 $Y2=2.91
r72 10 17 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.645 $Y=1.86
+ $X2=1.775 $Y2=1.775
r73 10 12 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=1.645 $Y=1.86
+ $X2=1.645 $Y2=1.98
r74 3 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.91
r75 3 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=1.98
r76 2 14 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.835 $X2=1.61 $Y2=2.91
r77 2 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.835 $X2=1.61 $Y2=1.98
r78 1 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.91
+ $Y=0.235 $X2=3.05 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r43 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r46 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r47 30 39 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.557
+ $Y2=0
r48 30 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=4.08
+ $Y2=0
r49 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r50 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r52 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r53 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.18
+ $Y2=0
r55 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.68
+ $Y2=0
r56 22 39 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.557
+ $Y2=0
r57 22 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.12
+ $Y2=0
r58 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r59 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r60 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.18
+ $Y2=0
r61 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.72
+ $Y2=0
r62 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r63 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r64 11 39 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.557 $Y=0.085
+ $X2=3.557 $Y2=0
r65 11 13 16.1342 $w=2.73e-07 $l=3.85e-07 $layer=LI1_cond $X=3.557 $Y=0.085
+ $X2=3.557 $Y2=0.47
r66 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085 $X2=1.18
+ $Y2=0
r67 7 9 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.52
r68 2 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.26 $X2=3.57 $Y2=0.47
r69 1 9 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=0.885
+ $Y=0.655 $X2=1.18 $Y2=0.52
.ends

