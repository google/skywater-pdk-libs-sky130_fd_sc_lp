* File: sky130_fd_sc_lp__or4b_lp.pex.spice
* Created: Fri Aug 28 11:26:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4B_LP%D_N 3 7 11 15 17 18 19 23
c39 23 0 2.79151e-19 $X=0.62 $Y=1.34
r40 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=1.34 $X2=0.62 $Y2=1.34
r41 19 24 9.85642 $w=3.78e-07 $l=3.25e-07 $layer=LI1_cond $X=0.645 $Y=1.665
+ $X2=0.645 $Y2=1.34
r42 18 24 1.36474 $w=3.78e-07 $l=4.5e-08 $layer=LI1_cond $X=0.645 $Y=1.295
+ $X2=0.645 $Y2=1.34
r43 16 23 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=0.597 $Y=1.658
+ $X2=0.597 $Y2=1.34
r44 16 17 33.0732 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.597 $Y=1.658
+ $X2=0.597 $Y2=1.845
r45 15 23 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.597 $Y=1.325
+ $X2=0.597 $Y2=1.34
r46 7 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.545 $Y=2.545
+ $X2=0.545 $Y2=1.845
r47 1 15 24.6308 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.665 $Y=1.175
+ $X2=0.665 $Y2=1.325
r48 1 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.845 $Y=1.175
+ $X2=0.845 $Y2=0.495
r49 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.485 $Y=1.175
+ $X2=0.485 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%A_27_57# 1 2 7 9 10 12 15 19 25 27 31 33 34
+ 36 40
c69 36 0 2.64321e-19 $X=1.34 $Y=0.99
r70 37 40 31.8098 $w=4.47e-07 $l=2.95e-07 $layer=POLY_cond $X=1.34 $Y=1.16
+ $X2=1.635 $Y2=1.16
r71 37 38 7.00895 $w=4.47e-07 $l=6.5e-08 $layer=POLY_cond $X=1.34 $Y=1.16
+ $X2=1.275 $Y2=1.16
r72 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.34
+ $Y=0.99 $X2=1.34 $Y2=0.99
r73 33 34 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=2.19
+ $X2=0.275 $Y2=2.025
r74 28 31 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=0.91
+ $X2=0.27 $Y2=0.91
r75 27 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=0.91
+ $X2=1.34 $Y2=0.91
r76 27 28 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.175 $Y=0.91
+ $X2=0.435 $Y2=0.91
r77 23 33 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.275 $Y=2.195
+ $X2=0.275 $Y2=2.19
r78 23 25 23.8962 $w=3.38e-07 $l=7.05e-07 $layer=LI1_cond $X=0.275 $Y=2.195
+ $X2=0.275 $Y2=2.9
r79 21 31 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.19 $Y=0.995
+ $X2=0.27 $Y2=0.91
r80 21 34 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.19 $Y=0.995
+ $X2=0.19 $Y2=2.025
r81 17 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=0.825
+ $X2=0.27 $Y2=0.91
r82 17 19 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.27 $Y=0.825
+ $X2=0.27 $Y2=0.495
r83 13 40 37.7405 $w=4.47e-07 $l=4.89643e-07 $layer=POLY_cond $X=1.985 $Y=1.495
+ $X2=1.635 $Y2=1.16
r84 13 15 270.814 $w=2.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.985 $Y=1.495
+ $X2=1.985 $Y2=2.585
r85 10 40 28.6003 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.635 $Y=0.825
+ $X2=1.635 $Y2=1.16
r86 10 12 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.635 $Y=0.825
+ $X2=1.635 $Y2=0.495
r87 7 38 28.6003 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.275 $Y=0.825
+ $X2=1.275 $Y2=1.16
r88 7 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.275 $Y=0.825
+ $X2=1.275 $Y2=0.495
r89 2 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r90 2 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r91 1 19 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.27 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%C 1 3 4 5 6 8 13 15 17 18 19 20 21 22 23 37
+ 38
c61 5 0 6.47666e-20 $X=2.14 $Y=0.855
r62 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.515
+ $Y=1.42 $X2=2.515 $Y2=1.42
r63 22 23 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.4 $Y=2.405 $X2=2.4
+ $Y2=2.775
r64 21 22 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.4 $Y=2.035 $X2=2.4
+ $Y2=2.405
r65 20 21 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.4 $Y=1.665 $X2=2.4
+ $Y2=2.035
r66 20 38 4.12731 $w=7.08e-07 $l=2.45e-07 $layer=LI1_cond $X=2.4 $Y=1.665
+ $X2=2.4 $Y2=1.42
r67 18 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.515 $Y=1.76
+ $X2=2.515 $Y2=1.42
r68 18 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.76
+ $X2=2.515 $Y2=1.925
r69 17 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.255
+ $X2=2.515 $Y2=1.42
r70 13 19 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.475 $Y=2.585
+ $X2=2.475 $Y2=1.925
r71 9 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=0.93
+ $X2=2.425 $Y2=0.855
r72 9 17 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.425 $Y=0.93
+ $X2=2.425 $Y2=1.255
r73 6 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=0.78
+ $X2=2.425 $Y2=0.855
r74 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.425 $Y=0.78 $X2=2.425
+ $Y2=0.495
r75 4 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.35 $Y=0.855
+ $X2=2.425 $Y2=0.855
r76 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.35 $Y=0.855 $X2=2.14
+ $Y2=0.855
r77 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.065 $Y=0.78
+ $X2=2.14 $Y2=0.855
r78 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.065 $Y=0.78 $X2=2.065
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%B 1 3 7 10 12 14 18 20 21 22 23 24 30 31 32
r56 30 32 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.092 $Y=1.42
+ $X2=3.092 $Y2=1.255
r57 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.1 $Y=1.42
+ $X2=3.1 $Y2=1.42
r58 23 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=2.405 $X2=3.1
+ $Y2=2.775
r59 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=2.035 $X2=3.1
+ $Y2=2.405
r60 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=1.665 $X2=3.1
+ $Y2=2.035
r61 21 31 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.1 $Y=1.665
+ $X2=3.1 $Y2=1.42
r62 17 18 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.995 $Y=0.855
+ $X2=3.215 $Y2=0.855
r63 15 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.855 $Y=0.855
+ $X2=2.995 $Y2=0.855
r64 12 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.215 $Y=0.78
+ $X2=3.215 $Y2=0.855
r65 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.215 $Y=0.78
+ $X2=3.215 $Y2=0.495
r66 10 20 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.045 $Y=2.585
+ $X2=3.045 $Y2=1.925
r67 7 20 33.2433 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=3.092 $Y=1.753
+ $X2=3.092 $Y2=1.925
r68 6 30 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=3.092 $Y=1.427
+ $X2=3.092 $Y2=1.42
r69 6 7 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=3.092 $Y=1.427
+ $X2=3.092 $Y2=1.753
r70 4 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.995 $Y=0.93
+ $X2=2.995 $Y2=0.855
r71 4 32 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.995 $Y=0.93
+ $X2=2.995 $Y2=1.255
r72 1 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.855 $Y=0.78
+ $X2=2.855 $Y2=0.855
r73 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.855 $Y=0.78 $X2=2.855
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%A 3 5 7 10 12 14 16 17 18 19 20 21 25
r61 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.695
+ $Y=1.42 $X2=3.695 $Y2=1.42
r62 21 26 6.87299 $w=6.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.08 $Y=1.59
+ $X2=3.695 $Y2=1.59
r63 20 26 1.69593 $w=6.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.6 $Y=1.59
+ $X2=3.695 $Y2=1.59
r64 17 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.695 $Y=1.76
+ $X2=3.695 $Y2=1.42
r65 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.76
+ $X2=3.695 $Y2=1.925
r66 16 25 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.255
+ $X2=3.695 $Y2=1.42
r67 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.005 $Y=0.78
+ $X2=4.005 $Y2=0.495
r68 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.72 $Y=0.855
+ $X2=3.645 $Y2=0.855
r69 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.93 $Y=0.855
+ $X2=4.005 $Y2=0.78
r70 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.93 $Y=0.855
+ $X2=3.72 $Y2=0.855
r71 8 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.645 $Y=0.93
+ $X2=3.645 $Y2=0.855
r72 8 16 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.645 $Y=0.93
+ $X2=3.645 $Y2=1.255
r73 5 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.645 $Y=0.78
+ $X2=3.645 $Y2=0.855
r74 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.645 $Y=0.78 $X2=3.645
+ $Y2=0.495
r75 3 18 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.655 $Y=2.585
+ $X2=3.655 $Y2=1.925
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%A_311_417# 1 2 3 10 12 15 19 21 24 27 31 35
+ 39 41 45 46 48 49 50
r111 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.54
+ $Y=1.335 $X2=4.54 $Y2=1.335
r112 43 45 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=4.54 $Y=1.075
+ $X2=4.54 $Y2=1.335
r113 42 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0.99
+ $X2=3.43 $Y2=0.99
r114 41 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.375 $Y=0.99
+ $X2=4.54 $Y2=1.075
r115 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.375 $Y=0.99
+ $X2=3.595 $Y2=0.99
r116 37 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=0.905
+ $X2=3.43 $Y2=0.99
r117 37 39 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.43 $Y=0.905
+ $X2=3.43 $Y2=0.495
r118 36 49 2.83584 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=0.99
+ $X2=1.85 $Y2=0.99
r119 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0.99
+ $X2=3.43 $Y2=0.99
r120 35 36 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.265 $Y=0.99
+ $X2=2.015 $Y2=0.99
r121 33 49 3.64284 $w=2.55e-07 $l=1.16619e-07 $layer=LI1_cond $X=1.775 $Y=1.075
+ $X2=1.85 $Y2=0.99
r122 33 48 61 $w=1.78e-07 $l=9.9e-07 $layer=LI1_cond $X=1.775 $Y=1.075 $X2=1.775
+ $Y2=2.065
r123 29 49 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.85 $Y=0.905
+ $X2=1.85 $Y2=0.99
r124 29 31 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.85 $Y=0.905
+ $X2=1.85 $Y2=0.495
r125 27 48 8.12648 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=2.23
+ $X2=1.7 $Y2=2.065
r126 24 46 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=4.477 $Y=1.32
+ $X2=4.477 $Y2=1.335
r127 21 46 33.9804 $w=4.55e-07 $l=2.78e-07 $layer=POLY_cond $X=4.477 $Y=1.613
+ $X2=4.477 $Y2=1.335
r128 13 24 24.7927 $w=4.55e-07 $l=1.5e-07 $layer=POLY_cond $X=4.56 $Y=1.17
+ $X2=4.56 $Y2=1.32
r129 13 19 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=4.795 $Y=1.17
+ $X2=4.795 $Y2=0.495
r130 13 15 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=4.435 $Y=1.17
+ $X2=4.435 $Y2=0.495
r131 10 21 44.4147 $w=3.82e-07 $l=4.41597e-07 $layer=POLY_cond $X=4.275 $Y=1.965
+ $X2=4.477 $Y2=1.613
r132 10 12 119.536 $w=2.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.275 $Y=1.965
+ $X2=4.275 $Y2=2.585
r133 3 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.555
+ $Y=2.085 $X2=1.7 $Y2=2.23
r134 2 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.285 $X2=3.43 $Y2=0.495
r135 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.71
+ $Y=0.285 $X2=1.85 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%VPWR 1 2 11 17 19 21 31 32 35 38
r48 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r52 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=3.33
+ $X2=3.92 $Y2=3.33
r53 29 31 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.085 $Y=3.33
+ $X2=5.04 $Y2=3.33
r54 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 25 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 24 27 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 24 25 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 22 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r60 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 21 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.92 $Y2=3.33
r62 21 27 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 19 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 19 25 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 15 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=3.245
+ $X2=3.92 $Y2=3.33
r66 15 17 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=3.92 $Y=3.245
+ $X2=3.92 $Y2=2.27
r67 11 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19 $X2=0.81
+ $Y2=2.9
r68 9 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245 $X2=0.81
+ $Y2=3.33
r69 9 14 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r70 2 17 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=3.78
+ $Y=2.085 $X2=3.92 $Y2=2.27
r71 1 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r72 1 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%X 1 2 7 8 9 10 11 12 13 32
r22 32 39 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=5.05 $Y=2.035 $X2=5.05
+ $Y2=2.065
r23 12 13 5.53186 $w=7.98e-07 $l=3.7e-07 $layer=LI1_cond $X=4.775 $Y=2.405
+ $X2=4.775 $Y2=2.775
r24 12 41 2.61642 $w=7.98e-07 $l=1.75e-07 $layer=LI1_cond $X=4.775 $Y=2.405
+ $X2=4.775 $Y2=2.23
r25 11 41 2.06324 $w=7.98e-07 $l=1.38e-07 $layer=LI1_cond $X=4.775 $Y=2.092
+ $X2=4.775 $Y2=2.23
r26 11 39 6.56939 $w=7.98e-07 $l=2.7e-08 $layer=LI1_cond $X=4.775 $Y=2.092
+ $X2=4.775 $Y2=2.065
r27 11 32 1.29074 $w=2.48e-07 $l=2.8e-08 $layer=LI1_cond $X=5.05 $Y=2.007
+ $X2=5.05 $Y2=2.035
r28 10 11 15.7654 $w=2.48e-07 $l=3.42e-07 $layer=LI1_cond $X=5.05 $Y=1.665
+ $X2=5.05 $Y2=2.007
r29 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=5.05 $Y=1.295
+ $X2=5.05 $Y2=1.665
r30 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=5.05 $Y=0.925 $X2=5.05
+ $Y2=1.295
r31 8 37 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=5.05 $Y=0.925 $X2=5.05
+ $Y2=0.725
r32 7 37 8.73685 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.01 $Y=0.495
+ $X2=5.01 $Y2=0.725
r33 2 41 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.4
+ $Y=2.085 $X2=4.54 $Y2=2.23
r34 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.285 $X2=5.01 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_LP%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r73 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r74 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r75 42 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r76 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r77 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=0 $X2=4.22
+ $Y2=0
r78 39 41 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.385 $Y=0 $X2=5.04
+ $Y2=0
r79 38 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r80 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r81 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.64
+ $Y2=0
r82 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=3.12
+ $Y2=0
r83 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=0 $X2=4.22
+ $Y2=0
r84 34 37 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=4.055 $Y=0 $X2=3.12
+ $Y2=0
r85 33 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r86 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r87 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.06
+ $Y2=0
r88 30 32 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=2.16
+ $Y2=0
r89 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.64
+ $Y2=0
r90 29 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.16
+ $Y2=0
r91 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r92 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r93 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.06
+ $Y2=0
r94 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.72
+ $Y2=0
r95 22 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r96 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r97 22 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r98 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.22 $Y=0.085
+ $X2=4.22 $Y2=0
r99 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.22 $Y=0.085
+ $X2=4.22 $Y2=0.495
r100 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0
r101 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0.495
r102 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0
r103 10 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0.455
r104 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.08
+ $Y=0.285 $X2=4.22 $Y2=0.495
r105 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.285 $X2=2.64 $Y2=0.495
r106 1 12 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.92
+ $Y=0.285 $X2=1.06 $Y2=0.455
.ends

