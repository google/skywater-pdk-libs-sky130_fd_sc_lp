# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o2bb2a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o2bb2a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.210000 1.380000 2.165000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.550000 1.755000 2.000000 2.140000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 1.920000 3.685000 2.210000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.010000 1.110000 3.755000 1.750000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.255000 0.355000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.525000  0.085000 0.875000 0.690000 ;
      RECT 0.525000  0.860000 1.320000 1.030000 ;
      RECT 0.525000  1.030000 0.865000 1.515000 ;
      RECT 0.525000  1.815000 0.855000 2.505000 ;
      RECT 0.525000  2.505000 1.265000 3.245000 ;
      RECT 1.045000  0.280000 2.370000 0.530000 ;
      RECT 1.045000  0.530000 1.320000 0.860000 ;
      RECT 1.435000  2.350000 2.500000 2.480000 ;
      RECT 1.435000  2.480000 1.675000 2.835000 ;
      RECT 1.485000  2.310000 2.500000 2.350000 ;
      RECT 1.550000  0.700000 1.880000 1.405000 ;
      RECT 1.550000  1.405000 2.500000 1.575000 ;
      RECT 1.970000  2.650000 2.300000 3.245000 ;
      RECT 2.075000  0.530000 2.370000 0.620000 ;
      RECT 2.175000  0.620000 2.370000 1.055000 ;
      RECT 2.175000  1.055000 2.840000 1.225000 ;
      RECT 2.240000  1.575000 2.500000 2.310000 ;
      RECT 2.505000  2.650000 2.840000 2.920000 ;
      RECT 2.540000  0.280000 2.765000 0.715000 ;
      RECT 2.540000  0.715000 3.695000 0.885000 ;
      RECT 2.670000  1.225000 2.840000 2.650000 ;
      RECT 2.935000  0.085000 3.265000 0.545000 ;
      RECT 3.325000  2.510000 3.655000 3.245000 ;
      RECT 3.435000  0.280000 3.695000 0.715000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__o2bb2a_1
END LIBRARY
