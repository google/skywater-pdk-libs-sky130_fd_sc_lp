# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xnor3_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__xnor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.180000 7.185000 1.510000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.729000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.345000 3.845000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.345000 1.315000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.575400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.255000 0.440000 1.125000 ;
        RECT 0.100000 1.125000 0.270000 1.815000 ;
        RECT 0.100000 1.815000 0.350000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.440000  1.295000 0.780000 1.625000 ;
      RECT 0.530000  2.290000 0.780000 3.245000 ;
      RECT 0.610000  0.535000 2.575000 0.705000 ;
      RECT 0.610000  0.705000 0.780000 1.295000 ;
      RECT 0.610000  1.625000 0.780000 1.950000 ;
      RECT 0.610000  1.950000 1.120000 2.120000 ;
      RECT 0.650000  0.085000 0.980000 0.365000 ;
      RECT 0.950000  2.120000 1.120000 2.865000 ;
      RECT 0.950000  2.865000 2.505000 3.035000 ;
      RECT 1.195000  0.875000 1.655000 1.125000 ;
      RECT 1.290000  1.950000 1.655000 2.495000 ;
      RECT 1.485000  1.125000 1.655000 1.555000 ;
      RECT 1.485000  1.555000 2.665000 1.885000 ;
      RECT 1.485000  1.885000 1.655000 1.950000 ;
      RECT 1.825000  0.875000 2.075000 1.180000 ;
      RECT 1.825000  1.180000 3.005000 1.385000 ;
      RECT 1.825000  2.235000 2.075000 2.525000 ;
      RECT 1.825000  2.525000 5.210000 2.540000 ;
      RECT 1.825000  2.540000 3.345000 2.695000 ;
      RECT 2.245000  0.525000 2.575000 0.535000 ;
      RECT 2.245000  0.705000 2.575000 1.010000 ;
      RECT 2.745000  0.525000 3.075000 0.615000 ;
      RECT 2.745000  0.615000 6.445000 0.765000 ;
      RECT 2.745000  0.765000 5.080000 0.785000 ;
      RECT 2.745000  0.785000 3.345000 1.010000 ;
      RECT 2.835000  1.385000 3.005000 2.355000 ;
      RECT 3.175000  1.010000 3.345000 2.370000 ;
      RECT 3.175000  2.370000 5.210000 2.525000 ;
      RECT 3.305000  0.085000 3.635000 0.445000 ;
      RECT 3.315000  2.865000 3.645000 3.245000 ;
      RECT 3.745000  1.950000 4.185000 2.030000 ;
      RECT 3.745000  2.030000 4.660000 2.200000 ;
      RECT 3.850000  0.955000 4.185000 1.125000 ;
      RECT 4.015000  1.125000 4.185000 1.950000 ;
      RECT 4.335000  2.710000 4.665000 2.895000 ;
      RECT 4.335000  2.895000 6.945000 3.065000 ;
      RECT 4.410000  0.255000 6.945000 0.425000 ;
      RECT 4.410000  0.425000 4.740000 0.445000 ;
      RECT 4.490000  1.375000 4.785000 1.705000 ;
      RECT 4.490000  1.705000 4.660000 2.030000 ;
      RECT 4.880000  1.875000 5.210000 2.370000 ;
      RECT 4.880000  2.540000 5.210000 2.725000 ;
      RECT 4.910000  0.595000 6.445000 0.615000 ;
      RECT 4.925000  0.955000 5.285000 1.205000 ;
      RECT 4.955000  1.205000 5.285000 1.455000 ;
      RECT 4.955000  1.455000 6.105000 1.625000 ;
      RECT 5.425000  1.845000 5.755000 2.515000 ;
      RECT 5.425000  2.515000 6.445000 2.685000 ;
      RECT 5.455000  0.935000 5.785000 1.115000 ;
      RECT 5.455000  1.115000 6.565000 1.285000 ;
      RECT 5.935000  1.625000 6.105000 2.345000 ;
      RECT 6.115000  0.765000 6.445000 0.940000 ;
      RECT 6.275000  1.285000 6.565000 1.675000 ;
      RECT 6.275000  1.675000 6.445000 2.515000 ;
      RECT 6.615000  0.425000 6.945000 0.775000 ;
      RECT 6.615000  0.775000 7.525000 0.945000 ;
      RECT 6.615000  1.845000 7.525000 2.175000 ;
      RECT 6.615000  2.175000 6.945000 2.895000 ;
      RECT 7.115000  0.085000 7.445000 0.605000 ;
      RECT 7.160000  2.345000 7.490000 3.245000 ;
      RECT 7.355000  0.945000 7.525000 1.190000 ;
      RECT 7.355000  1.190000 7.645000 1.520000 ;
      RECT 7.355000  1.520000 7.525000 1.845000 ;
      RECT 7.695000  0.340000 8.075000 1.020000 ;
      RECT 7.695000  1.895000 8.075000 2.935000 ;
      RECT 7.835000  1.020000 8.075000 1.895000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.210000 2.725000 1.380000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  1.210000 5.125000 1.380000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  2.320000 5.605000 2.490000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  2.320000 8.005000 2.490000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
    LAYER met1 ;
      RECT 2.495000 1.180000 2.785000 1.225000 ;
      RECT 2.495000 1.225000 5.185000 1.365000 ;
      RECT 2.495000 1.365000 2.785000 1.410000 ;
      RECT 4.895000 1.180000 5.185000 1.225000 ;
      RECT 4.895000 1.365000 5.185000 1.410000 ;
      RECT 5.375000 2.290000 5.665000 2.335000 ;
      RECT 5.375000 2.335000 8.065000 2.475000 ;
      RECT 5.375000 2.475000 5.665000 2.520000 ;
      RECT 7.775000 2.290000 8.065000 2.335000 ;
      RECT 7.775000 2.475000 8.065000 2.520000 ;
  END
END sky130_fd_sc_lp__xnor3_1
