* File: sky130_fd_sc_lp__a41oi_1.pxi.spice
* Created: Wed Sep  2 09:29:34 2020
* 
x_PM_SKY130_FD_SC_LP__A41OI_1%B1 N_B1_c_54_n N_B1_M1007_g N_B1_M1001_g
+ N_B1_c_56_n N_B1_c_57_n B1 PM_SKY130_FD_SC_LP__A41OI_1%B1
x_PM_SKY130_FD_SC_LP__A41OI_1%A4 N_A4_M1004_g N_A4_M1009_g A4 A4 N_A4_c_84_n
+ PM_SKY130_FD_SC_LP__A41OI_1%A4
x_PM_SKY130_FD_SC_LP__A41OI_1%A3 N_A3_M1002_g N_A3_M1000_g A3 A3 N_A3_c_125_n
+ PM_SKY130_FD_SC_LP__A41OI_1%A3
x_PM_SKY130_FD_SC_LP__A41OI_1%A2 N_A2_M1008_g N_A2_M1006_g A2 A2 N_A2_c_161_n
+ N_A2_c_162_n PM_SKY130_FD_SC_LP__A41OI_1%A2
x_PM_SKY130_FD_SC_LP__A41OI_1%A1 N_A1_M1003_g N_A1_M1005_g A1 A1 N_A1_c_195_n
+ N_A1_c_196_n PM_SKY130_FD_SC_LP__A41OI_1%A1
x_PM_SKY130_FD_SC_LP__A41OI_1%Y N_Y_M1007_s N_Y_M1003_d N_Y_M1001_s N_Y_c_218_n
+ N_Y_c_223_n N_Y_c_219_n N_Y_c_220_n Y Y Y N_Y_c_225_n Y N_Y_c_222_n
+ PM_SKY130_FD_SC_LP__A41OI_1%Y
x_PM_SKY130_FD_SC_LP__A41OI_1%A_128_367# N_A_128_367#_M1001_d
+ N_A_128_367#_M1000_d N_A_128_367#_M1005_d N_A_128_367#_c_278_n
+ N_A_128_367#_c_279_n N_A_128_367#_c_281_n N_A_128_367#_c_315_p
+ N_A_128_367#_c_294_n N_A_128_367#_c_276_n N_A_128_367#_c_277_n
+ N_A_128_367#_c_283_n N_A_128_367#_c_286_n N_A_128_367#_c_291_n
+ PM_SKY130_FD_SC_LP__A41OI_1%A_128_367#
x_PM_SKY130_FD_SC_LP__A41OI_1%VPWR N_VPWR_M1004_d N_VPWR_M1008_d N_VPWR_c_335_n
+ N_VPWR_c_324_n N_VPWR_c_325_n VPWR N_VPWR_c_326_n N_VPWR_c_327_n
+ N_VPWR_c_328_n N_VPWR_c_323_n N_VPWR_c_330_n N_VPWR_c_331_n
+ PM_SKY130_FD_SC_LP__A41OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A41OI_1%VGND N_VGND_M1007_d VGND N_VGND_c_373_n
+ N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n PM_SKY130_FD_SC_LP__A41OI_1%VGND
cc_1 VNB N_B1_c_54_n 0.0250732f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.185
cc_2 VNB N_B1_M1001_g 0.0109075f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_3 VNB N_B1_c_56_n 0.0388165f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.35
cc_4 VNB N_B1_c_57_n 0.0106698f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.35
cc_5 VNB B1 0.017405f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A4_M1004_g 0.00744465f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.655
cc_7 VNB N_A4_M1009_g 0.0207574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A4 0.00423003f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.35
cc_9 VNB N_A4_c_84_n 0.0543649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A3_M1002_g 0.0188544f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.655
cc_11 VNB N_A3_M1000_g 0.00723896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A3 0.00704458f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.35
cc_13 VNB N_A3_c_125_n 0.0307152f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.35
cc_14 VNB N_A2_M1008_g 0.00614389f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.655
cc_15 VNB A2 0.0069502f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.35
cc_16 VNB N_A2_c_161_n 0.0307309f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.35
cc_17 VNB N_A2_c_162_n 0.0178391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1005_g 0.00900329f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_19 VNB A1 0.0209376f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.35
cc_20 VNB N_A1_c_195_n 0.0395145f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.35
cc_21 VNB N_A1_c_196_n 0.0224093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_218_n 0.0218244f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.35
cc_23 VNB N_Y_c_219_n 0.00755746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_220_n 0.0223155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB Y 0.00513794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_222_n 0.00784917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_323_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_373_n 0.0605948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_374_n 0.19226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_375_n 0.0182809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_376_n 0.0151186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_B1_M1001_g 0.0251186f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.465
cc_33 VPB N_A4_M1004_g 0.0259292f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.655
cc_34 VPB A4 0.00291351f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.35
cc_35 VPB N_A3_M1000_g 0.0255137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB A3 0.00452261f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.35
cc_37 VPB N_A2_M1008_g 0.019662f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.655
cc_38 VPB A2 0.00438532f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.35
cc_39 VPB N_A1_M1005_g 0.0265838f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.465
cc_40 VPB A1 0.00705314f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.35
cc_41 VPB N_Y_c_223_n 0.0459084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB Y 9.5111e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_Y_c_225_n 0.0119377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_128_367#_c_276_n 0.00755006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_128_367#_c_277_n 0.0376446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_324_n 0.00274626f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_47 VPB N_VPWR_c_325_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.35
cc_48 VPB N_VPWR_c_326_n 0.0300411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_327_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_328_n 0.0158241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_323_n 0.0484002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_330_n 0.0139417f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_331_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 N_B1_M1001_g N_A4_M1004_g 0.0148706f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_55 N_B1_c_57_n A4 3.96174e-19 $X=0.565 $Y=1.35 $X2=0 $Y2=0
cc_56 N_B1_c_57_n N_A4_c_84_n 0.0148706f $X=0.565 $Y=1.35 $X2=0 $Y2=0
cc_57 N_B1_c_54_n Y 0.0111978f $X=0.565 $Y=1.185 $X2=0 $Y2=0
cc_58 N_B1_M1001_g Y 0.0103169f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_59 N_B1_c_57_n Y 0.0102109f $X=0.565 $Y=1.35 $X2=0 $Y2=0
cc_60 B1 Y 0.0244747f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_B1_M1001_g N_Y_c_225_n 0.0167354f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_62 N_B1_c_56_n N_Y_c_225_n 0.00803968f $X=0.49 $Y=1.35 $X2=0 $Y2=0
cc_63 B1 N_Y_c_225_n 0.0158375f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_64 N_B1_c_54_n N_Y_c_222_n 0.0140582f $X=0.565 $Y=1.185 $X2=0 $Y2=0
cc_65 N_B1_c_56_n N_Y_c_222_n 0.00712992f $X=0.49 $Y=1.35 $X2=0 $Y2=0
cc_66 B1 N_Y_c_222_n 0.0163665f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B1_M1001_g N_A_128_367#_c_278_n 0.00214926f $X=0.565 $Y=2.465 $X2=0
+ $Y2=0
cc_68 N_B1_M1001_g N_A_128_367#_c_279_n 0.00962096f $X=0.565 $Y=2.465 $X2=0
+ $Y2=0
cc_69 N_B1_M1001_g N_VPWR_c_324_n 0.00112429f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_70 N_B1_M1001_g N_VPWR_c_326_n 0.0054895f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_71 N_B1_M1001_g N_VPWR_c_323_n 0.0110726f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_72 N_B1_c_54_n N_VGND_c_374_n 0.00551899f $X=0.565 $Y=1.185 $X2=0 $Y2=0
cc_73 N_B1_c_54_n N_VGND_c_375_n 0.00486043f $X=0.565 $Y=1.185 $X2=0 $Y2=0
cc_74 N_B1_c_54_n N_VGND_c_376_n 0.0148328f $X=0.565 $Y=1.185 $X2=0 $Y2=0
cc_75 N_A4_M1009_g N_A3_M1002_g 0.052499f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_76 A4 N_A3_M1000_g 7.05268e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A4_M1004_g A3 9.72917e-19 $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A4_M1009_g A3 0.00323109f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_79 A4 A3 0.0481628f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 A4 N_A3_c_125_n 2.23812e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A4_c_84_n N_A3_c_125_n 0.021098f $X=1.445 $Y=1.375 $X2=0 $Y2=0
cc_82 N_A4_M1009_g N_Y_c_219_n 0.0180202f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_83 A4 N_Y_c_219_n 0.02416f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A4_c_84_n N_Y_c_219_n 0.00454693f $X=1.445 $Y=1.375 $X2=0 $Y2=0
cc_85 N_A4_M1009_g Y 0.00418852f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_86 A4 Y 0.0407529f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A4_c_84_n Y 0.0040325f $X=1.445 $Y=1.375 $X2=0 $Y2=0
cc_88 N_A4_M1004_g N_Y_c_225_n 0.0038605f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_89 A4 N_Y_c_225_n 0.0045419f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A4_M1009_g N_Y_c_222_n 2.59997e-19 $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_91 N_A4_M1004_g N_A_128_367#_c_279_n 0.00440279f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A4_M1004_g N_A_128_367#_c_281_n 0.011864f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_93 A4 N_A_128_367#_c_281_n 0.00367087f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A4_M1004_g N_A_128_367#_c_283_n 0.00789197f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_95 A4 N_A_128_367#_c_283_n 0.0117465f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A4_c_84_n N_A_128_367#_c_283_n 6.2048e-19 $X=1.445 $Y=1.375 $X2=0 $Y2=0
cc_97 N_A4_M1004_g N_A_128_367#_c_286_n 8.70195e-19 $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_98 A4 N_A_128_367#_c_286_n 0.00553776f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A4_c_84_n N_A_128_367#_c_286_n 0.00573337f $X=1.445 $Y=1.375 $X2=0 $Y2=0
cc_100 N_A4_M1004_g N_VPWR_c_335_n 0.00863723f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A4_M1004_g N_VPWR_c_324_n 0.010705f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A4_M1004_g N_VPWR_c_326_n 0.00388479f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A4_M1004_g N_VPWR_c_323_n 0.00685293f $X=1.05 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A4_M1009_g N_VGND_c_373_n 0.00486043f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_105 N_A4_M1009_g N_VGND_c_374_n 0.00461704f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_106 N_A4_M1009_g N_VGND_c_376_n 0.0179082f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_107 A3 N_A2_M1008_g 2.68115e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_108 N_A3_c_125_n N_A2_M1008_g 0.0248457f $X=1.895 $Y=1.375 $X2=0 $Y2=0
cc_109 A3 A2 0.0401175f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A3_c_125_n A2 0.00253346f $X=1.895 $Y=1.375 $X2=0 $Y2=0
cc_111 N_A3_M1002_g N_A2_c_161_n 8.829e-19 $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_112 A3 N_A2_c_161_n 0.00124423f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_113 N_A3_c_125_n N_A2_c_161_n 0.0185869f $X=1.895 $Y=1.375 $X2=0 $Y2=0
cc_114 N_A3_M1002_g N_A2_c_162_n 0.0357776f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_115 N_A3_M1002_g N_Y_c_219_n 0.0126288f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_116 A3 N_Y_c_219_n 0.0366419f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A3_c_125_n N_Y_c_219_n 9.02157e-19 $X=1.895 $Y=1.375 $X2=0 $Y2=0
cc_118 N_A3_M1000_g N_A_128_367#_c_283_n 0.00244005f $X=1.985 $Y=2.465 $X2=0
+ $Y2=0
cc_119 A3 N_A_128_367#_c_286_n 0.00871239f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_120 N_A3_M1000_g N_A_128_367#_c_291_n 0.0142423f $X=1.985 $Y=2.465 $X2=0
+ $Y2=0
cc_121 A3 N_A_128_367#_c_291_n 0.0317112f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A3_c_125_n N_A_128_367#_c_291_n 6.89016e-19 $X=1.895 $Y=1.375 $X2=0
+ $Y2=0
cc_123 N_A3_M1000_g N_VPWR_c_335_n 0.0103032f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A3_M1000_g N_VPWR_c_324_n 0.00831425f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A3_M1000_g N_VPWR_c_325_n 6.54575e-19 $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A3_M1000_g N_VPWR_c_327_n 0.00486043f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A3_M1000_g N_VPWR_c_323_n 0.0082726f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A3_M1002_g N_VGND_c_373_n 0.00585385f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_129 N_A3_M1002_g N_VGND_c_374_n 0.00689897f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A3_M1002_g N_VGND_c_376_n 0.00317246f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_131 N_A2_M1008_g N_A1_M1005_g 0.0370494f $X=2.415 $Y=2.465 $X2=0 $Y2=0
cc_132 A2 A1 0.0462774f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A2_c_161_n A1 2.62349e-19 $X=2.435 $Y=1.35 $X2=0 $Y2=0
cc_134 N_A2_c_161_n N_A1_c_195_n 0.0205067f $X=2.435 $Y=1.35 $X2=0 $Y2=0
cc_135 A2 N_A1_c_196_n 0.00465077f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A2_c_162_n N_A1_c_196_n 0.0488851f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_137 A2 N_Y_c_219_n 0.033994f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A2_c_161_n N_Y_c_219_n 9.7882e-19 $X=2.435 $Y=1.35 $X2=0 $Y2=0
cc_139 N_A2_c_162_n N_Y_c_219_n 0.0126873f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_140 N_A2_c_162_n N_Y_c_220_n 0.00276498f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A2_M1008_g N_A_128_367#_c_294_n 0.0129889f $X=2.415 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A2_c_161_n N_A_128_367#_c_294_n 3.71353e-19 $X=2.435 $Y=1.35 $X2=0
+ $Y2=0
cc_143 A2 N_A_128_367#_c_291_n 0.0339619f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A2_c_161_n N_A_128_367#_c_291_n 2.04278e-19 $X=2.435 $Y=1.35 $X2=0
+ $Y2=0
cc_145 N_A2_M1008_g N_VPWR_c_324_n 5.52132e-19 $X=2.415 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A2_M1008_g N_VPWR_c_325_n 0.0130514f $X=2.415 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A2_M1008_g N_VPWR_c_327_n 0.00564095f $X=2.415 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A2_M1008_g N_VPWR_c_323_n 0.00950825f $X=2.415 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A2_c_162_n N_VGND_c_373_n 0.00585385f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_150 N_A2_c_162_n N_VGND_c_374_n 0.00692489f $X=2.435 $Y=1.185 $X2=0 $Y2=0
cc_151 A1 N_Y_c_219_n 0.0261078f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A1_c_195_n N_Y_c_219_n 0.00147112f $X=3.005 $Y=1.35 $X2=0 $Y2=0
cc_153 N_A1_c_196_n N_Y_c_219_n 0.0127848f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_154 N_A1_c_196_n N_Y_c_220_n 0.0127134f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_155 N_A1_M1005_g N_A_128_367#_c_294_n 0.0163836f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_156 A1 N_A_128_367#_c_294_n 0.00402539f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_157 A1 N_A_128_367#_c_276_n 0.0240081f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A1_c_195_n N_A_128_367#_c_276_n 8.00916e-19 $X=3.005 $Y=1.35 $X2=0
+ $Y2=0
cc_159 N_A1_M1005_g N_VPWR_c_325_n 0.0148711f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A1_M1005_g N_VPWR_c_328_n 0.00564095f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A1_M1005_g N_VPWR_c_323_n 0.0104155f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A1_c_196_n N_VGND_c_373_n 0.00549284f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_163 N_A1_c_196_n N_VGND_c_374_n 0.0072441f $X=2.99 $Y=1.185 $X2=0 $Y2=0
cc_164 N_Y_c_225_n N_A_128_367#_M1001_d 0.00227021f $X=0.722 $Y=1.695 $X2=-0.19
+ $Y2=-0.245
cc_165 N_Y_c_225_n N_A_128_367#_c_278_n 0.0159373f $X=0.722 $Y=1.695 $X2=0 $Y2=0
cc_166 N_Y_c_223_n N_VPWR_c_326_n 0.0178111f $X=0.35 $Y=1.98 $X2=0 $Y2=0
cc_167 N_Y_M1001_s N_VPWR_c_323_n 0.00371702f $X=0.225 $Y=1.835 $X2=0 $Y2=0
cc_168 N_Y_c_223_n N_VPWR_c_323_n 0.0100304f $X=0.35 $Y=1.98 $X2=0 $Y2=0
cc_169 N_Y_c_219_n N_VGND_M1007_d 0.0146631f $X=2.935 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_170 Y N_VGND_M1007_d 0.00163933f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_171 N_Y_c_222_n N_VGND_M1007_d 0.00298607f $X=0.87 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_172 N_Y_c_220_n N_VGND_c_373_n 0.0197852f $X=3.1 $Y=0.43 $X2=0 $Y2=0
cc_173 N_Y_M1007_s N_VGND_c_374_n 0.00244875f $X=0.225 $Y=0.235 $X2=0 $Y2=0
cc_174 N_Y_M1003_d N_VGND_c_374_n 0.00215406f $X=2.96 $Y=0.235 $X2=0 $Y2=0
cc_175 N_Y_c_218_n N_VGND_c_374_n 0.0099354f $X=0.35 $Y=0.43 $X2=0 $Y2=0
cc_176 N_Y_c_219_n N_VGND_c_374_n 0.049492f $X=2.935 $Y=0.92 $X2=0 $Y2=0
cc_177 N_Y_c_220_n N_VGND_c_374_n 0.012508f $X=3.1 $Y=0.43 $X2=0 $Y2=0
cc_178 N_Y_c_222_n N_VGND_c_374_n 0.00755245f $X=0.87 $Y=0.925 $X2=0 $Y2=0
cc_179 N_Y_c_218_n N_VGND_c_375_n 0.0165299f $X=0.35 $Y=0.43 $X2=0 $Y2=0
cc_180 N_Y_c_222_n N_VGND_c_376_n 0.0524082f $X=0.87 $Y=0.925 $X2=0 $Y2=0
cc_181 N_Y_c_219_n A_304_47# 0.00505953f $X=2.935 $Y=0.92 $X2=-0.19 $Y2=-0.245
cc_182 N_Y_c_219_n A_390_47# 0.0155644f $X=2.935 $Y=0.92 $X2=-0.19 $Y2=-0.245
cc_183 N_Y_c_219_n A_504_47# 0.00530001f $X=2.935 $Y=0.92 $X2=-0.19 $Y2=-0.245
cc_184 N_A_128_367#_c_283_n N_VPWR_M1004_d 0.0044121f $X=1.2 $Y=2.01 $X2=-0.19
+ $Y2=1.655
cc_185 N_A_128_367#_c_286_n N_VPWR_M1004_d 0.0119631f $X=1.635 $Y=2.007
+ $X2=-0.19 $Y2=1.655
cc_186 N_A_128_367#_c_291_n N_VPWR_M1004_d 0.00535514f $X=2.315 $Y=2.007
+ $X2=-0.19 $Y2=1.655
cc_187 N_A_128_367#_c_294_n N_VPWR_M1008_d 0.00425838f $X=2.985 $Y=2.005 $X2=0
+ $Y2=0
cc_188 N_A_128_367#_c_279_n N_VPWR_c_335_n 0.0388485f $X=0.78 $Y=2.525 $X2=0
+ $Y2=0
cc_189 N_A_128_367#_c_281_n N_VPWR_c_335_n 0.00304701f $X=1.115 $Y=2.12 $X2=0
+ $Y2=0
cc_190 N_A_128_367#_c_283_n N_VPWR_c_335_n 0.00930091f $X=1.2 $Y=2.01 $X2=0
+ $Y2=0
cc_191 N_A_128_367#_c_286_n N_VPWR_c_335_n 0.043809f $X=1.635 $Y=2.007 $X2=0
+ $Y2=0
cc_192 N_A_128_367#_c_279_n N_VPWR_c_324_n 0.0218986f $X=0.78 $Y=2.525 $X2=0
+ $Y2=0
cc_193 N_A_128_367#_c_294_n N_VPWR_c_325_n 0.017285f $X=2.985 $Y=2.005 $X2=0
+ $Y2=0
cc_194 N_A_128_367#_c_279_n N_VPWR_c_326_n 0.0181806f $X=0.78 $Y=2.525 $X2=0
+ $Y2=0
cc_195 N_A_128_367#_c_315_p N_VPWR_c_327_n 0.0131621f $X=2.2 $Y=2.46 $X2=0 $Y2=0
cc_196 N_A_128_367#_c_277_n N_VPWR_c_328_n 0.0185207f $X=3.1 $Y=2.46 $X2=0 $Y2=0
cc_197 N_A_128_367#_M1001_d N_VPWR_c_323_n 0.00511301f $X=0.64 $Y=1.835 $X2=0
+ $Y2=0
cc_198 N_A_128_367#_M1000_d N_VPWR_c_323_n 0.00467071f $X=2.06 $Y=1.835 $X2=0
+ $Y2=0
cc_199 N_A_128_367#_M1005_d N_VPWR_c_323_n 0.00302127f $X=2.96 $Y=1.835 $X2=0
+ $Y2=0
cc_200 N_A_128_367#_c_279_n N_VPWR_c_323_n 0.0110138f $X=0.78 $Y=2.525 $X2=0
+ $Y2=0
cc_201 N_A_128_367#_c_315_p N_VPWR_c_323_n 0.00808656f $X=2.2 $Y=2.46 $X2=0
+ $Y2=0
cc_202 N_A_128_367#_c_277_n N_VPWR_c_323_n 0.010808f $X=3.1 $Y=2.46 $X2=0 $Y2=0
cc_203 N_VGND_c_374_n A_304_47# 0.00408795f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_204 N_VGND_c_374_n A_390_47# 0.0061521f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_205 N_VGND_c_374_n A_504_47# 0.00423395f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
