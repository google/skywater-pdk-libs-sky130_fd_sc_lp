# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrtn_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrtn_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.460000 1.110000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.030000 2.055000 7.565000 3.065000 ;
        RECT 7.235000 0.265000 7.565000 2.055000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.205000 6.500000 1.875000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.030000 1.120000 1.360000 1.790000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.110000  0.265000 0.445000 0.675000 ;
      RECT 0.110000  0.675000 0.280000 2.055000 ;
      RECT 0.110000  2.055000 0.565000 2.495000 ;
      RECT 0.110000  2.495000 1.445000 2.665000 ;
      RECT 0.110000  2.665000 0.565000 3.065000 ;
      RECT 0.765000  2.845000 1.095000 3.245000 ;
      RECT 0.905000  0.085000 1.235000 0.675000 ;
      RECT 1.275000  2.665000 2.575000 2.835000 ;
      RECT 1.295000  2.055000 1.875000 2.315000 ;
      RECT 1.570000  0.295000 2.055000 0.485000 ;
      RECT 1.570000  0.485000 1.875000 2.055000 ;
      RECT 2.055000  0.665000 4.645000 0.835000 ;
      RECT 2.055000  0.835000 2.225000 2.485000 ;
      RECT 2.315000  0.265000 2.645000 0.665000 ;
      RECT 2.405000  1.585000 3.230000 1.915000 ;
      RECT 2.405000  1.915000 2.575000 2.665000 ;
      RECT 2.440000  1.015000 4.130000 1.345000 ;
      RECT 2.755000  2.095000 3.005000 3.245000 ;
      RECT 3.105000  0.085000 3.435000 0.485000 ;
      RECT 3.440000  1.585000 4.480000 1.755000 ;
      RECT 3.440000  1.755000 3.770000 1.915000 ;
      RECT 3.950000  2.055000 4.995000 2.225000 ;
      RECT 3.950000  2.225000 4.280000 3.065000 ;
      RECT 4.035000  0.295000 4.995000 0.485000 ;
      RECT 4.310000  0.835000 4.645000 1.435000 ;
      RECT 4.310000  1.435000 4.480000 1.585000 ;
      RECT 4.825000  0.485000 4.995000 1.425000 ;
      RECT 4.825000  1.425000 5.705000 1.755000 ;
      RECT 4.825000  1.755000 4.995000 2.055000 ;
      RECT 5.175000  0.085000 5.425000 0.675000 ;
      RECT 5.175000  0.855000 7.040000 1.025000 ;
      RECT 5.175000  1.025000 5.505000 1.185000 ;
      RECT 5.175000  2.055000 5.505000 3.245000 ;
      RECT 5.655000  0.265000 5.985000 0.855000 ;
      RECT 5.865000  2.055000 6.850000 2.225000 ;
      RECT 5.865000  2.225000 6.195000 3.065000 ;
      RECT 6.395000  2.405000 6.725000 3.245000 ;
      RECT 6.445000  0.085000 6.775000 0.675000 ;
      RECT 6.680000  1.025000 7.040000 1.525000 ;
      RECT 6.680000  1.525000 6.850000 2.055000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrtn_lp
