* NGSPICE file created from sky130_fd_sc_lp__ha_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__ha_2 A B VGND VNB VPB VPWR COUT SUM
M1000 VGND a_227_397# SUM VNB nshort w=840000u l=150000u
+  ad=9.996e+11p pd=8.71e+06u as=2.352e+11p ps=2.24e+06u
M1001 VGND A a_492_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1002 SUM a_227_397# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.7551e+12p ps=1.389e+07u
M1003 VPWR a_270_95# a_227_397# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.496e+11p ps=2.06e+06u
M1004 a_492_131# B a_270_95# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VGND a_270_95# COUT VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 a_227_397# B a_155_397# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1007 VPWR A a_270_95# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1008 VPWR a_270_95# COUT VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1009 a_45_121# B VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1010 VGND A a_45_121# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_227_397# a_270_95# a_45_121# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1012 SUM a_227_397# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_155_397# A VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_270_95# B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 COUT a_270_95# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 COUT a_270_95# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_227_397# SUM VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

