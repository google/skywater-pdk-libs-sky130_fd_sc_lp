* File: sky130_fd_sc_lp__o311a_0.spice
* Created: Wed Sep  2 10:22:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311a_0.pex.spice"
.subckt sky130_fd_sc_lp__o311a_0  VNB VPB A1 A2 A3 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_96_161#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.2541 PD=0.74 PS=2.05 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.5
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1011 N_A_292_55#_M1011_d N_A1_M1011_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_292_55#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_292_55#_M1004_d N_A3_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.9
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_564_55# N_B1_M1008_g N_A_292_55#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_96_161#_M1010_d N_C1_M1010_g A_564_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_96_161#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.1696 PD=1.03 PS=1.81 NRD=16.9223 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1003 A_270_481# N_A1_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64 AD=0.096
+ AS=0.1248 PD=0.94 PS=1.03 NRD=29.2348 NRS=16.9223 M=1 R=4.26667 SA=75000.7
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1006 A_360_481# N_A2_M1006_g A_270_481# VPB PHIGHVT L=0.15 W=0.64 AD=0.096
+ AS=0.096 PD=0.94 PS=0.94 NRD=29.2348 NRS=29.2348 M=1 R=4.26667 SA=75001.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_96_161#_M1007_d N_A3_M1007_g A_360_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0992 AS=0.096 PD=0.95 PS=0.94 NRD=4.6098 NRS=29.2348 M=1 R=4.26667
+ SA=75001.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g N_A_96_161#_M1007_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.112 AS=0.0992 PD=0.99 PS=0.95 NRD=16.9223 NRS=4.6098 M=1 R=4.26667
+ SA=75002.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1001 N_A_96_161#_M1001_d N_C1_M1001_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.112 PD=1.81 PS=0.99 NRD=0 NRS=4.6098 M=1 R=4.26667 SA=75002.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o311a_0.pxi.spice"
*
.ends
*
*
