* NGSPICE file created from sky130_fd_sc_lp__a2111o_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111o_m A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_503_47# A1 a_85_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_85_21# D1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4.389e+11p ps=4.61e+06u
M1002 VGND A2 a_503_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_339_369# C1 a_267_369# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1004 a_411_369# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.457e+11p ps=2.85e+06u
M1005 VPWR A1 a_411_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C1 a_85_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_85_21# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_411_369# B1 a_339_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_85_21# B1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_85_21# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 a_267_369# D1 a_85_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

