* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_m A B VGND VNB VPB VPWR X
X0 a_124_535# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_41_535# B a_124_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_282_535# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR A a_282_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_357_156# B X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_41_535# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND B a_41_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_282_535# a_41_535# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_41_535# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND A a_357_156# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
