* File: sky130_fd_sc_lp__sdlclkp_1.spice
* Created: Fri Aug 28 11:31:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdlclkp_1.pex.spice"
.subckt sky130_fd_sc_lp__sdlclkp_1  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1011 N_A_154_69#_M1011_d N_SCE_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.126 PD=0.7 PS=1.44 NRD=0 NRS=7.14 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_GATE_M1018_g N_A_154_69#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_334_69#_M1016_d N_A_254_357#_M1016_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_623_133#_M1019_d N_A_254_357#_M1019_g N_A_154_69#_M1019_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0714 AS=0.1281 PD=0.76 PS=1.45 NRD=17.136 NRS=5.712 M=1
+ R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 A_721_133# N_A_334_69#_M1006_g N_A_623_133#_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0714 PD=0.63 PS=0.76 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_737_329#_M1000_g A_721_133# VNB NSHORT L=0.15 W=0.42
+ AD=0.123333 AS=0.0441 PD=0.926667 PS=0.63 NRD=68.184 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1021 N_A_737_329#_M1021_d N_A_623_133#_M1021_g N_VGND_M1000_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.246667 PD=2.25 PS=1.85333 NRD=0 NRS=12.132 M=1
+ R=5.6 SA=75001 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_CLK_M1003_g N_A_254_357#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1012 A_1194_52# N_CLK_M1012_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_1231_367#_M1013_d N_A_737_329#_M1013_g A_1194_52# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_GCLK_M1005_d N_A_1231_367#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 A_110_468# N_SCE_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1015 N_A_154_69#_M1015_d N_GATE_M1015_g A_110_468# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_334_69#_M1004_d N_A_254_357#_M1004_g N_VPWR_M1004_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.3296 PD=1.85 PS=2.31 NRD=3.0732 NRS=73.8553 M=1
+ R=4.26667 SA=75000.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_623_133#_M1001_d N_A_334_69#_M1001_g N_A_154_69#_M1001_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1017 A_736_463# N_A_254_357#_M1017_g N_A_623_133#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_737_329#_M1009_g A_736_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09765 AS=0.0441 PD=0.83 PS=0.63 NRD=56.2829 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1014 N_A_737_329#_M1014_d N_A_623_133#_M1014_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.29295 PD=3.05 PS=2.49 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_CLK_M1007_g N_A_254_357#_M1007_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.18575 AS=0.1824 PD=1.39 PS=1.85 NRD=72.3975 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_1231_367#_M1002_d N_CLK_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.18575 PD=0.92 PS=1.39 NRD=0 NRS=72.3975 M=1 R=4.26667
+ SA=75000.8 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_737_329#_M1008_g N_A_1231_367#_M1002_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.132952 AS=0.0896 PD=1.09137 PS=0.92 NRD=24.6053 NRS=0 M=1
+ R=4.26667 SA=75001.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1010 N_GCLK_M1010_d N_A_1231_367#_M1010_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.261748 PD=3.05 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.0631 P=19.91
*
.include "sky130_fd_sc_lp__sdlclkp_1.pxi.spice"
*
.ends
*
*
