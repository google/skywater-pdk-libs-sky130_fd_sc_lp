* File: sky130_fd_sc_lp__fa_2.spice
* Created: Fri Aug 28 10:34:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fa_2.pex.spice"
.subckt sky130_fd_sc_lp__fa_2  VNB VPB A CIN B VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* B	B
* CIN	CIN
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_84_21#_M1007_g N_SUM_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A_84_21#_M1008_g N_SUM_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1904 AS=0.1176 PD=1.64667 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1023 N_A_309_131#_M1023_d N_B_M1023_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.123675 AS=0.0952 PD=1.06 PS=0.823333 NRD=34.284 NRS=49.044 M=1 R=2.8
+ SA=75001.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1018 N_A_395_398#_M1018_d N_CIN_M1018_g N_A_309_131#_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.123675 PD=1.37 PS=1.06 NRD=0 NRS=68.412 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_309_131#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75005.5
+ A=0.063 P=1.14 MULT=1
MM1002 A_710_119# N_A_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6 SB=75005.1
+ A=0.063 P=1.14 MULT=1
MM1029 A_782_119# N_B_M1029_g A_710_119# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001 SB=75004.7
+ A=0.063 P=1.14 MULT=1
MM1019 N_A_84_21#_M1019_d N_CIN_M1019_g A_782_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1022 N_A_940_119#_M1022_d N_A_395_398#_M1022_g N_A_84_21#_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.8 SB=75004 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_CIN_M1015_g N_A_940_119#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.13755 AS=0.0588 PD=1.075 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1024 N_A_940_119#_M1024_d N_B_M1024_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.13755 PD=0.7 PS=1.075 NRD=0 NRS=0 M=1 R=2.8 SA=75003 SB=75002.7
+ A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_M1026_g N_A_940_119#_M1024_d VNB NSHORT L=0.15 W=0.42
+ AD=0.130167 AS=0.0588 PD=0.963333 PS=0.7 NRD=72.828 NRS=0 M=1 R=2.8 SA=75003.4
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1004 N_COUT_M1004_d N_A_395_398#_M1004_g N_VGND_M1026_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.260333 PD=1.12 PS=1.92667 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75002.2 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1016 N_COUT_M1004_d N_A_395_398#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.321933 PD=1.12 PS=2.22 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75002.6 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1009 A_1653_137# N_A_M1009_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.160967 PD=0.63 PS=1.11 NRD=14.28 NRS=93.78 M=1 R=2.8 SA=75004.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_395_398#_M1006_d N_B_M1006_g A_1653_137# VNB NSHORT L=0.15 W=0.42
+ AD=0.1512 AS=0.0441 PD=1.56 PS=0.63 NRD=27.132 NRS=14.28 M=1 R=2.8 SA=75004.9
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1020 N_SUM_M1020_d N_A_84_21#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1030 N_SUM_M1020_d N_A_84_21#_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.276603 PD=1.54 PS=2.19505 NRD=0 NRS=3.5066 M=1 R=8.4 SA=75000.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1027 N_A_309_398#_M1027_d N_B_M1027_g N_VPWR_M1030_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.140497 PD=0.92 PS=1.11495 NRD=0 NRS=21.5321 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_395_398#_M1011_d N_CIN_M1011_g N_A_309_398#_M1027_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g N_A_309_398#_M1012_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.1696 PD=1 PS=1.81 NRD=24.6053 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004.6 A=0.096 P=1.58 MULT=1
MM1010 A_710_419# N_A_M1010_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1152 PD=0.85 PS=1 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.7 SB=75004.1
+ A=0.096 P=1.58 MULT=1
MM1013 A_782_419# N_B_M1013_g A_710_419# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0672 PD=0.85 PS=0.85 NRD=15.3857 NRS=15.3857 M=1 R=4.26667 SA=75001.1
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1017 N_A_84_21#_M1017_d N_CIN_M1017_g A_782_419# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0912 AS=0.0672 PD=0.925 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75001.4 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1031 N_A_941_419#_M1031_d N_A_395_398#_M1031_g N_A_84_21#_M1017_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.181325 AS=0.0912 PD=1.275 PS=0.925 NRD=36.1495 NRS=1.5366
+ M=1 R=4.26667 SA=75001.9 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_CIN_M1005_g N_A_941_419#_M1031_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.181325 PD=0.96 PS=1.275 NRD=4.6098 NRS=35.3812 M=1
+ R=4.26667 SA=75002.1 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_941_419#_M1000_d N_B_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=7.683 M=1 R=4.26667 SA=75002.6
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_A_941_419#_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.225819 AS=0.0896 PD=1.28337 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1003 N_COUT_M1003_d N_A_395_398#_M1003_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.444581 PD=1.54 PS=2.52663 NRD=0 NRS=57.0512 M=1 R=8.4
+ SA=75002.1 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1028 N_COUT_M1003_d N_A_395_398#_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.37422 PD=1.54 PS=2.50011 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.5 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1025 A_1653_367# N_A_M1025_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.19008 PD=0.85 PS=1.26989 NRD=15.3857 NRS=74.4857 M=1 R=4.26667
+ SA=75003 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_A_395_398#_M1014_d N_B_M1014_g A_1653_367# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=6.1464 NRS=15.3857 M=1 R=4.26667
+ SA=75003.4 SB=75000.2 A=0.096 P=1.58 MULT=1
DX32_noxref VNB VPB NWDIODE A=17.7175 P=22.73
*
.include "sky130_fd_sc_lp__fa_2.pxi.spice"
*
.ends
*
*
