* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_511_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_673_49# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_403_367# B1 a_511_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR A2 a_511_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_325_367# C1 a_403_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_105_239# A1 a_673_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 X a_105_239# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 X a_105_239# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_105_239# D1 a_325_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND D1 a_105_239# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_105_239# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND B1 a_105_239# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
