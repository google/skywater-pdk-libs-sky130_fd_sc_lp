* NGSPICE file created from sky130_fd_sc_lp__srsdfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__srsdfstp_1 CLK D SCD SCE SET_B SLEEP_B KAPWR VGND VNB VPB
+ VPWR Q
M1000 VPWR SCD a_27_481# VPB phighvt w=640000u l=150000u
+  ad=1.6054e+12p pd=1.277e+07u as=3.456e+11p ps=3.64e+06u
M1001 a_111_119# SCD VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.5248e+12p ps=1.521e+07u
M1002 VGND a_1068_21# a_996_73# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.694e+11p ps=1.82e+06u
M1003 VGND SET_B a_1336_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.029e+11p ps=1.33e+06u
M1004 Q a_3466_403# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.465e+11p pd=3.07e+06u as=0p ps=0u
M1005 a_887_139# a_689_139# a_189_119# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=3.283e+11p ps=3.39e+06u
M1006 a_2074_125# a_1972_99# a_2002_125# VNB nshort w=420000u l=150000u
+  ad=2.331e+11p pd=2.79e+06u as=8.82e+10p ps=1.26e+06u
M1007 VGND a_1728_125# a_3466_403# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1008 VGND SET_B a_2074_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1068_21# a_887_139# VPWR VPB phighvt w=420000u l=150000u
+  ad=2.541e+11p pd=2.47e+06u as=0p ps=0u
M1010 a_689_139# a_659_113# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1011 KAPWR a_1972_99# a_2862_414# VPB phighvt w=1e+06u l=250000u
+  ad=1.30002e+12p pd=9.18e+06u as=2.7e+11p ps=2.54e+06u
M1012 a_189_119# D a_213_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1013 a_189_119# SCE a_111_119# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1014 a_3134_72# SLEEP_B a_3056_72# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.008e+11p ps=1.32e+06u
M1015 a_3056_72# CLK a_659_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.8105e+11p ps=1.73e+06u
M1016 a_275_119# D a_189_119# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1017 a_1728_125# a_689_139# a_1656_125# VNB nshort w=640000u l=150000u
+  ad=5.339e+11p pd=3e+06u as=1.344e+11p ps=1.7e+06u
M1018 KAPWR a_1728_125# a_1972_99# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=8.55e+11p ps=3.71e+06u
M1019 VPWR a_1728_125# a_3466_403# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1020 a_3292_72# SLEEP_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1021 a_2862_414# a_689_139# a_1728_125# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.194e+11p ps=4.81e+06u
M1022 a_2216_99# SLEEP_B a_3292_72# VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1023 VGND a_339_93# a_275_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_2658_414# a_2216_99# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1025 a_1656_125# a_689_139# a_1541_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.72e+11p ps=2.13e+06u
M1026 KAPWR SLEEP_B a_659_113# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1027 VPWR SET_B a_1068_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_689_139# a_659_113# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1029 VGND SCE a_339_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1030 a_1712_451# a_659_113# a_1541_125# VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=5.922e+11p ps=3.09e+06u
M1031 a_996_73# a_689_139# a_887_139# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.2695e+11p ps=2.29e+06u
M1032 a_1541_125# a_887_139# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q a_3466_403# VGND VNB nshort w=840000u l=150000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1034 a_1132_535# a_659_113# a_887_139# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1035 VPWR a_1068_21# a_1132_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR SCE a_339_93# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1037 a_1728_125# a_659_113# a_1712_451# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1336_97# a_887_139# a_1068_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1039 a_659_113# CLK KAPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1541_125# a_887_139# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1972_99# a_1728_125# a_2463_119# VNB nshort w=420000u l=150000u
+  ad=2.282e+11p pd=2.08e+06u as=8.82e+10p ps=1.26e+06u
M1042 a_213_481# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1728_125# SET_B a_2658_414# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_2074_125# a_2216_99# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_2216_99# SLEEP_B KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1046 a_2002_125# a_1972_99# a_1930_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1047 a_887_139# a_659_113# a_189_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_27_481# a_339_93# a_189_119# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND SLEEP_B a_3134_72# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_1930_125# a_659_113# a_1728_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_2463_119# a_1728_125# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

