* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
X0 a_470_367# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND a_1418_21# a_110_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 Y A1 a_470_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR a_1418_21# a_470_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND S a_470_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_470_69# S VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_126_367# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_110_69# A0 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 Y A1 a_470_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_110_69# a_1418_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 Y A0 a_110_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND S a_1418_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_470_367# a_1418_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_110_69# A0 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y A0 a_126_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y A1 a_470_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_470_367# a_1418_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR a_1418_21# a_470_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_470_69# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VGND a_1418_21# a_110_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 Y A0 a_126_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_126_367# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_110_69# a_1418_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_126_367# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VPWR S a_126_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_470_69# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 Y A1 a_470_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 Y A0 a_110_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_470_367# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 VPWR S a_126_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_126_367# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 VGND S a_470_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 VPWR S a_1418_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_470_69# S VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
