* File: sky130_fd_sc_lp__o211ai_0.pxi.spice
* Created: Wed Sep  2 10:14:22 2020
* 
x_PM_SKY130_FD_SC_LP__O211AI_0%A1 N_A1_c_58_n N_A1_M1004_g N_A1_M1002_g
+ N_A1_c_60_n N_A1_c_61_n A1 A1 N_A1_c_62_n PM_SKY130_FD_SC_LP__O211AI_0%A1
x_PM_SKY130_FD_SC_LP__O211AI_0%A2 N_A2_c_92_n N_A2_M1000_g N_A2_c_93_n
+ N_A2_M1007_g N_A2_c_94_n N_A2_c_95_n A2 A2 N_A2_c_97_n N_A2_c_98_n
+ PM_SKY130_FD_SC_LP__O211AI_0%A2
x_PM_SKY130_FD_SC_LP__O211AI_0%B1 N_B1_c_145_n N_B1_M1005_g N_B1_c_146_n
+ N_B1_M1003_g N_B1_c_147_n N_B1_c_142_n N_B1_c_149_n B1 B1 N_B1_c_144_n
+ PM_SKY130_FD_SC_LP__O211AI_0%B1
x_PM_SKY130_FD_SC_LP__O211AI_0%C1 N_C1_M1001_g N_C1_c_193_n N_C1_M1006_g C1 C1
+ C1 PM_SKY130_FD_SC_LP__O211AI_0%C1
x_PM_SKY130_FD_SC_LP__O211AI_0%VPWR N_VPWR_M1002_s N_VPWR_M1005_d N_VPWR_c_221_n
+ N_VPWR_c_222_n N_VPWR_c_223_n VPWR N_VPWR_c_224_n N_VPWR_c_225_n
+ N_VPWR_c_220_n N_VPWR_c_227_n PM_SKY130_FD_SC_LP__O211AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O211AI_0%Y N_Y_M1001_d N_Y_M1000_d N_Y_M1006_d N_Y_c_254_n
+ N_Y_c_255_n N_Y_c_252_n Y Y Y Y Y N_Y_c_258_n PM_SKY130_FD_SC_LP__O211AI_0%Y
x_PM_SKY130_FD_SC_LP__O211AI_0%A_36_47# N_A_36_47#_M1004_s N_A_36_47#_M1007_d
+ N_A_36_47#_c_299_n N_A_36_47#_c_300_n N_A_36_47#_c_301_n N_A_36_47#_c_302_n
+ PM_SKY130_FD_SC_LP__O211AI_0%A_36_47#
x_PM_SKY130_FD_SC_LP__O211AI_0%VGND N_VGND_M1004_d VGND N_VGND_c_333_n
+ N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n PM_SKY130_FD_SC_LP__O211AI_0%VGND
cc_1 VNB N_A1_c_58_n 0.0344456f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.915
cc_2 VNB N_A1_M1004_g 0.0313959f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.445
cc_3 VNB N_A1_c_60_n 0.0271175f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.585
cc_4 VNB N_A1_c_61_n 0.00561606f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.75
cc_5 VNB N_A1_c_62_n 0.0288046f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_6 VNB N_A2_c_92_n 0.0204783f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.445
cc_7 VNB N_A2_c_93_n 0.0187175f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_8 VNB N_A2_c_94_n 6.64879e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A2_c_95_n 0.0194222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A2 0.00624538f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_11 VNB N_A2_c_97_n 0.0179605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_98_n 0.0140514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1003_g 0.0349648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_142_n 0.0216264f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_15 VNB B1 0.00755075f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_16 VNB N_B1_c_144_n 0.0157492f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.665
cc_17 VNB N_C1_M1001_g 0.0241273f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.445
cc_18 VNB N_C1_c_193_n 0.101884f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.75
cc_19 VNB N_C1_M1006_g 0.00828029f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.645
cc_20 VNB C1 0.0414111f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_21 VNB N_VPWR_c_220_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_252_n 0.0139405f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_23 VNB Y 0.00905166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_36_47#_c_299_n 0.0186284f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.245
cc_25 VNB N_A_36_47#_c_300_n 0.0216299f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.75
cc_26 VNB N_A_36_47#_c_301_n 0.00984039f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_A_36_47#_c_302_n 7.92356e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_333_n 0.0463179f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_VGND_c_334_n 0.174538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_335_n 0.0162959f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.245
cc_31 VNB N_VGND_c_336_n 0.0123937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_A1_M1002_g 0.0560772f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.645
cc_33 VPB N_A1_c_61_n 0.0127594f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.75
cc_34 VPB N_A1_c_62_n 0.0170586f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_35 VPB N_A2_M1000_g 0.0363722f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.75
cc_36 VPB N_A2_c_94_n 0.0171387f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_37 VPB A2 0.00122413f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_38 VPB N_B1_c_145_n 0.0201759f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=0.915
cc_39 VPB N_B1_c_146_n 0.013944f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.75
cc_40 VPB N_B1_c_147_n 0.0202884f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_41 VPB N_B1_c_142_n 5.91602e-19 $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_42 VPB N_B1_c_149_n 0.0157918f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_43 VPB B1 0.00119541f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_44 VPB N_C1_M1006_g 0.0578994f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.645
cc_45 VPB C1 0.0105342f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_46 VPB N_VPWR_c_221_n 0.0146748f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.645
cc_47 VPB N_VPWR_c_222_n 0.0390517f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_48 VPB N_VPWR_c_223_n 0.0175814f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_49 VPB N_VPWR_c_224_n 0.0269762f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.245
cc_50 VPB N_VPWR_c_225_n 0.0239584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_220_n 0.0644373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_227_n 0.0113226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_Y_c_254_n 0.00197461f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.585
cc_54 VPB N_Y_c_255_n 0.00428965f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_55 VPB Y 0.0268324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB Y 0.0514376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_258_n 0.0174978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 N_A1_c_60_n N_A2_c_92_n 0.0292735f $X=0.49 $Y=1.585 $X2=0 $Y2=0
cc_59 N_A1_M1002_g N_A2_M1000_g 0.0292735f $X=0.58 $Y=2.645 $X2=0 $Y2=0
cc_60 N_A1_M1004_g N_A2_c_93_n 0.0046625f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_61 N_A1_c_61_n N_A2_c_94_n 0.0292735f $X=0.49 $Y=1.75 $X2=0 $Y2=0
cc_62 N_A1_c_58_n N_A2_c_95_n 0.00776863f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_63 N_A1_M1004_g N_A2_c_95_n 0.00305918f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_64 N_A1_c_58_n A2 0.00276853f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_65 N_A1_c_62_n A2 0.0319291f $X=0.49 $Y=1.245 $X2=0 $Y2=0
cc_66 N_A1_c_58_n N_A2_c_97_n 0.0292735f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_67 N_A1_c_62_n N_A2_c_97_n 0.00246911f $X=0.49 $Y=1.245 $X2=0 $Y2=0
cc_68 N_A1_M1002_g N_VPWR_c_222_n 0.0168604f $X=0.58 $Y=2.645 $X2=0 $Y2=0
cc_69 N_A1_c_61_n N_VPWR_c_222_n 0.00103504f $X=0.49 $Y=1.75 $X2=0 $Y2=0
cc_70 N_A1_c_62_n N_VPWR_c_222_n 0.0152575f $X=0.49 $Y=1.245 $X2=0 $Y2=0
cc_71 N_A1_M1002_g N_VPWR_c_224_n 0.00386543f $X=0.58 $Y=2.645 $X2=0 $Y2=0
cc_72 N_A1_M1002_g N_VPWR_c_220_n 0.0076021f $X=0.58 $Y=2.645 $X2=0 $Y2=0
cc_73 N_A1_M1002_g N_Y_c_254_n 9.1846e-19 $X=0.58 $Y=2.645 $X2=0 $Y2=0
cc_74 N_A1_M1002_g N_Y_c_255_n 0.00270302f $X=0.58 $Y=2.645 $X2=0 $Y2=0
cc_75 N_A1_M1004_g N_A_36_47#_c_299_n 0.00375589f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A1_c_58_n N_A_36_47#_c_300_n 0.00329468f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_77 N_A1_M1004_g N_A_36_47#_c_300_n 0.0149092f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_78 N_A1_c_62_n N_A_36_47#_c_300_n 0.013385f $X=0.49 $Y=1.245 $X2=0 $Y2=0
cc_79 N_A1_c_58_n N_A_36_47#_c_301_n 5.8044e-19 $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_80 N_A1_c_62_n N_A_36_47#_c_301_n 0.0238827f $X=0.49 $Y=1.245 $X2=0 $Y2=0
cc_81 N_A1_M1004_g N_VGND_c_334_n 0.0054391f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A1_M1004_g N_VGND_c_335_n 0.00365758f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A1_M1004_g N_VGND_c_336_n 0.0114124f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A2_c_93_n N_B1_M1003_g 0.0194252f $X=1.29 $Y=0.77 $X2=0 $Y2=0
cc_85 A2 N_B1_M1003_g 2.11463e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A2_c_98_n N_B1_M1003_g 0.00763927f $X=1.045 $Y=1.155 $X2=0 $Y2=0
cc_87 N_A2_M1000_g N_B1_c_147_n 0.0168071f $X=0.94 $Y=2.645 $X2=0 $Y2=0
cc_88 N_A2_c_92_n N_B1_c_142_n 0.0119167f $X=1.045 $Y=1.645 $X2=0 $Y2=0
cc_89 N_A2_M1000_g N_B1_c_149_n 0.0067428f $X=0.94 $Y=2.645 $X2=0 $Y2=0
cc_90 N_A2_c_94_n N_B1_c_149_n 0.0119167f $X=1.045 $Y=1.825 $X2=0 $Y2=0
cc_91 N_A2_c_94_n B1 2.10841e-19 $X=1.045 $Y=1.825 $X2=0 $Y2=0
cc_92 A2 B1 0.0546014f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A2_c_97_n B1 6.49174e-19 $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_94 N_A2_c_98_n B1 2.67888e-19 $X=1.045 $Y=1.155 $X2=0 $Y2=0
cc_95 A2 N_B1_c_144_n 0.0036216f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A2_c_97_n N_B1_c_144_n 0.0119167f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_97 N_A2_M1000_g N_VPWR_c_222_n 0.00243681f $X=0.94 $Y=2.645 $X2=0 $Y2=0
cc_98 N_A2_M1000_g N_VPWR_c_224_n 0.00438034f $X=0.94 $Y=2.645 $X2=0 $Y2=0
cc_99 N_A2_M1000_g N_VPWR_c_220_n 0.00829237f $X=0.94 $Y=2.645 $X2=0 $Y2=0
cc_100 N_A2_M1000_g N_Y_c_254_n 0.00658702f $X=0.94 $Y=2.645 $X2=0 $Y2=0
cc_101 N_A2_c_94_n N_Y_c_254_n 0.00611986f $X=1.045 $Y=1.825 $X2=0 $Y2=0
cc_102 A2 N_Y_c_254_n 0.0238075f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A2_M1000_g N_Y_c_255_n 0.0160361f $X=0.94 $Y=2.645 $X2=0 $Y2=0
cc_104 N_A2_c_93_n N_A_36_47#_c_300_n 0.0048244f $X=1.29 $Y=0.77 $X2=0 $Y2=0
cc_105 N_A2_c_95_n N_A_36_47#_c_300_n 0.0148684f $X=1.29 $Y=0.845 $X2=0 $Y2=0
cc_106 A2 N_A_36_47#_c_300_n 0.0320702f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A2_c_97_n N_A_36_47#_c_300_n 0.00220741f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_108 N_A2_c_93_n N_A_36_47#_c_302_n 0.00224886f $X=1.29 $Y=0.77 $X2=0 $Y2=0
cc_109 N_A2_c_93_n N_VGND_c_333_n 0.00365758f $X=1.29 $Y=0.77 $X2=0 $Y2=0
cc_110 N_A2_c_93_n N_VGND_c_334_n 0.00441909f $X=1.29 $Y=0.77 $X2=0 $Y2=0
cc_111 N_A2_c_93_n N_VGND_c_336_n 0.0103009f $X=1.29 $Y=0.77 $X2=0 $Y2=0
cc_112 N_A2_c_95_n N_VGND_c_336_n 8.40465e-19 $X=1.29 $Y=0.845 $X2=0 $Y2=0
cc_113 N_B1_M1003_g N_C1_M1001_g 0.0345446f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_114 B1 N_C1_c_193_n 0.00266976f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B1_c_144_n N_C1_c_193_n 0.0485846f $X=1.63 $Y=1.325 $X2=0 $Y2=0
cc_116 N_B1_c_145_n N_C1_M1006_g 0.00375989f $X=1.37 $Y=2.215 $X2=0 $Y2=0
cc_117 N_B1_c_146_n N_C1_M1006_g 0.00924478f $X=1.54 $Y=2.065 $X2=0 $Y2=0
cc_118 N_B1_c_142_n N_C1_M1006_g 0.01404f $X=1.63 $Y=1.665 $X2=0 $Y2=0
cc_119 N_B1_c_145_n N_VPWR_c_223_n 0.00439863f $X=1.37 $Y=2.215 $X2=0 $Y2=0
cc_120 N_B1_c_147_n N_VPWR_c_223_n 0.00458496f $X=1.54 $Y=2.14 $X2=0 $Y2=0
cc_121 N_B1_c_145_n N_VPWR_c_224_n 0.00465548f $X=1.37 $Y=2.215 $X2=0 $Y2=0
cc_122 N_B1_c_145_n N_VPWR_c_220_n 0.00919736f $X=1.37 $Y=2.215 $X2=0 $Y2=0
cc_123 N_B1_c_147_n N_Y_c_255_n 0.00518245f $X=1.54 $Y=2.14 $X2=0 $Y2=0
cc_124 N_B1_M1003_g N_Y_c_252_n 0.0011034f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_125 N_B1_c_146_n Y 0.00210604f $X=1.54 $Y=2.065 $X2=0 $Y2=0
cc_126 N_B1_M1003_g Y 0.00228375f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_127 N_B1_c_149_n Y 0.00104456f $X=1.63 $Y=1.83 $X2=0 $Y2=0
cc_128 B1 Y 0.0563126f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B1_c_144_n Y 0.00157111f $X=1.63 $Y=1.325 $X2=0 $Y2=0
cc_130 N_B1_c_146_n N_Y_c_258_n 0.00736809f $X=1.54 $Y=2.065 $X2=0 $Y2=0
cc_131 N_B1_c_147_n N_Y_c_258_n 0.0152855f $X=1.54 $Y=2.14 $X2=0 $Y2=0
cc_132 N_B1_c_149_n N_Y_c_258_n 0.00502306f $X=1.63 $Y=1.83 $X2=0 $Y2=0
cc_133 B1 N_Y_c_258_n 0.0296966f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B1_M1003_g N_A_36_47#_c_300_n 0.00467555f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_135 B1 N_A_36_47#_c_300_n 0.01882f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B1_c_144_n N_A_36_47#_c_300_n 0.0011256f $X=1.63 $Y=1.325 $X2=0 $Y2=0
cc_137 N_B1_M1003_g N_A_36_47#_c_302_n 0.00738847f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_138 N_B1_M1003_g N_VGND_c_333_n 0.0054978f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_139 N_B1_M1003_g N_VGND_c_334_n 0.00995168f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_140 N_B1_M1003_g N_VGND_c_336_n 0.00124576f $X=1.72 $Y=0.445 $X2=0 $Y2=0
cc_141 N_C1_M1006_g N_VPWR_c_223_n 0.00439863f $X=2.14 $Y=2.645 $X2=0 $Y2=0
cc_142 N_C1_M1006_g N_VPWR_c_225_n 0.00465548f $X=2.14 $Y=2.645 $X2=0 $Y2=0
cc_143 N_C1_M1006_g N_VPWR_c_220_n 0.00928042f $X=2.14 $Y=2.645 $X2=0 $Y2=0
cc_144 N_C1_M1001_g N_Y_c_252_n 0.0090404f $X=2.08 $Y=0.445 $X2=0 $Y2=0
cc_145 N_C1_c_193_n N_Y_c_252_n 0.00818614f $X=2.14 $Y=1.51 $X2=0 $Y2=0
cc_146 C1 N_Y_c_252_n 0.00502908f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_147 N_C1_M1001_g Y 0.00877248f $X=2.08 $Y=0.445 $X2=0 $Y2=0
cc_148 N_C1_c_193_n Y 0.0359378f $X=2.14 $Y=1.51 $X2=0 $Y2=0
cc_149 N_C1_M1006_g Y 0.0323648f $X=2.14 $Y=2.645 $X2=0 $Y2=0
cc_150 C1 Y 0.109398f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_151 N_C1_M1006_g Y 0.00905102f $X=2.14 $Y=2.645 $X2=0 $Y2=0
cc_152 N_C1_M1001_g N_A_36_47#_c_300_n 4.78309e-19 $X=2.08 $Y=0.445 $X2=0 $Y2=0
cc_153 N_C1_M1001_g N_A_36_47#_c_302_n 0.00116829f $X=2.08 $Y=0.445 $X2=0 $Y2=0
cc_154 N_C1_M1001_g N_VGND_c_333_n 0.0037047f $X=2.08 $Y=0.445 $X2=0 $Y2=0
cc_155 N_C1_M1001_g N_VGND_c_334_n 0.00683579f $X=2.08 $Y=0.445 $X2=0 $Y2=0
cc_156 C1 N_VGND_c_334_n 0.0139442f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_157 N_VPWR_c_222_n N_Y_c_255_n 0.0225862f $X=0.365 $Y=2.47 $X2=0 $Y2=0
cc_158 N_VPWR_c_223_n N_Y_c_255_n 0.00328429f $X=1.925 $Y=2.47 $X2=0 $Y2=0
cc_159 N_VPWR_c_224_n N_Y_c_255_n 0.0134967f $X=1.46 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_220_n N_Y_c_255_n 0.0109236f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_161 N_VPWR_c_223_n Y 0.00360736f $X=1.925 $Y=2.47 $X2=0 $Y2=0
cc_162 N_VPWR_c_223_n Y 0.00344526f $X=1.925 $Y=2.47 $X2=0 $Y2=0
cc_163 N_VPWR_c_225_n Y 0.0260909f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_c_220_n Y 0.0212262f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_c_223_n N_Y_c_258_n 0.0460092f $X=1.925 $Y=2.47 $X2=0 $Y2=0
cc_166 Y N_A_36_47#_c_300_n 0.00750115f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_167 N_Y_c_252_n N_A_36_47#_c_302_n 0.0144673f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_168 Y N_A_36_47#_c_302_n 0.00508407f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_169 N_Y_c_252_n N_VGND_c_333_n 0.0240041f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_170 N_Y_M1001_d N_VGND_c_334_n 0.0021695f $X=2.155 $Y=0.235 $X2=0 $Y2=0
cc_171 N_Y_c_252_n N_VGND_c_334_n 0.0162595f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_172 N_A_36_47#_c_300_n N_VGND_c_333_n 0.00226785f $X=1.41 $Y=0.825 $X2=0
+ $Y2=0
cc_173 N_A_36_47#_c_302_n N_VGND_c_333_n 0.0134701f $X=1.505 $Y=0.445 $X2=0
+ $Y2=0
cc_174 N_A_36_47#_M1004_s N_VGND_c_334_n 0.00239031f $X=0.18 $Y=0.235 $X2=0
+ $Y2=0
cc_175 N_A_36_47#_M1007_d N_VGND_c_334_n 0.00248289f $X=1.365 $Y=0.235 $X2=0
+ $Y2=0
cc_176 N_A_36_47#_c_299_n N_VGND_c_334_n 0.00988702f $X=0.305 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_36_47#_c_300_n N_VGND_c_334_n 0.0101907f $X=1.41 $Y=0.825 $X2=0 $Y2=0
cc_178 N_A_36_47#_c_302_n N_VGND_c_334_n 0.0097649f $X=1.505 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_36_47#_c_299_n N_VGND_c_335_n 0.0152657f $X=0.305 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_36_47#_c_300_n N_VGND_c_335_n 0.00226785f $X=1.41 $Y=0.825 $X2=0
+ $Y2=0
cc_181 N_A_36_47#_c_300_n N_VGND_c_336_n 0.0477084f $X=1.41 $Y=0.825 $X2=0 $Y2=0
cc_182 N_VGND_c_334_n A_359_47# 0.00899413f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
