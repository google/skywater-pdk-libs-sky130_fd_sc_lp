* File: sky130_fd_sc_lp__xnor2_2.pex.spice
* Created: Fri Aug 28 11:35:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR2_2%A 3 7 11 15 19 23 27 31 34 35 36 38 39 41 44
+ 45 53 61 63
c142 61 0 1.88077e-19 $X=3.545 $Y=1.49
c143 53 0 1.00558e-19 $X=1.185 $Y=1.51
c144 41 0 5.16709e-20 $X=2.97 $Y=1.49
c145 39 0 1.97098e-19 $X=2.635 $Y=1.49
c146 38 0 7.0048e-20 $X=2.55 $Y=1.405
c147 23 0 1.91591e-19 $X=3.08 $Y=2.465
r148 60 61 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.115 $Y=1.49
+ $X2=3.545 $Y2=1.49
r149 59 60 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.08 $Y=1.49
+ $X2=3.115 $Y2=1.49
r150 53 55 3.44286 $w=2.8e-07 $l=2e-08 $layer=POLY_cond $X=1.185 $Y=1.51
+ $X2=1.205 $Y2=1.51
r151 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.185
+ $Y=1.51 $X2=1.185 $Y2=1.51
r152 51 53 3.44286 $w=2.8e-07 $l=2e-08 $layer=POLY_cond $X=1.165 $Y=1.51
+ $X2=1.185 $Y2=1.51
r153 50 51 74.0214 $w=2.8e-07 $l=4.3e-07 $layer=POLY_cond $X=0.735 $Y=1.51
+ $X2=1.165 $Y2=1.51
r154 45 63 2.65806 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=1.587
+ $X2=1.655 $Y2=1.587
r155 45 63 1.06379 $w=3.23e-07 $l=3e-08 $layer=LI1_cond $X=1.625 $Y=1.587
+ $X2=1.655 $Y2=1.587
r156 44 45 15.0704 $w=3.23e-07 $l=4.25e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.625 $Y2=1.587
r157 44 54 0.531897 $w=3.23e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.185 $Y2=1.587
r158 42 59 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.97 $Y=1.49
+ $X2=3.08 $Y2=1.49
r159 42 56 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=2.97 $Y=1.49
+ $X2=2.65 $Y2=1.49
r160 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.97
+ $Y=1.49 $X2=2.97 $Y2=1.49
r161 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.635 $Y=1.49
+ $X2=2.97 $Y2=1.49
r162 38 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.55 $Y=1.405
+ $X2=2.635 $Y2=1.49
r163 37 38 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.55 $Y=1.175
+ $X2=2.55 $Y2=1.405
r164 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.465 $Y=1.09
+ $X2=2.55 $Y2=1.175
r165 35 36 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.465 $Y=1.09
+ $X2=1.825 $Y2=1.09
r166 34 45 5.06595 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=1.74 $Y=1.425
+ $X2=1.74 $Y2=1.587
r167 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.74 $Y=1.175
+ $X2=1.825 $Y2=1.09
r168 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.74 $Y=1.175
+ $X2=1.74 $Y2=1.425
r169 29 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=1.325
+ $X2=3.545 $Y2=1.49
r170 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.545 $Y=1.325
+ $X2=3.545 $Y2=0.745
r171 25 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.325
+ $X2=3.115 $Y2=1.49
r172 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.115 $Y=1.325
+ $X2=3.115 $Y2=0.745
r173 21 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.655
+ $X2=3.08 $Y2=1.49
r174 21 23 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.08 $Y=1.655
+ $X2=3.08 $Y2=2.465
r175 17 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.655
+ $X2=2.65 $Y2=1.49
r176 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.65 $Y=1.655
+ $X2=2.65 $Y2=2.465
r177 13 55 17.3521 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.345
+ $X2=1.205 $Y2=1.51
r178 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.205 $Y=1.345
+ $X2=1.205 $Y2=0.655
r179 9 51 17.3521 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.675
+ $X2=1.165 $Y2=1.51
r180 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.165 $Y=1.675
+ $X2=1.165 $Y2=2.465
r181 5 50 17.3521 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.675
+ $X2=0.735 $Y2=1.51
r182 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.735 $Y=1.675
+ $X2=0.735 $Y2=2.465
r183 1 50 44.7571 $w=2.8e-07 $l=3.32415e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.735 $Y2=1.51
r184 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%B 3 7 11 15 19 23 27 31 33 34 37 42 43 46 47
+ 48 49 54
c142 54 0 7.61574e-20 $X=4.335 $Y=1.51
c143 43 0 4.63394e-19 $X=2.09 $Y=1.51
c144 42 0 1.00558e-19 $X=2.09 $Y=1.51
c145 33 0 3.89867e-19 $X=4.05 $Y=1.51
c146 31 0 8.77403e-20 $X=4.905 $Y=2.465
c147 27 0 7.76303e-20 $X=4.835 $Y=0.745
c148 3 0 8.28055e-20 $X=1.635 $Y=0.655
r149 55 57 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.635 $Y=1.51
+ $X2=2.065 $Y2=1.51
r150 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.335
+ $Y=1.51 $X2=4.335 $Y2=1.51
r151 49 54 8.51806 $w=3.43e-07 $l=2.55e-07 $layer=LI1_cond $X=4.08 $Y=1.577
+ $X2=4.335 $Y2=1.577
r152 48 49 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.577
+ $X2=4.08 $Y2=1.577
r153 47 48 4.17552 $w=3.43e-07 $l=1.25e-07 $layer=LI1_cond $X=3.475 $Y=1.577
+ $X2=3.6 $Y2=1.577
r154 46 47 8.64642 $w=3.43e-07 $l=1.7e-07 $layer=LI1_cond $X=3.305 $Y=1.66
+ $X2=3.475 $Y2=1.66
r155 43 57 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.09 $Y=1.51
+ $X2=2.065 $Y2=1.51
r156 42 44 16.3347 $w=2.39e-07 $l=3.2e-07 $layer=LI1_cond $X=2.14 $Y=1.51
+ $X2=2.14 $Y2=1.83
r157 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.51 $X2=2.09 $Y2=1.51
r158 40 44 2.73298 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.285 $Y=1.83
+ $X2=2.14 $Y2=1.83
r159 40 46 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.285 $Y=1.83
+ $X2=3.305 $Y2=1.83
r160 36 37 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.835 $Y=1.51
+ $X2=4.905 $Y2=1.51
r161 35 36 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.475 $Y=1.51
+ $X2=4.835 $Y2=1.51
r162 34 53 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=4.4 $Y=1.51
+ $X2=4.335 $Y2=1.51
r163 34 35 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.4 $Y=1.51
+ $X2=4.475 $Y2=1.51
r164 33 53 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=4.05 $Y=1.51
+ $X2=4.335 $Y2=1.51
r165 29 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.675
+ $X2=4.905 $Y2=1.51
r166 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.905 $Y=1.675
+ $X2=4.905 $Y2=2.465
r167 25 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.345
+ $X2=4.835 $Y2=1.51
r168 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.835 $Y=1.345
+ $X2=4.835 $Y2=0.745
r169 21 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.475 $Y=1.675
+ $X2=4.475 $Y2=1.51
r170 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.475 $Y=1.675
+ $X2=4.475 $Y2=2.465
r171 17 33 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.975 $Y=1.345
+ $X2=4.05 $Y2=1.51
r172 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.975 $Y=1.345
+ $X2=3.975 $Y2=0.745
r173 13 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.675
+ $X2=2.065 $Y2=1.51
r174 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.065 $Y=1.675
+ $X2=2.065 $Y2=2.465
r175 9 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.345
+ $X2=2.065 $Y2=1.51
r176 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.065 $Y=1.345
+ $X2=2.065 $Y2=0.655
r177 5 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.675
+ $X2=1.635 $Y2=1.51
r178 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.635 $Y=1.675
+ $X2=1.635 $Y2=2.465
r179 1 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.345
+ $X2=1.635 $Y2=1.51
r180 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.635 $Y=1.345
+ $X2=1.635 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%A_162_367# 1 2 3 12 16 20 24 27 30 32 33 34
+ 37 38 40 42 44 46 48 51 52 54 58 63 72
c147 72 0 7.61574e-20 $X=5.765 $Y=1.51
c148 63 0 1.46605e-19 $X=3.75 $Y=2.005
c149 40 0 1.96248e-19 $X=1.85 $Y=0.71
r150 71 72 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.695 $Y=1.51
+ $X2=5.765 $Y2=1.51
r151 67 69 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.265 $Y=1.51
+ $X2=5.335 $Y2=1.51
r152 63 65 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.75 $Y=2.005
+ $X2=3.75 $Y2=2.17
r153 61 62 4.41277 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=2.085
+ $X2=1.88 $Y2=2.17
r154 59 61 4.15319 $w=2.35e-07 $l=8e-08 $layer=LI1_cond $X=1.88 $Y=2.005
+ $X2=1.88 $Y2=2.085
r155 55 71 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=5.55 $Y=1.51
+ $X2=5.695 $Y2=1.51
r156 55 69 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.55 $Y=1.51
+ $X2=5.335 $Y2=1.51
r157 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=1.51 $X2=5.55 $Y2=1.51
r158 52 54 38.5409 $w=1.98e-07 $l=6.95e-07 $layer=LI1_cond $X=4.855 $Y=1.505
+ $X2=5.55 $Y2=1.505
r159 50 52 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.77 $Y=1.605
+ $X2=4.855 $Y2=1.505
r160 50 51 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.77 $Y=1.605
+ $X2=4.77 $Y2=1.92
r161 49 63 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.855 $Y=2.005
+ $X2=3.75 $Y2=2.005
r162 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.685 $Y=2.005
+ $X2=4.77 $Y2=1.92
r163 48 49 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.685 $Y=2.005
+ $X2=3.855 $Y2=2.005
r164 47 62 2.6346 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.015 $Y=2.17
+ $X2=1.88 $Y2=2.17
r165 46 65 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.645 $Y=2.17
+ $X2=3.75 $Y2=2.17
r166 46 47 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=3.645 $Y=2.17
+ $X2=2.015 $Y2=2.17
r167 42 62 4.07826 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=2.255
+ $X2=1.88 $Y2=2.17
r168 42 44 27.9574 $w=2.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.88 $Y=2.255
+ $X2=1.88 $Y2=2.91
r169 38 40 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.485 $Y=0.715
+ $X2=1.85 $Y2=0.715
r170 36 38 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.4 $Y=0.815
+ $X2=1.485 $Y2=0.715
r171 36 37 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.4 $Y=0.815
+ $X2=1.4 $Y2=1.075
r172 35 58 2.11342 $w=1.7e-07 $l=1.95484e-07 $layer=LI1_cond $X=1.065 $Y=2.005
+ $X2=0.872 $Y2=2.01
r173 34 59 2.6346 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=2.005
+ $X2=1.88 $Y2=2.005
r174 34 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.745 $Y=2.005
+ $X2=1.065 $Y2=2.005
r175 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.315 $Y=1.16
+ $X2=1.4 $Y2=1.075
r176 32 33 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.315 $Y=1.16
+ $X2=0.85 $Y2=1.16
r177 28 58 4.3182 $w=2.1e-07 $l=1.19248e-07 $layer=LI1_cond $X=0.94 $Y=2.1
+ $X2=0.872 $Y2=2.01
r178 28 30 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=0.94 $Y=2.1
+ $X2=0.94 $Y2=2.475
r179 27 58 4.3182 $w=2.1e-07 $l=1.45186e-07 $layer=LI1_cond $X=0.765 $Y=1.92
+ $X2=0.872 $Y2=2.01
r180 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.765 $Y=1.245
+ $X2=0.85 $Y2=1.16
r181 26 27 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.765 $Y=1.245
+ $X2=0.765 $Y2=1.92
r182 22 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=1.675
+ $X2=5.765 $Y2=1.51
r183 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.765 $Y=1.675
+ $X2=5.765 $Y2=2.465
r184 18 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.345
+ $X2=5.695 $Y2=1.51
r185 18 20 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.695 $Y=1.345
+ $X2=5.695 $Y2=0.745
r186 14 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.335 $Y=1.675
+ $X2=5.335 $Y2=1.51
r187 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.335 $Y=1.675
+ $X2=5.335 $Y2=2.465
r188 10 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.345
+ $X2=5.265 $Y2=1.51
r189 10 12 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.265 $Y=1.345
+ $X2=5.265 $Y2=0.745
r190 3 61 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.835 $X2=1.85 $Y2=2.085
r191 3 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.835 $X2=1.85 $Y2=2.91
r192 2 58 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=0.81
+ $Y=1.835 $X2=0.95 $Y2=2.015
r193 2 30 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=0.81
+ $Y=1.835 $X2=0.95 $Y2=2.475
r194 1 40 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=1.71
+ $Y=0.235 $X2=1.85 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%VPWR 1 2 3 4 5 18 23 26 30 34 38 44 45 47 48
+ 50 51 53 54 55 69 78 79 82 90
r95 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r96 79 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r97 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r98 76 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=3.33
+ $X2=5.55 $Y2=3.33
r99 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.715 $Y=3.33 $X2=6
+ $Y2=3.33
r100 75 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r101 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r102 72 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 72 90 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.36 $Y2=3.33
r104 71 74 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r105 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r106 69 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=5.55 $Y2=3.33
r107 69 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 55 90 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.36 $Y2=3.33
r114 55 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 55 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 53 67 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.2 $Y=3.33 $X2=3.12
+ $Y2=3.33
r117 53 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.2 $Y=3.33 $X2=3.33
+ $Y2=3.33
r118 52 71 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 52 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.33 $Y2=3.33
r120 50 64 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.36 $Y2=3.33
r122 49 67 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=3.12 $Y2=3.33
r123 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.36 $Y2=3.33
r124 47 61 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=1.4 $Y2=3.33
r126 46 64 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.4 $Y2=3.33
r128 44 58 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=3.33 $X2=0.24
+ $Y2=3.33
r129 44 45 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=0.3 $Y=3.33
+ $X2=0.472 $Y2=3.33
r130 43 61 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 43 45 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.472 $Y2=3.33
r132 38 41 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=5.55 $Y=2.2
+ $X2=5.55 $Y2=2.97
r133 36 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=3.245
+ $X2=5.55 $Y2=3.33
r134 36 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.55 $Y=3.245
+ $X2=5.55 $Y2=2.97
r135 32 54 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=3.33
r136 32 34 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=2.94
r137 28 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=3.245
+ $X2=2.36 $Y2=3.33
r138 28 30 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=2.36 $Y=3.245
+ $X2=2.36 $Y2=2.54
r139 24 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=3.245 $X2=1.4
+ $Y2=3.33
r140 24 26 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=1.4 $Y=3.245
+ $X2=1.4 $Y2=2.385
r141 21 45 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.472 $Y=3.245
+ $X2=0.472 $Y2=3.33
r142 21 23 26.0552 $w=3.43e-07 $l=7.8e-07 $layer=LI1_cond $X=0.472 $Y=3.245
+ $X2=0.472 $Y2=2.465
r143 20 42 7.49751 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=0.472 $Y=2.442
+ $X2=0.472 $Y2=2.27
r144 20 23 0.768295 $w=3.43e-07 $l=2.3e-08 $layer=LI1_cond $X=0.472 $Y=2.442
+ $X2=0.472 $Y2=2.465
r145 18 42 15.316 $w=2.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.405 $Y=1.98
+ $X2=0.405 $Y2=2.27
r146 5 41 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.835 $X2=5.55 $Y2=2.97
r147 5 38 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.835 $X2=5.55 $Y2=2.2
r148 4 34 600 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=1.835 $X2=3.295 $Y2=2.94
r149 3 30 300 $w=1.7e-07 $l=8.07543e-07 $layer=licon1_PDIFF $count=2 $X=2.14
+ $Y=1.835 $X2=2.36 $Y2=2.54
r150 2 26 300 $w=1.7e-07 $l=6.249e-07 $layer=licon1_PDIFF $count=2 $X=1.24
+ $Y=1.835 $X2=1.4 $Y2=2.385
r151 1 23 300 $w=1.7e-07 $l=7.40338e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=1.835 $X2=0.52 $Y2=2.465
r152 1 18 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.28
+ $Y=1.835 $X2=0.425 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%A_545_367# 1 2 9 12 13 14 16 18
c43 13 0 8.77403e-20 $X=4.525 $Y=2.98
r44 18 20 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.69 $Y=2.725
+ $X2=4.69 $Y2=2.98
r45 13 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=2.98
+ $X2=4.69 $Y2=2.98
r46 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.525 $Y=2.98
+ $X2=3.855 $Y2=2.98
r47 12 14 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.742 $Y=2.895
+ $X2=3.855 $Y2=2.98
r48 11 12 14.8537 $w=2.23e-07 $l=2.9e-07 $layer=LI1_cond $X=3.742 $Y=2.605
+ $X2=3.742 $Y2=2.895
r49 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=2.52
+ $X2=2.865 $Y2=2.52
r50 9 11 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.63 $Y=2.52
+ $X2=3.742 $Y2=2.605
r51 9 10 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.63 $Y=2.52 $X2=3.03
+ $Y2=2.52
r52 2 18 600 $w=1.7e-07 $l=9.57445e-07 $layer=licon1_PDIFF $count=1 $X=4.55
+ $Y=1.835 $X2=4.69 $Y2=2.725
r53 1 16 300 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.835 $X2=2.865 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%Y 1 2 3 4 13 21 23 24 25 26 27 36 37 38 39
+ 40 41 42 51 55 57
c61 26 0 7.76303e-20 $X=5.645 $Y=1.15
r62 55 57 2.56098 $w=2.68e-07 $l=6e-08 $layer=LI1_cond $X=6.02 $Y=1.235 $X2=6.02
+ $Y2=1.295
r63 42 69 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.02 $Y=2.775
+ $X2=6.02 $Y2=2.91
r64 41 42 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.02 $Y=2.405
+ $X2=6.02 $Y2=2.775
r65 40 41 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.02 $Y=1.98
+ $X2=6.02 $Y2=2.405
r66 38 55 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=1.15 $X2=6.02
+ $Y2=1.235
r67 38 39 15.2805 $w=2.68e-07 $l=3.58e-07 $layer=LI1_cond $X=6.02 $Y=1.307
+ $X2=6.02 $Y2=1.665
r68 38 57 0.512197 $w=2.68e-07 $l=1.2e-08 $layer=LI1_cond $X=6.02 $Y=1.307
+ $X2=6.02 $Y2=1.295
r69 37 51 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=5.48 $Y=0.925
+ $X2=5.48 $Y2=0.68
r70 35 40 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.02 $Y=1.945
+ $X2=6.02 $Y2=1.98
r71 35 36 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=1.945
+ $X2=6.02 $Y2=1.86
r72 34 39 4.69514 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.02 $Y=1.775
+ $X2=6.02 $Y2=1.665
r73 34 36 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=1.775
+ $X2=6.02 $Y2=1.86
r74 33 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.48 $Y=1.065
+ $X2=5.48 $Y2=0.925
r75 27 30 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=4.225 $Y=2.345
+ $X2=4.225 $Y2=2.425
r76 26 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.645 $Y=1.15
+ $X2=5.48 $Y2=1.065
r77 25 38 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.885 $Y=1.15
+ $X2=6.02 $Y2=1.15
r78 25 26 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.885 $Y=1.15
+ $X2=5.645 $Y2=1.15
r79 23 36 3.05049 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.885 $Y=1.86
+ $X2=6.02 $Y2=1.86
r80 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.885 $Y=1.86
+ $X2=5.215 $Y2=1.86
r81 19 32 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.43 $X2=5.12
+ $Y2=2.345
r82 19 21 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=5.12 $Y=2.43
+ $X2=5.12 $Y2=2.455
r83 16 32 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.26 $X2=5.12
+ $Y2=2.345
r84 16 18 16.3445 $w=1.88e-07 $l=2.8e-07 $layer=LI1_cond $X=5.12 $Y=2.26
+ $X2=5.12 $Y2=1.98
r85 15 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.12 $Y=1.945
+ $X2=5.215 $Y2=1.86
r86 15 18 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=5.12 $Y=1.945
+ $X2=5.12 $Y2=1.98
r87 14 27 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.355 $Y=2.345
+ $X2=4.225 $Y2=2.345
r88 13 32 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.025 $Y=2.345
+ $X2=5.12 $Y2=2.345
r89 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.025 $Y=2.345
+ $X2=4.355 $Y2=2.345
r90 4 69 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.84
+ $Y=1.835 $X2=5.98 $Y2=2.91
r91 4 40 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.84
+ $Y=1.835 $X2=5.98 $Y2=1.98
r92 3 21 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=4.98
+ $Y=1.835 $X2=5.12 $Y2=2.455
r93 3 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.835 $X2=5.12 $Y2=1.98
r94 2 30 600 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.835 $X2=4.26 $Y2=2.425
r95 1 51 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.325 $X2=5.48 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%A_27_47# 1 2 3 12 14 15 17 18 19 25
c52 25 0 1.88077e-19 $X=2.35 $Y=0.38
c53 15 0 1.37872e-19 $X=0.425 $Y=0.82
c54 14 0 8.28055e-20 $X=0.975 $Y=0.82
r55 19 21 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.145 $Y=0.35
+ $X2=1.42 $Y2=0.35
r56 18 25 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0.35
+ $X2=2.35 $Y2=0.35
r57 18 21 44.6555 $w=1.88e-07 $l=7.65e-07 $layer=LI1_cond $X=2.185 $Y=0.35
+ $X2=1.42 $Y2=0.35
r58 16 19 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.06 $Y=0.445
+ $X2=1.145 $Y2=0.35
r59 16 17 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.06 $Y=0.445
+ $X2=1.06 $Y2=0.735
r60 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=0.82
+ $X2=1.06 $Y2=0.735
r61 14 15 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.975 $Y=0.82
+ $X2=0.425 $Y2=0.82
r62 10 15 7.68211 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=0.735
+ $X2=0.425 $Y2=0.82
r63 10 12 11.3444 $w=3.18e-07 $l=3.15e-07 $layer=LI1_cond $X=0.255 $Y=0.735
+ $X2=0.255 $Y2=0.42
r64 3 25 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.14
+ $Y=0.235 $X2=2.35 $Y2=0.38
r65 2 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.235 $X2=1.42 $Y2=0.36
r66 1 12 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%VGND 1 2 3 12 16 18 22 24 25 26 28 45 46 49
+ 52 62
c80 28 0 1.37872e-19 $X=0.585 $Y=0
r81 55 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.36
+ $Y2=0
r82 53 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r83 52 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r84 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r85 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r87 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r88 43 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r89 42 45 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6 $Y2=0
r90 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r91 40 52 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=4.405
+ $Y2=0
r92 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=5.04
+ $Y2=0
r93 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r94 35 38 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r95 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r96 33 49 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.695
+ $Y2=0
r97 33 35 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=1.2
+ $Y2=0
r98 31 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r99 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r100 28 49 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.695
+ $Y2=0
r101 28 30 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r102 26 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=3.36 $Y2=0
r103 26 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=1.2
+ $Y2=0
r104 26 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r105 24 38 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.12
+ $Y2=0
r106 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.33
+ $Y2=0
r107 20 52 3.03114 $w=7.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=0.085
+ $X2=4.405 $Y2=0
r108 20 22 5.74432 $w=7.58e-07 $l=3.65e-07 $layer=LI1_cond $X=4.405 $Y=0.085
+ $X2=4.405 $Y2=0.45
r109 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.33
+ $Y2=0
r110 18 52 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=4.405
+ $Y2=0
r111 18 19 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=3.495 $Y2=0
r112 14 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0.085
+ $X2=3.33 $Y2=0
r113 14 16 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.33 $Y=0.085
+ $X2=3.33 $Y2=0.45
r114 10 49 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r115 10 12 16.5009 $w=2.18e-07 $l=3.15e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.4
r116 3 22 45.5 $w=1.7e-07 $l=6.29404e-07 $layer=licon1_NDIFF $count=4 $X=4.05
+ $Y=0.325 $X2=4.62 $Y2=0.45
r117 2 16 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.19
+ $Y=0.325 $X2=3.33 $Y2=0.45
r118 1 12 182 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.72 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_2%A_555_65# 1 2 3 4 15 17 18 21 23 29 30 33 35
r64 31 33 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.98 $Y=0.425
+ $X2=5.98 $Y2=0.47
r65 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.815 $Y=0.34
+ $X2=5.98 $Y2=0.425
r66 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.815 $Y=0.34
+ $X2=5.145 $Y2=0.34
r67 26 28 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=5.05 $Y=1.065
+ $X2=5.05 $Y2=0.47
r68 25 30 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.05 $Y=0.425
+ $X2=5.145 $Y2=0.34
r69 25 28 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=5.05 $Y=0.425
+ $X2=5.05 $Y2=0.47
r70 24 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.855 $Y=1.15
+ $X2=3.76 $Y2=1.15
r71 23 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.955 $Y=1.15
+ $X2=5.05 $Y2=1.065
r72 23 24 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=4.955 $Y=1.15
+ $X2=3.855 $Y2=1.15
r73 19 35 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=1.065
+ $X2=3.76 $Y2=1.15
r74 19 21 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=3.76 $Y=1.065
+ $X2=3.76 $Y2=0.47
r75 17 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.665 $Y=1.15
+ $X2=3.76 $Y2=1.15
r76 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.665 $Y=1.15
+ $X2=2.995 $Y2=1.15
r77 13 18 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.9 $Y=1.065
+ $X2=2.995 $Y2=1.15
r78 13 15 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=2.9 $Y=1.065
+ $X2=2.9 $Y2=0.47
r79 4 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.77
+ $Y=0.325 $X2=5.98 $Y2=0.47
r80 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.325 $X2=5.05 $Y2=0.47
r81 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.62
+ $Y=0.325 $X2=3.76 $Y2=0.47
r82 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.325 $X2=2.9 $Y2=0.47
.ends

