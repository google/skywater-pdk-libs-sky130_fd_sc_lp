* File: sky130_fd_sc_lp__a21o_2.pxi.spice
* Created: Fri Aug 28 09:50:54 2020
* 
x_PM_SKY130_FD_SC_LP__A21O_2%A_86_269# N_A_86_269#_M1003_d N_A_86_269#_M1000_s
+ N_A_86_269#_M1002_g N_A_86_269#_M1001_g N_A_86_269#_M1006_g
+ N_A_86_269#_M1009_g N_A_86_269#_c_62_n N_A_86_269#_c_63_n N_A_86_269#_c_113_p
+ N_A_86_269#_c_70_n N_A_86_269#_c_71_n N_A_86_269#_c_72_n N_A_86_269#_c_73_n
+ N_A_86_269#_c_93_p N_A_86_269#_c_64_n N_A_86_269#_c_65_n N_A_86_269#_c_66_n
+ PM_SKY130_FD_SC_LP__A21O_2%A_86_269#
x_PM_SKY130_FD_SC_LP__A21O_2%B1 N_B1_M1003_g N_B1_M1000_g B1 N_B1_c_140_n
+ N_B1_c_141_n PM_SKY130_FD_SC_LP__A21O_2%B1
x_PM_SKY130_FD_SC_LP__A21O_2%A1 N_A1_M1005_g N_A1_M1007_g A1 A1 A1 N_A1_c_179_n
+ N_A1_c_180_n PM_SKY130_FD_SC_LP__A21O_2%A1
x_PM_SKY130_FD_SC_LP__A21O_2%A2 N_A2_c_214_n N_A2_M1008_g N_A2_M1004_g A2
+ N_A2_c_217_n PM_SKY130_FD_SC_LP__A21O_2%A2
x_PM_SKY130_FD_SC_LP__A21O_2%VPWR N_VPWR_M1002_s N_VPWR_M1006_s N_VPWR_M1007_d
+ N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n
+ N_VPWR_c_243_n VPWR N_VPWR_c_244_n N_VPWR_c_245_n N_VPWR_c_237_n
+ N_VPWR_c_247_n PM_SKY130_FD_SC_LP__A21O_2%VPWR
x_PM_SKY130_FD_SC_LP__A21O_2%X N_X_M1001_d N_X_M1002_d N_X_c_303_p N_X_c_285_n X
+ X X X X PM_SKY130_FD_SC_LP__A21O_2%X
x_PM_SKY130_FD_SC_LP__A21O_2%A_392_367# N_A_392_367#_M1000_d
+ N_A_392_367#_M1004_d N_A_392_367#_c_321_n N_A_392_367#_c_306_n
+ N_A_392_367#_c_307_n N_A_392_367#_c_325_n
+ PM_SKY130_FD_SC_LP__A21O_2%A_392_367#
x_PM_SKY130_FD_SC_LP__A21O_2%VGND N_VGND_M1001_s N_VGND_M1009_s N_VGND_M1008_d
+ N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n
+ N_VGND_c_332_n N_VGND_c_333_n VGND N_VGND_c_334_n N_VGND_c_335_n
+ N_VGND_c_336_n PM_SKY130_FD_SC_LP__A21O_2%VGND
cc_1 VNB N_A_86_269#_M1002_g 0.0127435f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_2 VNB N_A_86_269#_M1001_g 0.0279042f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.655
cc_3 VNB N_A_86_269#_M1009_g 0.0238406f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.655
cc_4 VNB N_A_86_269#_c_62_n 8.55094e-19 $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.93
cc_5 VNB N_A_86_269#_c_63_n 0.0086267f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.07
cc_6 VNB N_A_86_269#_c_64_n 0.0010458f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.51
cc_7 VNB N_A_86_269#_c_65_n 0.00183661f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.345
cc_8 VNB N_A_86_269#_c_66_n 0.0493127f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.585
cc_9 VNB N_B1_M1003_g 0.0279881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_140_n 0.0323445f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.655
cc_11 VNB N_B1_c_141_n 0.00359659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1007_g 0.00777322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A1 0.00900496f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_14 VNB N_A1_c_179_n 0.0309412f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.655
cc_15 VNB N_A1_c_180_n 0.0179801f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.515
cc_16 VNB N_A2_c_214_n 0.0226082f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=0.235
cc_17 VNB N_A2_M1004_g 0.0116295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A2 0.0204241f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_19 VNB N_A2_c_217_n 0.0451421f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.655
cc_20 VNB N_VPWR_c_237_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.345
cc_21 VNB N_X_c_285_n 0.00718784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB X 0.010912f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_23 VNB N_VGND_c_327_n 0.0265527f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.655
cc_24 VNB N_VGND_c_328_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_329_n 0.00274225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_330_n 0.0132956f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.655
cc_27 VNB N_VGND_c_331_n 0.0348057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_332_n 0.0115308f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.93
cc_29 VNB N_VGND_c_333_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.155
cc_30 VNB N_VGND_c_334_n 0.0377663f $X=-0.19 $Y=-0.245 $X2=1.662 $Y2=2.1
cc_31 VNB N_VGND_c_335_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.51
cc_32 VNB N_VGND_c_336_n 0.199517f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=2.095
cc_33 VPB N_A_86_269#_M1002_g 0.0272177f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_34 VPB N_A_86_269#_M1006_g 0.0222235f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_35 VPB N_A_86_269#_c_62_n 0.00291991f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.93
cc_36 VPB N_A_86_269#_c_70_n 0.0131344f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=2.015
cc_37 VPB N_A_86_269#_c_71_n 0.00108717f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=2.015
cc_38 VPB N_A_86_269#_c_72_n 5.52007e-19 $X=-0.19 $Y=1.655 $X2=1.662 $Y2=2.1
cc_39 VPB N_A_86_269#_c_73_n 0.0100398f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=2.91
cc_40 VPB N_A_86_269#_c_66_n 0.00917678f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.585
cc_41 VPB N_B1_M1000_g 0.0233895f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.495
cc_42 VPB N_B1_c_140_n 0.00984439f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.655
cc_43 VPB N_B1_c_141_n 0.00365378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A1_M1007_g 0.018992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A2_M1004_g 0.0247156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_238_n 0.0117405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_239_n 0.0653449f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.655
cc_48 VPB N_VPWR_c_240_n 0.0106046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_241_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_242_n 0.0277741f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=1.07
cc_51 VPB N_VPWR_c_243_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=1.07
cc_52 VPB N_VPWR_c_244_n 0.0148832f $X=-0.19 $Y=1.655 $X2=1.662 $Y2=2.1
cc_53 VPB N_VPWR_c_245_n 0.0195708f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.51
cc_54 VPB N_VPWR_c_237_n 0.0590296f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.345
cc_55 VPB N_VPWR_c_247_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.585
cc_56 VPB X 0.00394414f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_57 VPB N_A_392_367#_c_306_n 0.0108567f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.655
cc_58 VPB N_A_392_367#_c_307_n 0.00582179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 N_A_86_269#_M1009_g N_B1_M1003_g 0.0282574f $X=1.105 $Y=0.655 $X2=0 $Y2=0
cc_60 N_A_86_269#_c_63_n N_B1_M1003_g 0.0144425f $X=1.705 $Y=1.07 $X2=0 $Y2=0
cc_61 N_A_86_269#_c_65_n N_B1_M1003_g 0.00388731f $X=1.155 $Y=1.345 $X2=0 $Y2=0
cc_62 N_A_86_269#_c_62_n N_B1_M1000_g 0.00283713f $X=1.155 $Y=1.93 $X2=0 $Y2=0
cc_63 N_A_86_269#_c_72_n N_B1_M1000_g 0.00166559f $X=1.662 $Y=2.1 $X2=0 $Y2=0
cc_64 N_A_86_269#_c_73_n N_B1_M1000_g 0.00961377f $X=1.67 $Y=2.91 $X2=0 $Y2=0
cc_65 N_A_86_269#_c_63_n N_B1_c_140_n 0.00435593f $X=1.705 $Y=1.07 $X2=0 $Y2=0
cc_66 N_A_86_269#_c_72_n N_B1_c_140_n 0.00168846f $X=1.662 $Y=2.1 $X2=0 $Y2=0
cc_67 N_A_86_269#_c_64_n N_B1_c_140_n 0.00105401f $X=1.115 $Y=1.51 $X2=0 $Y2=0
cc_68 N_A_86_269#_c_66_n N_B1_c_140_n 0.018208f $X=1.105 $Y=1.585 $X2=0 $Y2=0
cc_69 N_A_86_269#_M1006_g N_B1_c_141_n 3.21246e-19 $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_86_269#_c_63_n N_B1_c_141_n 0.0232879f $X=1.705 $Y=1.07 $X2=0 $Y2=0
cc_71 N_A_86_269#_c_70_n N_B1_c_141_n 6.92291e-19 $X=1.505 $Y=2.015 $X2=0 $Y2=0
cc_72 N_A_86_269#_c_72_n N_B1_c_141_n 0.0252087f $X=1.662 $Y=2.1 $X2=0 $Y2=0
cc_73 N_A_86_269#_c_64_n N_B1_c_141_n 0.0345441f $X=1.115 $Y=1.51 $X2=0 $Y2=0
cc_74 N_A_86_269#_c_66_n N_B1_c_141_n 9.99602e-19 $X=1.105 $Y=1.585 $X2=0 $Y2=0
cc_75 N_A_86_269#_M1003_d A1 0.00774813f $X=1.67 $Y=0.235 $X2=0 $Y2=0
cc_76 N_A_86_269#_c_63_n A1 0.0155216f $X=1.705 $Y=1.07 $X2=0 $Y2=0
cc_77 N_A_86_269#_c_93_p A1 0.0545642f $X=1.81 $Y=0.42 $X2=0 $Y2=0
cc_78 N_A_86_269#_c_63_n N_A1_c_180_n 6.1033e-19 $X=1.705 $Y=1.07 $X2=0 $Y2=0
cc_79 N_A_86_269#_c_93_p N_A1_c_180_n 0.00319208f $X=1.81 $Y=0.42 $X2=0 $Y2=0
cc_80 N_A_86_269#_c_62_n N_VPWR_M1006_s 3.48153e-19 $X=1.155 $Y=1.93 $X2=0 $Y2=0
cc_81 N_A_86_269#_c_71_n N_VPWR_M1006_s 0.00310159f $X=1.325 $Y=2.015 $X2=0
+ $Y2=0
cc_82 N_A_86_269#_M1002_g N_VPWR_c_239_n 0.0076281f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_83 N_A_86_269#_M1002_g N_VPWR_c_240_n 6.93887e-19 $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_84 N_A_86_269#_M1006_g N_VPWR_c_240_n 0.0171543f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_85 N_A_86_269#_c_71_n N_VPWR_c_240_n 0.0243971f $X=1.325 $Y=2.015 $X2=0 $Y2=0
cc_86 N_A_86_269#_c_73_n N_VPWR_c_240_n 0.0617695f $X=1.67 $Y=2.91 $X2=0 $Y2=0
cc_87 N_A_86_269#_c_66_n N_VPWR_c_240_n 8.18092e-19 $X=1.105 $Y=1.585 $X2=0
+ $Y2=0
cc_88 N_A_86_269#_c_73_n N_VPWR_c_242_n 0.0200241f $X=1.67 $Y=2.91 $X2=0 $Y2=0
cc_89 N_A_86_269#_M1002_g N_VPWR_c_244_n 0.00585385f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_90 N_A_86_269#_M1006_g N_VPWR_c_244_n 0.00486043f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_91 N_A_86_269#_M1000_s N_VPWR_c_237_n 0.00215158f $X=1.545 $Y=1.835 $X2=0
+ $Y2=0
cc_92 N_A_86_269#_M1002_g N_VPWR_c_237_n 0.0114959f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_93 N_A_86_269#_M1006_g N_VPWR_c_237_n 0.00824727f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_A_86_269#_c_73_n N_VPWR_c_237_n 0.0120544f $X=1.67 $Y=2.91 $X2=0 $Y2=0
cc_95 N_A_86_269#_M1001_g N_X_c_285_n 0.0117891f $X=0.675 $Y=0.655 $X2=0 $Y2=0
cc_96 N_A_86_269#_M1009_g N_X_c_285_n 6.07664e-19 $X=1.105 $Y=0.655 $X2=0 $Y2=0
cc_97 N_A_86_269#_c_113_p N_X_c_285_n 0.0104823f $X=1.325 $Y=1.07 $X2=0 $Y2=0
cc_98 N_A_86_269#_c_66_n N_X_c_285_n 0.00412479f $X=1.105 $Y=1.585 $X2=0 $Y2=0
cc_99 N_A_86_269#_M1002_g X 0.00947569f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_86_269#_M1001_g X 0.00675591f $X=0.675 $Y=0.655 $X2=0 $Y2=0
cc_101 N_A_86_269#_M1009_g X 0.00134296f $X=1.105 $Y=0.655 $X2=0 $Y2=0
cc_102 N_A_86_269#_c_64_n X 0.0406171f $X=1.115 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A_86_269#_c_65_n X 0.00828283f $X=1.155 $Y=1.345 $X2=0 $Y2=0
cc_104 N_A_86_269#_c_66_n X 0.0173837f $X=1.105 $Y=1.585 $X2=0 $Y2=0
cc_105 N_A_86_269#_c_62_n N_A_392_367#_c_307_n 0.00282906f $X=1.155 $Y=1.93
+ $X2=0 $Y2=0
cc_106 N_A_86_269#_c_63_n N_VGND_M1009_s 0.00145634f $X=1.705 $Y=1.07 $X2=0
+ $Y2=0
cc_107 N_A_86_269#_c_113_p N_VGND_M1009_s 9.73829e-19 $X=1.325 $Y=1.07 $X2=0
+ $Y2=0
cc_108 N_A_86_269#_M1001_g N_VGND_c_327_n 0.0110384f $X=0.675 $Y=0.655 $X2=0
+ $Y2=0
cc_109 N_A_86_269#_M1009_g N_VGND_c_327_n 6.0835e-19 $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_110 N_A_86_269#_c_66_n N_VGND_c_327_n 0.00446639f $X=1.105 $Y=1.585 $X2=0
+ $Y2=0
cc_111 N_A_86_269#_M1001_g N_VGND_c_328_n 0.00486043f $X=0.675 $Y=0.655 $X2=0
+ $Y2=0
cc_112 N_A_86_269#_M1009_g N_VGND_c_328_n 0.00486043f $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_113 N_A_86_269#_M1001_g N_VGND_c_329_n 6.0835e-19 $X=0.675 $Y=0.655 $X2=0
+ $Y2=0
cc_114 N_A_86_269#_M1009_g N_VGND_c_329_n 0.0099551f $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_115 N_A_86_269#_c_63_n N_VGND_c_329_n 0.011191f $X=1.705 $Y=1.07 $X2=0 $Y2=0
cc_116 N_A_86_269#_c_113_p N_VGND_c_329_n 0.00992353f $X=1.325 $Y=1.07 $X2=0
+ $Y2=0
cc_117 N_A_86_269#_c_66_n N_VGND_c_329_n 2.8405e-19 $X=1.105 $Y=1.585 $X2=0
+ $Y2=0
cc_118 N_A_86_269#_c_93_p N_VGND_c_334_n 0.0124873f $X=1.81 $Y=0.42 $X2=0 $Y2=0
cc_119 N_A_86_269#_M1003_d N_VGND_c_336_n 0.0112763f $X=1.67 $Y=0.235 $X2=0
+ $Y2=0
cc_120 N_A_86_269#_M1001_g N_VGND_c_336_n 0.00824727f $X=0.675 $Y=0.655 $X2=0
+ $Y2=0
cc_121 N_A_86_269#_M1009_g N_VGND_c_336_n 0.00824727f $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_122 N_A_86_269#_c_93_p N_VGND_c_336_n 0.00730901f $X=1.81 $Y=0.42 $X2=0 $Y2=0
cc_123 N_B1_c_140_n N_A1_M1007_g 0.0260523f $X=1.685 $Y=1.51 $X2=0 $Y2=0
cc_124 N_B1_c_141_n N_A1_M1007_g 8.62894e-19 $X=1.685 $Y=1.51 $X2=0 $Y2=0
cc_125 N_B1_M1003_g A1 0.00464548f $X=1.595 $Y=0.655 $X2=0 $Y2=0
cc_126 N_B1_c_140_n A1 0.00135506f $X=1.685 $Y=1.51 $X2=0 $Y2=0
cc_127 N_B1_c_141_n A1 0.0108529f $X=1.685 $Y=1.51 $X2=0 $Y2=0
cc_128 N_B1_c_140_n N_A1_c_179_n 0.006166f $X=1.685 $Y=1.51 $X2=0 $Y2=0
cc_129 N_B1_M1003_g N_A1_c_180_n 0.0171617f $X=1.595 $Y=0.655 $X2=0 $Y2=0
cc_130 N_B1_M1000_g N_VPWR_c_240_n 0.00363414f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B1_M1000_g N_VPWR_c_241_n 0.0013327f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_132 N_B1_M1000_g N_VPWR_c_242_n 0.00571722f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_133 N_B1_M1000_g N_VPWR_c_237_n 0.0117938f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B1_M1000_g N_A_392_367#_c_307_n 0.0019217f $X=1.885 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_B1_c_141_n N_A_392_367#_c_307_n 0.00631736f $X=1.685 $Y=1.51 $X2=0
+ $Y2=0
cc_136 N_B1_M1003_g N_VGND_c_329_n 0.00612025f $X=1.595 $Y=0.655 $X2=0 $Y2=0
cc_137 N_B1_M1003_g N_VGND_c_334_n 0.00585385f $X=1.595 $Y=0.655 $X2=0 $Y2=0
cc_138 N_B1_M1003_g N_VGND_c_336_n 0.0113398f $X=1.595 $Y=0.655 $X2=0 $Y2=0
cc_139 A1 N_A2_c_214_n 0.028804f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_140 N_A1_c_180_n N_A2_c_214_n 0.0321041f $X=2.335 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A1_M1007_g N_A2_M1004_g 0.0233828f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_142 A1 A2 0.0263479f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A1_c_179_n A2 2.04525e-19 $X=2.335 $Y=1.35 $X2=0 $Y2=0
cc_144 A1 N_A2_c_217_n 0.0087931f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_145 N_A1_c_179_n N_A2_c_217_n 0.0214455f $X=2.335 $Y=1.35 $X2=0 $Y2=0
cc_146 N_A1_M1007_g N_VPWR_c_241_n 0.0145911f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A1_M1007_g N_VPWR_c_242_n 0.00564095f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A1_M1007_g N_VPWR_c_237_n 0.00950825f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A1_M1007_g N_A_392_367#_c_306_n 0.0144298f $X=2.315 $Y=2.465 $X2=0
+ $Y2=0
cc_150 A1 N_A_392_367#_c_306_n 0.041742f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_151 N_A1_c_179_n N_A_392_367#_c_306_n 9.47144e-19 $X=2.335 $Y=1.35 $X2=0
+ $Y2=0
cc_152 A1 N_A_392_367#_c_307_n 0.0137565f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_153 N_A1_c_179_n N_A_392_367#_c_307_n 3.51912e-19 $X=2.335 $Y=1.35 $X2=0
+ $Y2=0
cc_154 A1 N_VGND_c_334_n 0.0293282f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A1_c_180_n N_VGND_c_334_n 0.00369917f $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_156 A1 N_VGND_c_336_n 0.0243531f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A1_c_180_n N_VGND_c_336_n 0.00623646f $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_158 A1 A_464_47# 0.00420714f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_159 N_A2_M1004_g N_VPWR_c_241_n 0.0154114f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_M1004_g N_VPWR_c_245_n 0.00564095f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A2_M1004_g N_VPWR_c_237_n 0.0104973f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A2_M1004_g N_A_392_367#_c_306_n 0.019714f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_163 A2 N_A_392_367#_c_306_n 0.0168667f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A2_c_217_n N_A_392_367#_c_306_n 0.00646977f $X=2.99 $Y=1.35 $X2=0 $Y2=0
cc_165 N_A2_c_214_n N_VGND_c_331_n 0.00615214f $X=2.785 $Y=1.185 $X2=0 $Y2=0
cc_166 A2 N_VGND_c_331_n 0.0217847f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A2_c_217_n N_VGND_c_331_n 0.0057671f $X=2.99 $Y=1.35 $X2=0 $Y2=0
cc_168 N_A2_c_214_n N_VGND_c_334_n 0.0055091f $X=2.785 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A2_c_214_n N_VGND_c_336_n 0.0111429f $X=2.785 $Y=1.185 $X2=0 $Y2=0
cc_170 N_VPWR_c_237_n N_X_M1002_d 0.00397496f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_239_n X 0.00152359f $X=0.29 $Y=1.98 $X2=0 $Y2=0
cc_172 N_VPWR_c_244_n X 0.0138717f $X=0.985 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_c_237_n X 0.00886411f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_c_237_n N_A_392_367#_M1000_d 0.0041489f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_175 N_VPWR_c_237_n N_A_392_367#_M1004_d 0.00375181f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_242_n N_A_392_367#_c_321_n 0.0136943f $X=2.385 $Y=3.33 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_237_n N_A_392_367#_c_321_n 0.00866972f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_178 N_VPWR_M1007_d N_A_392_367#_c_306_n 0.00218982f $X=2.39 $Y=1.835 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_241_n N_A_392_367#_c_306_n 0.017285f $X=2.55 $Y=2.11 $X2=0 $Y2=0
cc_180 N_VPWR_c_245_n N_A_392_367#_c_325_n 0.0142484f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_237_n N_A_392_367#_c_325_n 0.00847534f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_182 N_X_c_285_n N_VGND_c_327_n 0.00178608f $X=0.89 $Y=1.07 $X2=0 $Y2=0
cc_183 N_X_c_303_p N_VGND_c_328_n 0.0124525f $X=0.89 $Y=0.42 $X2=0 $Y2=0
cc_184 N_X_M1001_d N_VGND_c_336_n 0.00536646f $X=0.75 $Y=0.235 $X2=0 $Y2=0
cc_185 N_X_c_303_p N_VGND_c_336_n 0.00730901f $X=0.89 $Y=0.42 $X2=0 $Y2=0
cc_186 N_VGND_c_336_n A_464_47# 0.00320415f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
