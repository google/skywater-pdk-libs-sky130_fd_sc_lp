* File: sky130_fd_sc_lp__iso0p_lp2.pex.spice
* Created: Fri Aug 28 10:40:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%SLEEP 1 3 6 8 10 11 12 16 17
c30 16 0 7.63997e-20 $X=0.71 $Y=1.175
r31 16 18 67.4279 $w=5.1e-07 $l=5.1e-07 $layer=POLY_cond $X=0.665 $Y=1.175
+ $X2=0.665 $Y2=1.685
r32 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=1.175 $X2=0.71 $Y2=1.175
r33 11 12 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.732 $Y=1.295
+ $X2=0.732 $Y2=1.665
r34 11 17 3.68782 $w=3.73e-07 $l=1.2e-07 $layer=LI1_cond $X=0.732 $Y=1.295
+ $X2=0.732 $Y2=1.175
r35 8 16 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.845 $Y=1.01
+ $X2=0.665 $Y2=1.175
r36 8 10 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.845 $Y=1.01
+ $X2=0.845 $Y2=0.675
r37 6 18 223.608 $w=2.5e-07 $l=9e-07 $layer=POLY_cond $X=0.535 $Y=2.585
+ $X2=0.535 $Y2=1.685
r38 1 16 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.485 $Y=1.01
+ $X2=0.665 $Y2=1.175
r39 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.485 $Y=1.01
+ $X2=0.485 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%A_27_93# 1 2 7 9 11 13 16 20 24 28 31
c59 24 0 1.32657e-19 $X=1.2 $Y=2.035
c60 11 0 4.20716e-20 $X=1.625 $Y=1.01
c61 9 0 7.63997e-20 $X=1.585 $Y=2.585
r62 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.43
+ $Y=1.175 $X2=1.43 $Y2=1.175
r63 26 28 22.6112 $w=3.93e-07 $l=7.75e-07 $layer=LI1_cond $X=1.397 $Y=1.95
+ $X2=1.397 $Y2=1.175
r64 25 31 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.375 $Y=2.035
+ $X2=0.265 $Y2=2.035
r65 24 26 8.32734 $w=1.7e-07 $l=2.35699e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=1.397 $Y2=1.95
r66 24 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=0.375 $Y2=2.035
r67 20 22 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=0.265 $Y=2.23
+ $X2=0.265 $Y2=2.91
r68 18 31 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.12
+ $X2=0.265 $Y2=2.035
r69 18 20 5.76222 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=0.265 $Y=2.12
+ $X2=0.265 $Y2=2.23
r70 14 31 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=1.95
+ $X2=0.265 $Y2=2.035
r71 14 16 64.432 $w=2.18e-07 $l=1.23e-06 $layer=LI1_cond $X=0.265 $Y=1.95
+ $X2=0.265 $Y2=0.72
r72 11 29 42.0549 $w=5.05e-07 $l=2.38642e-07 $layer=POLY_cond $X=1.625 $Y=1.01
+ $X2=1.455 $Y2=1.175
r73 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.625 $Y=1.01
+ $X2=1.625 $Y2=0.675
r74 7 29 60.4941 $w=5.05e-07 $l=5.66282e-07 $layer=POLY_cond $X=1.585 $Y=1.68
+ $X2=1.455 $Y2=1.175
r75 7 9 224.851 $w=2.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.585 $Y=1.68
+ $X2=1.585 $Y2=2.585
r76 2 22 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.27 $Y2=2.91
r77 2 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.27 $Y2=2.23
r78 1 16 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.27 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%A 3 5 8 10 11 12 13 18 22
c46 22 0 1.57318e-19 $X=2.145 $Y=1.48
c47 8 0 1.32657e-19 $X=2.135 $Y=2.585
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.145
+ $Y=1.48 $X2=2.145 $Y2=1.48
r49 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.48 $X2=2.485 $Y2=1.48
r50 16 22 1.50692 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.26 $Y=1.48
+ $X2=2.12 $Y2=1.48
r51 16 18 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.26 $Y=1.48
+ $X2=2.485 $Y2=1.48
r52 13 19 5.03179 $w=3.53e-07 $l=1.55e-07 $layer=LI1_cond $X=2.64 $Y=1.572
+ $X2=2.485 $Y2=1.572
r53 12 19 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=2.16 $Y=1.572
+ $X2=2.485 $Y2=1.572
r54 12 23 0.486948 $w=3.53e-07 $l=1.5e-08 $layer=LI1_cond $X=2.16 $Y=1.572
+ $X2=2.145 $Y2=1.572
r55 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.02 $Y=0.995
+ $X2=2.02 $Y2=1.145
r56 6 22 30.2679 $w=2e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.135 $Y=1.645
+ $X2=2.12 $Y2=1.48
r57 6 8 233.546 $w=2.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.135 $Y=1.645
+ $X2=2.135 $Y2=2.585
r58 5 22 30.2679 $w=2e-07 $l=1.94808e-07 $layer=POLY_cond $X=2.055 $Y=1.315
+ $X2=2.12 $Y2=1.48
r59 5 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.055 $Y=1.315
+ $X2=2.055 $Y2=1.145
r60 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.985 $Y=0.675
+ $X2=1.985 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%A_342_417# 1 2 7 9 12 14 16 19 23 24 27 29
+ 30 31 32 35
c64 27 0 4.20716e-20 $X=2.2 $Y=0.72
c65 23 0 1.57318e-19 $X=2.925 $Y=2.04
r66 35 37 67.9525 $w=5.1e-07 $l=5.15e-07 $layer=POLY_cond $X=3.115 $Y=1.17
+ $X2=3.115 $Y2=1.685
r67 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.06
+ $Y=1.17 $X2=3.06 $Y2=1.17
r68 31 34 2.96055 $w=3.05e-07 $l=1.1e-07 $layer=LI1_cond $X=3.077 $Y=1.225
+ $X2=3.077 $Y2=1.115
r69 31 32 27.5831 $w=3.03e-07 $l=7.3e-07 $layer=LI1_cond $X=3.077 $Y=1.225
+ $X2=3.077 $Y2=1.955
r70 29 34 4.09094 $w=2.2e-07 $l=1.52e-07 $layer=LI1_cond $X=2.925 $Y=1.115
+ $X2=3.077 $Y2=1.115
r71 29 30 32.4779 $w=2.18e-07 $l=6.2e-07 $layer=LI1_cond $X=2.925 $Y=1.115
+ $X2=2.305 $Y2=1.115
r72 25 30 6.82129 $w=2.2e-07 $l=1.53786e-07 $layer=LI1_cond $X=2.2 $Y=1.005
+ $X2=2.305 $Y2=1.115
r73 25 27 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.2 $Y=1.005
+ $X2=2.2 $Y2=0.72
r74 23 32 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=2.925 $Y=2.04
+ $X2=3.077 $Y2=1.955
r75 23 24 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.925 $Y=2.04
+ $X2=1.975 $Y2=2.04
r76 19 21 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=1.87 $Y=2.23
+ $X2=1.87 $Y2=2.91
r77 17 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.87 $Y=2.125
+ $X2=1.975 $Y2=2.04
r78 17 19 5.54545 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=1.87 $Y=2.125
+ $X2=1.87 $Y2=2.23
r79 14 35 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=3.295 $Y=1.005
+ $X2=3.115 $Y2=1.17
r80 14 16 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.295 $Y=1.005
+ $X2=3.295 $Y2=0.675
r81 12 37 223.608 $w=2.5e-07 $l=9e-07 $layer=POLY_cond $X=3.245 $Y=2.585
+ $X2=3.245 $Y2=1.685
r82 7 35 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.935 $Y=1.005
+ $X2=3.115 $Y2=1.17
r83 7 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.935 $Y=1.005
+ $X2=2.935 $Y2=0.675
r84 2 21 400 $w=1.7e-07 $l=9.01457e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.87 $Y2=2.91
r85 2 19 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.87 $Y2=2.23
r86 1 27 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.465 $X2=2.2 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%KAPWR 1 2 7 10 17 21
r35 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.98 $Y=2.775
+ $X2=2.98 $Y2=2.775
r36 17 20 5.09451 $w=9.08e-07 $l=3.8e-07 $layer=LI1_cond $X=2.69 $Y=2.395
+ $X2=2.69 $Y2=2.775
r37 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.32 $Y=2.775
+ $X2=1.32 $Y2=2.775
r38 10 13 5.45412 $w=8.48e-07 $l=3.8e-07 $layer=LI1_cond $X=1.06 $Y=2.395
+ $X2=1.06 $Y2=2.775
r39 7 21 0.680101 $w=2.3e-07 $l=1.06e-06 $layer=MET1_cond $X=1.92 $Y=2.775
+ $X2=2.98 $Y2=2.775
r40 7 14 0.384963 $w=2.3e-07 $l=6e-07 $layer=MET1_cond $X=1.92 $Y=2.775 $X2=1.32
+ $Y2=2.775
r41 2 17 150 $w=1.7e-07 $l=8.61162e-07 $layer=licon1_PDIFF $count=4 $X=2.26
+ $Y=2.085 $X2=2.98 $Y2=2.395
r42 1 10 150 $w=1.7e-07 $l=8.00125e-07 $layer=licon1_PDIFF $count=4 $X=0.66
+ $Y=2.085 $X2=1.32 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%X 1 2 7 8 9 10 11 18
r14 11 33 16.3939 $w=3.53e-07 $l=5.05e-07 $layer=LI1_cond $X=3.577 $Y=2.405
+ $X2=3.577 $Y2=2.91
r15 11 29 5.68106 $w=3.53e-07 $l=1.75e-07 $layer=LI1_cond $X=3.577 $Y=2.405
+ $X2=3.577 $Y2=2.23
r16 10 29 6.33032 $w=3.53e-07 $l=1.95e-07 $layer=LI1_cond $X=3.577 $Y=2.035
+ $X2=3.577 $Y2=2.23
r17 9 10 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.577 $Y=1.665
+ $X2=3.577 $Y2=2.035
r18 8 9 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.577 $Y=1.295
+ $X2=3.577 $Y2=1.665
r19 7 8 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.577 $Y=0.925
+ $X2=3.577 $Y2=1.295
r20 7 18 6.65495 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=3.577 $Y=0.925
+ $X2=3.577 $Y2=0.72
r21 2 33 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=2.085 $X2=3.51 $Y2=2.91
r22 2 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=2.085 $X2=3.51 $Y2=2.23
r23 1 18 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.465 $X2=3.51 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%VGND 1 2 9 13 15 17 22 29 30 33 36
r40 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r43 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 27 36 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.717
+ $Y2=0
r45 27 29 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.6
+ $Y2=0
r46 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r47 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 23 33 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.235
+ $Y2=0
r49 23 25 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=2.16
+ $Y2=0
r50 22 36 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.717
+ $Y2=0
r51 22 25 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.16
+ $Y2=0
r52 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r53 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 17 33 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.235
+ $Y2=0
r55 17 19 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.72
+ $Y2=0
r56 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r57 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r58 11 36 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.717 $Y=0.085
+ $X2=2.717 $Y2=0
r59 11 13 21.8448 $w=3.33e-07 $l=6.35e-07 $layer=LI1_cond $X=2.717 $Y=0.085
+ $X2=2.717 $Y2=0.72
r60 7 33 2.80049 $w=6.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r61 7 9 10.3777 $w=6.78e-07 $l=5.9e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.675
r62 2 13 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.465 $X2=2.72 $Y2=0.72
r63 1 9 91 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.465 $X2=1.41 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0P_LP2%VPWR 1 8 14
r28 5 14 0.00390625 $w=3.84e-06 $l=1.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.92 $Y2=3.21
r29 5 8 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r30 4 8 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=3.6
+ $Y2=3.33
r31 4 5 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 1 14 9.76563e-05 $w=3.84e-06 $l=3e-09 $layer=MET1_cond $X=1.92 $Y=3.207
+ $X2=1.92 $Y2=3.21
.ends

