* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o31ai_m A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_226_535# A2 a_154_535# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1001 Y A3 a_226_535# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1002 a_154_535# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.74e+06u
M1003 a_126_129# A3 VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=2.289e+11p ps=2.77e+06u
M1004 Y B1 a_126_129# VNB nshort w=420000u l=150000u
+  ad=1.449e+11p pd=1.53e+06u as=0p ps=0u
M1005 VGND A2 a_126_129# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_126_129# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
