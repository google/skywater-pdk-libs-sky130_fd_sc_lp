* NGSPICE file created from sky130_fd_sc_lp__o32a_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_355_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=1.449e+12p ps=9.86e+06u
M1001 a_341_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=7.224e+11p pd=6.76e+06u as=1.1634e+12p ps=7.81e+06u
M1002 VPWR B1 a_643_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=4.914e+11p ps=3.3e+06u
M1003 a_341_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A2 a_341_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_85_21# A3 a_427_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.914e+11p pd=3.3e+06u as=4.914e+11p ps=3.3e+06u
M1006 X a_85_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1007 a_341_47# B1 a_85_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.32e+06u
M1008 a_427_367# A2 a_355_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_85_21# B2 a_341_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_643_367# B2 a_85_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_85_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1012 VPWR a_85_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_85_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

