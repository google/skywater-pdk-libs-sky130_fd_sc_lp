* File: sky130_fd_sc_lp__or3_0.spice
* Created: Wed Sep  2 10:30:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3_0.pex.spice"
.subckt sky130_fd_sc_lp__or3_0  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_29_55#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1575 AS=0.1113 PD=1.17 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_29_55#_M1007_d N_B_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1575 PD=0.7 PS=1.17 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_29_55#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_29_55#_M1006_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1281 AS=0.0588 PD=1.45 PS=0.7 NRD=11.424 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_191_481# N_C_M1000_g N_A_29_55#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 A_263_481# N_B_M1002_g A_191_481# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_263_481# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.128021 AS=0.0441 PD=0.998491 PS=0.63 NRD=80.9079 NRS=23.443 M=1 R=2.8
+ SA=75000.9 SB=75001 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_29_55#_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.195079 PD=1.81 PS=1.52151 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__or3_0.pxi.spice"
*
.ends
*
*
