* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__maj3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_275_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_275_391# B a_30_57# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_30_57# B a_479_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND A a_315_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_117_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_30_57# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_30_57# B a_479_389# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_479_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_30_57# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_117_391# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_479_389# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_315_57# B a_30_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_30_57# C a_117_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_30_57# C a_117_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
