* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41oi_lp A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_326_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A3 a_27_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VPWR A1 a_27_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 Y B1 a_514_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_409# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_27_409# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_514_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_170_47# A3 a_248_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_27_409# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_248_47# A2 a_326_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND A4 a_170_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
