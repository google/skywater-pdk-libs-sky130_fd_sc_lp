* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4bb_m A_N B_N C D VGND VNB VPB VPWR X
X0 a_332_125# a_223_55# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_332_125# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR B_N a_223_55# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_54_55# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_415_125# a_223_55# a_487_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_595_125# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_332_125# a_54_55# a_415_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_332_125# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_54_55# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_487_125# C a_595_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_54_55# a_332_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_332_125# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VGND B_N a_223_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR C a_332_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
