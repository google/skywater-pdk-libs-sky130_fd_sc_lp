* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32a_lp A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_31_101# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_134_101# A3 a_376_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_151_419# B2 a_134_101# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_376_419# A2 a_474_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VPWR a_134_101# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_31_101# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_134_101# a_612_89# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_474_419# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VGND A2 a_31_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_31_101# B1 a_134_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_134_101# B2 a_31_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR B1 a_151_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_612_89# a_134_101# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
