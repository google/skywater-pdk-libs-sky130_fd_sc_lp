* File: sky130_fd_sc_lp__nand3_0.pxi.spice
* Created: Wed Sep  2 10:04:02 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3_0%C N_C_c_45_n N_C_M1001_g N_C_M1000_g N_C_c_47_n
+ N_C_c_48_n N_C_c_53_n C C C C N_C_c_50_n PM_SKY130_FD_SC_LP__NAND3_0%C
x_PM_SKY130_FD_SC_LP__NAND3_0%B N_B_M1004_g N_B_M1003_g B B B N_B_c_84_n
+ PM_SKY130_FD_SC_LP__NAND3_0%B
x_PM_SKY130_FD_SC_LP__NAND3_0%A N_A_M1005_g N_A_M1002_g N_A_c_122_n N_A_c_123_n
+ A A A N_A_c_125_n PM_SKY130_FD_SC_LP__NAND3_0%A
x_PM_SKY130_FD_SC_LP__NAND3_0%VPWR N_VPWR_M1001_s N_VPWR_M1003_d N_VPWR_c_156_n
+ N_VPWR_c_157_n N_VPWR_c_158_n N_VPWR_c_159_n N_VPWR_c_160_n VPWR
+ N_VPWR_c_161_n N_VPWR_c_155_n PM_SKY130_FD_SC_LP__NAND3_0%VPWR
x_PM_SKY130_FD_SC_LP__NAND3_0%Y N_Y_M1005_d N_Y_M1001_d N_Y_M1002_d N_Y_c_182_n
+ N_Y_c_183_n Y Y Y N_Y_c_187_n N_Y_c_188_n N_Y_c_189_n
+ PM_SKY130_FD_SC_LP__NAND3_0%Y
x_PM_SKY130_FD_SC_LP__NAND3_0%VGND N_VGND_M1000_s N_VGND_c_223_n N_VGND_c_224_n
+ VGND N_VGND_c_225_n N_VGND_c_226_n PM_SKY130_FD_SC_LP__NAND3_0%VGND
cc_1 VNB N_C_c_45_n 0.00967017f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.77
cc_2 VNB N_C_M1000_g 0.0252447f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.445
cc_3 VNB N_C_c_47_n 0.0308874f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.99
cc_4 VNB N_C_c_48_n 0.0185661f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_5 VNB C 0.0350269f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_C_c_50_n 0.0298297f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_B_M1004_g 0.0367405f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.92
cc_8 VNB N_B_M1003_g 0.00656382f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.84
cc_9 VNB B 0.00893108f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.445
cc_10 VNB N_B_c_84_n 0.0319875f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.845
cc_11 VNB N_A_M1005_g 0.023721f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.92
cc_12 VNB N_A_M1002_g 0.00834029f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.84
cc_13 VNB N_A_c_122_n 0.0234523f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_14 VNB N_A_c_123_n 0.0166109f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.84
cc_15 VNB A 0.00970139f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.99
cc_16 VNB N_A_c_125_n 0.0165751f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_17 VNB N_VPWR_c_155_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_182_n 0.0511151f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_19 VNB N_Y_c_183_n 0.0180143f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_20 VNB N_VGND_c_223_n 0.0114569f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.63
cc_21 VNB N_VGND_c_224_n 0.0173648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_225_n 0.0431266f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_23 VNB N_VGND_c_226_n 0.129088f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.845
cc_24 VPB N_C_c_45_n 0.00775879f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.77
cc_25 VPB N_C_M1001_g 0.037398f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.63
cc_26 VPB N_C_c_53_n 0.0239576f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.845
cc_27 VPB C 0.0222776f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_28 VPB N_B_M1003_g 0.0439431f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_29 VPB B 0.00386797f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.445
cc_30 VPB N_A_M1002_g 0.0515692f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_31 VPB A 0.00358728f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.99
cc_32 VPB N_VPWR_c_156_n 0.0116772f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_33 VPB N_VPWR_c_157_n 0.0409712f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.445
cc_34 VPB N_VPWR_c_158_n 0.011379f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.99
cc_35 VPB N_VPWR_c_159_n 0.01683f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.845
cc_36 VPB N_VPWR_c_160_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_161_n 0.0198171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_155_n 0.0597606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_Y_c_182_n 0.0132955f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_40 VPB Y 0.00394514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB Y 0.0150759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_Y_c_187_n 0.00849134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_Y_c_188_n 0.00648803f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=0.925
cc_44 VPB N_Y_c_189_n 0.0424242f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.665
cc_45 N_C_M1000_g N_B_M1004_g 0.0492605f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_46 C N_B_M1004_g 2.65381e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_47 N_C_c_50_n N_B_M1004_g 0.00557585f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_48 N_C_c_45_n N_B_M1003_g 0.00553293f $X=0.36 $Y=1.77 $X2=0 $Y2=0
cc_49 N_C_c_53_n N_B_M1003_g 0.0271677f $X=0.5 $Y=1.845 $X2=0 $Y2=0
cc_50 C N_B_M1003_g 8.88572e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_51 N_C_M1000_g B 0.00162428f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_52 N_C_c_47_n B 0.00450397f $X=0.345 $Y=0.99 $X2=0 $Y2=0
cc_53 C B 0.0630964f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_54 N_C_c_50_n B 0.00615104f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_55 C N_B_c_84_n 3.10182e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_56 N_C_c_50_n N_B_c_84_n 0.0171887f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_57 N_C_M1001_g N_VPWR_c_157_n 0.00425278f $X=0.5 $Y=2.63 $X2=0 $Y2=0
cc_58 N_C_c_53_n N_VPWR_c_157_n 0.00268809f $X=0.5 $Y=1.845 $X2=0 $Y2=0
cc_59 C N_VPWR_c_157_n 0.0218313f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_60 N_C_M1001_g N_VPWR_c_159_n 0.00570944f $X=0.5 $Y=2.63 $X2=0 $Y2=0
cc_61 N_C_M1001_g N_VPWR_c_155_n 0.00542671f $X=0.5 $Y=2.63 $X2=0 $Y2=0
cc_62 N_C_M1001_g Y 0.00204032f $X=0.5 $Y=2.63 $X2=0 $Y2=0
cc_63 C Y 0.0140859f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_64 N_C_M1001_g N_Y_c_188_n 0.00493193f $X=0.5 $Y=2.63 $X2=0 $Y2=0
cc_65 N_C_M1000_g N_VGND_c_224_n 0.0139429f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_66 N_C_c_47_n N_VGND_c_224_n 0.00386217f $X=0.345 $Y=0.99 $X2=0 $Y2=0
cc_67 C N_VGND_c_224_n 0.0199694f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_68 N_C_M1000_g N_VGND_c_225_n 0.00486043f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_69 N_C_M1000_g N_VGND_c_226_n 0.00784452f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_70 C N_VGND_c_226_n 0.00276004f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_71 N_B_M1004_g N_A_M1005_g 0.0583182f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_72 B N_A_M1005_g 3.44374e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_73 N_B_c_84_n N_A_M1002_g 0.0389455f $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_74 N_B_c_84_n N_A_c_122_n 0.0191562f $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_75 N_B_M1004_g A 0.00220398f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_76 B A 0.0731345f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_77 N_B_c_84_n A 0.00378217f $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_78 B N_A_c_125_n 6.05905e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_79 N_B_M1003_g N_VPWR_c_158_n 0.00191103f $X=0.93 $Y=2.63 $X2=0 $Y2=0
cc_80 N_B_M1003_g N_VPWR_c_159_n 0.00570944f $X=0.93 $Y=2.63 $X2=0 $Y2=0
cc_81 N_B_M1003_g N_VPWR_c_155_n 0.00542671f $X=0.93 $Y=2.63 $X2=0 $Y2=0
cc_82 N_B_M1004_g N_Y_c_183_n 0.00161915f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_83 B Y 0.0238924f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_B_c_84_n Y 7.91292e-19 $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_85 N_B_M1003_g N_Y_c_187_n 0.0184271f $X=0.93 $Y=2.63 $X2=0 $Y2=0
cc_86 B N_Y_c_187_n 0.00655788f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 N_B_M1003_g N_Y_c_188_n 0.00271737f $X=0.93 $Y=2.63 $X2=0 $Y2=0
cc_88 N_B_M1004_g N_VGND_c_224_n 0.00294663f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_89 N_B_M1004_g N_VGND_c_225_n 0.00585385f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_90 N_B_M1004_g N_VGND_c_226_n 0.00778255f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_91 B N_VGND_c_226_n 0.0137968f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A_M1002_g N_VPWR_c_158_n 0.00330548f $X=1.36 $Y=2.63 $X2=0 $Y2=0
cc_93 N_A_M1002_g N_VPWR_c_161_n 0.00570944f $X=1.36 $Y=2.63 $X2=0 $Y2=0
cc_94 N_A_M1002_g N_VPWR_c_155_n 0.00542671f $X=1.36 $Y=2.63 $X2=0 $Y2=0
cc_95 N_A_M1005_g N_Y_c_182_n 0.00662634f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_M1002_g N_Y_c_182_n 0.0071756f $X=1.36 $Y=2.63 $X2=0 $Y2=0
cc_97 A N_Y_c_182_n 0.0706474f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_98 N_A_c_125_n N_Y_c_182_n 0.0163177f $X=1.38 $Y=1.005 $X2=0 $Y2=0
cc_99 N_A_M1005_g N_Y_c_183_n 0.0067103f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_100 A N_Y_c_183_n 0.00633558f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_101 N_A_c_125_n N_Y_c_183_n 0.00351543f $X=1.38 $Y=1.005 $X2=0 $Y2=0
cc_102 N_A_c_123_n Y 0.00279892f $X=1.38 $Y=1.51 $X2=0 $Y2=0
cc_103 A Y 0.00318565f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_104 N_A_M1002_g N_Y_c_187_n 0.0181842f $X=1.36 $Y=2.63 $X2=0 $Y2=0
cc_105 N_A_c_123_n N_Y_c_187_n 3.04466e-19 $X=1.38 $Y=1.51 $X2=0 $Y2=0
cc_106 A N_Y_c_187_n 0.0280855f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_107 N_A_M1002_g N_Y_c_189_n 0.00623196f $X=1.36 $Y=2.63 $X2=0 $Y2=0
cc_108 N_A_M1005_g N_VGND_c_225_n 0.0054833f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_M1005_g N_VGND_c_226_n 0.0073966f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_110 A N_VGND_c_226_n 0.00892327f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_111 N_VPWR_c_158_n N_Y_c_187_n 0.0220348f $X=1.145 $Y=2.455 $X2=0 $Y2=0
cc_112 N_VPWR_c_157_n N_Y_c_188_n 0.00307479f $X=0.285 $Y=2.455 $X2=0 $Y2=0
cc_113 N_VPWR_c_158_n N_Y_c_188_n 0.00304534f $X=1.145 $Y=2.455 $X2=0 $Y2=0
cc_114 N_VPWR_c_159_n N_Y_c_188_n 0.0108533f $X=1.01 $Y=3.33 $X2=0 $Y2=0
cc_115 N_VPWR_c_155_n N_Y_c_188_n 0.00928771f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_116 N_VPWR_c_158_n N_Y_c_189_n 0.00314943f $X=1.145 $Y=2.455 $X2=0 $Y2=0
cc_117 N_VPWR_c_161_n N_Y_c_189_n 0.0168591f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_118 N_VPWR_c_155_n N_Y_c_189_n 0.0144272f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_119 N_Y_c_183_n N_VGND_c_225_n 0.0269737f $X=1.74 $Y=0.445 $X2=0 $Y2=0
cc_120 N_Y_M1005_d N_VGND_c_226_n 0.0021695f $X=1.365 $Y=0.235 $X2=0 $Y2=0
cc_121 N_Y_c_183_n N_VGND_c_226_n 0.0185031f $X=1.74 $Y=0.445 $X2=0 $Y2=0
cc_122 N_VGND_c_226_n A_117_47# 0.00330251f $X=1.68 $Y=0 $X2=-0.19 $Y2=-0.245
cc_123 N_VGND_c_226_n A_195_47# 0.00692683f $X=1.68 $Y=0 $X2=-0.19 $Y2=-0.245
