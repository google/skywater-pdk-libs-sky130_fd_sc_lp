* File: sky130_fd_sc_lp__sdfstp_4.pxi.spice
* Created: Fri Aug 28 11:29:51 2020
* 
x_PM_SKY130_FD_SC_LP__SDFSTP_4%SCD N_SCD_M1038_g N_SCD_c_286_n N_SCD_M1014_g
+ N_SCD_c_287_n N_SCD_c_288_n SCD SCD N_SCD_c_289_n N_SCD_c_290_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%SCD
x_PM_SKY130_FD_SC_LP__SDFSTP_4%D N_D_M1017_g N_D_M1013_g N_D_c_323_n D D D D D
+ N_D_c_327_n N_D_c_324_n D N_D_c_330_n PM_SKY130_FD_SC_LP__SDFSTP_4%D
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_346_93# N_A_346_93#_M1001_d N_A_346_93#_M1039_d
+ N_A_346_93#_M1000_g N_A_346_93#_M1031_g N_A_346_93#_c_382_n
+ N_A_346_93#_c_383_n N_A_346_93#_c_377_n N_A_346_93#_c_378_n
+ N_A_346_93#_c_379_n N_A_346_93#_c_386_n N_A_346_93#_c_387_n
+ N_A_346_93#_c_388_n PM_SKY130_FD_SC_LP__SDFSTP_4%A_346_93#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%SCE N_SCE_M1012_g N_SCE_M1009_g N_SCE_c_452_n
+ N_SCE_c_453_n N_SCE_M1001_g N_SCE_c_455_n N_SCE_c_465_n N_SCE_M1039_g
+ N_SCE_c_456_n N_SCE_c_457_n N_SCE_c_458_n N_SCE_c_468_n N_SCE_c_459_n
+ N_SCE_c_460_n N_SCE_c_461_n SCE SCE SCE SCE N_SCE_c_463_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%SCE
x_PM_SKY130_FD_SC_LP__SDFSTP_4%CLK N_CLK_c_552_n N_CLK_M1042_g N_CLK_M1037_g
+ N_CLK_c_555_n CLK CLK CLK N_CLK_c_557_n PM_SKY130_FD_SC_LP__SDFSTP_4%CLK
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_961_491# N_A_961_491#_M1005_d
+ N_A_961_491#_M1023_d N_A_961_491#_M1033_g N_A_961_491#_M1008_g
+ N_A_961_491#_M1035_g N_A_961_491#_M1026_g N_A_961_491#_c_607_n
+ N_A_961_491#_c_599_n N_A_961_491#_c_600_n N_A_961_491#_c_664_p
+ N_A_961_491#_c_608_n N_A_961_491#_c_609_n N_A_961_491#_c_610_n
+ N_A_961_491#_c_611_n N_A_961_491#_c_612_n N_A_961_491#_c_613_n
+ N_A_961_491#_c_614_n N_A_961_491#_c_615_n N_A_961_491#_c_616_n
+ N_A_961_491#_c_628_p N_A_961_491#_c_601_n N_A_961_491#_c_602_n
+ N_A_961_491#_c_702_p N_A_961_491#_c_617_n N_A_961_491#_c_618_n
+ N_A_961_491#_c_603_n N_A_961_491#_c_620_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_961_491#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_1339_331# N_A_1339_331#_M1027_s
+ N_A_1339_331#_M1029_d N_A_1339_331#_M1025_g N_A_1339_331#_M1011_g
+ N_A_1339_331#_c_787_n N_A_1339_331#_c_780_n N_A_1339_331#_c_781_n
+ N_A_1339_331#_c_782_n N_A_1339_331#_c_789_n N_A_1339_331#_c_783_n
+ N_A_1339_331#_c_784_n N_A_1339_331#_c_785_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_1339_331#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_1211_463# N_A_1211_463#_M1041_d
+ N_A_1211_463#_M1033_d N_A_1211_463#_M1029_g N_A_1211_463#_c_850_n
+ N_A_1211_463#_M1027_g N_A_1211_463#_M1010_g N_A_1211_463#_c_852_n
+ N_A_1211_463#_c_853_n N_A_1211_463#_M1028_g N_A_1211_463#_c_854_n
+ N_A_1211_463#_c_862_n N_A_1211_463#_c_863_n N_A_1211_463#_c_855_n
+ N_A_1211_463#_c_895_n N_A_1211_463#_c_856_n N_A_1211_463#_c_857_n
+ N_A_1211_463#_c_858_n N_A_1211_463#_c_859_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_1211_463#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%SET_B N_SET_B_M1018_g N_SET_B_c_974_n
+ N_SET_B_c_975_n N_SET_B_c_966_n N_SET_B_M1032_g N_SET_B_M1024_g
+ N_SET_B_M1003_g N_SET_B_c_969_n N_SET_B_c_978_n N_SET_B_c_970_n
+ N_SET_B_c_971_n N_SET_B_c_972_n SET_B SET_B SET_B SET_B SET_B
+ PM_SKY130_FD_SC_LP__SDFSTP_4%SET_B
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_773_409# N_A_773_409#_M1037_s
+ N_A_773_409#_M1042_s N_A_773_409#_M1023_g N_A_773_409#_M1005_g
+ N_A_773_409#_c_1064_n N_A_773_409#_c_1065_n N_A_773_409#_c_1075_n
+ N_A_773_409#_c_1076_n N_A_773_409#_c_1077_n N_A_773_409#_c_1078_n
+ N_A_773_409#_c_1066_n N_A_773_409#_M1041_g N_A_773_409#_M1022_g
+ N_A_773_409#_c_1080_n N_A_773_409#_M1002_g N_A_773_409#_c_1067_n
+ N_A_773_409#_c_1068_n N_A_773_409#_M1020_g N_A_773_409#_c_1084_n
+ N_A_773_409#_c_1085_n N_A_773_409#_c_1070_n N_A_773_409#_c_1071_n
+ N_A_773_409#_c_1088_n N_A_773_409#_c_1089_n N_A_773_409#_c_1072_n
+ N_A_773_409#_c_1073_n PM_SKY130_FD_SC_LP__SDFSTP_4%A_773_409#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_2205_231# N_A_2205_231#_M1043_d
+ N_A_2205_231#_M1015_d N_A_2205_231#_M1016_g N_A_2205_231#_M1019_g
+ N_A_2205_231#_c_1228_n N_A_2205_231#_c_1229_n N_A_2205_231#_c_1230_n
+ N_A_2205_231#_c_1231_n N_A_2205_231#_c_1232_n N_A_2205_231#_c_1233_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_2205_231#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_1960_125# N_A_1960_125#_M1035_d
+ N_A_1960_125#_M1026_d N_A_1960_125#_M1003_d N_A_1960_125#_M1043_g
+ N_A_1960_125#_c_1283_n N_A_1960_125#_M1015_g N_A_1960_125#_c_1284_n
+ N_A_1960_125#_M1007_g N_A_1960_125#_c_1291_n N_A_1960_125#_M1040_g
+ N_A_1960_125#_c_1286_n N_A_1960_125#_c_1293_n N_A_1960_125#_c_1287_n
+ N_A_1960_125#_c_1295_n N_A_1960_125#_c_1296_n N_A_1960_125#_c_1297_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_1960_125#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_2638_53# N_A_2638_53#_M1007_s
+ N_A_2638_53#_M1040_s N_A_2638_53#_M1004_g N_A_2638_53#_M1006_g
+ N_A_2638_53#_M1030_g N_A_2638_53#_M1021_g N_A_2638_53#_M1036_g
+ N_A_2638_53#_M1034_g N_A_2638_53#_M1045_g N_A_2638_53#_M1044_g
+ N_A_2638_53#_c_1384_n N_A_2638_53#_c_1392_n N_A_2638_53#_c_1385_n
+ N_A_2638_53#_c_1386_n N_A_2638_53#_c_1387_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_2638_53#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_27_479# N_A_27_479#_M1038_s N_A_27_479#_M1031_d
+ N_A_27_479#_c_1485_n N_A_27_479#_c_1486_n N_A_27_479#_c_1487_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_27_479#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%VPWR N_VPWR_M1038_d N_VPWR_M1039_s N_VPWR_M1042_d
+ N_VPWR_M1025_d N_VPWR_M1018_d N_VPWR_M1019_d N_VPWR_M1015_s N_VPWR_M1040_d
+ N_VPWR_M1021_d N_VPWR_M1044_d N_VPWR_c_1513_n N_VPWR_c_1514_n N_VPWR_c_1515_n
+ N_VPWR_c_1516_n N_VPWR_c_1517_n N_VPWR_c_1518_n N_VPWR_c_1519_n
+ N_VPWR_c_1520_n N_VPWR_c_1521_n N_VPWR_c_1522_n N_VPWR_c_1523_n
+ N_VPWR_c_1524_n N_VPWR_c_1525_n N_VPWR_c_1526_n N_VPWR_c_1527_n
+ N_VPWR_c_1528_n N_VPWR_c_1529_n VPWR N_VPWR_c_1530_n N_VPWR_c_1531_n
+ N_VPWR_c_1532_n N_VPWR_c_1533_n N_VPWR_c_1534_n N_VPWR_c_1535_n
+ N_VPWR_c_1536_n N_VPWR_c_1537_n N_VPWR_c_1538_n N_VPWR_c_1539_n
+ N_VPWR_c_1540_n N_VPWR_c_1541_n N_VPWR_c_1542_n N_VPWR_c_1512_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%VPWR
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_218_119# N_A_218_119#_M1009_d
+ N_A_218_119#_M1041_s N_A_218_119#_M1017_d N_A_218_119#_M1033_s
+ N_A_218_119#_c_1713_n N_A_218_119#_c_1697_n N_A_218_119#_c_1698_n
+ N_A_218_119#_c_1702_n N_A_218_119#_c_1703_n N_A_218_119#_c_1699_n
+ N_A_218_119#_c_1705_n N_A_218_119#_c_1706_n N_A_218_119#_c_1763_n
+ N_A_218_119#_c_1707_n N_A_218_119#_c_1708_n N_A_218_119#_c_1752_n
+ N_A_218_119#_c_1709_n N_A_218_119#_c_1710_n N_A_218_119#_c_1700_n
+ N_A_218_119#_c_1712_n N_A_218_119#_c_1701_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_218_119#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_1751_379# N_A_1751_379#_M1010_d
+ N_A_1751_379#_M1002_d N_A_1751_379#_c_1843_n N_A_1751_379#_c_1840_n
+ N_A_1751_379#_c_1841_n PM_SKY130_FD_SC_LP__SDFSTP_4%A_1751_379#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%A_1858_463# N_A_1858_463#_M1026_s
+ N_A_1858_463#_M1019_s N_A_1858_463#_c_1870_n N_A_1858_463#_c_1871_n
+ PM_SKY130_FD_SC_LP__SDFSTP_4%A_1858_463#
x_PM_SKY130_FD_SC_LP__SDFSTP_4%Q N_Q_M1004_s N_Q_M1036_s N_Q_M1006_s N_Q_M1034_s
+ N_Q_c_1931_n N_Q_c_1889_n N_Q_c_1890_n N_Q_c_1891_n N_Q_c_1895_n N_Q_c_1896_n
+ N_Q_c_1892_n N_Q_c_1936_n N_Q_c_1897_n Q Q PM_SKY130_FD_SC_LP__SDFSTP_4%Q
x_PM_SKY130_FD_SC_LP__SDFSTP_4%VGND N_VGND_M1014_s N_VGND_M1000_d N_VGND_M1037_d
+ N_VGND_M1011_d N_VGND_M1032_d N_VGND_M1024_d N_VGND_M1007_d N_VGND_M1030_d
+ N_VGND_M1045_d N_VGND_c_1953_n N_VGND_c_1954_n N_VGND_c_1955_n N_VGND_c_1956_n
+ N_VGND_c_1957_n N_VGND_c_1958_n N_VGND_c_1959_n N_VGND_c_1960_n
+ N_VGND_c_1961_n N_VGND_c_1962_n N_VGND_c_1963_n N_VGND_c_1964_n
+ N_VGND_c_1965_n N_VGND_c_1966_n N_VGND_c_1967_n N_VGND_c_1968_n VGND
+ N_VGND_c_1969_n N_VGND_c_1970_n N_VGND_c_1971_n N_VGND_c_1972_n
+ N_VGND_c_1973_n N_VGND_c_1974_n N_VGND_c_1975_n N_VGND_c_1976_n
+ N_VGND_c_1977_n N_VGND_c_1978_n N_VGND_c_1979_n N_VGND_c_1980_n
+ N_VGND_c_1981_n N_VGND_c_1982_n PM_SKY130_FD_SC_LP__SDFSTP_4%VGND
cc_1 VNB N_SCD_c_286_n 0.0210117f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.125
cc_2 VNB N_SCD_c_287_n 0.0325633f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.2
cc_3 VNB N_SCD_c_288_n 0.00205046f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.795
cc_4 VNB N_SCD_c_289_n 0.0301776f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_5 VNB N_SCD_c_290_n 0.0254176f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_6 VNB N_D_M1013_g 0.0242263f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_7 VNB N_D_c_323_n 0.00757936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D_c_324_n 0.00688124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_346_93#_M1000_g 0.0455458f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_10 VNB N_A_346_93#_c_377_n 0.0174107f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_11 VNB N_A_346_93#_c_378_n 0.00827725f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_12 VNB N_A_346_93#_c_379_n 0.0439437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_M1009_g 0.0491807f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.2
cc_14 VNB N_SCE_c_452_n 0.0765232f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_15 VNB N_SCE_c_453_n 0.0125466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_M1001_g 0.041559f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.63
cc_17 VNB N_SCE_c_455_n 0.0988678f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_SCE_c_456_n 0.0317385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_SCE_c_457_n 0.0167577f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_20 VNB N_SCE_c_458_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_459_n 0.0152377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_460_n 0.0294732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_461_n 0.0212061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB SCE 0.00524288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_SCE_c_463_n 0.0236731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_CLK_c_552_n 0.0183586f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.795
cc_27 VNB N_CLK_M1042_g 0.00836477f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.715
cc_28 VNB N_CLK_M1037_g 0.0205583f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.805
cc_29 VNB N_CLK_c_555_n 0.0255043f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.2
cc_30 VNB CLK 0.0115811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_CLK_c_557_n 0.0161151f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_32 VNB N_A_961_491#_M1008_g 0.0349625f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.63
cc_33 VNB N_A_961_491#_M1035_g 0.0343851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_961_491#_c_599_n 0.0152493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_961_491#_c_600_n 0.00104173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_961_491#_c_601_n 0.00223031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_961_491#_c_602_n 0.0048558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_961_491#_c_603_n 0.0690268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1339_331#_c_780_n 0.0041882f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_40 VNB N_A_1339_331#_c_781_n 0.021395f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_41 VNB N_A_1339_331#_c_782_n 0.0353113f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.295
cc_42 VNB N_A_1339_331#_c_783_n 0.00313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1339_331#_c_784_n 0.0209196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1339_331#_c_785_n 0.0188105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1211_463#_M1029_g 0.00268514f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_46 VNB N_A_1211_463#_c_850_n 0.0200942f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.2
cc_47 VNB N_A_1211_463#_M1027_g 0.0259334f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_48 VNB N_A_1211_463#_c_852_n 0.0303559f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_49 VNB N_A_1211_463#_c_853_n 0.0194881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1211_463#_c_854_n 0.00757723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1211_463#_c_855_n 7.80901e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1211_463#_c_856_n 0.00794761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1211_463#_c_857_n 0.0328202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1211_463#_c_858_n 0.0340297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1211_463#_c_859_n 0.0262469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_SET_B_c_966_n 0.05499f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.805
cc_57 VNB N_SET_B_M1032_g 0.043527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_M1024_g 0.035414f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.63
cc_59 VNB N_SET_B_c_969_n 0.00446475f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_60 VNB N_SET_B_c_970_n 0.00929652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_SET_B_c_971_n 0.0139266f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_62 VNB N_SET_B_c_972_n 0.0418803f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_63 VNB N_A_773_409#_M1005_g 0.0269604f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.63
cc_64 VNB N_A_773_409#_c_1064_n 0.0812553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_773_409#_c_1065_n 0.0144833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_773_409#_c_1066_n 0.0191538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_773_409#_c_1067_n 0.0193632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_773_409#_c_1068_n 0.00983532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_773_409#_M1020_g 0.0331426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_773_409#_c_1070_n 0.00533974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_773_409#_c_1071_n 0.0180962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_773_409#_c_1072_n 0.00486811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_773_409#_c_1073_n 0.0359318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_2205_231#_M1019_g 0.00856611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_2205_231#_c_1228_n 0.0210455f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.795
cc_76 VNB N_A_2205_231#_c_1229_n 0.0332599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_2205_231#_c_1230_n 0.0264134f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_78 VNB N_A_2205_231#_c_1231_n 0.0109283f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_79 VNB N_A_2205_231#_c_1232_n 0.00319433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_2205_231#_c_1233_n 0.0179223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1960_125#_M1043_g 0.0484158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1960_125#_c_1283_n 0.0150987f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.795
cc_83 VNB N_A_1960_125#_c_1284_n 0.0290609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1960_125#_M1007_g 0.0392339f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.29
cc_85 VNB N_A_1960_125#_c_1286_n 0.00362067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1960_125#_c_1287_n 0.00807407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2638_53#_M1004_g 0.0228903f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_88 VNB N_A_2638_53#_M1030_g 0.0213867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2638_53#_M1036_g 0.0213652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2638_53#_M1045_g 0.0262458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2638_53#_c_1384_n 0.0335089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2638_53#_c_1385_n 0.00521674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2638_53#_c_1386_n 0.00324131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2638_53#_c_1387_n 0.0721789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VPWR_c_1512_n 0.661241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_218_119#_c_1697_n 0.0326239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_218_119#_c_1698_n 0.00251249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_218_119#_c_1699_n 0.00239036f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.295
cc_99 VNB N_A_218_119#_c_1700_n 0.0166265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_218_119#_c_1701_n 0.00287881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_Q_c_1889_n 0.0015362f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_102 VNB N_Q_c_1890_n 0.00320529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_Q_c_1891_n 0.00304786f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_104 VNB N_Q_c_1892_n 0.0015362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB Q 0.0119302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB Q 0.019342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1953_n 0.0383409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1954_n 0.00831555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1955_n 0.00653261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1956_n 0.0210438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1957_n 0.016308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1958_n 0.00105389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1959_n 0.00828717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1960_n 0.031794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1961_n 0.00403121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1962_n 7.97178e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1963_n 0.0142614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1964_n 0.0291522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1965_n 0.0108943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1966_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1967_n 0.0223217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1968_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1969_n 0.0372213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1970_n 0.0618353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1971_n 0.0589607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1972_n 0.0906641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1973_n 0.0434415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1974_n 0.0133348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1975_n 0.0133348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1976_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1977_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1978_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1979_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1980_n 0.00476075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1981_n 0.00476075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1982_n 0.887509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VPB N_SCD_M1038_g 0.0556934f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.715
cc_138 VPB N_SCD_c_288_n 0.0169143f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.795
cc_139 VPB N_SCD_c_290_n 0.00553174f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_140 VPB N_D_M1017_g 0.0193167f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.715
cc_141 VPB D 0.020374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_D_c_327_n 0.0286158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_D_c_324_n 0.013415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB D 0.0194795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_D_c_330_n 0.00477283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_346_93#_M1000_g 0.00620135f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_147 VPB N_A_346_93#_M1031_g 0.0427292f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.63
cc_148 VPB N_A_346_93#_c_382_n 0.0725692f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_149 VPB N_A_346_93#_c_383_n 0.00491573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_346_93#_c_378_n 5.20702e-19 $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_151 VPB N_A_346_93#_c_379_n 0.00816673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_346_93#_c_386_n 0.0197065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_346_93#_c_387_n 0.00471757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_346_93#_c_388_n 0.00988152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_SCE_M1012_g 0.0450281f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.715
cc_156 VPB N_SCE_c_465_n 0.0228696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_SCE_c_456_n 0.0301333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_SCE_c_457_n 0.00429693f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_159 VPB N_SCE_c_468_n 0.0293059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB SCE 0.00395404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_CLK_M1042_g 0.0607318f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.715
cc_162 VPB CLK 0.00639381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_961_491#_M1033_g 0.0316187f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_164 VPB N_A_961_491#_M1035_g 0.00850255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_961_491#_M1026_g 0.0276457f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_166 VPB N_A_961_491#_c_607_n 0.0150543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_961_491#_c_608_n 0.00353162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_961_491#_c_609_n 0.0105088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_961_491#_c_610_n 8.35868e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_961_491#_c_611_n 0.0145974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_961_491#_c_612_n 0.0034399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_961_491#_c_613_n 7.80494e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_961_491#_c_614_n 0.0115411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_961_491#_c_615_n 0.0023525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_961_491#_c_616_n 0.00379662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_961_491#_c_617_n 7.47086e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_961_491#_c_618_n 0.0198763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_961_491#_c_603_n 0.0592605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_961_491#_c_620_n 0.0504438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1339_331#_M1025_g 0.0290101f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.275
cc_181 VPB N_A_1339_331#_c_787_n 0.0131277f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_182 VPB N_A_1339_331#_c_780_n 0.0317235f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_183 VPB N_A_1339_331#_c_789_n 0.00671821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1211_463#_M1029_g 0.0453172f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.275
cc_185 VPB N_A_1211_463#_M1010_g 0.0233775f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_186 VPB N_A_1211_463#_c_862_n 0.00113714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1211_463#_c_863_n 0.00432117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1211_463#_c_859_n 0.00850748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_SET_B_M1018_g 0.0373144f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.715
cc_190 VPB N_SET_B_c_974_n 0.0214462f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.125
cc_191 VPB N_SET_B_c_975_n 0.00845722f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=0.805
cc_192 VPB N_SET_B_M1032_g 9.04807e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_SET_B_M1003_g 0.0540476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_SET_B_c_978_n 3.7562e-19 $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_195 VPB N_SET_B_c_970_n 0.00587837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_SET_B_c_971_n 0.0156757f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.295
cc_197 VPB N_A_773_409#_M1023_g 0.0207113f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_198 VPB N_A_773_409#_c_1075_n 0.0272656f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_199 VPB N_A_773_409#_c_1076_n 0.0478741f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.29
cc_200 VPB N_A_773_409#_c_1077_n 0.0700111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_773_409#_c_1078_n 0.0098971f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.295
cc_202 VPB N_A_773_409#_M1022_g 0.030607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_773_409#_c_1080_n 0.316034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_773_409#_M1002_g 0.0184764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_773_409#_c_1067_n 0.00571568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_773_409#_c_1068_n 0.00130694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_773_409#_c_1084_n 0.0712704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_773_409#_c_1085_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_773_409#_c_1070_n 0.00126008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_773_409#_c_1071_n 0.0121394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_773_409#_c_1088_n 0.0136486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_773_409#_c_1089_n 0.0272956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_773_409#_c_1073_n 0.0205949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_2205_231#_M1019_g 0.0607266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_2205_231#_c_1232_n 0.019085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1960_125#_c_1283_n 0.0703092f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.795
cc_217 VPB N_A_1960_125#_M1015_g 0.0229525f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_218 VPB N_A_1960_125#_c_1284_n 0.0266317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1960_125#_c_1291_n 0.0194818f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.295
cc_220 VPB N_A_1960_125#_c_1286_n 0.0026819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_1960_125#_c_1293_n 0.00231006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_1960_125#_c_1287_n 0.00560889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_1960_125#_c_1295_n 0.0216409f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1960_125#_c_1296_n 0.0172378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1960_125#_c_1297_n 0.0130474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_2638_53#_M1006_g 0.0190324f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.63
cc_227 VPB N_A_2638_53#_M1021_g 0.0179096f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_228 VPB N_A_2638_53#_M1034_g 0.0178867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_2638_53#_M1044_g 0.0215411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_2638_53#_c_1392_n 0.0154541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_2638_53#_c_1387_n 0.0138076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_27_479#_c_1485_n 0.0227749f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_233 VPB N_A_27_479#_c_1486_n 0.0103825f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.2
cc_234 VPB N_A_27_479#_c_1487_n 0.00955727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1513_n 0.00203383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1514_n 0.00654408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1515_n 0.00239351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1516_n 0.0521466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1517_n 0.00956215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1518_n 0.0136035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1519_n 0.00732807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1520_n 0.019412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1521_n 0.0180353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1522_n 0.00727196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1523_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1524_n 0.0130511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1525_n 0.0412014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1526_n 0.0457167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1527_n 0.00401372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1528_n 0.0684221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1529_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1530_n 0.0159091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1531_n 0.0347933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1532_n 0.0302021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1533_n 0.0311697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1534_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1535_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1536_n 0.00510102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1537_n 0.00375621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1538_n 0.00250432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1539_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1540_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1541_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1542_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1512_n 0.103928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_218_119#_c_1702_n 0.0135244f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.29
cc_267 VPB N_A_218_119#_c_1703_n 0.00872032f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.29
cc_268 VPB N_A_218_119#_c_1699_n 0.0155095f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.295
cc_269 VPB N_A_218_119#_c_1705_n 0.00709585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_218_119#_c_1706_n 0.00729732f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.665
cc_271 VPB N_A_218_119#_c_1707_n 0.0136194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_218_119#_c_1708_n 0.00133753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_218_119#_c_1709_n 0.00509263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_218_119#_c_1710_n 4.9691e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_218_119#_c_1700_n 0.0180174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_218_119#_c_1712_n 0.00304074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_1751_379#_c_1840_n 0.00343151f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.21
cc_278 VPB N_A_1751_379#_c_1841_n 0.0127575f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_279 VPB N_A_1858_463#_c_1870_n 0.0104242f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.275
cc_280 VPB N_A_1858_463#_c_1871_n 0.00875105f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.795
cc_281 VPB N_Q_c_1895_n 0.00320221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_Q_c_1896_n 0.00260607f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_283 VPB N_Q_c_1897_n 0.00965916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB Q 0.00598624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 N_SCD_M1038_g D 0.0141927f $X=0.475 $Y=2.715 $X2=0 $Y2=0
cc_286 N_SCD_c_287_n D 0.00422265f $X=0.655 $Y=1.2 $X2=0 $Y2=0
cc_287 N_SCD_c_288_n D 0.00486318f $X=0.385 $Y=1.795 $X2=0 $Y2=0
cc_288 N_SCD_c_290_n D 0.0374759f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_289 N_SCD_M1038_g N_D_c_330_n 0.0017625f $X=0.475 $Y=2.715 $X2=0 $Y2=0
cc_290 N_SCD_c_287_n N_D_c_330_n 2.81031e-19 $X=0.655 $Y=1.2 $X2=0 $Y2=0
cc_291 N_SCD_c_288_n N_SCE_M1012_g 0.0517403f $X=0.385 $Y=1.795 $X2=0 $Y2=0
cc_292 N_SCD_c_290_n N_SCE_M1012_g 6.20955e-19 $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_293 N_SCD_c_286_n N_SCE_M1009_g 0.0483781f $X=0.655 $Y=1.125 $X2=0 $Y2=0
cc_294 N_SCD_c_289_n N_SCE_M1009_g 0.00670961f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_295 N_SCD_c_290_n N_SCE_M1009_g 0.00123789f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_296 N_SCD_c_289_n N_SCE_c_457_n 0.00824046f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_297 N_SCD_c_290_n N_SCE_c_457_n 9.52378e-19 $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_298 N_SCD_M1038_g N_A_27_479#_c_1485_n 2.21843e-19 $X=0.475 $Y=2.715 $X2=0
+ $Y2=0
cc_299 N_SCD_M1038_g N_A_27_479#_c_1486_n 0.0109678f $X=0.475 $Y=2.715 $X2=0
+ $Y2=0
cc_300 N_SCD_M1038_g N_VPWR_c_1513_n 0.0104114f $X=0.475 $Y=2.715 $X2=0 $Y2=0
cc_301 N_SCD_M1038_g N_VPWR_c_1530_n 0.00437283f $X=0.475 $Y=2.715 $X2=0 $Y2=0
cc_302 N_SCD_M1038_g N_VPWR_c_1512_n 0.00487376f $X=0.475 $Y=2.715 $X2=0 $Y2=0
cc_303 N_SCD_c_286_n N_A_218_119#_c_1713_n 0.00201294f $X=0.655 $Y=1.125 $X2=0
+ $Y2=0
cc_304 N_SCD_c_290_n N_A_218_119#_c_1713_n 0.00232057f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_305 N_SCD_c_287_n N_A_218_119#_c_1698_n 2.03909e-19 $X=0.655 $Y=1.2 $X2=0
+ $Y2=0
cc_306 N_SCD_c_289_n N_A_218_119#_c_1698_n 8.90737e-19 $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_307 N_SCD_c_290_n N_A_218_119#_c_1698_n 0.010687f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_308 N_SCD_c_286_n N_VGND_c_1953_n 0.0128514f $X=0.655 $Y=1.125 $X2=0 $Y2=0
cc_309 N_SCD_c_287_n N_VGND_c_1953_n 0.00797474f $X=0.655 $Y=1.2 $X2=0 $Y2=0
cc_310 N_SCD_c_290_n N_VGND_c_1953_n 0.0226101f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_311 N_SCD_c_286_n N_VGND_c_1969_n 0.0035863f $X=0.655 $Y=1.125 $X2=0 $Y2=0
cc_312 N_SCD_c_286_n N_VGND_c_1982_n 0.00401353f $X=0.655 $Y=1.125 $X2=0 $Y2=0
cc_313 N_D_M1013_g N_A_346_93#_M1000_g 0.0637093f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_314 N_D_c_324_n N_A_346_93#_M1000_g 0.0233949f $X=1.355 $Y=1.905 $X2=0 $Y2=0
cc_315 N_D_M1017_g N_A_346_93#_M1031_g 0.0169158f $X=1.265 $Y=2.715 $X2=0 $Y2=0
cc_316 D N_A_346_93#_M1031_g 0.0130635f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_317 N_D_c_327_n N_A_346_93#_M1031_g 0.0217398f $X=1.355 $Y=2.07 $X2=0 $Y2=0
cc_318 D N_A_346_93#_c_382_n 0.0142173f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_319 D N_A_346_93#_c_383_n 0.00385004f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_320 D N_SCE_M1012_g 0.0126603f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_321 N_D_c_327_n N_SCE_M1012_g 0.0794227f $X=1.355 $Y=2.07 $X2=0 $Y2=0
cc_322 N_D_c_324_n N_SCE_M1012_g 0.00939796f $X=1.355 $Y=1.905 $X2=0 $Y2=0
cc_323 N_D_c_330_n N_SCE_M1012_g 0.00564086f $X=0.862 $Y=2.012 $X2=0 $Y2=0
cc_324 N_D_M1013_g N_SCE_M1009_g 0.0237811f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_325 N_D_c_323_n N_SCE_M1009_g 0.00822116f $X=1.43 $Y=1.515 $X2=0 $Y2=0
cc_326 N_D_M1013_g N_SCE_c_452_n 0.0103162f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_327 D N_SCE_c_457_n 0.00426321f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_328 N_D_c_324_n N_SCE_c_457_n 0.00822116f $X=1.355 $Y=1.905 $X2=0 $Y2=0
cc_329 N_D_c_330_n N_SCE_c_457_n 0.00105237f $X=0.862 $Y=2.012 $X2=0 $Y2=0
cc_330 N_D_M1017_g N_A_27_479#_c_1486_n 0.0126426f $X=1.265 $Y=2.715 $X2=0 $Y2=0
cc_331 D N_A_27_479#_c_1486_n 0.0220506f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_332 N_D_c_327_n N_A_27_479#_c_1486_n 0.00508121f $X=1.355 $Y=2.07 $X2=0 $Y2=0
cc_333 D N_A_27_479#_c_1486_n 0.112741f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_334 D N_A_27_479#_c_1487_n 0.0224562f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_335 N_D_M1017_g N_VPWR_c_1513_n 0.00187574f $X=1.265 $Y=2.715 $X2=0 $Y2=0
cc_336 N_D_M1017_g N_VPWR_c_1526_n 0.00526658f $X=1.265 $Y=2.715 $X2=0 $Y2=0
cc_337 N_D_M1017_g N_VPWR_c_1512_n 0.00592517f $X=1.265 $Y=2.715 $X2=0 $Y2=0
cc_338 N_D_M1013_g N_A_218_119#_c_1713_n 0.0123524f $X=1.445 $Y=0.805 $X2=0
+ $Y2=0
cc_339 N_D_M1013_g N_A_218_119#_c_1697_n 0.00896488f $X=1.445 $Y=0.805 $X2=0
+ $Y2=0
cc_340 N_D_c_323_n N_A_218_119#_c_1697_n 0.00327863f $X=1.43 $Y=1.515 $X2=0
+ $Y2=0
cc_341 D N_A_218_119#_c_1697_n 0.0410229f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_342 N_D_c_324_n N_A_218_119#_c_1697_n 0.00233826f $X=1.355 $Y=1.905 $X2=0
+ $Y2=0
cc_343 N_D_M1013_g N_A_218_119#_c_1698_n 0.00208912f $X=1.445 $Y=0.805 $X2=0
+ $Y2=0
cc_344 N_D_c_323_n N_A_218_119#_c_1698_n 0.00312041f $X=1.43 $Y=1.515 $X2=0
+ $Y2=0
cc_345 D N_A_218_119#_c_1698_n 0.0176069f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_346 N_D_c_327_n N_A_218_119#_c_1698_n 0.00101355f $X=1.355 $Y=2.07 $X2=0
+ $Y2=0
cc_347 N_D_c_324_n N_A_218_119#_c_1698_n 0.00152516f $X=1.355 $Y=1.905 $X2=0
+ $Y2=0
cc_348 D N_A_218_119#_c_1699_n 0.0236205f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_349 N_D_M1017_g N_A_218_119#_c_1712_n 8.74829e-19 $X=1.265 $Y=2.715 $X2=0
+ $Y2=0
cc_350 N_D_M1013_g N_VGND_c_1954_n 0.00177594f $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_351 N_D_M1013_g N_VGND_c_1982_n 9.39239e-19 $X=1.445 $Y=0.805 $X2=0 $Y2=0
cc_352 N_A_346_93#_M1000_g N_SCE_c_452_n 0.0103107f $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_353 N_A_346_93#_M1000_g N_SCE_M1001_g 0.0138939f $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_354 N_A_346_93#_c_382_n N_SCE_M1001_g 0.00181362f $X=2.695 $Y=1.83 $X2=0
+ $Y2=0
cc_355 N_A_346_93#_c_378_n N_SCE_M1001_g 0.00427933f $X=2.86 $Y=1.4 $X2=0 $Y2=0
cc_356 N_A_346_93#_c_377_n N_SCE_c_455_n 0.0117094f $X=2.765 $Y=0.805 $X2=0
+ $Y2=0
cc_357 N_A_346_93#_c_388_n N_SCE_c_465_n 0.00414277f $X=3.46 $Y=2.57 $X2=0 $Y2=0
cc_358 N_A_346_93#_c_378_n N_SCE_c_456_n 0.00342232f $X=2.86 $Y=1.4 $X2=0 $Y2=0
cc_359 N_A_346_93#_c_379_n N_SCE_c_456_n 0.0183657f $X=2.86 $Y=1.4 $X2=0 $Y2=0
cc_360 N_A_346_93#_c_386_n N_SCE_c_456_n 0.00926152f $X=3.365 $Y=2.015 $X2=0
+ $Y2=0
cc_361 N_A_346_93#_c_388_n N_SCE_c_456_n 0.00104853f $X=3.46 $Y=2.57 $X2=0 $Y2=0
cc_362 N_A_346_93#_c_386_n N_SCE_c_468_n 0.00849751f $X=3.365 $Y=2.015 $X2=0
+ $Y2=0
cc_363 N_A_346_93#_c_388_n N_SCE_c_468_n 0.0168602f $X=3.46 $Y=2.57 $X2=0 $Y2=0
cc_364 N_A_346_93#_c_377_n N_SCE_c_460_n 0.00658837f $X=2.765 $Y=0.805 $X2=0
+ $Y2=0
cc_365 N_A_346_93#_c_378_n N_SCE_c_460_n 0.00478834f $X=2.86 $Y=1.4 $X2=0 $Y2=0
cc_366 N_A_346_93#_c_377_n SCE 0.014215f $X=2.765 $Y=0.805 $X2=0 $Y2=0
cc_367 N_A_346_93#_c_378_n SCE 0.0290988f $X=2.86 $Y=1.4 $X2=0 $Y2=0
cc_368 N_A_346_93#_c_379_n SCE 0.00222157f $X=2.86 $Y=1.4 $X2=0 $Y2=0
cc_369 N_A_346_93#_c_386_n SCE 0.0163609f $X=3.365 $Y=2.015 $X2=0 $Y2=0
cc_370 N_A_346_93#_c_386_n N_CLK_M1042_g 3.98864e-19 $X=3.365 $Y=2.015 $X2=0
+ $Y2=0
cc_371 N_A_346_93#_c_388_n N_CLK_M1042_g 0.00511763f $X=3.46 $Y=2.57 $X2=0 $Y2=0
cc_372 N_A_346_93#_c_386_n N_A_773_409#_c_1071_n 0.0131015f $X=3.365 $Y=2.015
+ $X2=0 $Y2=0
cc_373 N_A_346_93#_c_388_n N_A_773_409#_c_1071_n 0.0143077f $X=3.46 $Y=2.57
+ $X2=0 $Y2=0
cc_374 N_A_346_93#_M1031_g N_A_27_479#_c_1486_n 0.0162507f $X=1.805 $Y=2.715
+ $X2=0 $Y2=0
cc_375 N_A_346_93#_c_382_n N_A_27_479#_c_1486_n 0.0010981f $X=2.695 $Y=1.83
+ $X2=0 $Y2=0
cc_376 N_A_346_93#_M1031_g N_VPWR_c_1526_n 0.00319878f $X=1.805 $Y=2.715 $X2=0
+ $Y2=0
cc_377 N_A_346_93#_M1031_g N_VPWR_c_1512_n 0.00571272f $X=1.805 $Y=2.715 $X2=0
+ $Y2=0
cc_378 N_A_346_93#_M1000_g N_A_218_119#_c_1713_n 0.0021239f $X=1.805 $Y=0.805
+ $X2=0 $Y2=0
cc_379 N_A_346_93#_M1000_g N_A_218_119#_c_1697_n 0.0246399f $X=1.805 $Y=0.805
+ $X2=0 $Y2=0
cc_380 N_A_346_93#_c_382_n N_A_218_119#_c_1697_n 0.0102497f $X=2.695 $Y=1.83
+ $X2=0 $Y2=0
cc_381 N_A_346_93#_c_377_n N_A_218_119#_c_1697_n 0.0153932f $X=2.765 $Y=0.805
+ $X2=0 $Y2=0
cc_382 N_A_346_93#_c_378_n N_A_218_119#_c_1697_n 0.0270462f $X=2.86 $Y=1.4 $X2=0
+ $Y2=0
cc_383 N_A_346_93#_c_379_n N_A_218_119#_c_1697_n 0.00773539f $X=2.86 $Y=1.4
+ $X2=0 $Y2=0
cc_384 N_A_346_93#_M1031_g N_A_218_119#_c_1702_n 0.0111005f $X=1.805 $Y=2.715
+ $X2=0 $Y2=0
cc_385 N_A_346_93#_M1031_g N_A_218_119#_c_1703_n 0.00251804f $X=1.805 $Y=2.715
+ $X2=0 $Y2=0
cc_386 N_A_346_93#_M1000_g N_A_218_119#_c_1699_n 0.00495338f $X=1.805 $Y=0.805
+ $X2=0 $Y2=0
cc_387 N_A_346_93#_M1031_g N_A_218_119#_c_1699_n 0.00500329f $X=1.805 $Y=2.715
+ $X2=0 $Y2=0
cc_388 N_A_346_93#_c_382_n N_A_218_119#_c_1699_n 0.0176128f $X=2.695 $Y=1.83
+ $X2=0 $Y2=0
cc_389 N_A_346_93#_c_378_n N_A_218_119#_c_1699_n 0.0282091f $X=2.86 $Y=1.4 $X2=0
+ $Y2=0
cc_390 N_A_346_93#_c_379_n N_A_218_119#_c_1699_n 0.0052118f $X=2.86 $Y=1.4 $X2=0
+ $Y2=0
cc_391 N_A_346_93#_c_387_n N_A_218_119#_c_1699_n 0.0143583f $X=3.025 $Y=2.015
+ $X2=0 $Y2=0
cc_392 N_A_346_93#_c_382_n N_A_218_119#_c_1705_n 0.00613425f $X=2.695 $Y=1.83
+ $X2=0 $Y2=0
cc_393 N_A_346_93#_c_386_n N_A_218_119#_c_1705_n 0.00987934f $X=3.365 $Y=2.015
+ $X2=0 $Y2=0
cc_394 N_A_346_93#_c_387_n N_A_218_119#_c_1705_n 0.0152872f $X=3.025 $Y=2.015
+ $X2=0 $Y2=0
cc_395 N_A_346_93#_c_388_n N_A_218_119#_c_1705_n 0.00792678f $X=3.46 $Y=2.57
+ $X2=0 $Y2=0
cc_396 N_A_346_93#_M1031_g N_A_218_119#_c_1706_n 3.41139e-19 $X=1.805 $Y=2.715
+ $X2=0 $Y2=0
cc_397 N_A_346_93#_c_382_n N_A_218_119#_c_1706_n 0.00339692f $X=2.695 $Y=1.83
+ $X2=0 $Y2=0
cc_398 N_A_346_93#_M1039_d N_A_218_119#_c_1707_n 0.00268105f $X=3.32 $Y=2.405
+ $X2=0 $Y2=0
cc_399 N_A_346_93#_c_388_n N_A_218_119#_c_1707_n 0.0189128f $X=3.46 $Y=2.57
+ $X2=0 $Y2=0
cc_400 N_A_346_93#_c_388_n N_A_218_119#_c_1752_n 0.00532669f $X=3.46 $Y=2.57
+ $X2=0 $Y2=0
cc_401 N_A_346_93#_c_388_n N_A_218_119#_c_1710_n 0.00899858f $X=3.46 $Y=2.57
+ $X2=0 $Y2=0
cc_402 N_A_346_93#_M1031_g N_A_218_119#_c_1712_n 3.15561e-19 $X=1.805 $Y=2.715
+ $X2=0 $Y2=0
cc_403 N_A_346_93#_M1000_g N_VGND_c_1954_n 0.0106103f $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_404 N_A_346_93#_c_377_n N_VGND_c_1970_n 0.0126564f $X=2.765 $Y=0.805 $X2=0
+ $Y2=0
cc_405 N_A_346_93#_M1000_g N_VGND_c_1982_n 7.88961e-19 $X=1.805 $Y=0.805 $X2=0
+ $Y2=0
cc_406 N_A_346_93#_c_377_n N_VGND_c_1982_n 0.0172104f $X=2.765 $Y=0.805 $X2=0
+ $Y2=0
cc_407 N_SCE_c_456_n N_CLK_M1042_g 0.00905238f $X=3.51 $Y=2.145 $X2=0 $Y2=0
cc_408 N_SCE_c_455_n N_CLK_M1037_g 0.00414758f $X=3.435 $Y=0.18 $X2=0 $Y2=0
cc_409 N_SCE_c_463_n N_CLK_M1037_g 0.00447524f $X=3.6 $Y=0.635 $X2=0 $Y2=0
cc_410 N_SCE_c_456_n N_CLK_c_555_n 0.00555499f $X=3.51 $Y=2.145 $X2=0 $Y2=0
cc_411 N_SCE_c_461_n N_CLK_c_555_n 0.00394057f $X=3.6 $Y=1.14 $X2=0 $Y2=0
cc_412 N_SCE_c_460_n N_CLK_c_557_n 0.00394057f $X=3.6 $Y=0.975 $X2=0 $Y2=0
cc_413 N_SCE_c_456_n N_A_773_409#_c_1071_n 0.00703704f $X=3.51 $Y=2.145 $X2=0
+ $Y2=0
cc_414 N_SCE_c_460_n N_A_773_409#_c_1071_n 0.00427351f $X=3.6 $Y=0.975 $X2=0
+ $Y2=0
cc_415 SCE N_A_773_409#_c_1071_n 0.0836267f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_416 N_SCE_c_459_n N_A_773_409#_c_1072_n 0.00173675f $X=3.6 $Y=0.47 $X2=0
+ $Y2=0
cc_417 SCE N_A_773_409#_c_1072_n 0.0215294f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_418 N_SCE_c_463_n N_A_773_409#_c_1072_n 0.00194184f $X=3.6 $Y=0.635 $X2=0
+ $Y2=0
cc_419 N_SCE_M1012_g N_A_27_479#_c_1486_n 0.011145f $X=0.905 $Y=2.715 $X2=0
+ $Y2=0
cc_420 N_SCE_M1012_g N_VPWR_c_1513_n 0.0117081f $X=0.905 $Y=2.715 $X2=0 $Y2=0
cc_421 N_SCE_c_465_n N_VPWR_c_1514_n 0.00400482f $X=3.245 $Y=2.295 $X2=0 $Y2=0
cc_422 N_SCE_M1012_g N_VPWR_c_1526_n 0.00437283f $X=0.905 $Y=2.715 $X2=0 $Y2=0
cc_423 N_SCE_c_465_n N_VPWR_c_1531_n 0.00325872f $X=3.245 $Y=2.295 $X2=0 $Y2=0
cc_424 N_SCE_M1012_g N_VPWR_c_1512_n 0.00420388f $X=0.905 $Y=2.715 $X2=0 $Y2=0
cc_425 N_SCE_c_465_n N_VPWR_c_1512_n 0.00666855f $X=3.245 $Y=2.295 $X2=0 $Y2=0
cc_426 N_SCE_M1009_g N_A_218_119#_c_1713_n 0.0124842f $X=1.015 $Y=0.805 $X2=0
+ $Y2=0
cc_427 N_SCE_c_452_n N_A_218_119#_c_1713_n 0.00339678f $X=2.16 $Y=0.18 $X2=0
+ $Y2=0
cc_428 N_SCE_M1001_g N_A_218_119#_c_1697_n 0.00459898f $X=2.235 $Y=0.805 $X2=0
+ $Y2=0
cc_429 N_SCE_M1009_g N_A_218_119#_c_1698_n 0.00860733f $X=1.015 $Y=0.805 $X2=0
+ $Y2=0
cc_430 N_SCE_c_457_n N_A_218_119#_c_1698_n 0.00109349f $X=1.015 $Y=1.59 $X2=0
+ $Y2=0
cc_431 N_SCE_c_465_n N_A_218_119#_c_1703_n 8.80021e-19 $X=3.245 $Y=2.295 $X2=0
+ $Y2=0
cc_432 N_SCE_c_468_n N_A_218_119#_c_1699_n 0.00581425f $X=3.51 $Y=2.22 $X2=0
+ $Y2=0
cc_433 N_SCE_c_465_n N_A_218_119#_c_1705_n 0.00627918f $X=3.245 $Y=2.295 $X2=0
+ $Y2=0
cc_434 N_SCE_c_465_n N_A_218_119#_c_1763_n 0.0147423f $X=3.245 $Y=2.295 $X2=0
+ $Y2=0
cc_435 N_SCE_c_465_n N_A_218_119#_c_1707_n 0.0124112f $X=3.245 $Y=2.295 $X2=0
+ $Y2=0
cc_436 N_SCE_c_468_n N_A_218_119#_c_1707_n 6.17753e-19 $X=3.51 $Y=2.22 $X2=0
+ $Y2=0
cc_437 N_SCE_c_465_n N_A_218_119#_c_1708_n 0.00351746f $X=3.245 $Y=2.295 $X2=0
+ $Y2=0
cc_438 N_SCE_c_465_n N_A_218_119#_c_1752_n 0.00359974f $X=3.245 $Y=2.295 $X2=0
+ $Y2=0
cc_439 N_SCE_M1009_g N_VGND_c_1953_n 0.00177594f $X=1.015 $Y=0.805 $X2=0 $Y2=0
cc_440 N_SCE_c_453_n N_VGND_c_1953_n 0.0101515f $X=1.09 $Y=0.18 $X2=0 $Y2=0
cc_441 N_SCE_c_452_n N_VGND_c_1954_n 0.0183681f $X=2.16 $Y=0.18 $X2=0 $Y2=0
cc_442 N_SCE_M1001_g N_VGND_c_1954_n 0.0263848f $X=2.235 $Y=0.805 $X2=0 $Y2=0
cc_443 N_SCE_c_458_n N_VGND_c_1954_n 0.00460513f $X=2.235 $Y=0.18 $X2=0 $Y2=0
cc_444 N_SCE_c_453_n N_VGND_c_1969_n 0.0296617f $X=1.09 $Y=0.18 $X2=0 $Y2=0
cc_445 N_SCE_c_458_n N_VGND_c_1970_n 0.0419271f $X=2.235 $Y=0.18 $X2=0 $Y2=0
cc_446 SCE N_VGND_c_1970_n 0.00949566f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_447 N_SCE_c_463_n N_VGND_c_1970_n 0.0024933f $X=3.6 $Y=0.635 $X2=0 $Y2=0
cc_448 N_SCE_c_452_n N_VGND_c_1982_n 0.0277107f $X=2.16 $Y=0.18 $X2=0 $Y2=0
cc_449 N_SCE_c_453_n N_VGND_c_1982_n 0.0108126f $X=1.09 $Y=0.18 $X2=0 $Y2=0
cc_450 N_SCE_c_455_n N_VGND_c_1982_n 0.0493858f $X=3.435 $Y=0.18 $X2=0 $Y2=0
cc_451 N_SCE_c_458_n N_VGND_c_1982_n 0.00749832f $X=2.235 $Y=0.18 $X2=0 $Y2=0
cc_452 SCE N_VGND_c_1982_n 0.00856505f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_453 N_SCE_c_463_n N_VGND_c_1982_n 0.00222868f $X=3.6 $Y=0.635 $X2=0 $Y2=0
cc_454 N_CLK_M1037_g N_A_773_409#_M1005_g 0.0135363f $X=4.32 $Y=0.495 $X2=0
+ $Y2=0
cc_455 CLK N_A_773_409#_M1005_g 0.00642798f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_456 N_CLK_c_557_n N_A_773_409#_M1005_g 0.00792343f $X=4.3 $Y=1.005 $X2=0
+ $Y2=0
cc_457 N_CLK_c_555_n N_A_773_409#_c_1065_n 0.00792343f $X=4.3 $Y=1.345 $X2=0
+ $Y2=0
cc_458 CLK N_A_773_409#_c_1065_n 0.00949179f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_459 N_CLK_M1042_g N_A_773_409#_c_1071_n 0.00500009f $X=4.3 $Y=2.775 $X2=0
+ $Y2=0
cc_460 N_CLK_M1037_g N_A_773_409#_c_1071_n 0.00354596f $X=4.32 $Y=0.495 $X2=0
+ $Y2=0
cc_461 CLK N_A_773_409#_c_1071_n 0.0752975f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_462 N_CLK_c_557_n N_A_773_409#_c_1071_n 0.0064365f $X=4.3 $Y=1.005 $X2=0
+ $Y2=0
cc_463 N_CLK_c_552_n N_A_773_409#_c_1088_n 0.00281214f $X=4.3 $Y=1.51 $X2=0
+ $Y2=0
cc_464 N_CLK_M1042_g N_A_773_409#_c_1088_n 0.0188705f $X=4.3 $Y=2.775 $X2=0
+ $Y2=0
cc_465 CLK N_A_773_409#_c_1088_n 0.0489848f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_466 N_CLK_M1042_g N_A_773_409#_c_1089_n 0.044374f $X=4.3 $Y=2.775 $X2=0 $Y2=0
cc_467 CLK N_A_773_409#_c_1089_n 0.00337774f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_468 N_CLK_c_557_n N_A_773_409#_c_1072_n 0.0027288f $X=4.3 $Y=1.005 $X2=0
+ $Y2=0
cc_469 N_CLK_M1042_g N_A_773_409#_c_1073_n 0.0105893f $X=4.3 $Y=2.775 $X2=0
+ $Y2=0
cc_470 N_CLK_c_555_n N_A_773_409#_c_1073_n 0.0118069f $X=4.3 $Y=1.345 $X2=0
+ $Y2=0
cc_471 CLK N_A_773_409#_c_1073_n 0.0112125f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_472 N_CLK_M1042_g N_VPWR_c_1515_n 0.00837679f $X=4.3 $Y=2.775 $X2=0 $Y2=0
cc_473 N_CLK_M1042_g N_VPWR_c_1531_n 0.00361815f $X=4.3 $Y=2.775 $X2=0 $Y2=0
cc_474 N_CLK_M1042_g N_VPWR_c_1512_n 0.00573574f $X=4.3 $Y=2.775 $X2=0 $Y2=0
cc_475 N_CLK_M1042_g N_A_218_119#_c_1709_n 0.0131124f $X=4.3 $Y=2.775 $X2=0
+ $Y2=0
cc_476 CLK N_A_218_119#_c_1700_n 0.0332304f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_477 N_CLK_M1037_g N_VGND_c_1955_n 0.00318388f $X=4.32 $Y=0.495 $X2=0 $Y2=0
cc_478 CLK N_VGND_c_1955_n 0.0185201f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_479 N_CLK_c_557_n N_VGND_c_1955_n 2.89144e-19 $X=4.3 $Y=1.005 $X2=0 $Y2=0
cc_480 N_CLK_M1037_g N_VGND_c_1970_n 0.0053602f $X=4.32 $Y=0.495 $X2=0 $Y2=0
cc_481 N_CLK_M1037_g N_VGND_c_1982_n 0.00621991f $X=4.32 $Y=0.495 $X2=0 $Y2=0
cc_482 CLK N_VGND_c_1982_n 0.0105942f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_483 N_A_961_491#_c_609_n N_A_1339_331#_M1025_g 0.00140192f $X=6.54 $Y=2.94
+ $X2=0 $Y2=0
cc_484 N_A_961_491#_c_610_n N_A_1339_331#_M1025_g 0.0101321f $X=6.63 $Y=2.805
+ $X2=0 $Y2=0
cc_485 N_A_961_491#_c_611_n N_A_1339_331#_M1025_g 0.0120325f $X=7.25 $Y=2.18
+ $X2=0 $Y2=0
cc_486 N_A_961_491#_c_612_n N_A_1339_331#_M1025_g 0.00244027f $X=6.72 $Y=2.18
+ $X2=0 $Y2=0
cc_487 N_A_961_491#_c_613_n N_A_1339_331#_M1025_g 0.00169781f $X=7.335 $Y=2.785
+ $X2=0 $Y2=0
cc_488 N_A_961_491#_c_611_n N_A_1339_331#_c_787_n 0.0531931f $X=7.25 $Y=2.18
+ $X2=0 $Y2=0
cc_489 N_A_961_491#_c_612_n N_A_1339_331#_c_787_n 0.0019325f $X=6.72 $Y=2.18
+ $X2=0 $Y2=0
cc_490 N_A_961_491#_c_628_p N_A_1339_331#_c_787_n 0.0115465f $X=8.12 $Y=1.88
+ $X2=0 $Y2=0
cc_491 N_A_961_491#_c_603_n N_A_1339_331#_c_787_n 9.51236e-19 $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_492 N_A_961_491#_M1033_g N_A_1339_331#_c_780_n 0.00233043f $X=5.98 $Y=2.525
+ $X2=0 $Y2=0
cc_493 N_A_961_491#_c_611_n N_A_1339_331#_c_780_n 0.00496257f $X=7.25 $Y=2.18
+ $X2=0 $Y2=0
cc_494 N_A_961_491#_c_603_n N_A_1339_331#_c_780_n 0.0159205f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_495 N_A_961_491#_M1008_g N_A_1339_331#_c_781_n 8.2089e-19 $X=6.5 $Y=0.615
+ $X2=0 $Y2=0
cc_496 N_A_961_491#_c_611_n N_A_1339_331#_c_789_n 0.0136934f $X=7.25 $Y=2.18
+ $X2=0 $Y2=0
cc_497 N_A_961_491#_c_613_n N_A_1339_331#_c_789_n 0.0137027f $X=7.335 $Y=2.785
+ $X2=0 $Y2=0
cc_498 N_A_961_491#_c_614_n N_A_1339_331#_c_789_n 0.0144329f $X=7.95 $Y=2.87
+ $X2=0 $Y2=0
cc_499 N_A_961_491#_c_616_n N_A_1339_331#_c_789_n 0.046466f $X=8.035 $Y=2.785
+ $X2=0 $Y2=0
cc_500 N_A_961_491#_c_628_p N_A_1339_331#_c_789_n 0.00318366f $X=8.12 $Y=1.88
+ $X2=0 $Y2=0
cc_501 N_A_961_491#_M1008_g N_A_1339_331#_c_784_n 0.0079817f $X=6.5 $Y=0.615
+ $X2=0 $Y2=0
cc_502 N_A_961_491#_c_603_n N_A_1339_331#_c_784_n 0.00584114f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_503 N_A_961_491#_M1008_g N_A_1339_331#_c_785_n 0.0595692f $X=6.5 $Y=0.615
+ $X2=0 $Y2=0
cc_504 N_A_961_491#_c_610_n N_A_1211_463#_M1029_g 2.04393e-19 $X=6.63 $Y=2.805
+ $X2=0 $Y2=0
cc_505 N_A_961_491#_c_611_n N_A_1211_463#_M1029_g 0.00526024f $X=7.25 $Y=2.18
+ $X2=0 $Y2=0
cc_506 N_A_961_491#_c_613_n N_A_1211_463#_M1029_g 0.0128602f $X=7.335 $Y=2.785
+ $X2=0 $Y2=0
cc_507 N_A_961_491#_c_614_n N_A_1211_463#_M1029_g 0.00793408f $X=7.95 $Y=2.87
+ $X2=0 $Y2=0
cc_508 N_A_961_491#_c_615_n N_A_1211_463#_M1029_g 0.00126155f $X=7.42 $Y=2.87
+ $X2=0 $Y2=0
cc_509 N_A_961_491#_c_616_n N_A_1211_463#_M1029_g 6.62752e-19 $X=8.035 $Y=2.785
+ $X2=0 $Y2=0
cc_510 N_A_961_491#_c_614_n N_A_1211_463#_M1010_g 2.00646e-19 $X=7.95 $Y=2.87
+ $X2=0 $Y2=0
cc_511 N_A_961_491#_c_616_n N_A_1211_463#_M1010_g 0.00319635f $X=8.035 $Y=2.785
+ $X2=0 $Y2=0
cc_512 N_A_961_491#_c_617_n N_A_1211_463#_M1010_g 2.43762e-19 $X=9.525 $Y=1.93
+ $X2=0 $Y2=0
cc_513 N_A_961_491#_c_618_n N_A_1211_463#_M1010_g 0.0166017f $X=9.36 $Y=1.905
+ $X2=0 $Y2=0
cc_514 N_A_961_491#_c_620_n N_A_1211_463#_M1010_g 0.00601788f $X=9.725 $Y=1.93
+ $X2=0 $Y2=0
cc_515 N_A_961_491#_c_617_n N_A_1211_463#_c_852_n 5.69189e-19 $X=9.525 $Y=1.93
+ $X2=0 $Y2=0
cc_516 N_A_961_491#_c_618_n N_A_1211_463#_c_852_n 0.00966534f $X=9.36 $Y=1.905
+ $X2=0 $Y2=0
cc_517 N_A_961_491#_c_620_n N_A_1211_463#_c_852_n 0.00499186f $X=9.725 $Y=1.93
+ $X2=0 $Y2=0
cc_518 N_A_961_491#_M1035_g N_A_1211_463#_c_853_n 0.0646104f $X=9.725 $Y=0.945
+ $X2=0 $Y2=0
cc_519 N_A_961_491#_M1008_g N_A_1211_463#_c_854_n 0.0102639f $X=6.5 $Y=0.615
+ $X2=0 $Y2=0
cc_520 N_A_961_491#_c_600_n N_A_1211_463#_c_854_n 0.0242571f $X=5.89 $Y=1.425
+ $X2=0 $Y2=0
cc_521 N_A_961_491#_c_603_n N_A_1211_463#_c_854_n 0.00725476f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_522 N_A_961_491#_c_608_n N_A_1211_463#_c_862_n 0.011547f $X=5.845 $Y=2.795
+ $X2=0 $Y2=0
cc_523 N_A_961_491#_c_609_n N_A_1211_463#_c_862_n 0.0185084f $X=6.54 $Y=2.94
+ $X2=0 $Y2=0
cc_524 N_A_961_491#_c_603_n N_A_1211_463#_c_862_n 0.00327113f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_525 N_A_961_491#_M1033_g N_A_1211_463#_c_863_n 0.00317912f $X=5.98 $Y=2.525
+ $X2=0 $Y2=0
cc_526 N_A_961_491#_c_664_p N_A_1211_463#_c_863_n 0.0294834f $X=5.845 $Y=1.46
+ $X2=0 $Y2=0
cc_527 N_A_961_491#_c_608_n N_A_1211_463#_c_863_n 0.0177472f $X=5.845 $Y=2.795
+ $X2=0 $Y2=0
cc_528 N_A_961_491#_c_610_n N_A_1211_463#_c_863_n 0.0151626f $X=6.63 $Y=2.805
+ $X2=0 $Y2=0
cc_529 N_A_961_491#_c_612_n N_A_1211_463#_c_863_n 0.0141085f $X=6.72 $Y=2.18
+ $X2=0 $Y2=0
cc_530 N_A_961_491#_c_603_n N_A_1211_463#_c_863_n 0.021599f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_531 N_A_961_491#_M1008_g N_A_1211_463#_c_855_n 0.00666485f $X=6.5 $Y=0.615
+ $X2=0 $Y2=0
cc_532 N_A_961_491#_c_602_n N_A_1211_463#_c_855_n 0.0242571f $X=5.89 $Y=1.295
+ $X2=0 $Y2=0
cc_533 N_A_961_491#_c_603_n N_A_1211_463#_c_855_n 0.00121914f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_534 N_A_961_491#_c_600_n N_A_1211_463#_c_895_n 0.0148734f $X=5.89 $Y=1.425
+ $X2=0 $Y2=0
cc_535 N_A_961_491#_c_603_n N_A_1211_463#_c_895_n 0.00597466f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_536 N_A_961_491#_c_618_n N_A_1211_463#_c_856_n 0.0238638f $X=9.36 $Y=1.905
+ $X2=0 $Y2=0
cc_537 N_A_961_491#_c_612_n N_A_1211_463#_c_857_n 0.00582769f $X=6.72 $Y=2.18
+ $X2=0 $Y2=0
cc_538 N_A_961_491#_c_628_p N_A_1211_463#_c_857_n 0.0102061f $X=8.12 $Y=1.88
+ $X2=0 $Y2=0
cc_539 N_A_961_491#_c_618_n N_A_1211_463#_c_857_n 0.0265901f $X=9.36 $Y=1.905
+ $X2=0 $Y2=0
cc_540 N_A_961_491#_c_603_n N_A_1211_463#_c_857_n 0.0155274f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_541 N_A_961_491#_M1035_g N_A_1211_463#_c_859_n 0.00333788f $X=9.725 $Y=0.945
+ $X2=0 $Y2=0
cc_542 N_A_961_491#_c_618_n N_A_1211_463#_c_859_n 0.0044365f $X=9.36 $Y=1.905
+ $X2=0 $Y2=0
cc_543 N_A_961_491#_c_613_n N_SET_B_M1018_g 5.30342e-19 $X=7.335 $Y=2.785 $X2=0
+ $Y2=0
cc_544 N_A_961_491#_c_614_n N_SET_B_M1018_g 0.00739051f $X=7.95 $Y=2.87 $X2=0
+ $Y2=0
cc_545 N_A_961_491#_c_616_n N_SET_B_M1018_g 0.0213579f $X=8.035 $Y=2.785 $X2=0
+ $Y2=0
cc_546 N_A_961_491#_c_628_p N_SET_B_M1018_g 0.00462269f $X=8.12 $Y=1.88 $X2=0
+ $Y2=0
cc_547 N_A_961_491#_c_628_p N_SET_B_c_974_n 0.00384434f $X=8.12 $Y=1.88 $X2=0
+ $Y2=0
cc_548 N_A_961_491#_c_618_n N_SET_B_c_974_n 0.00805473f $X=9.36 $Y=1.905 $X2=0
+ $Y2=0
cc_549 N_A_961_491#_c_628_p N_SET_B_c_975_n 9.72533e-19 $X=8.12 $Y=1.88 $X2=0
+ $Y2=0
cc_550 N_A_961_491#_M1035_g N_SET_B_c_972_n 0.0181831f $X=9.725 $Y=0.945 $X2=0
+ $Y2=0
cc_551 N_A_961_491#_c_607_n N_A_773_409#_M1023_g 0.00336422f $X=5.76 $Y=2.935
+ $X2=0 $Y2=0
cc_552 N_A_961_491#_c_601_n N_A_773_409#_M1005_g 0.00100807f $X=4.95 $Y=0.34
+ $X2=0 $Y2=0
cc_553 N_A_961_491#_c_599_n N_A_773_409#_c_1064_n 0.0115587f $X=5.85 $Y=0.34
+ $X2=0 $Y2=0
cc_554 N_A_961_491#_c_600_n N_A_773_409#_c_1064_n 5.87425e-19 $X=5.89 $Y=1.425
+ $X2=0 $Y2=0
cc_555 N_A_961_491#_c_602_n N_A_773_409#_c_1064_n 0.00892864f $X=5.89 $Y=1.295
+ $X2=0 $Y2=0
cc_556 N_A_961_491#_c_603_n N_A_773_409#_c_1064_n 0.0328218f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_557 N_A_961_491#_c_601_n N_A_773_409#_c_1065_n 0.0056879f $X=4.95 $Y=0.34
+ $X2=0 $Y2=0
cc_558 N_A_961_491#_M1033_g N_A_773_409#_c_1075_n 0.00944831f $X=5.98 $Y=2.525
+ $X2=0 $Y2=0
cc_559 N_A_961_491#_c_607_n N_A_773_409#_c_1076_n 0.0175803f $X=5.76 $Y=2.935
+ $X2=0 $Y2=0
cc_560 N_A_961_491#_c_608_n N_A_773_409#_c_1076_n 0.00357261f $X=5.845 $Y=2.795
+ $X2=0 $Y2=0
cc_561 N_A_961_491#_M1033_g N_A_773_409#_c_1077_n 0.00895246f $X=5.98 $Y=2.525
+ $X2=0 $Y2=0
cc_562 N_A_961_491#_c_607_n N_A_773_409#_c_1077_n 0.0089456f $X=5.76 $Y=2.935
+ $X2=0 $Y2=0
cc_563 N_A_961_491#_c_609_n N_A_773_409#_c_1077_n 0.00541734f $X=6.54 $Y=2.94
+ $X2=0 $Y2=0
cc_564 N_A_961_491#_c_702_p N_A_773_409#_c_1077_n 0.00378523f $X=5.845 $Y=2.935
+ $X2=0 $Y2=0
cc_565 N_A_961_491#_M1008_g N_A_773_409#_c_1066_n 0.0204558f $X=6.5 $Y=0.615
+ $X2=0 $Y2=0
cc_566 N_A_961_491#_c_599_n N_A_773_409#_c_1066_n 0.00694974f $X=5.85 $Y=0.34
+ $X2=0 $Y2=0
cc_567 N_A_961_491#_c_602_n N_A_773_409#_c_1066_n 0.0146948f $X=5.89 $Y=1.295
+ $X2=0 $Y2=0
cc_568 N_A_961_491#_M1033_g N_A_773_409#_M1022_g 0.0137097f $X=5.98 $Y=2.525
+ $X2=0 $Y2=0
cc_569 N_A_961_491#_c_608_n N_A_773_409#_M1022_g 6.29904e-19 $X=5.845 $Y=2.795
+ $X2=0 $Y2=0
cc_570 N_A_961_491#_c_609_n N_A_773_409#_M1022_g 0.0209799f $X=6.54 $Y=2.94
+ $X2=0 $Y2=0
cc_571 N_A_961_491#_c_610_n N_A_773_409#_M1022_g 0.00245818f $X=6.63 $Y=2.805
+ $X2=0 $Y2=0
cc_572 N_A_961_491#_c_612_n N_A_773_409#_M1022_g 5.69522e-19 $X=6.72 $Y=2.18
+ $X2=0 $Y2=0
cc_573 N_A_961_491#_c_603_n N_A_773_409#_M1022_g 0.00640448f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_574 N_A_961_491#_M1026_g N_A_773_409#_c_1080_n 0.00880325f $X=9.725 $Y=2.525
+ $X2=0 $Y2=0
cc_575 N_A_961_491#_c_609_n N_A_773_409#_c_1080_n 0.00465661f $X=6.54 $Y=2.94
+ $X2=0 $Y2=0
cc_576 N_A_961_491#_c_614_n N_A_773_409#_c_1080_n 0.0113689f $X=7.95 $Y=2.87
+ $X2=0 $Y2=0
cc_577 N_A_961_491#_c_615_n N_A_773_409#_c_1080_n 0.00359016f $X=7.42 $Y=2.87
+ $X2=0 $Y2=0
cc_578 N_A_961_491#_c_620_n N_A_773_409#_M1002_g 0.0187232f $X=9.725 $Y=1.93
+ $X2=0 $Y2=0
cc_579 N_A_961_491#_M1035_g N_A_773_409#_c_1068_n 0.0187232f $X=9.725 $Y=0.945
+ $X2=0 $Y2=0
cc_580 N_A_961_491#_c_603_n N_A_773_409#_c_1073_n 0.00682635f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_581 N_A_961_491#_c_617_n N_A_1960_125#_c_1293_n 0.00653633f $X=9.525 $Y=1.93
+ $X2=0 $Y2=0
cc_582 N_A_961_491#_c_620_n N_A_1960_125#_c_1293_n 0.00453357f $X=9.725 $Y=1.93
+ $X2=0 $Y2=0
cc_583 N_A_961_491#_M1035_g N_A_1960_125#_c_1287_n 0.0282089f $X=9.725 $Y=0.945
+ $X2=0 $Y2=0
cc_584 N_A_961_491#_c_617_n N_A_1960_125#_c_1287_n 0.0117173f $X=9.525 $Y=1.93
+ $X2=0 $Y2=0
cc_585 N_A_961_491#_c_613_n N_VPWR_M1025_d 0.00442123f $X=7.335 $Y=2.785 $X2=0
+ $Y2=0
cc_586 N_A_961_491#_c_616_n N_VPWR_M1018_d 0.00404792f $X=8.035 $Y=2.785 $X2=0
+ $Y2=0
cc_587 N_A_961_491#_c_618_n N_VPWR_M1018_d 0.00221108f $X=9.36 $Y=1.905 $X2=0
+ $Y2=0
cc_588 N_A_961_491#_c_607_n N_VPWR_c_1516_n 0.0627333f $X=5.76 $Y=2.935 $X2=0
+ $Y2=0
cc_589 N_A_961_491#_c_609_n N_VPWR_c_1516_n 0.0523249f $X=6.54 $Y=2.94 $X2=0
+ $Y2=0
cc_590 N_A_961_491#_c_702_p N_VPWR_c_1516_n 0.0115893f $X=5.845 $Y=2.935 $X2=0
+ $Y2=0
cc_591 N_A_961_491#_c_609_n N_VPWR_c_1517_n 0.0227047f $X=6.54 $Y=2.94 $X2=0
+ $Y2=0
cc_592 N_A_961_491#_c_610_n N_VPWR_c_1517_n 0.0152563f $X=6.63 $Y=2.805 $X2=0
+ $Y2=0
cc_593 N_A_961_491#_c_611_n N_VPWR_c_1517_n 0.015052f $X=7.25 $Y=2.18 $X2=0
+ $Y2=0
cc_594 N_A_961_491#_c_613_n N_VPWR_c_1517_n 0.0257323f $X=7.335 $Y=2.785 $X2=0
+ $Y2=0
cc_595 N_A_961_491#_c_615_n N_VPWR_c_1517_n 0.0144673f $X=7.42 $Y=2.87 $X2=0
+ $Y2=0
cc_596 N_A_961_491#_c_614_n N_VPWR_c_1518_n 0.0144403f $X=7.95 $Y=2.87 $X2=0
+ $Y2=0
cc_597 N_A_961_491#_c_616_n N_VPWR_c_1518_n 0.048239f $X=8.035 $Y=2.785 $X2=0
+ $Y2=0
cc_598 N_A_961_491#_c_618_n N_VPWR_c_1518_n 0.0220024f $X=9.36 $Y=1.905 $X2=0
+ $Y2=0
cc_599 N_A_961_491#_c_614_n N_VPWR_c_1532_n 0.0262848f $X=7.95 $Y=2.87 $X2=0
+ $Y2=0
cc_600 N_A_961_491#_c_615_n N_VPWR_c_1532_n 0.0068857f $X=7.42 $Y=2.87 $X2=0
+ $Y2=0
cc_601 N_A_961_491#_M1023_d N_VPWR_c_1512_n 0.00212318f $X=4.805 $Y=2.455 $X2=0
+ $Y2=0
cc_602 N_A_961_491#_c_607_n N_VPWR_c_1512_n 0.0344959f $X=5.76 $Y=2.935 $X2=0
+ $Y2=0
cc_603 N_A_961_491#_c_609_n N_VPWR_c_1512_n 0.0267577f $X=6.54 $Y=2.94 $X2=0
+ $Y2=0
cc_604 N_A_961_491#_c_614_n N_VPWR_c_1512_n 0.0217828f $X=7.95 $Y=2.87 $X2=0
+ $Y2=0
cc_605 N_A_961_491#_c_615_n N_VPWR_c_1512_n 0.00550129f $X=7.42 $Y=2.87 $X2=0
+ $Y2=0
cc_606 N_A_961_491#_c_702_p N_VPWR_c_1512_n 0.00583135f $X=5.845 $Y=2.935 $X2=0
+ $Y2=0
cc_607 N_A_961_491#_c_599_n N_A_218_119#_M1041_s 0.00614391f $X=5.85 $Y=0.34
+ $X2=0 $Y2=0
cc_608 N_A_961_491#_c_602_n N_A_218_119#_M1041_s 0.008944f $X=5.89 $Y=1.295
+ $X2=0 $Y2=0
cc_609 N_A_961_491#_c_608_n N_A_218_119#_M1033_s 0.00452284f $X=5.845 $Y=2.795
+ $X2=0 $Y2=0
cc_610 N_A_961_491#_M1023_d N_A_218_119#_c_1709_n 0.00465233f $X=4.805 $Y=2.455
+ $X2=0 $Y2=0
cc_611 N_A_961_491#_c_607_n N_A_218_119#_c_1709_n 0.0358781f $X=5.76 $Y=2.935
+ $X2=0 $Y2=0
cc_612 N_A_961_491#_M1033_g N_A_218_119#_c_1700_n 0.00238461f $X=5.98 $Y=2.525
+ $X2=0 $Y2=0
cc_613 N_A_961_491#_c_607_n N_A_218_119#_c_1700_n 0.0204747f $X=5.76 $Y=2.935
+ $X2=0 $Y2=0
cc_614 N_A_961_491#_c_600_n N_A_218_119#_c_1700_n 0.0884388f $X=5.89 $Y=1.425
+ $X2=0 $Y2=0
cc_615 N_A_961_491#_c_608_n N_A_218_119#_c_1700_n 0.0138309f $X=5.845 $Y=2.795
+ $X2=0 $Y2=0
cc_616 N_A_961_491#_c_602_n N_A_218_119#_c_1700_n 0.0269683f $X=5.89 $Y=1.295
+ $X2=0 $Y2=0
cc_617 N_A_961_491#_c_603_n N_A_218_119#_c_1700_n 0.0097916f $X=5.98 $Y=1.63
+ $X2=0 $Y2=0
cc_618 N_A_961_491#_c_599_n N_A_218_119#_c_1701_n 0.025217f $X=5.85 $Y=0.34
+ $X2=0 $Y2=0
cc_619 N_A_961_491#_c_601_n N_A_218_119#_c_1701_n 0.00373916f $X=4.95 $Y=0.34
+ $X2=0 $Y2=0
cc_620 N_A_961_491#_c_602_n N_A_218_119#_c_1701_n 0.0160861f $X=5.89 $Y=1.295
+ $X2=0 $Y2=0
cc_621 N_A_961_491#_c_618_n N_A_1751_379#_M1010_d 0.0033259f $X=9.36 $Y=1.905
+ $X2=-0.19 $Y2=-0.245
cc_622 N_A_961_491#_M1026_g N_A_1751_379#_c_1843_n 0.00374726f $X=9.725 $Y=2.525
+ $X2=0 $Y2=0
cc_623 N_A_961_491#_c_618_n N_A_1751_379#_c_1843_n 0.00882135f $X=9.36 $Y=1.905
+ $X2=0 $Y2=0
cc_624 N_A_961_491#_M1026_g N_A_1751_379#_c_1840_n 2.29152e-19 $X=9.725 $Y=2.525
+ $X2=0 $Y2=0
cc_625 N_A_961_491#_M1026_g N_A_1751_379#_c_1841_n 0.0171911f $X=9.725 $Y=2.525
+ $X2=0 $Y2=0
cc_626 N_A_961_491#_c_617_n N_A_1751_379#_c_1841_n 0.0165057f $X=9.525 $Y=1.93
+ $X2=0 $Y2=0
cc_627 N_A_961_491#_c_618_n N_A_1751_379#_c_1841_n 0.0171207f $X=9.36 $Y=1.905
+ $X2=0 $Y2=0
cc_628 N_A_961_491#_c_620_n N_A_1751_379#_c_1841_n 0.00663534f $X=9.725 $Y=1.93
+ $X2=0 $Y2=0
cc_629 N_A_961_491#_M1026_g N_A_1858_463#_c_1870_n 0.011795f $X=9.725 $Y=2.525
+ $X2=0 $Y2=0
cc_630 N_A_961_491#_M1026_g N_A_1858_463#_c_1871_n 0.00203065f $X=9.725 $Y=2.525
+ $X2=0 $Y2=0
cc_631 N_A_961_491#_c_601_n N_VGND_c_1955_n 0.00230656f $X=4.95 $Y=0.34 $X2=0
+ $Y2=0
cc_632 N_A_961_491#_M1008_g N_VGND_c_1956_n 0.00197091f $X=6.5 $Y=0.615 $X2=0
+ $Y2=0
cc_633 N_A_961_491#_M1035_g N_VGND_c_1959_n 9.91921e-19 $X=9.725 $Y=0.945 $X2=0
+ $Y2=0
cc_634 N_A_961_491#_c_618_n N_VGND_c_1959_n 0.010898f $X=9.36 $Y=1.905 $X2=0
+ $Y2=0
cc_635 N_A_961_491#_M1008_g N_VGND_c_1971_n 0.00530021f $X=6.5 $Y=0.615 $X2=0
+ $Y2=0
cc_636 N_A_961_491#_c_599_n N_VGND_c_1971_n 0.0624039f $X=5.85 $Y=0.34 $X2=0
+ $Y2=0
cc_637 N_A_961_491#_c_601_n N_VGND_c_1971_n 0.0164155f $X=4.95 $Y=0.34 $X2=0
+ $Y2=0
cc_638 N_A_961_491#_M1035_g N_VGND_c_1972_n 5.34712e-19 $X=9.725 $Y=0.945 $X2=0
+ $Y2=0
cc_639 N_A_961_491#_M1008_g N_VGND_c_1982_n 0.00534666f $X=6.5 $Y=0.615 $X2=0
+ $Y2=0
cc_640 N_A_961_491#_c_599_n N_VGND_c_1982_n 0.0359315f $X=5.85 $Y=0.34 $X2=0
+ $Y2=0
cc_641 N_A_961_491#_c_601_n N_VGND_c_1982_n 0.00913237f $X=4.95 $Y=0.34 $X2=0
+ $Y2=0
cc_642 N_A_1339_331#_M1025_g N_A_1211_463#_M1029_g 0.012444f $X=6.77 $Y=2.525
+ $X2=0 $Y2=0
cc_643 N_A_1339_331#_c_787_n N_A_1211_463#_M1029_g 0.016151f $X=7.59 $Y=1.82
+ $X2=0 $Y2=0
cc_644 N_A_1339_331#_c_789_n N_A_1211_463#_M1029_g 0.00596385f $X=7.685 $Y=2.45
+ $X2=0 $Y2=0
cc_645 N_A_1339_331#_c_784_n N_A_1211_463#_M1029_g 0.0128236f $X=6.86 $Y=1.655
+ $X2=0 $Y2=0
cc_646 N_A_1339_331#_c_787_n N_A_1211_463#_c_850_n 7.50437e-19 $X=7.59 $Y=1.82
+ $X2=0 $Y2=0
cc_647 N_A_1339_331#_c_783_n N_A_1211_463#_M1027_g 0.00309709f $X=7.7 $Y=0.9
+ $X2=0 $Y2=0
cc_648 N_A_1339_331#_c_781_n N_A_1211_463#_c_854_n 0.0095158f $X=7.595 $Y=1.067
+ $X2=0 $Y2=0
cc_649 N_A_1339_331#_c_784_n N_A_1211_463#_c_854_n 2.51581e-19 $X=6.86 $Y=1.655
+ $X2=0 $Y2=0
cc_650 N_A_1339_331#_M1025_g N_A_1211_463#_c_863_n 6.10694e-19 $X=6.77 $Y=2.525
+ $X2=0 $Y2=0
cc_651 N_A_1339_331#_c_787_n N_A_1211_463#_c_863_n 0.00944586f $X=7.59 $Y=1.82
+ $X2=0 $Y2=0
cc_652 N_A_1339_331#_c_780_n N_A_1211_463#_c_863_n 0.00348457f $X=6.86 $Y=1.82
+ $X2=0 $Y2=0
cc_653 N_A_1339_331#_c_784_n N_A_1211_463#_c_863_n 5.53506e-19 $X=6.86 $Y=1.655
+ $X2=0 $Y2=0
cc_654 N_A_1339_331#_c_785_n N_A_1211_463#_c_855_n 0.00109603f $X=6.95 $Y=0.935
+ $X2=0 $Y2=0
cc_655 N_A_1339_331#_c_787_n N_A_1211_463#_c_857_n 0.0815007f $X=7.59 $Y=1.82
+ $X2=0 $Y2=0
cc_656 N_A_1339_331#_c_780_n N_A_1211_463#_c_857_n 0.00338934f $X=6.86 $Y=1.82
+ $X2=0 $Y2=0
cc_657 N_A_1339_331#_c_781_n N_A_1211_463#_c_857_n 0.0601404f $X=7.595 $Y=1.067
+ $X2=0 $Y2=0
cc_658 N_A_1339_331#_c_782_n N_A_1211_463#_c_857_n 0.00313427f $X=6.95 $Y=1.1
+ $X2=0 $Y2=0
cc_659 N_A_1339_331#_c_783_n N_A_1211_463#_c_857_n 0.0147152f $X=7.7 $Y=0.9
+ $X2=0 $Y2=0
cc_660 N_A_1339_331#_c_784_n N_A_1211_463#_c_857_n 0.0118384f $X=6.86 $Y=1.655
+ $X2=0 $Y2=0
cc_661 N_A_1339_331#_c_787_n N_A_1211_463#_c_858_n 0.00447463f $X=7.59 $Y=1.82
+ $X2=0 $Y2=0
cc_662 N_A_1339_331#_c_781_n N_A_1211_463#_c_858_n 0.00731873f $X=7.595 $Y=1.067
+ $X2=0 $Y2=0
cc_663 N_A_1339_331#_c_783_n N_A_1211_463#_c_858_n 0.00424918f $X=7.7 $Y=0.9
+ $X2=0 $Y2=0
cc_664 N_A_1339_331#_c_784_n N_A_1211_463#_c_858_n 0.0154804f $X=6.86 $Y=1.655
+ $X2=0 $Y2=0
cc_665 N_A_1339_331#_c_789_n N_SET_B_M1018_g 0.00357862f $X=7.685 $Y=2.45 $X2=0
+ $Y2=0
cc_666 N_A_1339_331#_c_787_n N_SET_B_c_975_n 0.00366687f $X=7.59 $Y=1.82 $X2=0
+ $Y2=0
cc_667 N_A_1339_331#_M1025_g N_A_773_409#_M1022_g 0.039927f $X=6.77 $Y=2.525
+ $X2=0 $Y2=0
cc_668 N_A_1339_331#_M1025_g N_A_773_409#_c_1080_n 0.0103024f $X=6.77 $Y=2.525
+ $X2=0 $Y2=0
cc_669 N_A_1339_331#_M1025_g N_VPWR_c_1517_n 0.00135426f $X=6.77 $Y=2.525 $X2=0
+ $Y2=0
cc_670 N_A_1339_331#_M1025_g N_VPWR_c_1512_n 7.82699e-19 $X=6.77 $Y=2.525 $X2=0
+ $Y2=0
cc_671 N_A_1339_331#_c_781_n N_VGND_c_1956_n 0.0243489f $X=7.595 $Y=1.067 $X2=0
+ $Y2=0
cc_672 N_A_1339_331#_c_782_n N_VGND_c_1956_n 0.00445138f $X=6.95 $Y=1.1 $X2=0
+ $Y2=0
cc_673 N_A_1339_331#_c_783_n N_VGND_c_1956_n 0.00209319f $X=7.7 $Y=0.9 $X2=0
+ $Y2=0
cc_674 N_A_1339_331#_c_785_n N_VGND_c_1956_n 0.0121736f $X=6.95 $Y=0.935 $X2=0
+ $Y2=0
cc_675 N_A_1339_331#_c_783_n N_VGND_c_1958_n 0.0192076f $X=7.7 $Y=0.9 $X2=0
+ $Y2=0
cc_676 N_A_1339_331#_c_783_n N_VGND_c_1967_n 0.0028554f $X=7.7 $Y=0.9 $X2=0
+ $Y2=0
cc_677 N_A_1339_331#_c_785_n N_VGND_c_1971_n 0.0045897f $X=6.95 $Y=0.935 $X2=0
+ $Y2=0
cc_678 N_A_1339_331#_c_783_n N_VGND_c_1982_n 0.00518644f $X=7.7 $Y=0.9 $X2=0
+ $Y2=0
cc_679 N_A_1339_331#_c_785_n N_VGND_c_1982_n 0.0044912f $X=6.95 $Y=0.935 $X2=0
+ $Y2=0
cc_680 N_A_1211_463#_M1010_g N_SET_B_M1018_g 0.00969536f $X=8.68 $Y=2.315 $X2=0
+ $Y2=0
cc_681 N_A_1211_463#_M1010_g N_SET_B_c_974_n 0.0120041f $X=8.68 $Y=2.315 $X2=0
+ $Y2=0
cc_682 N_A_1211_463#_M1029_g N_SET_B_c_975_n 0.0285944f $X=7.47 $Y=2.525 $X2=0
+ $Y2=0
cc_683 N_A_1211_463#_c_850_n N_SET_B_c_975_n 0.00695688f $X=7.84 $Y=1.355 $X2=0
+ $Y2=0
cc_684 N_A_1211_463#_c_857_n N_SET_B_c_975_n 0.00690956f $X=8.605 $Y=1.49 $X2=0
+ $Y2=0
cc_685 N_A_1211_463#_M1027_g N_SET_B_c_966_n 0.0295317f $X=7.915 $Y=0.835 $X2=0
+ $Y2=0
cc_686 N_A_1211_463#_c_853_n N_SET_B_c_966_n 2.33609e-19 $X=9.365 $Y=1.375 $X2=0
+ $Y2=0
cc_687 N_A_1211_463#_M1029_g N_SET_B_M1032_g 0.00125061f $X=7.47 $Y=2.525 $X2=0
+ $Y2=0
cc_688 N_A_1211_463#_c_850_n N_SET_B_M1032_g 0.0295317f $X=7.84 $Y=1.355 $X2=0
+ $Y2=0
cc_689 N_A_1211_463#_c_856_n N_SET_B_M1032_g 5.06407e-19 $X=8.77 $Y=1.54 $X2=0
+ $Y2=0
cc_690 N_A_1211_463#_c_857_n N_SET_B_M1032_g 0.0122059f $X=8.605 $Y=1.49 $X2=0
+ $Y2=0
cc_691 N_A_1211_463#_c_858_n N_SET_B_M1032_g 0.00396309f $X=7.49 $Y=1.355 $X2=0
+ $Y2=0
cc_692 N_A_1211_463#_c_859_n N_SET_B_M1032_g 0.0120041f $X=8.77 $Y=1.45 $X2=0
+ $Y2=0
cc_693 N_A_1211_463#_c_853_n N_SET_B_c_972_n 0.0172321f $X=9.365 $Y=1.375 $X2=0
+ $Y2=0
cc_694 N_A_1211_463#_c_854_n N_A_773_409#_c_1064_n 0.00107106f $X=6.28 $Y=1.355
+ $X2=0 $Y2=0
cc_695 N_A_1211_463#_c_855_n N_A_773_409#_c_1066_n 0.00107106f $X=6.285 $Y=0.7
+ $X2=0 $Y2=0
cc_696 N_A_1211_463#_c_862_n N_A_773_409#_M1022_g 0.00407671f $X=6.195 $Y=2.47
+ $X2=0 $Y2=0
cc_697 N_A_1211_463#_c_863_n N_A_773_409#_M1022_g 0.00247018f $X=6.235 $Y=2.305
+ $X2=0 $Y2=0
cc_698 N_A_1211_463#_c_857_n N_A_773_409#_M1022_g 0.00173918f $X=8.605 $Y=1.49
+ $X2=0 $Y2=0
cc_699 N_A_1211_463#_M1029_g N_A_773_409#_c_1080_n 0.00885705f $X=7.47 $Y=2.525
+ $X2=0 $Y2=0
cc_700 N_A_1211_463#_M1010_g N_A_773_409#_c_1080_n 0.0103107f $X=8.68 $Y=2.315
+ $X2=0 $Y2=0
cc_701 N_A_1211_463#_M1029_g N_VPWR_c_1517_n 0.00118842f $X=7.47 $Y=2.525 $X2=0
+ $Y2=0
cc_702 N_A_1211_463#_M1010_g N_VPWR_c_1518_n 0.0183005f $X=8.68 $Y=2.315 $X2=0
+ $Y2=0
cc_703 N_A_1211_463#_M1010_g N_VPWR_c_1512_n 7.88961e-19 $X=8.68 $Y=2.315 $X2=0
+ $Y2=0
cc_704 N_A_1211_463#_M1010_g N_A_1858_463#_c_1871_n 0.00365079f $X=8.68 $Y=2.315
+ $X2=0 $Y2=0
cc_705 N_A_1211_463#_M1027_g N_VGND_c_1956_n 0.00547746f $X=7.915 $Y=0.835 $X2=0
+ $Y2=0
cc_706 N_A_1211_463#_c_855_n N_VGND_c_1956_n 0.00805003f $X=6.285 $Y=0.7 $X2=0
+ $Y2=0
cc_707 N_A_1211_463#_M1027_g N_VGND_c_1957_n 0.0131998f $X=7.915 $Y=0.835 $X2=0
+ $Y2=0
cc_708 N_A_1211_463#_M1027_g N_VGND_c_1958_n 0.00732386f $X=7.915 $Y=0.835 $X2=0
+ $Y2=0
cc_709 N_A_1211_463#_c_857_n N_VGND_c_1958_n 0.0142171f $X=8.605 $Y=1.49 $X2=0
+ $Y2=0
cc_710 N_A_1211_463#_c_852_n N_VGND_c_1959_n 0.00808422f $X=9.29 $Y=1.45 $X2=0
+ $Y2=0
cc_711 N_A_1211_463#_c_853_n N_VGND_c_1959_n 0.00698752f $X=9.365 $Y=1.375 $X2=0
+ $Y2=0
cc_712 N_A_1211_463#_c_857_n N_VGND_c_1959_n 0.0636517f $X=8.605 $Y=1.49 $X2=0
+ $Y2=0
cc_713 N_A_1211_463#_c_859_n N_VGND_c_1959_n 0.00231231f $X=8.77 $Y=1.45 $X2=0
+ $Y2=0
cc_714 N_A_1211_463#_M1027_g N_VGND_c_1967_n 0.00345209f $X=7.915 $Y=0.835 $X2=0
+ $Y2=0
cc_715 N_A_1211_463#_c_855_n N_VGND_c_1971_n 0.00542506f $X=6.285 $Y=0.7 $X2=0
+ $Y2=0
cc_716 N_A_1211_463#_c_853_n N_VGND_c_1972_n 5.34712e-19 $X=9.365 $Y=1.375 $X2=0
+ $Y2=0
cc_717 N_A_1211_463#_M1027_g N_VGND_c_1982_n 0.00394323f $X=7.915 $Y=0.835 $X2=0
+ $Y2=0
cc_718 N_A_1211_463#_c_855_n N_VGND_c_1982_n 0.00830702f $X=6.285 $Y=0.7 $X2=0
+ $Y2=0
cc_719 N_SET_B_M1018_g N_A_773_409#_c_1080_n 0.0088568f $X=7.94 $Y=2.525 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_978_n N_A_773_409#_M1002_g 2.31323e-19 $X=10.855 $Y=1.675 $X2=0
+ $Y2=0
cc_721 N_SET_B_c_969_n N_A_773_409#_M1020_g 0.0224783f $X=10.77 $Y=1.585 $X2=0
+ $Y2=0
cc_722 N_SET_B_c_972_n N_A_773_409#_M1020_g 0.0109354f $X=10.685 $Y=0.46 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_978_n N_A_773_409#_c_1084_n 0.00461719f $X=10.855 $Y=1.675
+ $X2=0 $Y2=0
cc_724 N_SET_B_c_969_n N_A_773_409#_c_1070_n 0.0031045f $X=10.77 $Y=1.585 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_978_n N_A_773_409#_c_1070_n 0.00447487f $X=10.855 $Y=1.675
+ $X2=0 $Y2=0
cc_726 N_SET_B_M1024_g N_A_2205_231#_M1019_g 0.0186422f $X=11.64 $Y=0.835 $X2=0
+ $Y2=0
cc_727 N_SET_B_M1003_g N_A_2205_231#_M1019_g 0.041381f $X=11.66 $Y=2.795 $X2=0
+ $Y2=0
cc_728 N_SET_B_c_969_n N_A_2205_231#_M1019_g 0.00180151f $X=10.77 $Y=1.585 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_970_n N_A_2205_231#_M1019_g 0.0110041f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_730 N_SET_B_M1024_g N_A_2205_231#_c_1228_n 0.0180619f $X=11.64 $Y=0.835 $X2=0
+ $Y2=0
cc_731 N_SET_B_c_969_n N_A_2205_231#_c_1228_n 0.01902f $X=10.77 $Y=1.585 $X2=0
+ $Y2=0
cc_732 N_SET_B_c_970_n N_A_2205_231#_c_1228_n 0.0638402f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_971_n N_A_2205_231#_c_1228_n 0.00456089f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_734 N_SET_B_M1024_g N_A_2205_231#_c_1229_n 0.0218326f $X=11.64 $Y=0.835 $X2=0
+ $Y2=0
cc_735 N_SET_B_c_969_n N_A_2205_231#_c_1229_n 0.00257422f $X=10.77 $Y=1.585
+ $X2=0 $Y2=0
cc_736 N_SET_B_c_970_n N_A_2205_231#_c_1229_n 0.00466614f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_737 N_SET_B_M1024_g N_A_2205_231#_c_1233_n 0.0268481f $X=11.64 $Y=0.835 $X2=0
+ $Y2=0
cc_738 N_SET_B_c_969_n N_A_2205_231#_c_1233_n 0.00318042f $X=10.77 $Y=1.585
+ $X2=0 $Y2=0
cc_739 N_SET_B_c_972_n N_A_2205_231#_c_1233_n 0.00340416f $X=10.685 $Y=0.46
+ $X2=0 $Y2=0
cc_740 N_SET_B_c_972_n N_A_1960_125#_M1035_d 0.0126957f $X=10.685 $Y=0.46
+ $X2=-0.19 $Y2=-0.245
cc_741 N_SET_B_M1024_g N_A_1960_125#_M1043_g 0.0180524f $X=11.64 $Y=0.835 $X2=0
+ $Y2=0
cc_742 N_SET_B_c_971_n N_A_1960_125#_M1043_g 0.0150183f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_743 N_SET_B_M1003_g N_A_1960_125#_c_1283_n 0.0110494f $X=11.66 $Y=2.795 $X2=0
+ $Y2=0
cc_744 N_SET_B_c_970_n N_A_1960_125#_c_1283_n 6.08674e-19 $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_745 N_SET_B_c_971_n N_A_1960_125#_c_1283_n 0.00593204f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_746 N_SET_B_c_969_n N_A_1960_125#_c_1287_n 0.0586921f $X=10.77 $Y=1.585 $X2=0
+ $Y2=0
cc_747 N_SET_B_c_978_n N_A_1960_125#_c_1287_n 0.0153729f $X=10.855 $Y=1.675
+ $X2=0 $Y2=0
cc_748 N_SET_B_c_972_n N_A_1960_125#_c_1287_n 0.0541695f $X=10.685 $Y=0.46 $X2=0
+ $Y2=0
cc_749 N_SET_B_M1003_g N_A_1960_125#_c_1295_n 0.0165091f $X=11.66 $Y=2.795 $X2=0
+ $Y2=0
cc_750 N_SET_B_c_978_n N_A_1960_125#_c_1295_n 0.0133834f $X=10.855 $Y=1.675
+ $X2=0 $Y2=0
cc_751 N_SET_B_c_970_n N_A_1960_125#_c_1295_n 0.0672205f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_752 N_SET_B_c_971_n N_A_1960_125#_c_1295_n 0.00142553f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_753 N_SET_B_M1003_g N_A_1960_125#_c_1296_n 0.00635818f $X=11.66 $Y=2.795
+ $X2=0 $Y2=0
cc_754 N_SET_B_c_970_n N_A_1960_125#_c_1296_n 0.0221632f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_755 N_SET_B_c_971_n N_A_1960_125#_c_1296_n 0.00510576f $X=11.73 $Y=1.67 $X2=0
+ $Y2=0
cc_756 N_SET_B_M1003_g N_A_1960_125#_c_1297_n 0.0142092f $X=11.66 $Y=2.795 $X2=0
+ $Y2=0
cc_757 N_SET_B_M1018_g N_VPWR_c_1518_n 0.00246998f $X=7.94 $Y=2.525 $X2=0 $Y2=0
cc_758 N_SET_B_c_974_n N_VPWR_c_1518_n 2.70818e-19 $X=8.2 $Y=1.745 $X2=0 $Y2=0
cc_759 N_SET_B_M1003_g N_VPWR_c_1519_n 0.00316325f $X=11.66 $Y=2.795 $X2=0 $Y2=0
cc_760 N_SET_B_M1003_g N_VPWR_c_1520_n 0.00499542f $X=11.66 $Y=2.795 $X2=0 $Y2=0
cc_761 N_SET_B_M1003_g N_VPWR_c_1521_n 0.00436568f $X=11.66 $Y=2.795 $X2=0 $Y2=0
cc_762 N_SET_B_M1003_g N_VPWR_c_1512_n 0.0102719f $X=11.66 $Y=2.795 $X2=0 $Y2=0
cc_763 N_SET_B_c_972_n N_VGND_M1032_d 0.00965879f $X=10.685 $Y=0.46 $X2=0 $Y2=0
cc_764 N_SET_B_c_966_n N_VGND_c_1957_n 0.0112014f $X=8.275 $Y=0.515 $X2=0 $Y2=0
cc_765 N_SET_B_c_972_n N_VGND_c_1957_n 0.0330034f $X=10.685 $Y=0.46 $X2=0 $Y2=0
cc_766 N_SET_B_c_966_n N_VGND_c_1959_n 0.00141836f $X=8.275 $Y=0.515 $X2=0 $Y2=0
cc_767 N_SET_B_M1032_g N_VGND_c_1959_n 0.0166381f $X=8.275 $Y=0.835 $X2=0 $Y2=0
cc_768 N_SET_B_c_972_n N_VGND_c_1959_n 0.0711012f $X=10.685 $Y=0.46 $X2=0 $Y2=0
cc_769 N_SET_B_M1024_g N_VGND_c_1960_n 0.00391968f $X=11.64 $Y=0.835 $X2=0 $Y2=0
cc_770 N_SET_B_c_966_n N_VGND_c_1972_n 0.00976578f $X=8.275 $Y=0.515 $X2=0 $Y2=0
cc_771 N_SET_B_M1024_g N_VGND_c_1972_n 0.00415323f $X=11.64 $Y=0.835 $X2=0 $Y2=0
cc_772 N_SET_B_c_972_n N_VGND_c_1972_n 0.174288f $X=10.685 $Y=0.46 $X2=0 $Y2=0
cc_773 N_SET_B_c_966_n N_VGND_c_1982_n 0.0135145f $X=8.275 $Y=0.515 $X2=0 $Y2=0
cc_774 N_SET_B_M1024_g N_VGND_c_1982_n 0.00469432f $X=11.64 $Y=0.835 $X2=0 $Y2=0
cc_775 N_SET_B_c_972_n N_VGND_c_1982_n 0.0963884f $X=10.685 $Y=0.46 $X2=0 $Y2=0
cc_776 N_SET_B_c_972_n A_1888_125# 0.00407361f $X=10.685 $Y=0.46 $X2=-0.19
+ $Y2=-0.245
cc_777 N_A_773_409#_c_1070_n N_A_2205_231#_M1019_g 0.0557873f $X=10.74 $Y=1.59
+ $X2=0 $Y2=0
cc_778 N_A_773_409#_M1020_g N_A_2205_231#_c_1228_n 2.755e-19 $X=10.74 $Y=0.835
+ $X2=0 $Y2=0
cc_779 N_A_773_409#_M1020_g N_A_2205_231#_c_1229_n 0.0210755f $X=10.74 $Y=0.835
+ $X2=0 $Y2=0
cc_780 N_A_773_409#_M1020_g N_A_2205_231#_c_1233_n 0.0277652f $X=10.74 $Y=0.835
+ $X2=0 $Y2=0
cc_781 N_A_773_409#_M1002_g N_A_1960_125#_c_1293_n 0.00748127f $X=10.25 $Y=2.315
+ $X2=0 $Y2=0
cc_782 N_A_773_409#_M1002_g N_A_1960_125#_c_1287_n 0.00888687f $X=10.25 $Y=2.315
+ $X2=0 $Y2=0
cc_783 N_A_773_409#_c_1067_n N_A_1960_125#_c_1287_n 0.01325f $X=10.665 $Y=1.59
+ $X2=0 $Y2=0
cc_784 N_A_773_409#_c_1068_n N_A_1960_125#_c_1287_n 0.00912423f $X=10.325
+ $Y=1.59 $X2=0 $Y2=0
cc_785 N_A_773_409#_M1020_g N_A_1960_125#_c_1287_n 0.0132222f $X=10.74 $Y=0.835
+ $X2=0 $Y2=0
cc_786 N_A_773_409#_c_1084_n N_A_1960_125#_c_1287_n 0.00420414f $X=10.74
+ $Y=3.075 $X2=0 $Y2=0
cc_787 N_A_773_409#_c_1067_n N_A_1960_125#_c_1295_n 0.00198902f $X=10.665
+ $Y=1.59 $X2=0 $Y2=0
cc_788 N_A_773_409#_c_1084_n N_A_1960_125#_c_1295_n 0.0145293f $X=10.74 $Y=3.075
+ $X2=0 $Y2=0
cc_789 N_A_773_409#_M1023_g N_VPWR_c_1515_n 0.00289494f $X=4.73 $Y=2.775 $X2=0
+ $Y2=0
cc_790 N_A_773_409#_M1023_g N_VPWR_c_1516_n 0.00422236f $X=4.73 $Y=2.775 $X2=0
+ $Y2=0
cc_791 N_A_773_409#_c_1078_n N_VPWR_c_1516_n 0.039746f $X=5.295 $Y=3.15 $X2=0
+ $Y2=0
cc_792 N_A_773_409#_M1022_g N_VPWR_c_1517_n 8.99742e-19 $X=6.41 $Y=2.525 $X2=0
+ $Y2=0
cc_793 N_A_773_409#_c_1080_n N_VPWR_c_1517_n 0.018118f $X=10.665 $Y=3.15 $X2=0
+ $Y2=0
cc_794 N_A_773_409#_c_1080_n N_VPWR_c_1518_n 0.025796f $X=10.665 $Y=3.15 $X2=0
+ $Y2=0
cc_795 N_A_773_409#_c_1084_n N_VPWR_c_1519_n 0.00171883f $X=10.74 $Y=3.075 $X2=0
+ $Y2=0
cc_796 N_A_773_409#_c_1080_n N_VPWR_c_1528_n 0.0533117f $X=10.665 $Y=3.15 $X2=0
+ $Y2=0
cc_797 N_A_773_409#_c_1080_n N_VPWR_c_1532_n 0.0312107f $X=10.665 $Y=3.15 $X2=0
+ $Y2=0
cc_798 N_A_773_409#_M1042_s N_VPWR_c_1512_n 0.00316316f $X=3.865 $Y=2.045 $X2=0
+ $Y2=0
cc_799 N_A_773_409#_M1023_g N_VPWR_c_1512_n 0.00594684f $X=4.73 $Y=2.775 $X2=0
+ $Y2=0
cc_800 N_A_773_409#_c_1077_n N_VPWR_c_1512_n 0.0244405f $X=6.335 $Y=3.15 $X2=0
+ $Y2=0
cc_801 N_A_773_409#_c_1078_n N_VPWR_c_1512_n 0.00472465f $X=5.295 $Y=3.15 $X2=0
+ $Y2=0
cc_802 N_A_773_409#_c_1080_n N_VPWR_c_1512_n 0.109306f $X=10.665 $Y=3.15 $X2=0
+ $Y2=0
cc_803 N_A_773_409#_c_1085_n N_VPWR_c_1512_n 0.00370846f $X=6.41 $Y=3.15 $X2=0
+ $Y2=0
cc_804 N_A_773_409#_M1042_s N_A_218_119#_c_1707_n 0.00754581f $X=3.865 $Y=2.045
+ $X2=0 $Y2=0
cc_805 N_A_773_409#_c_1071_n N_A_218_119#_c_1707_n 0.00402227f $X=3.95 $Y=1.945
+ $X2=0 $Y2=0
cc_806 N_A_773_409#_M1042_s N_A_218_119#_c_1752_n 0.00650858f $X=3.865 $Y=2.045
+ $X2=0 $Y2=0
cc_807 N_A_773_409#_M1023_g N_A_218_119#_c_1709_n 0.0121747f $X=4.73 $Y=2.775
+ $X2=0 $Y2=0
cc_808 N_A_773_409#_c_1075_n N_A_218_119#_c_1709_n 0.00235412f $X=5.145 $Y=2.2
+ $X2=0 $Y2=0
cc_809 N_A_773_409#_c_1076_n N_A_218_119#_c_1709_n 0.0154769f $X=5.22 $Y=3.075
+ $X2=0 $Y2=0
cc_810 N_A_773_409#_c_1088_n N_A_218_119#_c_1709_n 0.0530915f $X=4.82 $Y=2.11
+ $X2=0 $Y2=0
cc_811 N_A_773_409#_c_1089_n N_A_218_119#_c_1709_n 6.08979e-19 $X=4.82 $Y=2.11
+ $X2=0 $Y2=0
cc_812 N_A_773_409#_M1042_s N_A_218_119#_c_1710_n 0.00553125f $X=3.865 $Y=2.045
+ $X2=0 $Y2=0
cc_813 N_A_773_409#_c_1071_n N_A_218_119#_c_1710_n 0.00716387f $X=3.95 $Y=1.945
+ $X2=0 $Y2=0
cc_814 N_A_773_409#_c_1088_n N_A_218_119#_c_1710_n 0.0118144f $X=4.82 $Y=2.11
+ $X2=0 $Y2=0
cc_815 N_A_773_409#_c_1064_n N_A_218_119#_c_1700_n 0.0212561f $X=5.995 $Y=1.01
+ $X2=0 $Y2=0
cc_816 N_A_773_409#_c_1075_n N_A_218_119#_c_1700_n 0.00779828f $X=5.145 $Y=2.2
+ $X2=0 $Y2=0
cc_817 N_A_773_409#_c_1066_n N_A_218_119#_c_1700_n 6.51386e-19 $X=6.07 $Y=0.935
+ $X2=0 $Y2=0
cc_818 N_A_773_409#_c_1088_n N_A_218_119#_c_1700_n 0.0160161f $X=4.82 $Y=2.11
+ $X2=0 $Y2=0
cc_819 N_A_773_409#_c_1089_n N_A_218_119#_c_1700_n 5.23956e-19 $X=4.82 $Y=2.11
+ $X2=0 $Y2=0
cc_820 N_A_773_409#_c_1073_n N_A_218_119#_c_1700_n 0.0105883f $X=4.82 $Y=1.945
+ $X2=0 $Y2=0
cc_821 N_A_773_409#_M1005_g N_A_218_119#_c_1701_n 0.00577127f $X=4.75 $Y=0.495
+ $X2=0 $Y2=0
cc_822 N_A_773_409#_c_1064_n N_A_218_119#_c_1701_n 0.00326982f $X=5.995 $Y=1.01
+ $X2=0 $Y2=0
cc_823 N_A_773_409#_c_1066_n N_A_218_119#_c_1701_n 0.00111095f $X=6.07 $Y=0.935
+ $X2=0 $Y2=0
cc_824 N_A_773_409#_c_1080_n N_A_1751_379#_c_1843_n 0.00342666f $X=10.665
+ $Y=3.15 $X2=0 $Y2=0
cc_825 N_A_773_409#_M1002_g N_A_1751_379#_c_1840_n 0.00202342f $X=10.25 $Y=2.315
+ $X2=0 $Y2=0
cc_826 N_A_773_409#_c_1067_n N_A_1751_379#_c_1840_n 3.77055e-19 $X=10.665
+ $Y=1.59 $X2=0 $Y2=0
cc_827 N_A_773_409#_c_1084_n N_A_1751_379#_c_1840_n 0.00735469f $X=10.74
+ $Y=3.075 $X2=0 $Y2=0
cc_828 N_A_773_409#_c_1080_n N_A_1751_379#_c_1841_n 0.00586836f $X=10.665
+ $Y=3.15 $X2=0 $Y2=0
cc_829 N_A_773_409#_M1002_g N_A_1751_379#_c_1841_n 0.00825059f $X=10.25 $Y=2.315
+ $X2=0 $Y2=0
cc_830 N_A_773_409#_M1002_g N_A_1858_463#_c_1870_n 0.0104736f $X=10.25 $Y=2.315
+ $X2=0 $Y2=0
cc_831 N_A_773_409#_c_1084_n N_A_1858_463#_c_1870_n 0.019496f $X=10.74 $Y=3.075
+ $X2=0 $Y2=0
cc_832 N_A_773_409#_c_1080_n N_A_1858_463#_c_1871_n 0.0262438f $X=10.665 $Y=3.15
+ $X2=0 $Y2=0
cc_833 N_A_773_409#_M1005_g N_VGND_c_1955_n 0.00262871f $X=4.75 $Y=0.495 $X2=0
+ $Y2=0
cc_834 N_A_773_409#_c_1072_n N_VGND_c_1970_n 0.0158654f $X=4.105 $Y=0.495 $X2=0
+ $Y2=0
cc_835 N_A_773_409#_M1005_g N_VGND_c_1971_n 0.0053602f $X=4.75 $Y=0.495 $X2=0
+ $Y2=0
cc_836 N_A_773_409#_c_1066_n N_VGND_c_1971_n 0.0047553f $X=6.07 $Y=0.935 $X2=0
+ $Y2=0
cc_837 N_A_773_409#_M1020_g N_VGND_c_1972_n 5.5016e-19 $X=10.74 $Y=0.835 $X2=0
+ $Y2=0
cc_838 N_A_773_409#_M1005_g N_VGND_c_1982_n 0.00801313f $X=4.75 $Y=0.495 $X2=0
+ $Y2=0
cc_839 N_A_773_409#_c_1066_n N_VGND_c_1982_n 0.00445555f $X=6.07 $Y=0.935 $X2=0
+ $Y2=0
cc_840 N_A_773_409#_c_1072_n N_VGND_c_1982_n 0.0136931f $X=4.105 $Y=0.495 $X2=0
+ $Y2=0
cc_841 N_A_2205_231#_c_1228_n N_A_1960_125#_M1043_g 0.0214621f $X=12.265
+ $Y=1.295 $X2=0 $Y2=0
cc_842 N_A_2205_231#_c_1231_n N_A_1960_125#_M1043_g 0.0058203f $X=12.395 $Y=0.84
+ $X2=0 $Y2=0
cc_843 N_A_2205_231#_c_1232_n N_A_1960_125#_M1043_g 0.00437521f $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_844 N_A_2205_231#_c_1230_n N_A_1960_125#_c_1283_n 0.0135756f $X=12.412
+ $Y=1.175 $X2=0 $Y2=0
cc_845 N_A_2205_231#_c_1232_n N_A_1960_125#_c_1283_n 0.0219311f $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_846 N_A_2205_231#_c_1232_n N_A_1960_125#_c_1284_n 0.0202013f $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_847 N_A_2205_231#_c_1232_n N_A_1960_125#_M1007_g 5.8321e-19 $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_848 N_A_2205_231#_M1019_g N_A_1960_125#_c_1287_n 7.66396e-19 $X=11.23
+ $Y=2.795 $X2=0 $Y2=0
cc_849 N_A_2205_231#_M1019_g N_A_1960_125#_c_1295_n 0.0161942f $X=11.23 $Y=2.795
+ $X2=0 $Y2=0
cc_850 N_A_2205_231#_c_1228_n N_A_1960_125#_c_1296_n 0.0204949f $X=12.265
+ $Y=1.295 $X2=0 $Y2=0
cc_851 N_A_2205_231#_c_1230_n N_A_1960_125#_c_1296_n 0.0178133f $X=12.412
+ $Y=1.175 $X2=0 $Y2=0
cc_852 N_A_2205_231#_c_1232_n N_A_1960_125#_c_1296_n 0.0427257f $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_853 N_A_2205_231#_c_1232_n N_A_1960_125#_c_1297_n 0.00586341f $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_854 N_A_2205_231#_c_1230_n N_A_2638_53#_c_1384_n 0.0177724f $X=12.412
+ $Y=1.175 $X2=0 $Y2=0
cc_855 N_A_2205_231#_c_1231_n N_A_2638_53#_c_1384_n 0.016806f $X=12.395 $Y=0.84
+ $X2=0 $Y2=0
cc_856 N_A_2205_231#_c_1232_n N_A_2638_53#_c_1384_n 7.27691e-19 $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_857 N_A_2205_231#_c_1232_n N_A_2638_53#_c_1392_n 0.0973414f $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_858 N_A_2205_231#_c_1232_n N_A_2638_53#_c_1386_n 0.0147472f $X=12.825
+ $Y=2.625 $X2=0 $Y2=0
cc_859 N_A_2205_231#_M1019_g N_VPWR_c_1519_n 0.0028524f $X=11.23 $Y=2.795 $X2=0
+ $Y2=0
cc_860 N_A_2205_231#_M1019_g N_VPWR_c_1528_n 0.00499542f $X=11.23 $Y=2.795 $X2=0
+ $Y2=0
cc_861 N_A_2205_231#_c_1232_n N_VPWR_c_1533_n 0.00655356f $X=12.825 $Y=2.625
+ $X2=0 $Y2=0
cc_862 N_A_2205_231#_M1019_g N_VPWR_c_1512_n 0.00983483f $X=11.23 $Y=2.795 $X2=0
+ $Y2=0
cc_863 N_A_2205_231#_c_1232_n N_VPWR_c_1512_n 0.00952812f $X=12.825 $Y=2.625
+ $X2=0 $Y2=0
cc_864 N_A_2205_231#_c_1228_n N_VGND_c_1960_n 0.0254551f $X=12.265 $Y=1.295
+ $X2=0 $Y2=0
cc_865 N_A_2205_231#_c_1233_n N_VGND_c_1972_n 0.00415323f $X=11.19 $Y=1.155
+ $X2=0 $Y2=0
cc_866 N_A_2205_231#_c_1231_n N_VGND_c_1973_n 0.00481978f $X=12.395 $Y=0.84
+ $X2=0 $Y2=0
cc_867 N_A_2205_231#_c_1231_n N_VGND_c_1982_n 0.00863262f $X=12.395 $Y=0.84
+ $X2=0 $Y2=0
cc_868 N_A_2205_231#_c_1233_n N_VGND_c_1982_n 0.00469432f $X=11.19 $Y=1.155
+ $X2=0 $Y2=0
cc_869 N_A_1960_125#_M1007_g N_A_2638_53#_M1004_g 0.0246651f $X=13.53 $Y=0.685
+ $X2=0 $Y2=0
cc_870 N_A_1960_125#_c_1286_n N_A_2638_53#_M1006_g 0.0210225f $X=13.545 $Y=1.65
+ $X2=0 $Y2=0
cc_871 N_A_1960_125#_M1007_g N_A_2638_53#_c_1384_n 0.0142962f $X=13.53 $Y=0.685
+ $X2=0 $Y2=0
cc_872 N_A_1960_125#_M1015_g N_A_2638_53#_c_1392_n 0.0041278f $X=12.61 $Y=2.625
+ $X2=0 $Y2=0
cc_873 N_A_1960_125#_c_1284_n N_A_2638_53#_c_1392_n 0.0110427f $X=13.455 $Y=1.65
+ $X2=0 $Y2=0
cc_874 N_A_1960_125#_c_1291_n N_A_2638_53#_c_1392_n 0.00678313f $X=13.56
+ $Y=1.725 $X2=0 $Y2=0
cc_875 N_A_1960_125#_c_1286_n N_A_2638_53#_c_1392_n 0.00235753f $X=13.545
+ $Y=1.65 $X2=0 $Y2=0
cc_876 N_A_1960_125#_M1007_g N_A_2638_53#_c_1385_n 0.00809938f $X=13.53 $Y=0.685
+ $X2=0 $Y2=0
cc_877 N_A_1960_125#_c_1286_n N_A_2638_53#_c_1385_n 0.0077815f $X=13.545 $Y=1.65
+ $X2=0 $Y2=0
cc_878 N_A_1960_125#_c_1284_n N_A_2638_53#_c_1386_n 0.00578208f $X=13.455
+ $Y=1.65 $X2=0 $Y2=0
cc_879 N_A_1960_125#_M1007_g N_A_2638_53#_c_1386_n 0.00463588f $X=13.53 $Y=0.685
+ $X2=0 $Y2=0
cc_880 N_A_1960_125#_M1007_g N_A_2638_53#_c_1387_n 0.0130981f $X=13.53 $Y=0.685
+ $X2=0 $Y2=0
cc_881 N_A_1960_125#_c_1286_n N_A_2638_53#_c_1387_n 0.00757265f $X=13.545
+ $Y=1.65 $X2=0 $Y2=0
cc_882 N_A_1960_125#_c_1295_n N_VPWR_c_1519_n 0.0070708f $X=11.77 $Y=2.03 $X2=0
+ $Y2=0
cc_883 N_A_1960_125#_c_1297_n N_VPWR_c_1520_n 0.0112322f $X=11.875 $Y=2.795
+ $X2=0 $Y2=0
cc_884 N_A_1960_125#_c_1283_n N_VPWR_c_1521_n 0.00344961f $X=12.61 $Y=2.255
+ $X2=0 $Y2=0
cc_885 N_A_1960_125#_M1015_g N_VPWR_c_1521_n 0.00427376f $X=12.61 $Y=2.625 $X2=0
+ $Y2=0
cc_886 N_A_1960_125#_c_1296_n N_VPWR_c_1521_n 0.0177319f $X=11.915 $Y=2.255
+ $X2=0 $Y2=0
cc_887 N_A_1960_125#_c_1297_n N_VPWR_c_1521_n 0.0408809f $X=11.875 $Y=2.795
+ $X2=0 $Y2=0
cc_888 N_A_1960_125#_c_1291_n N_VPWR_c_1522_n 0.00417057f $X=13.56 $Y=1.725
+ $X2=0 $Y2=0
cc_889 N_A_1960_125#_M1015_g N_VPWR_c_1533_n 0.00490845f $X=12.61 $Y=2.625 $X2=0
+ $Y2=0
cc_890 N_A_1960_125#_c_1291_n N_VPWR_c_1533_n 0.00585385f $X=13.56 $Y=1.725
+ $X2=0 $Y2=0
cc_891 N_A_1960_125#_M1015_g N_VPWR_c_1512_n 0.00506877f $X=12.61 $Y=2.625 $X2=0
+ $Y2=0
cc_892 N_A_1960_125#_c_1291_n N_VPWR_c_1512_n 0.0118611f $X=13.56 $Y=1.725 $X2=0
+ $Y2=0
cc_893 N_A_1960_125#_c_1297_n N_VPWR_c_1512_n 0.0105077f $X=11.875 $Y=2.795
+ $X2=0 $Y2=0
cc_894 N_A_1960_125#_c_1293_n N_A_1751_379#_M1002_d 0.00146434f $X=10.192
+ $Y=1.935 $X2=0 $Y2=0
cc_895 N_A_1960_125#_c_1287_n N_A_1751_379#_M1002_d 5.24516e-19 $X=10.43 $Y=1
+ $X2=0 $Y2=0
cc_896 N_A_1960_125#_c_1295_n N_A_1751_379#_M1002_d 0.00210204f $X=11.77 $Y=2.03
+ $X2=0 $Y2=0
cc_897 N_A_1960_125#_c_1295_n N_A_1751_379#_c_1840_n 0.00869108f $X=11.77
+ $Y=2.03 $X2=0 $Y2=0
cc_898 N_A_1960_125#_M1026_d N_A_1751_379#_c_1841_n 0.00515281f $X=9.8 $Y=2.315
+ $X2=0 $Y2=0
cc_899 N_A_1960_125#_c_1293_n N_A_1751_379#_c_1841_n 0.0427257f $X=10.192
+ $Y=1.935 $X2=0 $Y2=0
cc_900 N_A_1960_125#_M1026_d N_A_1858_463#_c_1870_n 0.00320957f $X=9.8 $Y=2.315
+ $X2=0 $Y2=0
cc_901 N_A_1960_125#_c_1295_n N_A_1858_463#_c_1870_n 0.0149747f $X=11.77 $Y=2.03
+ $X2=0 $Y2=0
cc_902 N_A_1960_125#_c_1287_n N_VGND_c_1959_n 0.0118833f $X=10.43 $Y=1 $X2=0
+ $Y2=0
cc_903 N_A_1960_125#_M1043_g N_VGND_c_1960_n 0.00391968f $X=12.18 $Y=0.835 $X2=0
+ $Y2=0
cc_904 N_A_1960_125#_M1007_g N_VGND_c_1961_n 0.0170097f $X=13.53 $Y=0.685 $X2=0
+ $Y2=0
cc_905 N_A_1960_125#_M1043_g N_VGND_c_1973_n 0.00415323f $X=12.18 $Y=0.835 $X2=0
+ $Y2=0
cc_906 N_A_1960_125#_M1007_g N_VGND_c_1973_n 0.00461019f $X=13.53 $Y=0.685 $X2=0
+ $Y2=0
cc_907 N_A_1960_125#_M1043_g N_VGND_c_1982_n 0.00469432f $X=12.18 $Y=0.835 $X2=0
+ $Y2=0
cc_908 N_A_1960_125#_M1007_g N_VGND_c_1982_n 0.00930161f $X=13.53 $Y=0.685 $X2=0
+ $Y2=0
cc_909 N_A_2638_53#_c_1392_n N_VPWR_c_1521_n 0.00857149f $X=13.345 $Y=1.98 $X2=0
+ $Y2=0
cc_910 N_A_2638_53#_M1006_g N_VPWR_c_1522_n 0.00268145f $X=13.99 $Y=2.465 $X2=0
+ $Y2=0
cc_911 N_A_2638_53#_c_1392_n N_VPWR_c_1522_n 0.00154474f $X=13.345 $Y=1.98 $X2=0
+ $Y2=0
cc_912 N_A_2638_53#_c_1385_n N_VPWR_c_1522_n 0.0172614f $X=14.69 $Y=1.51 $X2=0
+ $Y2=0
cc_913 N_A_2638_53#_c_1387_n N_VPWR_c_1522_n 0.00140804f $X=15.28 $Y=1.51 $X2=0
+ $Y2=0
cc_914 N_A_2638_53#_M1006_g N_VPWR_c_1523_n 7.40567e-19 $X=13.99 $Y=2.465 $X2=0
+ $Y2=0
cc_915 N_A_2638_53#_M1021_g N_VPWR_c_1523_n 0.0142699f $X=14.42 $Y=2.465 $X2=0
+ $Y2=0
cc_916 N_A_2638_53#_M1034_g N_VPWR_c_1523_n 0.0141781f $X=14.85 $Y=2.465 $X2=0
+ $Y2=0
cc_917 N_A_2638_53#_M1044_g N_VPWR_c_1523_n 7.24342e-19 $X=15.28 $Y=2.465 $X2=0
+ $Y2=0
cc_918 N_A_2638_53#_M1034_g N_VPWR_c_1525_n 7.24342e-19 $X=14.85 $Y=2.465 $X2=0
+ $Y2=0
cc_919 N_A_2638_53#_M1044_g N_VPWR_c_1525_n 0.0152818f $X=15.28 $Y=2.465 $X2=0
+ $Y2=0
cc_920 N_A_2638_53#_c_1392_n N_VPWR_c_1533_n 0.0206641f $X=13.345 $Y=1.98 $X2=0
+ $Y2=0
cc_921 N_A_2638_53#_M1006_g N_VPWR_c_1534_n 0.00585385f $X=13.99 $Y=2.465 $X2=0
+ $Y2=0
cc_922 N_A_2638_53#_M1021_g N_VPWR_c_1534_n 0.00486043f $X=14.42 $Y=2.465 $X2=0
+ $Y2=0
cc_923 N_A_2638_53#_M1034_g N_VPWR_c_1535_n 0.00486043f $X=14.85 $Y=2.465 $X2=0
+ $Y2=0
cc_924 N_A_2638_53#_M1044_g N_VPWR_c_1535_n 0.00486043f $X=15.28 $Y=2.465 $X2=0
+ $Y2=0
cc_925 N_A_2638_53#_M1040_s N_VPWR_c_1512_n 0.00232552f $X=13.22 $Y=1.835 $X2=0
+ $Y2=0
cc_926 N_A_2638_53#_M1006_g N_VPWR_c_1512_n 0.0105614f $X=13.99 $Y=2.465 $X2=0
+ $Y2=0
cc_927 N_A_2638_53#_M1021_g N_VPWR_c_1512_n 0.00824727f $X=14.42 $Y=2.465 $X2=0
+ $Y2=0
cc_928 N_A_2638_53#_M1034_g N_VPWR_c_1512_n 0.00824727f $X=14.85 $Y=2.465 $X2=0
+ $Y2=0
cc_929 N_A_2638_53#_M1044_g N_VPWR_c_1512_n 0.00824727f $X=15.28 $Y=2.465 $X2=0
+ $Y2=0
cc_930 N_A_2638_53#_c_1392_n N_VPWR_c_1512_n 0.0123631f $X=13.345 $Y=1.98 $X2=0
+ $Y2=0
cc_931 N_A_2638_53#_M1004_g N_Q_c_1889_n 7.99655e-19 $X=13.96 $Y=0.685 $X2=0
+ $Y2=0
cc_932 N_A_2638_53#_M1030_g N_Q_c_1889_n 7.99655e-19 $X=14.39 $Y=0.685 $X2=0
+ $Y2=0
cc_933 N_A_2638_53#_M1030_g N_Q_c_1890_n 0.0139613f $X=14.39 $Y=0.685 $X2=0
+ $Y2=0
cc_934 N_A_2638_53#_M1036_g N_Q_c_1890_n 0.0147289f $X=14.82 $Y=0.685 $X2=0
+ $Y2=0
cc_935 N_A_2638_53#_c_1385_n N_Q_c_1890_n 0.0410179f $X=14.69 $Y=1.51 $X2=0
+ $Y2=0
cc_936 N_A_2638_53#_c_1387_n N_Q_c_1890_n 0.00259709f $X=15.28 $Y=1.51 $X2=0
+ $Y2=0
cc_937 N_A_2638_53#_M1004_g N_Q_c_1891_n 0.00230792f $X=13.96 $Y=0.685 $X2=0
+ $Y2=0
cc_938 N_A_2638_53#_c_1384_n N_Q_c_1891_n 0.00405716f $X=13.315 $Y=0.42 $X2=0
+ $Y2=0
cc_939 N_A_2638_53#_c_1385_n N_Q_c_1891_n 0.0153308f $X=14.69 $Y=1.51 $X2=0
+ $Y2=0
cc_940 N_A_2638_53#_c_1387_n N_Q_c_1891_n 0.00269667f $X=15.28 $Y=1.51 $X2=0
+ $Y2=0
cc_941 N_A_2638_53#_M1021_g N_Q_c_1895_n 0.0129589f $X=14.42 $Y=2.465 $X2=0
+ $Y2=0
cc_942 N_A_2638_53#_M1034_g N_Q_c_1895_n 0.0137842f $X=14.85 $Y=2.465 $X2=0
+ $Y2=0
cc_943 N_A_2638_53#_c_1385_n N_Q_c_1895_n 0.0388002f $X=14.69 $Y=1.51 $X2=0
+ $Y2=0
cc_944 N_A_2638_53#_c_1387_n N_Q_c_1895_n 0.00259366f $X=15.28 $Y=1.51 $X2=0
+ $Y2=0
cc_945 N_A_2638_53#_M1006_g N_Q_c_1896_n 0.00102666f $X=13.99 $Y=2.465 $X2=0
+ $Y2=0
cc_946 N_A_2638_53#_c_1392_n N_Q_c_1896_n 0.00182356f $X=13.345 $Y=1.98 $X2=0
+ $Y2=0
cc_947 N_A_2638_53#_c_1385_n N_Q_c_1896_n 0.0185589f $X=14.69 $Y=1.51 $X2=0
+ $Y2=0
cc_948 N_A_2638_53#_c_1387_n N_Q_c_1896_n 0.00269667f $X=15.28 $Y=1.51 $X2=0
+ $Y2=0
cc_949 N_A_2638_53#_M1036_g N_Q_c_1892_n 7.99655e-19 $X=14.82 $Y=0.685 $X2=0
+ $Y2=0
cc_950 N_A_2638_53#_M1045_g N_Q_c_1892_n 7.99655e-19 $X=15.25 $Y=0.685 $X2=0
+ $Y2=0
cc_951 N_A_2638_53#_M1044_g N_Q_c_1897_n 0.0135498f $X=15.28 $Y=2.465 $X2=0
+ $Y2=0
cc_952 N_A_2638_53#_c_1387_n N_Q_c_1897_n 6.28182e-19 $X=15.28 $Y=1.51 $X2=0
+ $Y2=0
cc_953 N_A_2638_53#_M1045_g Q 0.0149335f $X=15.25 $Y=0.685 $X2=0 $Y2=0
cc_954 N_A_2638_53#_c_1387_n Q 0.00169954f $X=15.28 $Y=1.51 $X2=0 $Y2=0
cc_955 N_A_2638_53#_M1036_g Q 0.00248442f $X=14.82 $Y=0.685 $X2=0 $Y2=0
cc_956 N_A_2638_53#_M1034_g Q 0.0025759f $X=14.85 $Y=2.465 $X2=0 $Y2=0
cc_957 N_A_2638_53#_M1045_g Q 0.00371777f $X=15.25 $Y=0.685 $X2=0 $Y2=0
cc_958 N_A_2638_53#_M1044_g Q 0.00374525f $X=15.28 $Y=2.465 $X2=0 $Y2=0
cc_959 N_A_2638_53#_c_1385_n Q 0.0134665f $X=14.69 $Y=1.51 $X2=0 $Y2=0
cc_960 N_A_2638_53#_c_1387_n Q 0.0313201f $X=15.28 $Y=1.51 $X2=0 $Y2=0
cc_961 N_A_2638_53#_M1004_g N_VGND_c_1961_n 0.0153316f $X=13.96 $Y=0.685 $X2=0
+ $Y2=0
cc_962 N_A_2638_53#_M1030_g N_VGND_c_1961_n 6.47063e-19 $X=14.39 $Y=0.685 $X2=0
+ $Y2=0
cc_963 N_A_2638_53#_c_1384_n N_VGND_c_1961_n 0.0341485f $X=13.315 $Y=0.42 $X2=0
+ $Y2=0
cc_964 N_A_2638_53#_c_1385_n N_VGND_c_1961_n 0.0182975f $X=14.69 $Y=1.51 $X2=0
+ $Y2=0
cc_965 N_A_2638_53#_c_1387_n N_VGND_c_1961_n 9.56069e-19 $X=15.28 $Y=1.51 $X2=0
+ $Y2=0
cc_966 N_A_2638_53#_M1004_g N_VGND_c_1962_n 5.72142e-19 $X=13.96 $Y=0.685 $X2=0
+ $Y2=0
cc_967 N_A_2638_53#_M1030_g N_VGND_c_1962_n 0.0109899f $X=14.39 $Y=0.685 $X2=0
+ $Y2=0
cc_968 N_A_2638_53#_M1036_g N_VGND_c_1962_n 0.0109899f $X=14.82 $Y=0.685 $X2=0
+ $Y2=0
cc_969 N_A_2638_53#_M1045_g N_VGND_c_1962_n 5.72142e-19 $X=15.25 $Y=0.685 $X2=0
+ $Y2=0
cc_970 N_A_2638_53#_M1036_g N_VGND_c_1964_n 5.72142e-19 $X=14.82 $Y=0.685 $X2=0
+ $Y2=0
cc_971 N_A_2638_53#_M1045_g N_VGND_c_1964_n 0.0119765f $X=15.25 $Y=0.685 $X2=0
+ $Y2=0
cc_972 N_A_2638_53#_c_1384_n N_VGND_c_1973_n 0.0177783f $X=13.315 $Y=0.42 $X2=0
+ $Y2=0
cc_973 N_A_2638_53#_M1004_g N_VGND_c_1974_n 0.00461019f $X=13.96 $Y=0.685 $X2=0
+ $Y2=0
cc_974 N_A_2638_53#_M1030_g N_VGND_c_1974_n 0.00461019f $X=14.39 $Y=0.685 $X2=0
+ $Y2=0
cc_975 N_A_2638_53#_M1036_g N_VGND_c_1975_n 0.00461019f $X=14.82 $Y=0.685 $X2=0
+ $Y2=0
cc_976 N_A_2638_53#_M1045_g N_VGND_c_1975_n 0.00461019f $X=15.25 $Y=0.685 $X2=0
+ $Y2=0
cc_977 N_A_2638_53#_M1004_g N_VGND_c_1982_n 0.00820187f $X=13.96 $Y=0.685 $X2=0
+ $Y2=0
cc_978 N_A_2638_53#_M1030_g N_VGND_c_1982_n 0.00820187f $X=14.39 $Y=0.685 $X2=0
+ $Y2=0
cc_979 N_A_2638_53#_M1036_g N_VGND_c_1982_n 0.00820187f $X=14.82 $Y=0.685 $X2=0
+ $Y2=0
cc_980 N_A_2638_53#_M1045_g N_VGND_c_1982_n 0.00820187f $X=15.25 $Y=0.685 $X2=0
+ $Y2=0
cc_981 N_A_2638_53#_c_1384_n N_VGND_c_1982_n 0.00964167f $X=13.315 $Y=0.42 $X2=0
+ $Y2=0
cc_982 N_A_27_479#_c_1486_n N_VPWR_M1038_d 0.00174003f $X=1.87 $Y=2.41 $X2=-0.19
+ $Y2=1.655
cc_983 N_A_27_479#_c_1485_n N_VPWR_c_1513_n 0.0146197f $X=0.26 $Y=2.54 $X2=0
+ $Y2=0
cc_984 N_A_27_479#_c_1486_n N_VPWR_c_1513_n 0.0166947f $X=1.87 $Y=2.41 $X2=0
+ $Y2=0
cc_985 N_A_27_479#_c_1485_n N_VPWR_c_1530_n 0.0156069f $X=0.26 $Y=2.54 $X2=0
+ $Y2=0
cc_986 N_A_27_479#_c_1485_n N_VPWR_c_1512_n 0.0098998f $X=0.26 $Y=2.54 $X2=0
+ $Y2=0
cc_987 N_A_27_479#_c_1486_n N_VPWR_c_1512_n 0.0229403f $X=1.87 $Y=2.41 $X2=0
+ $Y2=0
cc_988 N_A_27_479#_c_1486_n A_196_479# 0.00192185f $X=1.87 $Y=2.41 $X2=-0.19
+ $Y2=1.655
cc_989 N_A_27_479#_c_1486_n N_A_218_119#_M1017_d 0.00305746f $X=1.87 $Y=2.41
+ $X2=0 $Y2=0
cc_990 N_A_27_479#_M1031_d N_A_218_119#_c_1702_n 0.00312078f $X=1.88 $Y=2.395
+ $X2=0 $Y2=0
cc_991 N_A_27_479#_c_1486_n N_A_218_119#_c_1702_n 0.0189886f $X=1.87 $Y=2.41
+ $X2=0 $Y2=0
cc_992 N_A_27_479#_c_1486_n N_A_218_119#_c_1703_n 0.0137631f $X=1.87 $Y=2.41
+ $X2=0 $Y2=0
cc_993 N_A_27_479#_c_1486_n N_A_218_119#_c_1699_n 0.0032276f $X=1.87 $Y=2.41
+ $X2=0 $Y2=0
cc_994 N_A_27_479#_c_1486_n N_A_218_119#_c_1706_n 0.0143997f $X=1.87 $Y=2.41
+ $X2=0 $Y2=0
cc_995 N_A_27_479#_c_1486_n N_A_218_119#_c_1712_n 0.021058f $X=1.87 $Y=2.41
+ $X2=0 $Y2=0
cc_996 N_VPWR_c_1514_n N_A_218_119#_c_1702_n 0.0143733f $X=2.76 $Y=2.89 $X2=0
+ $Y2=0
cc_997 N_VPWR_c_1526_n N_A_218_119#_c_1702_n 0.0504536f $X=2.645 $Y=3.33 $X2=0
+ $Y2=0
cc_998 N_VPWR_c_1512_n N_A_218_119#_c_1702_n 0.0286242f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_999 N_VPWR_c_1514_n N_A_218_119#_c_1703_n 0.0134868f $X=2.76 $Y=2.89 $X2=0
+ $Y2=0
cc_1000 N_VPWR_M1039_s N_A_218_119#_c_1705_n 0.00853092f $X=2.635 $Y=2.405 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1514_n N_A_218_119#_c_1705_n 0.0164692f $X=2.76 $Y=2.89 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1512_n N_A_218_119#_c_1705_n 0.0069784f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1512_n N_A_218_119#_c_1706_n 0.00626065f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1004 N_VPWR_M1039_s N_A_218_119#_c_1763_n 0.00489953f $X=2.635 $Y=2.405 $X2=0
+ $Y2=0
cc_1005 N_VPWR_c_1514_n N_A_218_119#_c_1763_n 0.013248f $X=2.76 $Y=2.89 $X2=0
+ $Y2=0
cc_1006 N_VPWR_c_1531_n N_A_218_119#_c_1707_n 0.0637482f $X=4.35 $Y=3.33 $X2=0
+ $Y2=0
cc_1007 N_VPWR_c_1512_n N_A_218_119#_c_1707_n 0.0367243f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1008 N_VPWR_M1039_s N_A_218_119#_c_1708_n 0.00155309f $X=2.635 $Y=2.405 $X2=0
+ $Y2=0
cc_1009 N_VPWR_c_1514_n N_A_218_119#_c_1708_n 0.0141252f $X=2.76 $Y=2.89 $X2=0
+ $Y2=0
cc_1010 N_VPWR_c_1531_n N_A_218_119#_c_1708_n 0.0121122f $X=4.35 $Y=3.33 $X2=0
+ $Y2=0
cc_1011 N_VPWR_c_1512_n N_A_218_119#_c_1708_n 0.00649737f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1012 N_VPWR_M1042_d N_A_218_119#_c_1709_n 0.00348485f $X=4.375 $Y=2.455 $X2=0
+ $Y2=0
cc_1013 N_VPWR_c_1515_n N_A_218_119#_c_1709_n 0.0146238f $X=4.515 $Y=2.96 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1516_n N_A_218_119#_c_1709_n 0.0021031f $X=6.89 $Y=3.33 $X2=0
+ $Y2=0
cc_1015 N_VPWR_c_1531_n N_A_218_119#_c_1709_n 0.0021031f $X=4.35 $Y=3.33 $X2=0
+ $Y2=0
cc_1016 N_VPWR_c_1512_n N_A_218_119#_c_1709_n 0.00986362f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1017 N_VPWR_c_1513_n N_A_218_119#_c_1712_n 0.00696143f $X=0.69 $Y=2.79 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1526_n N_A_218_119#_c_1712_n 0.0226434f $X=2.645 $Y=3.33 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1512_n N_A_218_119#_c_1712_n 0.0125895f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1528_n N_A_1751_379#_c_1843_n 0.00311321f $X=11.34 $Y=3.33
+ $X2=0 $Y2=0
cc_1021 N_VPWR_c_1512_n N_A_1751_379#_c_1843_n 0.00479434f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1512_n N_A_1751_379#_c_1841_n 0.00925731f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1519_n N_A_1858_463#_c_1870_n 0.00128496f $X=11.445 $Y=2.795
+ $X2=0 $Y2=0
cc_1024 N_VPWR_c_1518_n N_A_1858_463#_c_1871_n 0.0125451f $X=8.465 $Y=2.22 $X2=0
+ $Y2=0
cc_1025 N_VPWR_c_1528_n N_A_1858_463#_c_1871_n 0.0957128f $X=11.34 $Y=3.33 $X2=0
+ $Y2=0
cc_1026 N_VPWR_c_1512_n N_A_1858_463#_c_1871_n 0.0629926f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1027 N_VPWR_c_1512_n N_Q_M1006_s 0.00397496f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1028 N_VPWR_c_1512_n N_Q_M1034_s 0.00536646f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1029 N_VPWR_c_1534_n N_Q_c_1931_n 0.0138717f $X=14.47 $Y=3.33 $X2=0 $Y2=0
cc_1030 N_VPWR_c_1512_n N_Q_c_1931_n 0.00886411f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1031 N_VPWR_M1021_d N_Q_c_1895_n 0.00176461f $X=14.495 $Y=1.835 $X2=0 $Y2=0
cc_1032 N_VPWR_c_1523_n N_Q_c_1895_n 0.0170777f $X=14.635 $Y=2.19 $X2=0 $Y2=0
cc_1033 N_VPWR_c_1522_n N_Q_c_1896_n 0.00164686f $X=13.775 $Y=1.98 $X2=0 $Y2=0
cc_1034 N_VPWR_c_1535_n N_Q_c_1936_n 0.0124525f $X=15.33 $Y=3.33 $X2=0 $Y2=0
cc_1035 N_VPWR_c_1512_n N_Q_c_1936_n 0.00730901f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1036 N_VPWR_M1044_d N_Q_c_1897_n 0.00277226f $X=15.355 $Y=1.835 $X2=0 $Y2=0
cc_1037 N_VPWR_c_1525_n N_Q_c_1897_n 0.0243971f $X=15.495 $Y=2.19 $X2=0 $Y2=0
cc_1038 N_A_218_119#_c_1713_n N_VGND_c_1953_n 0.0110409f $X=1.23 $Y=0.805 $X2=0
+ $Y2=0
cc_1039 N_A_218_119#_c_1713_n N_VGND_c_1954_n 0.0110409f $X=1.23 $Y=0.805 $X2=0
+ $Y2=0
cc_1040 N_A_218_119#_c_1697_n N_VGND_c_1954_n 0.017615f $X=2.425 $Y=1.377 $X2=0
+ $Y2=0
cc_1041 N_A_218_119#_c_1713_n N_VGND_c_1969_n 0.00510213f $X=1.23 $Y=0.805 $X2=0
+ $Y2=0
cc_1042 N_A_218_119#_c_1713_n N_VGND_c_1982_n 0.00852361f $X=1.23 $Y=0.805 $X2=0
+ $Y2=0
cc_1043 N_A_1751_379#_c_1841_n N_A_1858_463#_M1026_s 0.00451829f $X=10.3 $Y=2.41
+ $X2=-0.19 $Y2=1.655
cc_1044 N_A_1751_379#_M1002_d N_A_1858_463#_c_1870_n 0.00225132f $X=10.325
+ $Y=1.895 $X2=0 $Y2=0
cc_1045 N_A_1751_379#_c_1840_n N_A_1858_463#_c_1870_n 0.0206917f $X=10.465
+ $Y=2.41 $X2=0 $Y2=0
cc_1046 N_A_1751_379#_c_1841_n N_A_1858_463#_c_1870_n 0.0318747f $X=10.3 $Y=2.41
+ $X2=0 $Y2=0
cc_1047 N_A_1751_379#_c_1841_n N_A_1858_463#_c_1871_n 0.0251505f $X=10.3 $Y=2.41
+ $X2=0 $Y2=0
cc_1048 N_Q_c_1890_n N_VGND_M1030_d 0.00176773f $X=14.94 $Y=1.165 $X2=0 $Y2=0
cc_1049 Q N_VGND_M1045_d 0.00244292f $X=15.035 $Y=1.21 $X2=0 $Y2=0
cc_1050 N_Q_c_1889_n N_VGND_c_1961_n 0.0311127f $X=14.175 $Y=0.42 $X2=0 $Y2=0
cc_1051 N_Q_c_1891_n N_VGND_c_1961_n 0.0031924f $X=14.27 $Y=1.165 $X2=0 $Y2=0
cc_1052 N_Q_c_1889_n N_VGND_c_1962_n 0.0247339f $X=14.175 $Y=0.42 $X2=0 $Y2=0
cc_1053 N_Q_c_1890_n N_VGND_c_1962_n 0.0171443f $X=14.94 $Y=1.165 $X2=0 $Y2=0
cc_1054 N_Q_c_1892_n N_VGND_c_1962_n 0.0247339f $X=15.035 $Y=0.42 $X2=0 $Y2=0
cc_1055 N_Q_c_1892_n N_VGND_c_1964_n 0.0247339f $X=15.035 $Y=0.42 $X2=0 $Y2=0
cc_1056 Q N_VGND_c_1964_n 0.0243971f $X=15.035 $Y=1.21 $X2=0 $Y2=0
cc_1057 N_Q_c_1889_n N_VGND_c_1974_n 0.0134771f $X=14.175 $Y=0.42 $X2=0 $Y2=0
cc_1058 N_Q_c_1892_n N_VGND_c_1975_n 0.0134771f $X=15.035 $Y=0.42 $X2=0 $Y2=0
cc_1059 N_Q_c_1889_n N_VGND_c_1982_n 0.00730901f $X=14.175 $Y=0.42 $X2=0 $Y2=0
cc_1060 N_Q_c_1892_n N_VGND_c_1982_n 0.00730901f $X=15.035 $Y=0.42 $X2=0 $Y2=0
cc_1061 N_VGND_c_1957_n A_1598_125# 0.0021897f $X=8.05 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
