* File: sky130_fd_sc_lp__sdfxbp_lp.pex.spice
* Created: Fri Aug 28 11:30:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_27_409# 1 2 7 9 12 14 15 18 22 26 30 32
+ 33
c61 33 0 1.52718e-19 $X=1.52 $Y=1.33
c62 32 0 1.98757e-19 $X=1.52 $Y=1.33
r63 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.33 $X2=1.52 $Y2=1.33
r64 27 30 4.19346 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.58 $Y=1.25 $X2=0.34
+ $Y2=1.25
r65 26 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.25
+ $X2=1.52 $Y2=1.25
r66 26 27 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.355 $Y=1.25
+ $X2=0.58 $Y2=1.25
r67 22 24 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.225 $Y=2.19
+ $X2=0.225 $Y2=2.9
r68 20 30 2.63236 $w=3.65e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.225 $Y=1.335
+ $X2=0.34 $Y2=1.25
r69 20 22 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=0.225 $Y=1.335
+ $X2=0.225 $Y2=2.19
r70 16 30 2.63236 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=1.165
+ $X2=0.34 $Y2=1.25
r71 16 18 8.22304 $w=4.78e-07 $l=3.3e-07 $layer=LI1_cond $X=0.34 $Y=1.165
+ $X2=0.34 $Y2=0.835
r72 15 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.52 $Y=1.67
+ $X2=1.52 $Y2=1.33
r73 14 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.165
+ $X2=1.52 $Y2=1.33
r74 12 14 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.61 $Y=0.835
+ $X2=1.61 $Y2=1.165
r75 7 15 47.383 $w=2.95e-07 $l=3.2311e-07 $layer=POLY_cond $X=1.59 $Y=1.96
+ $X2=1.52 $Y2=1.67
r76 7 9 120.5 $w=2.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.59 $Y=1.96 $X2=1.59
+ $Y2=2.585
r77 2 24 400 $w=1.7e-07 $l=9.17701e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.265 $Y2=2.9
r78 2 22 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.265 $Y2=2.19
r79 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.625 $X2=0.415 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%D 3 7 11 12 13 16 17
c41 17 0 1.52718e-19 $X=2.09 $Y=1.38
r42 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.09
+ $Y=1.38 $X2=2.09 $Y2=1.38
r43 13 17 9.38418 $w=3.48e-07 $l=2.85e-07 $layer=LI1_cond $X=2.1 $Y=1.665
+ $X2=2.1 $Y2=1.38
r44 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.09 $Y=1.72
+ $X2=2.09 $Y2=1.38
r45 11 12 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.72
+ $X2=2.09 $Y2=1.885
r46 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.215
+ $X2=2.09 $Y2=1.38
r47 7 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.12 $Y=2.585 $X2=2.12
+ $Y2=1.885
r48 3 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2 $Y=0.835 $X2=2
+ $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%SCE 3 7 12 13 14 18 19 21 24 29
c73 29 0 1.98757e-19 $X=0.695 $Y=1.68
r74 27 29 11.6903 $w=2.68e-07 $l=6.5e-08 $layer=POLY_cond $X=0.63 $Y=1.68
+ $X2=0.695 $Y2=1.68
r75 26 27 17.9851 $w=2.68e-07 $l=1e-07 $layer=POLY_cond $X=0.53 $Y=1.68 $X2=0.63
+ $Y2=1.68
r76 24 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.695
+ $Y=1.68 $X2=0.695 $Y2=1.68
r77 19 23 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.59 $Y=1.76
+ $X2=2.59 $Y2=1.635
r78 19 21 204.974 $w=2.5e-07 $l=8.25e-07 $layer=POLY_cond $X=2.59 $Y=1.76
+ $X2=2.59 $Y2=2.585
r79 18 23 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.54 $Y=0.835 $X2=2.54
+ $Y2=1.635
r80 15 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.54 $Y=0.255
+ $X2=2.54 $Y2=0.835
r81 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.465 $Y=0.18
+ $X2=2.54 $Y2=0.255
r82 13 14 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=2.465 $Y=0.18
+ $X2=1.095 $Y2=0.18
r83 10 29 58.4515 $w=2.68e-07 $l=3.99061e-07 $layer=POLY_cond $X=1.02 $Y=1.515
+ $X2=0.695 $Y2=1.68
r84 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.02 $Y=1.515
+ $X2=1.02 $Y2=0.835
r85 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.02 $Y=0.255
+ $X2=1.095 $Y2=0.18
r86 9 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.02 $Y=0.255
+ $X2=1.02 $Y2=0.835
r87 5 27 16.3317 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.515
+ $X2=0.63 $Y2=1.68
r88 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.63 $Y=1.515 $X2=0.63
+ $Y2=0.835
r89 1 26 4.4917 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.845
+ $X2=0.53 $Y2=1.68
r90 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.53 $Y=1.845 $X2=0.53
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%SCD 3 5 7 11 13 16 17
r42 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.12
+ $Y=1.41 $X2=3.12 $Y2=1.41
r43 13 17 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.41
r44 12 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.12 $Y=1.75
+ $X2=3.12 $Y2=1.41
r45 11 16 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.12 $Y=1.395
+ $X2=3.12 $Y2=1.41
r46 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.055 $Y=1.245
+ $X2=3.055 $Y2=1.395
r47 5 12 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.915
+ $X2=3.12 $Y2=1.75
r48 5 7 166.464 $w=2.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.12 $Y=1.915 $X2=3.12
+ $Y2=2.585
r49 3 10 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.9 $Y=0.835 $X2=2.9
+ $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%CLK 3 7 11 13 14 23
c41 7 0 1.86192e-19 $X=4.22 $Y=2.235
r42 22 23 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.22 $Y=1.345 $X2=4.23
+ $Y2=1.345
r43 20 22 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=3.96 $Y=1.345
+ $X2=4.22 $Y2=1.345
r44 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.96
+ $Y=1.345 $X2=3.96 $Y2=1.345
r45 17 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.87 $Y=1.345 $X2=3.96
+ $Y2=1.345
r46 14 21 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.08 $Y=1.345
+ $X2=3.96 $Y2=1.345
r47 13 21 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.6 $Y=1.345
+ $X2=3.96 $Y2=1.345
r48 9 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.18
+ $X2=4.23 $Y2=1.345
r49 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.23 $Y=1.18 $X2=4.23
+ $Y2=0.54
r50 5 22 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.22 $Y=1.51
+ $X2=4.22 $Y2=1.345
r51 5 7 180.129 $w=2.5e-07 $l=7.25e-07 $layer=POLY_cond $X=4.22 $Y=1.51 $X2=4.22
+ $Y2=2.235
r52 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.87 $Y=1.18
+ $X2=3.87 $Y2=1.345
r53 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.87 $Y=1.18 $X2=3.87
+ $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1530_231# 1 2 3 12 16 17 22 25 29 31 33
+ 36 37 39
c94 37 0 1.71737e-19 $X=8.89 $Y=0.98
c95 36 0 8.2274e-20 $X=7.815 $Y=1.32
c96 25 0 1.99622e-19 $X=8.91 $Y=1.88
c97 22 0 1.23651e-19 $X=8.87 $Y=0.835
r98 36 40 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.815 $Y=1.32
+ $X2=7.815 $Y2=1.485
r99 36 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.815 $Y=1.32
+ $X2=7.815 $Y2=1.155
r100 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.815
+ $Y=1.32 $X2=7.815 $Y2=1.32
r101 33 35 16.0154 $w=2.59e-07 $l=3.4e-07 $layer=LI1_cond $X=7.815 $Y=0.98
+ $X2=7.815 $Y2=1.32
r102 29 31 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=9.075 $Y=0.35
+ $X2=10.41 $Y2=0.35
r103 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.91 $Y=1.88
+ $X2=8.91 $Y2=2.59
r104 23 37 2.73602 $w=3.5e-07 $l=9.44722e-08 $layer=LI1_cond $X=8.91 $Y=1.065
+ $X2=8.89 $Y2=0.98
r105 23 25 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=8.91 $Y=1.065
+ $X2=8.91 $Y2=1.88
r106 20 37 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=0.895
+ $X2=8.89 $Y2=0.98
r107 20 22 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=8.89 $Y=0.895
+ $X2=8.89 $Y2=0.835
r108 19 29 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=8.89 $Y=0.435
+ $X2=9.075 $Y2=0.35
r109 19 22 12.4588 $w=3.68e-07 $l=4e-07 $layer=LI1_cond $X=8.89 $Y=0.435
+ $X2=8.89 $Y2=0.835
r110 18 33 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.98 $Y=0.98
+ $X2=7.815 $Y2=0.98
r111 17 37 4.03347 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.705 $Y=0.98
+ $X2=8.89 $Y2=0.98
r112 17 18 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.705 $Y=0.98
+ $X2=7.98 $Y2=0.98
r113 16 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.735 $Y=0.835
+ $X2=7.735 $Y2=1.155
r114 12 40 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=7.775 $Y=2.235
+ $X2=7.775 $Y2=1.485
r115 3 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.735 $X2=8.91 $Y2=2.59
r116 3 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.735 $X2=8.91 $Y2=1.88
r117 2 31 182 $w=1.7e-07 $l=5.17446e-07 $layer=licon1_NDIFF $count=1 $X=10.205
+ $Y=0.775 $X2=10.41 $Y2=0.35
r118 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.73
+ $Y=0.625 $X2=8.87 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1278_155# 1 2 9 13 17 21 25 29 30 33 42
c79 33 0 1.03056e-19 $X=8.385 $Y=1.41
c80 30 0 8.2274e-20 $X=7.185 $Y=1.75
r81 41 42 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=8.645 $Y=1.41
+ $X2=8.655 $Y2=1.41
r82 34 41 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=8.385 $Y=1.41
+ $X2=8.645 $Y2=1.41
r83 34 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.385 $Y=1.41
+ $X2=8.295 $Y2=1.41
r84 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.385
+ $Y=1.41 $X2=8.385 $Y2=1.41
r85 31 33 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=8.385 $Y=1.665
+ $X2=8.385 $Y2=1.41
r86 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.22 $Y=1.75
+ $X2=8.385 $Y2=1.665
r87 29 30 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=8.22 $Y=1.75
+ $X2=7.185 $Y2=1.75
r88 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.02 $Y=1.88 $X2=7.02
+ $Y2=2.59
r89 23 30 9.0585 $w=2.8e-07 $l=2.5446e-07 $layer=LI1_cond $X=7.02 $Y=1.565
+ $X2=7.185 $Y2=1.75
r90 23 25 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.02 $Y=1.835
+ $X2=7.02 $Y2=1.88
r91 19 23 20.9143 $w=2.8e-07 $l=4.8e-07 $layer=LI1_cond $X=6.54 $Y=1.565
+ $X2=7.02 $Y2=1.565
r92 19 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.54 $Y=1.395
+ $X2=6.54 $Y2=1.05
r93 15 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=1.245
+ $X2=8.655 $Y2=1.41
r94 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.655 $Y=1.245
+ $X2=8.655 $Y2=0.835
r95 11 41 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.575
+ $X2=8.645 $Y2=1.41
r96 11 13 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.645 $Y=1.575
+ $X2=8.645 $Y2=2.235
r97 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.295 $Y=1.245
+ $X2=8.295 $Y2=1.41
r98 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.295 $Y=1.245
+ $X2=8.295 $Y2=0.835
r99 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.88
+ $Y=1.735 $X2=7.02 $Y2=2.59
r100 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.88
+ $Y=1.735 $X2=7.02 $Y2=1.88
r101 1 21 182 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_NDIFF $count=1 $X=6.39
+ $Y=0.775 $X2=6.54 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_706_66# 1 2 7 9 12 17 18 19 22 24 26 28
+ 32 35 38 40 42 43 44 45 49 53 55 59 60 62 67
c157 59 0 1.87063e-19 $X=4.375 $Y=0.915
c158 40 0 3.23273e-19 $X=9.635 $Y=1.27
c159 35 0 1.03056e-19 $X=9.145 $Y=1.27
c160 22 0 1.25733e-20 $X=6.755 $Y=0.985
r161 67 70 66.9034 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=4.84 $Y=1.025
+ $X2=4.84 $Y2=1.53
r162 66 68 17.3374 $w=5.33e-07 $l=5.05e-07 $layer=LI1_cond $X=4.642 $Y=1.025
+ $X2=4.642 $Y2=1.53
r163 66 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.75
+ $Y=1.025 $X2=4.75 $Y2=1.025
r164 62 68 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.46 $Y=1.715
+ $X2=4.46 $Y2=1.53
r165 59 66 2.45923 $w=5.33e-07 $l=1.1e-07 $layer=LI1_cond $X=4.642 $Y=0.915
+ $X2=4.642 $Y2=1.025
r166 59 60 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.375 $Y=0.915
+ $X2=3.82 $Y2=0.915
r167 55 62 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.375 $Y=1.845
+ $X2=4.46 $Y2=1.715
r168 55 57 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=4.375 $Y=1.845
+ $X2=3.955 $Y2=1.845
r169 51 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.655 $Y=0.83
+ $X2=3.82 $Y2=0.915
r170 51 53 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.655 $Y=0.83
+ $X2=3.655 $Y2=0.54
r171 40 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.635 $Y=1.27
+ $X2=9.635 $Y2=1.345
r172 40 42 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.635 $Y=1.27
+ $X2=9.635 $Y2=0.985
r173 36 49 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=9.385 $Y=1.345
+ $X2=9.635 $Y2=1.345
r174 36 46 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.385 $Y=1.345
+ $X2=9.145 $Y2=1.345
r175 36 38 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.385 $Y=1.42
+ $X2=9.385 $Y2=2.235
r176 35 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.145 $Y=1.27
+ $X2=9.145 $Y2=1.345
r177 34 35 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=9.145 $Y=0.255
+ $X2=9.145 $Y2=1.27
r178 33 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.32 $Y=0.18
+ $X2=7.245 $Y2=0.18
r179 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.07 $Y=0.18
+ $X2=9.145 $Y2=0.255
r180 32 33 897.34 $w=1.5e-07 $l=1.75e-06 $layer=POLY_cond $X=9.07 $Y=0.18
+ $X2=7.32 $Y2=0.18
r181 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.245 $Y=0.255
+ $X2=7.245 $Y2=0.18
r182 30 44 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=7.245 $Y=0.255
+ $X2=7.245 $Y2=1.27
r183 26 44 39.2742 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.285 $Y=1.395
+ $X2=7.285 $Y2=1.27
r184 26 28 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.285 $Y=1.395
+ $X2=7.285 $Y2=2.235
r185 25 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.83 $Y=0.18
+ $X2=6.755 $Y2=0.18
r186 24 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.17 $Y=0.18
+ $X2=7.245 $Y2=0.18
r187 24 25 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.17 $Y=0.18
+ $X2=6.83 $Y2=0.18
r188 20 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.755 $Y=0.255
+ $X2=6.755 $Y2=0.18
r189 20 22 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=6.755 $Y=0.255
+ $X2=6.755 $Y2=0.985
r190 18 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.68 $Y=0.18
+ $X2=6.755 $Y2=0.18
r191 18 19 812.734 $w=1.5e-07 $l=1.585e-06 $layer=POLY_cond $X=6.68 $Y=0.18
+ $X2=5.095 $Y2=0.18
r192 15 67 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=5.02 $Y=0.86
+ $X2=4.84 $Y2=1.025
r193 15 17 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.02 $Y=0.86
+ $X2=5.02 $Y2=0.54
r194 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.02 $Y=0.255
+ $X2=5.095 $Y2=0.18
r195 14 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.02 $Y=0.255
+ $X2=5.02 $Y2=0.54
r196 12 70 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=4.75 $Y=2.235
+ $X2=4.75 $Y2=1.53
r197 7 67 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=4.66 $Y=0.86
+ $X2=4.84 $Y2=1.025
r198 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.66 $Y=0.86 $X2=4.66
+ $Y2=0.54
r199 2 57 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.735 $X2=3.955 $Y2=1.885
r200 1 53 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.53
+ $Y=0.33 $X2=3.655 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_975_347# 1 2 8 9 10 11 12 13 15 18 20 25
+ 28 32 33 35 36 43 47 48 49
c102 36 0 1.86192e-19 $X=5.23 $Y=1.845
c103 25 0 1.53485e-19 $X=10.075 $Y=2.26
c104 10 0 1.87063e-19 $X=5.665 $Y=1.38
r105 47 50 10.0504 $w=4.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.445 $Y=1.47
+ $X2=5.445 $Y2=1.845
r106 47 49 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.445 $Y=1.47
+ $X2=5.445 $Y2=1.305
r107 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.5
+ $Y=1.47 $X2=5.5 $Y2=1.47
r108 45 49 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.315 $Y=0.65
+ $X2=5.315 $Y2=1.305
r109 43 45 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.235 $Y=0.48
+ $X2=5.235 $Y2=0.65
r110 36 50 3.68054 $w=2.6e-07 $l=2.15e-07 $layer=LI1_cond $X=5.23 $Y=1.845
+ $X2=5.445 $Y2=1.845
r111 36 38 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=5.23 $Y=1.845
+ $X2=5.015 $Y2=1.845
r112 34 35 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=10.077 $Y=1.4
+ $X2=10.077 $Y2=1.55
r113 31 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.5 $Y=1.81 $X2=5.5
+ $Y2=1.47
r114 31 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.81
+ $X2=5.5 $Y2=1.975
r115 30 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.5 $Y=1.455
+ $X2=5.5 $Y2=1.47
r116 28 34 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=10.13 $Y=0.985
+ $X2=10.13 $Y2=1.4
r117 25 35 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=10.075 $Y=2.26
+ $X2=10.075 $Y2=1.55
r118 23 25 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=10.075 $Y=3.075
+ $X2=10.075 $Y2=2.26
r119 21 33 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.88 $Y=3.15
+ $X2=6.755 $Y2=3.15
r120 20 23 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=9.95 $Y=3.15
+ $X2=10.075 $Y2=3.075
r121 20 21 1574.19 $w=1.5e-07 $l=3.07e-06 $layer=POLY_cond $X=9.95 $Y=3.15
+ $X2=6.88 $Y2=3.15
r122 16 33 1.63566 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.755 $Y=3.075
+ $X2=6.755 $Y2=3.15
r123 16 18 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.755 $Y=3.075
+ $X2=6.755 $Y2=2.235
r124 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.315 $Y=1.305
+ $X2=6.315 $Y2=0.985
r125 11 33 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.63 $Y=3.15
+ $X2=6.755 $Y2=3.15
r126 11 12 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=6.63 $Y=3.15
+ $X2=5.665 $Y2=3.15
r127 10 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.665 $Y=1.38
+ $X2=5.5 $Y2=1.455
r128 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.24 $Y=1.38
+ $X2=6.315 $Y2=1.305
r129 9 10 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.24 $Y=1.38
+ $X2=5.665 $Y2=1.38
r130 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.59 $Y=3.075
+ $X2=5.665 $Y2=3.15
r131 8 32 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=5.59 $Y=3.075
+ $X2=5.59 $Y2=1.975
r132 2 38 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=4.875
+ $Y=1.735 $X2=5.015 $Y2=1.885
r133 1 43 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=5.095
+ $Y=0.33 $X2=5.235 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_2089_254# 1 2 9 12 13 14 17 21 25 29 33
+ 37 41 45 48 49 53 57 58 59 63 69 73 75 77 80 85 96
c170 77 0 6.64951e-20 $X=11.815 $Y=0.945
c171 45 0 1.53485e-19 $X=10.73 $Y=1.435
c172 21 0 4.93603e-20 $X=12.915 $Y=2.505
r173 93 94 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=13.445 $Y=1.64
+ $X2=13.68 $Y2=1.64
r174 87 89 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=12.89 $Y=1.64
+ $X2=12.915 $Y2=1.64
r175 81 91 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=12.98 $Y=1.64
+ $X2=13.25 $Y2=1.64
r176 81 89 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=12.98 $Y=1.64
+ $X2=12.915 $Y2=1.64
r177 80 81 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.98
+ $Y=1.64 $X2=12.98 $Y2=1.64
r178 73 75 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.525 $Y=2.215
+ $X2=11.815 $Y2=2.215
r179 70 96 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=14 $Y=1.64 $X2=14.04
+ $Y2=1.64
r180 70 94 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=14 $Y=1.64
+ $X2=13.68 $Y2=1.64
r181 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=14
+ $Y=1.64 $X2=14 $Y2=1.64
r182 67 93 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=13.32 $Y=1.64
+ $X2=13.445 $Y2=1.64
r183 67 91 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=13.32 $Y=1.64
+ $X2=13.25 $Y2=1.64
r184 66 69 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.32 $Y=1.64
+ $X2=14 $Y2=1.64
r185 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.32
+ $Y=1.64 $X2=13.32 $Y2=1.64
r186 64 80 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.11 $Y=1.64
+ $X2=13.025 $Y2=1.64
r187 64 66 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=13.11 $Y=1.64
+ $X2=13.32 $Y2=1.64
r188 63 80 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.025 $Y=1.475
+ $X2=13.025 $Y2=1.64
r189 62 63 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=13.025 $Y=0.435
+ $X2=13.025 $Y2=1.475
r190 58 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.94 $Y=0.35
+ $X2=13.025 $Y2=0.435
r191 58 59 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=12.94 $Y=0.35
+ $X2=12.32 $Y2=0.35
r192 55 77 18.5179 $w=2.24e-07 $l=3.4e-07 $layer=LI1_cond $X=12.155 $Y=0.945
+ $X2=11.815 $Y2=0.945
r193 55 57 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=12.155 $Y=0.775
+ $X2=12.155 $Y2=0.495
r194 54 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.155 $Y=0.435
+ $X2=12.32 $Y2=0.35
r195 54 57 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=12.155 $Y=0.435
+ $X2=12.155 $Y2=0.495
r196 53 75 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.815 $Y=2.13
+ $X2=11.815 $Y2=2.215
r197 52 77 2.3549 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.815 $Y=1.135
+ $X2=11.815 $Y2=0.945
r198 52 53 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=11.815 $Y=1.135
+ $X2=11.815 $Y2=2.13
r199 48 77 5.36773 $w=2.24e-07 $l=1.41244e-07 $layer=LI1_cond $X=11.73 $Y=1.05
+ $X2=11.815 $Y2=0.945
r200 48 49 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=11.73 $Y=1.05
+ $X2=10.895 $Y2=1.05
r201 46 85 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.73 $Y=1.435
+ $X2=10.82 $Y2=1.435
r202 46 82 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=10.73 $Y=1.435
+ $X2=10.57 $Y2=1.435
r203 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.73
+ $Y=1.435 $X2=10.73 $Y2=1.435
r204 43 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.73 $Y=1.135
+ $X2=10.895 $Y2=1.05
r205 43 45 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=10.73 $Y=1.135
+ $X2=10.73 $Y2=1.435
r206 39 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.04 $Y=1.475
+ $X2=14.04 $Y2=1.64
r207 39 41 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=14.04 $Y=1.475
+ $X2=14.04 $Y2=0.845
r208 35 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.68 $Y=1.475
+ $X2=13.68 $Y2=1.64
r209 35 37 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=13.68 $Y=1.475
+ $X2=13.68 $Y2=0.845
r210 31 93 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.445 $Y=1.805
+ $X2=13.445 $Y2=1.64
r211 31 33 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=13.445 $Y=1.805
+ $X2=13.445 $Y2=2.505
r212 27 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.25 $Y=1.475
+ $X2=13.25 $Y2=1.64
r213 27 29 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=13.25 $Y=1.475
+ $X2=13.25 $Y2=0.845
r214 23 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.89 $Y=1.475
+ $X2=12.89 $Y2=1.64
r215 23 25 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=12.89 $Y=1.475
+ $X2=12.89 $Y2=0.845
r216 19 89 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.915 $Y=1.805
+ $X2=12.915 $Y2=1.64
r217 19 21 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=12.915 $Y=1.805
+ $X2=12.915 $Y2=2.505
r218 15 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.15 $Y=0.925
+ $X2=11.15 $Y2=0.495
r219 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.075 $Y=1
+ $X2=11.15 $Y2=0.925
r220 13 14 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=11.075 $Y=1
+ $X2=10.895 $Y2=1
r221 12 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.82 $Y=1.27
+ $X2=10.82 $Y2=1.435
r222 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.82 $Y=1.075
+ $X2=10.895 $Y2=1
r223 11 12 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=10.82 $Y=1.075
+ $X2=10.82 $Y2=1.27
r224 7 82 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.57 $Y=1.6
+ $X2=10.57 $Y2=1.435
r225 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.57 $Y=1.6
+ $X2=10.57 $Y2=2.26
r226 2 73 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=11.385
+ $Y=1.805 $X2=11.525 $Y2=2.295
r227 1 57 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.015
+ $Y=0.285 $X2=12.155 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1902_347# 1 2 9 11 13 15 16 18 20 21 24
+ 28 30 34 41 45
c91 11 0 1.74055e-19 $X=11.58 $Y=0.78
r92 35 45 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=11.385 $Y=1.48
+ $X2=11.58 $Y2=1.48
r93 35 42 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=11.385 $Y=1.48
+ $X2=11.26 $Y2=1.48
r94 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.385
+ $Y=1.48 $X2=11.385 $Y2=1.48
r95 32 34 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=11.385 $Y=1.78
+ $X2=11.385 $Y2=1.48
r96 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.22 $Y=1.865
+ $X2=11.385 $Y2=1.78
r97 30 41 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=11.22 $Y=1.865
+ $X2=10.08 $Y2=1.865
r98 26 41 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=9.915 $Y=1.832
+ $X2=10.08 $Y2=1.832
r99 26 38 9.07242 $w=2.33e-07 $l=1.85e-07 $layer=LI1_cond $X=9.915 $Y=1.832
+ $X2=9.73 $Y2=1.832
r100 26 28 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=9.915 $Y=1.715
+ $X2=9.915 $Y2=1.05
r101 24 38 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=9.73 $Y=2.615
+ $X2=9.73 $Y2=1.95
r102 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.94 $Y=0.78
+ $X2=11.94 $Y2=0.495
r103 17 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.655 $Y=0.855
+ $X2=11.58 $Y2=0.855
r104 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.865 $Y=0.855
+ $X2=11.94 $Y2=0.78
r105 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=11.865 $Y=0.855
+ $X2=11.655 $Y2=0.855
r106 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.58 $Y=1.315
+ $X2=11.58 $Y2=1.48
r107 14 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.58 $Y=0.93
+ $X2=11.58 $Y2=0.855
r108 14 15 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=11.58 $Y=0.93
+ $X2=11.58 $Y2=1.315
r109 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.58 $Y=0.78
+ $X2=11.58 $Y2=0.855
r110 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.58 $Y=0.78
+ $X2=11.58 $Y2=0.495
r111 7 42 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.26 $Y=1.645
+ $X2=11.26 $Y2=1.48
r112 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.26 $Y=1.645
+ $X2=11.26 $Y2=2.305
r113 2 38 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=9.51
+ $Y=1.735 $X2=9.73 $Y2=1.88
r114 2 24 400 $w=1.7e-07 $l=9.8387e-07 $layer=licon1_PDIFF $count=1 $X=9.51
+ $Y=1.735 $X2=9.73 $Y2=2.615
r115 1 28 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=9.71
+ $Y=0.775 $X2=9.915 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_2714_401# 1 2 9 13 15 19 21 23 25 27 28
+ 30 38 39
c64 21 0 4.93603e-20 $X=13.71 $Y=2.155
r65 39 40 40.8095 $w=5.85e-07 $l=7.5e-08 $layer=POLY_cond $X=14.782 $Y=0.98
+ $X2=14.782 $Y2=0.905
r66 37 42 64.0993 $w=5.85e-07 $l=5.05e-07 $layer=POLY_cond $X=14.782 $Y=1.07
+ $X2=14.782 $Y2=1.575
r67 37 39 8.23122 $w=5.85e-07 $l=9e-08 $layer=POLY_cond $X=14.782 $Y=1.07
+ $X2=14.782 $Y2=0.98
r68 30 38 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=14.43 $Y=1.985
+ $X2=14.43 $Y2=1.575
r69 28 38 11.2652 $w=4.78e-07 $l=2.4e-07 $layer=LI1_cond $X=14.585 $Y=1.335
+ $X2=14.585 $Y2=1.575
r70 27 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.66
+ $Y=1.07 $X2=14.66 $Y2=1.07
r71 27 34 13.42 $w=3e-07 $l=4.61357e-07 $layer=LI1_cond $X=14.585 $Y=1.075
+ $X2=14.255 $Y2=0.76
r72 27 28 6.47876 $w=4.78e-07 $l=2.6e-07 $layer=LI1_cond $X=14.585 $Y=1.075
+ $X2=14.585 $Y2=1.335
r73 26 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.875 $Y=2.07
+ $X2=13.71 $Y2=2.07
r74 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.345 $Y=2.07
+ $X2=14.43 $Y2=1.985
r75 25 26 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=14.345 $Y=2.07
+ $X2=13.875 $Y2=2.07
r76 21 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.71 $Y=2.155
+ $X2=13.71 $Y2=2.07
r77 21 23 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=13.71 $Y=2.155
+ $X2=13.71 $Y2=2.86
r78 17 19 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=15.36 $Y=0.905
+ $X2=15.36 $Y2=0.495
r79 16 39 35.4195 $w=1.5e-07 $l=2.93e-07 $layer=POLY_cond $X=15.075 $Y=0.98
+ $X2=14.782 $Y2=0.98
r80 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.285 $Y=0.98
+ $X2=15.36 $Y2=0.905
r81 15 16 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=15.285 $Y=0.98
+ $X2=15.075 $Y2=0.98
r82 13 40 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=15 $Y=0.495 $X2=15
+ $Y2=0.905
r83 9 42 241 $w=2.5e-07 $l=9.7e-07 $layer=POLY_cond $X=14.615 $Y=2.545
+ $X2=14.615 $Y2=1.575
r84 2 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.57
+ $Y=2.005 $X2=13.71 $Y2=2.15
r85 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=13.57
+ $Y=2.005 $X2=13.71 $Y2=2.86
r86 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.115
+ $Y=0.635 $X2=14.255 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%VPWR 1 2 3 4 5 6 7 24 30 34 38 42 46 52 55
+ 56 58 59 60 62 74 81 86 91 107 108 111 114 117 120 123
r133 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r134 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r135 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r138 105 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.6 $Y2=3.33
r139 104 107 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=14.64 $Y=3.33
+ $X2=15.6 $Y2=3.33
r140 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r141 102 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r142 102 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.2 $Y2=3.33
r143 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r144 99 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.345 $Y=3.33
+ $X2=13.18 $Y2=3.33
r145 99 101 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=13.345 $Y=3.33
+ $X2=14.16 $Y2=3.33
r146 98 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r147 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r148 95 98 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.72 $Y2=3.33
r149 95 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r150 94 97 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.72 $Y2=3.33
r151 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r152 92 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.08 $Y=3.33
+ $X2=10.915 $Y2=3.33
r153 92 94 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=11.08 $Y=3.33
+ $X2=11.28 $Y2=3.33
r154 91 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.015 $Y=3.33
+ $X2=13.18 $Y2=3.33
r155 91 97 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.015 $Y=3.33
+ $X2=12.72 $Y2=3.33
r156 90 121 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r157 89 90 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r158 87 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=3.33
+ $X2=8.04 $Y2=3.33
r159 87 89 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.205 $Y=3.33
+ $X2=8.4 $Y2=3.33
r160 86 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.75 $Y=3.33
+ $X2=10.915 $Y2=3.33
r161 86 89 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=10.75 $Y=3.33
+ $X2=8.4 $Y2=3.33
r162 85 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r163 84 85 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r164 82 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=4.485 $Y2=3.33
r165 82 84 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=5.04 $Y2=3.33
r166 81 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=3.33
+ $X2=8.04 $Y2=3.33
r167 81 84 184.957 $w=1.68e-07 $l=2.835e-06 $layer=LI1_cond $X=7.875 $Y=3.33
+ $X2=5.04 $Y2=3.33
r168 80 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r169 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r170 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r171 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r172 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r173 74 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.485 $Y2=3.33
r174 74 79 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r176 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r177 70 73 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r178 70 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 69 72 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r180 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r181 67 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=0.795 $Y2=3.33
r182 67 69 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r183 65 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r185 62 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=3.33
+ $X2=0.795 $Y2=3.33
r186 62 64 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=3.33
+ $X2=0.24 $Y2=3.33
r187 60 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r188 60 85 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=5.04 $Y2=3.33
r189 60 117 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r190 58 101 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=14.185 $Y=3.33
+ $X2=14.16 $Y2=3.33
r191 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.185 $Y=3.33
+ $X2=14.35 $Y2=3.33
r192 57 104 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=14.515 $Y=3.33
+ $X2=14.64 $Y2=3.33
r193 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.515 $Y=3.33
+ $X2=14.35 $Y2=3.33
r194 55 72 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=3.33 $X2=2.64
+ $Y2=3.33
r195 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.855 $Y2=3.33
r196 54 76 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=3.33 $X2=3.12
+ $Y2=3.33
r197 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.855 $Y2=3.33
r198 50 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.35 $Y=3.245
+ $X2=14.35 $Y2=3.33
r199 50 52 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=14.35 $Y=3.245
+ $X2=14.35 $Y2=2.5
r200 46 49 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=13.18 $Y=2.15
+ $X2=13.18 $Y2=2.86
r201 44 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.18 $Y=3.245
+ $X2=13.18 $Y2=3.33
r202 44 49 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=13.18 $Y=3.245
+ $X2=13.18 $Y2=2.86
r203 40 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.915 $Y=3.245
+ $X2=10.915 $Y2=3.33
r204 40 42 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=10.915 $Y=3.245
+ $X2=10.915 $Y2=2.295
r205 36 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=3.245
+ $X2=8.04 $Y2=3.33
r206 36 38 37.1925 $w=3.28e-07 $l=1.065e-06 $layer=LI1_cond $X=8.04 $Y=3.245
+ $X2=8.04 $Y2=2.18
r207 32 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=3.33
r208 32 34 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=2.59
r209 28 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=3.33
r210 28 30 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=2.94
r211 24 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.795 $Y=2.19
+ $X2=0.795 $Y2=2.9
r212 22 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=3.245
+ $X2=0.795 $Y2=3.33
r213 22 27 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.795 $Y=3.245
+ $X2=0.795 $Y2=2.9
r214 7 52 300 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=2 $X=14.205
+ $Y=2.045 $X2=14.35 $Y2=2.5
r215 6 49 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=13.04
+ $Y=2.005 $X2=13.18 $Y2=2.86
r216 6 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.04
+ $Y=2.005 $X2=13.18 $Y2=2.15
r217 5 42 300 $w=1.7e-07 $l=6.35551e-07 $layer=licon1_PDIFF $count=2 $X=10.695
+ $Y=1.76 $X2=10.915 $Y2=2.295
r218 4 38 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=7.9
+ $Y=1.735 $X2=8.04 $Y2=2.18
r219 3 34 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.735 $X2=4.485 $Y2=2.59
r220 2 30 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=2.085 $X2=2.855 $Y2=2.94
r221 1 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=2.045 $X2=0.795 $Y2=2.9
r222 1 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=2.045 $X2=0.795 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_239_417# 1 2 9 13 17 19
r41 15 17 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.385 $Y=2.675
+ $X2=3.385 $Y2=2.785
r42 14 19 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=2.59
+ $X2=1.325 $Y2=2.59
r43 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.22 $Y=2.59
+ $X2=3.385 $Y2=2.675
r44 13 14 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=3.22 $Y=2.59
+ $X2=1.49 $Y2=2.59
r45 7 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=2.505
+ $X2=1.325 $Y2=2.59
r46 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.325 $Y=2.505
+ $X2=1.325 $Y2=2.23
r47 2 17 600 $w=1.7e-07 $l=7.66812e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=2.085 $X2=3.385 $Y2=2.785
r48 1 9 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=1.195
+ $Y=2.085 $X2=1.325 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_343_417# 1 2 3 4 13 18 19 23 24 27 32 34
+ 36 37
c99 37 0 1.25733e-20 $X=6.34 $Y=1.745
c100 24 0 1.33018e-19 $X=6.195 $Y=0.7
r101 38 40 6.64488 $w=6.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.34 $Y=2.24
+ $X2=6.34 $Y2=2.59
r102 36 38 6.26517 $w=6.28e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=1.91
+ $X2=6.34 $Y2=2.24
r103 36 37 10.3517 $w=6.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=1.91
+ $X2=6.34 $Y2=1.745
r104 30 32 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.325 $Y=0.82
+ $X2=2.54 $Y2=0.82
r105 25 27 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=7.01 $Y=0.785
+ $X2=7.01 $Y2=0.985
r106 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.885 $Y=0.7
+ $X2=7.01 $Y2=0.785
r107 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.885 $Y=0.7
+ $X2=6.195 $Y2=0.7
r108 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.11 $Y=0.785
+ $X2=6.195 $Y2=0.7
r109 21 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.11 $Y=0.785
+ $X2=6.11 $Y2=1.745
r110 20 34 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=2.625 $Y=2.24
+ $X2=2.54 $Y2=2.195
r111 19 38 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=6.025 $Y=2.24
+ $X2=6.34 $Y2=2.24
r112 19 20 221.818 $w=1.68e-07 $l=3.4e-06 $layer=LI1_cond $X=6.025 $Y=2.24
+ $X2=2.625 $Y2=2.24
r113 18 34 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=2.065
+ $X2=2.54 $Y2=2.195
r114 17 32 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.54 $Y=1.035
+ $X2=2.54 $Y2=0.82
r115 17 18 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.54 $Y=1.035
+ $X2=2.54 $Y2=2.065
r116 13 34 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=2.195
+ $X2=2.54 $Y2=2.195
r117 13 15 26.5948 $w=2.58e-07 $l=6e-07 $layer=LI1_cond $X=2.455 $Y=2.195
+ $X2=1.855 $Y2=2.195
r118 4 40 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=1.735 $X2=6.49 $Y2=2.59
r119 4 36 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=1.735 $X2=6.49 $Y2=1.91
r120 3 15 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=2.085 $X2=1.855 $Y2=2.235
r121 2 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.83
+ $Y=0.775 $X2=6.97 $Y2=0.985
r122 1 30 182 $w=1.7e-07 $l=3.33542e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.625 $X2=2.325 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%Q 1 2 9 10 13 15 16 24 25
r35 24 25 10.8692 $w=7.08e-07 $l=1.65e-07 $layer=LI1_cond $X=12.48 $Y=2.15
+ $X2=12.48 $Y2=1.985
r36 15 16 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=12.48 $Y=2.405
+ $X2=12.48 $Y2=2.775
r37 15 24 4.29577 $w=7.08e-07 $l=2.55e-07 $layer=LI1_cond $X=12.48 $Y=2.405
+ $X2=12.48 $Y2=2.15
r38 11 13 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=12.635 $Y=1.125
+ $X2=12.635 $Y2=0.845
r39 9 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.51 $Y=1.21
+ $X2=12.635 $Y2=1.125
r40 9 10 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=12.51 $Y=1.21
+ $X2=12.295 $Y2=1.21
r41 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.21 $Y=1.295
+ $X2=12.295 $Y2=1.21
r42 7 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.21 $Y=1.295
+ $X2=12.21 $Y2=1.985
r43 2 16 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.505
+ $Y=2.005 $X2=12.65 $Y2=2.86
r44 2 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.505
+ $Y=2.005 $X2=12.65 $Y2=2.15
r45 1 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=12.55
+ $Y=0.635 $X2=12.675 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%Q_N 1 2 9 11 12 13
r21 13 36 1.4878 $w=1.023e-06 $l=1.25e-07 $layer=LI1_cond $X=15.227 $Y=2.775
+ $X2=15.227 $Y2=2.9
r22 12 13 4.4039 $w=1.023e-06 $l=3.7e-07 $layer=LI1_cond $X=15.227 $Y=2.405
+ $X2=15.227 $Y2=2.775
r23 12 28 2.55902 $w=1.023e-06 $l=2.15e-07 $layer=LI1_cond $X=15.227 $Y=2.405
+ $X2=15.227 $Y2=2.19
r24 11 28 1.84488 $w=1.023e-06 $l=1.55e-07 $layer=LI1_cond $X=15.227 $Y=2.035
+ $X2=15.227 $Y2=2.19
r25 11 24 7.44224 $w=1.023e-06 $l=1.15e-07 $layer=LI1_cond $X=15.227 $Y=2.035
+ $X2=15.227 $Y2=1.92
r26 9 24 49.7646 $w=3.28e-07 $l=1.425e-06 $layer=LI1_cond $X=15.575 $Y=0.495
+ $X2=15.575 $Y2=1.92
r27 2 36 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=14.74
+ $Y=2.045 $X2=14.88 $Y2=2.9
r28 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.74
+ $Y=2.045 $X2=14.88 $Y2=2.19
r29 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.435
+ $Y=0.285 $X2=15.575 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%VGND 1 2 3 4 5 6 7 24 28 32 34 38 42 46 50
+ 53 54 55 57 62 70 75 87 93 94 97 100 103 106 109 112
r158 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r159 109 110 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r160 103 104 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r161 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r162 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r163 94 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=14.64 $Y2=0
r164 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0 $X2=15.6
+ $Y2=0
r165 91 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.95 $Y=0
+ $X2=14.785 $Y2=0
r166 91 93 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=14.95 $Y=0 $X2=15.6
+ $Y2=0
r167 90 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.64 $Y2=0
r168 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r169 87 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.62 $Y=0
+ $X2=14.785 $Y2=0
r170 87 89 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=14.62 $Y=0
+ $X2=13.68 $Y2=0
r171 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r172 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r173 83 86 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r174 83 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r175 82 85 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r176 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r177 80 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.53 $Y=0
+ $X2=11.405 $Y2=0
r178 80 82 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.53 $Y=0
+ $X2=11.76 $Y2=0
r179 79 110 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=11.28 $Y2=0
r180 78 79 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r181 76 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.18 $Y=0
+ $X2=8.015 $Y2=0
r182 76 78 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.18 $Y=0 $X2=8.4
+ $Y2=0
r183 75 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=11.405 $Y2=0
r184 75 78 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=11.28 $Y=0 $X2=8.4
+ $Y2=0
r185 74 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r186 74 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=3.12 $Y2=0
r187 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r188 71 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=0
+ $X2=3.115 $Y2=0
r189 71 73 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=4.08
+ $Y2=0
r190 70 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.28 $Y=0
+ $X2=4.445 $Y2=0
r191 70 73 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.28 $Y=0 $X2=4.08
+ $Y2=0
r192 69 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r193 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r194 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r195 66 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r196 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r197 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r198 63 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.315
+ $Y2=0
r199 63 65 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.68
+ $Y2=0
r200 62 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=0
+ $X2=3.115 $Y2=0
r201 62 68 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.95 $Y=0 $X2=2.64
+ $Y2=0
r202 60 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r203 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r204 57 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.315
+ $Y2=0
r205 57 59 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=0.24
+ $Y2=0
r206 55 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r207 55 104 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=4.56 $Y2=0
r208 55 106 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r209 53 85 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=13.3 $Y=0 $X2=13.2
+ $Y2=0
r210 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.3 $Y=0
+ $X2=13.465 $Y2=0
r211 52 89 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=13.63 $Y=0 $X2=13.68
+ $Y2=0
r212 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.63 $Y=0
+ $X2=13.465 $Y2=0
r213 48 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.785 $Y=0.085
+ $X2=14.785 $Y2=0
r214 48 50 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=14.785 $Y=0.085
+ $X2=14.785 $Y2=0.495
r215 44 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.465 $Y=0.085
+ $X2=13.465 $Y2=0
r216 44 46 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=13.465 $Y=0.085
+ $X2=13.465 $Y2=0.845
r217 40 109 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.405 $Y=0.085
+ $X2=11.405 $Y2=0
r218 40 42 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=11.405 $Y=0.085
+ $X2=11.405 $Y2=0.43
r219 36 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=0.085
+ $X2=8.015 $Y2=0
r220 36 38 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.015 $Y=0.085
+ $X2=8.015 $Y2=0.55
r221 35 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.61 $Y=0
+ $X2=4.445 $Y2=0
r222 34 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.85 $Y=0
+ $X2=8.015 $Y2=0
r223 34 35 211.38 $w=1.68e-07 $l=3.24e-06 $layer=LI1_cond $X=7.85 $Y=0 $X2=4.61
+ $Y2=0
r224 30 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.445 $Y=0.085
+ $X2=4.445 $Y2=0
r225 30 32 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.445 $Y=0.085
+ $X2=4.445 $Y2=0.48
r226 26 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0
r227 26 28 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0.835
r228 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=0.085
+ $X2=1.315 $Y2=0
r229 22 24 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.315 $Y=0.085
+ $X2=1.315 $Y2=0.795
r230 7 50 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=14.655
+ $Y=0.285 $X2=14.785 $Y2=0.495
r231 6 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.325
+ $Y=0.635 $X2=13.465 $Y2=0.845
r232 5 42 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.225
+ $Y=0.285 $X2=11.365 $Y2=0.43
r233 4 38 182 $w=1.7e-07 $l=2.39583e-07 $layer=licon1_NDIFF $count=1 $X=7.81
+ $Y=0.625 $X2=8.015 $Y2=0.55
r234 3 32 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.33 $X2=4.445 $Y2=0.48
r235 2 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.625 $X2=3.115 $Y2=0.835
r236 1 24 182 $w=1.7e-07 $l=2.92916e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.625 $X2=1.315 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1127_155# 1 2 9 11 12 15
c33 1 0 1.33018e-19 $X=5.635 $Y=0.775
r34 13 15 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=7.48 $Y=0.435
+ $X2=7.48 $Y2=0.79
r35 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.355 $Y=0.35
+ $X2=7.48 $Y2=0.435
r36 11 12 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=7.355 $Y=0.35
+ $X2=5.845 $Y2=0.35
r37 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.72 $Y=0.435
+ $X2=5.845 $Y2=0.35
r38 7 9 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=5.72 $Y=0.435
+ $X2=5.72 $Y2=0.94
r39 2 15 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=7.395
+ $Y=0.625 $X2=7.52 $Y2=0.79
r40 1 9 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=5.635
+ $Y=0.775 $X2=5.76 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_LP%A_1859_155# 1 2 9 11 12 15
c35 15 0 1.0756e-19 $X=10.935 $Y=0.495
r36 13 15 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=10.935 $Y=0.615
+ $X2=10.935 $Y2=0.495
r37 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.77 $Y=0.7
+ $X2=10.935 $Y2=0.615
r38 11 12 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=10.77 $Y=0.7
+ $X2=9.505 $Y2=0.7
r39 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.38 $Y=0.785
+ $X2=9.505 $Y2=0.7
r40 7 9 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=9.38 $Y=0.785 $X2=9.38
+ $Y2=0.985
r41 2 15 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=10.805
+ $Y=0.285 $X2=10.935 $Y2=0.495
r42 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=0.775 $X2=9.42 $Y2=0.985
.ends

