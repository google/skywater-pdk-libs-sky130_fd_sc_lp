* File: sky130_fd_sc_lp__o31a_0.spice
* Created: Wed Sep  2 10:24:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31a_0.pex.spice"
.subckt sky130_fd_sc_lp__o31a_0  VNB VPB A1 A2 A3 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_90_309#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1113 PD=0.84 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_270_55#_M1000_d N_A1_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0882 PD=0.78 PS=0.84 NRD=11.424 NRS=19.992 M=1 R=2.8 SA=75000.8
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_270_55#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0756 PD=0.74 PS=0.78 NRD=5.712 NRS=11.424 M=1 R=2.8 SA=75001.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_A_270_55#_M1003_d N_A3_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_90_309#_M1007_d N_B1_M1007_g N_A_270_55#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_90_309#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1424 AS=0.1696 PD=1.085 PS=1.81 NRD=26.1616 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1004 A_270_481# N_A1_M1004_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1424 PD=0.91 PS=1.085 NRD=24.625 NRS=24.6053 M=1 R=4.26667
+ SA=75000.8 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 A_354_481# N_A2_M1002_g A_270_481# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=24.625 M=1 R=4.26667 SA=75001.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_A_90_309#_M1009_d N_A3_M1009_g A_354_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1056 AS=0.0672 PD=0.97 PS=0.85 NRD=3.0732 NRS=15.3857 M=1 R=4.26667
+ SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_A_90_309#_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1888 AS=0.1056 PD=1.87 PS=0.97 NRD=9.2196 NRS=12.2928 M=1 R=4.26667
+ SA=75002 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o31a_0.pxi.spice"
*
.ends
*
*
