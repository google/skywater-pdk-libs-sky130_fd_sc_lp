* NGSPICE file created from sky130_fd_sc_lp__iso1p_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__iso1p_lp2 A SLEEP KAPWR VGND VNB VPB VPWR X
M1000 a_137_409# A a_147_57# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.008e+11p ps=1.32e+06u
M1001 a_469_57# a_137_409# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.373e+11p ps=2.81e+06u
M1002 X a_137_409# a_469_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 a_240_409# A a_137_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.1e+11p pd=2.42e+06u as=2.65e+11p ps=2.53e+06u
M1004 KAPWR SLEEP a_240_409# VPB phighvt w=1e+06u l=250000u
+  ad=6.2e+11p pd=3.24e+06u as=0p ps=0u
M1005 X a_137_409# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1006 a_147_57# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_311_57# SLEEP a_137_409# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 VGND SLEEP a_311_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

