* File: sky130_fd_sc_lp__a31o_0.spice
* Created: Fri Aug 28 09:58:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31o_0.pex.spice"
.subckt sky130_fd_sc_lp__a31o_0  VNB VPB A3 A2 A1 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_86_241#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1006 A_272_50# N_A3_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.06195
+ AS=0.1113 PD=0.715 PS=0.95 NRD=26.424 NRS=48.564 M=1 R=2.8 SA=75000.9
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 A_361_50# N_A2_M1000_g A_272_50# VNB NSHORT L=0.15 W=0.42 AD=0.06405
+ AS=0.06195 PD=0.725 PS=0.715 NRD=27.852 NRS=26.424 M=1 R=2.8 SA=75001.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_86_241#_M1009_d N_A1_M1009_g A_361_50# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.06405 PD=0.81 PS=0.725 NRD=11.424 NRS=27.852 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_A_86_241#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_86_241#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1001 N_A_266_483#_M1001_d N_A3_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_266_483#_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1003 N_A_266_483#_M1003_d N_A1_M1003_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_86_241#_M1007_d N_B1_M1007_g N_A_266_483#_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a31o_0.pxi.spice"
*
.ends
*
*
