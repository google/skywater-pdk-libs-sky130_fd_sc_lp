* File: sky130_fd_sc_lp__dfrbp_lp.pex.spice
* Created: Wed Sep  2 09:43:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%D 3 5 6 10 13 17 19 20 21 22 23 34
c64 34 0 4.84792e-20 $X=2.15 $Y=1.295
r65 23 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.295 $X2=2.15 $Y2=1.295
r66 22 23 5.90065 $w=7.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.94 $Y=0.925
+ $X2=1.94 $Y2=1.295
r67 21 22 5.90065 $w=7.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.94 $Y=0.555
+ $X2=1.94 $Y2=0.925
r68 19 34 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.15 $Y=1.24
+ $X2=2.15 $Y2=1.295
r69 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.24
+ $X2=2.15 $Y2=1.075
r70 17 34 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.15 $Y=1.47
+ $X2=2.15 $Y2=1.295
r71 14 17 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.805 $Y=1.545
+ $X2=2.15 $Y2=1.545
r72 13 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.06 $Y=0.79 $X2=2.06
+ $Y2=1.075
r73 8 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.805 $Y=3.075
+ $X2=1.805 $Y2=2.68
r74 7 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=1.62
+ $X2=1.805 $Y2=1.545
r75 7 10 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.805 $Y=1.62
+ $X2=1.805 $Y2=2.68
r76 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.73 $Y=3.15
+ $X2=1.805 $Y2=3.075
r77 5 6 602.5 $w=1.5e-07 $l=1.175e-06 $layer=POLY_cond $X=1.73 $Y=3.15 $X2=0.555
+ $Y2=3.15
r78 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.48 $Y=3.075
+ $X2=0.555 $Y2=3.15
r79 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.48 $Y=3.075 $X2=0.48
+ $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_662_90# 1 2 7 9 12 14 16 18 20 22 25 26
+ 28 29 31 32 33 35 36 37 40 44 46 50 53
c166 37 0 1.05935e-19 $X=6.73 $Y=1.26
c167 20 0 7.06823e-20 $X=9.38 $Y=0.985
c168 16 0 3.0878e-19 $X=8.92 $Y=2.105
c169 14 0 5.56669e-20 $X=8.92 $Y=1.345
r170 51 60 22.7066 $w=4.67e-07 $l=2.2e-07 $layer=POLY_cond $X=8.702 $Y=0.84
+ $X2=8.702 $Y2=1.06
r171 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.575
+ $Y=0.84 $X2=8.575 $Y2=0.84
r172 48 50 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.575 $Y=1.175
+ $X2=8.575 $Y2=0.84
r173 47 53 4.96294 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.145 $Y=1.26
+ $X2=7.98 $Y2=1.26
r174 46 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.41 $Y=1.26
+ $X2=8.575 $Y2=1.175
r175 46 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.41 $Y=1.26
+ $X2=8.145 $Y2=1.26
r176 42 53 1.49777 $w=2.75e-07 $l=9.80051e-08 $layer=LI1_cond $X=7.952 $Y=1.345
+ $X2=7.98 $Y2=1.26
r177 42 44 14.877 $w=2.73e-07 $l=3.55e-07 $layer=LI1_cond $X=7.952 $Y=1.345
+ $X2=7.952 $Y2=1.7
r178 38 53 1.49777 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=1.175
+ $X2=7.98 $Y2=1.26
r179 38 40 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.98 $Y=1.175
+ $X2=7.98 $Y2=0.765
r180 36 53 4.96294 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=1.26
+ $X2=7.98 $Y2=1.26
r181 36 37 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=7.815 $Y=1.26
+ $X2=6.73 $Y2=1.26
r182 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.645 $Y=1.175
+ $X2=6.73 $Y2=1.26
r183 34 35 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.645 $Y=0.435
+ $X2=6.645 $Y2=1.175
r184 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.56 $Y=0.35
+ $X2=6.645 $Y2=0.435
r185 32 33 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=6.56 $Y=0.35
+ $X2=5.395 $Y2=0.35
r186 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.31 $Y=0.435
+ $X2=5.395 $Y2=0.35
r187 30 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.31 $Y=0.435
+ $X2=5.31 $Y2=0.75
r188 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.225 $Y=0.835
+ $X2=5.31 $Y2=0.75
r189 28 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.225 $Y=0.835
+ $X2=3.845 $Y2=0.835
r190 26 56 31.0579 $w=3.85e-07 $l=2.15e-07 $layer=POLY_cond $X=3.68 $Y=1.267
+ $X2=3.465 $Y2=1.267
r191 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.295 $X2=3.68 $Y2=1.295
r192 23 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.68 $Y=0.92
+ $X2=3.845 $Y2=0.835
r193 23 25 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=3.68 $Y=0.92
+ $X2=3.68 $Y2=1.295
r194 20 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.38 $Y=0.985
+ $X2=9.38 $Y2=0.555
r195 19 60 29.6916 $w=1.5e-07 $l=2.93e-07 $layer=POLY_cond $X=8.995 $Y=1.06
+ $X2=8.702 $Y2=1.06
r196 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.305 $Y=1.06
+ $X2=9.38 $Y2=0.985
r197 18 19 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=9.305 $Y=1.06
+ $X2=8.995 $Y2=1.06
r198 14 60 53.4773 $w=4.67e-07 $l=3.78622e-07 $layer=POLY_cond $X=8.92 $Y=1.345
+ $X2=8.702 $Y2=1.06
r199 14 16 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.92 $Y=1.345
+ $X2=8.92 $Y2=2.105
r200 10 56 24.9301 $w=1.5e-07 $l=1.93e-07 $layer=POLY_cond $X=3.465 $Y=1.46
+ $X2=3.465 $Y2=1.267
r201 10 12 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.465 $Y=1.46
+ $X2=3.465 $Y2=2.265
r202 7 56 11.5564 $w=3.85e-07 $l=8e-08 $layer=POLY_cond $X=3.385 $Y=1.267
+ $X2=3.465 $Y2=1.267
r203 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.385 $Y=1.075
+ $X2=3.385 $Y2=0.79
r204 2 44 600 $w=1.7e-07 $l=4.71858e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.065 $X2=8.005 $Y2=1.7
r205 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.84
+ $Y=0.555 $X2=7.98 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_817_90# 1 2 3 4 15 17 19 24 29 30 32 33
+ 36 40 43 44 45 48 51 52 54 57 58
r164 52 54 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.25 $Y=2.04
+ $X2=9.67 $Y2=2.04
r165 51 52 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.165 $Y=1.875
+ $X2=9.25 $Y2=2.04
r166 50 58 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=9.165 $Y=1.695
+ $X2=9.085 $Y2=1.61
r167 50 51 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=9.165 $Y=1.695
+ $X2=9.165 $Y2=1.875
r168 46 58 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.085 $Y=1.525
+ $X2=9.085 $Y2=1.61
r169 46 48 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=9.085 $Y=1.525
+ $X2=9.085 $Y2=0.58
r170 44 58 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.92 $Y=1.61
+ $X2=9.085 $Y2=1.61
r171 44 45 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.92 $Y=1.61
+ $X2=8.44 $Y2=1.61
r172 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.355 $Y=1.695
+ $X2=8.44 $Y2=1.61
r173 42 43 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.355 $Y=1.695
+ $X2=8.355 $Y2=2.045
r174 41 57 5.27292 $w=1.7e-07 $l=1.85257e-07 $layer=LI1_cond $X=6.38 $Y=2.13
+ $X2=6.215 $Y2=2.087
r175 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.27 $Y=2.13
+ $X2=8.355 $Y2=2.045
r176 40 41 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=8.27 $Y=2.13
+ $X2=6.38 $Y2=2.13
r177 34 57 1.30193 $w=3.3e-07 $l=1.27e-07 $layer=LI1_cond $X=6.215 $Y=1.96
+ $X2=6.215 $Y2=2.087
r178 34 36 41.7324 $w=3.28e-07 $l=1.195e-06 $layer=LI1_cond $X=6.215 $Y=1.96
+ $X2=6.215 $Y2=0.765
r179 32 57 5.27292 $w=1.7e-07 $l=1.84811e-07 $layer=LI1_cond $X=6.05 $Y=2.045
+ $X2=6.215 $Y2=2.087
r180 32 33 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=6.05 $Y=2.045
+ $X2=4.705 $Y2=2.045
r181 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.54
+ $Y=1.62 $X2=4.54 $Y2=1.62
r182 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.705 $Y2=2.045
r183 27 29 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.54 $Y2=1.62
r184 26 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.54 $Y=1.96
+ $X2=4.54 $Y2=1.62
r185 24 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.54 $Y=1.605
+ $X2=4.54 $Y2=1.62
r186 21 24 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.16 $Y=1.53
+ $X2=4.54 $Y2=1.53
r187 17 26 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=2.125
+ $X2=4.54 $Y2=1.96
r188 17 19 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.54 $Y=2.125
+ $X2=4.54 $Y2=2.495
r189 13 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.16 $Y=1.455
+ $X2=4.16 $Y2=1.53
r190 13 15 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=4.16 $Y=1.455
+ $X2=4.16 $Y2=0.79
r191 4 54 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.53
+ $Y=1.895 $X2=9.67 $Y2=2.04
r192 3 57 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=6.085
+ $Y=1.865 $X2=6.215 $Y2=2.01
r193 2 48 182 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_NDIFF $count=1 $X=8.94
+ $Y=0.235 $X2=9.085 $Y2=0.58
r194 1 36 182 $w=1.7e-07 $l=4.97242e-07 $layer=licon1_NDIFF $count=1 $X=6.07
+ $Y=0.335 $X2=6.215 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%RESET_B 1 3 7 9 10 14 15 16 20 21 22 25 27
+ 28 30 33 35 39 43 49 51 53 55 56 57 58 65 66 69 70 72 75 76
c249 76 0 1.0799e-19 $X=12.29 $Y=1.275
c250 70 0 1.56469e-19 $X=1.15 $Y=1.275
c251 53 0 1.68525e-19 $X=12.36 $Y=1.63
c252 43 0 5.70993e-20 $X=12.54 $Y=2.195
c253 35 0 6.56506e-20 $X=12.18 $Y=2.195
r254 76 88 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=12.29 $Y=1.275
+ $X2=12.29 $Y2=1.665
r255 75 77 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=12.285 $Y=1.275
+ $X2=12.285 $Y2=1.11
r256 75 76 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.29
+ $Y=1.275 $X2=12.29 $Y2=1.275
r257 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.275 $X2=1.15 $Y2=1.275
r258 66 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=1.665
+ $X2=12.24 $Y2=1.665
r259 65 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.11
+ $Y=1.615 $X2=5.11 $Y2=1.615
r260 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r261 61 70 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.275
r262 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r263 58 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r264 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=12.24 $Y2=1.665
r265 57 58 8.55196 $w=1.4e-07 $l=6.91e-06 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=5.185 $Y2=1.665
r266 56 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r267 55 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=5.04 $Y2=1.665
r268 55 56 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=1.345 $Y2=1.665
r269 51 72 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=5.11 $Y=1.845
+ $X2=5.11 $Y2=1.615
r270 49 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.11 $Y=1.45
+ $X2=5.11 $Y2=1.615
r271 46 69 26.2269 $w=5.1e-07 $l=2.5e-07 $layer=POLY_cond $X=1.09 $Y=1.525
+ $X2=1.09 $Y2=1.275
r272 45 69 1.57362 $w=5.1e-07 $l=1.5e-08 $layer=POLY_cond $X=1.09 $Y=1.26
+ $X2=1.09 $Y2=1.275
r273 39 77 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=12.39 $Y=0.465
+ $X2=12.39 $Y2=1.11
r274 33 53 25.8164 $w=3.6e-07 $l=1.5e-07 $layer=POLY_cond $X=12.36 $Y=1.78
+ $X2=12.36 $Y2=1.63
r275 33 43 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=12.54 $Y=1.78
+ $X2=12.54 $Y2=2.195
r276 33 35 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=12.18 $Y=1.78
+ $X2=12.18 $Y2=2.195
r277 31 75 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=12.285 $Y=1.29
+ $X2=12.285 $Y2=1.275
r278 31 53 54.4984 $w=3.6e-07 $l=3.4e-07 $layer=POLY_cond $X=12.285 $Y=1.29
+ $X2=12.285 $Y2=1.63
r279 28 51 79.5963 $w=2.18e-07 $l=4.31833e-07 $layer=POLY_cond $X=5.47 $Y=2.16
+ $X2=5.11 $Y2=2.002
r280 28 30 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.47 $Y=2.16
+ $X2=5.47 $Y2=2.495
r281 25 51 11.5617 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=5.11 $Y=2.16
+ $X2=5.11 $Y2=2.002
r282 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.11 $Y=2.16
+ $X2=5.11 $Y2=2.495
r283 23 49 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=5.02 $Y=1.225
+ $X2=5.02 $Y2=1.45
r284 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.945 $Y=1.15
+ $X2=5.02 $Y2=1.225
r285 21 22 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.945 $Y=1.15
+ $X2=4.625 $Y2=1.15
r286 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.55 $Y=1.075
+ $X2=4.625 $Y2=1.15
r287 18 20 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.55 $Y=1.075
+ $X2=4.55 $Y2=0.79
r288 17 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.55 $Y=0.24
+ $X2=4.55 $Y2=0.79
r289 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.475 $Y=0.165
+ $X2=4.55 $Y2=0.24
r290 15 16 1399.85 $w=1.5e-07 $l=2.73e-06 $layer=POLY_cond $X=4.475 $Y=0.165
+ $X2=1.745 $Y2=0.165
r291 12 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.67 $Y=1.11
+ $X2=1.67 $Y2=0.79
r292 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.67 $Y=0.24
+ $X2=1.745 $Y2=0.165
r293 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.67 $Y=0.24
+ $X2=1.67 $Y2=0.79
r294 10 45 38.9973 $w=1.5e-07 $l=2.90086e-07 $layer=POLY_cond $X=1.345 $Y=1.185
+ $X2=1.09 $Y2=1.26
r295 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.595 $Y=1.185
+ $X2=1.67 $Y2=1.11
r296 9 10 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.595 $Y=1.185
+ $X2=1.345 $Y2=1.185
r297 1 46 35.748 $w=5.1e-07 $l=2.55e-07 $layer=POLY_cond $X=1.09 $Y=1.78
+ $X2=1.09 $Y2=1.525
r298 1 7 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.27 $Y=1.78
+ $X2=1.27 $Y2=2.495
r299 1 3 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=0.91 $Y=1.78
+ $X2=0.91 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_590_116# 1 2 3 10 11 12 14 17 19 21 23 26
+ 29 30 32 35 37 40 42 43 44 45 46 50 53 54 55 61 62
c177 30 0 1.05935e-19 $X=6.79 $Y=1.175
r178 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.705
+ $Y=1.265 $X2=5.705 $Y2=1.265
r179 55 58 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.685 $Y=2.395
+ $X2=5.685 $Y2=2.515
r180 50 52 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.17 $Y=0.79
+ $X2=3.17 $Y2=1
r181 45 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=2.395
+ $X2=5.685 $Y2=2.395
r182 45 46 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=5.52 $Y=2.395
+ $X2=4.195 $Y2=2.395
r183 43 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=1.185
+ $X2=5.705 $Y2=1.185
r184 43 44 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.54 $Y=1.185
+ $X2=4.195 $Y2=1.185
r185 42 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.11 $Y=2.31
+ $X2=4.195 $Y2=2.395
r186 41 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=1.855
+ $X2=4.11 $Y2=1.77
r187 41 42 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=4.11 $Y=1.855
+ $X2=4.11 $Y2=2.31
r188 40 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=1.685
+ $X2=4.11 $Y2=1.77
r189 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.11 $Y=1.27
+ $X2=4.195 $Y2=1.185
r190 39 40 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.11 $Y=1.27
+ $X2=4.11 $Y2=1.685
r191 38 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.77
+ $X2=3.25 $Y2=1.77
r192 37 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=1.77
+ $X2=4.11 $Y2=1.77
r193 37 38 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.025 $Y=1.77
+ $X2=3.335 $Y2=1.77
r194 33 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=1.855
+ $X2=3.25 $Y2=1.77
r195 33 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.25 $Y=1.855
+ $X2=3.25 $Y2=2.2
r196 32 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=1.685
+ $X2=3.25 $Y2=1.77
r197 32 52 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.25 $Y=1.685
+ $X2=3.25 $Y2=1
r198 28 62 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.705 $Y=1.25
+ $X2=5.705 $Y2=1.265
r199 24 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.79 $Y=1.25
+ $X2=6.79 $Y2=1.175
r200 24 26 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=6.79 $Y=1.25
+ $X2=6.79 $Y2=2.285
r201 21 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.79 $Y=1.1
+ $X2=6.79 $Y2=1.175
r202 21 23 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.79 $Y=1.1
+ $X2=6.79 $Y2=0.655
r203 20 29 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.505 $Y=1.175
+ $X2=6.43 $Y2=1.175
r204 19 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.715 $Y=1.175
+ $X2=6.79 $Y2=1.175
r205 19 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.715 $Y=1.175
+ $X2=6.505 $Y2=1.175
r206 15 29 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.43 $Y=1.25 $X2=6.43
+ $Y2=1.175
r207 15 17 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=6.43 $Y=1.25
+ $X2=6.43 $Y2=2.285
r208 12 29 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.43 $Y=1.1 $X2=6.43
+ $Y2=1.175
r209 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.43 $Y=1.1
+ $X2=6.43 $Y2=0.655
r210 11 28 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.87 $Y=1.175
+ $X2=5.705 $Y2=1.25
r211 10 29 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.355 $Y=1.175
+ $X2=6.43 $Y2=1.175
r212 10 11 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.355 $Y=1.175
+ $X2=5.87 $Y2=1.175
r213 3 58 600 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=1 $X=5.545
+ $Y=2.285 $X2=5.685 $Y2=2.515
r214 2 35 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.055 $X2=3.25 $Y2=2.2
r215 1 50 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=2.95
+ $Y=0.58 $X2=3.17 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_560_90# 1 2 9 14 15 16 20 23 25 30 33 35
+ 40 41 42 45 49 55 57 60 63 64 66 67 69 70 71 75 76 79 80 81 82 84
c242 67 0 7.06823e-20 $X=10.27 $Y=0.75
r243 83 84 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=15.25 $Y=0.9
+ $X2=15.25 $Y2=1.94
r244 81 84 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.165 $Y=2.025
+ $X2=15.25 $Y2=1.94
r245 81 82 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=15.165 $Y=2.025
+ $X2=14.03 $Y2=2.025
r246 79 83 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.165 $Y=0.815
+ $X2=15.25 $Y2=0.9
r247 79 80 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=15.165 $Y=0.815
+ $X2=14 $Y2=0.815
r248 76 82 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.865 $Y=2.11
+ $X2=14.03 $Y2=2.025
r249 76 78 3.88182 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=13.865 $Y=2.11
+ $X2=13.865 $Y2=2.215
r250 73 80 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.835 $Y=0.73
+ $X2=14 $Y2=0.815
r251 73 75 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=13.835 $Y=0.73
+ $X2=13.835 $Y2=0.47
r252 72 75 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=13.835 $Y=0.435
+ $X2=13.835 $Y2=0.47
r253 70 72 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.67 $Y=0.35
+ $X2=13.835 $Y2=0.435
r254 70 71 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=13.67 $Y=0.35
+ $X2=11.315 $Y2=0.35
r255 68 71 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.23 $Y=0.435
+ $X2=11.315 $Y2=0.35
r256 68 69 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.23 $Y=0.435
+ $X2=11.23 $Y2=0.665
r257 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.145 $Y=0.75
+ $X2=11.23 $Y2=0.665
r258 66 67 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=11.145 $Y=0.75
+ $X2=10.27 $Y2=0.75
r259 64 87 35.7527 $w=4.2e-07 $l=2.7e-07 $layer=POLY_cond $X=10.06 $Y=1.18
+ $X2=10.06 $Y2=1.45
r260 64 86 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.06 $Y=1.18
+ $X2=10.06 $Y2=1.015
r261 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.105
+ $Y=1.18 $X2=10.105 $Y2=1.18
r262 61 67 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.105 $Y=0.835
+ $X2=10.27 $Y2=0.75
r263 61 63 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=10.105 $Y=0.835
+ $X2=10.105 $Y2=1.18
r264 57 58 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.325 $Y=2.92
+ $X2=7.325 $Y2=3.15
r265 54 55 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.685 $Y=1.405
+ $X2=7.765 $Y2=1.405
r266 53 54 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.405 $Y=1.405
+ $X2=7.685 $Y2=1.405
r267 51 53 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.325 $Y=1.405
+ $X2=7.405 $Y2=1.405
r268 47 49 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.875 $Y=1.87
+ $X2=3.035 $Y2=1.87
r269 45 86 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=9.925 $Y=0.465
+ $X2=9.925 $Y2=1.015
r270 41 87 27.059 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.85 $Y=1.45
+ $X2=10.06 $Y2=1.45
r271 41 42 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.85 $Y=1.45
+ $X2=9.53 $Y2=1.45
r272 38 40 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.455 $Y=2.845
+ $X2=9.455 $Y2=2.315
r273 37 42 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.455 $Y=1.525
+ $X2=9.53 $Y2=1.45
r274 37 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.455 $Y=1.525
+ $X2=9.455 $Y2=2.315
r275 36 60 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.76 $Y=2.92
+ $X2=7.685 $Y2=2.92
r276 35 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.38 $Y=2.92
+ $X2=9.455 $Y2=2.845
r277 35 36 830.681 $w=1.5e-07 $l=1.62e-06 $layer=POLY_cond $X=9.38 $Y=2.92
+ $X2=7.76 $Y2=2.92
r278 31 55 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.765 $Y=1.33
+ $X2=7.765 $Y2=1.405
r279 31 33 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=7.765 $Y=1.33
+ $X2=7.765 $Y2=0.765
r280 28 60 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.685 $Y=2.845
+ $X2=7.685 $Y2=2.92
r281 28 30 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.685 $Y=2.845
+ $X2=7.685 $Y2=2.385
r282 27 54 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.685 $Y=1.48
+ $X2=7.685 $Y2=1.405
r283 27 30 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=7.685 $Y=1.48
+ $X2=7.685 $Y2=2.385
r284 26 57 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.4 $Y=2.92
+ $X2=7.325 $Y2=2.92
r285 25 60 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.61 $Y=2.92
+ $X2=7.685 $Y2=2.92
r286 25 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.61 $Y=2.92
+ $X2=7.4 $Y2=2.92
r287 21 53 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.405 $Y=1.33
+ $X2=7.405 $Y2=1.405
r288 21 23 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=7.405 $Y=1.33
+ $X2=7.405 $Y2=0.765
r289 18 57 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.325 $Y=2.845
+ $X2=7.325 $Y2=2.92
r290 18 20 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.325 $Y=2.845
+ $X2=7.325 $Y2=2.385
r291 17 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.325 $Y=1.48
+ $X2=7.325 $Y2=1.405
r292 17 20 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=7.325 $Y=1.48
+ $X2=7.325 $Y2=2.385
r293 15 58 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.25 $Y=3.15
+ $X2=7.325 $Y2=3.15
r294 15 16 2122.85 $w=1.5e-07 $l=4.14e-06 $layer=POLY_cond $X=7.25 $Y=3.15
+ $X2=3.11 $Y2=3.15
r295 12 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.035 $Y=3.075
+ $X2=3.11 $Y2=3.15
r296 12 14 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.035 $Y=3.075
+ $X2=3.035 $Y2=2.265
r297 11 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.035 $Y=1.945
+ $X2=3.035 $Y2=1.87
r298 11 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.035 $Y=1.945
+ $X2=3.035 $Y2=2.265
r299 7 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=1.795
+ $X2=2.875 $Y2=1.87
r300 7 9 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=2.875 $Y=1.795
+ $X2=2.875 $Y2=0.79
r301 2 78 600 $w=1.7e-07 $l=4.4238e-07 $layer=licon1_PDIFF $count=1 $X=13.73
+ $Y=1.835 $X2=13.865 $Y2=2.215
r302 1 75 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=13.69
+ $Y=0.24 $X2=13.835 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_2102_25# 1 2 9 13 15 18 21 23 25 27 31 33
r76 31 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.675 $Y=1.18
+ $X2=10.675 $Y2=1.345
r77 31 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.675 $Y=1.18
+ $X2=10.675 $Y2=1.015
r78 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.675
+ $Y=1.18 $X2=10.675 $Y2=1.18
r79 27 30 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.675 $Y=1.1
+ $X2=10.675 $Y2=1.18
r80 23 25 54.1648 $w=2.48e-07 $l=1.175e-06 $layer=LI1_cond $X=11.935 $Y=0.74
+ $X2=13.11 $Y2=0.74
r81 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.85 $Y=1.185
+ $X2=11.85 $Y2=1.1
r82 19 21 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=11.85 $Y=1.185
+ $X2=11.85 $Y2=2.165
r83 18 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.85 $Y=1.015
+ $X2=11.85 $Y2=1.1
r84 17 23 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.85 $Y=0.865
+ $X2=11.935 $Y2=0.74
r85 17 18 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=11.85 $Y=0.865
+ $X2=11.85 $Y2=1.015
r86 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.84 $Y=1.1
+ $X2=10.675 $Y2=1.1
r87 15 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.765 $Y=1.1
+ $X2=11.85 $Y2=1.1
r88 15 16 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=11.765 $Y=1.1
+ $X2=10.84 $Y2=1.1
r89 13 36 789.66 $w=1.5e-07 $l=1.54e-06 $layer=POLY_cond $X=10.585 $Y=2.885
+ $X2=10.585 $Y2=1.345
r90 9 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.585 $Y=0.465
+ $X2=10.585 $Y2=1.015
r91 2 21 600 $w=1.7e-07 $l=3.33054e-07 $layer=licon1_PDIFF $count=1 $X=11.595
+ $Y=1.985 $X2=11.85 $Y2=2.165
r92 1 25 182 $w=1.7e-07 $l=5.58122e-07 $layer=licon1_NDIFF $count=1 $X=12.855
+ $Y=0.255 $X2=13.11 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_1799_379# 1 2 9 13 15 16 21 25 29 31 35
+ 39 41 45 49 51 55 59 61 62 63 64 70 72 73 75 79 80 81 83 84 85 86 87 88 90 94
+ 95 99 101 108 111 116
c249 88 0 1.39319e-19 $X=14.725 $Y=1.675
c250 86 0 1.68525e-19 $X=13.205 $Y=1.76
c251 73 0 1.81705e-19 $X=9.76 $Y=1.61
c252 70 0 1.27075e-19 $X=9.595 $Y=0.58
c253 35 0 1.69072e-19 $X=15.465 $Y=0.66
r254 115 116 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=15.105 $Y=1.51
+ $X2=15.18 $Y2=1.51
r255 102 115 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=14.89 $Y=1.51
+ $X2=15.105 $Y2=1.51
r256 101 104 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=14.855 $Y=1.51
+ $X2=14.855 $Y2=1.675
r257 101 102 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.89
+ $Y=1.51 $X2=14.89 $Y2=1.51
r258 99 112 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.205 $Y=1.755
+ $X2=13.205 $Y2=1.92
r259 99 111 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.205 $Y=1.755
+ $X2=13.205 $Y2=1.59
r260 98 99 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.205
+ $Y=1.755 $X2=13.205 $Y2=1.755
r261 93 108 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=11.38 $Y=1.53
+ $X2=11.52 $Y2=1.53
r262 92 95 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=11.38 $Y=1.53
+ $X2=11.5 $Y2=1.53
r263 92 94 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.38 $Y=1.53
+ $X2=11.215 $Y2=1.53
r264 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.38
+ $Y=1.53 $X2=11.38 $Y2=1.53
r265 89 98 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.37 $Y=1.675
+ $X2=13.205 $Y2=1.675
r266 88 104 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=14.725 $Y=1.675
+ $X2=14.855 $Y2=1.675
r267 88 89 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=14.725 $Y=1.675
+ $X2=13.37 $Y2=1.675
r268 86 98 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=1.76
+ $X2=13.205 $Y2=1.675
r269 86 87 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=13.205 $Y=1.76
+ $X2=13.205 $Y2=1.96
r270 84 87 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.04 $Y=2.045
+ $X2=13.205 $Y2=1.96
r271 84 85 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=13.04 $Y=2.045
+ $X2=12.285 $Y2=2.045
r272 82 85 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.2 $Y=2.13
+ $X2=12.285 $Y2=2.045
r273 82 83 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=12.2 $Y=2.13
+ $X2=12.2 $Y2=2.545
r274 80 83 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.115 $Y=2.63
+ $X2=12.2 $Y2=2.545
r275 80 81 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=12.115 $Y=2.63
+ $X2=11.585 $Y2=2.63
r276 79 81 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.5 $Y=2.545
+ $X2=11.585 $Y2=2.63
r277 78 95 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.5 $Y=1.695
+ $X2=11.5 $Y2=1.53
r278 78 79 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=11.5 $Y=1.695
+ $X2=11.5 $Y2=2.545
r279 77 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.105 $Y=1.61
+ $X2=10.02 $Y2=1.61
r280 77 94 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=10.105 $Y=1.61
+ $X2=11.215 $Y2=1.61
r281 74 90 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.02 $Y=1.695
+ $X2=10.02 $Y2=1.61
r282 74 75 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.02 $Y=1.695
+ $X2=10.02 $Y2=2.385
r283 72 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.935 $Y=1.61
+ $X2=10.02 $Y2=1.61
r284 72 73 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.935 $Y=1.61
+ $X2=9.76 $Y2=1.61
r285 68 73 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.595 $Y=1.525
+ $X2=9.76 $Y2=1.61
r286 68 70 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=9.595 $Y=1.525
+ $X2=9.595 $Y2=0.58
r287 64 75 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.935 $Y=2.55
+ $X2=10.02 $Y2=2.385
r288 64 66 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.935 $Y=2.55
+ $X2=9.24 $Y2=2.55
r289 57 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.83 $Y=1.495
+ $X2=16.83 $Y2=1.42
r290 57 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=16.83 $Y=1.495
+ $X2=16.83 $Y2=2.155
r291 53 63 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.83 $Y=1.345
+ $X2=16.83 $Y2=1.42
r292 53 55 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=16.83 $Y=1.345
+ $X2=16.83 $Y2=0.895
r293 52 62 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.545 $Y=1.42
+ $X2=16.47 $Y2=1.42
r294 51 63 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.755 $Y=1.42
+ $X2=16.83 $Y2=1.42
r295 51 52 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=16.755 $Y=1.42
+ $X2=16.545 $Y2=1.42
r296 47 62 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.47 $Y=1.495
+ $X2=16.47 $Y2=1.42
r297 47 49 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=16.47 $Y=1.495
+ $X2=16.47 $Y2=2.155
r298 43 62 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.47 $Y=1.345
+ $X2=16.47 $Y2=1.42
r299 43 45 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=16.47 $Y=1.345
+ $X2=16.47 $Y2=0.895
r300 42 61 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.54 $Y=1.42
+ $X2=15.465 $Y2=1.42
r301 41 62 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.395 $Y=1.42
+ $X2=16.47 $Y2=1.42
r302 41 42 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=16.395 $Y=1.42
+ $X2=15.54 $Y2=1.42
r303 37 61 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.465 $Y=1.495
+ $X2=15.465 $Y2=1.42
r304 37 39 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=15.465 $Y=1.495
+ $X2=15.465 $Y2=2.465
r305 33 61 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.465 $Y=1.345
+ $X2=15.465 $Y2=1.42
r306 33 35 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=15.465 $Y=1.345
+ $X2=15.465 $Y2=0.66
r307 31 61 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.39 $Y=1.42
+ $X2=15.465 $Y2=1.42
r308 31 116 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=15.39 $Y=1.42
+ $X2=15.18 $Y2=1.42
r309 27 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.105 $Y=1.675
+ $X2=15.105 $Y2=1.51
r310 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=15.105 $Y=1.675
+ $X2=15.105 $Y2=2.465
r311 23 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.105 $Y=1.345
+ $X2=15.105 $Y2=1.51
r312 23 25 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=15.105 $Y=1.345
+ $X2=15.105 $Y2=0.66
r313 21 112 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=13.115 $Y=2.76
+ $X2=13.115 $Y2=1.92
r314 17 111 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=13.115 $Y=1.07
+ $X2=13.115 $Y2=1.59
r315 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.04 $Y=0.995
+ $X2=13.115 $Y2=1.07
r316 15 16 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=13.04 $Y=0.995
+ $X2=12.855 $Y2=0.995
r317 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.78 $Y=0.92
+ $X2=12.855 $Y2=0.995
r318 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=12.78 $Y=0.92
+ $X2=12.78 $Y2=0.465
r319 7 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.52 $Y=1.695
+ $X2=11.52 $Y2=1.53
r320 7 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=11.52 $Y=1.695
+ $X2=11.52 $Y2=2.195
r321 2 66 600 $w=1.7e-07 $l=7.67789e-07 $layer=licon1_PDIFF $count=1 $X=8.995
+ $Y=1.895 $X2=9.24 $Y2=2.55
r322 1 70 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=9.455
+ $Y=0.235 $X2=9.595 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%CLK 3 7 9 13 17 19 20 21 24
c57 9 0 1.39319e-19 $X=14.365 $Y=1.155
r58 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.99 $Y=1.245
+ $X2=13.99 $Y2=1.41
r59 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.99
+ $Y=1.245 $X2=13.99 $Y2=1.245
r60 24 27 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.99 $Y=1.155
+ $X2=13.99 $Y2=1.245
r61 24 25 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=13.99 $Y=1.155
+ $X2=13.99 $Y2=1.08
r62 21 28 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=14.16 $Y=1.245
+ $X2=13.99 $Y2=1.245
r63 20 28 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=13.68 $Y=1.245
+ $X2=13.99 $Y2=1.245
r64 15 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.44 $Y=1.23
+ $X2=14.44 $Y2=1.155
r65 15 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=14.44 $Y=1.23
+ $X2=14.44 $Y2=2.155
r66 11 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.44 $Y=1.08
+ $X2=14.44 $Y2=1.155
r67 11 13 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=14.44 $Y=1.08
+ $X2=14.44 $Y2=0.45
r68 10 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.155 $Y=1.155
+ $X2=13.99 $Y2=1.155
r69 9 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.365 $Y=1.155
+ $X2=14.44 $Y2=1.155
r70 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=14.365 $Y=1.155
+ $X2=14.155 $Y2=1.155
r71 7 29 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=14.08 $Y=2.155
+ $X2=14.08 $Y2=1.41
r72 3 25 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=14.05 $Y=0.45
+ $X2=14.05 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_3222_137# 1 2 9 13 17 21 25 29 33 36 40
c62 36 0 1.69072e-19 $X=16.255 $Y=1.47
c63 29 0 1.59406e-19 $X=16.255 $Y=1.98
r64 34 40 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=17.44 $Y=1.47
+ $X2=17.735 $Y2=1.47
r65 34 37 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=17.44 $Y=1.47
+ $X2=17.375 $Y2=1.47
r66 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.44
+ $Y=1.47 $X2=17.44 $Y2=1.47
r67 31 36 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.42 $Y=1.47
+ $X2=16.255 $Y2=1.47
r68 31 33 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=16.42 $Y=1.47
+ $X2=17.44 $Y2=1.47
r69 27 36 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.255 $Y=1.635
+ $X2=16.255 $Y2=1.47
r70 27 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=16.255 $Y=1.635
+ $X2=16.255 $Y2=1.98
r71 23 36 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.255 $Y=1.305
+ $X2=16.255 $Y2=1.47
r72 23 25 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=16.255 $Y=1.305
+ $X2=16.255 $Y2=0.895
r73 19 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.735 $Y=1.635
+ $X2=17.735 $Y2=1.47
r74 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=17.735 $Y=1.635
+ $X2=17.735 $Y2=2.465
r75 15 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.735 $Y=1.305
+ $X2=17.735 $Y2=1.47
r76 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=17.735 $Y=1.305
+ $X2=17.735 $Y2=0.685
r77 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.375 $Y=1.635
+ $X2=17.375 $Y2=1.47
r78 11 13 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=17.375 $Y=1.635
+ $X2=17.375 $Y2=2.465
r79 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.375 $Y=1.305
+ $X2=17.375 $Y2=1.47
r80 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=17.375 $Y=1.305
+ $X2=17.375 $Y2=0.685
r81 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.11
+ $Y=1.835 $X2=16.255 $Y2=1.98
r82 1 25 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=16.11
+ $Y=0.685 $X2=16.255 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_27_457# 1 2 9 11 12 14 15 16 19
r41 17 19 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=2.06 $Y=2.48 $X2=2.06
+ $Y2=2.68
r42 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.935 $Y=2.395
+ $X2=2.06 $Y2=2.48
r43 15 16 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.935 $Y=2.395
+ $X2=1.21 $Y2=2.395
r44 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.125 $Y=2.48
+ $X2=1.21 $Y2=2.395
r45 13 14 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.125 $Y=2.48
+ $X2=1.125 $Y2=2.895
r46 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.04 $Y=2.98
+ $X2=1.125 $Y2=2.895
r47 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.04 $Y=2.98 $X2=0.35
+ $Y2=2.98
r48 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.225 $Y=2.895
+ $X2=0.35 $Y2=2.98
r49 7 9 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.225 $Y=2.895 $X2=0.225
+ $Y2=2.495
r50 2 19 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=2.47 $X2=2.02 $Y2=2.68
r51 1 9 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.285 $X2=0.265 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_111_457# 1 2 3 12 14 15 18 21 22 23 26 28
r74 24 26 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.68 $Y=2.545
+ $X2=3.68 $Y2=2.265
r75 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.515 $Y=2.63
+ $X2=3.68 $Y2=2.545
r76 22 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.515 $Y=2.63
+ $X2=2.985 $Y2=2.63
r77 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.9 $Y=2.545
+ $X2=2.985 $Y2=2.63
r78 20 28 3.70735 $w=2.5e-07 $l=1.9799e-07 $layer=LI1_cond $X=2.9 $Y=2.13
+ $X2=2.74 $Y2=2.045
r79 20 21 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.9 $Y=2.13 $X2=2.9
+ $Y2=2.545
r80 16 28 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.66 $Y=1.96
+ $X2=2.74 $Y2=2.045
r81 16 18 40.8593 $w=3.28e-07 $l=1.17e-06 $layer=LI1_cond $X=2.66 $Y=1.96
+ $X2=2.66 $Y2=0.79
r82 14 28 2.76166 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.495 $Y=2.045
+ $X2=2.74 $Y2=2.045
r83 14 15 106.668 $w=1.68e-07 $l=1.635e-06 $layer=LI1_cond $X=2.495 $Y=2.045
+ $X2=0.86 $Y2=2.045
r84 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.695 $Y=2.13
+ $X2=0.86 $Y2=2.045
r85 10 12 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.695 $Y=2.13
+ $X2=0.695 $Y2=2.49
r86 3 26 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=2.055 $X2=3.68 $Y2=2.265
r87 2 12 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=2.285 $X2=0.695 $Y2=2.49
r88 1 18 182 $w=1.7e-07 $l=6.21188e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.58 $X2=2.66 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48 53
+ 54 56 57 59 60 61 63 75 82 103 109 110 113 116 119 122
r153 122 123 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r154 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r155 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r156 113 114 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r157 110 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18 $Y=3.33
+ $X2=17.04 $Y2=3.33
r158 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18 $Y=3.33
+ $X2=18 $Y2=3.33
r159 107 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.325 $Y=3.33
+ $X2=17.16 $Y2=3.33
r160 107 109 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=17.325 $Y=3.33
+ $X2=18 $Y2=3.33
r161 106 123 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=17.04 $Y2=3.33
r162 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r163 103 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.995 $Y=3.33
+ $X2=17.16 $Y2=3.33
r164 103 105 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=16.995 $Y=3.33
+ $X2=15.12 $Y2=3.33
r165 102 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r166 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r167 99 102 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=14.64 $Y2=3.33
r168 98 101 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=13.2 $Y=3.33
+ $X2=14.64 $Y2=3.33
r169 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r170 96 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r171 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r172 93 96 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.72 $Y2=3.33
r173 93 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r174 92 95 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.72 $Y2=3.33
r175 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r176 90 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.885 $Y=3.33
+ $X2=10.76 $Y2=3.33
r177 90 92 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.885 $Y=3.33
+ $X2=11.28 $Y2=3.33
r178 89 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r179 88 89 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r180 86 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r181 85 88 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=10.32 $Y2=3.33
r182 85 86 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r183 83 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=7.005 $Y2=3.33
r184 83 85 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=7.44 $Y2=3.33
r185 82 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.76 $Y2=3.33
r186 82 88 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.32 $Y2=3.33
r187 81 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r188 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r189 78 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r191 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r192 75 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.84 $Y=3.33
+ $X2=7.005 $Y2=3.33
r193 75 80 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.84 $Y=3.33
+ $X2=6.48 $Y2=3.33
r194 74 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r195 74 114 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=1.68 $Y2=3.33
r196 73 74 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r197 71 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.59 $Y2=3.33
r198 71 73 183 $w=1.68e-07 $l=2.805e-06 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=4.56 $Y2=3.33
r199 70 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r200 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r201 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r202 65 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r203 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r204 63 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.59 $Y2=3.33
r205 63 69 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r206 61 89 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=10.32 $Y2=3.33
r207 61 86 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=7.44 $Y2=3.33
r208 59 101 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=14.715 $Y=3.33
+ $X2=14.64 $Y2=3.33
r209 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.715 $Y=3.33
+ $X2=14.88 $Y2=3.33
r210 58 105 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=15.045 $Y=3.33
+ $X2=15.12 $Y2=3.33
r211 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.045 $Y=3.33
+ $X2=14.88 $Y2=3.33
r212 56 95 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=12.815 $Y=3.33
+ $X2=12.72 $Y2=3.33
r213 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.815 $Y=3.33
+ $X2=12.9 $Y2=3.33
r214 55 98 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=12.985 $Y=3.33
+ $X2=13.2 $Y2=3.33
r215 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.985 $Y=3.33
+ $X2=12.9 $Y2=3.33
r216 53 73 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.66 $Y=3.33 $X2=4.56
+ $Y2=3.33
r217 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=4.825 $Y2=3.33
r218 52 77 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.99 $Y=3.33 $X2=5.04
+ $Y2=3.33
r219 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=3.33
+ $X2=4.825 $Y2=3.33
r220 48 51 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=17.16 $Y=1.98
+ $X2=17.16 $Y2=2.465
r221 46 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.16 $Y=3.245
+ $X2=17.16 $Y2=3.33
r222 46 51 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=17.16 $Y=3.245
+ $X2=17.16 $Y2=2.465
r223 42 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.88 $Y=3.245
+ $X2=14.88 $Y2=3.33
r224 42 44 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=14.88 $Y=3.245
+ $X2=14.88 $Y2=2.455
r225 38 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.9 $Y=3.245
+ $X2=12.9 $Y2=3.33
r226 38 40 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=12.9 $Y=3.245
+ $X2=12.9 $Y2=2.825
r227 34 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.76 $Y2=3.33
r228 34 36 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.76 $Y2=2.885
r229 30 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.005 $Y=3.245
+ $X2=7.005 $Y2=3.33
r230 30 32 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=7.005 $Y=3.245
+ $X2=7.005 $Y2=2.56
r231 26 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.825 $Y=3.245
+ $X2=4.825 $Y2=3.33
r232 26 28 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.825 $Y=3.245
+ $X2=4.825 $Y2=2.825
r233 22 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=3.33
r234 22 24 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=2.745
r235 7 51 300 $w=1.7e-07 $l=7.46693e-07 $layer=licon1_PDIFF $count=2 $X=16.905
+ $Y=1.835 $X2=17.16 $Y2=2.465
r236 7 48 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=16.905
+ $Y=1.835 $X2=17.16 $Y2=1.98
r237 6 44 300 $w=1.7e-07 $l=7.81473e-07 $layer=licon1_PDIFF $count=2 $X=14.515
+ $Y=1.835 $X2=14.88 $Y2=2.455
r238 5 40 600 $w=1.7e-07 $l=9.72111e-07 $layer=licon1_PDIFF $count=1 $X=12.615
+ $Y=1.985 $X2=12.9 $Y2=2.825
r239 4 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.66
+ $Y=2.675 $X2=10.8 $Y2=2.885
r240 3 32 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=1.865 $X2=7.005 $Y2=2.56
r241 2 28 600 $w=1.7e-07 $l=6.36396e-07 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=2.285 $X2=4.825 $Y2=2.825
r242 1 24 600 $w=1.7e-07 $l=5.69473e-07 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=2.285 $X2=1.59 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_484_411# 1 2 9 11 12 14
r40 14 16 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.22 $Y=2.825
+ $X2=4.22 $Y2=2.98
r41 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=2.98
+ $X2=4.22 $Y2=2.98
r42 11 12 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=4.055 $Y=2.98
+ $X2=2.635 $Y2=2.98
r43 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.51 $Y=2.895
+ $X2=2.635 $Y2=2.98
r44 7 9 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=2.51 $Y=2.895 $X2=2.51
+ $Y2=2.475
r45 2 14 600 $w=1.7e-07 $l=6.03738e-07 $layer=licon1_PDIFF $count=1 $X=4.085
+ $Y=2.285 $X2=4.22 $Y2=2.825
r46 1 9 600 $w=1.7e-07 $l=4.80625e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=2.055 $X2=2.55 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_1712_379# 1 2 9 11 12 14
r27 14 16 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=10.37 $Y=2.86
+ $X2=10.37 $Y2=2.98
r28 11 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=2.98
+ $X2=10.37 $Y2=2.98
r29 11 12 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=10.285 $Y=2.98
+ $X2=8.87 $Y2=2.98
r30 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.745 $Y=2.895
+ $X2=8.87 $Y2=2.98
r31 7 9 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.745 $Y=2.895
+ $X2=8.745 $Y2=2.105
r32 2 14 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=10.225
+ $Y=2.675 $X2=10.37 $Y2=2.86
r33 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=1.895 $X2=8.705 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%A_2185_397# 1 2 8 9 10 12 13 14 17 20
c51 17 0 5.70993e-20 $X=13.33 $Y=2.76
c52 12 0 6.56506e-20 $X=12.55 $Y=2.895
r53 20 22 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=11.07 $Y=2.195
+ $X2=11.07 $Y2=2.425
r54 15 17 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=13.33 $Y=2.48
+ $X2=13.33 $Y2=2.76
r55 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.165 $Y=2.395
+ $X2=13.33 $Y2=2.48
r56 13 14 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=13.165 $Y=2.395
+ $X2=12.635 $Y2=2.395
r57 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.55 $Y=2.48
+ $X2=12.635 $Y2=2.395
r58 11 12 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=12.55 $Y=2.48
+ $X2=12.55 $Y2=2.895
r59 9 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.465 $Y=2.98
+ $X2=12.55 $Y2=2.895
r60 9 10 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=12.465 $Y=2.98
+ $X2=11.235 $Y2=2.98
r61 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.15 $Y=2.895
+ $X2=11.235 $Y2=2.98
r62 8 22 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=11.15 $Y=2.895
+ $X2=11.15 $Y2=2.425
r63 2 17 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=13.19
+ $Y=2.55 $X2=13.33 $Y2=2.76
r64 1 20 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=10.925
+ $Y=1.985 $X2=11.07 $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%Q_N 1 2 7 8 9 10 11 12 13 22
r22 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=15.68 $Y=2.775
+ $X2=15.68 $Y2=2.9
r23 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=15.68 $Y=2.405
+ $X2=15.68 $Y2=2.775
r24 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=15.68 $Y=1.98
+ $X2=15.68 $Y2=2.405
r25 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=15.68 $Y=1.665
+ $X2=15.68 $Y2=1.98
r26 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=15.68 $Y=1.295
+ $X2=15.68 $Y2=1.665
r27 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=15.68 $Y=0.925
+ $X2=15.68 $Y2=1.295
r28 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=15.68 $Y=0.555
+ $X2=15.68 $Y2=0.925
r29 7 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=15.68 $Y=0.555
+ $X2=15.68 $Y2=0.43
r30 2 40 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=15.54
+ $Y=1.835 $X2=15.68 $Y2=2.9
r31 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.54
+ $Y=1.835 $X2=15.68 $Y2=1.98
r32 1 22 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=15.54
+ $Y=0.24 $X2=15.68 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%Q 1 2 7 8 9 10 11 12 13 22
r15 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=17.95 $Y=2.775
+ $X2=17.95 $Y2=2.9
r16 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.95 $Y=2.405
+ $X2=17.95 $Y2=2.775
r17 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=17.95 $Y=1.98
+ $X2=17.95 $Y2=2.405
r18 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=17.95 $Y=1.665
+ $X2=17.95 $Y2=1.98
r19 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.95 $Y=1.295
+ $X2=17.95 $Y2=1.665
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.95 $Y=0.925
+ $X2=17.95 $Y2=1.295
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.95 $Y=0.555
+ $X2=17.95 $Y2=0.925
r22 7 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=17.95 $Y=0.555
+ $X2=17.95 $Y2=0.43
r23 2 40 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=17.81
+ $Y=1.835 $X2=17.95 $Y2=2.9
r24 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=17.81
+ $Y=1.835 $X2=17.95 $Y2=1.98
r25 1 22 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=17.81
+ $Y=0.265 $X2=17.95 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_LP%VGND 1 2 3 4 5 6 20 23 25 29 33 37 41 47 49
+ 54 62 70 78 85 86 89 92 95 98 101 104
c152 86 0 5.56669e-20 $X=18 $Y=0
r153 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r154 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r155 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r156 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r157 93 96 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r158 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r159 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r160 86 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18 $Y=0 $X2=17.04
+ $Y2=0
r161 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18 $Y=0 $X2=18
+ $Y2=0
r162 83 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.325 $Y=0
+ $X2=17.16 $Y2=0
r163 83 85 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=17.325 $Y=0 $X2=18
+ $Y2=0
r164 82 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=17.04 $Y2=0
r165 82 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=14.64 $Y2=0
r166 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r167 79 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.82 $Y=0
+ $X2=14.655 $Y2=0
r168 79 81 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=14.82 $Y=0 $X2=15.12
+ $Y2=0
r169 78 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.995 $Y=0
+ $X2=17.16 $Y2=0
r170 78 81 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=16.995 $Y=0
+ $X2=15.12 $Y2=0
r171 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r172 76 77 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r173 74 77 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=14.16 $Y2=0
r174 74 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r175 73 76 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=14.16 $Y2=0
r176 73 74 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r177 71 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.965 $Y=0
+ $X2=10.8 $Y2=0
r178 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.965 $Y=0
+ $X2=11.28 $Y2=0
r179 70 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.49 $Y=0
+ $X2=14.655 $Y2=0
r180 70 76 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=14.49 $Y=0
+ $X2=14.16 $Y2=0
r181 69 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r182 68 69 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r183 66 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r184 65 68 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=7.44 $Y=0
+ $X2=10.32 $Y2=0
r185 65 66 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r186 63 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=0 $X2=7.075
+ $Y2=0
r187 63 65 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.24 $Y=0 $X2=7.44
+ $Y2=0
r188 62 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.8 $Y2=0
r189 62 68 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.32 $Y2=0
r190 61 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r191 60 61 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r192 58 61 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=4.56 $Y2=0
r193 58 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r194 57 60 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=4.56
+ $Y2=0
r195 57 58 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r196 55 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r197 55 57 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r198 54 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.88
+ $Y2=0
r199 54 60 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.56 $Y2=0
r200 52 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r201 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r202 49 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r203 49 51 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r204 47 69 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=10.32 $Y2=0
r205 47 66 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=7.44 $Y2=0
r206 41 43 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=17.16 $Y=0.41
+ $X2=17.16 $Y2=0.96
r207 39 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.16 $Y=0.085
+ $X2=17.16 $Y2=0
r208 39 41 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=17.16 $Y=0.085
+ $X2=17.16 $Y2=0.41
r209 35 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.655 $Y=0.085
+ $X2=14.655 $Y2=0
r210 35 37 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=14.655 $Y=0.085
+ $X2=14.655 $Y2=0.385
r211 31 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.8 $Y2=0
r212 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.8 $Y2=0.4
r213 27 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=0.085
+ $X2=7.075 $Y2=0
r214 27 29 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=7.075 $Y=0.085
+ $X2=7.075 $Y2=0.48
r215 26 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=4.88
+ $Y2=0
r216 25 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.91 $Y=0 $X2=7.075
+ $Y2=0
r217 25 26 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=6.91 $Y=0
+ $X2=5.045 $Y2=0
r218 21 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r219 21 23 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.405
r220 20 46 9.10249 $w=3.3e-07 $l=2.4e-07 $layer=LI1_cond $X=1.22 $Y=0.535
+ $X2=1.22 $Y2=0.775
r221 19 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r222 19 20 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.535
r223 6 43 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=16.905
+ $Y=0.685 $X2=17.16 $Y2=0.96
r224 6 41 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=16.905
+ $Y=0.685 $X2=17.16 $Y2=0.41
r225 5 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=14.515
+ $Y=0.24 $X2=14.655 $Y2=0.385
r226 4 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=10.66
+ $Y=0.255 $X2=10.8 $Y2=0.4
r227 3 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.865
+ $Y=0.335 $X2=7.075 $Y2=0.48
r228 2 23 182 $w=1.7e-07 $l=3.31134e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.58 $X2=4.88 $Y2=0.405
r229 1 46 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.58 $X2=1.22 $Y2=0.775
.ends

