* File: sky130_fd_sc_lp__or4_2.spice
* Created: Fri Aug 28 11:25:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4_2.pex.spice"
.subckt sky130_fd_sc_lp__or4_2  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1010 N_A_72_367#_M1010_d N_D_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_C_M1002_g N_A_72_367#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0903 AS=0.0588 PD=0.85 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_72_367#_M1000_d N_B_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0903 PD=0.7 PS=0.85 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_72_367#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.14 AS=0.0588 PD=0.973333 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1006_d N_A_72_367#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.28 AS=0.1176 PD=1.94667 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A_72_367#_M1011_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 A_155_367# N_D_M1008_g N_A_72_367#_M1008_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1005 A_227_367# N_C_M1005_g A_155_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=65.6601 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1001 A_335_367# N_B_M1001_g A_227_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0819 PD=0.81 PS=0.81 NRD=65.6601 NRS=65.6601 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_335_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.120225 AS=0.0819 PD=0.9375 PS=0.81 NRD=68.0044 NRS=65.6601 M=1 R=2.8
+ SA=75001.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_72_367#_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.17955 AS=0.360675 PD=1.545 PS=2.8125 NRD=0 NRS=9.8894 M=1 R=8.4
+ SA=75000.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_X_M1004_d N_A_72_367#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.17955 AS=0.3339 PD=1.545 PS=3.05 NRD=0.7683 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__or4_2.pxi.spice"
*
.ends
*
*
