* File: sky130_fd_sc_lp__einvn_4.pex.spice
* Created: Wed Sep  2 09:51:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVN_4%A 1 3 6 8 10 13 17 21 23 24 27 31 33 34 35
+ 36 37
r92 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.51 $X2=1.6 $Y2=1.51
r93 46 48 42.175 $w=3.6e-07 $l=3.15e-07 $layer=POLY_cond $X=1.285 $Y=1.485
+ $X2=1.6 $Y2=1.485
r94 45 49 13.652 $w=3.23e-07 $l=3.85e-07 $layer=LI1_cond $X=1.215 $Y=1.587
+ $X2=1.6 $Y2=1.587
r95 44 46 9.37222 $w=3.6e-07 $l=7e-08 $layer=POLY_cond $X=1.215 $Y=1.485
+ $X2=1.285 $Y2=1.485
r96 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=1.51 $X2=1.215 $Y2=1.51
r97 42 44 58.9111 $w=3.6e-07 $l=4.4e-07 $layer=POLY_cond $X=0.775 $Y=1.485
+ $X2=1.215 $Y2=1.485
r98 37 49 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.587 $X2=1.6
+ $Y2=1.587
r99 36 45 0.531897 $w=3.23e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.215 $Y2=1.587
r100 35 36 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=1.2 $Y2=1.587
r101 34 35 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.587
+ $X2=0.72 $Y2=1.587
r102 29 33 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.675
+ $X2=2.225 $Y2=1.51
r103 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.225 $Y=1.675
+ $X2=2.225 $Y2=2.465
r104 25 33 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.345
+ $X2=2.225 $Y2=1.51
r105 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.225 $Y=1.345
+ $X2=2.225 $Y2=0.765
r106 23 33 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=1.51
+ $X2=2.225 $Y2=1.51
r107 23 24 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.15 $Y=1.51
+ $X2=1.79 $Y2=1.51
r108 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.715 $Y=1.675
+ $X2=1.715 $Y2=2.465
r109 15 24 10.4642 $w=3.6e-07 $l=8.66025e-08 $layer=POLY_cond $X=1.715 $Y=1.485
+ $X2=1.79 $Y2=1.51
r110 15 19 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.715 $Y=1.485
+ $X2=1.715 $Y2=1.675
r111 15 48 15.3972 $w=3.6e-07 $l=1.15e-07 $layer=POLY_cond $X=1.715 $Y=1.485
+ $X2=1.6 $Y2=1.485
r112 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.715 $Y=1.345
+ $X2=1.715 $Y2=0.765
r113 11 46 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.285 $Y=1.675
+ $X2=1.285 $Y2=1.485
r114 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.285 $Y=1.675
+ $X2=1.285 $Y2=2.465
r115 8 46 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.285 $Y=1.295
+ $X2=1.285 $Y2=1.485
r116 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.285 $Y=1.295
+ $X2=1.285 $Y2=0.765
r117 4 42 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.775 $Y=1.675
+ $X2=0.775 $Y2=1.485
r118 4 6 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.775 $Y=1.675
+ $X2=0.775 $Y2=2.465
r119 1 42 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.775 $Y=1.295
+ $X2=0.775 $Y2=1.485
r120 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.775 $Y=1.295
+ $X2=0.775 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_4%A_555_201# 1 2 7 9 11 12 14 16 17 19 21 22
+ 24 26 27 28 29 30 34 40 43 44 48
r98 44 51 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.94 $Y=1.17 $X2=2.94
+ $Y2=1.26
r99 43 46 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.94 $Y=1.17
+ $X2=2.94 $Y2=1.485
r100 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.17 $X2=2.94 $Y2=1.17
r101 38 48 3.49899 $w=2.82e-07 $l=1.00846e-07 $layer=LI1_cond $X=5.525 $Y=1.395
+ $X2=5.502 $Y2=1.485
r102 38 40 43.2166 $w=2.58e-07 $l=9.75e-07 $layer=LI1_cond $X=5.525 $Y=1.395
+ $X2=5.525 $Y2=0.42
r103 34 36 35.1401 $w=3.03e-07 $l=9.3e-07 $layer=LI1_cond $X=5.502 $Y=1.98
+ $X2=5.502 $Y2=2.91
r104 32 48 3.49899 $w=2.82e-07 $l=9e-08 $layer=LI1_cond $X=5.502 $Y=1.575
+ $X2=5.502 $Y2=1.485
r105 32 34 15.3029 $w=3.03e-07 $l=4.05e-07 $layer=LI1_cond $X=5.502 $Y=1.575
+ $X2=5.502 $Y2=1.98
r106 31 46 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=1.485
+ $X2=2.94 $Y2=1.485
r107 30 48 3.00573 $w=1.8e-07 $l=1.52e-07 $layer=LI1_cond $X=5.35 $Y=1.485
+ $X2=5.502 $Y2=1.485
r108 30 31 138.328 $w=1.78e-07 $l=2.245e-06 $layer=LI1_cond $X=5.35 $Y=1.485
+ $X2=3.105 $Y2=1.485
r109 24 26 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.845 $Y=1.185
+ $X2=4.845 $Y2=0.655
r110 23 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.49 $Y=1.26
+ $X2=4.415 $Y2=1.26
r111 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.77 $Y=1.26
+ $X2=4.845 $Y2=1.185
r112 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.77 $Y=1.26
+ $X2=4.49 $Y2=1.26
r113 19 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.415 $Y=1.185
+ $X2=4.415 $Y2=1.26
r114 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.415 $Y=1.185
+ $X2=4.415 $Y2=0.655
r115 18 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.06 $Y=1.26
+ $X2=3.985 $Y2=1.26
r116 17 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.34 $Y=1.26
+ $X2=4.415 $Y2=1.26
r117 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.34 $Y=1.26
+ $X2=4.06 $Y2=1.26
r118 14 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.985 $Y=1.185
+ $X2=3.985 $Y2=1.26
r119 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.985 $Y=1.185
+ $X2=3.985 $Y2=0.655
r120 13 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.63 $Y=1.26
+ $X2=3.555 $Y2=1.26
r121 12 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.91 $Y=1.26
+ $X2=3.985 $Y2=1.26
r122 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.91 $Y=1.26
+ $X2=3.63 $Y2=1.26
r123 9 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.555 $Y=1.185
+ $X2=3.555 $Y2=1.26
r124 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.555 $Y=1.185
+ $X2=3.555 $Y2=0.655
r125 8 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.26
+ $X2=2.94 $Y2=1.26
r126 7 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.48 $Y=1.26
+ $X2=3.555 $Y2=1.26
r127 7 8 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=3.48 $Y=1.26
+ $X2=3.105 $Y2=1.26
r128 2 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.835 $X2=5.49 $Y2=2.91
r129 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.835 $X2=5.49 $Y2=1.98
r130 1 40 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.35
+ $Y=0.235 $X2=5.49 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_4%TE_B 1 3 4 5 6 8 9 11 13 14 16 18 19 21 25
+ 27 29 30 31 32 34 35 36 37 38 43 44
c90 25 0 1.07959e-19 $X=5.275 $Y=0.655
c91 1 0 8.21527e-20 $X=2.655 $Y=1.725
r92 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.61
+ $Y=1.91 $X2=4.61 $Y2=1.91
r93 37 38 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=4.597 $Y=2.405
+ $X2=4.597 $Y2=2.775
r94 36 37 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=4.597 $Y=2.035
+ $X2=4.597 $Y2=2.405
r95 36 44 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=4.597 $Y=2.035
+ $X2=4.597 $Y2=1.91
r96 33 43 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=4.61 $Y=1.725
+ $X2=4.61 $Y2=1.91
r97 33 34 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.61 $Y=1.725
+ $X2=4.61 $Y2=1.65
r98 27 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.275 $Y=1.725
+ $X2=5.275 $Y2=1.65
r99 27 29 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.275 $Y=1.725
+ $X2=5.275 $Y2=2.465
r100 23 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.275 $Y=1.575
+ $X2=5.275 $Y2=1.65
r101 23 25 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=5.275 $Y=1.575
+ $X2=5.275 $Y2=0.655
r102 22 34 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.775 $Y=1.65
+ $X2=4.61 $Y2=1.65
r103 21 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.2 $Y=1.65
+ $X2=5.275 $Y2=1.65
r104 21 22 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=5.2 $Y=1.65
+ $X2=4.775 $Y2=1.65
r105 20 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.02 $Y=1.65
+ $X2=3.945 $Y2=1.65
r106 19 34 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.65
+ $X2=4.61 $Y2=1.65
r107 19 20 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.445 $Y=1.65
+ $X2=4.02 $Y2=1.65
r108 16 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.945 $Y=1.725
+ $X2=3.945 $Y2=1.65
r109 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.945 $Y=1.725
+ $X2=3.945 $Y2=2.465
r110 15 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.59 $Y=1.65
+ $X2=3.515 $Y2=1.65
r111 14 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.87 $Y=1.65
+ $X2=3.945 $Y2=1.65
r112 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.87 $Y=1.65
+ $X2=3.59 $Y2=1.65
r113 11 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.515 $Y=1.725
+ $X2=3.515 $Y2=1.65
r114 11 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.515 $Y=1.725
+ $X2=3.515 $Y2=2.465
r115 10 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.16 $Y=1.65
+ $X2=3.085 $Y2=1.65
r116 9 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.44 $Y=1.65
+ $X2=3.515 $Y2=1.65
r117 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.44 $Y=1.65
+ $X2=3.16 $Y2=1.65
r118 6 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.085 $Y=1.725
+ $X2=3.085 $Y2=1.65
r119 6 8 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.085 $Y=1.725
+ $X2=3.085 $Y2=2.465
r120 4 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.01 $Y=1.65
+ $X2=3.085 $Y2=1.65
r121 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.01 $Y=1.65 $X2=2.73
+ $Y2=1.65
r122 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.655 $Y=1.725
+ $X2=2.73 $Y2=1.65
r123 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.655 $Y=1.725
+ $X2=2.655 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_4%A_87_367# 1 2 3 4 5 16 18 20 24 26 29 32 33
+ 36 40 44 50 53
r66 44 46 45.6073 $w=2.33e-07 $l=9.3e-07 $layer=LI1_cond $X=4.182 $Y=1.98
+ $X2=4.182 $Y2=2.91
r67 42 44 2.69721 $w=2.33e-07 $l=5.5e-08 $layer=LI1_cond $X=4.182 $Y=1.925
+ $X2=4.182 $Y2=1.98
r68 41 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.395 $Y=1.84 $X2=3.3
+ $Y2=1.84
r69 40 42 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=4.065 $Y=1.84
+ $X2=4.182 $Y2=1.925
r70 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.065 $Y=1.84
+ $X2=3.395 $Y2=1.84
r71 36 38 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.3 $Y=1.98 $X2=3.3
+ $Y2=2.91
r72 34 53 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=1.925 $X2=3.3
+ $Y2=1.84
r73 34 36 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=3.3 $Y=1.925 $X2=3.3
+ $Y2=1.98
r74 32 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.205 $Y=1.84 $X2=3.3
+ $Y2=1.84
r75 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.205 $Y=1.84
+ $X2=2.535 $Y2=1.84
r76 29 52 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=2.905
+ $X2=2.44 $Y2=2.99
r77 29 31 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=2.44 $Y=2.905
+ $X2=2.44 $Y2=1.98
r78 28 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.44 $Y=1.925
+ $X2=2.535 $Y2=1.84
r79 28 31 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=2.44 $Y=1.925
+ $X2=2.44 $Y2=1.98
r80 27 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.675 $Y=2.99
+ $X2=1.54 $Y2=2.99
r81 26 52 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.345 $Y=2.99
+ $X2=2.44 $Y2=2.99
r82 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.345 $Y=2.99
+ $X2=1.675 $Y2=2.99
r83 22 50 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.905
+ $X2=1.54 $Y2=2.99
r84 22 24 20.4879 $w=2.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.54 $Y=2.905
+ $X2=1.54 $Y2=2.425
r85 21 49 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.665 $Y=2.99
+ $X2=0.53 $Y2=2.99
r86 20 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.405 $Y=2.99
+ $X2=1.54 $Y2=2.99
r87 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.405 $Y=2.99
+ $X2=0.665 $Y2=2.99
r88 16 49 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.53 $Y=2.905
+ $X2=0.53 $Y2=2.99
r89 16 18 34.1465 $w=2.68e-07 $l=8e-07 $layer=LI1_cond $X=0.53 $Y=2.905 $X2=0.53
+ $Y2=2.105
r90 5 46 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=2.91
r91 5 44 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=1.98
r92 4 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.835 $X2=3.3 $Y2=2.91
r93 4 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.835 $X2=3.3 $Y2=1.98
r94 3 52 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.835 $X2=2.44 $Y2=2.91
r95 3 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.835 $X2=2.44 $Y2=1.98
r96 2 24 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.425
r97 1 49 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.435
+ $Y=1.835 $X2=0.56 $Y2=2.91
r98 1 18 400 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=0.435
+ $Y=1.835 $X2=0.56 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_4%Z 1 2 3 4 15 19 21 22 23 24 27 29 30 31 32
+ 33 38
c61 30 0 8.21527e-20 $X=2.06 $Y=1.92
r62 36 42 2.90198 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=1.075
+ $X2=2.045 $Y2=1.16
r63 33 42 4.84412 $w=3.4e-07 $l=1.35e-07 $layer=LI1_cond $X=2.045 $Y=1.295
+ $X2=2.045 $Y2=1.16
r64 32 36 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.045 $Y=0.925
+ $X2=2.045 $Y2=1.075
r65 32 38 7.05871 $w=3.98e-07 $l=2.45e-07 $layer=LI1_cond $X=2.045 $Y=0.925
+ $X2=2.045 $Y2=0.68
r66 30 31 3.351 $w=2.8e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.06 $Y=1.92
+ $X2=2.01 $Y2=2.005
r67 29 33 8.6392 $w=3.4e-07 $l=2.12368e-07 $layer=LI1_cond $X=2.06 $Y=1.5
+ $X2=2.045 $Y2=1.295
r68 29 30 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.06 $Y=1.5 $X2=2.06
+ $Y2=1.92
r69 25 31 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=2.09 $X2=2.01
+ $Y2=2.005
r70 25 27 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.01 $Y=2.09 $X2=2.01
+ $Y2=2.095
r71 23 31 3.18746 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.005
+ $X2=2.01 $Y2=2.005
r72 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.845 $Y=2.005
+ $X2=1.235 $Y2=2.005
r73 21 42 4.80115 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.845 $Y=1.16 $X2=2.045
+ $Y2=1.16
r74 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.845 $Y=1.16
+ $X2=1.155 $Y2=1.16
r75 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.07 $Y=2.09
+ $X2=1.235 $Y2=2.005
r76 17 19 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.07 $Y=2.09 $X2=1.07
+ $Y2=2.095
r77 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.99 $Y=1.075
+ $X2=1.155 $Y2=1.16
r78 13 15 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.99 $Y=1.075
+ $X2=0.99 $Y2=0.68
r79 4 27 300 $w=1.7e-07 $l=3.5327e-07 $layer=licon1_PDIFF $count=2 $X=1.79
+ $Y=1.835 $X2=2.01 $Y2=2.095
r80 3 19 300 $w=1.7e-07 $l=3.5327e-07 $layer=licon1_PDIFF $count=2 $X=0.85
+ $Y=1.835 $X2=1.07 $Y2=2.095
r81 2 38 91 $w=1.7e-07 $l=4.3119e-07 $layer=licon1_NDIFF $count=2 $X=1.79
+ $Y=0.345 $X2=2.01 $Y2=0.68
r82 1 15 91 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=2 $X=0.85
+ $Y=0.345 $X2=0.99 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_4%VPWR 1 2 3 12 16 20 26 30 31 32 41 48 49 52
+ 55
r74 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r76 49 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 46 55 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.037 $Y2=3.33
r79 46 48 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 45 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r82 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r83 42 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=3.73 $Y2=3.33
r84 42 44 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=4.56 $Y2=3.33
r85 41 55 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=5.037 $Y2=3.33
r86 41 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 36 40 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 35 39 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r91 32 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r92 32 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 30 39 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.87 $Y2=3.33
r95 26 29 39.2235 $w=2.83e-07 $l=9.7e-07 $layer=LI1_cond $X=5.037 $Y=1.98
+ $X2=5.037 $Y2=2.95
r96 24 55 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.037 $Y=3.245
+ $X2=5.037 $Y2=3.33
r97 24 29 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=5.037 $Y=3.245
+ $X2=5.037 $Y2=2.95
r98 20 23 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.73 $Y=2.18
+ $X2=3.73 $Y2=2.95
r99 18 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=3.245
+ $X2=3.73 $Y2=3.33
r100 18 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.73 $Y=3.245
+ $X2=3.73 $Y2=2.95
r101 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.87 $Y2=3.33
r102 16 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=3.33
+ $X2=3.73 $Y2=3.33
r103 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.565 $Y=3.33
+ $X2=3.035 $Y2=3.33
r104 12 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.87 $Y=2.18
+ $X2=2.87 $Y2=2.95
r105 10 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=3.33
r106 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=2.95
r107 3 29 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=1.835 $X2=5.06 $Y2=2.95
r108 3 26 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=1.835 $X2=5.06 $Y2=1.98
r109 2 23 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.95
r110 2 20 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.18
r111 1 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.835 $X2=2.87 $Y2=2.95
r112 1 12 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.835 $X2=2.87 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_4%A_83_69# 1 2 3 4 5 18 20 21 24 26 31 34 36
+ 41 44 46 47 50 52 53 54
c95 46 0 1.07959e-19 $X=4.535 $Y=1.14
r96 48 50 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=4.63 $Y=1.055
+ $X2=4.63 $Y2=0.42
r97 46 48 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.535 $Y=1.14
+ $X2=4.63 $Y2=1.055
r98 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.535 $Y=1.14
+ $X2=3.865 $Y2=1.14
r99 42 54 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.77 $Y=0.725
+ $X2=3.735 $Y2=0.81
r100 42 44 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.77 $Y=0.725
+ $X2=3.77 $Y2=0.42
r101 39 47 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.735 $Y=1.055
+ $X2=3.865 $Y2=1.14
r102 39 41 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=3.735 $Y=1.055
+ $X2=3.735 $Y2=0.93
r103 38 54 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.895
+ $X2=3.735 $Y2=0.81
r104 38 41 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=3.735 $Y=0.895
+ $X2=3.735 $Y2=0.93
r105 37 53 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.675 $Y=0.81
+ $X2=2.545 $Y2=0.81
r106 36 54 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.605 $Y=0.81
+ $X2=3.735 $Y2=0.81
r107 36 37 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.605 $Y=0.81
+ $X2=2.675 $Y2=0.81
r108 32 53 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=2.51 $Y=0.895
+ $X2=2.545 $Y2=0.81
r109 32 34 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.51 $Y=0.895
+ $X2=2.51 $Y2=1.04
r110 29 53 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0.725
+ $X2=2.545 $Y2=0.81
r111 29 31 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=2.545 $Y=0.725
+ $X2=2.545 $Y2=0.49
r112 28 31 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=2.545 $Y=0.425
+ $X2=2.545 $Y2=0.49
r113 27 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=0.34
+ $X2=1.5 $Y2=0.34
r114 26 28 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.415 $Y=0.34
+ $X2=2.545 $Y2=0.425
r115 26 27 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.415 $Y=0.34
+ $X2=1.665 $Y2=0.34
r116 22 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=0.425 $X2=1.5
+ $Y2=0.34
r117 22 24 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.5 $Y=0.425
+ $X2=1.5 $Y2=0.47
r118 20 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=0.34
+ $X2=1.5 $Y2=0.34
r119 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.335 $Y=0.34
+ $X2=0.645 $Y2=0.34
r120 16 21 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.51 $Y=0.425
+ $X2=0.645 $Y2=0.34
r121 16 18 2.7744 $w=2.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.51 $Y=0.425
+ $X2=0.51 $Y2=0.49
r122 5 50 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.49
+ $Y=0.235 $X2=4.63 $Y2=0.42
r123 4 44 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.235 $X2=3.77 $Y2=0.42
r124 4 41 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.235 $X2=3.77 $Y2=0.93
r125 3 34 182 $w=1.7e-07 $l=7.93079e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.345 $X2=2.51 $Y2=1.04
r126 3 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.345 $X2=2.51 $Y2=0.49
r127 2 24 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.36
+ $Y=0.345 $X2=1.5 $Y2=0.47
r128 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.415
+ $Y=0.345 $X2=0.54 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_4%VGND 1 2 3 12 14 18 22 24 25 26 35 42 43 46
+ 49
r70 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r71 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r72 43 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r73 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r74 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.06
+ $Y2=0
r75 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.52
+ $Y2=0
r76 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r77 39 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r78 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r79 36 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=0 $X2=4.2
+ $Y2=0
r80 36 38 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.365 $Y=0 $X2=4.56
+ $Y2=0
r81 35 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=0 $X2=5.06
+ $Y2=0
r82 35 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.56
+ $Y2=0
r83 34 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r84 33 34 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r85 29 33 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r86 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r87 26 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.12
+ $Y2=0
r88 26 30 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.24
+ $Y2=0
r89 24 33 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.12
+ $Y2=0
r90 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.34
+ $Y2=0
r91 20 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0
r92 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0.38
r93 16 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=0.085 $X2=4.2
+ $Y2=0
r94 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.2 $Y=0.085
+ $X2=4.2 $Y2=0.36
r95 15 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.34
+ $Y2=0
r96 14 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=4.2
+ $Y2=0
r97 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=3.505
+ $Y2=0
r98 10 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.34 $Y=0.085
+ $X2=3.34 $Y2=0
r99 10 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.34 $Y=0.085
+ $X2=3.34 $Y2=0.425
r100 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.92
+ $Y=0.235 $X2=5.06 $Y2=0.38
r101 2 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.06
+ $Y=0.235 $X2=4.2 $Y2=0.36
r102 1 12 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.235 $X2=3.34 $Y2=0.425
.ends

