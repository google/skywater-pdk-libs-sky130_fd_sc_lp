* File: sky130_fd_sc_lp__nor4_m.pex.spice
* Created: Fri Aug 28 10:57:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4_M%A 3 6 9 13 14 17 19 20 24
r39 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.355 $X2=0.525 $Y2=1.355
r40 20 25 9.78787 $w=3.63e-07 $l=3.1e-07 $layer=LI1_cond $X=0.622 $Y=1.665
+ $X2=0.622 $Y2=1.355
r41 19 25 1.89443 $w=3.63e-07 $l=6e-08 $layer=LI1_cond $X=0.622 $Y=1.295
+ $X2=0.622 $Y2=1.355
r42 15 17 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.615 $Y=2.175
+ $X2=0.795 $Y2=2.175
r43 13 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=1.695
+ $X2=0.525 $Y2=1.355
r44 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.695
+ $X2=0.525 $Y2=1.86
r45 12 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.19
+ $X2=0.525 $Y2=1.355
r46 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.795 $Y=2.25
+ $X2=0.795 $Y2=2.175
r47 7 9 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.795 $Y=2.25
+ $X2=0.795 $Y2=2.625
r48 6 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=2.1
+ $X2=0.615 $Y2=2.175
r49 6 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.615 $Y=2.1
+ $X2=0.615 $Y2=1.86
r50 3 12 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.615 $Y=0.56
+ $X2=0.615 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_M%B 3 7 11 12 13 14 18
r38 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.095
+ $Y=1.355 $X2=1.095 $Y2=1.355
r39 14 19 12.9912 $w=2.73e-07 $l=3.1e-07 $layer=LI1_cond $X=1.147 $Y=1.665
+ $X2=1.147 $Y2=1.355
r40 13 19 2.51442 $w=2.73e-07 $l=6e-08 $layer=LI1_cond $X=1.147 $Y=1.295
+ $X2=1.147 $Y2=1.355
r41 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.095 $Y=1.695
+ $X2=1.095 $Y2=1.355
r42 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.695
+ $X2=1.095 $Y2=1.86
r43 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.19
+ $X2=1.095 $Y2=1.355
r44 7 12 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.185 $Y=2.625
+ $X2=1.185 $Y2=1.86
r45 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.045 $Y=0.56
+ $X2=1.045 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_M%C 3 7 11 12 13 14 18
c37 3 0 1.08685e-19 $X=1.575 $Y=2.625
r38 13 14 22.1818 $w=1.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.672 $Y=1.295
+ $X2=1.672 $Y2=1.665
r39 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.665
+ $Y=1.355 $X2=1.665 $Y2=1.355
r40 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.665 $Y=1.695
+ $X2=1.665 $Y2=1.355
r41 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.695
+ $X2=1.665 $Y2=1.86
r42 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.19
+ $X2=1.665 $Y2=1.355
r43 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.715 $Y=0.56
+ $X2=1.715 $Y2=1.19
r44 3 12 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.575 $Y=2.625
+ $X2=1.575 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_M%D 3 7 9 12 14 15 16 21 23
r34 21 24 80.0222 $w=5.9e-07 $l=5.05e-07 $layer=POLY_cond $X=2.365 $Y=1.045
+ $X2=2.365 $Y2=1.55
r35 21 23 49.19 $w=5.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.045
+ $X2=2.365 $Y2=0.88
r36 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.495
+ $Y=1.045 $X2=2.495 $Y2=1.045
r37 15 16 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.567 $Y=1.295
+ $X2=2.567 $Y2=1.665
r38 15 22 9.14637 $w=3.13e-07 $l=2.5e-07 $layer=LI1_cond $X=2.567 $Y=1.295
+ $X2=2.567 $Y2=1.045
r39 14 22 4.39026 $w=3.13e-07 $l=1.2e-07 $layer=LI1_cond $X=2.567 $Y=0.925
+ $X2=2.567 $Y2=1.045
r40 10 12 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.965 $Y=2.175
+ $X2=2.145 $Y2=2.175
r41 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.145 $Y=2.1
+ $X2=2.145 $Y2=2.175
r42 9 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.145 $Y=2.1
+ $X2=2.145 $Y2=1.55
r43 7 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.145 $Y=0.56
+ $X2=2.145 $Y2=0.88
r44 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=2.25
+ $X2=1.965 $Y2=2.175
r45 1 3 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.965 $Y=2.25
+ $X2=1.965 $Y2=2.625
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_M%VPWR 1 6 9 10 11 21 22
r19 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r20 18 21 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r21 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r22 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 11 22 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r25 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 9 14 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 9 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.58 $Y2=3.33
r28 8 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.685 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 8 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.685 $Y=3.33
+ $X2=0.58 $Y2=3.33
r30 4 10 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.58 $Y=3.245
+ $X2=0.58 $Y2=3.33
r31 4 6 32.4805 $w=2.08e-07 $l=6.15e-07 $layer=LI1_cond $X=0.58 $Y=3.245
+ $X2=0.58 $Y2=2.63
r32 1 6 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.455
+ $Y=2.415 $X2=0.58 $Y2=2.63
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_M%Y 1 2 3 11 12 13 16 20 22 23 24 25 26 39
c59 20 0 1.08685e-19 $X=2.18 $Y=2.62
r60 25 26 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.925
+ $X2=1.68 $Y2=0.925
r61 25 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=0.925
+ $X2=0.935 $Y2=0.925
r62 24 32 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.785 $Y=0.925
+ $X2=0.935 $Y2=0.925
r63 24 39 7.03072 $w=4.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.785 $Y=0.84
+ $X2=0.785 $Y2=0.625
r64 23 26 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=0.925
+ $X2=1.68 $Y2=0.925
r65 22 24 14.1504 $w=3.38e-07 $l=3.75e-07 $layer=LI1_cond $X=0.26 $Y=0.925
+ $X2=0.635 $Y2=0.925
r66 18 20 20.8615 $w=2.08e-07 $l=3.95e-07 $layer=LI1_cond $X=2.18 $Y=2.225
+ $X2=2.18 $Y2=2.62
r67 14 23 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.93 $Y=0.84
+ $X2=1.825 $Y2=0.925
r68 14 16 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.93 $Y=0.84
+ $X2=1.93 $Y2=0.625
r69 12 18 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.075 $Y=2.14
+ $X2=2.18 $Y2=2.225
r70 12 13 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=2.075 $Y=2.14
+ $X2=0.26 $Y2=2.14
r71 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.175 $Y=2.055
+ $X2=0.26 $Y2=2.14
r72 10 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.175 $Y=1.01
+ $X2=0.26 $Y2=0.925
r73 10 11 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=0.175 $Y=1.01
+ $X2=0.175 $Y2=2.055
r74 3 20 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=2.415 $X2=2.18 $Y2=2.62
r75 2 16 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.35 $X2=1.93 $Y2=0.625
r76 1 39 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.35 $X2=0.83 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_M%VGND 1 2 3 10 12 16 20 23 24 25 27 37 38 44
r38 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r39 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 35 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r42 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r43 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r44 32 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=2.16
+ $Y2=0
r45 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r46 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r47 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 28 41 3.6162 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r49 28 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r50 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r51 27 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r52 25 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r53 25 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r54 23 34 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.16
+ $Y2=0
r55 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.36
+ $Y2=0
r56 22 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.64
+ $Y2=0
r57 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.36
+ $Y2=0
r58 18 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0
r59 18 20 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.495
r60 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r61 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.495
r62 10 41 3.29899 $w=2.1e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.227 $Y2=0
r63 10 12 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.35 $Y2=0.495
r64 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.22
+ $Y=0.35 $X2=2.36 $Y2=0.495
r65 2 16 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.35 $X2=1.28 $Y2=0.495
r66 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.35 $X2=0.35 $Y2=0.495
.ends

