* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__clkinv_1 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phighvt w=840000u l=150000u
+  ad=4.452e+11p pd=4.42e+06u as=2.352e+11p ps=2.24e+06u
M1001 VGND A Y VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.113e+11p ps=1.37e+06u
M1002 Y A VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
