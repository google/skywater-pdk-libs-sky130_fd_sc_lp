* File: sky130_fd_sc_lp__fa_4.spice
* Created: Fri Aug 28 10:35:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fa_4.pex.spice"
.subckt sky130_fd_sc_lp__fa_4  VNB VPB A CIN B VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* B	B
* CIN	CIN
* A	A
* VPB	VPB
* VNB	VNB
MM1030 N_VGND_M1030_d N_A_M1030_g N_A_37_131#_M1030_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75008.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_37_131#_M1005_d N_B_M1005_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0756 PD=0.8 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.7
+ SB=75008.3 A=0.063 P=1.14 MULT=1
MM1025 N_A_328_131#_M1025_d N_CIN_M1025_g N_A_37_131#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0798 PD=0.7 PS=0.8 NRD=0 NRS=28.56 M=1 R=2.8 SA=75001.2
+ SB=75007.7 A=0.063 P=1.14 MULT=1
MM1028 A_414_131# N_B_M1028_g N_A_328_131#_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75007.3 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_M1016_g A_414_131# VNB NSHORT L=0.15 W=0.42 AD=0.0924
+ AS=0.0441 PD=0.86 PS=0.63 NRD=5.712 NRS=14.28 M=1 R=2.8 SA=75002 SB=75007
+ A=0.063 P=1.14 MULT=1
MM1032 N_A_604_131#_M1032_d N_CIN_M1032_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=39.996 M=1 R=2.8
+ SA=75002.6 SB=75006.4 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_B_M1033_g N_A_604_131#_M1032_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0588 PD=0.81 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75003
+ SB=75005.9 A=0.063 P=1.14 MULT=1
MM1035 N_A_604_131#_M1035_d N_A_M1035_g N_VGND_M1033_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=25.704 M=1 R=2.8 SA=75003.6
+ SB=75005.4 A=0.063 P=1.14 MULT=1
MM1039 N_A_884_131#_M1039_d N_A_328_131#_M1039_g N_A_604_131#_M1035_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=11.424 NRS=0 M=1 R=2.8
+ SA=75004 SB=75005 A=0.063 P=1.14 MULT=1
MM1001 A_978_131# N_CIN_M1001_g N_A_884_131#_M1039_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.5
+ SB=75004.5 A=0.063 P=1.14 MULT=1
MM1008 A_1050_131# N_B_M1008_g A_978_131# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75004.8 SB=75004.1
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g A_1050_131# VNB NSHORT L=0.15 W=0.42 AD=0.0994
+ AS=0.0441 PD=0.843333 PS=0.63 NRD=51.9 NRS=14.28 M=1 R=2.8 SA=75005.2
+ SB=75003.8 A=0.063 P=1.14 MULT=1
MM1004 N_SUM_M1004_d N_A_884_131#_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1988 PD=1.12 PS=1.68667 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75003 SB=75003.2 A=0.126 P=1.98 MULT=1
MM1017 N_SUM_M1004_d N_A_884_131#_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.4
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1018 N_SUM_M1018_d N_A_884_131#_M1018_g N_VGND_M1017_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.9
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1021 N_SUM_M1018_d N_A_884_131#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.3
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1021_s N_A_328_131#_M1014_g N_COUT_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_A_328_131#_M1015_g N_COUT_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1034 N_VGND_M1015_d N_A_328_131#_M1034_g N_COUT_M1034_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1036 N_VGND_M1036_d N_A_328_131#_M1036_g N_COUT_M1034_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1038 N_VPWR_M1038_d N_A_M1038_g N_A_27_440#_M1038_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75007.5 A=0.096 P=1.58 MULT=1
MM1011 N_A_27_440#_M1011_d N_B_M1011_g N_VPWR_M1038_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.176325 AS=0.0896 PD=1.255 PS=0.92 NRD=29.2348 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75007.1 A=0.096 P=1.58 MULT=1
MM1024 N_A_328_131#_M1024_d N_CIN_M1024_g N_A_27_440#_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1392 AS=0.176325 PD=1.075 PS=1.255 NRD=47.6937 NRS=41.5473 M=1
+ R=4.26667 SA=75001.1 SB=75007.7 A=0.096 P=1.58 MULT=1
MM1019 A_445_419# N_B_M1019_g N_A_328_131#_M1024_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1392 PD=0.85 PS=1.075 NRD=15.3857 NRS=0 M=1 R=4.26667
+ SA=75001.7 SB=75007.2 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_445_419# VPB PHIGHVT L=0.15 W=0.64 AD=0.0912
+ AS=0.0672 PD=0.925 PS=0.85 NRD=1.5366 NRS=15.3857 M=1 R=4.26667 SA=75002.1
+ SB=75006.8 A=0.096 P=1.58 MULT=1
MM1026 N_A_604_419#_M1026_d N_CIN_M1026_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0912 PD=0.92 PS=0.925 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.5 SB=75006.4 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_B_M1009_g N_A_604_419#_M1026_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0896 PD=1.03 PS=0.92 NRD=16.9223 NRS=0 M=1 R=4.26667 SA=75002.9
+ SB=75005.9 A=0.096 P=1.58 MULT=1
MM1031 N_A_604_419#_M1031_d N_A_M1031_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1248 PD=0.92 PS=1.03 NRD=0 NRS=16.9223 M=1 R=4.26667 SA=75003.5
+ SB=75005.4 A=0.096 P=1.58 MULT=1
MM1012 N_A_884_131#_M1012_d N_A_328_131#_M1012_g N_A_604_419#_M1031_d VPB
+ PHIGHVT L=0.15 W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=6.1464 NRS=0 M=1
+ R=4.26667 SA=75003.9 SB=75005 A=0.096 P=1.58 MULT=1
MM1007 A_978_419# N_CIN_M1007_g N_A_884_131#_M1012_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1024 PD=0.85 PS=0.96 NRD=15.3857 NRS=6.1464 M=1 R=4.26667
+ SA=75004.4 SB=75004.5 A=0.096 P=1.58 MULT=1
MM1002 A_1050_419# N_B_M1002_g A_978_419# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0672 PD=0.85 PS=0.85 NRD=15.3857 NRS=15.3857 M=1 R=4.26667 SA=75004.7
+ SB=75004.1 A=0.096 P=1.58 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g A_1050_419# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.146964 AS=0.0672 PD=1.13516 PS=0.85 NRD=44.6205 NRS=15.3857 M=1 R=4.26667
+ SA=75005.1 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1029_d N_A_884_131#_M1000_g N_SUM_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.289336 AS=0.1764 PD=2.23484 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_884_131#_M1013_g N_SUM_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1020 N_VPWR_M1013_d N_A_884_131#_M1020_g N_SUM_M1020_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1027 N_VPWR_M1027_d N_A_884_131#_M1027_g N_SUM_M1020_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1027_d N_A_328_131#_M1010_g N_COUT_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.7
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_328_131#_M1022_g N_COUT_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1022_d N_A_328_131#_M1023_g N_COUT_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1037_d N_A_328_131#_M1037_g N_COUT_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=18.6127 P=23.69
*
.include "sky130_fd_sc_lp__fa_4.pxi.spice"
*
.ends
*
*
