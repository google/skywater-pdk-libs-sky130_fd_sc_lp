* File: sky130_fd_sc_lp__einvp_4.spice
* Created: Fri Aug 28 10:33:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvp_4.pex.spice"
.subckt sky130_fd_sc_lp__einvp_4  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_TE_M1016_g N_A_35_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1016_d N_TE_M1005_g N_A_204_47#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_TE_M1006_g N_A_204_47#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1006_d N_TE_M1014_g N_A_204_47#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_TE_M1017_g N_A_204_47#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_Z_M1003_d N_A_M1003_g N_A_204_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2898 AS=0.1176 PD=2.37 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.3
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1008 N_Z_M1008_d N_A_M1008_g N_A_204_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1011 N_Z_M1008_d N_A_M1011_g N_A_204_47#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=1.428 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1013 N_Z_M1013_d N_A_M1013_g N_A_204_47#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_TE_M1004_g N_A_35_47#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A_35_47#_M1000_g N_A_301_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1000_d N_A_35_47#_M1007_g N_A_301_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A_35_47#_M1012_g N_A_301_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1012_d N_A_35_47#_M1015_g N_A_301_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3969 PD=1.54 PS=1.89 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1001 N_A_301_367#_M1015_s N_A_M1001_g N_Z_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3969 AS=0.1764 PD=1.89 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 N_A_301_367#_M1002_d N_A_M1002_g N_Z_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_A_301_367#_M1002_d N_A_M1009_g N_Z_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_301_367#_M1010_d N_A_M1010_g N_Z_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__einvp_4.pxi.spice"
*
.ends
*
*
