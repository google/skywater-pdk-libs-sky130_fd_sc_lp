* File: sky130_fd_sc_lp__inv_m.pxi.spice
* Created: Wed Sep  2 09:56:19 2020
* 
x_PM_SKY130_FD_SC_LP__INV_M%A N_A_M1000_g N_A_M1001_g A A A A N_A_c_21_n
+ N_A_c_22_n N_A_c_23_n PM_SKY130_FD_SC_LP__INV_M%A
x_PM_SKY130_FD_SC_LP__INV_M%VPWR N_VPWR_M1001_s N_VPWR_c_41_n N_VPWR_c_42_n VPWR
+ N_VPWR_c_43_n N_VPWR_c_40_n PM_SKY130_FD_SC_LP__INV_M%VPWR
x_PM_SKY130_FD_SC_LP__INV_M%Y N_Y_M1000_d N_Y_M1001_d Y Y Y Y Y Y N_Y_c_53_n
+ PM_SKY130_FD_SC_LP__INV_M%Y
x_PM_SKY130_FD_SC_LP__INV_M%VGND N_VGND_M1000_s N_VGND_c_63_n N_VGND_c_64_n VGND
+ N_VGND_c_65_n N_VGND_c_66_n PM_SKY130_FD_SC_LP__INV_M%VGND
cc_1 VNB N_A_M1000_g 0.0286097f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.56
cc_2 VNB N_A_M1001_g 0.00169337f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.52
cc_3 VNB N_A_c_21_n 0.106199f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_4 VNB N_A_c_22_n 0.00124579f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_5 VNB N_A_c_23_n 0.00673884f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.055
cc_6 VNB N_VPWR_c_40_n 0.0442671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_Y_c_53_n 0.0439506f $X=-0.19 $Y=-0.245 $X2=0.332 $Y2=0.955
cc_8 VNB N_VGND_c_63_n 0.0111188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_64_n 0.0105254f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.52
cc_10 VNB N_VGND_c_65_n 0.0200473f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_11 VNB N_VGND_c_66_n 0.0980881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VPB N_A_M1001_g 0.0550429f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.52
cc_13 VPB N_A_c_22_n 0.0238206f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_14 VPB N_VPWR_c_41_n 0.0114776f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_15 VPB N_VPWR_c_42_n 0.0291231f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.52
cc_16 VPB N_VPWR_c_43_n 0.0191968f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_17 VPB N_VPWR_c_40_n 0.0560048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB N_Y_c_53_n 0.046411f $X=-0.19 $Y=1.655 $X2=0.332 $Y2=0.955
cc_19 N_A_M1001_g N_VPWR_c_42_n 0.00385941f $X=0.485 $Y=2.52 $X2=0 $Y2=0
cc_20 N_A_c_21_n N_VPWR_c_42_n 0.00113233f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_21 N_A_c_22_n N_VPWR_c_42_n 0.0169111f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_22 N_A_M1001_g N_VPWR_c_43_n 0.00428744f $X=0.485 $Y=2.52 $X2=0 $Y2=0
cc_23 N_A_M1001_g N_VPWR_c_40_n 0.00476395f $X=0.485 $Y=2.52 $X2=0 $Y2=0
cc_24 N_A_M1000_g N_Y_c_53_n 0.0481793f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_25 N_A_c_22_n N_Y_c_53_n 0.0625068f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_26 N_A_c_23_n N_Y_c_53_n 0.0121009f $X=0.255 $Y=1.055 $X2=0 $Y2=0
cc_27 N_A_M1000_g N_VGND_c_64_n 0.00494422f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_28 N_A_c_21_n N_VGND_c_64_n 0.00114553f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_29 N_A_c_23_n N_VGND_c_64_n 0.0152344f $X=0.255 $Y=1.055 $X2=0 $Y2=0
cc_30 N_A_M1000_g N_VGND_c_65_n 0.00478016f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_31 N_A_M1000_g N_VGND_c_66_n 0.00976615f $X=0.485 $Y=0.56 $X2=0 $Y2=0
cc_32 N_A_c_23_n N_VGND_c_66_n 0.00102874f $X=0.255 $Y=1.055 $X2=0 $Y2=0
cc_33 N_VPWR_c_42_n N_Y_c_53_n 0.0154405f $X=0.27 $Y=2.525 $X2=0 $Y2=0
cc_34 N_VPWR_c_43_n N_Y_c_53_n 0.00859063f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_35 N_VPWR_c_40_n N_Y_c_53_n 0.0075889f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_36 N_Y_c_53_n N_VGND_c_65_n 0.00617369f $X=0.7 $Y=0.61 $X2=0 $Y2=0
cc_37 N_Y_c_53_n N_VGND_c_66_n 0.00722785f $X=0.7 $Y=0.61 $X2=0 $Y2=0
