* File: sky130_fd_sc_lp__a31oi_m.pex.spice
* Created: Wed Sep  2 09:27:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31OI_M%A3 2 3 4 5 6 7 9 10 12 15 16 17 18 19 20 27
r36 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.105 $X2=0.27 $Y2=1.105
r37 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r38 18 19 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r39 17 18 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r40 17 28 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.105
r41 16 28 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.105
r42 14 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.445
+ $X2=0.27 $Y2=1.105
r43 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.445
+ $X2=0.27 $Y2=1.61
r44 13 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.09
+ $X2=0.27 $Y2=1.105
r45 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.87 $Y=0.94
+ $X2=0.87 $Y2=0.62
r46 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.77 $Y=2.39 $X2=0.77
+ $Y2=2.71
r47 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.695 $Y=2.315
+ $X2=0.77 $Y2=2.39
r48 5 6 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=0.695 $Y=2.315
+ $X2=0.435 $Y2=2.315
r49 4 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=1.015
+ $X2=0.27 $Y2=1.09
r50 3 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.795 $Y=1.015
+ $X2=0.87 $Y2=0.94
r51 3 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=0.795 $Y=1.015
+ $X2=0.435 $Y2=1.015
r52 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.36 $Y=2.24
+ $X2=0.435 $Y2=2.315
r53 2 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.24 $X2=0.36
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_M%A2 3 7 11 12 13 14 15 16 17 24
c44 3 0 1.44336e-19 $X=1.2 $Y=2.71
r45 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.495 $X2=1.14 $Y2=1.495
r46 16 17 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=2.035
r47 16 25 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.495
r48 15 25 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=1.17 $Y=1.295 $X2=1.17
+ $Y2=1.495
r49 14 15 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=0.925
+ $X2=1.17 $Y2=1.295
r50 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=0.555
+ $X2=1.17 $Y2=0.925
r51 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.14 $Y=1.835
+ $X2=1.14 $Y2=1.495
r52 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.835
+ $X2=1.14 $Y2=2
r53 10 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.33
+ $X2=1.14 $Y2=1.495
r54 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.23 $Y=0.62 $X2=1.23
+ $Y2=1.33
r55 3 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.2 $Y=2.71 $X2=1.2
+ $Y2=2
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_M%A1 3 7 11 12 13 14 15 16 17 24
c51 13 0 1.44336e-19 $X=1.68 $Y=0.555
c52 3 0 1.30505e-19 $X=1.59 $Y=0.62
r53 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.495 $X2=1.68 $Y2=1.495
r54 16 17 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=2.035
r55 16 25 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.495
r56 15 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.68 $Y=1.295 $X2=1.68
+ $Y2=1.495
r57 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=0.925
+ $X2=1.68 $Y2=1.295
r58 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=0.555
+ $X2=1.68 $Y2=0.925
r59 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.68 $Y=1.835
+ $X2=1.68 $Y2=1.495
r60 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.835
+ $X2=1.68 $Y2=2
r61 10 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.33
+ $X2=1.68 $Y2=1.495
r62 7 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.63 $Y=2.71 $X2=1.63
+ $Y2=2
r63 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.59 $Y=0.62 $X2=1.59
+ $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_M%B1 1 3 5 8 12 16 17 18 19 20 25
c49 18 0 1.30505e-19 $X=2.16 $Y=1.295
r50 20 27 14.7455 $w=2.3e-07 $l=2.7e-07 $layer=LI1_cond $X=2.19 $Y=2.035
+ $X2=2.19 $Y2=1.765
r51 19 27 5.01062 $w=2.28e-07 $l=1e-07 $layer=LI1_cond $X=2.19 $Y=1.665 $X2=2.19
+ $Y2=1.765
r52 18 19 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=1.295
+ $X2=2.19 $Y2=1.665
r53 18 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.22
+ $Y=1.375 $X2=2.22 $Y2=1.375
r54 16 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.22 $Y=1.715
+ $X2=2.22 $Y2=1.375
r55 16 17 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.715
+ $X2=2.22 $Y2=1.88
r56 15 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.21
+ $X2=2.22 $Y2=1.375
r57 10 12 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.06 $Y=2.315 $X2=2.16
+ $Y2=2.315
r58 8 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.31 $Y=0.62 $X2=2.31
+ $Y2=1.21
r59 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=2.24 $X2=2.16
+ $Y2=2.315
r60 5 17 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.16 $Y=2.24 $X2=2.16
+ $Y2=1.88
r61 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=2.39 $X2=2.06
+ $Y2=2.315
r62 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.06 $Y=2.39 $X2=2.06
+ $Y2=2.71
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_M%VPWR 1 2 9 13 16 17 19 20 21 34 35
r34 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r37 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 21 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 21 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 19 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.25 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.415 $Y2=3.33
r45 18 31 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.58 $Y=3.33 $X2=1.68
+ $Y2=3.33
r46 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=3.33
+ $X2=1.415 $Y2=3.33
r47 16 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.39 $Y=3.33 $X2=0.24
+ $Y2=3.33
r48 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.555 $Y2=3.33
r49 15 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=0.555 $Y2=3.33
r51 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=3.245
+ $X2=1.415 $Y2=3.33
r52 11 13 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.415 $Y=3.245
+ $X2=1.415 $Y2=2.795
r53 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.555 $Y=3.245
+ $X2=0.555 $Y2=3.33
r54 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.555 $Y=3.245
+ $X2=0.555 $Y2=2.775
r55 2 13 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=2.5 $X2=1.415 $Y2=2.795
r56 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.43
+ $Y=2.5 $X2=0.555 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_M%A_169_500# 1 2 9 11 12 15
r22 13 15 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=1.855 $Y=2.51
+ $X2=1.855 $Y2=2.625
r23 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.76 $Y=2.425
+ $X2=1.855 $Y2=2.51
r24 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.76 $Y=2.425
+ $X2=1.07 $Y2=2.425
r25 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.985 $Y=2.51
+ $X2=1.07 $Y2=2.425
r26 7 9 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.985 $Y=2.51
+ $X2=0.985 $Y2=2.625
r27 2 15 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=2.5 $X2=1.845 $Y2=2.625
r28 1 9 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.845
+ $Y=2.5 $X2=0.985 $Y2=2.625
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_M%Y 1 2 9 11 15 16 19
c33 9 0 1.64292e-19 $X=2.075 $Y=0.685
r34 18 19 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=2.64 $Y=2.48
+ $X2=2.64 $Y2=1.295
r35 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.64 $Y=1.01
+ $X2=2.64 $Y2=1.295
r36 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.555 $Y=0.925
+ $X2=2.64 $Y2=1.01
r37 15 16 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.555 $Y=0.925
+ $X2=2.18 $Y2=0.925
r38 11 18 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.555 $Y=2.645
+ $X2=2.64 $Y2=2.48
r39 11 13 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.555 $Y=2.645
+ $X2=2.275 $Y2=2.645
r40 7 16 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.075 $Y=0.84
+ $X2=2.18 $Y2=0.925
r41 7 9 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=2.075 $Y=0.84
+ $X2=2.075 $Y2=0.685
r42 2 13 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=2.5 $X2=2.275 $Y2=2.645
r43 1 9 182 $w=1.7e-07 $l=5.29953e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.41 $X2=2.075 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_M%VGND 1 2 9 11 13 15 17 22 31 35
r31 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r32 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r34 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r36 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r37 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.655
+ $Y2=0
r39 23 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.2
+ $Y2=0
r40 22 34 4.5891 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.62
+ $Y2=0
r41 22 28 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.16
+ $Y2=0
r42 20 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r43 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.49 $Y=0 $X2=0.655
+ $Y2=0
r45 17 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.49 $Y=0 $X2=0.24
+ $Y2=0
r46 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r47 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r48 11 34 3.17707 $w=3.3e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.62 $Y2=0
r49 11 13 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0.555
r50 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.655 $Y=0.085
+ $X2=0.655 $Y2=0
r51 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.655 $Y=0.085
+ $X2=0.655 $Y2=0.555
r52 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.41 $X2=2.525 $Y2=0.555
r53 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.53
+ $Y=0.41 $X2=0.655 $Y2=0.555
.ends

