* File: sky130_fd_sc_lp__and4_m.spice
* Created: Wed Sep  2 09:33:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4_m.pex.spice"
.subckt sky130_fd_sc_lp__and4_m  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_136_47# N_A_M1002_g N_A_53_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1008 A_208_47# N_B_M1008_g A_136_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1000 A_316_47# N_C_M1000_g A_208_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_D_M1003_g A_316_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=8.568 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_53_47#_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=22.848 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_53_47#_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_53_47#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_53_47#_M1009_d N_C_M1009_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_D_M1006_g N_A_53_47#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_53_47#_M1004_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__and4_m.pxi.spice"
*
.ends
*
*
