* File: sky130_fd_sc_lp__dfsbp_2.pex.spice
* Created: Wed Sep  2 09:44:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFSBP_2%CLK 3 7 9 10 14 15
r26 14 17 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.467 $Y=1.65
+ $X2=0.467 $Y2=1.815
r27 14 16 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.467 $Y=1.65
+ $X2=0.467 $Y2=1.485
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.455
+ $Y=1.65 $X2=0.455 $Y2=1.65
r29 9 10 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=2.035
r30 9 15 0.394312 $w=4.53e-07 $l=1.5e-08 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=1.65
r31 7 17 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.57 $Y=2.295
+ $X2=0.57 $Y2=1.815
r32 3 16 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.57 $Y=1.105
+ $X2=0.57 $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_129_179# 1 2 7 11 12 14 17 19 20 23 27 31
+ 36 39 40 41 44 45 47 50 51 52 54 57 58 60 63 64 65 67 68 69 70 77 78 83 84 88
+ 89 90 91 96 97 105
c265 97 0 8.27457e-20 $X=6.815 $Y=1.52
c266 96 0 1.54738e-19 $X=6.815 $Y=1.52
c267 88 0 1.52427e-19 $X=1.51 $Y=1.32
c268 68 0 7.7085e-20 $X=6.025 $Y=1.25
c269 64 0 4.60718e-20 $X=4.975 $Y=0.617
c270 54 0 5.68328e-20 $X=3.555 $Y=1.125
c271 23 0 1.26652e-19 $X=3.43 $Y=2.885
c272 20 0 1.38789e-19 $X=2.965 $Y=1.49
c273 17 0 4.45677e-20 $X=2.89 $Y=0.835
c274 12 0 1.23604e-19 $X=1.86 $Y=3.075
r275 96 97 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.815
+ $Y=1.52 $X2=6.815 $Y2=1.52
r276 91 93 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.11 $Y=1.25
+ $X2=6.11 $Y2=1.44
r277 88 105 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.51 $Y=1.32
+ $X2=1.51 $Y2=1.155
r278 87 89 8.94374 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=1.25
+ $X2=1.675 $Y2=1.25
r279 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.32 $X2=1.51 $Y2=1.32
r280 84 102 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.05 $Y=2.94
+ $X2=1.05 $Y2=3.15
r281 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=2.94 $X2=1.05 $Y2=2.94
r282 80 83 8.25918 $w=2.98e-07 $l=2.15e-07 $layer=LI1_cond $X=0.835 $Y=2.925
+ $X2=1.05 $Y2=2.925
r283 77 79 7.93859 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=0.82 $Y=2.455
+ $X2=0.82 $Y2=2.63
r284 77 78 7.49534 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=2.455
+ $X2=0.82 $Y2=2.29
r285 71 93 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=1.44
+ $X2=6.11 $Y2=1.44
r286 70 96 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.65 $Y=1.44
+ $X2=6.78 $Y2=1.44
r287 70 71 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.65 $Y=1.44
+ $X2=6.195 $Y2=1.44
r288 68 91 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=1.25
+ $X2=6.11 $Y2=1.25
r289 68 69 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=6.025 $Y=1.25
+ $X2=5.145 $Y2=1.25
r290 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.06 $Y=1.165
+ $X2=5.145 $Y2=1.25
r291 66 67 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.06 $Y=0.72
+ $X2=5.06 $Y2=1.165
r292 64 66 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=4.975 $Y=0.617
+ $X2=5.06 $Y2=0.72
r293 64 65 29.7561 $w=2.03e-07 $l=5.5e-07 $layer=LI1_cond $X=4.975 $Y=0.617
+ $X2=4.425 $Y2=0.617
r294 62 65 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=4.34 $Y=0.72
+ $X2=4.425 $Y2=0.617
r295 62 63 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.34 $Y=0.72
+ $X2=4.34 $Y2=1.125
r296 61 90 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.655 $Y=1.21
+ $X2=3.56 $Y2=1.21
r297 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.255 $Y=1.21
+ $X2=4.34 $Y2=1.125
r298 60 61 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.255 $Y=1.21
+ $X2=3.655 $Y2=1.21
r299 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.56
+ $Y=1.68 $X2=3.56 $Y2=1.68
r300 55 90 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=1.295
+ $X2=3.56 $Y2=1.21
r301 55 57 22.4737 $w=1.88e-07 $l=3.85e-07 $layer=LI1_cond $X=3.56 $Y=1.295
+ $X2=3.56 $Y2=1.68
r302 54 90 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=3.555 $Y=1.125
+ $X2=3.56 $Y2=1.21
r303 53 54 43.1313 $w=1.78e-07 $l=7e-07 $layer=LI1_cond $X=3.555 $Y=0.425
+ $X2=3.555 $Y2=1.125
r304 51 53 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.465 $Y=0.34
+ $X2=3.555 $Y2=0.425
r305 51 52 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=3.465 $Y=0.34
+ $X2=2.41 $Y2=0.34
r306 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.325 $Y=0.425
+ $X2=2.41 $Y2=0.34
r307 49 50 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.325 $Y=0.425
+ $X2=2.325 $Y2=1.015
r308 47 50 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.24 $Y=1.105
+ $X2=2.325 $Y2=1.015
r309 47 89 34.8131 $w=1.78e-07 $l=5.65e-07 $layer=LI1_cond $X=2.24 $Y=1.105
+ $X2=1.675 $Y2=1.105
r310 46 75 2.90196 $w=4.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=1.25
+ $X2=0.785 $Y2=1.25
r311 45 87 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=1.44 $Y=1.25 $X2=1.51
+ $Y2=1.25
r312 45 46 12.4698 $w=4.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.44 $Y=1.25
+ $X2=0.95 $Y2=1.25
r313 44 80 2.29563 $w=2.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.835 $Y=2.775
+ $X2=0.835 $Y2=2.925
r314 44 79 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.835 $Y=2.775
+ $X2=0.835 $Y2=2.63
r315 41 75 5.01248 $w=2.3e-07 $l=2.58795e-07 $layer=LI1_cond $X=0.835 $Y=1.485
+ $X2=0.785 $Y2=1.25
r316 41 78 40.3355 $w=2.28e-07 $l=8.05e-07 $layer=LI1_cond $X=0.835 $Y=1.485
+ $X2=0.835 $Y2=2.29
r317 39 97 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.815 $Y=1.86
+ $X2=6.815 $Y2=1.52
r318 39 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.86
+ $X2=6.815 $Y2=2.025
r319 38 97 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.355
+ $X2=6.815 $Y2=1.52
r320 35 58 49.9064 $w=3.7e-07 $l=3.2e-07 $layer=POLY_cond $X=3.54 $Y=2 $X2=3.54
+ $Y2=1.68
r321 35 36 49.8761 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.54 $Y=2 $X2=3.54
+ $Y2=2.185
r322 34 58 2.33936 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=3.54 $Y=1.665
+ $X2=3.54 $Y2=1.68
r323 31 38 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.74 $Y=1.005
+ $X2=6.74 $Y2=1.355
r324 27 40 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=6.725 $Y=2.675
+ $X2=6.725 $Y2=2.025
r325 23 36 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=3.43 $Y=2.885
+ $X2=3.43 $Y2=2.185
r326 19 34 80.1144 $w=1.81e-07 $l=3.19022e-07 $layer=POLY_cond $X=3.245 $Y=1.49
+ $X2=3.54 $Y2=1.54
r327 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.245 $Y=1.49
+ $X2=2.965 $Y2=1.49
r328 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.89 $Y=1.415
+ $X2=2.965 $Y2=1.49
r329 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.89 $Y=1.415
+ $X2=2.89 $Y2=0.835
r330 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.86 $Y=3.075
+ $X2=1.86 $Y2=2.645
r331 11 105 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.6 $Y=0.835
+ $X2=1.6 $Y2=1.155
r332 8 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=3.15
+ $X2=1.05 $Y2=3.15
r333 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.785 $Y=3.15
+ $X2=1.86 $Y2=3.075
r334 7 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.785 $Y=3.15
+ $X2=1.215 $Y2=3.15
r335 2 77 600 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.975 $X2=0.785 $Y2=2.455
r336 1 75 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.895 $X2=0.785 $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%D 3 7 9 10 11 16 20
c46 20 0 1.10806e-19 $X=2.51 $Y=2.35
c47 16 0 7.7582e-21 $X=2.08 $Y=1.45
c48 11 0 3.35784e-19 $X=2.16 $Y=2.405
r49 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=2.35
+ $X2=2.51 $Y2=2.515
r50 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=2.35 $X2=2.51 $Y2=2.35
r51 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.45 $X2=2.08 $Y2=1.45
r52 11 21 1.10726 $w=6.06e-07 $l=5.5e-08 $layer=LI1_cond $X=2.255 $Y=2.405
+ $X2=2.255 $Y2=2.35
r53 10 21 6.34158 $w=6.06e-07 $l=3.15e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=2.255 $Y2=2.35
r54 9 10 7.44884 $w=6.06e-07 $l=3.7e-07 $layer=LI1_cond $X=2.255 $Y=1.665
+ $X2=2.255 $Y2=2.035
r55 9 17 4.32838 $w=6.06e-07 $l=2.89569e-07 $layer=LI1_cond $X=2.255 $Y=1.665
+ $X2=2.08 $Y2=1.45
r56 7 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.53 $Y=2.885
+ $X2=2.53 $Y2=2.515
r57 1 16 74.7592 $w=2.45e-07 $l=4.55082e-07 $layer=POLY_cond $X=2.46 $Y=1.285
+ $X2=2.08 $Y2=1.45
r58 1 3 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.46 $Y=1.285 $X2=2.46
+ $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_721_99# 1 2 7 9 12 14 15 16 17 22 25 29 30
+ 32 33 36 40 42 49 51
c102 49 0 2.62346e-19 $X=4.13 $Y=1.715
c103 40 0 1.53526e-19 $X=5.625 $Y=2.885
c104 33 0 4.20846e-20 $X=4.345 $Y=2.58
c105 29 0 8.45674e-20 $X=4.26 $Y=2.35
c106 25 0 7.3458e-20 $X=4.13 $Y=1.55
c107 22 0 2.62794e-20 $X=4.595 $Y=1.555
c108 7 0 1.46742e-19 $X=3.68 $Y=1.155
r109 49 51 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.17 $Y=1.715 $X2=4.17
+ $Y2=2.185
r110 42 45 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.995 $Y=2.58
+ $X2=4.995 $Y2=2.885
r111 38 45 0.460977 $w=2.98e-07 $l=1.2e-08 $layer=LI1_cond $X=4.995 $Y=2.897
+ $X2=4.995 $Y2=2.885
r112 38 40 15.5823 $w=3.53e-07 $l=4.8e-07 $layer=LI1_cond $X=5.145 $Y=2.897
+ $X2=5.625 $Y2=2.897
r113 34 36 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=4.695 $Y=1.465
+ $X2=4.695 $Y2=1.055
r114 32 42 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.845 $Y=2.58
+ $X2=4.995 $Y2=2.58
r115 32 33 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.845 $Y=2.58
+ $X2=4.345 $Y2=2.58
r116 30 52 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=4.26 $Y=2.35
+ $X2=4.26 $Y2=2.47
r117 30 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.26 $Y=2.35
+ $X2=4.26 $Y2=2.185
r118 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.26
+ $Y=2.35 $X2=4.26 $Y2=2.35
r119 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.26 $Y=2.495
+ $X2=4.345 $Y2=2.58
r120 27 29 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.26 $Y=2.495
+ $X2=4.26 $Y2=2.35
r121 25 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.55
+ $X2=4.13 $Y2=1.715
r122 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.55 $X2=4.13 $Y2=1.55
r123 22 34 6.84108 $w=1.8e-07 $l=1.3784e-07 $layer=LI1_cond $X=4.595 $Y=1.555
+ $X2=4.695 $Y2=1.465
r124 22 24 28.6515 $w=1.78e-07 $l=4.65e-07 $layer=LI1_cond $X=4.595 $Y=1.555
+ $X2=4.13 $Y2=1.555
r125 18 25 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=4.13 $Y=1.305
+ $X2=4.13 $Y2=1.55
r126 16 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=2.47
+ $X2=4.26 $Y2=2.47
r127 16 17 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.095 $Y=2.47
+ $X2=3.865 $Y2=2.47
r128 14 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.965 $Y=1.23
+ $X2=4.13 $Y2=1.305
r129 14 15 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.965 $Y=1.23
+ $X2=3.755 $Y2=1.23
r130 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.79 $Y=2.545
+ $X2=3.865 $Y2=2.47
r131 10 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.79 $Y=2.545
+ $X2=3.79 $Y2=2.885
r132 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.68 $Y=1.155
+ $X2=3.755 $Y2=1.23
r133 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.68 $Y=1.155
+ $X2=3.68 $Y2=0.835
r134 2 45 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=2.675 $X2=4.94 $Y2=2.885
r135 2 40 600 $w=1.7e-07 $l=9.24054e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=2.675 $X2=5.625 $Y2=2.885
r136 1 36 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.565
+ $Y=0.845 $X2=4.69 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_593_125# 1 2 9 13 15 17 18 19 21 24 26 29
+ 31 34 36 39 40 41 44 45 48 54 56 58 60 62 70
c172 58 0 1.48864e-19 $X=4.897 $Y=1.815
c173 45 0 1.8694e-19 $X=5.145 $Y=1.59
c174 31 0 1.545e-19 $X=3.205 $Y=2.365
c175 19 0 5.22007e-20 $X=5.865 $Y=1.45
r176 52 54 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.105 $Y=0.835
+ $X2=3.205 $Y2=0.835
r177 49 70 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=6.245 $Y=1.87
+ $X2=6.365 $Y2=1.87
r178 49 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.245 $Y=1.87
+ $X2=6.155 $Y2=1.87
r179 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.245
+ $Y=1.87 $X2=6.245 $Y2=1.87
r180 46 62 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.76 $Y=1.87
+ $X2=5.76 $Y2=1.59
r181 46 48 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.845 $Y=1.87
+ $X2=6.245 $Y2=1.87
r182 44 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=1.59
+ $X2=5.76 $Y2=1.59
r183 44 45 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.675 $Y=1.59
+ $X2=5.145 $Y2=1.59
r184 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.06 $Y=1.675
+ $X2=5.145 $Y2=1.59
r185 42 58 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.06 $Y=1.675
+ $X2=5.06 $Y2=1.815
r186 40 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.815
+ $Y=1.9 $X2=4.815 $Y2=1.9
r187 40 58 7.55351 $w=4.93e-07 $l=8.5e-08 $layer=LI1_cond $X=4.897 $Y=1.9
+ $X2=4.897 $Y2=1.815
r188 40 41 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.65 $Y=1.9
+ $X2=3.995 $Y2=1.9
r189 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.91 $Y=1.985
+ $X2=3.995 $Y2=1.9
r190 38 39 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.91 $Y=1.985
+ $X2=3.91 $Y2=2.365
r191 37 56 2.28545 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.375 $Y=2.45
+ $X2=3.245 $Y2=2.45
r192 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.825 $Y=2.45
+ $X2=3.91 $Y2=2.365
r193 36 37 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.825 $Y=2.45
+ $X2=3.375 $Y2=2.45
r194 32 56 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=2.535
+ $X2=3.245 $Y2=2.45
r195 32 34 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=3.245 $Y=2.535
+ $X2=3.245 $Y2=2.88
r196 31 56 4.14756 $w=2.2e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.205 $Y=2.365
+ $X2=3.245 $Y2=2.45
r197 30 54 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=1
+ $X2=3.205 $Y2=0.835
r198 30 31 84.1061 $w=1.78e-07 $l=1.365e-06 $layer=LI1_cond $X=3.205 $Y=1
+ $X2=3.205 $Y2=2.365
r199 28 60 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=4.815 $Y=2.25
+ $X2=4.815 $Y2=1.9
r200 28 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=2.25
+ $X2=4.815 $Y2=2.415
r201 26 60 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=4.815 $Y=1.77
+ $X2=4.815 $Y2=1.9
r202 26 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.77
+ $X2=4.815 $Y2=1.605
r203 22 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=2.035
+ $X2=6.365 $Y2=1.87
r204 22 24 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.365 $Y=2.035
+ $X2=6.365 $Y2=2.675
r205 21 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.155 $Y=1.705
+ $X2=6.155 $Y2=1.87
r206 20 21 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.155 $Y=1.525
+ $X2=6.155 $Y2=1.705
r207 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.08 $Y=1.45
+ $X2=6.155 $Y2=1.525
r208 18 19 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.08 $Y=1.45
+ $X2=5.865 $Y2=1.45
r209 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.79 $Y=1.375
+ $X2=5.865 $Y2=1.45
r210 15 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.79 $Y=1.375
+ $X2=5.79 $Y2=0.945
r211 13 27 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.905 $Y=1.055
+ $X2=4.905 $Y2=1.605
r212 9 29 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.725 $Y=2.885 $X2=4.725
+ $Y2=2.415
r213 2 34 600 $w=1.7e-07 $l=2.79106e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=2.675 $X2=3.21 $Y2=2.88
r214 1 52 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.965
+ $Y=0.625 $X2=3.105 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%SET_B 3 5 7 11 13 17 19 21 22 24 28 29 30 32
+ 33 35 38 39 43 49
c120 38 0 5.22007e-20 $X=6.435 $Y=2.347
c121 5 0 2.30611e-19 $X=5.84 $Y=2.425
c122 3 0 7.23512e-20 $X=5.265 $Y=1.055
r123 47 49 0.606549 $w=2.83e-07 $l=1.5e-08 $layer=LI1_cond $X=5.505 $Y=2.347
+ $X2=5.52 $Y2=2.347
r124 39 47 2.87695 $w=2.85e-07 $l=9.5e-08 $layer=LI1_cond $X=5.41 $Y=2.347
+ $X2=5.505 $Y2=2.347
r125 39 49 1.41528 $w=2.83e-07 $l=3.5e-08 $layer=LI1_cond $X=5.555 $Y=2.347
+ $X2=5.52 $Y2=2.347
r126 38 39 35.5842 $w=2.83e-07 $l=8.8e-07 $layer=LI1_cond $X=6.435 $Y=2.347
+ $X2=5.555 $Y2=2.347
r127 36 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.26 $Y=1.93
+ $X2=8.26 $Y2=2.095
r128 36 43 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.26 $Y=1.93 $X2=8.26
+ $Y2=1.84
r129 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.26
+ $Y=1.93 $X2=8.26 $Y2=1.93
r130 33 35 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=7.62 $Y=1.93
+ $X2=8.26 $Y2=1.93
r131 31 33 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.525 $Y=2.095
+ $X2=7.62 $Y2=1.93
r132 31 32 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=7.525 $Y=2.095
+ $X2=7.525 $Y2=2.905
r133 29 32 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.43 $Y=2.99
+ $X2=7.525 $Y2=2.905
r134 29 30 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=7.43 $Y=2.99
+ $X2=6.605 $Y2=2.99
r135 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.52 $Y=2.905
+ $X2=6.605 $Y2=2.99
r136 27 38 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=6.52 $Y=2.49
+ $X2=6.435 $Y2=2.347
r137 27 28 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.52 $Y=2.49
+ $X2=6.52 $Y2=2.905
r138 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.41
+ $Y=2.01 $X2=5.41 $Y2=2.01
r139 22 39 4.30028 $w=1.9e-07 $l=1.42e-07 $layer=LI1_cond $X=5.41 $Y=2.205
+ $X2=5.41 $Y2=2.347
r140 22 24 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=5.41 $Y=2.205
+ $X2=5.41 $Y2=2.01
r141 21 25 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=5.695 $Y=2.01
+ $X2=5.41 $Y2=2.01
r142 19 25 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.34 $Y=2.01 $X2=5.41
+ $Y2=2.01
r143 15 17 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=8.67 $Y=1.765
+ $X2=8.67 $Y2=0.665
r144 14 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.425 $Y=1.84
+ $X2=8.26 $Y2=1.84
r145 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.595 $Y=1.84
+ $X2=8.67 $Y2=1.765
r146 13 14 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=8.595 $Y=1.84
+ $X2=8.425 $Y2=1.84
r147 11 46 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.17 $Y=2.465
+ $X2=8.17 $Y2=2.095
r148 5 21 119.73 $w=1.68e-07 $l=4.32146e-07 $layer=POLY_cond $X=5.84 $Y=2.425
+ $X2=5.805 $Y2=2.01
r149 5 7 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=5.84 $Y=2.425
+ $X2=5.84 $Y2=2.885
r150 1 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.265 $Y=1.845
+ $X2=5.34 $Y2=2.01
r151 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.265 $Y=1.845
+ $X2=5.265 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_191_21# 1 2 8 9 11 12 15 19 21 25 27 29 31
+ 39 42 49
c131 42 0 1.23604e-19 $X=1.612 $Y=2.475
c132 25 0 1.54738e-19 $X=7.265 $Y=0.895
r133 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.38
+ $Y=1.89 $X2=1.38 $Y2=1.89
r134 37 42 15.1358 $w=1.68e-07 $l=2.32e-07 $layer=LI1_cond $X=1.38 $Y=2.39
+ $X2=1.612 $Y2=2.39
r135 37 39 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.38 $Y=2.305
+ $X2=1.38 $Y2=1.89
r136 32 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=0.35
+ $X2=1.12 $Y2=0.515
r137 32 49 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.12 $Y=0.35
+ $X2=1.12 $Y2=0.18
r138 31 35 8.04086 $w=5.93e-07 $l=4e-07 $layer=LI1_cond $X=1.252 $Y=0.35
+ $X2=1.252 $Y2=0.75
r139 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=0.35 $X2=1.12 $Y2=0.35
r140 25 27 805.043 $w=1.5e-07 $l=1.57e-06 $layer=POLY_cond $X=7.265 $Y=0.895
+ $X2=7.265 $Y2=2.465
r141 23 25 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.265 $Y=0.255
+ $X2=7.265 $Y2=0.895
r142 22 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.395 $Y=0.18
+ $X2=3.32 $Y2=0.18
r143 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.19 $Y=0.18
+ $X2=7.265 $Y2=0.255
r144 21 22 1945.95 $w=1.5e-07 $l=3.795e-06 $layer=POLY_cond $X=7.19 $Y=0.18
+ $X2=3.395 $Y2=0.18
r145 17 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.32 $Y=0.255
+ $X2=3.32 $Y2=0.18
r146 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.32 $Y=0.255
+ $X2=3.32 $Y2=0.835
r147 13 15 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.96 $Y=1.975
+ $X2=2.96 $Y2=2.885
r148 12 40 39.2615 $w=2.56e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.545 $Y=1.9
+ $X2=1.38 $Y2=1.89
r149 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.885 $Y=1.9
+ $X2=2.96 $Y2=1.975
r150 11 12 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=2.885 $Y=1.9
+ $X2=1.545 $Y2=1.9
r151 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=0.18
+ $X2=1.12 $Y2=0.18
r152 9 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.245 $Y=0.18
+ $X2=3.32 $Y2=0.18
r153 9 10 1005.02 $w=1.5e-07 $l=1.96e-06 $layer=POLY_cond $X=3.245 $Y=0.18
+ $X2=1.285 $Y2=0.18
r154 8 40 60.25 $w=2.56e-07 $l=3.93954e-07 $layer=POLY_cond $X=1.06 $Y=1.725
+ $X2=1.38 $Y2=1.89
r155 8 52 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=1.06 $Y=1.725
+ $X2=1.06 $Y2=0.515
r156 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.52
+ $Y=2.325 $X2=1.645 $Y2=2.47
r157 1 35 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.24
+ $Y=0.625 $X2=1.385 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_1533_258# 1 2 9 11 12 15 16 19 21 23 26 27
+ 33 39
r85 35 36 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=9.405 $Y=1.11 $X2=9.405
+ $Y2=1.15
r86 33 35 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=9.405 $Y=0.865
+ $X2=9.405 $Y2=1.11
r87 27 30 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=9.365 $Y=1.9
+ $X2=9.365 $Y2=2.045
r88 25 26 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=9.92 $Y=1.235
+ $X2=9.92 $Y2=1.815
r89 24 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.57 $Y=1.15
+ $X2=9.405 $Y2=1.15
r90 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.835 $Y=1.15
+ $X2=9.92 $Y2=1.235
r91 23 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.835 $Y=1.15
+ $X2=9.57 $Y2=1.15
r92 22 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.53 $Y=1.9
+ $X2=9.365 $Y2=1.9
r93 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.835 $Y=1.9
+ $X2=9.92 $Y2=1.815
r94 21 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.835 $Y=1.9
+ $X2=9.53 $Y2=1.9
r95 19 40 34.4622 $w=3.6e-07 $l=2.15e-07 $layer=POLY_cond $X=8.205 $Y=1.15
+ $X2=8.205 $Y2=1.365
r96 19 39 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=8.205 $Y=1.15
+ $X2=8.205 $Y2=0.985
r97 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.19
+ $Y=1.15 $X2=8.19 $Y2=1.15
r98 16 35 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.24 $Y=1.11
+ $X2=9.405 $Y2=1.11
r99 16 18 48.4026 $w=2.48e-07 $l=1.05e-06 $layer=LI1_cond $X=9.24 $Y=1.11
+ $X2=8.19 $Y2=1.11
r100 15 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.31 $Y=0.665
+ $X2=8.31 $Y2=0.985
r101 11 40 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.025 $Y=1.365
+ $X2=8.205 $Y2=1.365
r102 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.025 $Y=1.365
+ $X2=7.815 $Y2=1.365
r103 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.74 $Y=1.44
+ $X2=7.815 $Y2=1.365
r104 7 9 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=7.74 $Y=1.44
+ $X2=7.74 $Y2=2.465
r105 2 30 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=9.24
+ $Y=1.835 $X2=9.365 $Y2=2.045
r106 1 33 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.28
+ $Y=0.655 $X2=9.405 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_1360_451# 1 2 3 10 12 16 18 22 26 28 32 36
+ 38 42 46 48 49 50 52 54 55 58 61 67 72 74 78 80
r156 76 78 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=8.385 $Y=2.44
+ $X2=8.61 $Y2=2.44
r157 70 72 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7 $Y=1.075 $X2=7.165
+ $Y2=1.075
r158 65 67 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=6.95 $Y=2.57
+ $X2=7.165 $Y2=2.57
r159 62 81 12.4655 $w=3.48e-07 $l=9e-08 $layer=POLY_cond $X=9.51 $Y=1.5 $X2=9.51
+ $Y2=1.41
r160 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.49
+ $Y=1.5 $X2=9.49 $Y2=1.5
r161 59 80 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.695 $Y=1.525
+ $X2=8.61 $Y2=1.525
r162 59 61 38.1747 $w=2.38e-07 $l=7.95e-07 $layer=LI1_cond $X=8.695 $Y=1.525
+ $X2=9.49 $Y2=1.525
r163 58 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.61 $Y=2.275
+ $X2=8.61 $Y2=2.44
r164 57 80 2.11342 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=8.61 $Y=1.645
+ $X2=8.61 $Y2=1.525
r165 57 58 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=8.61 $Y=1.645
+ $X2=8.61 $Y2=2.275
r166 56 74 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.25 $Y=1.495
+ $X2=7.165 $Y2=1.495
r167 55 80 4.3182 $w=2.1e-07 $l=9.88686e-08 $layer=LI1_cond $X=8.525 $Y=1.495
+ $X2=8.61 $Y2=1.525
r168 55 56 78.5606 $w=1.78e-07 $l=1.275e-06 $layer=LI1_cond $X=8.525 $Y=1.495
+ $X2=7.25 $Y2=1.495
r169 54 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=2.405
+ $X2=7.165 $Y2=2.57
r170 53 74 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.165 $Y=1.585
+ $X2=7.165 $Y2=1.495
r171 53 54 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=7.165 $Y=1.585
+ $X2=7.165 $Y2=2.405
r172 52 74 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.165 $Y=1.405
+ $X2=7.165 $Y2=1.495
r173 51 72 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.165 $Y=1.175
+ $X2=7.165 $Y2=1.075
r174 51 52 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.165 $Y=1.175
+ $X2=7.165 $Y2=1.405
r175 44 50 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=11.1 $Y=1.335
+ $X2=11.08 $Y2=1.41
r176 44 46 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=11.1 $Y=1.335 $X2=11.1
+ $Y2=0.865
r177 40 50 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=11.06 $Y=1.485
+ $X2=11.08 $Y2=1.41
r178 40 42 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=11.06 $Y=1.485
+ $X2=11.06 $Y2=2.155
r179 39 49 12.05 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=10.65 $Y=1.41
+ $X2=10.555 $Y2=1.41
r180 38 50 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=11.08 $Y2=1.41
r181 38 39 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=10.65 $Y2=1.41
r182 34 49 12.05 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=10.575 $Y=1.335
+ $X2=10.555 $Y2=1.41
r183 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.575 $Y=1.335
+ $X2=10.575 $Y2=0.655
r184 30 49 12.05 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=10.535 $Y=1.485
+ $X2=10.555 $Y2=1.41
r185 30 32 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=10.535 $Y=1.485
+ $X2=10.535 $Y2=2.465
r186 29 48 12.05 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=10.22 $Y=1.41
+ $X2=10.125 $Y2=1.41
r187 28 49 12.05 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=10.46 $Y=1.41
+ $X2=10.555 $Y2=1.41
r188 28 29 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.46 $Y=1.41
+ $X2=10.22 $Y2=1.41
r189 24 48 12.05 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=10.145 $Y=1.335
+ $X2=10.125 $Y2=1.41
r190 24 26 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.145 $Y=1.335
+ $X2=10.145 $Y2=0.655
r191 20 48 12.05 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=10.105 $Y=1.485
+ $X2=10.125 $Y2=1.41
r192 20 22 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=10.105 $Y=1.485
+ $X2=10.105 $Y2=2.465
r193 19 81 22.4912 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=9.695 $Y=1.41
+ $X2=9.51 $Y2=1.41
r194 18 48 12.05 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=10.03 $Y=1.41
+ $X2=10.125 $Y2=1.41
r195 18 19 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.03 $Y=1.41
+ $X2=9.695 $Y2=1.41
r196 14 81 26.2957 $w=3.48e-07 $l=1.42653e-07 $layer=POLY_cond $X=9.62 $Y=1.335
+ $X2=9.51 $Y2=1.41
r197 14 16 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=9.62 $Y=1.335 $X2=9.62
+ $Y2=0.865
r198 10 62 38.7612 $w=3.48e-07 $l=1.96914e-07 $layer=POLY_cond $X=9.58 $Y=1.665
+ $X2=9.51 $Y2=1.5
r199 10 12 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.58 $Y=1.665
+ $X2=9.58 $Y2=2.045
r200 3 76 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=2.255 $X2=8.385 $Y2=2.44
r201 2 65 600 $w=1.7e-07 $l=3.82721e-07 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=2.255 $X2=6.95 $Y2=2.57
r202 1 70 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=6.815
+ $Y=0.795 $X2=7 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_2227_367# 1 2 9 12 14 16 18 21 23 26 30 34
+ 37 38 39
r53 38 39 33.1619 $w=4e-07 $l=7.5e-08 $layer=POLY_cond $X=11.925 $Y=1.42
+ $X2=11.925 $Y2=1.345
r54 35 41 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=11.925 $Y=1.51
+ $X2=11.925 $Y2=1.675
r55 35 38 12.5135 $w=4e-07 $l=9e-08 $layer=POLY_cond $X=11.925 $Y=1.51
+ $X2=11.925 $Y2=1.42
r56 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.89
+ $Y=1.51 $X2=11.89 $Y2=1.51
r57 32 37 1.25991 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=11.48 $Y=1.51
+ $X2=11.315 $Y2=1.51
r58 32 34 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=11.48 $Y=1.51
+ $X2=11.89 $Y2=1.51
r59 28 37 5.2656 $w=3.22e-07 $l=1.68953e-07 $layer=LI1_cond $X=11.307 $Y=1.675
+ $X2=11.315 $Y2=1.51
r60 28 30 11.1586 $w=3.13e-07 $l=3.05e-07 $layer=LI1_cond $X=11.307 $Y=1.675
+ $X2=11.307 $Y2=1.98
r61 24 37 5.2656 $w=3.22e-07 $l=1.65e-07 $layer=LI1_cond $X=11.315 $Y=1.345
+ $X2=11.315 $Y2=1.51
r62 24 26 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=11.315 $Y=1.345
+ $X2=11.315 $Y2=0.865
r63 19 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.48 $Y=1.495
+ $X2=12.48 $Y2=1.42
r64 19 21 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=12.48 $Y=1.495
+ $X2=12.48 $Y2=2.465
r65 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.48 $Y=1.345
+ $X2=12.48 $Y2=1.42
r66 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=12.48 $Y=1.345
+ $X2=12.48 $Y2=0.815
r67 15 38 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=12.125 $Y=1.42
+ $X2=11.925 $Y2=1.42
r68 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.405 $Y=1.42
+ $X2=12.48 $Y2=1.42
r69 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.405 $Y=1.42
+ $X2=12.125 $Y2=1.42
r70 12 41 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=12.05 $Y=2.465
+ $X2=12.05 $Y2=1.675
r71 9 39 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=12.05 $Y=0.815
+ $X2=12.05 $Y2=1.345
r72 2 30 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=11.135
+ $Y=1.835 $X2=11.275 $Y2=1.98
r73 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.175
+ $Y=0.655 $X2=11.315 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 52
+ 58 62 64 68 70 86 91 99 107 112 117 126 130 134 136 139 142 145 148 152
c154 34 0 1.10806e-19 $X=2.195 $Y=2.82
r155 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r156 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r157 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r158 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r159 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r160 136 137 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r161 132 134 8.99479 $w=5.78e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=3.125
+ $X2=4.675 $Y2=3.125
r162 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r163 129 132 1.0311 $w=5.78e-07 $l=5e-08 $layer=LI1_cond $X=4.51 $Y=3.125
+ $X2=4.56 $Y2=3.125
r164 129 130 20.44 $w=5.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.51 $Y=3.125
+ $X2=3.84 $Y2=3.125
r165 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r166 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r167 121 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r168 121 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r169 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r170 118 148 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=11.975 $Y=3.33
+ $X2=11.822 $Y2=3.33
r171 118 120 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.975 $Y=3.33
+ $X2=12.24 $Y2=3.33
r172 117 151 4.48816 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=12.56 $Y=3.33
+ $X2=12.76 $Y2=3.33
r173 117 120 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.56 $Y=3.33
+ $X2=12.24 $Y2=3.33
r174 116 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r175 116 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r176 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r177 113 145 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=10.98 $Y=3.33
+ $X2=10.812 $Y2=3.33
r178 113 115 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.98 $Y=3.33
+ $X2=11.28 $Y2=3.33
r179 112 148 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=11.67 $Y=3.33
+ $X2=11.822 $Y2=3.33
r180 112 115 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.67 $Y=3.33
+ $X2=11.28 $Y2=3.33
r181 111 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r182 111 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r183 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r184 108 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.055 $Y=3.33
+ $X2=9.89 $Y2=3.33
r185 108 110 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.055 $Y=3.33
+ $X2=10.32 $Y2=3.33
r186 107 145 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=10.645 $Y=3.33
+ $X2=10.812 $Y2=3.33
r187 107 110 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.645 $Y=3.33
+ $X2=10.32 $Y2=3.33
r188 106 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r189 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r190 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r191 103 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r192 102 105 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r193 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 100 139 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=7.937 $Y2=3.33
r195 100 102 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=8.4 $Y2=3.33
r196 99 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.725 $Y=3.33
+ $X2=9.89 $Y2=3.33
r197 99 105 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.725 $Y=3.33
+ $X2=9.36 $Y2=3.33
r198 98 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r199 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r200 94 97 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r201 92 136 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6.125 $Y2=3.33
r202 92 94 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6.48 $Y2=3.33
r203 91 139 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.79 $Y=3.33
+ $X2=7.937 $Y2=3.33
r204 91 97 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.79 $Y=3.33
+ $X2=7.44 $Y2=3.33
r205 90 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r206 90 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r207 89 134 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=4.675 $Y2=3.33
r208 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r209 86 136 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.985 $Y=3.33
+ $X2=6.125 $Y2=3.33
r210 86 89 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=5.985 $Y=3.33
+ $X2=5.04 $Y2=3.33
r211 85 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r212 84 130 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=3.84 $Y2=3.33
r213 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r214 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r215 82 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r216 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r217 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r218 79 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.195 $Y2=3.33
r219 79 81 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r220 77 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r221 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r222 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r223 74 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r224 73 76 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r226 71 123 4.5891 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=0.52 $Y=3.33
+ $X2=0.26 $Y2=3.33
r227 71 73 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.52 $Y=3.33 $X2=0.72
+ $Y2=3.33
r228 70 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=3.33
+ $X2=2.195 $Y2=3.33
r229 70 76 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=3.33
+ $X2=1.68 $Y2=3.33
r230 68 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r231 68 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r232 68 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r233 64 67 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=12.71 $Y=1.98
+ $X2=12.71 $Y2=2.95
r234 62 151 3.02951 $w=3e-07 $l=1.07121e-07 $layer=LI1_cond $X=12.71 $Y=3.245
+ $X2=12.76 $Y2=3.33
r235 62 67 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=12.71 $Y=3.245
+ $X2=12.71 $Y2=2.95
r236 58 61 35.5179 $w=3.03e-07 $l=9.4e-07 $layer=LI1_cond $X=11.822 $Y=2.01
+ $X2=11.822 $Y2=2.95
r237 56 148 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.822 $Y=3.245
+ $X2=11.822 $Y2=3.33
r238 56 61 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=11.822 $Y=3.245
+ $X2=11.822 $Y2=2.95
r239 52 55 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=10.812 $Y=1.98
+ $X2=10.812 $Y2=2.46
r240 50 145 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=10.812 $Y=3.245
+ $X2=10.812 $Y2=3.33
r241 50 55 27.005 $w=3.33e-07 $l=7.85e-07 $layer=LI1_cond $X=10.812 $Y=3.245
+ $X2=10.812 $Y2=2.46
r242 46 49 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.89 $Y=2.24
+ $X2=9.89 $Y2=2.95
r243 44 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.89 $Y=3.245
+ $X2=9.89 $Y2=3.33
r244 44 49 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.89 $Y=3.245
+ $X2=9.89 $Y2=2.95
r245 40 139 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.937 $Y=3.245
+ $X2=7.937 $Y2=3.33
r246 40 42 31.448 $w=2.93e-07 $l=8.05e-07 $layer=LI1_cond $X=7.937 $Y=3.245
+ $X2=7.937 $Y2=2.44
r247 36 136 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=3.245
+ $X2=6.125 $Y2=3.33
r248 36 38 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=6.125 $Y=3.245
+ $X2=6.125 $Y2=2.825
r249 32 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=3.245
+ $X2=2.195 $Y2=3.33
r250 32 34 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.195 $Y=3.245
+ $X2=2.195 $Y2=2.82
r251 28 123 3.17707 $w=3.3e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.355 $Y=3.245
+ $X2=0.26 $Y2=3.33
r252 28 30 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=0.355 $Y=3.245
+ $X2=0.355 $Y2=2.41
r253 9 67 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=12.555
+ $Y=1.835 $X2=12.695 $Y2=2.95
r254 9 64 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.555
+ $Y=1.835 $X2=12.695 $Y2=1.98
r255 8 61 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=11.71
+ $Y=1.835 $X2=11.835 $Y2=2.95
r256 8 58 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=11.71
+ $Y=1.835 $X2=11.835 $Y2=2.01
r257 7 55 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=10.61
+ $Y=1.835 $X2=10.75 $Y2=2.46
r258 7 52 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=10.61
+ $Y=1.835 $X2=10.845 $Y2=1.98
r259 6 49 400 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=9.655
+ $Y=1.835 $X2=9.89 $Y2=2.95
r260 6 46 400 $w=1.7e-07 $l=5.09117e-07 $layer=licon1_PDIFF $count=1 $X=9.655
+ $Y=1.835 $X2=9.89 $Y2=2.24
r261 5 42 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=7.815
+ $Y=2.255 $X2=7.955 $Y2=2.44
r262 4 38 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=5.915
+ $Y=2.675 $X2=6.15 $Y2=2.825
r263 3 129 300 $w=1.7e-07 $l=7.68228e-07 $layer=licon1_PDIFF $count=2 $X=3.865
+ $Y=2.675 $X2=4.51 $Y2=2.945
r264 2 34 600 $w=1.7e-07 $l=6.11331e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=2.325 $X2=2.195 $Y2=2.82
r265 1 30 600 $w=1.7e-07 $l=4.93559e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.975 $X2=0.355 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_507_125# 1 2 9 12 15 20
c34 9 0 5.68328e-20 $X=2.675 $Y=0.835
r35 18 20 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.745 $Y=2.86
+ $X2=2.855 $Y2=2.86
r36 12 20 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=2.695
+ $X2=2.855 $Y2=2.86
r37 11 15 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=1.435
+ $X2=2.855 $Y2=1.35
r38 11 12 77.6364 $w=1.78e-07 $l=1.26e-06 $layer=LI1_cond $X=2.855 $Y=1.435
+ $X2=2.855 $Y2=2.695
r39 7 15 10.308 $w=1.68e-07 $l=1.58e-07 $layer=LI1_cond $X=2.697 $Y=1.35
+ $X2=2.855 $Y2=1.35
r40 7 9 21.0873 $w=2.33e-07 $l=4.3e-07 $layer=LI1_cond $X=2.697 $Y=1.265
+ $X2=2.697 $Y2=0.835
r41 2 18 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=2.605
+ $Y=2.675 $X2=2.745 $Y2=2.86
r42 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.625 $X2=2.675 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%Q_N 1 2 7 8 9 10 11 12 13 22
r20 13 40 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=10.345 $Y=2.775
+ $X2=10.345 $Y2=2.91
r21 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=2.405
+ $X2=10.345 $Y2=2.775
r22 11 12 18.7272 $w=2.38e-07 $l=3.9e-07 $layer=LI1_cond $X=10.345 $Y=2.015
+ $X2=10.345 $Y2=2.405
r23 10 11 16.8065 $w=2.38e-07 $l=3.5e-07 $layer=LI1_cond $X=10.345 $Y=1.665
+ $X2=10.345 $Y2=2.015
r24 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=1.295
+ $X2=10.345 $Y2=1.665
r25 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=0.925
+ $X2=10.345 $Y2=1.295
r26 7 8 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=0.555
+ $X2=10.345 $Y2=0.925
r27 7 22 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=10.345 $Y=0.555
+ $X2=10.345 $Y2=0.42
r28 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.18
+ $Y=1.835 $X2=10.32 $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=10.18
+ $Y=1.835 $X2=10.32 $Y2=2.015
r30 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=10.22
+ $Y=0.235 $X2=10.36 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%Q 1 2 7 10
r17 15 17 44.6866 $w=2.43e-07 $l=9.5e-07 $layer=LI1_cond $X=12.267 $Y=1.96
+ $X2=12.267 $Y2=2.91
r18 7 15 31.2806 $w=2.43e-07 $l=6.65e-07 $layer=LI1_cond $X=12.267 $Y=1.295
+ $X2=12.267 $Y2=1.96
r19 7 10 35.5141 $w=2.43e-07 $l=7.55e-07 $layer=LI1_cond $X=12.267 $Y=1.295
+ $X2=12.267 $Y2=0.54
r20 2 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=12.125
+ $Y=1.835 $X2=12.265 $Y2=2.91
r21 2 15 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=12.125
+ $Y=1.835 $X2=12.265 $Y2=1.96
r22 1 10 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.125
+ $Y=0.395 $X2=12.265 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 48
+ 52 56 62 64 66 69 70 72 73 74 89 96 104 109 114 123 126 129 132 135 139
r146 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r147 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r148 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r149 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r150 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.84 $Y2=0
r151 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r152 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r153 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r154 118 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r155 118 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r156 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r157 115 135 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=11.975 $Y=0
+ $X2=11.822 $Y2=0
r158 115 117 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.975 $Y=0
+ $X2=12.24 $Y2=0
r159 114 138 4.48816 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=12.56 $Y=0 $X2=12.76
+ $Y2=0
r160 114 117 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.56 $Y=0
+ $X2=12.24 $Y2=0
r161 113 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r162 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r163 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r164 110 132 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=10.98 $Y=0
+ $X2=10.807 $Y2=0
r165 110 112 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.98 $Y=0
+ $X2=11.28 $Y2=0
r166 109 135 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=11.67 $Y=0
+ $X2=11.822 $Y2=0
r167 109 112 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.67 $Y=0
+ $X2=11.28 $Y2=0
r168 108 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r169 108 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r170 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r171 105 129 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.055 $Y=0
+ $X2=9.91 $Y2=0
r172 105 107 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.055 $Y=0
+ $X2=10.32 $Y2=0
r173 104 132 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.807 $Y2=0
r174 104 107 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.32 $Y2=0
r175 103 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r176 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r177 100 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r178 99 102 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.4
+ $Y2=0
r179 99 100 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r180 97 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.74 $Y=0
+ $X2=5.575 $Y2=0
r181 97 99 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.74 $Y=0 $X2=6
+ $Y2=0
r182 96 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.72 $Y=0
+ $X2=8.885 $Y2=0
r183 96 102 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.72 $Y=0 $X2=8.4
+ $Y2=0
r184 95 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r185 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r186 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r187 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r188 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r189 89 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.41 $Y=0
+ $X2=5.575 $Y2=0
r190 89 94 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.04
+ $Y2=0
r191 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r192 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r193 85 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r194 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r195 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r196 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r197 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r198 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r199 79 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r200 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r201 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r202 76 120 4.05675 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=0
+ $X2=0.225 $Y2=0
r203 76 78 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.72
+ $Y2=0
r204 74 103 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=8.4 $Y2=0
r205 74 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r206 72 87 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.6
+ $Y2=0
r207 72 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.945
+ $Y2=0
r208 71 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.075 $Y=0 $X2=4.08
+ $Y2=0
r209 71 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.075 $Y=0 $X2=3.945
+ $Y2=0
r210 69 81 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.68
+ $Y2=0
r211 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.895
+ $Y2=0
r212 68 84 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=2.16
+ $Y2=0
r213 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=1.895
+ $Y2=0
r214 64 138 3.02951 $w=3e-07 $l=1.07121e-07 $layer=LI1_cond $X=12.71 $Y=0.085
+ $X2=12.76 $Y2=0
r215 64 66 17.4787 $w=2.98e-07 $l=4.55e-07 $layer=LI1_cond $X=12.71 $Y=0.085
+ $X2=12.71 $Y2=0.54
r216 60 135 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.822 $Y=0.085
+ $X2=11.822 $Y2=0
r217 60 62 17.1922 $w=3.03e-07 $l=4.55e-07 $layer=LI1_cond $X=11.822 $Y=0.085
+ $X2=11.822 $Y2=0.54
r218 56 58 18.3723 $w=3.43e-07 $l=5.5e-07 $layer=LI1_cond $X=10.807 $Y=0.38
+ $X2=10.807 $Y2=0.93
r219 54 132 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.807 $Y=0.085
+ $X2=10.807 $Y2=0
r220 54 56 9.85422 $w=3.43e-07 $l=2.95e-07 $layer=LI1_cond $X=10.807 $Y=0.085
+ $X2=10.807 $Y2=0.38
r221 50 129 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.91 $Y=0.085
+ $X2=9.91 $Y2=0
r222 50 52 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=9.91 $Y=0.085
+ $X2=9.91 $Y2=0.38
r223 49 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.05 $Y=0
+ $X2=8.885 $Y2=0
r224 48 129 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.765 $Y=0
+ $X2=9.91 $Y2=0
r225 48 49 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.765 $Y=0
+ $X2=9.05 $Y2=0
r226 44 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=0.085
+ $X2=8.885 $Y2=0
r227 44 46 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=8.885 $Y=0.085
+ $X2=8.885 $Y2=0.665
r228 40 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0
r229 40 42 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0.87
r230 36 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=3.945 $Y2=0
r231 36 38 31.2489 $w=2.58e-07 $l=7.05e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=3.945 $Y2=0.79
r232 32 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.085
+ $X2=1.895 $Y2=0
r233 32 34 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.895 $Y=0.085
+ $X2=1.895 $Y2=0.75
r234 28 120 3.19131 $w=2.65e-07 $l=1.27609e-07 $layer=LI1_cond $X=0.317 $Y=0.085
+ $X2=0.225 $Y2=0
r235 28 30 44.3582 $w=2.63e-07 $l=1.02e-06 $layer=LI1_cond $X=0.317 $Y=0.085
+ $X2=0.317 $Y2=1.105
r236 9 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.555
+ $Y=0.395 $X2=12.695 $Y2=0.54
r237 8 62 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=11.71
+ $Y=0.395 $X2=11.835 $Y2=0.54
r238 7 58 182 $w=1.7e-07 $l=8.03959e-07 $layer=licon1_NDIFF $count=1 $X=10.65
+ $Y=0.235 $X2=10.885 $Y2=0.93
r239 7 56 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=10.65
+ $Y=0.235 $X2=10.79 $Y2=0.38
r240 6 52 91 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=2 $X=9.695
+ $Y=0.655 $X2=9.93 $Y2=0.38
r241 5 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.745
+ $Y=0.455 $X2=8.885 $Y2=0.665
r242 4 42 182 $w=1.7e-07 $l=2.47184e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.845 $X2=5.575 $Y2=0.87
r243 3 38 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=3.755
+ $Y=0.625 $X2=3.9 $Y2=0.79
r244 2 34 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.625 $X2=1.895 $Y2=0.75
r245 1 30 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.895 $X2=0.35 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_1173_125# 1 2 9 11 13
r27 11 13 77.9136 $w=1.98e-07 $l=1.405e-06 $layer=LI1_cond $X=6.17 $Y=0.365
+ $X2=7.575 $Y2=0.365
r28 7 11 6.96842 $w=2e-07 $l=1.72916e-07 $layer=LI1_cond $X=6.04 $Y=0.465
+ $X2=6.17 $Y2=0.365
r29 7 9 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=6.04 $Y=0.465
+ $X2=6.04 $Y2=0.83
r30 2 13 182 $w=1.7e-07 $l=3.21559e-07 $layer=licon1_NDIFF $count=1 $X=7.34
+ $Y=0.575 $X2=7.575 $Y2=0.37
r31 1 9 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.865
+ $Y=0.625 $X2=6.005 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_2%A_1280_159# 1 2 9 12 14 15
c31 15 0 8.27457e-20 $X=7.93 $Y=0.652
r32 14 15 8.47458 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=0.652
+ $X2=7.93 $Y2=0.652
r33 12 15 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=6.665 $Y=0.72
+ $X2=7.93 $Y2=0.72
r34 7 12 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.515 $Y=0.805
+ $X2=6.665 $Y2=0.72
r35 7 9 7.68295 $w=2.98e-07 $l=2e-07 $layer=LI1_cond $X=6.515 $Y=0.805 $X2=6.515
+ $Y2=1.005
r36 2 14 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=7.97
+ $Y=0.455 $X2=8.095 $Y2=0.665
r37 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.4
+ $Y=0.795 $X2=6.525 $Y2=1.005
.ends

