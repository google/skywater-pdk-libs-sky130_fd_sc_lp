* File: sky130_fd_sc_lp__dfstp_1.spice
* Created: Wed Sep  2 09:44:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfstp_1.pex.spice"
.subckt sky130_fd_sc_lp__dfstp_1  VNB VPB CLK D SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_CLK_M1017_g N_A_33_463#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1018 N_A_202_463#_M1018_d N_A_33_463#_M1018_g N_VGND_M1017_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_400_119#_M1005_d N_D_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1028 N_A_486_119#_M1028_d N_A_33_463#_M1028_g N_A_400_119#_M1005_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1030 A_572_119# N_A_202_463#_M1030_g N_A_486_119#_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_614_93#_M1022_g A_572_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1687 AS=0.0441 PD=1.7 PS=0.63 NRD=28.56 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1027 A_853_47# N_A_486_119#_M1027_g N_A_614_93#_M1027_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_SET_B_M1016_g A_853_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.159917 AS=0.0441 PD=1.12132 PS=0.63 NRD=142.848 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1029 A_1110_47# N_A_486_119#_M1029_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.243683 PD=0.85 PS=1.70868 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1031 N_A_1175_417#_M1031_d N_A_202_463#_M1031_g A_1110_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=5.148 NRS=9.372 M=1
+ R=4.26667 SA=75001.4 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1014 A_1287_91# N_A_33_463#_M1014_g N_A_1175_417#_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0855057 PD=0.63 PS=0.80434 NRD=14.28 NRS=19.992 M=1
+ R=2.8 SA=75001.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1015 A_1359_91# N_A_1329_65#_M1015_g A_1287_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_SET_B_M1008_g A_1359_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0441 PD=0.78 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_A_1329_65#_M1019_d N_A_1175_417#_M1019_g N_VGND_M1008_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=5.712 NRS=22.848 M=1
+ R=2.8 SA=75003 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_1175_417#_M1011_g N_A_1832_131#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0875 AS=0.1113 PD=0.8 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_Q_M1000_d N_A_1832_131#_M1000_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.175 PD=2.21 PS=1.6 NRD=0 NRS=4.284 M=1 R=5.6 SA=75000.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_33_463#_M1012_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1024 N_A_202_463#_M1024_d N_A_33_463#_M1024_g N_VPWR_M1012_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_400_119#_M1009_d N_D_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.1
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_486_119#_M1001_d N_A_202_463#_M1001_g N_A_400_119#_M1009_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1020 A_582_463# N_A_33_463#_M1020_g N_A_486_119#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_614_93#_M1023_g A_582_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75001.4
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_614_93#_M1003_d N_A_486_119#_M1003_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=28.1316 M=1 R=2.8
+ SA=75001.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_SET_B_M1025_g N_A_614_93#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.112 AS=0.0588 PD=0.916667 PS=0.7 NRD=60.9715 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1007 N_A_985_379#_M1007_d N_A_486_119#_M1007_g N_VPWR_M1025_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.224 PD=2.21 PS=1.83333 NRD=0 NRS=29.8849 M=1
+ R=5.6 SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_A_1175_417#_M1013_d N_A_202_463#_M1013_g N_A_1092_417#_M1013_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=32.8202 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_985_379#_M1004_d N_A_33_463#_M1004_g N_A_1175_417#_M1013_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.3399 AS=0.1792 PD=2.7 PS=1.62 NRD=23.443 NRS=5.8509
+ M=1 R=5.6 SA=75000.5 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_1329_65#_M1002_g N_A_1092_417#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_A_1175_417#_M1021_d N_SET_B_M1021_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_1329_65#_M1010_d N_A_1175_417#_M1010_g N_VPWR_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_VPWR_M1026_d N_A_1175_417#_M1026_g N_A_1832_131#_M1026_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.14912 AS=0.1696 PD=1.14189 PS=1.81 NRD=33.8446 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1006 N_Q_M1006_d N_A_1832_131#_M1006_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.29358 PD=3.05 PS=2.24811 NRD=0 NRS=4.9447 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.6423 P=26.07
c_110 VNB 0 1.94585e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfstp_1.pxi.spice"
*
.ends
*
*
