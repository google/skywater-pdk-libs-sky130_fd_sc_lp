* File: sky130_fd_sc_lp__o22ai_4.pxi.spice
* Created: Wed Sep  2 10:20:50 2020
* 
x_PM_SKY130_FD_SC_LP__O22AI_4%A1 N_A1_M1001_g N_A1_M1002_g N_A1_M1006_g
+ N_A1_M1005_g N_A1_M1016_g N_A1_M1012_g N_A1_M1017_g N_A1_M1025_g N_A1_c_124_n
+ N_A1_c_125_n N_A1_c_126_n N_A1_c_127_n N_A1_c_128_n N_A1_c_140_p A1 A1 A1 A1
+ A1 N_A1_c_130_n PM_SKY130_FD_SC_LP__O22AI_4%A1
x_PM_SKY130_FD_SC_LP__O22AI_4%A2 N_A2_M1011_g N_A2_M1003_g N_A2_M1014_g
+ N_A2_M1010_g N_A2_M1023_g N_A2_M1019_g N_A2_M1026_g N_A2_M1022_g A2 A2 A2
+ N_A2_c_254_n PM_SKY130_FD_SC_LP__O22AI_4%A2
x_PM_SKY130_FD_SC_LP__O22AI_4%B1 N_B1_M1007_g N_B1_M1000_g N_B1_M1015_g
+ N_B1_M1009_g N_B1_M1024_g N_B1_M1020_g N_B1_M1027_g N_B1_M1029_g N_B1_c_341_n
+ N_B1_c_342_n N_B1_c_343_n B1 B1 B1 N_B1_c_344_n N_B1_c_345_n N_B1_c_346_n
+ N_B1_c_347_n B1 N_B1_c_348_n PM_SKY130_FD_SC_LP__O22AI_4%B1
x_PM_SKY130_FD_SC_LP__O22AI_4%B2 N_B2_M1008_g N_B2_M1004_g N_B2_M1018_g
+ N_B2_M1013_g N_B2_M1030_g N_B2_M1021_g N_B2_M1031_g N_B2_M1028_g N_B2_c_482_n
+ B2 N_B2_c_472_n N_B2_c_467_n PM_SKY130_FD_SC_LP__O22AI_4%B2
x_PM_SKY130_FD_SC_LP__O22AI_4%VPWR N_VPWR_M1002_s N_VPWR_M1005_s N_VPWR_M1025_s
+ N_VPWR_M1009_s N_VPWR_M1029_s N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n
+ N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n
+ N_VPWR_c_556_n N_VPWR_c_557_n VPWR N_VPWR_c_558_n N_VPWR_c_559_n
+ N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_547_n PM_SKY130_FD_SC_LP__O22AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O22AI_4%A_119_367# N_A_119_367#_M1002_d
+ N_A_119_367#_M1012_d N_A_119_367#_M1010_s N_A_119_367#_M1022_s
+ N_A_119_367#_c_655_n N_A_119_367#_c_665_n N_A_119_367#_c_670_n
+ N_A_119_367#_c_684_n N_A_119_367#_c_671_n N_A_119_367#_c_688_n
+ PM_SKY130_FD_SC_LP__O22AI_4%A_119_367#
x_PM_SKY130_FD_SC_LP__O22AI_4%Y N_Y_M1007_s N_Y_M1024_s N_Y_M1018_d N_Y_M1031_d
+ N_Y_M1003_d N_Y_M1019_d N_Y_M1004_d N_Y_M1021_d N_Y_c_706_n N_Y_c_709_n
+ N_Y_c_698_n N_Y_c_699_n N_Y_c_696_n N_Y_c_700_n N_Y_c_774_n N_Y_c_777_n
+ N_Y_c_701_n N_Y_c_787_n N_Y_c_702_n N_Y_c_697_n N_Y_c_714_n N_Y_c_715_n Y Y
+ N_Y_c_755_n Y N_Y_c_760_n PM_SKY130_FD_SC_LP__O22AI_4%Y
x_PM_SKY130_FD_SC_LP__O22AI_4%A_821_367# N_A_821_367#_M1000_d
+ N_A_821_367#_M1020_d N_A_821_367#_M1013_s N_A_821_367#_M1028_s
+ N_A_821_367#_c_872_n N_A_821_367#_c_854_n N_A_821_367#_c_844_n
+ N_A_821_367#_c_874_n N_A_821_367#_c_846_n N_A_821_367#_c_860_n
+ N_A_821_367#_c_877_n N_A_821_367#_c_848_n N_A_821_367#_c_864_n
+ N_A_821_367#_c_880_n N_A_821_367#_c_866_n
+ PM_SKY130_FD_SC_LP__O22AI_4%A_821_367#
x_PM_SKY130_FD_SC_LP__O22AI_4%A_33_47# N_A_33_47#_M1001_d N_A_33_47#_M1006_d
+ N_A_33_47#_M1011_d N_A_33_47#_M1023_d N_A_33_47#_M1017_d N_A_33_47#_M1015_d
+ N_A_33_47#_M1008_s N_A_33_47#_M1030_s N_A_33_47#_M1027_d N_A_33_47#_c_881_n
+ N_A_33_47#_c_882_n N_A_33_47#_c_883_n N_A_33_47#_c_954_p N_A_33_47#_c_884_n
+ N_A_33_47#_c_955_p N_A_33_47#_c_885_n N_A_33_47#_c_956_p N_A_33_47#_c_886_n
+ N_A_33_47#_c_958_p N_A_33_47#_c_922_n N_A_33_47#_c_887_n N_A_33_47#_c_888_n
+ N_A_33_47#_c_889_n N_A_33_47#_c_890_n PM_SKY130_FD_SC_LP__O22AI_4%A_33_47#
x_PM_SKY130_FD_SC_LP__O22AI_4%VGND N_VGND_M1001_s N_VGND_M1016_s N_VGND_M1014_s
+ N_VGND_M1026_s N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n
+ N_VGND_c_979_n N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n
+ N_VGND_c_984_n VGND N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n
+ N_VGND_c_988_n PM_SKY130_FD_SC_LP__O22AI_4%VGND
cc_1 VNB N_A1_M1001_g 0.0284365f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_2 VNB N_A1_M1002_g 0.00212106f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.465
cc_3 VNB N_A1_M1006_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_4 VNB N_A1_M1005_g 0.00134439f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.465
cc_5 VNB N_A1_M1016_g 0.0209507f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.655
cc_6 VNB N_A1_M1012_g 0.00124287f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=2.465
cc_7 VNB N_A1_M1017_g 0.0208017f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=0.655
cc_8 VNB N_A1_M1025_g 0.00249937f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_9 VNB N_A1_c_124_n 0.018975f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.487
cc_10 VNB N_A1_c_125_n 3.10976e-19 $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=1.95
cc_11 VNB N_A1_c_126_n 0.00232718f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.63
cc_12 VNB N_A1_c_127_n 0.002369f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=1.44
cc_13 VNB N_A1_c_128_n 0.0306239f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=1.44
cc_14 VNB A1 2.42494e-19 $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_15 VNB N_A1_c_130_n 0.0913342f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.46
cc_16 VNB N_A2_M1011_g 0.0235502f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_17 VNB N_A2_M1014_g 0.023273f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_18 VNB N_A2_M1023_g 0.023273f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.655
cc_19 VNB N_A2_M1026_g 0.0234281f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=0.655
cc_20 VNB A2 0.00236206f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_21 VNB N_A2_c_254_n 0.064737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_M1007_g 0.021536f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_23 VNB N_B1_M1000_g 0.00269364f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.465
cc_24 VNB N_B1_M1015_g 0.0202411f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_25 VNB N_B1_M1009_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.465
cc_26 VNB N_B1_M1024_g 0.0197358f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.655
cc_27 VNB N_B1_M1020_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=2.465
cc_28 VNB N_B1_M1029_g 0.00813779f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_29 VNB N_B1_c_341_n 0.0130822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_c_342_n 0.00423877f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_31 VNB N_B1_c_343_n 0.033272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B1_c_344_n 0.0575871f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.95
cc_33 VNB N_B1_c_345_n 0.019576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B1_c_346_n 0.00467605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B1_c_347_n 0.00154988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B1_c_348_n 0.00444237f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.46
cc_37 VNB N_B2_M1008_g 0.0201095f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_38 VNB N_B2_M1004_g 0.00257191f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.465
cc_39 VNB N_B2_M1018_g 0.0199088f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_40 VNB N_B2_M1013_g 0.00228709f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.465
cc_41 VNB N_B2_M1030_g 0.0199122f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.655
cc_42 VNB N_B2_M1021_g 0.00228709f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=2.465
cc_43 VNB N_B2_M1031_g 0.0201064f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=0.655
cc_44 VNB N_B2_M1028_g 0.00257136f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_45 VNB N_B2_c_467_n 0.0802356f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.95
cc_46 VNB N_VPWR_c_547_n 0.322901f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=1.605
cc_47 VNB N_Y_c_696_n 0.0110107f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_48 VNB N_Y_c_697_n 0.0370652f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.95
cc_49 VNB N_A_33_47#_c_881_n 0.0284746f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_50 VNB N_A_33_47#_c_882_n 0.00289934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_33_47#_c_883_n 0.00901278f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.487
cc_52 VNB N_A_33_47#_c_884_n 0.0099995f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.487
cc_53 VNB N_A_33_47#_c_885_n 0.00306278f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.487
cc_54 VNB N_A_33_47#_c_886_n 0.0126689f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=1.44
cc_55 VNB N_A_33_47#_c_887_n 0.00936708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_33_47#_c_888_n 0.00144427f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_57 VNB N_A_33_47#_c_889_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_33_47#_c_890_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.46
cc_59 VNB N_VGND_c_975_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.465
cc_60 VNB N_VGND_c_976_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.655
cc_61 VNB N_VGND_c_977_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=2.465
cc_62 VNB N_VGND_c_978_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=0.655
cc_63 VNB N_VGND_c_979_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_64 VNB N_VGND_c_980_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=2.465
cc_65 VNB N_VGND_c_981_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.487
cc_66 VNB N_VGND_c_982_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.487
cc_67 VNB N_VGND_c_983_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_68 VNB N_VGND_c_984_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_985_n 0.0163305f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_70 VNB N_VGND_c_986_n 0.0982923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_987_n 0.373079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_988_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VPB N_A1_M1002_g 0.0272599f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.465
cc_74 VPB N_A1_M1005_g 0.0195346f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.465
cc_75 VPB N_A1_M1012_g 0.0191536f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=2.465
cc_76 VPB N_A1_M1025_g 0.020213f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.465
cc_77 VPB N_A1_c_125_n 0.00143437f $X=-0.19 $Y=1.655 $X2=3.47 $Y2=1.95
cc_78 VPB A1 0.00182096f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_79 VPB N_A2_M1003_g 0.0187402f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.465
cc_80 VPB N_A2_M1010_g 0.0181378f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.465
cc_81 VPB N_A2_M1019_g 0.0181366f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=2.465
cc_82 VPB N_A2_M1022_g 0.0183228f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.465
cc_83 VPB A2 0.00919786f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_84 VPB N_A2_c_254_n 0.0127351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_B1_M1000_g 0.019392f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.465
cc_86 VPB N_B1_M1009_g 0.0184959f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.465
cc_87 VPB N_B1_M1020_g 0.018645f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=2.465
cc_88 VPB N_B1_M1029_g 0.0228733f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.465
cc_89 VPB N_B2_M1004_g 0.0188365f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.465
cc_90 VPB N_B2_M1013_g 0.0193316f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.465
cc_91 VPB N_B2_M1021_g 0.0193316f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=2.465
cc_92 VPB N_B2_M1028_g 0.0188168f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.465
cc_93 VPB N_B2_c_472_n 0.00260722f $X=-0.19 $Y=1.655 $X2=3.385 $Y2=2.035
cc_94 VPB N_VPWR_c_548_n 0.012219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_549_n 0.0554469f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.655
cc_96 VPB N_VPWR_c_550_n 4.06069e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_551_n 0.00269594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_552_n 0.0133881f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=2.465
cc_99 VPB N_VPWR_c_553_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.487
cc_100 VPB N_VPWR_c_554_n 0.015603f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_101 VPB N_VPWR_c_555_n 0.0413341f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.487
cc_102 VPB N_VPWR_c_556_n 0.0535028f $X=-0.19 $Y=1.655 $X2=3.47 $Y2=1.95
cc_103 VPB N_VPWR_c_557_n 0.00483875f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.63
cc_104 VPB N_VPWR_c_558_n 0.0148832f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.46
cc_105 VPB N_VPWR_c_559_n 0.0509662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_560_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=1.46
cc_107 VPB N_VPWR_c_561_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=1.46
cc_108 VPB N_VPWR_c_547_n 0.0528199f $X=-0.19 $Y=1.655 $X2=3.55 $Y2=1.605
cc_109 VPB N_A_119_367#_c_655_n 0.00251931f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.465
cc_110 VPB N_Y_c_698_n 0.00754068f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=1.487
cc_111 VPB N_Y_c_699_n 0.00612848f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.487
cc_112 VPB N_Y_c_700_n 0.00298266f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.63
cc_113 VPB N_Y_c_701_n 0.00298266f $X=-0.19 $Y=1.655 $X2=3.55 $Y2=1.44
cc_114 VPB N_Y_c_702_n 0.0218214f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_115 VPB N_Y_c_697_n 0.00247608f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.95
cc_116 N_A1_M1016_g N_A2_M1011_g 0.0225092f $X=1.365 $Y=0.655 $X2=0 $Y2=0
cc_117 N_A1_c_130_n N_A2_M1011_g 0.00971091f $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_118 N_A1_M1012_g N_A2_M1003_g 0.035354f $X=1.38 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A1_c_140_p N_A2_M1003_g 0.015106f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_120 A1 N_A2_M1003_g 0.00150758f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_121 N_A1_c_140_p N_A2_M1010_g 0.0106743f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_122 N_A1_c_140_p N_A2_M1019_g 0.0106743f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_123 N_A1_M1017_g N_A2_M1026_g 0.0214932f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_124 N_A1_c_128_n N_A2_M1026_g 0.0153566f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_125 N_A1_c_125_n N_A2_M1022_g 0.00394299f $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_126 N_A1_c_140_p N_A2_M1022_g 0.0106277f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_127 N_A1_M1012_g A2 3.49926e-19 $X=1.38 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A1_M1025_g A2 4.99531e-19 $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A1_c_125_n A2 0.0178591f $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_130 N_A1_c_126_n A2 0.0132261f $X=1.24 $Y=1.63 $X2=0 $Y2=0
cc_131 N_A1_c_127_n A2 0.0144452f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_132 N_A1_c_128_n A2 0.00121415f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_133 N_A1_c_140_p A2 0.0828357f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_134 A1 A2 0.00530552f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_135 N_A1_c_130_n A2 3.12103e-19 $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_136 N_A1_M1012_g N_A2_c_254_n 0.00971091f $X=1.38 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A1_M1025_g N_A2_c_254_n 0.0566206f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A1_c_125_n N_A2_c_254_n 5.17472e-19 $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_139 N_A1_c_126_n N_A2_c_254_n 0.00131758f $X=1.24 $Y=1.63 $X2=0 $Y2=0
cc_140 N_A1_c_127_n N_A2_c_254_n 2.03455e-19 $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_141 N_A1_c_128_n N_A2_c_254_n 0.00502885f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_142 N_A1_c_140_p N_A2_c_254_n 0.00170125f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_143 A1 N_A2_c_254_n 2.07027e-19 $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_144 N_A1_M1017_g N_B1_M1007_g 0.0156599f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_145 N_A1_M1025_g N_B1_M1000_g 0.0398062f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A1_c_125_n N_B1_M1000_g 2.35822e-19 $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_147 N_A1_c_125_n N_B1_c_344_n 9.34811e-19 $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_148 N_A1_c_127_n N_B1_c_344_n 4.52288e-19 $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_149 N_A1_c_128_n N_B1_c_344_n 0.0209981f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_150 N_A1_M1017_g N_B1_c_347_n 3.33682e-19 $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A1_c_125_n N_B1_c_347_n 3.81205e-19 $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_152 N_A1_c_127_n N_B1_c_347_n 0.0107485f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_153 N_A1_c_128_n N_B1_c_347_n 6.9215e-19 $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_154 A1 N_VPWR_M1005_s 0.00249603f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_155 N_A1_M1002_g N_VPWR_c_549_n 0.0076281f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A1_c_124_n N_VPWR_c_549_n 0.0237411f $X=1.025 $Y=1.487 $X2=0 $Y2=0
cc_157 N_A1_c_130_n N_VPWR_c_549_n 0.00222894f $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_158 N_A1_M1002_g N_VPWR_c_550_n 5.9204e-19 $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A1_M1005_g N_VPWR_c_550_n 0.0101807f $X=0.95 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A1_M1012_g N_VPWR_c_550_n 0.0112591f $X=1.38 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A1_M1025_g N_VPWR_c_551_n 0.00353939f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A1_M1012_g N_VPWR_c_556_n 0.00486043f $X=1.38 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A1_M1025_g N_VPWR_c_556_n 0.00547467f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A1_M1002_g N_VPWR_c_558_n 0.00585385f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A1_M1005_g N_VPWR_c_558_n 0.00486043f $X=0.95 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A1_M1002_g N_VPWR_c_547_n 0.0115086f $X=0.52 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A1_M1005_g N_VPWR_c_547_n 0.00824727f $X=0.95 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A1_M1012_g N_VPWR_c_547_n 0.0082726f $X=1.38 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A1_M1025_g N_VPWR_c_547_n 0.0063959f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A1_c_140_p N_A_119_367#_M1012_d 0.00809843f $X=3.385 $Y=2.035 $X2=0
+ $Y2=0
cc_171 N_A1_c_140_p N_A_119_367#_M1010_s 0.00345037f $X=3.385 $Y=2.035 $X2=0
+ $Y2=0
cc_172 N_A1_c_125_n N_A_119_367#_M1022_s 0.00136045f $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_173 N_A1_c_140_p N_A_119_367#_M1022_s 0.00755195f $X=3.385 $Y=2.035 $X2=0
+ $Y2=0
cc_174 N_A1_M1002_g N_A_119_367#_c_655_n 4.85227e-19 $X=0.52 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A1_M1005_g N_A_119_367#_c_655_n 4.69998e-19 $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A1_c_124_n N_A_119_367#_c_655_n 0.0208506f $X=1.025 $Y=1.487 $X2=0
+ $Y2=0
cc_177 A1 N_A_119_367#_c_655_n 0.00158296f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_178 N_A1_c_130_n N_A_119_367#_c_655_n 7.7261e-19 $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_179 N_A1_M1005_g N_A_119_367#_c_665_n 0.0144438f $X=0.95 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1012_g N_A_119_367#_c_665_n 0.0122068f $X=1.38 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A1_c_124_n N_A_119_367#_c_665_n 0.00370588f $X=1.025 $Y=1.487 $X2=0
+ $Y2=0
cc_182 A1 N_A_119_367#_c_665_n 0.0248978f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_183 N_A1_c_130_n N_A_119_367#_c_665_n 2.63801e-19 $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_184 N_A1_c_140_p N_A_119_367#_c_670_n 0.0135055f $X=3.385 $Y=2.035 $X2=0
+ $Y2=0
cc_185 N_A1_M1025_g N_A_119_367#_c_671_n 0.00358529f $X=3.53 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A1_c_140_p N_A_119_367#_c_671_n 0.00335247f $X=3.385 $Y=2.035 $X2=0
+ $Y2=0
cc_187 N_A1_c_140_p N_Y_M1003_d 0.00345037f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_188 N_A1_c_140_p N_Y_M1019_d 0.00345037f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_189 N_A1_M1025_g N_Y_c_706_n 0.0142086f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A1_c_128_n N_Y_c_706_n 0.00198469f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_191 N_A1_c_140_p N_Y_c_706_n 0.00852791f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_192 N_A1_M1025_g N_Y_c_709_n 0.00521948f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A1_c_125_n N_Y_c_709_n 0.00405209f $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_194 N_A1_c_140_p N_Y_c_709_n 0.0103974f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_195 N_A1_M1025_g N_Y_c_699_n 0.00134994f $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A1_c_125_n N_Y_c_699_n 0.0107026f $X=3.47 $Y=1.95 $X2=0 $Y2=0
cc_197 N_A1_c_140_p N_Y_c_714_n 0.0807147f $X=3.385 $Y=2.035 $X2=0 $Y2=0
cc_198 N_A1_M1025_g N_Y_c_715_n 7.2002e-19 $X=3.53 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A1_M1001_g N_A_33_47#_c_882_n 0.0142722f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A1_M1006_g N_A_33_47#_c_882_n 0.0134628f $X=0.935 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A1_c_124_n N_A_33_47#_c_882_n 0.0463719f $X=1.025 $Y=1.487 $X2=0 $Y2=0
cc_202 N_A1_c_126_n N_A_33_47#_c_882_n 0.00236015f $X=1.24 $Y=1.63 $X2=0 $Y2=0
cc_203 N_A1_c_130_n N_A_33_47#_c_882_n 0.00350824f $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_204 N_A1_c_124_n N_A_33_47#_c_883_n 0.0217074f $X=1.025 $Y=1.487 $X2=0 $Y2=0
cc_205 N_A1_c_130_n N_A_33_47#_c_883_n 0.00643463f $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_206 N_A1_M1016_g N_A_33_47#_c_884_n 0.0134101f $X=1.365 $Y=0.655 $X2=0 $Y2=0
cc_207 N_A1_c_126_n N_A_33_47#_c_884_n 0.0161841f $X=1.24 $Y=1.63 $X2=0 $Y2=0
cc_208 N_A1_c_130_n N_A_33_47#_c_884_n 4.18914e-19 $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_209 N_A1_M1017_g N_A_33_47#_c_886_n 0.0132546f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A1_c_127_n N_A_33_47#_c_886_n 0.0238342f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_211 N_A1_c_128_n N_A_33_47#_c_886_n 0.00452562f $X=3.55 $Y=1.44 $X2=0 $Y2=0
cc_212 N_A1_c_126_n N_A_33_47#_c_888_n 0.0169405f $X=1.24 $Y=1.63 $X2=0 $Y2=0
cc_213 N_A1_c_130_n N_A_33_47#_c_888_n 0.00253548f $X=1.38 $Y=1.46 $X2=0 $Y2=0
cc_214 N_A1_M1001_g N_VGND_c_975_n 0.0118416f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_215 N_A1_M1006_g N_VGND_c_975_n 0.010086f $X=0.935 $Y=0.655 $X2=0 $Y2=0
cc_216 N_A1_M1016_g N_VGND_c_975_n 6.11179e-19 $X=1.365 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A1_M1006_g N_VGND_c_976_n 6.11179e-19 $X=0.935 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A1_M1016_g N_VGND_c_976_n 0.0100502f $X=1.365 $Y=0.655 $X2=0 $Y2=0
cc_219 N_A1_M1017_g N_VGND_c_978_n 0.0112815f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_220 N_A1_M1006_g N_VGND_c_979_n 0.00486043f $X=0.935 $Y=0.655 $X2=0 $Y2=0
cc_221 N_A1_M1016_g N_VGND_c_979_n 0.00486043f $X=1.365 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A1_M1001_g N_VGND_c_985_n 0.00486043f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_223 N_A1_M1017_g N_VGND_c_986_n 0.00486043f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_224 N_A1_M1001_g N_VGND_c_987_n 0.00920706f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_225 N_A1_M1006_g N_VGND_c_987_n 0.00824727f $X=0.935 $Y=0.655 $X2=0 $Y2=0
cc_226 N_A1_M1016_g N_VGND_c_987_n 0.00824727f $X=1.365 $Y=0.655 $X2=0 $Y2=0
cc_227 N_A1_M1017_g N_VGND_c_987_n 0.00839973f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_228 N_A2_M1003_g N_VPWR_c_550_n 0.00109252f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A2_M1003_g N_VPWR_c_556_n 0.00357877f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A2_M1010_g N_VPWR_c_556_n 0.00357877f $X=2.24 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A2_M1019_g N_VPWR_c_556_n 0.00357877f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A2_M1022_g N_VPWR_c_556_n 0.00357877f $X=3.1 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A2_M1003_g N_VPWR_c_547_n 0.00537654f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A2_M1010_g N_VPWR_c_547_n 0.0053512f $X=2.24 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A2_M1019_g N_VPWR_c_547_n 0.0053512f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A2_M1022_g N_VPWR_c_547_n 0.00537654f $X=3.1 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A2_M1003_g N_A_119_367#_c_671_n 0.0130424f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A2_M1010_g N_A_119_367#_c_671_n 0.0106414f $X=2.24 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A2_M1019_g N_A_119_367#_c_671_n 0.0107199f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A2_M1022_g N_A_119_367#_c_671_n 0.0114335f $X=3.1 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A2_M1022_g N_Y_c_706_n 0.00824286f $X=3.1 $Y=2.465 $X2=0 $Y2=0
cc_242 N_A2_M1010_g N_Y_c_714_n 0.0127032f $X=2.24 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A2_M1019_g N_Y_c_714_n 0.0126123f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A2_M1022_g N_Y_c_715_n 0.00402437f $X=3.1 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A2_M1011_g N_A_33_47#_c_884_n 0.0161281f $X=1.795 $Y=0.655 $X2=0 $Y2=0
cc_246 A2 N_A_33_47#_c_884_n 0.00775529f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A2_M1014_g N_A_33_47#_c_885_n 0.0134628f $X=2.225 $Y=0.655 $X2=0 $Y2=0
cc_248 N_A2_M1023_g N_A_33_47#_c_885_n 0.0134628f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_249 A2 N_A_33_47#_c_885_n 0.0499611f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_250 N_A2_c_254_n N_A_33_47#_c_885_n 0.00230115f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_251 N_A2_M1026_g N_A_33_47#_c_886_n 0.0134162f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_252 A2 N_A_33_47#_c_886_n 0.0179166f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_253 A2 N_A_33_47#_c_889_n 0.0162531f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_254 N_A2_c_254_n N_A_33_47#_c_889_n 0.00238873f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_255 A2 N_A_33_47#_c_890_n 0.0162531f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_256 N_A2_c_254_n N_A_33_47#_c_890_n 0.00238873f $X=3.085 $Y=1.51 $X2=0 $Y2=0
cc_257 N_A2_M1011_g N_VGND_c_976_n 0.0100502f $X=1.795 $Y=0.655 $X2=0 $Y2=0
cc_258 N_A2_M1014_g N_VGND_c_976_n 6.11179e-19 $X=2.225 $Y=0.655 $X2=0 $Y2=0
cc_259 N_A2_M1011_g N_VGND_c_977_n 6.11179e-19 $X=1.795 $Y=0.655 $X2=0 $Y2=0
cc_260 N_A2_M1014_g N_VGND_c_977_n 0.010086f $X=2.225 $Y=0.655 $X2=0 $Y2=0
cc_261 N_A2_M1023_g N_VGND_c_977_n 0.010086f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A2_M1026_g N_VGND_c_977_n 6.11179e-19 $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_263 N_A2_M1023_g N_VGND_c_978_n 6.11179e-19 $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_264 N_A2_M1026_g N_VGND_c_978_n 0.0100502f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_265 N_A2_M1011_g N_VGND_c_981_n 0.00486043f $X=1.795 $Y=0.655 $X2=0 $Y2=0
cc_266 N_A2_M1014_g N_VGND_c_981_n 0.00486043f $X=2.225 $Y=0.655 $X2=0 $Y2=0
cc_267 N_A2_M1023_g N_VGND_c_983_n 0.00486043f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_268 N_A2_M1026_g N_VGND_c_983_n 0.00486043f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_269 N_A2_M1011_g N_VGND_c_987_n 0.00824727f $X=1.795 $Y=0.655 $X2=0 $Y2=0
cc_270 N_A2_M1014_g N_VGND_c_987_n 0.00824727f $X=2.225 $Y=0.655 $X2=0 $Y2=0
cc_271 N_A2_M1023_g N_VGND_c_987_n 0.00824727f $X=2.655 $Y=0.655 $X2=0 $Y2=0
cc_272 N_A2_M1026_g N_VGND_c_987_n 0.00824727f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_273 N_B1_M1024_g N_B2_M1008_g 0.0358959f $X=4.86 $Y=0.655 $X2=0 $Y2=0
cc_274 N_B1_c_341_n N_B2_M1008_g 0.01044f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_275 N_B1_c_348_n N_B2_M1008_g 0.00605565f $X=5.005 $Y=1.09 $X2=0 $Y2=0
cc_276 N_B1_M1020_g N_B2_M1004_g 0.0256206f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_277 N_B1_c_341_n N_B2_M1018_g 0.010446f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_278 N_B1_c_341_n N_B2_M1030_g 0.0104771f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_279 N_B1_c_341_n N_B2_M1031_g 0.010446f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_280 N_B1_c_342_n N_B2_M1031_g 0.00196985f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_281 N_B1_c_345_n N_B2_M1031_g 0.0363647f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_282 N_B1_c_341_n N_B2_c_482_n 0.0376261f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_283 N_B1_c_342_n N_B2_c_482_n 0.00954582f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_284 N_B1_c_343_n N_B2_c_482_n 2.04223e-19 $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_285 N_B1_c_341_n N_B2_c_472_n 0.0591438f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_286 N_B1_c_348_n N_B2_c_472_n 0.014415f $X=5.005 $Y=1.09 $X2=0 $Y2=0
cc_287 N_B1_M1029_g N_B2_c_467_n 0.0300728f $X=7.04 $Y=2.465 $X2=0 $Y2=0
cc_288 N_B1_c_341_n N_B2_c_467_n 0.00867291f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_289 N_B1_c_342_n N_B2_c_467_n 0.00270226f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_290 N_B1_c_343_n N_B2_c_467_n 0.0129091f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_291 N_B1_c_344_n N_B2_c_467_n 0.0186519f $X=4.86 $Y=1.44 $X2=0 $Y2=0
cc_292 N_B1_M1000_g N_VPWR_c_551_n 0.00834448f $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_293 N_B1_M1009_g N_VPWR_c_551_n 5.51453e-19 $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_294 N_B1_M1000_g N_VPWR_c_552_n 0.00564095f $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_295 N_B1_M1009_g N_VPWR_c_552_n 0.00486043f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_296 N_B1_M1000_g N_VPWR_c_553_n 6.50463e-19 $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_297 N_B1_M1009_g N_VPWR_c_553_n 0.0117756f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_298 N_B1_M1020_g N_VPWR_c_553_n 0.0129021f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_299 N_B1_M1029_g N_VPWR_c_555_n 0.0164126f $X=7.04 $Y=2.465 $X2=0 $Y2=0
cc_300 N_B1_M1020_g N_VPWR_c_559_n 0.00486043f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_301 N_B1_M1029_g N_VPWR_c_559_n 0.00486043f $X=7.04 $Y=2.465 $X2=0 $Y2=0
cc_302 N_B1_M1000_g N_VPWR_c_547_n 0.00948291f $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_303 N_B1_M1009_g N_VPWR_c_547_n 0.00824727f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_304 N_B1_M1020_g N_VPWR_c_547_n 0.0082726f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_305 N_B1_M1029_g N_VPWR_c_547_n 0.0082726f $X=7.04 $Y=2.465 $X2=0 $Y2=0
cc_306 N_B1_c_341_n N_Y_M1024_s 5.19434e-19 $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_307 N_B1_c_348_n N_Y_M1024_s 0.00161671f $X=5.005 $Y=1.09 $X2=0 $Y2=0
cc_308 N_B1_c_341_n N_Y_M1018_d 0.00176891f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_309 N_B1_c_341_n N_Y_M1031_d 0.00176891f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_310 N_B1_M1000_g N_Y_c_706_n 0.00410192f $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_311 N_B1_M1000_g N_Y_c_709_n 0.00860806f $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_312 N_B1_M1009_g N_Y_c_709_n 7.41383e-19 $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_313 N_B1_M1000_g N_Y_c_698_n 0.0126188f $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_314 N_B1_M1009_g N_Y_c_698_n 0.010446f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_315 N_B1_M1020_g N_Y_c_698_n 0.0104291f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_316 N_B1_c_341_n N_Y_c_698_n 0.00559513f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_317 N_B1_c_344_n N_Y_c_698_n 0.00512592f $X=4.86 $Y=1.44 $X2=0 $Y2=0
cc_318 N_B1_c_346_n N_Y_c_698_n 0.0537927f $X=4.885 $Y=1.372 $X2=0 $Y2=0
cc_319 N_B1_c_347_n N_Y_c_698_n 0.0141727f $X=4.157 $Y=1.372 $X2=0 $Y2=0
cc_320 N_B1_c_348_n N_Y_c_698_n 0.0190504f $X=5.005 $Y=1.09 $X2=0 $Y2=0
cc_321 N_B1_M1000_g N_Y_c_699_n 0.00173418f $X=4.03 $Y=2.465 $X2=0 $Y2=0
cc_322 N_B1_c_344_n N_Y_c_699_n 0.00129031f $X=4.86 $Y=1.44 $X2=0 $Y2=0
cc_323 N_B1_c_347_n N_Y_c_699_n 3.84502e-19 $X=4.157 $Y=1.372 $X2=0 $Y2=0
cc_324 N_B1_M1024_g N_Y_c_696_n 0.00968963f $X=4.86 $Y=0.655 $X2=0 $Y2=0
cc_325 N_B1_c_341_n N_Y_c_696_n 0.107389f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_326 N_B1_c_343_n N_Y_c_696_n 0.00262758f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_327 N_B1_c_345_n N_Y_c_696_n 0.0108522f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_328 N_B1_c_346_n N_Y_c_696_n 0.00573827f $X=4.885 $Y=1.372 $X2=0 $Y2=0
cc_329 N_B1_c_348_n N_Y_c_696_n 0.0142553f $X=5.005 $Y=1.09 $X2=0 $Y2=0
cc_330 N_B1_M1020_g N_Y_c_700_n 7.60491e-19 $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_331 N_B1_M1029_g N_Y_c_701_n 7.75429e-19 $X=7.04 $Y=2.465 $X2=0 $Y2=0
cc_332 N_B1_M1029_g N_Y_c_702_n 0.016109f $X=7.04 $Y=2.465 $X2=0 $Y2=0
cc_333 N_B1_c_341_n N_Y_c_702_n 0.00928473f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_334 N_B1_c_342_n N_Y_c_702_n 0.0183297f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_335 N_B1_c_343_n N_Y_c_702_n 0.0033578f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_336 N_B1_M1029_g N_Y_c_697_n 0.00593838f $X=7.04 $Y=2.465 $X2=0 $Y2=0
cc_337 N_B1_c_341_n N_Y_c_697_n 0.0141404f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_338 N_B1_c_342_n N_Y_c_697_n 0.0251291f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_339 N_B1_c_343_n N_Y_c_697_n 0.00803689f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_340 N_B1_c_345_n N_Y_c_697_n 0.00613674f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_341 N_B1_M1007_g N_Y_c_755_n 0.00928855f $X=4 $Y=0.655 $X2=0 $Y2=0
cc_342 N_B1_M1015_g N_Y_c_755_n 0.0147855f $X=4.43 $Y=0.655 $X2=0 $Y2=0
cc_343 N_B1_c_344_n N_Y_c_755_n 6.31585e-19 $X=4.86 $Y=1.44 $X2=0 $Y2=0
cc_344 N_B1_c_346_n N_Y_c_755_n 0.0404181f $X=4.885 $Y=1.372 $X2=0 $Y2=0
cc_345 N_B1_c_347_n N_Y_c_755_n 0.0110157f $X=4.157 $Y=1.372 $X2=0 $Y2=0
cc_346 N_B1_M1024_g N_Y_c_760_n 0.00554745f $X=4.86 $Y=0.655 $X2=0 $Y2=0
cc_347 N_B1_c_344_n N_Y_c_760_n 6.31585e-19 $X=4.86 $Y=1.44 $X2=0 $Y2=0
cc_348 N_B1_c_348_n N_Y_c_760_n 0.00274663f $X=5.005 $Y=1.09 $X2=0 $Y2=0
cc_349 N_B1_M1009_g N_A_821_367#_c_844_n 0.0125125f $X=4.46 $Y=2.465 $X2=0 $Y2=0
cc_350 N_B1_M1020_g N_A_821_367#_c_844_n 0.0124988f $X=4.89 $Y=2.465 $X2=0 $Y2=0
cc_351 N_B1_c_341_n N_A_33_47#_M1008_s 0.00176891f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_352 N_B1_c_341_n N_A_33_47#_M1030_s 0.00176891f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_353 N_B1_c_341_n N_A_33_47#_M1027_d 0.00134836f $X=6.93 $Y=1.09 $X2=0 $Y2=0
cc_354 N_B1_M1007_g N_A_33_47#_c_886_n 0.00406925f $X=4 $Y=0.655 $X2=0 $Y2=0
cc_355 N_B1_M1007_g N_A_33_47#_c_922_n 0.00461003f $X=4 $Y=0.655 $X2=0 $Y2=0
cc_356 N_B1_M1007_g N_A_33_47#_c_887_n 0.0108801f $X=4 $Y=0.655 $X2=0 $Y2=0
cc_357 N_B1_M1015_g N_A_33_47#_c_887_n 0.00900817f $X=4.43 $Y=0.655 $X2=0 $Y2=0
cc_358 N_B1_M1024_g N_A_33_47#_c_887_n 0.00894775f $X=4.86 $Y=0.655 $X2=0 $Y2=0
cc_359 N_B1_c_345_n N_A_33_47#_c_887_n 0.00894775f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_360 N_B1_M1007_g N_VGND_c_978_n 0.00101295f $X=4 $Y=0.655 $X2=0 $Y2=0
cc_361 N_B1_M1007_g N_VGND_c_986_n 0.00357877f $X=4 $Y=0.655 $X2=0 $Y2=0
cc_362 N_B1_M1015_g N_VGND_c_986_n 0.00357877f $X=4.43 $Y=0.655 $X2=0 $Y2=0
cc_363 N_B1_M1024_g N_VGND_c_986_n 0.00357877f $X=4.86 $Y=0.655 $X2=0 $Y2=0
cc_364 N_B1_c_345_n N_VGND_c_986_n 0.00357877f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_365 N_B1_M1007_g N_VGND_c_987_n 0.00550366f $X=4 $Y=0.655 $X2=0 $Y2=0
cc_366 N_B1_M1015_g N_VGND_c_987_n 0.0053512f $X=4.43 $Y=0.655 $X2=0 $Y2=0
cc_367 N_B1_M1024_g N_VGND_c_987_n 0.00537849f $X=4.86 $Y=0.655 $X2=0 $Y2=0
cc_368 N_B1_c_345_n N_VGND_c_987_n 0.00645063f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_369 N_B2_M1004_g N_VPWR_c_553_n 0.00109252f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_370 N_B2_M1028_g N_VPWR_c_555_n 0.00109252f $X=6.61 $Y=2.465 $X2=0 $Y2=0
cc_371 N_B2_M1004_g N_VPWR_c_559_n 0.00357877f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_372 N_B2_M1013_g N_VPWR_c_559_n 0.00357877f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_373 N_B2_M1021_g N_VPWR_c_559_n 0.00357877f $X=6.18 $Y=2.465 $X2=0 $Y2=0
cc_374 N_B2_M1028_g N_VPWR_c_559_n 0.00357877f $X=6.61 $Y=2.465 $X2=0 $Y2=0
cc_375 N_B2_M1004_g N_VPWR_c_547_n 0.00537654f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_376 N_B2_M1013_g N_VPWR_c_547_n 0.0053512f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_377 N_B2_M1021_g N_VPWR_c_547_n 0.0053512f $X=6.18 $Y=2.465 $X2=0 $Y2=0
cc_378 N_B2_M1028_g N_VPWR_c_547_n 0.00537654f $X=6.61 $Y=2.465 $X2=0 $Y2=0
cc_379 N_B2_M1004_g N_Y_c_698_n 0.0118156f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_380 N_B2_c_472_n N_Y_c_698_n 0.00440986f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_381 N_B2_c_467_n N_Y_c_698_n 9.85391e-19 $X=6.61 $Y=1.44 $X2=0 $Y2=0
cc_382 N_B2_M1008_g N_Y_c_696_n 0.00895939f $X=5.29 $Y=0.655 $X2=0 $Y2=0
cc_383 N_B2_M1018_g N_Y_c_696_n 0.00895939f $X=5.72 $Y=0.655 $X2=0 $Y2=0
cc_384 N_B2_M1030_g N_Y_c_696_n 0.00894563f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_385 N_B2_M1031_g N_Y_c_696_n 0.00895939f $X=6.58 $Y=0.655 $X2=0 $Y2=0
cc_386 N_B2_M1004_g N_Y_c_700_n 0.00579072f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_387 N_B2_M1013_g N_Y_c_700_n 0.00265591f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_388 N_B2_c_472_n N_Y_c_700_n 0.0280132f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_389 N_B2_c_467_n N_Y_c_700_n 0.00266387f $X=6.61 $Y=1.44 $X2=0 $Y2=0
cc_390 N_B2_M1004_g N_Y_c_774_n 0.00967335f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_391 N_B2_M1013_g N_Y_c_774_n 0.0109251f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_392 N_B2_M1021_g N_Y_c_774_n 5.66402e-19 $X=6.18 $Y=2.465 $X2=0 $Y2=0
cc_393 N_B2_M1013_g N_Y_c_777_n 0.0120127f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_394 N_B2_M1021_g N_Y_c_777_n 0.0120127f $X=6.18 $Y=2.465 $X2=0 $Y2=0
cc_395 N_B2_c_482_n N_Y_c_777_n 0.00379673f $X=6.49 $Y=1.44 $X2=0 $Y2=0
cc_396 N_B2_c_472_n N_Y_c_777_n 0.0240273f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_397 N_B2_c_467_n N_Y_c_777_n 4.80737e-19 $X=6.61 $Y=1.44 $X2=0 $Y2=0
cc_398 N_B2_M1021_g N_Y_c_701_n 0.00265591f $X=6.18 $Y=2.465 $X2=0 $Y2=0
cc_399 N_B2_M1028_g N_Y_c_701_n 0.00579985f $X=6.61 $Y=2.465 $X2=0 $Y2=0
cc_400 N_B2_c_482_n N_Y_c_701_n 0.0233953f $X=6.49 $Y=1.44 $X2=0 $Y2=0
cc_401 N_B2_c_472_n N_Y_c_701_n 0.00461783f $X=5.81 $Y=1.44 $X2=0 $Y2=0
cc_402 N_B2_c_467_n N_Y_c_701_n 0.00266387f $X=6.61 $Y=1.44 $X2=0 $Y2=0
cc_403 N_B2_M1013_g N_Y_c_787_n 5.66402e-19 $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_404 N_B2_M1021_g N_Y_c_787_n 0.0109251f $X=6.18 $Y=2.465 $X2=0 $Y2=0
cc_405 N_B2_M1028_g N_Y_c_787_n 0.00965235f $X=6.61 $Y=2.465 $X2=0 $Y2=0
cc_406 N_B2_M1028_g N_Y_c_702_n 0.0113688f $X=6.61 $Y=2.465 $X2=0 $Y2=0
cc_407 N_B2_c_482_n N_Y_c_702_n 0.00646083f $X=6.49 $Y=1.44 $X2=0 $Y2=0
cc_408 N_B2_M1004_g N_A_821_367#_c_846_n 0.0115031f $X=5.32 $Y=2.465 $X2=0 $Y2=0
cc_409 N_B2_M1013_g N_A_821_367#_c_846_n 0.0114565f $X=5.75 $Y=2.465 $X2=0 $Y2=0
cc_410 N_B2_M1021_g N_A_821_367#_c_848_n 0.0114565f $X=6.18 $Y=2.465 $X2=0 $Y2=0
cc_411 N_B2_M1028_g N_A_821_367#_c_848_n 0.0115031f $X=6.61 $Y=2.465 $X2=0 $Y2=0
cc_412 N_B2_M1008_g N_A_33_47#_c_887_n 0.00894775f $X=5.29 $Y=0.655 $X2=0 $Y2=0
cc_413 N_B2_M1018_g N_A_33_47#_c_887_n 0.00900817f $X=5.72 $Y=0.655 $X2=0 $Y2=0
cc_414 N_B2_M1030_g N_A_33_47#_c_887_n 0.00900817f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_415 N_B2_M1031_g N_A_33_47#_c_887_n 0.00894775f $X=6.58 $Y=0.655 $X2=0 $Y2=0
cc_416 N_B2_M1008_g N_VGND_c_986_n 0.00357877f $X=5.29 $Y=0.655 $X2=0 $Y2=0
cc_417 N_B2_M1018_g N_VGND_c_986_n 0.00357877f $X=5.72 $Y=0.655 $X2=0 $Y2=0
cc_418 N_B2_M1030_g N_VGND_c_986_n 0.00357877f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_419 N_B2_M1031_g N_VGND_c_986_n 0.00357877f $X=6.58 $Y=0.655 $X2=0 $Y2=0
cc_420 N_B2_M1008_g N_VGND_c_987_n 0.00537849f $X=5.29 $Y=0.655 $X2=0 $Y2=0
cc_421 N_B2_M1018_g N_VGND_c_987_n 0.0053512f $X=5.72 $Y=0.655 $X2=0 $Y2=0
cc_422 N_B2_M1030_g N_VGND_c_987_n 0.0053512f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_423 N_B2_M1031_g N_VGND_c_987_n 0.00537849f $X=6.58 $Y=0.655 $X2=0 $Y2=0
cc_424 N_VPWR_c_547_n N_A_119_367#_M1002_d 0.00397496f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_425 N_VPWR_c_547_n N_A_119_367#_M1012_d 0.00376626f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_547_n N_A_119_367#_M1010_s 0.00223577f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_547_n N_A_119_367#_M1022_s 0.00223577f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_549_n N_A_119_367#_c_655_n 0.00153539f $X=0.305 $Y=1.98 $X2=0
+ $Y2=0
cc_429 N_VPWR_M1005_s N_A_119_367#_c_665_n 0.00345322f $X=1.025 $Y=1.835 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_550_n N_A_119_367#_c_665_n 0.0170777f $X=1.165 $Y=2.795 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_556_n N_A_119_367#_c_684_n 0.0128782f $X=3.65 $Y=3.33 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_547_n N_A_119_367#_c_684_n 0.00777554f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_556_n N_A_119_367#_c_671_n 0.100562f $X=3.65 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_547_n N_A_119_367#_c_671_n 0.0644764f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_558_n N_A_119_367#_c_688_n 0.0138717f $X=1 $Y=3.33 $X2=0 $Y2=0
cc_436 N_VPWR_c_547_n N_A_119_367#_c_688_n 0.00886411f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_547_n N_Y_M1003_d 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_438 N_VPWR_c_547_n N_Y_M1019_d 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_c_547_n N_Y_M1004_d 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_440 N_VPWR_c_547_n N_Y_M1021_d 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_441 N_VPWR_M1025_s N_Y_c_706_n 0.00631592f $X=3.605 $Y=1.835 $X2=0 $Y2=0
cc_442 N_VPWR_c_551_n N_Y_c_706_n 0.0200148f $X=3.79 $Y=2.805 $X2=0 $Y2=0
cc_443 N_VPWR_c_547_n N_Y_c_706_n 0.00692128f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_444 N_VPWR_M1025_s N_Y_c_709_n 0.00429079f $X=3.605 $Y=1.835 $X2=0 $Y2=0
cc_445 N_VPWR_M1009_s N_Y_c_698_n 0.00176891f $X=4.535 $Y=1.835 $X2=0 $Y2=0
cc_446 N_VPWR_M1025_s N_Y_c_699_n 3.98562e-19 $X=3.605 $Y=1.835 $X2=0 $Y2=0
cc_447 N_VPWR_M1029_s N_Y_c_702_n 0.00270389f $X=7.115 $Y=1.835 $X2=0 $Y2=0
cc_448 N_VPWR_c_555_n N_Y_c_702_n 0.0179492f $X=7.255 $Y=2.19 $X2=0 $Y2=0
cc_449 N_VPWR_c_547_n N_A_821_367#_M1000_d 0.00467071f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_450 N_VPWR_c_547_n N_A_821_367#_M1020_d 0.00376627f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_547_n N_A_821_367#_M1013_s 0.00223565f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_547_n N_A_821_367#_M1028_s 0.00376627f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_552_n N_A_821_367#_c_854_n 0.0131621f $X=4.51 $Y=3.33 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_547_n N_A_821_367#_c_854_n 0.00808656f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_455 N_VPWR_M1009_s N_A_821_367#_c_844_n 0.00340214f $X=4.535 $Y=1.835 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_553_n N_A_821_367#_c_844_n 0.0171443f $X=4.675 $Y=2.515 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_559_n N_A_821_367#_c_846_n 0.0361172f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_547_n N_A_821_367#_c_846_n 0.023676f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_459 N_VPWR_c_559_n N_A_821_367#_c_860_n 0.0125234f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_547_n N_A_821_367#_c_860_n 0.00738676f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_559_n N_A_821_367#_c_848_n 0.0361172f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_547_n N_A_821_367#_c_848_n 0.023676f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_463 N_VPWR_c_559_n N_A_821_367#_c_864_n 0.0125234f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_547_n N_A_821_367#_c_864_n 0.00738676f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_559_n N_A_821_367#_c_866_n 0.0125234f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_547_n N_A_821_367#_c_866_n 0.00738676f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_467 N_A_119_367#_c_671_n N_Y_M1003_d 0.00338113f $X=3.315 $Y=2.915 $X2=0
+ $Y2=0
cc_468 N_A_119_367#_c_671_n N_Y_M1019_d 0.00338113f $X=3.315 $Y=2.915 $X2=0
+ $Y2=0
cc_469 N_A_119_367#_M1022_s N_Y_c_706_n 0.00408274f $X=3.175 $Y=1.835 $X2=0
+ $Y2=0
cc_470 N_A_119_367#_c_671_n N_Y_c_706_n 0.0129231f $X=3.315 $Y=2.915 $X2=0 $Y2=0
cc_471 N_A_119_367#_M1010_s N_Y_c_714_n 0.00347271f $X=2.315 $Y=1.835 $X2=0
+ $Y2=0
cc_472 N_A_119_367#_c_671_n N_Y_c_714_n 0.0608369f $X=3.315 $Y=2.915 $X2=0 $Y2=0
cc_473 N_Y_c_698_n N_A_821_367#_M1000_d 0.00176461f $X=5.37 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_474 N_Y_c_698_n N_A_821_367#_M1020_d 0.00176461f $X=5.37 $Y=1.79 $X2=0 $Y2=0
cc_475 N_Y_c_777_n N_A_821_367#_M1013_s 0.00335273f $X=6.23 $Y=2.015 $X2=0 $Y2=0
cc_476 N_Y_c_702_n N_A_821_367#_M1028_s 0.00176461f $X=7.365 $Y=1.79 $X2=0 $Y2=0
cc_477 N_Y_c_698_n N_A_821_367#_c_872_n 0.0135055f $X=5.37 $Y=1.79 $X2=0 $Y2=0
cc_478 N_Y_c_698_n N_A_821_367#_c_844_n 0.0324646f $X=5.37 $Y=1.79 $X2=0 $Y2=0
cc_479 N_Y_c_698_n N_A_821_367#_c_874_n 0.0135055f $X=5.37 $Y=1.79 $X2=0 $Y2=0
cc_480 N_Y_M1004_d N_A_821_367#_c_846_n 0.00332344f $X=5.395 $Y=1.835 $X2=0
+ $Y2=0
cc_481 N_Y_c_774_n N_A_821_367#_c_846_n 0.0159805f $X=5.535 $Y=2.615 $X2=0 $Y2=0
cc_482 N_Y_c_777_n N_A_821_367#_c_877_n 0.0135055f $X=6.23 $Y=2.015 $X2=0 $Y2=0
cc_483 N_Y_M1021_d N_A_821_367#_c_848_n 0.00332344f $X=6.255 $Y=1.835 $X2=0
+ $Y2=0
cc_484 N_Y_c_787_n N_A_821_367#_c_848_n 0.0159805f $X=6.395 $Y=2.615 $X2=0 $Y2=0
cc_485 N_Y_c_702_n N_A_821_367#_c_880_n 0.0135055f $X=7.365 $Y=1.79 $X2=0 $Y2=0
cc_486 N_Y_c_696_n N_A_33_47#_M1015_d 3.10352e-19 $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_487 N_Y_c_760_n N_A_33_47#_M1015_d 0.00558684f $X=4.715 $Y=0.842 $X2=0 $Y2=0
cc_488 N_Y_c_696_n N_A_33_47#_M1008_s 0.00334619f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_489 N_Y_c_696_n N_A_33_47#_M1030_s 0.00334619f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_490 N_Y_c_696_n N_A_33_47#_M1027_d 0.00867194f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_491 N_Y_c_697_n N_A_33_47#_M1027_d 0.00278247f $X=7.45 $Y=1.705 $X2=0 $Y2=0
cc_492 N_Y_c_699_n N_A_33_47#_c_886_n 0.00105962f $X=3.96 $Y=1.79 $X2=0 $Y2=0
cc_493 N_Y_c_755_n N_A_33_47#_c_886_n 0.00297172f $X=4.518 $Y=0.842 $X2=0 $Y2=0
cc_494 N_Y_c_755_n N_A_33_47#_c_922_n 0.0282929f $X=4.518 $Y=0.842 $X2=0 $Y2=0
cc_495 N_Y_M1007_s N_A_33_47#_c_887_n 0.00335431f $X=4.075 $Y=0.235 $X2=0 $Y2=0
cc_496 N_Y_M1024_s N_A_33_47#_c_887_n 0.00334357f $X=4.935 $Y=0.235 $X2=0 $Y2=0
cc_497 N_Y_M1018_d N_A_33_47#_c_887_n 0.00335431f $X=5.795 $Y=0.235 $X2=0 $Y2=0
cc_498 N_Y_M1031_d N_A_33_47#_c_887_n 0.00335431f $X=6.655 $Y=0.235 $X2=0 $Y2=0
cc_499 N_Y_c_696_n N_A_33_47#_c_887_n 0.00201845f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_500 N_Y_c_755_n N_A_33_47#_c_887_n 0.175391f $X=4.518 $Y=0.842 $X2=0 $Y2=0
cc_501 N_Y_c_696_n N_VGND_c_986_n 0.00287673f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_502 N_Y_M1007_s N_VGND_c_987_n 0.00225186f $X=4.075 $Y=0.235 $X2=0 $Y2=0
cc_503 N_Y_M1024_s N_VGND_c_987_n 0.00225186f $X=4.935 $Y=0.235 $X2=0 $Y2=0
cc_504 N_Y_M1018_d N_VGND_c_987_n 0.00225186f $X=5.795 $Y=0.235 $X2=0 $Y2=0
cc_505 N_Y_M1031_d N_VGND_c_987_n 0.00225186f $X=6.655 $Y=0.235 $X2=0 $Y2=0
cc_506 N_Y_c_696_n N_VGND_c_987_n 0.00443107f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_507 N_A_33_47#_c_882_n N_VGND_M1001_s 0.00180746f $X=1.055 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_508 N_A_33_47#_c_884_n N_VGND_M1016_s 0.00180746f $X=1.915 $Y=1.09 $X2=0
+ $Y2=0
cc_509 N_A_33_47#_c_885_n N_VGND_M1014_s 0.00180746f $X=2.775 $Y=1.09 $X2=0
+ $Y2=0
cc_510 N_A_33_47#_c_886_n N_VGND_M1026_s 0.00180746f $X=3.635 $Y=1.09 $X2=0
+ $Y2=0
cc_511 N_A_33_47#_c_882_n N_VGND_c_975_n 0.0163515f $X=1.055 $Y=1.09 $X2=0 $Y2=0
cc_512 N_A_33_47#_c_884_n N_VGND_c_976_n 0.0163515f $X=1.915 $Y=1.09 $X2=0 $Y2=0
cc_513 N_A_33_47#_c_885_n N_VGND_c_977_n 0.0163515f $X=2.775 $Y=1.09 $X2=0 $Y2=0
cc_514 N_A_33_47#_c_886_n N_VGND_c_978_n 0.0163515f $X=3.635 $Y=1.09 $X2=0 $Y2=0
cc_515 N_A_33_47#_c_954_p N_VGND_c_979_n 0.0124525f $X=1.15 $Y=0.42 $X2=0 $Y2=0
cc_516 N_A_33_47#_c_955_p N_VGND_c_981_n 0.0124525f $X=2.01 $Y=0.42 $X2=0 $Y2=0
cc_517 N_A_33_47#_c_956_p N_VGND_c_983_n 0.0124525f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_518 N_A_33_47#_c_881_n N_VGND_c_985_n 0.0178111f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_519 N_A_33_47#_c_958_p N_VGND_c_986_n 0.0122383f $X=3.725 $Y=0.475 $X2=0
+ $Y2=0
cc_520 N_A_33_47#_c_887_n N_VGND_c_986_n 0.201378f $X=7.225 $Y=0.37 $X2=0 $Y2=0
cc_521 N_A_33_47#_M1001_d N_VGND_c_987_n 0.00371702f $X=0.165 $Y=0.235 $X2=0
+ $Y2=0
cc_522 N_A_33_47#_M1006_d N_VGND_c_987_n 0.00536646f $X=1.01 $Y=0.235 $X2=0
+ $Y2=0
cc_523 N_A_33_47#_M1011_d N_VGND_c_987_n 0.00536646f $X=1.87 $Y=0.235 $X2=0
+ $Y2=0
cc_524 N_A_33_47#_M1023_d N_VGND_c_987_n 0.00536646f $X=2.73 $Y=0.235 $X2=0
+ $Y2=0
cc_525 N_A_33_47#_M1017_d N_VGND_c_987_n 0.0042086f $X=3.59 $Y=0.235 $X2=0 $Y2=0
cc_526 N_A_33_47#_M1015_d N_VGND_c_987_n 0.00223577f $X=4.505 $Y=0.235 $X2=0
+ $Y2=0
cc_527 N_A_33_47#_M1008_s N_VGND_c_987_n 0.00223577f $X=5.365 $Y=0.235 $X2=0
+ $Y2=0
cc_528 N_A_33_47#_M1030_s N_VGND_c_987_n 0.00223577f $X=6.225 $Y=0.235 $X2=0
+ $Y2=0
cc_529 N_A_33_47#_M1027_d N_VGND_c_987_n 0.00231933f $X=7.085 $Y=0.235 $X2=0
+ $Y2=0
cc_530 N_A_33_47#_c_881_n N_VGND_c_987_n 0.0100304f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_531 N_A_33_47#_c_954_p N_VGND_c_987_n 0.00730901f $X=1.15 $Y=0.42 $X2=0 $Y2=0
cc_532 N_A_33_47#_c_955_p N_VGND_c_987_n 0.00730901f $X=2.01 $Y=0.42 $X2=0 $Y2=0
cc_533 N_A_33_47#_c_956_p N_VGND_c_987_n 0.00730901f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_534 N_A_33_47#_c_958_p N_VGND_c_987_n 0.00699798f $X=3.725 $Y=0.475 $X2=0
+ $Y2=0
cc_535 N_A_33_47#_c_887_n N_VGND_c_987_n 0.12912f $X=7.225 $Y=0.37 $X2=0 $Y2=0
