* File: sky130_fd_sc_lp__inv_1.pxi.spice
* Created: Fri Aug 28 10:38:05 2020
* 
x_PM_SKY130_FD_SC_LP__INV_1%A N_A_M1000_g N_A_M1001_g A A N_A_c_20_n N_A_c_21_n
+ PM_SKY130_FD_SC_LP__INV_1%A
x_PM_SKY130_FD_SC_LP__INV_1%VPWR N_VPWR_M1001_s N_VPWR_c_37_n N_VPWR_c_38_n VPWR
+ N_VPWR_c_39_n N_VPWR_c_36_n PM_SKY130_FD_SC_LP__INV_1%VPWR
x_PM_SKY130_FD_SC_LP__INV_1%Y N_Y_M1000_d N_Y_M1001_d Y Y Y Y Y Y Y N_Y_c_49_n
+ PM_SKY130_FD_SC_LP__INV_1%Y
x_PM_SKY130_FD_SC_LP__INV_1%VGND N_VGND_M1000_s N_VGND_c_59_n N_VGND_c_60_n VGND
+ N_VGND_c_61_n N_VGND_c_62_n PM_SKY130_FD_SC_LP__INV_1%VGND
cc_1 VNB N_A_M1001_g 0.00750016f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_2 VNB A 0.0203343f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_20_n 0.0431243f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.375
cc_4 VNB N_A_c_21_n 0.0243431f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=1.21
cc_5 VNB N_VPWR_c_36_n 0.0442671f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=1.21
cc_6 VNB N_Y_c_49_n 0.0634045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_VGND_c_59_n 0.0108742f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.54
cc_8 VNB N_VGND_c_60_n 0.0345158f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_9 VNB N_VGND_c_61_n 0.0154464f $X=-0.19 $Y=-0.245 $X2=0.372 $Y2=1.375
cc_10 VNB N_VGND_c_62_n 0.0914566f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.375
cc_11 VPB N_A_M1001_g 0.0285014f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_12 VPB A 0.00735577f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_13 VPB N_VPWR_c_37_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.54
cc_14 VPB N_VPWR_c_38_n 0.0484529f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_15 VPB N_VPWR_c_39_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0.35 $Y2=1.375
cc_16 VPB N_VPWR_c_36_n 0.0437929f $X=-0.19 $Y=1.655 $X2=0.372 $Y2=1.21
cc_17 VPB N_Y_c_49_n 0.0573297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 N_A_M1001_g N_VPWR_c_38_n 0.0224724f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_19 A N_VPWR_c_38_n 0.026915f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_20 N_A_c_20_n N_VPWR_c_38_n 9.85169e-19 $X=0.35 $Y=1.375 $X2=0 $Y2=0
cc_21 N_A_M1001_g N_VPWR_c_39_n 0.00486043f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_22 N_A_M1001_g N_VPWR_c_36_n 0.00917987f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_23 A N_Y_c_49_n 0.0422022f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_24 N_A_c_21_n N_Y_c_49_n 0.0267988f $X=0.372 $Y=1.21 $X2=0 $Y2=0
cc_25 A N_VGND_c_60_n 0.0259278f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_26 N_A_c_20_n N_VGND_c_60_n 0.00160808f $X=0.35 $Y=1.375 $X2=0 $Y2=0
cc_27 N_A_c_21_n N_VGND_c_60_n 0.0179048f $X=0.372 $Y=1.21 $X2=0 $Y2=0
cc_28 N_A_c_21_n N_VGND_c_61_n 0.00465098f $X=0.372 $Y=1.21 $X2=0 $Y2=0
cc_29 N_A_c_21_n N_VGND_c_62_n 0.00905258f $X=0.372 $Y=1.21 $X2=0 $Y2=0
cc_30 N_VPWR_c_36_n N_Y_M1001_d 0.00371702f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_31 N_VPWR_c_39_n N_Y_c_49_n 0.018528f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_32 N_VPWR_c_36_n N_Y_c_49_n 0.0104192f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_33 N_Y_c_49_n N_VGND_c_60_n 0.0296165f $X=0.7 $Y=0.42 $X2=0 $Y2=0
cc_34 N_Y_c_49_n N_VGND_c_61_n 0.019212f $X=0.7 $Y=0.42 $X2=0 $Y2=0
cc_35 N_Y_c_49_n N_VGND_c_62_n 0.0104192f $X=0.7 $Y=0.42 $X2=0 $Y2=0
