* File: sky130_fd_sc_lp__and4_0.pxi.spice
* Created: Fri Aug 28 10:07:23 2020
* 
x_PM_SKY130_FD_SC_LP__AND4_0%A N_A_M1009_g N_A_M1002_g N_A_c_71_n N_A_c_72_n
+ N_A_c_73_n A A A A N_A_c_75_n PM_SKY130_FD_SC_LP__AND4_0%A
x_PM_SKY130_FD_SC_LP__AND4_0%B N_B_M1000_g N_B_M1003_g N_B_c_109_n N_B_c_114_n B
+ B N_B_c_111_n PM_SKY130_FD_SC_LP__AND4_0%B
x_PM_SKY130_FD_SC_LP__AND4_0%C N_C_M1006_g N_C_c_152_n N_C_M1007_g N_C_c_157_n C
+ C N_C_c_154_n PM_SKY130_FD_SC_LP__AND4_0%C
x_PM_SKY130_FD_SC_LP__AND4_0%D N_D_c_191_n N_D_M1008_g N_D_M1004_g N_D_c_192_n
+ N_D_c_197_n N_D_c_198_n N_D_c_193_n D D D N_D_c_195_n
+ PM_SKY130_FD_SC_LP__AND4_0%D
x_PM_SKY130_FD_SC_LP__AND4_0%A_84_58# N_A_84_58#_M1002_s N_A_84_58#_M1009_d
+ N_A_84_58#_M1007_d N_A_84_58#_M1005_g N_A_84_58#_M1001_g N_A_84_58#_c_241_n
+ N_A_84_58#_c_242_n N_A_84_58#_c_243_n N_A_84_58#_c_244_n N_A_84_58#_c_245_n
+ N_A_84_58#_c_253_n N_A_84_58#_c_246_n N_A_84_58#_c_254_n N_A_84_58#_c_255_n
+ N_A_84_58#_c_247_n N_A_84_58#_c_248_n N_A_84_58#_c_256_n N_A_84_58#_c_249_n
+ N_A_84_58#_c_250_n PM_SKY130_FD_SC_LP__AND4_0%A_84_58#
x_PM_SKY130_FD_SC_LP__AND4_0%VPWR N_VPWR_M1009_s N_VPWR_M1000_d N_VPWR_M1004_d
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n VPWR
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_335_n N_VPWR_c_344_n
+ N_VPWR_c_345_n PM_SKY130_FD_SC_LP__AND4_0%VPWR
x_PM_SKY130_FD_SC_LP__AND4_0%X N_X_M1005_d N_X_M1001_d X X X X X X X N_X_c_374_n
+ X PM_SKY130_FD_SC_LP__AND4_0%X
x_PM_SKY130_FD_SC_LP__AND4_0%VGND N_VGND_M1008_d VGND N_VGND_c_391_n
+ N_VGND_c_392_n N_VGND_c_393_n PM_SKY130_FD_SC_LP__AND4_0%VGND
cc_1 VNB N_A_M1009_g 0.00689828f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.6
cc_2 VNB N_A_c_71_n 0.0204222f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.82
cc_3 VNB N_A_c_72_n 0.038107f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.97
cc_4 VNB N_A_c_73_n 0.0307127f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.51
cc_5 VNB A 0.0338228f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A_c_75_n 0.028745f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.005
cc_7 VNB N_B_M1003_g 0.0336799f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.5
cc_8 VNB N_B_c_109_n 0.0173378f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.28
cc_9 VNB B 0.00551613f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_10 VNB N_B_c_111_n 0.0152537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_M1006_g 0.0324509f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.6
cc_12 VNB N_C_c_152_n 0.0201769f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.5
cc_13 VNB C 0.00533177f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.51
cc_14 VNB N_C_c_154_n 0.0171358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D_c_191_n 0.0177096f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.51
cc_16 VNB N_D_c_192_n 0.0225528f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.51
cc_17 VNB N_D_c_193_n 0.0332711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB D 0.00477914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_c_195_n 0.01222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_84_58#_M1001_g 0.0101266f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A_84_58#_c_241_n 0.0230014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_84_58#_c_242_n 0.0184424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_84_58#_c_243_n 0.0206873f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.005
cc_24 VNB N_A_84_58#_c_244_n 0.00377099f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.005
cc_25 VNB N_A_84_58#_c_245_n 0.00466697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_84_58#_c_246_n 0.0394855f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.665
cc_27 VNB N_A_84_58#_c_247_n 0.0135833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_84_58#_c_248_n 3.35665e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_84_58#_c_249_n 0.00548583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_84_58#_c_250_n 0.0290753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_335_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 0.0555347f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.97
cc_33 VNB N_X_c_374_n 0.0218129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_391_n 0.0765092f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.5
cc_35 VNB N_VGND_c_392_n 0.0239462f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_36 VNB N_VGND_c_393_n 0.206265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A_M1009_g 0.0533588f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.6
cc_38 VPB A 0.0376646f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_39 VPB N_B_M1000_g 0.037576f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.6
cc_40 VPB N_B_c_109_n 0.00366642f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.28
cc_41 VPB N_B_c_114_n 0.0152454f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.51
cc_42 VPB B 0.00395875f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_43 VPB N_C_c_152_n 5.87678e-19 $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.5
cc_44 VPB N_C_M1007_g 0.0409041f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.82
cc_45 VPB N_C_c_157_n 0.0171358f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.28
cc_46 VPB C 0.00388993f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.51
cc_47 VPB N_D_M1004_g 0.0230948f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.5
cc_48 VPB N_D_c_197_n 0.0281958f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_49 VPB N_D_c_198_n 0.0317735f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_50 VPB N_D_c_195_n 0.00523943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_84_58#_M1001_g 0.0609635f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_52 VPB N_A_84_58#_c_245_n 0.00300855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_84_58#_c_253_n 0.00219752f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.295
cc_54 VPB N_A_84_58#_c_254_n 0.012974f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=2.035
cc_55 VPB N_A_84_58#_c_255_n 0.00254375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_84_58#_c_256_n 0.00465237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_336_n 0.0139101f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.97
cc_58 VPB N_VPWR_c_337_n 0.0360731f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.51
cc_59 VPB N_VPWR_c_338_n 0.0138058f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_60 VPB N_VPWR_c_339_n 0.0319458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_340_n 0.0177099f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.925
cc_62 VPB N_VPWR_c_341_n 0.0180304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_342_n 0.0202963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_335_n 0.0706069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_344_n 0.00574453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_345_n 0.0129576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB X 0.0409371f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.97
cc_68 VPB X 0.0240689f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_69 VPB X 0.0160697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 N_A_M1009_g N_B_M1000_g 0.0273252f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_71 N_A_c_71_n N_B_M1003_g 0.0508524f $X=0.51 $Y=0.82 $X2=0 $Y2=0
cc_72 N_A_c_75_n N_B_M1003_g 0.00622968f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_73 N_A_c_73_n N_B_c_109_n 0.0129634f $X=0.415 $Y=1.51 $X2=0 $Y2=0
cc_74 N_A_M1009_g N_B_c_114_n 0.0129634f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_75 N_A_c_75_n B 7.245e-19 $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_76 N_A_c_75_n N_B_c_111_n 0.0129634f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_77 N_A_c_71_n N_A_84_58#_c_244_n 0.00615788f $X=0.51 $Y=0.82 $X2=0 $Y2=0
cc_78 N_A_M1009_g N_A_84_58#_c_245_n 0.00967451f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_79 N_A_c_73_n N_A_84_58#_c_245_n 0.00523435f $X=0.415 $Y=1.51 $X2=0 $Y2=0
cc_80 A N_A_84_58#_c_245_n 0.0788652f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A_c_75_n N_A_84_58#_c_245_n 0.00742513f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_82 N_A_M1009_g N_A_84_58#_c_253_n 0.00344968f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_83 N_A_c_72_n N_A_84_58#_c_246_n 0.00387262f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_84 N_A_c_71_n N_A_84_58#_c_247_n 0.00907807f $X=0.51 $Y=0.82 $X2=0 $Y2=0
cc_85 N_A_c_72_n N_A_84_58#_c_247_n 0.00949984f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_86 A N_A_84_58#_c_247_n 0.00439431f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A_c_72_n N_A_84_58#_c_248_n 0.00981017f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_88 A N_A_84_58#_c_248_n 0.0127464f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A_c_75_n N_A_84_58#_c_248_n 6.42966e-19 $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_90 N_A_M1009_g N_A_84_58#_c_256_n 0.00859156f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_91 A N_A_84_58#_c_256_n 0.0130631f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A_M1009_g N_VPWR_c_337_n 0.00421835f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_93 A N_VPWR_c_337_n 0.0185935f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_94 N_A_M1009_g N_VPWR_c_340_n 0.00475172f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_95 N_A_M1009_g N_VPWR_c_335_n 0.00499434f $X=0.57 $Y=2.6 $X2=0 $Y2=0
cc_96 N_A_c_71_n N_VGND_c_391_n 0.00401104f $X=0.51 $Y=0.82 $X2=0 $Y2=0
cc_97 N_A_c_71_n N_VGND_c_393_n 0.00580887f $X=0.51 $Y=0.82 $X2=0 $Y2=0
cc_98 N_A_c_72_n N_VGND_c_393_n 0.00501246f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_99 A N_VGND_c_393_n 0.0110114f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_100 N_B_M1003_g N_C_M1006_g 0.0270232f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_101 B N_C_M1006_g 0.0054017f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B_c_109_n N_C_c_152_n 0.0270232f $X=1.03 $Y=1.715 $X2=0 $Y2=0
cc_103 N_B_M1000_g N_C_M1007_g 0.0233381f $X=1 $Y=2.6 $X2=0 $Y2=0
cc_104 N_B_c_114_n N_C_c_157_n 0.0270232f $X=1.03 $Y=1.88 $X2=0 $Y2=0
cc_105 N_B_M1003_g C 5.48108e-19 $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_106 B C 0.0535368f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B_c_111_n N_C_c_154_n 0.0270232f $X=1.03 $Y=1.375 $X2=0 $Y2=0
cc_108 B D 0.0014156f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B_M1003_g N_A_84_58#_c_244_n 9.49655e-19 $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_110 N_B_M1000_g N_A_84_58#_c_245_n 0.00379347f $X=1 $Y=2.6 $X2=0 $Y2=0
cc_111 N_B_M1003_g N_A_84_58#_c_245_n 0.00341147f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_112 B N_A_84_58#_c_245_n 0.0549406f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B_c_111_n N_A_84_58#_c_245_n 0.00425229f $X=1.03 $Y=1.375 $X2=0 $Y2=0
cc_114 N_B_M1000_g N_A_84_58#_c_253_n 0.00190949f $X=1 $Y=2.6 $X2=0 $Y2=0
cc_115 N_B_M1003_g N_A_84_58#_c_246_n 0.0109865f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_116 B N_A_84_58#_c_246_n 0.0316778f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B_c_111_n N_A_84_58#_c_246_n 0.00376368f $X=1.03 $Y=1.375 $X2=0 $Y2=0
cc_118 N_B_M1000_g N_A_84_58#_c_254_n 0.0172878f $X=1 $Y=2.6 $X2=0 $Y2=0
cc_119 N_B_c_114_n N_A_84_58#_c_254_n 0.00123286f $X=1.03 $Y=1.88 $X2=0 $Y2=0
cc_120 B N_A_84_58#_c_254_n 0.0303744f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_121 N_B_M1003_g N_A_84_58#_c_247_n 0.00193367f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_122 N_B_c_114_n N_A_84_58#_c_256_n 0.00236819f $X=1.03 $Y=1.88 $X2=0 $Y2=0
cc_123 N_B_M1000_g N_VPWR_c_338_n 0.00207739f $X=1 $Y=2.6 $X2=0 $Y2=0
cc_124 N_B_M1000_g N_VPWR_c_340_n 0.00475172f $X=1 $Y=2.6 $X2=0 $Y2=0
cc_125 N_B_M1000_g N_VPWR_c_335_n 0.00499434f $X=1 $Y=2.6 $X2=0 $Y2=0
cc_126 N_B_M1003_g N_VGND_c_391_n 0.00531318f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_127 N_B_M1003_g N_VGND_c_393_n 0.00567101f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_128 N_C_M1006_g N_D_c_191_n 0.0509931f $X=1.48 $Y=0.5 $X2=-0.19 $Y2=-0.245
cc_129 C N_D_c_192_n 4.21152e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_C_M1007_g N_D_c_197_n 0.00681918f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_131 N_C_c_157_n N_D_c_197_n 0.0113687f $X=1.58 $Y=1.84 $X2=0 $Y2=0
cc_132 N_C_M1007_g N_D_c_198_n 0.0192115f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_133 N_C_M1006_g N_D_c_193_n 0.00666751f $X=1.48 $Y=0.5 $X2=0 $Y2=0
cc_134 C N_D_c_193_n 0.00380152f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_135 N_C_c_154_n N_D_c_193_n 0.0113687f $X=1.59 $Y=1.335 $X2=0 $Y2=0
cc_136 N_C_M1007_g D 0.00126181f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_137 C D 0.0528188f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_138 N_C_c_154_n D 7.38804e-19 $X=1.59 $Y=1.335 $X2=0 $Y2=0
cc_139 N_C_c_152_n N_D_c_195_n 0.0113687f $X=1.58 $Y=1.665 $X2=0 $Y2=0
cc_140 N_C_M1006_g N_A_84_58#_c_246_n 0.0141872f $X=1.48 $Y=0.5 $X2=0 $Y2=0
cc_141 C N_A_84_58#_c_246_n 0.0244333f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_C_c_154_n N_A_84_58#_c_246_n 0.00137591f $X=1.59 $Y=1.335 $X2=0 $Y2=0
cc_143 N_C_M1007_g N_A_84_58#_c_254_n 0.0194724f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_144 N_C_c_157_n N_A_84_58#_c_254_n 0.00150963f $X=1.58 $Y=1.84 $X2=0 $Y2=0
cc_145 C N_A_84_58#_c_254_n 0.0230831f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_C_M1007_g N_A_84_58#_c_255_n 0.00188399f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_147 N_C_M1007_g N_VPWR_c_338_n 0.0020518f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_148 N_C_M1007_g N_VPWR_c_341_n 0.00475172f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_149 N_C_M1007_g N_VPWR_c_335_n 0.00499434f $X=1.48 $Y=2.6 $X2=0 $Y2=0
cc_150 N_C_M1006_g N_VGND_c_391_n 0.00807867f $X=1.48 $Y=0.5 $X2=0 $Y2=0
cc_151 N_C_M1006_g N_VGND_c_393_n 0.00567101f $X=1.48 $Y=0.5 $X2=0 $Y2=0
cc_152 N_D_M1004_g N_A_84_58#_M1001_g 0.00410178f $X=1.91 $Y=2.6 $X2=0 $Y2=0
cc_153 N_D_c_193_n N_A_84_58#_M1001_g 0.00114647f $X=2.16 $Y=1.56 $X2=0 $Y2=0
cc_154 D N_A_84_58#_M1001_g 0.00330838f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_155 N_D_c_195_n N_A_84_58#_M1001_g 0.0231609f $X=2.16 $Y=1.725 $X2=0 $Y2=0
cc_156 N_D_c_191_n N_A_84_58#_c_241_n 0.00498624f $X=1.84 $Y=0.81 $X2=0 $Y2=0
cc_157 N_D_c_192_n N_A_84_58#_c_241_n 0.0023665f $X=2.07 $Y=0.885 $X2=0 $Y2=0
cc_158 N_D_c_193_n N_A_84_58#_c_242_n 0.0023665f $X=2.16 $Y=1.56 $X2=0 $Y2=0
cc_159 N_D_c_192_n N_A_84_58#_c_246_n 0.0160692f $X=2.07 $Y=0.885 $X2=0 $Y2=0
cc_160 N_D_c_193_n N_A_84_58#_c_246_n 0.00332034f $X=2.16 $Y=1.56 $X2=0 $Y2=0
cc_161 D N_A_84_58#_c_246_n 0.0264685f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_162 N_D_c_195_n N_A_84_58#_c_246_n 5.44562e-19 $X=2.16 $Y=1.725 $X2=0 $Y2=0
cc_163 N_D_c_198_n N_A_84_58#_c_254_n 0.00320636f $X=2.08 $Y=2.23 $X2=0 $Y2=0
cc_164 D N_A_84_58#_c_254_n 0.0126104f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_165 N_D_M1004_g N_A_84_58#_c_255_n 0.00322853f $X=1.91 $Y=2.6 $X2=0 $Y2=0
cc_166 N_D_c_193_n N_A_84_58#_c_249_n 0.00129416f $X=2.16 $Y=1.56 $X2=0 $Y2=0
cc_167 D N_A_84_58#_c_249_n 0.0197766f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_168 N_D_c_193_n N_A_84_58#_c_250_n 0.0139065f $X=2.16 $Y=1.56 $X2=0 $Y2=0
cc_169 D N_A_84_58#_c_250_n 0.00265045f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_170 N_D_M1004_g N_VPWR_c_339_n 0.00333812f $X=1.91 $Y=2.6 $X2=0 $Y2=0
cc_171 N_D_c_198_n N_VPWR_c_339_n 0.00912052f $X=2.08 $Y=2.23 $X2=0 $Y2=0
cc_172 D N_VPWR_c_339_n 0.0292419f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_D_M1004_g N_VPWR_c_341_n 0.00475172f $X=1.91 $Y=2.6 $X2=0 $Y2=0
cc_174 N_D_M1004_g N_VPWR_c_335_n 0.00499434f $X=1.91 $Y=2.6 $X2=0 $Y2=0
cc_175 D X 0.0201635f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_176 N_D_c_191_n N_VGND_c_391_n 0.0170449f $X=1.84 $Y=0.81 $X2=0 $Y2=0
cc_177 N_D_c_192_n N_VGND_c_391_n 0.00557411f $X=2.07 $Y=0.885 $X2=0 $Y2=0
cc_178 N_D_c_191_n N_VGND_c_393_n 0.00419263f $X=1.84 $Y=0.81 $X2=0 $Y2=0
cc_179 N_A_84_58#_c_254_n N_VPWR_c_338_n 0.0212864f $X=1.555 $Y=2.162 $X2=0
+ $Y2=0
cc_180 N_A_84_58#_M1001_g N_VPWR_c_339_n 0.00555287f $X=2.745 $Y=2.71 $X2=0
+ $Y2=0
cc_181 N_A_84_58#_c_255_n N_VPWR_c_339_n 7.80401e-19 $X=1.695 $Y=2.575 $X2=0
+ $Y2=0
cc_182 N_A_84_58#_c_253_n N_VPWR_c_340_n 0.00484442f $X=0.785 $Y=2.6 $X2=0 $Y2=0
cc_183 N_A_84_58#_c_255_n N_VPWR_c_341_n 0.00466515f $X=1.695 $Y=2.575 $X2=0
+ $Y2=0
cc_184 N_A_84_58#_M1001_g N_VPWR_c_342_n 0.00520454f $X=2.745 $Y=2.71 $X2=0
+ $Y2=0
cc_185 N_A_84_58#_M1001_g N_VPWR_c_335_n 0.01134f $X=2.745 $Y=2.71 $X2=0 $Y2=0
cc_186 N_A_84_58#_c_253_n N_VPWR_c_335_n 0.00824747f $X=0.785 $Y=2.6 $X2=0 $Y2=0
cc_187 N_A_84_58#_c_255_n N_VPWR_c_335_n 0.00840561f $X=1.695 $Y=2.575 $X2=0
+ $Y2=0
cc_188 N_A_84_58#_M1001_g X 0.0238502f $X=2.745 $Y=2.71 $X2=0 $Y2=0
cc_189 N_A_84_58#_c_241_n X 0.00494523f $X=2.715 $Y=0.82 $X2=0 $Y2=0
cc_190 N_A_84_58#_c_242_n X 0.0167595f $X=2.715 $Y=0.97 $X2=0 $Y2=0
cc_191 N_A_84_58#_c_249_n X 0.0523937f $X=2.73 $Y=0.985 $X2=0 $Y2=0
cc_192 N_A_84_58#_c_242_n N_X_c_374_n 0.00427806f $X=2.715 $Y=0.97 $X2=0 $Y2=0
cc_193 N_A_84_58#_c_249_n N_X_c_374_n 0.00771709f $X=2.73 $Y=0.985 $X2=0 $Y2=0
cc_194 N_A_84_58#_M1001_g X 9.17742e-19 $X=2.745 $Y=2.71 $X2=0 $Y2=0
cc_195 N_A_84_58#_c_241_n N_VGND_c_391_n 0.00410318f $X=2.715 $Y=0.82 $X2=0
+ $Y2=0
cc_196 N_A_84_58#_c_246_n N_VGND_c_391_n 0.0454452f $X=2.565 $Y=0.905 $X2=0
+ $Y2=0
cc_197 N_A_84_58#_c_247_n N_VGND_c_391_n 0.0168373f $X=0.695 $Y=0.495 $X2=0
+ $Y2=0
cc_198 N_A_84_58#_c_241_n N_VGND_c_392_n 0.00531318f $X=2.715 $Y=0.82 $X2=0
+ $Y2=0
cc_199 N_A_84_58#_c_241_n N_VGND_c_393_n 0.00677426f $X=2.715 $Y=0.82 $X2=0
+ $Y2=0
cc_200 N_A_84_58#_c_246_n N_VGND_c_393_n 0.0386806f $X=2.565 $Y=0.905 $X2=0
+ $Y2=0
cc_201 N_A_84_58#_c_247_n N_VGND_c_393_n 0.0143025f $X=0.695 $Y=0.495 $X2=0
+ $Y2=0
cc_202 N_A_84_58#_c_249_n N_VGND_c_393_n 0.0044267f $X=2.73 $Y=0.985 $X2=0 $Y2=0
cc_203 N_VPWR_c_342_n X 0.0253918f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_335_n X 0.0165413f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_c_339_n X 0.0312803f $X=2.53 $Y=2.545 $X2=0 $Y2=0
cc_206 N_X_c_374_n N_VGND_c_392_n 0.0265126f $X=3.13 $Y=0.485 $X2=0 $Y2=0
cc_207 N_X_c_374_n N_VGND_c_393_n 0.0213116f $X=3.13 $Y=0.485 $X2=0 $Y2=0
