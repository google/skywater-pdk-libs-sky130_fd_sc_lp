* File: sky130_fd_sc_lp__nand3_2.pxi.spice
* Created: Wed Sep  2 10:04:16 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3_2%A N_A_c_62_n N_A_M1009_g N_A_M1004_g N_A_c_64_n
+ N_A_c_65_n N_A_M1010_g N_A_M1008_g N_A_c_67_n A A N_A_c_69_n
+ PM_SKY130_FD_SC_LP__NAND3_2%A
x_PM_SKY130_FD_SC_LP__NAND3_2%B N_B_M1002_g N_B_M1005_g N_B_M1006_g N_B_M1003_g
+ N_B_c_116_n N_B_c_109_n N_B_c_110_n N_B_c_111_n B B B N_B_c_112_n N_B_c_113_n
+ N_B_c_127_p B PM_SKY130_FD_SC_LP__NAND3_2%B
x_PM_SKY130_FD_SC_LP__NAND3_2%C N_C_M1000_g N_C_M1001_g N_C_M1011_g N_C_M1007_g
+ C N_C_c_194_n PM_SKY130_FD_SC_LP__NAND3_2%C
x_PM_SKY130_FD_SC_LP__NAND3_2%VPWR N_VPWR_M1004_s N_VPWR_M1008_s N_VPWR_M1001_d
+ N_VPWR_M1006_d N_VPWR_c_244_n N_VPWR_c_245_n N_VPWR_c_246_n N_VPWR_c_247_n
+ N_VPWR_c_248_n N_VPWR_c_249_n VPWR N_VPWR_c_250_n N_VPWR_c_251_n
+ N_VPWR_c_252_n N_VPWR_c_253_n N_VPWR_c_254_n N_VPWR_c_243_n
+ PM_SKY130_FD_SC_LP__NAND3_2%VPWR
x_PM_SKY130_FD_SC_LP__NAND3_2%Y N_Y_M1009_d N_Y_M1004_d N_Y_M1005_s N_Y_M1011_s
+ N_Y_c_300_n N_Y_c_309_n N_Y_c_336_n N_Y_c_323_n N_Y_c_325_n N_Y_c_310_n
+ N_Y_c_312_n N_Y_c_326_n N_Y_c_328_n Y PM_SKY130_FD_SC_LP__NAND3_2%Y
x_PM_SKY130_FD_SC_LP__NAND3_2%A_43_65# N_A_43_65#_M1009_s N_A_43_65#_M1010_s
+ N_A_43_65#_M1003_d N_A_43_65#_c_348_n N_A_43_65#_c_349_n N_A_43_65#_c_350_n
+ N_A_43_65#_c_351_n N_A_43_65#_c_352_n N_A_43_65#_c_353_n
+ PM_SKY130_FD_SC_LP__NAND3_2%A_43_65#
x_PM_SKY130_FD_SC_LP__NAND3_2%A_298_65# N_A_298_65#_M1002_s N_A_298_65#_M1007_s
+ N_A_298_65#_c_393_n N_A_298_65#_c_396_n N_A_298_65#_c_397_n
+ N_A_298_65#_c_394_n PM_SKY130_FD_SC_LP__NAND3_2%A_298_65#
x_PM_SKY130_FD_SC_LP__NAND3_2%VGND N_VGND_M1000_d N_VGND_c_422_n VGND
+ N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n
+ PM_SKY130_FD_SC_LP__NAND3_2%VGND
cc_1 VNB N_A_c_62_n 0.0206343f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.275
cc_2 VNB N_A_M1004_g 0.00302368f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_3 VNB N_A_c_64_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.35
cc_4 VNB N_A_c_65_n 0.0159594f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.275
cc_5 VNB N_A_M1008_g 0.0103887f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_6 VNB N_A_c_67_n 0.00515988f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_7 VNB A 0.0248754f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_c_69_n 0.0458272f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.44
cc_9 VNB N_B_M1002_g 0.0204456f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.745
cc_10 VNB N_B_M1003_g 0.0265786f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_11 VNB N_B_c_109_n 0.00284919f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_B_c_110_n 0.0086712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_111_n 0.0302714f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_14 VNB N_B_c_112_n 0.0239558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_113_n 0.00289146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C_M1000_g 0.021488f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.745
cc_17 VNB N_C_M1007_g 0.0210196f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_18 VNB C 0.00152431f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_19 VNB N_C_c_194_n 0.0381655f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_20 VNB N_VPWR_c_243_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_300_n 0.00222248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_43_65#_c_348_n 0.0233564f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.745
cc_23 VNB N_A_43_65#_c_349_n 0.00484211f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_24 VNB N_A_43_65#_c_350_n 0.00928796f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_25 VNB N_A_43_65#_c_351_n 0.0228962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_43_65#_c_352_n 0.00246665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_43_65#_c_353_n 0.0316355f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_28 VNB N_A_298_65#_c_393_n 0.00245183f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.35
cc_29 VNB N_A_298_65#_c_394_n 0.00214535f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_30 VNB N_VGND_c_422_n 0.00809655f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_31 VNB N_VGND_c_423_n 0.0507622f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.275
cc_32 VNB N_VGND_c_424_n 0.0296704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_425_n 0.207691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_426_n 0.00632057f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.44
cc_35 VPB N_A_M1004_g 0.0251188f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_36 VPB N_A_M1008_g 0.0194686f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_37 VPB A 0.0100485f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_38 VPB N_B_M1005_g 0.0177081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_B_M1006_g 0.0249717f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.745
cc_40 VPB N_B_c_116_n 0.00145457f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_41 VPB N_B_c_111_n 0.00776298f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.44
cc_42 VPB N_B_c_112_n 0.00635135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_B_c_113_n 0.00251493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_C_M1001_g 0.0186851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_C_M1011_g 0.0192822f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.745
cc_46 VPB C 0.00370347f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.35
cc_47 VPB N_C_c_194_n 0.00622089f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.44
cc_48 VPB N_VPWR_c_244_n 0.0128916f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.425
cc_49 VPB N_VPWR_c_245_n 0.0482589f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_50 VPB N_VPWR_c_246_n 3.19588e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_247_n 0.00228457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_248_n 0.013074f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.44
cc_53 VPB N_VPWR_c_249_n 0.0555199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_250_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_251_n 0.0138364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_252_n 0.0170994f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_253_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_254_n 0.00522677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_243_n 0.050503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_Y_c_300_n 0.00166109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 N_A_c_65_n N_B_M1002_g 0.0202272f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_62 N_A_M1008_g N_B_M1005_g 0.0419717f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A_c_67_n N_B_c_112_n 0.020473f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_64 N_A_M1008_g N_B_c_113_n 0.00445928f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A_M1004_g N_VPWR_c_245_n 0.020423f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_M1008_g N_VPWR_c_245_n 8.25447e-19 $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_67 A N_VPWR_c_245_n 0.0269147f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_c_69_n N_VPWR_c_245_n 0.00156499f $X=0.63 $Y=1.44 $X2=0 $Y2=0
cc_69 N_A_M1004_g N_VPWR_c_246_n 5.5535e-19 $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_M1008_g N_VPWR_c_246_n 0.0093124f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_VPWR_c_250_n 0.00486043f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_72 N_A_M1008_g N_VPWR_c_250_n 0.00564095f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_VPWR_c_243_n 0.00824727f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A_M1008_g N_VPWR_c_243_n 0.00948291f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_75 N_A_c_62_n N_Y_c_300_n 0.0016362f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_76 N_A_c_64_n N_Y_c_300_n 0.0101622f $X=0.91 $Y=1.35 $X2=0 $Y2=0
cc_77 N_A_c_65_n N_Y_c_300_n 0.00318739f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_78 N_A_M1008_g N_Y_c_300_n 0.0147641f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_c_67_n N_Y_c_300_n 0.0026119f $X=0.985 $Y=1.35 $X2=0 $Y2=0
cc_80 A N_Y_c_300_n 0.0420231f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_c_69_n N_Y_c_300_n 0.00522533f $X=0.63 $Y=1.44 $X2=0 $Y2=0
cc_82 N_A_M1008_g N_Y_c_309_n 0.0149388f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_c_62_n N_Y_c_310_n 0.00750987f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_84 N_A_c_65_n N_Y_c_310_n 0.00512809f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_85 N_A_M1008_g N_Y_c_312_n 0.00157824f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_86 A N_A_43_65#_c_348_n 0.0228785f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A_c_69_n N_A_43_65#_c_348_n 0.00169228f $X=0.63 $Y=1.44 $X2=0 $Y2=0
cc_88 N_A_c_62_n N_A_43_65#_c_349_n 0.0125027f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_89 N_A_c_65_n N_A_43_65#_c_349_n 0.0118308f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_90 N_A_c_65_n N_A_43_65#_c_352_n 7.38449e-19 $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_91 N_A_c_62_n N_VGND_c_423_n 0.00302501f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_92 N_A_c_65_n N_VGND_c_423_n 0.00302501f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_93 N_A_c_62_n N_VGND_c_425_n 0.00473131f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_94 N_A_c_65_n N_VGND_c_425_n 0.00435646f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_95 N_B_M1002_g N_C_M1000_g 0.0180218f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_96 N_B_M1005_g N_C_M1001_g 0.0339219f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B_c_113_n N_C_M1001_g 0.00464493f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B_c_127_p N_C_M1001_g 0.0113188f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_99 N_B_M1006_g N_C_M1011_g 0.0209255f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B_c_127_p N_C_M1011_g 0.0137044f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_101 N_B_M1003_g N_C_M1007_g 0.0211296f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_102 N_B_c_116_n C 0.00829151f $X=2.617 $Y=1.92 $X2=0 $Y2=0
cc_103 N_B_c_109_n C 0.0185294f $X=2.745 $Y=1.535 $X2=0 $Y2=0
cc_104 N_B_c_111_n C 2.31952e-19 $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B_c_112_n C 8.66797e-19 $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_106 N_B_c_113_n C 0.0222131f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_107 N_B_c_127_p C 0.0347386f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_108 N_B_c_116_n N_C_c_194_n 0.00337497f $X=2.617 $Y=1.92 $X2=0 $Y2=0
cc_109 N_B_c_109_n N_C_c_194_n 0.00395807f $X=2.745 $Y=1.535 $X2=0 $Y2=0
cc_110 N_B_c_111_n N_C_c_194_n 0.0317876f $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_111 N_B_c_112_n N_C_c_194_n 0.0221004f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_112 N_B_c_113_n N_C_c_194_n 3.10277e-19 $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_113 N_B_c_127_p N_C_c_194_n 8.7831e-19 $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_114 N_B_c_113_n N_VPWR_M1008_s 0.00346286f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_115 N_B_c_127_p N_VPWR_M1001_d 0.00431729f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_116 N_B_M1005_g N_VPWR_c_246_n 0.00935629f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B_M1005_g N_VPWR_c_247_n 5.55001e-19 $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B_M1006_g N_VPWR_c_249_n 0.00734928f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B_c_116_n N_VPWR_c_249_n 0.00451364f $X=2.617 $Y=1.92 $X2=0 $Y2=0
cc_120 N_B_c_110_n N_VPWR_c_249_n 0.0109957f $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_121 N_B_c_111_n N_VPWR_c_249_n 0.00333442f $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_122 N_B_M1005_g N_VPWR_c_251_n 0.00564095f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B_M1006_g N_VPWR_c_252_n 0.0054895f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B_M1005_g N_VPWR_c_243_n 0.00950825f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B_M1006_g N_VPWR_c_243_n 0.0107983f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B_c_113_n N_Y_M1005_s 0.00178522f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_127 N_B_c_127_p N_Y_M1005_s 0.00533721f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_128 N_B_c_116_n N_Y_M1011_s 0.00183822f $X=2.617 $Y=1.92 $X2=0 $Y2=0
cc_129 N_B_M1002_g N_Y_c_300_n 5.25854e-19 $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_130 N_B_M1005_g N_Y_c_300_n 0.00113361f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B_c_112_n N_Y_c_300_n 6.22723e-19 $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_132 N_B_c_113_n N_Y_c_300_n 0.0431982f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_133 N_B_M1005_g N_Y_c_309_n 0.0129889f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B_c_112_n N_Y_c_309_n 2.5744e-19 $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_135 N_B_c_113_n N_Y_c_309_n 0.0282031f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_136 N_B_M1006_g N_Y_c_323_n 0.00247149f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B_c_116_n N_Y_c_323_n 0.0169838f $X=2.617 $Y=1.92 $X2=0 $Y2=0
cc_138 N_B_M1006_g N_Y_c_325_n 0.00785269f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B_c_113_n N_Y_c_326_n 0.00108369f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_140 N_B_c_127_p N_Y_c_326_n 0.0125855f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_141 N_B_c_127_p N_Y_c_328_n 0.0368552f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_142 N_B_M1002_g N_A_43_65#_c_349_n 8.65746e-19 $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_143 N_B_M1002_g N_A_43_65#_c_351_n 0.0138505f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_144 N_B_M1003_g N_A_43_65#_c_351_n 0.0139823f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_145 N_B_c_109_n N_A_43_65#_c_351_n 0.0212964f $X=2.745 $Y=1.535 $X2=0 $Y2=0
cc_146 N_B_c_110_n N_A_43_65#_c_351_n 0.022193f $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_147 N_B_c_111_n N_A_43_65#_c_351_n 0.0048013f $X=2.885 $Y=1.51 $X2=0 $Y2=0
cc_148 N_B_c_112_n N_A_43_65#_c_351_n 0.0035112f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_149 N_B_c_113_n N_A_43_65#_c_351_n 0.022136f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_150 N_B_c_127_p N_A_43_65#_c_351_n 0.00841499f $X=2.49 $Y=2.02 $X2=0 $Y2=0
cc_151 N_B_c_112_n N_A_43_65#_c_352_n 0.00115454f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_152 N_B_c_113_n N_A_43_65#_c_352_n 0.0194095f $X=1.435 $Y=1.51 $X2=0 $Y2=0
cc_153 N_B_M1003_g N_A_43_65#_c_353_n 0.00354556f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_154 N_B_M1002_g N_A_298_65#_c_393_n 0.00450378f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_155 N_B_M1003_g N_A_298_65#_c_396_n 0.00215054f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_156 N_B_M1002_g N_A_298_65#_c_397_n 0.00149101f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_157 N_B_M1003_g N_A_298_65#_c_394_n 0.00618917f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_158 N_B_M1002_g N_VGND_c_423_n 0.00494414f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_159 N_B_M1003_g N_VGND_c_424_n 0.0046877f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_160 N_B_M1002_g N_VGND_c_425_n 0.00977655f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_161 N_B_M1003_g N_VGND_c_425_n 0.00939295f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_162 N_C_M1001_g N_VPWR_c_246_n 5.63047e-19 $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_163 N_C_M1001_g N_VPWR_c_247_n 0.00842884f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_164 N_C_M1011_g N_VPWR_c_247_n 0.00242764f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_165 N_C_M1001_g N_VPWR_c_251_n 0.00564095f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_166 N_C_M1011_g N_VPWR_c_252_n 0.00585385f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_167 N_C_M1001_g N_VPWR_c_243_n 0.0052092f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_168 N_C_M1011_g N_VPWR_c_243_n 0.0063579f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_169 N_C_M1001_g N_Y_c_328_n 0.0110918f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_170 N_C_M1011_g N_Y_c_328_n 0.0111898f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_171 N_C_M1000_g N_A_43_65#_c_351_n 0.0113031f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_172 N_C_M1007_g N_A_43_65#_c_351_n 0.0127204f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_173 C N_A_43_65#_c_351_n 0.0377242f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_174 N_C_c_194_n N_A_43_65#_c_351_n 0.00572325f $X=2.365 $Y=1.51 $X2=0 $Y2=0
cc_175 N_C_M1000_g N_A_298_65#_c_393_n 0.00628737f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_176 N_C_M1007_g N_A_298_65#_c_393_n 5.71435e-19 $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_177 N_C_M1000_g N_A_298_65#_c_396_n 0.0105222f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_178 N_C_M1007_g N_A_298_65#_c_396_n 0.010086f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_179 N_C_M1000_g N_A_298_65#_c_394_n 4.23006e-19 $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_180 N_C_M1007_g N_A_298_65#_c_394_n 0.00705285f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_181 N_C_M1000_g N_VGND_c_422_n 0.00240631f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_182 N_C_M1007_g N_VGND_c_422_n 0.00415568f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_183 N_C_M1000_g N_VGND_c_423_n 0.00367927f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_184 N_C_M1007_g N_VGND_c_424_n 0.0035973f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_185 N_C_M1000_g N_VGND_c_425_n 0.00513392f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_186 N_C_M1007_g N_VGND_c_425_n 0.00506374f $X=2.435 $Y=0.745 $X2=0 $Y2=0
cc_187 N_VPWR_c_243_n N_Y_M1004_d 0.00467071f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_c_243_n N_Y_M1005_s 0.00325643f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_189 N_VPWR_c_243_n N_Y_M1011_s 0.00232041f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_190 N_VPWR_M1008_s N_Y_c_309_n 0.00433339f $X=1.06 $Y=1.835 $X2=0 $Y2=0
cc_191 N_VPWR_c_246_n N_Y_c_309_n 0.017285f $X=1.22 $Y=2.755 $X2=0 $Y2=0
cc_192 N_VPWR_c_251_n N_Y_c_336_n 0.0138717f $X=1.955 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_243_n N_Y_c_336_n 0.00886411f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_252_n N_Y_c_325_n 0.0167525f $X=2.915 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_243_n N_Y_c_325_n 0.0110138f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_250_n N_Y_c_312_n 0.0131621f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_243_n N_Y_c_312_n 0.00808656f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_M1001_d N_Y_c_328_n 0.00445762f $X=1.96 $Y=1.835 $X2=0 $Y2=0
cc_199 N_VPWR_c_247_n N_Y_c_328_n 0.0176325f $X=2.12 $Y=2.785 $X2=0 $Y2=0
cc_200 N_VPWR_c_243_n N_Y_c_328_n 0.01072f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_249_n N_A_43_65#_c_351_n 0.00505244f $X=3.01 $Y=1.98 $X2=0 $Y2=0
cc_202 N_Y_M1009_d N_A_43_65#_c_349_n 0.00176461f $X=0.63 $Y=0.325 $X2=0 $Y2=0
cc_203 N_Y_c_310_n N_A_43_65#_c_349_n 0.015935f $X=0.77 $Y=0.68 $X2=0 $Y2=0
cc_204 N_Y_c_300_n N_A_43_65#_c_352_n 0.0103283f $X=0.77 $Y=1.96 $X2=0 $Y2=0
cc_205 N_A_43_65#_c_351_n N_A_298_65#_M1002_s 0.00218982f $X=2.985 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_206 N_A_43_65#_c_351_n N_A_298_65#_M1007_s 0.00176461f $X=2.985 $Y=1.17 $X2=0
+ $Y2=0
cc_207 N_A_43_65#_c_349_n N_A_298_65#_c_393_n 0.00709621f $X=1.105 $Y=0.34 $X2=0
+ $Y2=0
cc_208 N_A_43_65#_c_351_n N_A_298_65#_c_396_n 0.0561298f $X=2.985 $Y=1.17 $X2=0
+ $Y2=0
cc_209 N_A_43_65#_c_351_n N_A_298_65#_c_397_n 0.0173303f $X=2.985 $Y=1.17 $X2=0
+ $Y2=0
cc_210 N_A_43_65#_c_353_n N_A_298_65#_c_394_n 0.0172348f $X=3.08 $Y=0.47 $X2=0
+ $Y2=0
cc_211 N_A_43_65#_c_351_n N_VGND_M1000_d 0.00322255f $X=2.985 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_212 N_A_43_65#_c_349_n N_VGND_c_422_n 9.92717e-19 $X=1.105 $Y=0.34 $X2=0
+ $Y2=0
cc_213 N_A_43_65#_c_349_n N_VGND_c_423_n 0.0572829f $X=1.105 $Y=0.34 $X2=0 $Y2=0
cc_214 N_A_43_65#_c_350_n N_VGND_c_423_n 0.0186386f $X=0.435 $Y=0.34 $X2=0 $Y2=0
cc_215 N_A_43_65#_c_353_n N_VGND_c_424_n 0.0140356f $X=3.08 $Y=0.47 $X2=0 $Y2=0
cc_216 N_A_43_65#_c_349_n N_VGND_c_425_n 0.0319816f $X=1.105 $Y=0.34 $X2=0 $Y2=0
cc_217 N_A_43_65#_c_350_n N_VGND_c_425_n 0.0101082f $X=0.435 $Y=0.34 $X2=0 $Y2=0
cc_218 N_A_43_65#_c_353_n N_VGND_c_425_n 0.00977851f $X=3.08 $Y=0.47 $X2=0 $Y2=0
cc_219 N_A_298_65#_c_396_n N_VGND_M1000_d 0.00608201f $X=2.485 $Y=0.83 $X2=-0.19
+ $Y2=-0.245
cc_220 N_A_298_65#_c_393_n N_VGND_c_422_n 0.0125041f $X=1.65 $Y=0.45 $X2=0 $Y2=0
cc_221 N_A_298_65#_c_396_n N_VGND_c_422_n 0.0224848f $X=2.485 $Y=0.83 $X2=0
+ $Y2=0
cc_222 N_A_298_65#_c_394_n N_VGND_c_422_n 0.0125041f $X=2.65 $Y=0.45 $X2=0 $Y2=0
cc_223 N_A_298_65#_c_393_n N_VGND_c_423_n 0.0196172f $X=1.65 $Y=0.45 $X2=0 $Y2=0
cc_224 N_A_298_65#_c_396_n N_VGND_c_423_n 0.00202826f $X=2.485 $Y=0.83 $X2=0
+ $Y2=0
cc_225 N_A_298_65#_c_396_n N_VGND_c_424_n 0.00191958f $X=2.485 $Y=0.83 $X2=0
+ $Y2=0
cc_226 N_A_298_65#_c_394_n N_VGND_c_424_n 0.0194846f $X=2.65 $Y=0.45 $X2=0 $Y2=0
cc_227 N_A_298_65#_c_393_n N_VGND_c_425_n 0.0124996f $X=1.65 $Y=0.45 $X2=0 $Y2=0
cc_228 N_A_298_65#_c_396_n N_VGND_c_425_n 0.00885632f $X=2.485 $Y=0.83 $X2=0
+ $Y2=0
cc_229 N_A_298_65#_c_394_n N_VGND_c_425_n 0.0123131f $X=2.65 $Y=0.45 $X2=0 $Y2=0
