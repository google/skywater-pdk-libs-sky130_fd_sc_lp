* File: sky130_fd_sc_lp__mux2_0.pxi.spice
* Created: Wed Sep  2 09:59:58 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_0%A_89_200# N_A_89_200#_M1008_d N_A_89_200#_M1005_d
+ N_A_89_200#_M1001_g N_A_89_200#_M1009_g N_A_89_200#_c_87_n N_A_89_200#_c_88_n
+ N_A_89_200#_c_89_n N_A_89_200#_c_90_n N_A_89_200#_c_91_n N_A_89_200#_c_92_n
+ N_A_89_200#_c_93_n N_A_89_200#_c_98_n N_A_89_200#_c_94_n N_A_89_200#_c_100_n
+ N_A_89_200#_c_118_p PM_SKY130_FD_SC_LP__MUX2_0%A_89_200#
x_PM_SKY130_FD_SC_LP__MUX2_0%S N_S_M1002_g N_S_c_165_n N_S_M1004_g N_S_M1007_g
+ N_S_M1000_g N_S_c_167_n N_S_c_168_n N_S_c_174_n N_S_c_175_n N_S_c_176_n
+ N_S_c_177_n N_S_c_178_n N_S_c_179_n N_S_c_180_n N_S_c_181_n N_S_c_182_n S S S
+ N_S_c_185_n N_S_c_170_n PM_SKY130_FD_SC_LP__MUX2_0%S
x_PM_SKY130_FD_SC_LP__MUX2_0%A1 N_A1_M1008_g N_A1_M1006_g N_A1_c_283_n
+ N_A1_c_284_n A1 N_A1_c_285_n N_A1_c_288_n N_A1_c_289_n N_A1_c_286_n
+ PM_SKY130_FD_SC_LP__MUX2_0%A1
x_PM_SKY130_FD_SC_LP__MUX2_0%A0 N_A0_M1005_g N_A0_c_347_n N_A0_c_342_n
+ N_A0_M1003_g N_A0_c_348_n A0 A0 N_A0_c_345_n PM_SKY130_FD_SC_LP__MUX2_0%A0
x_PM_SKY130_FD_SC_LP__MUX2_0%A_509_99# N_A_509_99#_M1007_d N_A_509_99#_M1000_d
+ N_A_509_99#_M1010_g N_A_509_99#_c_393_n N_A_509_99#_M1011_g
+ N_A_509_99#_c_401_n N_A_509_99#_c_394_n N_A_509_99#_c_395_n
+ N_A_509_99#_c_396_n N_A_509_99#_c_397_n N_A_509_99#_c_398_n
+ N_A_509_99#_c_404_n PM_SKY130_FD_SC_LP__MUX2_0%A_509_99#
x_PM_SKY130_FD_SC_LP__MUX2_0%X N_X_M1009_s N_X_M1001_s N_X_c_460_n X X X X X X X
+ N_X_c_455_n X PM_SKY130_FD_SC_LP__MUX2_0%X
x_PM_SKY130_FD_SC_LP__MUX2_0%VPWR N_VPWR_M1001_d N_VPWR_M1011_d N_VPWR_c_480_n
+ N_VPWR_c_481_n N_VPWR_c_482_n N_VPWR_c_483_n VPWR N_VPWR_c_484_n
+ N_VPWR_c_479_n N_VPWR_c_486_n PM_SKY130_FD_SC_LP__MUX2_0%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_0%VGND N_VGND_M1009_d N_VGND_M1010_d N_VGND_c_525_n
+ N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n
+ VGND N_VGND_c_531_n N_VGND_c_532_n PM_SKY130_FD_SC_LP__MUX2_0%VGND
cc_1 VNB N_A_89_200#_c_87_n 0.0216605f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1
cc_2 VNB N_A_89_200#_c_88_n 0.0231477f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.505
cc_3 VNB N_A_89_200#_c_89_n 0.0102727f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.67
cc_4 VNB N_A_89_200#_c_90_n 0.00475782f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_5 VNB N_A_89_200#_c_91_n 0.0164297f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_6 VNB N_A_89_200#_c_92_n 0.00801865f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=0.955
cc_7 VNB N_A_89_200#_c_93_n 0.00103295f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.955
cc_8 VNB N_A_89_200#_c_94_n 0.00863877f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.815
cc_9 VNB N_S_c_165_n 0.0164048f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.67
cc_10 VNB N_S_M1007_g 0.0471143f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.68
cc_11 VNB N_S_c_167_n 0.0181351f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_12 VNB N_S_c_168_n 0.0112697f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.955
cc_13 VNB S 0.00377321f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_14 VNB N_S_c_170_n 0.0274127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_283_n 0.0132602f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.775
cc_16 VNB N_A1_c_284_n 0.0448671f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1
cc_17 VNB N_A1_c_285_n 0.0171978f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.165
cc_18 VNB N_A1_c_286_n 0.00547443f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.625
cc_19 VNB N_A0_c_342_n 0.0366528f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.67
cc_20 VNB N_A0_M1003_g 0.028087f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1
cc_21 VNB A0 0.011473f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.04
cc_22 VNB N_A0_c_345_n 0.023624f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.625
cc_23 VNB N_A_509_99#_M1010_g 0.0190073f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.775
cc_24 VNB N_A_509_99#_c_393_n 0.0220041f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.68
cc_25 VNB N_A_509_99#_c_394_n 0.00723552f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_26 VNB N_A_509_99#_c_395_n 0.0385412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_509_99#_c_396_n 0.0152279f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=0.955
cc_28 VNB N_A_509_99#_c_397_n 0.00242643f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.985
cc_29 VNB N_A_509_99#_c_398_n 0.0167179f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.625
cc_30 VNB X 0.0483559f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.68
cc_31 VNB N_X_c_455_n 0.0140713f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.625
cc_32 VNB N_VPWR_c_479_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.9
cc_33 VNB N_VGND_c_525_n 0.0122996f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.775
cc_34 VNB N_VGND_c_526_n 0.0253736f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.68
cc_35 VNB N_VGND_c_527_n 0.0250726f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.505
cc_36 VNB N_VGND_c_528_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.67
cc_37 VNB N_VGND_c_529_n 0.0425027f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.165
cc_38 VNB N_VGND_c_530_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.165
cc_39 VNB N_VGND_c_531_n 0.0268053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_532_n 0.260934f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.835
cc_41 VPB N_A_89_200#_M1001_g 0.0612086f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.775
cc_42 VPB N_A_89_200#_c_89_n 0.00616441f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.67
cc_43 VPB N_A_89_200#_c_90_n 0.00748613f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.165
cc_44 VPB N_A_89_200#_c_98_n 0.0113763f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.625
cc_45 VPB N_A_89_200#_c_94_n 0.00362468f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.815
cc_46 VPB N_A_89_200#_c_100_n 0.0110183f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.9
cc_47 VPB N_S_M1002_g 0.0189977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_S_M1000_g 0.0362978f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.505
cc_49 VPB N_S_c_168_n 0.00625302f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.955
cc_50 VPB N_S_c_174_n 0.0176988f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.625
cc_51 VPB N_S_c_175_n 0.00690751f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.625
cc_52 VPB N_S_c_176_n 0.0331611f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.815
cc_53 VPB N_S_c_177_n 0.00340496f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.9
cc_54 VPB N_S_c_178_n 0.0129271f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_S_c_179_n 0.00235546f $X=-0.19 $Y=1.655 $X2=1.98 $Y2=0.835
cc_56 VPB N_S_c_180_n 9.84701e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_S_c_181_n 0.00728113f $X=-0.19 $Y=1.655 $X2=1.98 $Y2=0.955
cc_58 VPB N_S_c_182_n 4.25224e-19 $X=-0.19 $Y=1.655 $X2=1.98 $Y2=1.04
cc_59 VPB S 0.00623249f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.165
cc_60 VPB S 0.00449787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_S_c_185_n 0.0259076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_S_c_170_n 0.0178924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A1_M1006_g 0.023525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A1_c_288_n 0.0473217f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=0.955
cc_65 VPB N_A1_c_289_n 0.00303536f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.955
cc_66 VPB N_A1_c_286_n 0.00905331f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.625
cc_67 VPB N_A0_M1005_g 0.032838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A0_c_347_n 0.0121025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A0_c_348_n 0.0175152f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1
cc_70 VPB N_A0_c_345_n 0.00898924f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.625
cc_71 VPB N_A_509_99#_c_393_n 0.00107884f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.68
cc_72 VPB N_A_509_99#_M1011_g 0.0541578f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1
cc_73 VPB N_A_509_99#_c_401_n 0.0214872f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.67
cc_74 VPB N_A_509_99#_c_396_n 0.0466695f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=0.955
cc_75 VPB N_A_509_99#_c_397_n 7.11642e-19 $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.985
cc_76 VPB N_A_509_99#_c_404_n 0.0127871f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.9
cc_77 VPB X 0.0426083f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.68
cc_78 VPB X 0.0116396f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.505
cc_79 VPB X 0.018008f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.67
cc_80 VPB N_VPWR_c_480_n 0.0141908f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1
cc_81 VPB N_VPWR_c_481_n 0.00727313f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1
cc_82 VPB N_VPWR_c_482_n 0.047328f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=1.04
cc_83 VPB N_VPWR_c_483_n 0.00382106f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=1.165
cc_84 VPB N_VPWR_c_484_n 0.0204881f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.815
cc_85 VPB N_VPWR_c_479_n 0.0645684f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.9
cc_86 VPB N_VPWR_c_486_n 0.0258177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 N_A_89_200#_M1001_g N_S_M1002_g 0.0105481f $X=0.52 $Y=2.775 $X2=0 $Y2=0
cc_88 N_A_89_200#_c_87_n N_S_c_165_n 0.0156597f $X=0.61 $Y=1 $X2=0 $Y2=0
cc_89 N_A_89_200#_c_92_n N_S_c_165_n 0.011065f $X=1.845 $Y=0.955 $X2=0 $Y2=0
cc_90 N_A_89_200#_c_90_n N_S_c_167_n 0.00637714f $X=0.61 $Y=1.165 $X2=0 $Y2=0
cc_91 N_A_89_200#_c_91_n N_S_c_167_n 0.0201429f $X=0.61 $Y=1.165 $X2=0 $Y2=0
cc_92 N_A_89_200#_c_92_n N_S_c_167_n 0.00827684f $X=1.845 $Y=0.955 $X2=0 $Y2=0
cc_93 N_A_89_200#_M1001_g N_S_c_175_n 7.87709e-19 $X=0.52 $Y=2.775 $X2=0 $Y2=0
cc_94 N_A_89_200#_c_98_n N_S_c_175_n 0.0151111f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_95 N_A_89_200#_M1001_g N_S_c_176_n 0.0202971f $X=0.52 $Y=2.775 $X2=0 $Y2=0
cc_96 N_A_89_200#_c_98_n N_S_c_176_n 2.80815e-19 $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_97 N_A_89_200#_c_98_n N_S_c_177_n 0.0207794f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_98 N_A_89_200#_M1005_d N_S_c_178_n 0.00414818f $X=1.495 $Y=2.455 $X2=0 $Y2=0
cc_99 N_A_89_200#_c_98_n N_S_c_178_n 0.025017f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_100 N_A_89_200#_M1001_g N_S_c_170_n 0.00979707f $X=0.52 $Y=2.775 $X2=0 $Y2=0
cc_101 N_A_89_200#_c_88_n N_S_c_170_n 0.0201429f $X=0.61 $Y=1.505 $X2=0 $Y2=0
cc_102 N_A_89_200#_c_100_n N_S_c_170_n 7.56695e-19 $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_103 N_A_89_200#_c_92_n N_A1_c_283_n 0.00653538f $X=1.845 $Y=0.955 $X2=0 $Y2=0
cc_104 N_A_89_200#_c_118_p N_A1_c_283_n 0.0204956f $X=2.01 $Y=0.835 $X2=0 $Y2=0
cc_105 N_A_89_200#_c_118_p N_A1_c_284_n 0.00299988f $X=2.01 $Y=0.835 $X2=0 $Y2=0
cc_106 N_A_89_200#_c_92_n N_A1_c_285_n 0.0103983f $X=1.845 $Y=0.955 $X2=0 $Y2=0
cc_107 N_A_89_200#_c_94_n N_A1_c_285_n 0.00300054f $X=2.03 $Y=1.815 $X2=0 $Y2=0
cc_108 N_A_89_200#_c_98_n N_A1_c_288_n 0.00755841f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_109 N_A_89_200#_c_100_n N_A1_c_288_n 0.00340028f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_110 N_A_89_200#_c_98_n N_A1_c_289_n 0.0439033f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_111 N_A_89_200#_c_100_n N_A1_c_289_n 0.00381218f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_112 N_A_89_200#_c_98_n N_A1_c_286_n 0.00716858f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_113 N_A_89_200#_c_100_n N_A1_c_286_n 0.0133892f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_114 N_A_89_200#_c_118_p N_A1_c_286_n 0.0791877f $X=2.01 $Y=0.835 $X2=0 $Y2=0
cc_115 N_A_89_200#_c_98_n N_A0_M1005_g 0.00740321f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_116 N_A_89_200#_c_94_n N_A0_c_347_n 0.00278394f $X=2.03 $Y=1.815 $X2=0 $Y2=0
cc_117 N_A_89_200#_c_100_n N_A0_c_347_n 0.00419388f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_118 N_A_89_200#_c_94_n N_A0_c_342_n 0.0128999f $X=2.03 $Y=1.815 $X2=0 $Y2=0
cc_119 N_A_89_200#_c_100_n N_A0_c_342_n 0.00568724f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_120 N_A_89_200#_c_118_p N_A0_c_342_n 0.00290214f $X=2.01 $Y=0.835 $X2=0 $Y2=0
cc_121 N_A_89_200#_c_118_p N_A0_M1003_g 0.00713994f $X=2.01 $Y=0.835 $X2=0 $Y2=0
cc_122 N_A_89_200#_c_98_n N_A0_c_348_n 0.00334051f $X=1.73 $Y=2.625 $X2=0 $Y2=0
cc_123 N_A_89_200#_c_100_n N_A0_c_348_n 0.00321283f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_124 N_A_89_200#_c_88_n A0 5.24448e-19 $X=0.61 $Y=1.505 $X2=0 $Y2=0
cc_125 N_A_89_200#_c_90_n A0 0.0293385f $X=0.61 $Y=1.165 $X2=0 $Y2=0
cc_126 N_A_89_200#_c_92_n A0 0.0582733f $X=1.845 $Y=0.955 $X2=0 $Y2=0
cc_127 N_A_89_200#_c_94_n A0 0.0353265f $X=2.03 $Y=1.815 $X2=0 $Y2=0
cc_128 N_A_89_200#_c_100_n A0 0.0160897f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_129 N_A_89_200#_c_92_n N_A0_c_345_n 9.65602e-19 $X=1.845 $Y=0.955 $X2=0 $Y2=0
cc_130 N_A_89_200#_c_94_n N_A0_c_345_n 0.00328295f $X=2.03 $Y=1.815 $X2=0 $Y2=0
cc_131 N_A_89_200#_c_100_n N_A0_c_345_n 0.00438376f $X=2.03 $Y=1.9 $X2=0 $Y2=0
cc_132 N_A_89_200#_c_93_n N_X_M1009_s 6.98889e-19 $X=0.78 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_89_200#_c_87_n N_X_c_460_n 0.00304732f $X=0.61 $Y=1 $X2=0 $Y2=0
cc_134 N_A_89_200#_c_91_n N_X_c_460_n 0.00338816f $X=0.61 $Y=1.165 $X2=0 $Y2=0
cc_135 N_A_89_200#_c_93_n N_X_c_460_n 0.00548028f $X=0.78 $Y=0.955 $X2=0 $Y2=0
cc_136 N_A_89_200#_c_87_n X 0.00488269f $X=0.61 $Y=1 $X2=0 $Y2=0
cc_137 N_A_89_200#_c_90_n X 0.0480443f $X=0.61 $Y=1.165 $X2=0 $Y2=0
cc_138 N_A_89_200#_c_91_n X 0.0437006f $X=0.61 $Y=1.165 $X2=0 $Y2=0
cc_139 N_A_89_200#_c_93_n X 0.014578f $X=0.78 $Y=0.955 $X2=0 $Y2=0
cc_140 N_A_89_200#_M1001_g X 0.00360377f $X=0.52 $Y=2.775 $X2=0 $Y2=0
cc_141 N_A_89_200#_M1001_g X 0.0045279f $X=0.52 $Y=2.775 $X2=0 $Y2=0
cc_142 N_A_89_200#_M1001_g N_VPWR_c_480_n 0.00657308f $X=0.52 $Y=2.775 $X2=0
+ $Y2=0
cc_143 N_A_89_200#_M1001_g N_VPWR_c_479_n 0.0120391f $X=0.52 $Y=2.775 $X2=0
+ $Y2=0
cc_144 N_A_89_200#_M1001_g N_VPWR_c_486_n 0.00549943f $X=0.52 $Y=2.775 $X2=0
+ $Y2=0
cc_145 N_A_89_200#_c_92_n N_VGND_M1009_d 0.00261503f $X=1.845 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_89_200#_c_87_n N_VGND_c_525_n 0.00483713f $X=0.61 $Y=1 $X2=0 $Y2=0
cc_147 N_A_89_200#_c_92_n N_VGND_c_525_n 0.0218002f $X=1.845 $Y=0.955 $X2=0
+ $Y2=0
cc_148 N_A_89_200#_c_87_n N_VGND_c_527_n 0.00484939f $X=0.61 $Y=1 $X2=0 $Y2=0
cc_149 N_A_89_200#_c_87_n N_VGND_c_532_n 0.00514438f $X=0.61 $Y=1 $X2=0 $Y2=0
cc_150 N_A_89_200#_c_92_n A_257_94# 0.0111828f $X=1.845 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_151 N_S_c_178_n N_A1_M1006_g 0.0147663f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_152 N_S_c_180_n N_A1_M1006_g 0.00120917f $X=2.72 $Y=2.905 $X2=0 $Y2=0
cc_153 N_S_c_165_n N_A1_c_283_n 5.9531e-19 $X=1.21 $Y=1 $X2=0 $Y2=0
cc_154 N_S_c_165_n N_A1_c_284_n 0.0137853f $X=1.21 $Y=1 $X2=0 $Y2=0
cc_155 N_S_c_167_n N_A1_c_285_n 0.0137853f $X=1.21 $Y=1.075 $X2=0 $Y2=0
cc_156 N_S_c_170_n N_A1_c_285_n 7.20368e-19 $X=0.97 $Y=1.965 $X2=0 $Y2=0
cc_157 N_S_c_178_n N_A1_c_288_n 0.00100021f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_158 N_S_c_178_n N_A1_c_289_n 0.0221527f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_159 N_S_c_180_n N_A1_c_289_n 0.0162593f $X=2.72 $Y=2.905 $X2=0 $Y2=0
cc_160 N_S_c_182_n N_A1_c_289_n 0.0144749f $X=2.805 $Y=2.405 $X2=0 $Y2=0
cc_161 S N_A1_c_286_n 0.0178523f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_162 N_S_c_176_n N_A0_M1005_g 0.0304505f $X=0.97 $Y=2.13 $X2=0 $Y2=0
cc_163 N_S_c_177_n N_A0_M1005_g 0.00360313f $X=1.245 $Y=2.905 $X2=0 $Y2=0
cc_164 N_S_c_178_n N_A0_M1005_g 0.0126759f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_165 N_S_c_175_n N_A0_c_348_n 0.00193798f $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_166 N_S_c_170_n N_A0_c_348_n 0.0304505f $X=0.97 $Y=1.965 $X2=0 $Y2=0
cc_167 N_S_c_167_n A0 0.00459868f $X=1.21 $Y=1.075 $X2=0 $Y2=0
cc_168 N_S_c_175_n A0 0.0146366f $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_169 N_S_c_170_n A0 0.020301f $X=0.97 $Y=1.965 $X2=0 $Y2=0
cc_170 N_S_c_170_n N_A0_c_345_n 0.0230207f $X=0.97 $Y=1.965 $X2=0 $Y2=0
cc_171 N_S_M1007_g N_A_509_99#_M1010_g 0.0146706f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_172 N_S_c_168_n N_A_509_99#_c_393_n 0.0174953f $X=3.285 $Y=1.73 $X2=0 $Y2=0
cc_173 S N_A_509_99#_c_393_n 0.00229847f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_174 N_S_M1000_g N_A_509_99#_M1011_g 0.0152776f $X=3.295 $Y=2.785 $X2=0 $Y2=0
cc_175 N_S_c_178_n N_A_509_99#_M1011_g 0.00836889f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_176 N_S_c_180_n N_A_509_99#_M1011_g 0.0124466f $X=2.72 $Y=2.905 $X2=0 $Y2=0
cc_177 N_S_c_182_n N_A_509_99#_M1011_g 0.0090514f $X=2.805 $Y=2.405 $X2=0 $Y2=0
cc_178 S N_A_509_99#_M1011_g 0.00496252f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_179 N_S_c_185_n N_A_509_99#_M1011_g 0.0113058f $X=3.3 $Y=1.745 $X2=0 $Y2=0
cc_180 N_S_c_181_n N_A_509_99#_c_401_n 0.00246303f $X=2.985 $Y=2.405 $X2=0 $Y2=0
cc_181 N_S_c_182_n N_A_509_99#_c_401_n 2.69515e-19 $X=2.805 $Y=2.405 $X2=0 $Y2=0
cc_182 N_S_c_185_n N_A_509_99#_c_401_n 0.00598993f $X=3.3 $Y=1.745 $X2=0 $Y2=0
cc_183 N_S_M1007_g N_A_509_99#_c_394_n 0.0110116f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_184 S N_A_509_99#_c_394_n 0.0199195f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_185 N_S_M1007_g N_A_509_99#_c_395_n 0.0135657f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_186 N_S_c_168_n N_A_509_99#_c_395_n 0.00434654f $X=3.285 $Y=1.73 $X2=0 $Y2=0
cc_187 S N_A_509_99#_c_395_n 0.0135618f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_188 N_S_M1007_g N_A_509_99#_c_396_n 0.00532863f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_189 N_S_M1000_g N_A_509_99#_c_396_n 0.0059815f $X=3.295 $Y=2.785 $X2=0 $Y2=0
cc_190 N_S_c_168_n N_A_509_99#_c_396_n 0.0164304f $X=3.285 $Y=1.73 $X2=0 $Y2=0
cc_191 S N_A_509_99#_c_396_n 0.0592678f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_192 S N_A_509_99#_c_396_n 0.0137853f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_193 N_S_M1007_g N_A_509_99#_c_397_n 0.00112856f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_194 N_S_c_181_n N_A_509_99#_c_397_n 3.11741e-19 $X=2.985 $Y=2.405 $X2=0 $Y2=0
cc_195 N_S_c_182_n N_A_509_99#_c_397_n 0.00634827f $X=2.805 $Y=2.405 $X2=0 $Y2=0
cc_196 S N_A_509_99#_c_397_n 0.0253844f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_197 N_S_M1007_g N_A_509_99#_c_398_n 0.0174953f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_198 N_S_M1000_g N_A_509_99#_c_404_n 0.00352694f $X=3.295 $Y=2.785 $X2=0 $Y2=0
cc_199 N_S_c_174_n N_A_509_99#_c_404_n 0.00206735f $X=3.3 $Y=2.25 $X2=0 $Y2=0
cc_200 S N_A_509_99#_c_404_n 0.00254923f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_201 N_S_c_175_n X 0.00846523f $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_202 N_S_M1002_g X 2.23226e-19 $X=1.06 $Y=2.665 $X2=0 $Y2=0
cc_203 N_S_M1002_g N_VPWR_c_480_n 0.00783768f $X=1.06 $Y=2.665 $X2=0 $Y2=0
cc_204 N_S_c_175_n N_VPWR_c_480_n 0.0150805f $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_205 N_S_c_176_n N_VPWR_c_480_n 0.00434771f $X=0.97 $Y=2.13 $X2=0 $Y2=0
cc_206 N_S_c_177_n N_VPWR_c_480_n 0.0195633f $X=1.245 $Y=2.905 $X2=0 $Y2=0
cc_207 N_S_c_179_n N_VPWR_c_480_n 0.0146845f $X=1.33 $Y=2.99 $X2=0 $Y2=0
cc_208 N_S_M1000_g N_VPWR_c_481_n 0.00333864f $X=3.295 $Y=2.785 $X2=0 $Y2=0
cc_209 N_S_c_178_n N_VPWR_c_481_n 0.0101484f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_210 N_S_c_181_n N_VPWR_c_481_n 6.91618e-19 $X=2.985 $Y=2.405 $X2=0 $Y2=0
cc_211 S N_VPWR_c_481_n 0.0164075f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_212 N_S_M1002_g N_VPWR_c_482_n 0.0049872f $X=1.06 $Y=2.665 $X2=0 $Y2=0
cc_213 N_S_c_178_n N_VPWR_c_482_n 0.0952128f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_214 N_S_c_179_n N_VPWR_c_482_n 0.0121867f $X=1.33 $Y=2.99 $X2=0 $Y2=0
cc_215 N_S_M1000_g N_VPWR_c_484_n 0.00461917f $X=3.295 $Y=2.785 $X2=0 $Y2=0
cc_216 N_S_M1002_g N_VPWR_c_479_n 0.00505191f $X=1.06 $Y=2.665 $X2=0 $Y2=0
cc_217 N_S_M1000_g N_VPWR_c_479_n 0.00543698f $X=3.295 $Y=2.785 $X2=0 $Y2=0
cc_218 N_S_c_178_n N_VPWR_c_479_n 0.0542938f $X=2.635 $Y=2.99 $X2=0 $Y2=0
cc_219 N_S_c_179_n N_VPWR_c_479_n 0.00660921f $X=1.33 $Y=2.99 $X2=0 $Y2=0
cc_220 N_S_c_181_n N_VPWR_c_479_n 0.0059211f $X=2.985 $Y=2.405 $X2=0 $Y2=0
cc_221 S N_VPWR_c_479_n 0.00653049f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_222 N_S_c_177_n A_227_491# 0.00143999f $X=1.245 $Y=2.905 $X2=-0.19 $Y2=-0.245
cc_223 N_S_c_178_n A_423_515# 0.00729077f $X=2.635 $Y=2.99 $X2=-0.19 $Y2=-0.245
cc_224 N_S_c_165_n N_VGND_c_525_n 0.00905729f $X=1.21 $Y=1 $X2=0 $Y2=0
cc_225 N_S_c_167_n N_VGND_c_525_n 7.20696e-19 $X=1.21 $Y=1.075 $X2=0 $Y2=0
cc_226 N_S_M1007_g N_VGND_c_526_n 0.0059501f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_227 N_S_c_165_n N_VGND_c_529_n 0.00421418f $X=1.21 $Y=1 $X2=0 $Y2=0
cc_228 N_S_M1007_g N_VGND_c_531_n 0.00415323f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_229 N_S_c_165_n N_VGND_c_532_n 0.00432128f $X=1.21 $Y=1 $X2=0 $Y2=0
cc_230 N_S_M1007_g N_VGND_c_532_n 0.00469432f $X=3.18 $Y=0.835 $X2=0 $Y2=0
cc_231 N_A1_c_288_n N_A0_M1005_g 0.0175628f $X=2.24 $Y=2.25 $X2=0 $Y2=0
cc_232 N_A1_c_285_n N_A0_c_342_n 0.00168115f $X=1.81 $Y=0.515 $X2=0 $Y2=0
cc_233 N_A1_c_288_n N_A0_c_342_n 0.00827104f $X=2.24 $Y=2.25 $X2=0 $Y2=0
cc_234 N_A1_c_289_n N_A0_c_342_n 9.74816e-19 $X=2.24 $Y=2.25 $X2=0 $Y2=0
cc_235 N_A1_c_286_n N_A0_c_342_n 0.00415331f $X=2.265 $Y=2.155 $X2=0 $Y2=0
cc_236 N_A1_c_283_n N_A0_M1003_g 0.00789319f $X=2.295 $Y=0.382 $X2=0 $Y2=0
cc_237 N_A1_c_284_n N_A0_M1003_g 0.00129904f $X=1.81 $Y=0.35 $X2=0 $Y2=0
cc_238 N_A1_c_285_n N_A0_M1003_g 0.0120442f $X=1.81 $Y=0.515 $X2=0 $Y2=0
cc_239 N_A1_c_286_n N_A0_M1003_g 0.0167311f $X=2.265 $Y=2.155 $X2=0 $Y2=0
cc_240 N_A1_c_285_n A0 0.00110484f $X=1.81 $Y=0.515 $X2=0 $Y2=0
cc_241 N_A1_c_285_n N_A0_c_345_n 0.00784012f $X=1.81 $Y=0.515 $X2=0 $Y2=0
cc_242 N_A1_c_286_n N_A_509_99#_M1010_g 0.0171782f $X=2.265 $Y=2.155 $X2=0 $Y2=0
cc_243 N_A1_M1006_g N_A_509_99#_M1011_g 0.0144312f $X=2.04 $Y=2.785 $X2=0 $Y2=0
cc_244 N_A1_c_288_n N_A_509_99#_M1011_g 0.0194965f $X=2.24 $Y=2.25 $X2=0 $Y2=0
cc_245 N_A1_c_286_n N_A_509_99#_M1011_g 0.0108232f $X=2.265 $Y=2.155 $X2=0 $Y2=0
cc_246 N_A1_c_286_n N_A_509_99#_c_397_n 0.0493894f $X=2.265 $Y=2.155 $X2=0 $Y2=0
cc_247 N_A1_M1006_g N_VPWR_c_482_n 0.00296932f $X=2.04 $Y=2.785 $X2=0 $Y2=0
cc_248 N_A1_M1006_g N_VPWR_c_479_n 0.00470987f $X=2.04 $Y=2.785 $X2=0 $Y2=0
cc_249 N_A1_c_289_n A_423_515# 0.00539805f $X=2.24 $Y=2.25 $X2=-0.19 $Y2=-0.245
cc_250 N_A1_c_283_n N_VGND_c_525_n 0.00820812f $X=2.295 $Y=0.382 $X2=0 $Y2=0
cc_251 N_A1_c_284_n N_VGND_c_525_n 0.00319315f $X=1.81 $Y=0.35 $X2=0 $Y2=0
cc_252 N_A1_c_283_n N_VGND_c_526_n 0.0150468f $X=2.295 $Y=0.382 $X2=0 $Y2=0
cc_253 N_A1_c_286_n N_VGND_c_526_n 0.0164098f $X=2.265 $Y=2.155 $X2=0 $Y2=0
cc_254 N_A1_c_283_n N_VGND_c_529_n 0.0507531f $X=2.295 $Y=0.382 $X2=0 $Y2=0
cc_255 N_A1_c_284_n N_VGND_c_529_n 0.00651318f $X=1.81 $Y=0.35 $X2=0 $Y2=0
cc_256 N_A1_c_283_n N_VGND_c_532_n 0.0295296f $X=2.295 $Y=0.382 $X2=0 $Y2=0
cc_257 N_A1_c_284_n N_VGND_c_532_n 0.0101042f $X=1.81 $Y=0.35 $X2=0 $Y2=0
cc_258 N_A1_c_286_n A_467_125# 0.00420101f $X=2.265 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_259 N_A0_M1003_g N_A_509_99#_M1010_g 0.031868f $X=2.26 $Y=0.835 $X2=0 $Y2=0
cc_260 N_A0_c_342_n N_A_509_99#_c_398_n 0.031868f $X=2.185 $Y=1.49 $X2=0 $Y2=0
cc_261 N_A0_M1005_g N_VPWR_c_480_n 2.26373e-19 $X=1.42 $Y=2.665 $X2=0 $Y2=0
cc_262 N_A0_M1005_g N_VPWR_c_482_n 7.94855e-19 $X=1.42 $Y=2.665 $X2=0 $Y2=0
cc_263 N_A0_M1003_g N_VGND_c_529_n 5.58252e-19 $X=2.26 $Y=0.835 $X2=0 $Y2=0
cc_264 N_A_509_99#_M1011_g N_VPWR_c_481_n 0.00228847f $X=2.69 $Y=2.785 $X2=0
+ $Y2=0
cc_265 N_A_509_99#_M1011_g N_VPWR_c_482_n 0.00296793f $X=2.69 $Y=2.785 $X2=0
+ $Y2=0
cc_266 N_A_509_99#_c_404_n N_VPWR_c_484_n 0.0128164f $X=3.65 $Y=2.8 $X2=0 $Y2=0
cc_267 N_A_509_99#_M1011_g N_VPWR_c_479_n 0.00442969f $X=2.69 $Y=2.785 $X2=0
+ $Y2=0
cc_268 N_A_509_99#_c_404_n N_VPWR_c_479_n 0.0134797f $X=3.65 $Y=2.8 $X2=0 $Y2=0
cc_269 N_A_509_99#_M1010_g N_VGND_c_526_n 0.00359965f $X=2.62 $Y=0.835 $X2=0
+ $Y2=0
cc_270 N_A_509_99#_c_394_n N_VGND_c_526_n 0.0179894f $X=3.235 $Y=1.26 $X2=0
+ $Y2=0
cc_271 N_A_509_99#_c_397_n N_VGND_c_526_n 0.00566103f $X=2.73 $Y=1.34 $X2=0
+ $Y2=0
cc_272 N_A_509_99#_c_398_n N_VGND_c_526_n 0.00268111f $X=2.73 $Y=1.34 $X2=0
+ $Y2=0
cc_273 N_A_509_99#_M1010_g N_VGND_c_529_n 0.00415323f $X=2.62 $Y=0.835 $X2=0
+ $Y2=0
cc_274 N_A_509_99#_M1010_g N_VGND_c_532_n 0.00469432f $X=2.62 $Y=0.835 $X2=0
+ $Y2=0
cc_275 N_A_509_99#_c_395_n N_VGND_c_532_n 0.0131423f $X=3.65 $Y=1.345 $X2=0
+ $Y2=0
cc_276 X N_VPWR_c_480_n 0.0241942f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_277 N_X_M1001_s N_VPWR_c_479_n 0.00216391f $X=0.18 $Y=2.455 $X2=0 $Y2=0
cc_278 X N_VPWR_c_479_n 0.0144743f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_279 X N_VPWR_c_486_n 0.0209488f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_280 N_X_c_460_n N_VGND_c_527_n 0.00721265f $X=0.485 $Y=0.595 $X2=0 $Y2=0
cc_281 N_X_c_455_n N_VGND_c_527_n 0.00807944f $X=0.22 $Y=0.7 $X2=0 $Y2=0
cc_282 N_X_c_460_n N_VGND_c_532_n 0.00962361f $X=0.485 $Y=0.595 $X2=0 $Y2=0
cc_283 N_X_c_455_n N_VGND_c_532_n 0.0092236f $X=0.22 $Y=0.7 $X2=0 $Y2=0
