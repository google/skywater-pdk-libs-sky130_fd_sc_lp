* File: sky130_fd_sc_lp__a22o_0.pxi.spice
* Created: Wed Sep  2 09:22:21 2020
* 
x_PM_SKY130_FD_SC_LP__A22O_0%A_85_155# N_A_85_155#_M1009_d N_A_85_155#_M1000_d
+ N_A_85_155#_M1008_g N_A_85_155#_M1005_g N_A_85_155#_c_67_n N_A_85_155#_c_68_n
+ N_A_85_155#_c_69_n N_A_85_155#_c_70_n N_A_85_155#_c_71_n N_A_85_155#_c_72_n
+ N_A_85_155#_c_77_n N_A_85_155#_c_78_n N_A_85_155#_c_73_n N_A_85_155#_c_84_p
+ N_A_85_155#_c_95_p N_A_85_155#_c_79_n N_A_85_155#_c_74_n
+ PM_SKY130_FD_SC_LP__A22O_0%A_85_155#
x_PM_SKY130_FD_SC_LP__A22O_0%A2 N_A2_M1003_g N_A2_M1007_g N_A2_c_154_n
+ N_A2_c_159_n A2 A2 N_A2_c_156_n PM_SKY130_FD_SC_LP__A22O_0%A2
x_PM_SKY130_FD_SC_LP__A22O_0%A1 N_A1_M1009_g N_A1_M1002_g N_A1_c_199_n
+ N_A1_c_200_n A1 A1 A1 A1 N_A1_c_202_n N_A1_c_203_n N_A1_c_204_n
+ PM_SKY130_FD_SC_LP__A22O_0%A1
x_PM_SKY130_FD_SC_LP__A22O_0%B1 N_B1_M1000_g N_B1_M1001_g N_B1_c_246_n
+ N_B1_c_250_n B1 B1 N_B1_c_248_n PM_SKY130_FD_SC_LP__A22O_0%B1
x_PM_SKY130_FD_SC_LP__A22O_0%B2 N_B2_M1006_g N_B2_M1004_g B2 B2 N_B2_c_297_n
+ PM_SKY130_FD_SC_LP__A22O_0%B2
x_PM_SKY130_FD_SC_LP__A22O_0%X N_X_M1008_s N_X_M1005_s X X X X X X X N_X_c_333_n
+ N_X_c_335_n PM_SKY130_FD_SC_LP__A22O_0%X
x_PM_SKY130_FD_SC_LP__A22O_0%VPWR N_VPWR_M1005_d N_VPWR_M1002_d N_VPWR_c_352_n
+ N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n VPWR
+ N_VPWR_c_357_n N_VPWR_c_351_n PM_SKY130_FD_SC_LP__A22O_0%VPWR
x_PM_SKY130_FD_SC_LP__A22O_0%A_257_491# N_A_257_491#_M1007_d
+ N_A_257_491#_M1006_d N_A_257_491#_c_388_n N_A_257_491#_c_389_n
+ N_A_257_491#_c_394_n N_A_257_491#_c_387_n
+ PM_SKY130_FD_SC_LP__A22O_0%A_257_491#
x_PM_SKY130_FD_SC_LP__A22O_0%VGND N_VGND_M1008_d N_VGND_M1004_d N_VGND_c_411_n
+ N_VGND_c_412_n VGND N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n N_VGND_c_417_n PM_SKY130_FD_SC_LP__A22O_0%VGND
cc_1 VNB N_A_85_155#_M1005_g 0.0119285f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_2 VNB N_A_85_155#_c_67_n 0.0207705f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.775
cc_3 VNB N_A_85_155#_c_68_n 0.0240092f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.28
cc_4 VNB N_A_85_155#_c_69_n 0.0188793f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.445
cc_5 VNB N_A_85_155#_c_70_n 0.00107176f $X=-0.19 $Y=-0.245 $X2=0.632 $Y2=0.945
cc_6 VNB N_A_85_155#_c_71_n 0.00777416f $X=-0.19 $Y=-0.245 $X2=0.632 $Y2=2.155
cc_7 VNB N_A_85_155#_c_72_n 0.0132042f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.86
cc_8 VNB N_A_85_155#_c_73_n 0.00113254f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=0.775
cc_9 VNB N_A_85_155#_c_74_n 0.0169831f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.94
cc_10 VNB N_A2_M1003_g 0.0467913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_154_n 0.0100491f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_12 VNB A2 0.00719531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_156_n 0.0157889f $X=-0.19 $Y=-0.245 $X2=0.632 $Y2=0.945
cc_14 VNB N_A1_c_199_n 0.0261857f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.445
cc_15 VNB N_A1_c_200_n 0.0352859f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_16 VNB A1 0.033848f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.94
cc_17 VNB N_A1_c_202_n 0.0169118f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=2.24
cc_18 VNB N_A1_c_203_n 0.0325193f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=0.775
cc_19 VNB N_A1_c_204_n 0.0230201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_M1001_g 0.0443562f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.775
cc_21 VNB N_B1_c_246_n 0.0253773f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_22 VNB B1 0.00664377f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.28
cc_23 VNB N_B1_c_248_n 0.0117822f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.86
cc_24 VNB N_B2_M1004_g 0.0681697f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.775
cc_25 VNB B2 0.00808945f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.445
cc_26 VNB X 0.0540222f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.775
cc_27 VNB N_X_c_333_n 0.0149364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_351_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_411_n 0.00235386f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_30 VNB N_VGND_c_412_n 0.017485f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.775
cc_31 VNB N_VGND_c_413_n 0.0411613f $X=-0.19 $Y=-0.245 $X2=0.632 $Y2=2.155
cc_32 VNB N_VGND_c_414_n 0.0218729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_415_n 0.194928f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.325
cc_34 VNB N_VGND_c_416_n 0.0213286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_417_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.94
cc_36 VPB N_A_85_155#_M1005_g 0.061901f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_37 VPB N_A_85_155#_c_71_n 0.00890571f $X=-0.19 $Y=1.655 $X2=0.632 $Y2=2.155
cc_38 VPB N_A_85_155#_c_77_n 0.0309472f $X=-0.19 $Y=1.655 $X2=1.76 $Y2=2.24
cc_39 VPB N_A_85_155#_c_78_n 0.00331422f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.24
cc_40 VPB N_A_85_155#_c_79_n 0.0034039f $X=-0.19 $Y=1.655 $X2=1.925 $Y2=2.63
cc_41 VPB N_A2_M1007_g 0.0355542f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.775
cc_42 VPB N_A2_c_154_n 0.0120067f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_43 VPB N_A2_c_159_n 0.0155414f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_44 VPB A2 0.00236188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A1_M1002_g 0.0406944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB A1 0.0300959f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.94
cc_47 VPB N_A1_c_203_n 0.0524658f $X=-0.19 $Y=1.655 $X2=1.13 $Y2=0.775
cc_48 VPB N_B1_M1000_g 0.0353421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B1_c_250_n 0.0151826f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.775
cc_50 VPB B1 0.00236188f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.28
cc_51 VPB N_B1_c_248_n 0.0120848f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.86
cc_52 VPB N_B2_M1006_g 0.0368564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B2_M1004_g 0.00309336f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.775
cc_54 VPB B2 0.00339432f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.445
cc_55 VPB N_B2_c_297_n 0.0358568f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.94
cc_56 VPB X 0.0434765f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.775
cc_57 VPB N_X_c_335_n 0.0289193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_352_n 0.0055232f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.445
cc_59 VPB N_VPWR_c_353_n 0.0143797f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_60 VPB N_VPWR_c_354_n 0.0298975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_355_n 0.0214649f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.28
cc_62 VPB N_VPWR_c_356_n 0.00631455f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.445
cc_63 VPB N_VPWR_c_357_n 0.0405583f $X=-0.19 $Y=1.655 $X2=1.13 $Y2=0.61
cc_64 VPB N_VPWR_c_351_n 0.0509055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_257_491#_c_387_n 0.00877716f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.775
cc_66 N_A_85_155#_c_67_n N_A2_M1003_g 0.0142574f $X=0.59 $Y=0.775 $X2=0 $Y2=0
cc_67 N_A_85_155#_c_71_n N_A2_M1003_g 0.00451465f $X=0.632 $Y=2.155 $X2=0 $Y2=0
cc_68 N_A_85_155#_c_72_n N_A2_M1003_g 0.00769501f $X=1.045 $Y=0.86 $X2=0 $Y2=0
cc_69 N_A_85_155#_c_73_n N_A2_M1003_g 0.00470013f $X=1.13 $Y=0.775 $X2=0 $Y2=0
cc_70 N_A_85_155#_c_84_p N_A2_M1003_g 0.0104888f $X=1.215 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_85_155#_c_74_n N_A2_M1003_g 0.025535f $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_72 N_A_85_155#_M1005_g N_A2_M1007_g 0.0246702f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_73 N_A_85_155#_c_71_n N_A2_M1007_g 0.00274897f $X=0.632 $Y=2.155 $X2=0 $Y2=0
cc_74 N_A_85_155#_c_77_n N_A2_M1007_g 0.0148608f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_75 N_A_85_155#_c_77_n N_A2_c_159_n 0.00484128f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_76 N_A_85_155#_M1005_g A2 6.68332e-19 $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_77 N_A_85_155#_c_68_n A2 5.66277e-19 $X=0.59 $Y=1.28 $X2=0 $Y2=0
cc_78 N_A_85_155#_c_71_n A2 0.049656f $X=0.632 $Y=2.155 $X2=0 $Y2=0
cc_79 N_A_85_155#_c_72_n A2 0.0143027f $X=1.045 $Y=0.86 $X2=0 $Y2=0
cc_80 N_A_85_155#_c_77_n A2 0.0286025f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_81 N_A_85_155#_c_95_p A2 0.00442876f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_85_155#_M1005_g N_A2_c_156_n 0.0267527f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_83 N_A_85_155#_c_69_n N_A2_c_156_n 0.00586648f $X=0.59 $Y=1.445 $X2=0 $Y2=0
cc_84 N_A_85_155#_c_71_n N_A2_c_156_n 0.00438859f $X=0.632 $Y=2.155 $X2=0 $Y2=0
cc_85 N_A_85_155#_c_72_n N_A2_c_156_n 3.55524e-19 $X=1.045 $Y=0.86 $X2=0 $Y2=0
cc_86 N_A_85_155#_c_71_n N_A1_c_199_n 0.00207015f $X=0.632 $Y=2.155 $X2=0 $Y2=0
cc_87 N_A_85_155#_c_72_n N_A1_c_199_n 0.0146713f $X=1.045 $Y=0.86 $X2=0 $Y2=0
cc_88 N_A_85_155#_c_95_p N_A1_c_199_n 0.0265634f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_85_155#_c_72_n N_A1_c_200_n 7.80677e-19 $X=1.045 $Y=0.86 $X2=0 $Y2=0
cc_90 N_A_85_155#_c_95_p N_A1_c_200_n 0.00402428f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_85_155#_c_73_n N_A1_c_202_n 0.00247302f $X=1.13 $Y=0.775 $X2=0 $Y2=0
cc_92 N_A_85_155#_c_95_p N_A1_c_202_n 0.0110483f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_85_155#_c_77_n N_B1_M1000_g 0.0123873f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_94 N_A_85_155#_c_79_n N_B1_M1000_g 0.005305f $X=1.925 $Y=2.63 $X2=0 $Y2=0
cc_95 N_A_85_155#_c_95_p N_B1_M1001_g 0.00479244f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_85_155#_c_77_n N_B1_c_246_n 0.00471862f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_97 N_A_85_155#_c_77_n N_B1_c_250_n 0.00490231f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_98 N_A_85_155#_c_77_n B1 0.0296555f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_99 N_A_85_155#_c_77_n N_B2_M1006_g 0.00590752f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_100 N_A_85_155#_c_79_n N_B2_M1006_g 0.00367741f $X=1.925 $Y=2.63 $X2=0 $Y2=0
cc_101 N_A_85_155#_c_77_n B2 0.00222328f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_102 N_A_85_155#_M1005_g X 0.01021f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_103 N_A_85_155#_c_67_n X 0.00596091f $X=0.59 $Y=0.775 $X2=0 $Y2=0
cc_104 N_A_85_155#_c_70_n X 0.0139766f $X=0.632 $Y=0.945 $X2=0 $Y2=0
cc_105 N_A_85_155#_c_71_n X 0.0946364f $X=0.632 $Y=2.155 $X2=0 $Y2=0
cc_106 N_A_85_155#_c_78_n X 0.0147443f $X=0.76 $Y=2.24 $X2=0 $Y2=0
cc_107 N_A_85_155#_c_74_n X 0.0166276f $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_108 N_A_85_155#_c_74_n N_X_c_333_n 0.00153556f $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_109 N_A_85_155#_M1005_g N_X_c_335_n 0.00516732f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_110 N_A_85_155#_c_78_n N_X_c_335_n 0.00500698f $X=0.76 $Y=2.24 $X2=0 $Y2=0
cc_111 N_A_85_155#_M1005_g N_VPWR_c_352_n 0.00326553f $X=0.66 $Y=2.775 $X2=0
+ $Y2=0
cc_112 N_A_85_155#_c_77_n N_VPWR_c_352_n 0.0252372f $X=1.76 $Y=2.24 $X2=0 $Y2=0
cc_113 N_A_85_155#_M1005_g N_VPWR_c_355_n 0.00579312f $X=0.66 $Y=2.775 $X2=0
+ $Y2=0
cc_114 N_A_85_155#_M1000_d N_VPWR_c_351_n 0.0031466f $X=1.715 $Y=2.455 $X2=0
+ $Y2=0
cc_115 N_A_85_155#_M1005_g N_VPWR_c_351_n 0.011779f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_116 N_A_85_155#_c_77_n N_A_257_491#_c_388_n 0.020482f $X=1.76 $Y=2.24 $X2=0
+ $Y2=0
cc_117 N_A_85_155#_M1000_d N_A_257_491#_c_389_n 0.00580468f $X=1.715 $Y=2.455
+ $X2=0 $Y2=0
cc_118 N_A_85_155#_c_77_n N_A_257_491#_c_389_n 0.00377396f $X=1.76 $Y=2.24 $X2=0
+ $Y2=0
cc_119 N_A_85_155#_c_79_n N_A_257_491#_c_389_n 0.0207521f $X=1.925 $Y=2.63 $X2=0
+ $Y2=0
cc_120 N_A_85_155#_c_79_n N_A_257_491#_c_387_n 6.24934e-19 $X=1.925 $Y=2.63
+ $X2=0 $Y2=0
cc_121 N_A_85_155#_c_67_n N_VGND_c_411_n 0.00764514f $X=0.59 $Y=0.775 $X2=0
+ $Y2=0
cc_122 N_A_85_155#_c_70_n N_VGND_c_411_n 0.00530185f $X=0.632 $Y=0.945 $X2=0
+ $Y2=0
cc_123 N_A_85_155#_c_72_n N_VGND_c_411_n 0.00705394f $X=1.045 $Y=0.86 $X2=0
+ $Y2=0
cc_124 N_A_85_155#_c_84_p N_VGND_c_411_n 0.0212766f $X=1.215 $Y=0.445 $X2=0
+ $Y2=0
cc_125 N_A_85_155#_c_74_n N_VGND_c_411_n 5.84318e-19 $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_126 N_A_85_155#_c_95_p N_VGND_c_412_n 0.00959326f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_127 N_A_85_155#_c_84_p N_VGND_c_413_n 0.00883178f $X=1.215 $Y=0.445 $X2=0
+ $Y2=0
cc_128 N_A_85_155#_c_95_p N_VGND_c_413_n 0.0285494f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_129 N_A_85_155#_M1009_d N_VGND_c_415_n 0.00398687f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_130 N_A_85_155#_c_67_n N_VGND_c_415_n 0.0059772f $X=0.59 $Y=0.775 $X2=0 $Y2=0
cc_131 N_A_85_155#_c_70_n N_VGND_c_415_n 0.00526932f $X=0.632 $Y=0.945 $X2=0
+ $Y2=0
cc_132 N_A_85_155#_c_72_n N_VGND_c_415_n 0.00655975f $X=1.045 $Y=0.86 $X2=0
+ $Y2=0
cc_133 N_A_85_155#_c_84_p N_VGND_c_415_n 0.00592031f $X=1.215 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_A_85_155#_c_95_p N_VGND_c_415_n 0.0205527f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_135 N_A_85_155#_c_74_n N_VGND_c_415_n 6.43983e-19 $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_136 N_A_85_155#_c_67_n N_VGND_c_416_n 0.00564095f $X=0.59 $Y=0.775 $X2=0
+ $Y2=0
cc_137 N_A_85_155#_c_74_n N_VGND_c_416_n 5.09353e-19 $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_138 N_A_85_155#_c_95_p A_235_47# 0.00288179f $X=1.675 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_139 N_A2_M1003_g N_A1_c_199_n 4.63706e-19 $X=1.1 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A2_M1003_g N_A1_c_202_n 0.0634124f $X=1.1 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A2_M1007_g N_B1_M1000_g 0.0277908f $X=1.21 $Y=2.775 $X2=0 $Y2=0
cc_142 A2 N_B1_c_246_n 0.0020557f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A2_c_156_n N_B1_c_246_n 0.0123257f $X=1.16 $Y=1.5 $X2=0 $Y2=0
cc_144 N_A2_c_159_n N_B1_c_250_n 0.0123257f $X=1.16 $Y=2.005 $X2=0 $Y2=0
cc_145 N_A2_M1003_g B1 7.32324e-19 $X=1.1 $Y=0.445 $X2=0 $Y2=0
cc_146 A2 B1 0.06762f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A2_c_156_n B1 0.00205688f $X=1.16 $Y=1.5 $X2=0 $Y2=0
cc_148 N_A2_c_154_n N_B1_c_248_n 0.0123257f $X=1.16 $Y=1.84 $X2=0 $Y2=0
cc_149 N_A2_M1007_g N_VPWR_c_352_n 0.0066321f $X=1.21 $Y=2.775 $X2=0 $Y2=0
cc_150 N_A2_M1007_g N_VPWR_c_357_n 0.00547432f $X=1.21 $Y=2.775 $X2=0 $Y2=0
cc_151 N_A2_M1007_g N_VPWR_c_351_n 0.0101706f $X=1.21 $Y=2.775 $X2=0 $Y2=0
cc_152 N_A2_M1007_g N_A_257_491#_c_388_n 0.00444586f $X=1.21 $Y=2.775 $X2=0
+ $Y2=0
cc_153 N_A2_M1007_g N_A_257_491#_c_394_n 0.00195361f $X=1.21 $Y=2.775 $X2=0
+ $Y2=0
cc_154 N_A2_M1003_g N_VGND_c_411_n 0.00521725f $X=1.1 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A2_M1003_g N_VGND_c_413_n 0.00392525f $X=1.1 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A2_M1003_g N_VGND_c_415_n 0.00564108f $X=1.1 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A1_c_199_n N_B1_M1001_g 0.0171074f $X=2.795 $Y=0.897 $X2=0 $Y2=0
cc_158 N_A1_c_200_n N_B1_M1001_g 0.0218601f $X=1.55 $Y=0.93 $X2=0 $Y2=0
cc_159 N_A1_c_202_n N_B1_M1001_g 0.0144742f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_160 N_A1_c_199_n N_B1_c_246_n 0.00195789f $X=2.795 $Y=0.897 $X2=0 $Y2=0
cc_161 N_A1_c_200_n N_B1_c_246_n 0.00784828f $X=1.55 $Y=0.93 $X2=0 $Y2=0
cc_162 N_A1_c_199_n B1 0.0306225f $X=2.795 $Y=0.897 $X2=0 $Y2=0
cc_163 N_A1_c_200_n B1 0.00204224f $X=1.55 $Y=0.93 $X2=0 $Y2=0
cc_164 A1 N_B2_M1006_g 6.13893e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A1_c_203_n N_B2_M1006_g 0.0290513f $X=2.96 $Y=1.615 $X2=0 $Y2=0
cc_166 N_A1_c_199_n N_B2_M1004_g 0.0162908f $X=2.795 $Y=0.897 $X2=0 $Y2=0
cc_167 A1 N_B2_M1004_g 0.00741526f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A1_c_203_n N_B2_M1004_g 0.0148439f $X=2.96 $Y=1.615 $X2=0 $Y2=0
cc_169 N_A1_c_199_n B2 0.0330297f $X=2.795 $Y=0.897 $X2=0 $Y2=0
cc_170 A1 B2 0.0403864f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A1_c_203_n B2 0.00322652f $X=2.96 $Y=1.615 $X2=0 $Y2=0
cc_172 A1 N_B2_c_297_n 0.00114913f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A1_c_203_n N_B2_c_297_n 0.0216724f $X=2.96 $Y=1.615 $X2=0 $Y2=0
cc_174 N_A1_M1002_g N_VPWR_c_354_n 0.0115315f $X=2.75 $Y=2.775 $X2=0 $Y2=0
cc_175 A1 N_VPWR_c_354_n 0.0216553f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A1_c_203_n N_VPWR_c_354_n 0.00193108f $X=2.96 $Y=1.615 $X2=0 $Y2=0
cc_177 N_A1_M1002_g N_VPWR_c_357_n 0.00564095f $X=2.75 $Y=2.775 $X2=0 $Y2=0
cc_178 N_A1_M1002_g N_VPWR_c_351_n 0.00994131f $X=2.75 $Y=2.775 $X2=0 $Y2=0
cc_179 N_A1_M1002_g N_A_257_491#_c_387_n 0.00288292f $X=2.75 $Y=2.775 $X2=0
+ $Y2=0
cc_180 N_A1_c_199_n N_VGND_c_412_n 0.0243027f $X=2.795 $Y=0.897 $X2=0 $Y2=0
cc_181 N_A1_c_202_n N_VGND_c_413_n 0.00363059f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_182 N_A1_c_199_n N_VGND_c_415_n 0.02543f $X=2.795 $Y=0.897 $X2=0 $Y2=0
cc_183 N_A1_c_202_n N_VGND_c_415_n 0.00554824f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A1_c_204_n N_VGND_c_415_n 0.0199581f $X=3.035 $Y=1.015 $X2=0 $Y2=0
cc_185 N_B1_M1001_g N_B2_M1004_g 0.0879446f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_186 B1 N_B2_M1004_g 3.20853e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B1_c_248_n N_B2_M1004_g 0.00642384f $X=1.73 $Y=1.5 $X2=0 $Y2=0
cc_188 N_B1_M1001_g B2 0.002912f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_189 N_B1_c_246_n B2 0.00383036f $X=2 $Y=1.41 $X2=0 $Y2=0
cc_190 B1 B2 0.064006f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_191 N_B1_c_248_n B2 0.00340994f $X=1.73 $Y=1.5 $X2=0 $Y2=0
cc_192 N_B1_M1000_g N_B2_c_297_n 0.0293676f $X=1.64 $Y=2.775 $X2=0 $Y2=0
cc_193 B1 N_B2_c_297_n 2.98707e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_194 N_B1_c_248_n N_B2_c_297_n 0.017727f $X=1.73 $Y=1.5 $X2=0 $Y2=0
cc_195 N_B1_M1000_g N_VPWR_c_357_n 0.00357842f $X=1.64 $Y=2.775 $X2=0 $Y2=0
cc_196 N_B1_M1000_g N_VPWR_c_351_n 0.00566459f $X=1.64 $Y=2.775 $X2=0 $Y2=0
cc_197 N_B1_M1000_g N_A_257_491#_c_388_n 0.00606766f $X=1.64 $Y=2.775 $X2=0
+ $Y2=0
cc_198 N_B1_M1000_g N_A_257_491#_c_389_n 0.0088809f $X=1.64 $Y=2.775 $X2=0 $Y2=0
cc_199 N_B1_M1000_g N_A_257_491#_c_394_n 5.81207e-19 $X=1.64 $Y=2.775 $X2=0
+ $Y2=0
cc_200 N_B1_M1001_g N_VGND_c_412_n 0.00234139f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_201 N_B1_M1001_g N_VGND_c_413_n 0.00585385f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_202 N_B1_M1001_g N_VGND_c_415_n 0.00650373f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_203 N_B2_M1006_g N_VPWR_c_354_n 0.00110461f $X=2.18 $Y=2.775 $X2=0 $Y2=0
cc_204 N_B2_M1006_g N_VPWR_c_357_n 0.00357877f $X=2.18 $Y=2.775 $X2=0 $Y2=0
cc_205 N_B2_M1006_g N_VPWR_c_351_n 0.00606062f $X=2.18 $Y=2.775 $X2=0 $Y2=0
cc_206 N_B2_M1006_g N_A_257_491#_c_388_n 6.17513e-19 $X=2.18 $Y=2.775 $X2=0
+ $Y2=0
cc_207 N_B2_M1006_g N_A_257_491#_c_389_n 0.0152564f $X=2.18 $Y=2.775 $X2=0 $Y2=0
cc_208 N_B2_M1006_g N_A_257_491#_c_387_n 0.00277486f $X=2.18 $Y=2.775 $X2=0
+ $Y2=0
cc_209 B2 N_A_257_491#_c_387_n 0.00640836f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_210 N_B2_c_297_n N_A_257_491#_c_387_n 0.0036085f $X=2.3 $Y=1.89 $X2=0 $Y2=0
cc_211 N_B2_M1004_g N_VGND_c_412_n 0.0134198f $X=2.36 $Y=0.445 $X2=0 $Y2=0
cc_212 N_B2_M1004_g N_VGND_c_413_n 0.00486043f $X=2.36 $Y=0.445 $X2=0 $Y2=0
cc_213 N_B2_M1004_g N_VGND_c_415_n 0.00432544f $X=2.36 $Y=0.445 $X2=0 $Y2=0
cc_214 N_X_c_335_n N_VPWR_c_355_n 0.0334756f $X=0.425 $Y=2.61 $X2=0 $Y2=0
cc_215 N_X_M1005_s N_VPWR_c_351_n 0.00231914f $X=0.3 $Y=2.455 $X2=0 $Y2=0
cc_216 N_X_c_335_n N_VPWR_c_351_n 0.0194235f $X=0.425 $Y=2.61 $X2=0 $Y2=0
cc_217 N_X_M1008_s N_VGND_c_415_n 0.00277316f $X=0.195 $Y=0.235 $X2=0 $Y2=0
cc_218 N_X_c_333_n N_VGND_c_415_n 0.0148012f $X=0.36 $Y=0.43 $X2=0 $Y2=0
cc_219 N_X_c_333_n N_VGND_c_416_n 0.0235171f $X=0.36 $Y=0.43 $X2=0 $Y2=0
cc_220 N_VPWR_c_351_n N_A_257_491#_M1007_d 0.00223559f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_221 N_VPWR_c_351_n N_A_257_491#_M1006_d 0.00461528f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_357_n N_A_257_491#_c_389_n 0.0625908f $X=2.82 $Y=3.33 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_351_n N_A_257_491#_c_389_n 0.0385998f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_357_n N_A_257_491#_c_394_n 0.0188708f $X=2.82 $Y=3.33 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_351_n N_A_257_491#_c_394_n 0.0123968f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_354_n N_A_257_491#_c_387_n 0.0166895f $X=2.965 $Y=2.61 $X2=0
+ $Y2=0
cc_227 N_VGND_c_415_n A_235_47# 0.00169649f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_228 N_VGND_c_415_n A_415_47# 0.00289284f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
