* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21bo_lp A1 A2 B1_N VGND VNB VPB VPWR X
X0 X a_84_29# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR B1_N a_308_364# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VPWR A2 a_252_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_272_55# A1 a_84_29# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_252_409# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_594_55# B1_N a_308_364# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_84_29# a_308_364# a_436_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_114_55# a_84_29# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_84_29# a_114_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND A2 a_272_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_436_55# a_308_364# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND B1_N a_594_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_252_409# a_308_364# a_84_29# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
