* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR a_218_131# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1136e+12p pd=8.56e+06u as=3.528e+11p ps=3.08e+06u
M1001 VPWR B1 a_27_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.488e+11p ps=3.65e+06u
M1002 a_218_131# a_260_341# a_27_481# VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1003 X a_218_131# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_218_131# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=1.04695e+12p ps=8.86e+06u
M1005 a_480_367# A2_N a_260_341# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.696e+11p ps=1.81e+06u
M1006 a_260_341# A2_N VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1007 VGND A1_N a_260_341# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_481# B2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1_N a_480_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_218_131# B2 a_146_131# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1011 VGND a_260_341# a_218_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_218_131# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_146_131# B1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
