* File: sky130_fd_sc_lp__iso0n_lp2.pxi.spice
* Created: Fri Aug 28 10:40:25 2020
* 
x_PM_SKY130_FD_SC_LP__ISO0N_LP2%A N_A_c_46_n N_A_c_47_n N_A_c_48_n N_A_M1005_g
+ N_A_M1001_g A A N_A_c_51_n N_A_c_52_n PM_SKY130_FD_SC_LP__ISO0N_LP2%A
x_PM_SKY130_FD_SC_LP__ISO0N_LP2%SLEEP_B N_SLEEP_B_M1002_g N_SLEEP_B_M1000_g
+ SLEEP_B SLEEP_B N_SLEEP_B_c_89_n PM_SKY130_FD_SC_LP__ISO0N_LP2%SLEEP_B
x_PM_SKY130_FD_SC_LP__ISO0N_LP2%A_65_65# N_A_65_65#_M1001_s N_A_65_65#_M1005_d
+ N_A_65_65#_M1004_g N_A_65_65#_M1006_g N_A_65_65#_M1003_g N_A_65_65#_c_133_n
+ N_A_65_65#_c_140_n N_A_65_65#_c_134_n N_A_65_65#_c_135_n N_A_65_65#_c_136_n
+ N_A_65_65#_c_141_n N_A_65_65#_c_137_n N_A_65_65#_c_138_n
+ PM_SKY130_FD_SC_LP__ISO0N_LP2%A_65_65#
x_PM_SKY130_FD_SC_LP__ISO0N_LP2%VPWR N_VPWR_M1005_s N_VPWR_M1000_d
+ N_VPWR_c_208_n N_VPWR_c_209_n N_VPWR_c_210_n N_VPWR_c_211_n N_VPWR_c_212_n
+ VPWR N_VPWR_c_213_n N_VPWR_c_207_n PM_SKY130_FD_SC_LP__ISO0N_LP2%VPWR
x_PM_SKY130_FD_SC_LP__ISO0N_LP2%X N_X_M1003_d N_X_M1006_d N_X_c_236_n X X X X X
+ X X PM_SKY130_FD_SC_LP__ISO0N_LP2%X
x_PM_SKY130_FD_SC_LP__ISO0N_LP2%KAGND N_KAGND_M1002_d KAGND N_KAGND_c_260_n
+ PM_SKY130_FD_SC_LP__ISO0N_LP2%KAGND
x_PM_SKY130_FD_SC_LP__ISO0N_LP2%VGND VGND N_VGND_c_285_n N_VGND_c_286_n VGND
+ PM_SKY130_FD_SC_LP__ISO0N_LP2%VGND
cc_1 VNB N_A_c_46_n 0.0158885f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.03
cc_2 VNB N_A_c_47_n 0.0228007f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.03
cc_3 VNB N_A_c_48_n 0.0376152f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.625
cc_4 VNB N_A_M1005_g 0.00175608f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.545
cc_5 VNB N_A_M1001_g 0.0293808f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.535
cc_6 VNB N_A_c_51_n 0.0376278f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_7 VNB N_A_c_52_n 0.00518461f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_8 VNB N_SLEEP_B_M1002_g 0.0520069f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.625
cc_9 VNB SLEEP_B 0.00279774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_SLEEP_B_c_89_n 0.0129694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_65_65#_M1004_g 0.0210797f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.535
cc_12 VNB N_A_65_65#_M1006_g 0.0127966f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.475
cc_13 VNB N_A_65_65#_M1003_g 0.0247466f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_A_65_65#_c_133_n 0.00172021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_65_65#_c_134_n 0.0150724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_65_65#_c_135_n 0.0174385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_65_65#_c_136_n 0.00140514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_65_65#_c_137_n 0.0047913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_65_65#_c_138_n 0.0610127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_207_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_236_n 0.017334f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.535
cc_22 VNB X 0.0462956f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.55
cc_23 VNB KAGND 0.0263773f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.545
cc_24 VNB N_KAGND_c_260_n 0.00474886f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.955
cc_25 VNB N_VGND_c_285_n 0.155602f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.545
cc_26 VNB N_VGND_c_286_n 0.071067f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.535
cc_27 VPB N_A_M1005_g 0.0483436f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.545
cc_28 VPB N_A_c_52_n 0.00939201f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_29 VPB N_SLEEP_B_M1000_g 0.0280951f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.955
cc_30 VPB SLEEP_B 0.00349196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_SLEEP_B_c_89_n 0.0130627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_65_65#_M1006_g 0.0439168f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.475
cc_33 VPB N_A_65_65#_c_140_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_65_65#_c_141_n 0.00758198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_65_65#_c_137_n 0.00294098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_208_n 0.0129883f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.955
cc_37 VPB N_VPWR_c_209_n 0.0500396f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.535
cc_38 VPB N_VPWR_c_210_n 0.00432555f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.55
cc_39 VPB N_VPWR_c_211_n 0.020707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_212_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_41 VPB N_VPWR_c_213_n 0.0226325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_207_n 0.0538051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB X 0.0194633f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.55
cc_44 VPB X 0.0396102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB X 0.0201056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 N_A_c_48_n N_SLEEP_B_M1002_g 0.0100564f $X=0.635 $Y=1.625 $X2=0 $Y2=0
cc_47 N_A_M1001_g N_SLEEP_B_M1002_g 0.0489402f $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_48 N_A_c_51_n N_SLEEP_B_M1002_g 0.00279393f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_49 N_A_c_52_n N_SLEEP_B_M1002_g 4.10267e-19 $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_50 N_A_M1005_g N_SLEEP_B_M1000_g 0.014985f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_51 N_A_c_48_n SLEEP_B 3.67953e-19 $X=0.635 $Y=1.625 $X2=0 $Y2=0
cc_52 N_A_M1005_g N_SLEEP_B_c_89_n 0.0100564f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_53 N_A_M1001_g N_A_65_65#_c_133_n 0.00910508f $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_54 N_A_M1005_g N_A_65_65#_c_140_n 0.0171305f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_55 N_A_c_47_n N_A_65_65#_c_135_n 0.00699461f $X=0.455 $Y=1.03 $X2=0 $Y2=0
cc_56 N_A_M1001_g N_A_65_65#_c_135_n 0.01241f $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_57 N_A_c_52_n N_A_65_65#_c_135_n 0.010846f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_58 N_A_c_46_n N_A_65_65#_c_136_n 0.00708836f $X=0.61 $Y=1.03 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_A_65_65#_c_136_n 5.76998e-19 $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_60 N_A_c_51_n N_A_65_65#_c_136_n 8.02948e-19 $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_61 N_A_c_52_n N_A_65_65#_c_136_n 0.0236223f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_62 N_A_M1005_g N_A_65_65#_c_141_n 0.00421869f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_63 N_A_c_48_n N_A_65_65#_c_137_n 0.0059504f $X=0.635 $Y=1.625 $X2=0 $Y2=0
cc_64 N_A_M1005_g N_A_65_65#_c_137_n 0.0166116f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_65 N_A_c_51_n N_A_65_65#_c_137_n 9.98714e-19 $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_66 N_A_c_52_n N_A_65_65#_c_137_n 0.0336202f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_67 N_A_c_48_n N_VPWR_c_209_n 0.00219826f $X=0.635 $Y=1.625 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_VPWR_c_209_n 0.0270912f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_69 N_A_c_52_n N_VPWR_c_209_n 0.0226684f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_VPWR_c_210_n 9.45383e-19 $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_71 N_A_M1005_g N_VPWR_c_211_n 0.00741874f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_72 N_A_M1005_g N_VPWR_c_207_n 0.0131735f $X=0.635 $Y=2.545 $X2=0 $Y2=0
cc_73 N_A_M1001_g KAGND 0.00178747f $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_74 N_A_c_52_n KAGND 0.00897973f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_75 N_A_M1001_g N_KAGND_c_260_n 0.00117079f $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_VGND_c_285_n 0.0043929f $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_77 N_A_M1001_g N_VGND_c_286_n 0.00344318f $X=0.685 $Y=0.535 $X2=0 $Y2=0
cc_78 N_SLEEP_B_M1002_g N_A_65_65#_M1004_g 0.0172351f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_79 N_SLEEP_B_M1000_g N_A_65_65#_M1006_g 0.0166396f $X=1.165 $Y=2.545 $X2=0
+ $Y2=0
cc_80 SLEEP_B N_A_65_65#_M1006_g 0.0265505f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_81 N_SLEEP_B_c_89_n N_A_65_65#_M1006_g 0.0181444f $X=1.165 $Y=1.68 $X2=0
+ $Y2=0
cc_82 N_SLEEP_B_M1002_g N_A_65_65#_c_133_n 0.0035663f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_83 N_SLEEP_B_M1000_g N_A_65_65#_c_140_n 0.0144676f $X=1.165 $Y=2.545 $X2=0
+ $Y2=0
cc_84 N_SLEEP_B_M1002_g N_A_65_65#_c_134_n 0.0177824f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_85 SLEEP_B N_A_65_65#_c_134_n 0.0430509f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_86 N_SLEEP_B_c_89_n N_A_65_65#_c_134_n 0.00443904f $X=1.165 $Y=1.68 $X2=0
+ $Y2=0
cc_87 N_SLEEP_B_M1002_g N_A_65_65#_c_135_n 0.00193101f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_88 N_SLEEP_B_M1000_g N_A_65_65#_c_141_n 0.00408034f $X=1.165 $Y=2.545 $X2=0
+ $Y2=0
cc_89 SLEEP_B N_A_65_65#_c_141_n 0.00506068f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_90 N_SLEEP_B_c_89_n N_A_65_65#_c_141_n 0.00108331f $X=1.165 $Y=1.68 $X2=0
+ $Y2=0
cc_91 N_SLEEP_B_M1002_g N_A_65_65#_c_137_n 0.00637178f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_92 N_SLEEP_B_M1000_g N_A_65_65#_c_137_n 0.0035511f $X=1.165 $Y=2.545 $X2=0
+ $Y2=0
cc_93 SLEEP_B N_A_65_65#_c_137_n 0.0250969f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_94 N_SLEEP_B_c_89_n N_A_65_65#_c_137_n 0.00100302f $X=1.165 $Y=1.68 $X2=0
+ $Y2=0
cc_95 N_SLEEP_B_M1002_g N_A_65_65#_c_138_n 0.0267797f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_96 SLEEP_B N_A_65_65#_c_138_n 0.00482492f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_97 N_SLEEP_B_M1000_g N_VPWR_c_210_n 0.022456f $X=1.165 $Y=2.545 $X2=0 $Y2=0
cc_98 SLEEP_B N_VPWR_c_210_n 0.0272775f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_99 N_SLEEP_B_c_89_n N_VPWR_c_210_n 9.27233e-19 $X=1.165 $Y=1.68 $X2=0 $Y2=0
cc_100 N_SLEEP_B_M1000_g N_VPWR_c_211_n 0.00769046f $X=1.165 $Y=2.545 $X2=0
+ $Y2=0
cc_101 N_SLEEP_B_M1000_g N_VPWR_c_207_n 0.0134474f $X=1.165 $Y=2.545 $X2=0 $Y2=0
cc_102 SLEEP_B X 0.0200402f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_103 N_SLEEP_B_M1000_g X 2.76234e-19 $X=1.165 $Y=2.545 $X2=0 $Y2=0
cc_104 N_SLEEP_B_M1002_g KAGND 0.00276725f $X=1.075 $Y=0.535 $X2=0 $Y2=0
cc_105 N_SLEEP_B_M1002_g N_KAGND_c_260_n 0.00928031f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_106 N_SLEEP_B_M1002_g N_VGND_c_285_n 0.00419871f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_107 N_SLEEP_B_M1002_g N_VGND_c_286_n 0.00417651f $X=1.075 $Y=0.535 $X2=0
+ $Y2=0
cc_108 N_A_65_65#_c_141_n N_VPWR_c_209_n 0.0400865f $X=0.9 $Y=2.19 $X2=0 $Y2=0
cc_109 N_A_65_65#_M1006_g N_VPWR_c_210_n 0.0237304f $X=1.695 $Y=2.545 $X2=0
+ $Y2=0
cc_110 N_A_65_65#_c_141_n N_VPWR_c_210_n 0.069715f $X=0.9 $Y=2.19 $X2=0 $Y2=0
cc_111 N_A_65_65#_c_140_n N_VPWR_c_211_n 0.0273857f $X=0.9 $Y=2.9 $X2=0 $Y2=0
cc_112 N_A_65_65#_M1006_g N_VPWR_c_213_n 0.00769046f $X=1.695 $Y=2.545 $X2=0
+ $Y2=0
cc_113 N_A_65_65#_M1006_g N_VPWR_c_207_n 0.0141634f $X=1.695 $Y=2.545 $X2=0
+ $Y2=0
cc_114 N_A_65_65#_c_140_n N_VPWR_c_207_n 0.0153677f $X=0.9 $Y=2.9 $X2=0 $Y2=0
cc_115 N_A_65_65#_M1004_g N_X_c_236_n 0.00140521f $X=1.505 $Y=0.535 $X2=0 $Y2=0
cc_116 N_A_65_65#_M1003_g N_X_c_236_n 0.00933413f $X=1.895 $Y=0.535 $X2=0 $Y2=0
cc_117 N_A_65_65#_M1003_g X 0.0116481f $X=1.895 $Y=0.535 $X2=0 $Y2=0
cc_118 N_A_65_65#_c_134_n X 0.0164626f $X=1.555 $Y=1.11 $X2=0 $Y2=0
cc_119 N_A_65_65#_c_138_n X 0.022612f $X=1.695 $Y=1.202 $X2=0 $Y2=0
cc_120 N_A_65_65#_M1006_g X 0.0141811f $X=1.695 $Y=2.545 $X2=0 $Y2=0
cc_121 N_A_65_65#_M1006_g X 0.00574402f $X=1.695 $Y=2.545 $X2=0 $Y2=0
cc_122 N_A_65_65#_c_135_n A_152_65# 0.00131132f $X=0.47 $Y=0.535 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_65_65#_M1004_g KAGND 0.00366884f $X=1.505 $Y=0.535 $X2=0 $Y2=0
cc_124 N_A_65_65#_M1003_g KAGND 0.00721626f $X=1.895 $Y=0.535 $X2=0 $Y2=0
cc_125 N_A_65_65#_c_134_n KAGND 0.0244107f $X=1.555 $Y=1.11 $X2=0 $Y2=0
cc_126 N_A_65_65#_c_135_n KAGND 0.0434398f $X=0.47 $Y=0.535 $X2=0 $Y2=0
cc_127 N_A_65_65#_c_138_n KAGND 0.00160632f $X=1.695 $Y=1.202 $X2=0 $Y2=0
cc_128 N_A_65_65#_M1004_g N_KAGND_c_260_n 0.0080343f $X=1.505 $Y=0.535 $X2=0
+ $Y2=0
cc_129 N_A_65_65#_M1003_g N_KAGND_c_260_n 0.00140269f $X=1.895 $Y=0.535 $X2=0
+ $Y2=0
cc_130 N_A_65_65#_c_134_n N_KAGND_c_260_n 0.0270912f $X=1.555 $Y=1.11 $X2=0
+ $Y2=0
cc_131 N_A_65_65#_c_135_n N_KAGND_c_260_n 0.0162252f $X=0.47 $Y=0.535 $X2=0
+ $Y2=0
cc_132 N_A_65_65#_c_138_n N_KAGND_c_260_n 9.14374e-19 $X=1.695 $Y=1.202 $X2=0
+ $Y2=0
cc_133 N_A_65_65#_M1004_g N_VGND_c_285_n 0.00436071f $X=1.505 $Y=0.535 $X2=0
+ $Y2=0
cc_134 N_A_65_65#_M1003_g N_VGND_c_285_n 0.00472444f $X=1.895 $Y=0.535 $X2=0
+ $Y2=0
cc_135 N_A_65_65#_c_135_n N_VGND_c_285_n 0.00442112f $X=0.47 $Y=0.535 $X2=0
+ $Y2=0
cc_136 N_A_65_65#_M1004_g N_VGND_c_286_n 0.00468046f $X=1.505 $Y=0.535 $X2=0
+ $Y2=0
cc_137 N_A_65_65#_M1003_g N_VGND_c_286_n 0.0046928f $X=1.895 $Y=0.535 $X2=0
+ $Y2=0
cc_138 N_A_65_65#_c_135_n N_VGND_c_286_n 0.0206855f $X=0.47 $Y=0.535 $X2=0 $Y2=0
cc_139 N_VPWR_c_213_n X 0.0321458f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_140 N_VPWR_c_207_n X 0.0183848f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_141 N_VPWR_c_210_n X 0.0705123f $X=1.43 $Y=2.19 $X2=0 $Y2=0
cc_142 N_X_c_236_n KAGND 0.03854f $X=2.11 $Y=0.535 $X2=0 $Y2=0
cc_143 N_X_c_236_n N_KAGND_c_260_n 0.0110294f $X=2.11 $Y=0.535 $X2=0 $Y2=0
cc_144 N_X_c_236_n N_VGND_c_285_n 0.00355114f $X=2.11 $Y=0.535 $X2=0 $Y2=0
cc_145 N_X_c_236_n N_VGND_c_286_n 0.0176183f $X=2.11 $Y=0.535 $X2=0 $Y2=0
cc_146 A_152_65# KAGND 0.00339372f $X=0.76 $Y=0.325 $X2=0 $Y2=0
cc_147 KAGND A_316_65# 0.00642965f $X=0.07 $Y=0.44 $X2=-0.19 $Y2=-0.245
cc_148 KAGND N_VGND_c_285_n 0.205312f $X=0.07 $Y=0.44 $X2=0 $Y2=0
cc_149 N_KAGND_c_260_n N_VGND_c_285_n 0.00380629f $X=1.2 $Y=0.555 $X2=0 $Y2=0
cc_150 KAGND N_VGND_c_286_n 0.00684865f $X=0.07 $Y=0.44 $X2=0 $Y2=0
cc_151 N_KAGND_c_260_n N_VGND_c_286_n 0.0191853f $X=1.2 $Y=0.555 $X2=0 $Y2=0
