* NGSPICE file created from sky130_fd_sc_lp__a221o_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_334_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=8.001e+11p pd=6.31e+06u as=1.3104e+12p ps=9.64e+06u
M1001 VGND B2 a_739_49# VNB nshort w=840000u l=150000u
+  ad=1.1886e+12p pd=9.55e+06u as=2.688e+11p ps=2.32e+06u
M1002 a_653_367# B2 a_334_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=0p ps=0u
M1003 a_86_27# A1 a_356_53# VNB nshort w=840000u l=150000u
+  ad=4.578e+11p pd=4.45e+06u as=1.764e+11p ps=2.1e+06u
M1004 X a_86_27# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1005 a_334_367# B1 a_653_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_739_49# B1 a_86_27# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_334_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_356_53# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_86_27# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_653_367# C1 a_86_27# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1011 VGND a_86_27# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1012 X a_86_27# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_86_27# C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

