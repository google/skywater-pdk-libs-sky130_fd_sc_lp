# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__and3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.105000 0.815000 1.435000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.105000 1.340000 1.435000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 1.105000 1.775000 1.455000 ;
        RECT 1.515000 2.355000 1.775000 2.940000 ;
        RECT 1.575000 1.455000 1.775000 1.520000 ;
        RECT 1.595000 1.520000 1.775000 2.355000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 0.255000 2.795000 1.125000 ;
        RECT 2.495000 1.125000 2.795000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.145000  0.310000 0.620000 0.765000 ;
      RECT 0.145000  0.765000 2.125000 0.935000 ;
      RECT 0.145000  0.935000 0.315000 1.605000 ;
      RECT 0.145000  1.605000 1.425000 1.775000 ;
      RECT 0.145000  1.775000 0.565000 2.210000 ;
      RECT 0.735000  1.945000 1.015000 3.245000 ;
      RECT 1.185000  1.775000 1.425000 2.210000 ;
      RECT 1.740000  0.085000 2.070000 0.595000 ;
      RECT 1.945000  0.935000 2.125000 1.305000 ;
      RECT 1.945000  1.305000 2.325000 1.635000 ;
      RECT 1.945000  1.810000 2.325000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_lp__and3_1
END LIBRARY
