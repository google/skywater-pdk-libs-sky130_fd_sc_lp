* File: sky130_fd_sc_lp__mux4_1.pex.spice
* Created: Fri Aug 28 10:46:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX4_1%A1 2 5 9 11 12 13 14 19
c36 9 0 9.426e-20 $X=0.505 $Y=0.615
r37 19 21 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.4 $Y=1.375
+ $X2=0.4 $Y2=1.21
r38 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.375 $X2=0.385 $Y2=1.375
r39 13 14 9.51718 $w=4.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=2.035
r40 13 20 7.45941 $w=4.63e-07 $l=2.9e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=1.375
r41 12 20 2.05777 $w=4.63e-07 $l=8e-08 $layer=LI1_cond $X=0.317 $Y=1.295
+ $X2=0.317 $Y2=1.375
r42 9 21 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=0.505 $Y=0.615
+ $X2=0.505 $Y2=1.21
r43 5 11 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=2.805
+ $X2=0.475 $Y2=1.88
r44 2 11 44.5126 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.4 $Y=1.7 $X2=0.4
+ $Y2=1.88
r45 1 19 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=0.4 $Y=1.39 $X2=0.4
+ $Y2=1.375
r46 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=0.4 $Y=1.39 $X2=0.4
+ $Y2=1.7
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A0 3 7 11 12 13 14 15 20
r45 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.995
+ $Y=1.75 $X2=0.995 $Y2=1.75
r46 15 21 5.4981 $w=6.18e-07 $l=2.85e-07 $layer=LI1_cond $X=1.14 $Y=2.035
+ $X2=1.14 $Y2=1.75
r47 14 21 1.63978 $w=6.18e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.75
r48 13 14 7.13789 $w=6.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.14 $Y=1.295
+ $X2=1.14 $Y2=1.665
r49 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.995 $Y=2.09
+ $X2=0.995 $Y2=1.75
r50 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=2.09
+ $X2=0.995 $Y2=2.255
r51 10 20 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.585
+ $X2=0.995 $Y2=1.75
r52 7 10 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.985 $Y=0.615
+ $X2=0.985 $Y2=1.585
r53 3 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.905 $Y=2.805
+ $X2=0.905 $Y2=2.255
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_254_55# 1 2 9 11 12 15 17 22 25 29 31 34 37
+ 40 42 43 46 47 50 51
c150 51 0 1.71404e-19 $X=2.34 $Y=1.265
c151 47 0 1.82533e-19 $X=4.34 $Y=1.53
c152 46 0 4.96254e-20 $X=4.34 $Y=1.53
c153 42 0 3.86399e-20 $X=4.175 $Y=2.06
c154 40 0 8.85205e-20 $X=3.05 $Y=2.68
c155 17 0 3.8501e-19 $X=2.175 $Y=1.27
r156 50 53 17.1263 $w=5.63e-07 $l=5.05e-07 $layer=LI1_cond $X=2.537 $Y=1.265
+ $X2=2.537 $Y2=1.77
r157 50 52 7.0111 $w=5.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.537 $Y=1.265
+ $X2=2.537 $Y2=1.1
r158 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.34
+ $Y=1.265 $X2=2.34 $Y2=1.265
r159 47 59 49.3392 $w=5.95e-07 $l=1.65e-07 $layer=POLY_cond $X=4.472 $Y=1.53
+ $X2=4.472 $Y2=1.365
r160 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.34
+ $Y=1.53 $X2=4.34 $Y2=1.53
r161 44 46 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=4.305 $Y=1.975
+ $X2=4.305 $Y2=1.53
r162 42 44 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.175 $Y=2.06
+ $X2=4.305 $Y2=1.975
r163 42 43 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.175 $Y=2.06
+ $X2=3.175 $Y2=2.06
r164 38 43 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.03 $Y=2.06
+ $X2=3.175 $Y2=2.06
r165 38 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.03 $Y=2.06
+ $X2=2.735 $Y2=2.06
r166 38 40 21.2606 $w=2.88e-07 $l=5.35e-07 $layer=LI1_cond $X=3.03 $Y=2.145
+ $X2=3.03 $Y2=2.68
r167 37 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=1.975
+ $X2=2.735 $Y2=2.06
r168 37 53 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.735 $Y=1.975
+ $X2=2.735 $Y2=1.77
r169 34 52 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.69 $Y=0.805
+ $X2=2.69 $Y2=1.1
r170 27 29 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.765 $Y=2.14
+ $X2=4.765 $Y2=2.715
r171 25 59 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.32 $Y=0.795
+ $X2=4.32 $Y2=1.365
r172 22 27 20.4816 $w=3.53e-07 $l=3.60276e-07 $layer=POLY_cond $X=4.472 $Y=1.99
+ $X2=4.765 $Y2=2.14
r173 21 47 11.8696 $w=5.95e-07 $l=1.32e-07 $layer=POLY_cond $X=4.472 $Y=1.662
+ $X2=4.472 $Y2=1.53
r174 21 22 29.4941 $w=5.95e-07 $l=3.28e-07 $layer=POLY_cond $X=4.472 $Y=1.662
+ $X2=4.472 $Y2=1.99
r175 18 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.93 $Y=1.27
+ $X2=1.855 $Y2=1.27
r176 17 51 20.3982 $w=1.5e-07 $l=1.8747e-07 $layer=POLY_cond $X=2.175 $Y=1.27
+ $X2=2.34 $Y2=1.222
r177 17 18 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=2.175 $Y=1.27
+ $X2=1.93 $Y2=1.27
r178 13 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=1.27
r179 13 15 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=2.505
r180 11 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.78 $Y=1.27
+ $X2=1.855 $Y2=1.27
r181 11 12 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.78 $Y=1.27
+ $X2=1.42 $Y2=1.27
r182 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.345 $Y=1.195
+ $X2=1.42 $Y2=1.27
r183 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.345 $Y=1.195
+ $X2=1.345 $Y2=0.615
r184 2 40 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=2.47 $X2=3.05 $Y2=2.68
r185 1 34 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.595 $X2=2.725 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%S0 3 5 6 7 9 10 11 12 14 16 17 19 23 26 27 28
+ 32 33 35 36 37 40 43 44 49 50
c112 50 0 1.84933e-19 $X=3.565 $Y=1.29
r113 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.565
+ $Y=1.29 $X2=3.565 $Y2=1.29
r114 44 50 7.9441 $w=6.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.12 $Y=1.46
+ $X2=3.565 $Y2=1.46
r115 42 49 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.565 $Y=1.63
+ $X2=3.565 $Y2=1.29
r116 42 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.63
+ $X2=3.565 $Y2=1.795
r117 39 49 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.565 $Y=1.275
+ $X2=3.565 $Y2=1.29
r118 39 40 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.565 $Y=1.2
+ $X2=3.89 $Y2=1.2
r119 33 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.335 $Y=2.395
+ $X2=4.335 $Y2=2.715
r120 30 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.89 $Y=1.125
+ $X2=3.89 $Y2=1.2
r121 30 32 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.89 $Y=1.125
+ $X2=3.89 $Y2=0.795
r122 29 32 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.89 $Y=0.255
+ $X2=3.89 $Y2=0.795
r123 27 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.26 $Y=2.32
+ $X2=4.335 $Y2=2.395
r124 27 28 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.26 $Y=2.32
+ $X2=3.73 $Y2=2.32
r125 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.655 $Y=2.245
+ $X2=3.73 $Y2=2.32
r126 26 43 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.655 $Y=2.245
+ $X2=3.655 $Y2=1.795
r127 21 23 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.265 $Y=2.185
+ $X2=3.265 $Y2=2.68
r128 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=2.11
+ $X2=2.94 $Y2=2.11
r129 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.19 $Y=2.11
+ $X2=3.265 $Y2=2.185
r130 19 20 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.19 $Y=2.11
+ $X2=3.015 $Y2=2.11
r131 18 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=1.2
+ $X2=2.94 $Y2=1.2
r132 17 39 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.2
+ $X2=3.565 $Y2=1.2
r133 17 18 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.4 $Y=1.2
+ $X2=3.015 $Y2=1.2
r134 16 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=2.035
+ $X2=2.94 $Y2=2.11
r135 15 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=1.275
+ $X2=2.94 $Y2=1.2
r136 15 16 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.94 $Y=1.275
+ $X2=2.94 $Y2=2.035
r137 12 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=1.125
+ $X2=2.94 $Y2=1.2
r138 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.94 $Y=1.125
+ $X2=2.94 $Y2=0.805
r139 10 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=2.11
+ $X2=2.94 $Y2=2.11
r140 10 11 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.865 $Y=2.11
+ $X2=2.36 $Y2=2.11
r141 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.285 $Y=2.185
+ $X2=2.36 $Y2=2.11
r142 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.285 $Y=2.185
+ $X2=2.285 $Y2=2.505
r143 5 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.815 $Y=0.18
+ $X2=3.89 $Y2=0.255
r144 5 6 1007.59 $w=1.5e-07 $l=1.965e-06 $layer=POLY_cond $X=3.815 $Y=0.18
+ $X2=1.85 $Y2=0.18
r145 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.775 $Y=0.255
+ $X2=1.85 $Y2=0.18
r146 1 3 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.775 $Y=0.255
+ $X2=1.775 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A3 3 9 11 12 13 14 15 16 17 21 22
c54 22 0 3.81595e-20 $X=5.145 $Y=1.245
c55 3 0 3.35041e-19 $X=5.125 $Y=2.715
r56 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.145
+ $Y=1.245 $X2=5.145 $Y2=1.245
r57 16 17 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=5.087 $Y=1.295
+ $X2=5.087 $Y2=1.665
r58 16 22 2.02183 $w=2.83e-07 $l=5e-08 $layer=LI1_cond $X=5.087 $Y=1.295
+ $X2=5.087 $Y2=1.245
r59 14 15 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=5.252 $Y=0.77
+ $X2=5.252 $Y2=0.92
r60 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.145 $Y=1.585
+ $X2=5.145 $Y2=1.245
r61 12 13 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.585
+ $X2=5.145 $Y2=1.75
r62 11 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.08
+ $X2=5.145 $Y2=1.245
r63 11 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=5.235 $Y=1.08
+ $X2=5.235 $Y2=0.92
r64 9 14 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=5.27 $Y=0.445
+ $X2=5.27 $Y2=0.77
r65 3 13 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=5.125 $Y=2.715
+ $X2=5.125 $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A2 3 7 11 12 13 14 18
c45 18 0 1.62374e-19 $X=5.715 $Y=1.325
c46 13 0 5.41696e-20 $X=5.52 $Y=1.295
c47 12 0 3.81595e-20 $X=5.715 $Y=1.83
r48 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.715
+ $Y=1.325 $X2=5.715 $Y2=1.325
r49 14 19 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=5.64 $Y=1.665
+ $X2=5.64 $Y2=1.325
r50 13 19 0.747549 $w=4.78e-07 $l=3e-08 $layer=LI1_cond $X=5.64 $Y=1.295
+ $X2=5.64 $Y2=1.325
r51 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.715 $Y=1.665
+ $X2=5.715 $Y2=1.325
r52 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.665
+ $X2=5.715 $Y2=1.83
r53 10 18 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.16
+ $X2=5.715 $Y2=1.325
r54 7 10 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=5.78 $Y=0.445
+ $X2=5.78 $Y2=1.16
r55 3 12 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=5.625 $Y=2.715
+ $X2=5.625 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%S1 3 7 9 11 13 16 19 21 22 23 26 27
c69 9 0 1.22512e-19 $X=8.025 $Y=1.35
r70 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.96
+ $Y=1.44 $X2=6.96 $Y2=1.44
r71 23 27 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.44
r72 20 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.96 $Y=1.78
+ $X2=6.96 $Y2=1.44
r73 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.96 $Y=1.78
+ $X2=6.96 $Y2=1.945
r74 18 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.96 $Y=1.425
+ $X2=6.96 $Y2=1.44
r75 18 19 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=6.96 $Y=1.425
+ $X2=6.96 $Y2=1.35
r76 14 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.1 $Y=1.425 $X2=8.1
+ $Y2=1.35
r77 14 16 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.1 $Y=1.425 $X2=8.1
+ $Y2=2.045
r78 11 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.1 $Y=1.275 $X2=8.1
+ $Y2=1.35
r79 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.1 $Y=1.275 $X2=8.1
+ $Y2=0.955
r80 10 19 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=6.96 $Y2=1.35
r81 9 22 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.025 $Y=1.35 $X2=8.1
+ $Y2=1.35
r82 9 10 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=8.025 $Y=1.35 $X2=7.125
+ $Y2=1.35
r83 7 21 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=6.87 $Y=2.435
+ $X2=6.87 $Y2=1.945
r84 1 19 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.87 $Y=1.275
+ $X2=6.96 $Y2=1.35
r85 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=6.87 $Y=1.275 $X2=6.87
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_1245_21# 1 2 10 11 12 13 14 15 17 20 22 25
+ 27 28 29 30 33 34 36 37 40 44 46 48 49
c130 37 0 1.62374e-19 $X=6.555 $Y=1.1
c131 36 0 3.22935e-20 $X=7 $Y=1.1
c132 33 0 2.25236e-20 $X=6.39 $Y=1.29
r133 49 54 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.485 $Y=2.945
+ $X2=7.485 $Y2=3.06
r134 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.485
+ $Y=2.945 $X2=7.485 $Y2=2.945
r135 46 48 9.18048 $w=2.93e-07 $l=2.35e-07 $layer=LI1_cond $X=7.25 $Y=2.927
+ $X2=7.485 $Y2=2.927
r136 42 44 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=7.125 $Y=1.015
+ $X2=7.125 $Y2=0.805
r137 38 46 6.84433 $w=2.95e-07 $l=2.26892e-07 $layer=LI1_cond $X=7.085 $Y=2.78
+ $X2=7.25 $Y2=2.927
r138 38 40 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=7.085 $Y=2.78
+ $X2=7.085 $Y2=2.48
r139 36 42 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7 $Y=1.1
+ $X2=7.125 $Y2=1.015
r140 36 37 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7 $Y=1.1 $X2=6.555
+ $Y2=1.1
r141 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.39
+ $Y=1.29 $X2=6.39 $Y2=1.29
r142 31 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.555 $Y2=1.1
r143 31 33 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.39 $Y2=1.29
r144 28 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.39 $Y=1.63
+ $X2=6.39 $Y2=1.29
r145 28 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.39 $Y=1.63
+ $X2=6.39 $Y2=1.795
r146 27 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.39 $Y=1.125
+ $X2=6.39 $Y2=1.29
r147 24 25 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=9.02 $Y=0.255
+ $X2=9.02 $Y2=1.275
r148 23 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.605 $Y=1.35
+ $X2=8.53 $Y2=1.35
r149 22 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.945 $Y=1.35
+ $X2=9.02 $Y2=1.275
r150 22 23 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.945 $Y=1.35
+ $X2=8.605 $Y2=1.35
r151 18 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.53 $Y=1.425
+ $X2=8.53 $Y2=1.35
r152 18 20 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.53 $Y=1.425
+ $X2=8.53 $Y2=2.045
r153 15 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.53 $Y=1.275
+ $X2=8.53 $Y2=1.35
r154 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.53 $Y=1.275
+ $X2=8.53 $Y2=0.955
r155 13 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.32 $Y=3.06
+ $X2=7.485 $Y2=3.06
r156 13 14 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=7.32 $Y=3.06
+ $X2=6.375 $Y2=3.06
r157 11 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.945 $Y=0.18
+ $X2=9.02 $Y2=0.255
r158 11 12 1317.81 $w=1.5e-07 $l=2.57e-06 $layer=POLY_cond $X=8.945 $Y=0.18
+ $X2=6.375 $Y2=0.18
r159 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.3 $Y=2.985
+ $X2=6.375 $Y2=3.06
r160 10 29 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=6.3 $Y=2.985
+ $X2=6.3 $Y2=1.795
r161 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.3 $Y=0.255
+ $X2=6.375 $Y2=0.18
r162 7 27 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.3 $Y=0.255 $X2=6.3
+ $Y2=1.125
r163 2 40 600 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=2.225 $X2=7.085 $Y2=2.48
r164 1 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.945
+ $Y=0.595 $X2=7.085 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_1635_149# 1 2 9 12 16 20 24 25 27 29
r42 25 30 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.492 $Y=1.51
+ $X2=9.492 $Y2=1.675
r43 25 29 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.492 $Y=1.51
+ $X2=9.492 $Y2=1.345
r44 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.47
+ $Y=1.51 $X2=9.47 $Y2=1.51
r45 22 27 0.0301287 $w=3.3e-07 $l=1.13e-07 $layer=LI1_cond $X=8.445 $Y=1.51
+ $X2=8.332 $Y2=1.51
r46 22 24 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=8.445 $Y=1.51
+ $X2=9.47 $Y2=1.51
r47 18 27 7.07379 $w=2.22e-07 $l=1.65997e-07 $layer=LI1_cond $X=8.33 $Y=1.675
+ $X2=8.332 $Y2=1.51
r48 18 20 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=8.33 $Y=1.675
+ $X2=8.33 $Y2=2.045
r49 14 27 7.07379 $w=2.22e-07 $l=1.65e-07 $layer=LI1_cond $X=8.332 $Y=1.345
+ $X2=8.332 $Y2=1.51
r50 14 16 19.9757 $w=2.23e-07 $l=3.9e-07 $layer=LI1_cond $X=8.332 $Y=1.345
+ $X2=8.332 $Y2=0.955
r51 12 30 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.605 $Y=2.465
+ $X2=9.605 $Y2=1.675
r52 9 29 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.605 $Y=0.815
+ $X2=9.605 $Y2=1.345
r53 2 20 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.175
+ $Y=1.835 $X2=8.315 $Y2=2.045
r54 1 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.175
+ $Y=0.745 $X2=8.315 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_27_519# 1 2 9 11 12 13
r21 13 16 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=1.605 $Y=2.43
+ $X2=1.605 $Y2=2.51
r22 11 13 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.475 $Y=2.43
+ $X2=1.605 $Y2=2.43
r23 11 12 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=1.475 $Y=2.43
+ $X2=0.355 $Y2=2.43
r24 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=2.515
+ $X2=0.355 $Y2=2.43
r25 7 9 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.225 $Y=2.515
+ $X2=0.225 $Y2=2.805
r26 2 16 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=2.295 $X2=1.64 $Y2=2.51
r27 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.595 $X2=0.26 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%VPWR 1 2 3 4 5 18 22 26 28 32 36 40 42 47 55
+ 60 70 71 74 77 80 83 86
c98 32 0 2.25236e-20 $X=6.585 $Y=2.48
r99 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r100 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r102 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r103 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 71 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r106 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r107 68 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.555 $Y=3.33
+ $X2=9.39 $Y2=3.33
r108 68 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.555 $Y=3.33
+ $X2=9.84 $Y2=3.33
r109 67 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r110 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r111 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r112 64 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r114 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 61 83 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.75 $Y=3.33
+ $X2=6.58 $Y2=3.33
r116 61 63 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.75 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 60 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=9.39 $Y2=3.33
r118 60 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=8.88 $Y2=3.33
r119 56 77 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.495 $Y2=3.33
r120 56 58 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 55 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.285 $Y=3.33
+ $X2=5.41 $Y2=3.33
r122 55 58 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.285 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 54 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 51 54 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 51 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 50 53 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 48 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r130 48 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 47 77 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.495 $Y2=3.33
r132 47 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r133 45 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 42 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r136 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 40 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r138 40 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r139 40 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r140 36 39 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=9.39 $Y=1.98
+ $X2=9.39 $Y2=2.95
r141 34 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=3.33
r142 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=2.95
r143 30 83 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=3.245
+ $X2=6.58 $Y2=3.33
r144 30 32 25.93 $w=3.38e-07 $l=7.65e-07 $layer=LI1_cond $X=6.58 $Y=3.245
+ $X2=6.58 $Y2=2.48
r145 29 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.535 $Y=3.33
+ $X2=5.41 $Y2=3.33
r146 28 83 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.58 $Y2=3.33
r147 28 29 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=5.535 $Y2=3.33
r148 24 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.41 $Y2=3.33
r149 24 26 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.41 $Y2=2.78
r150 20 77 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=3.33
r151 20 22 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=2.68
r152 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r153 16 18 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.805
r154 5 39 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.835 $X2=9.39 $Y2=2.95
r155 5 36 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.835 $X2=9.39 $Y2=1.98
r156 4 32 600 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_PDIFF $count=1 $X=6.45
+ $Y=2.225 $X2=6.585 $Y2=2.48
r157 3 26 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=2.505 $X2=5.385 $Y2=2.78
r158 2 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.47 $X2=3.48 $Y2=2.68
r159 1 18 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.595 $X2=0.69 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_196_519# 1 2 7 11 14
c23 11 0 1.71404e-19 $X=2.5 $Y=2.505
r24 14 16 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=1.155 $Y=2.85
+ $X2=1.155 $Y2=2.95
r25 9 11 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=2.535 $Y=2.865
+ $X2=2.535 $Y2=2.505
r26 8 16 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.285 $Y=2.95
+ $X2=1.155 $Y2=2.95
r27 7 9 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.405 $Y=2.95
+ $X2=2.535 $Y2=2.865
r28 7 8 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=2.405 $Y=2.95
+ $X2=1.285 $Y2=2.95
r29 2 11 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=2.295 $X2=2.5 $Y2=2.505
r30 1 14 600 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.595 $X2=1.12 $Y2=2.85
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_284_81# 1 2 3 4 13 19 23 24 27 30 34 35 38
+ 41 42 45 48
c135 48 0 3.22935e-20 $X=7.915 $Y=1.88
c136 41 0 1.22512e-19 $X=7.92 $Y=2.035
c137 38 0 1.86083e-19 $X=2.16 $Y=2.035
c138 35 0 2.87447e-19 $X=2.305 $Y=2.035
r139 42 48 8.18908 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.915 $Y=2.035
+ $X2=7.915 $Y2=1.88
r140 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r141 38 46 4.27653 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.105 $Y2=2.17
r142 38 45 6.63084 $w=3.98e-07 $l=9.5e-08 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.105 $Y2=1.94
r143 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r144 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r145 34 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r146 34 35 6.76979 $w=1.4e-07 $l=5.47e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=2.305 $Y2=2.035
r147 30 32 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.56 $Y=0.7
+ $X2=1.56 $Y2=0.92
r148 25 27 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=8.762 $Y=0.62
+ $X2=8.762 $Y2=0.955
r149 23 25 6.95328 $w=2.3e-07 $l=1.9625e-07 $layer=LI1_cond $X=8.615 $Y=0.505
+ $X2=8.762 $Y2=0.62
r150 23 24 28.31 $w=2.28e-07 $l=5.65e-07 $layer=LI1_cond $X=8.615 $Y=0.505
+ $X2=8.05 $Y2=0.505
r151 21 24 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.965 $Y=0.62
+ $X2=8.05 $Y2=0.505
r152 21 48 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=7.965 $Y=0.62
+ $X2=7.965 $Y2=1.88
r153 19 46 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.07 $Y=2.505
+ $X2=2.07 $Y2=2.17
r154 15 45 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.99 $Y=1.005 $X2=1.99
+ $Y2=1.94
r155 14 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=0.92
+ $X2=1.56 $Y2=0.92
r156 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.905 $Y=0.92
+ $X2=1.99 $Y2=1.005
r157 13 14 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.905 $Y=0.92
+ $X2=1.725 $Y2=0.92
r158 4 42 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.835 $X2=7.885 $Y2=2.045
r159 3 19 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=2.295 $X2=2.07 $Y2=2.505
r160 2 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.605
+ $Y=0.745 $X2=8.745 $Y2=0.955
r161 1 30 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.42
+ $Y=0.405 $X2=1.56 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_799_501# 1 2 9 11 12 14 15 16 19
r47 17 19 10.372 $w=2.98e-07 $l=2.7e-07 $layer=LI1_cond $X=5.855 $Y=2.445
+ $X2=5.855 $Y2=2.715
r48 15 17 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=5.705 $Y=2.36
+ $X2=5.855 $Y2=2.445
r49 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.705 $Y=2.36
+ $X2=5.115 $Y2=2.36
r50 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.03 $Y=2.445
+ $X2=5.115 $Y2=2.36
r51 13 14 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.03 $Y=2.445
+ $X2=5.03 $Y2=2.905
r52 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.945 $Y=2.99
+ $X2=5.03 $Y2=2.905
r53 11 12 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.945 $Y=2.99
+ $X2=4.205 $Y2=2.99
r54 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.08 $Y=2.905
+ $X2=4.205 $Y2=2.99
r55 7 9 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=4.08 $Y=2.905
+ $X2=4.08 $Y2=2.71
r56 2 19 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=2.505 $X2=5.84 $Y2=2.715
r57 1 9 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=3.995
+ $Y=2.505 $X2=4.12 $Y2=2.71
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_793_117# 1 2 3 4 15 17 18 20 22 23 25 28 30
+ 31 32 35 40 42 43 50 52
c134 40 0 1.92606e-19 $X=4.69 $Y=2.63
c135 18 0 1.82533e-19 $X=4.2 $Y=1.1
c136 15 0 1.77638e-19 $X=4.105 $Y=0.79
r137 47 50 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=7.515 $Y=0.955
+ $X2=7.615 $Y2=0.955
r138 43 45 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.53 $Y=2.02 $X2=6.53
+ $Y2=2.12
r139 38 40 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=4.55 $Y=2.63
+ $X2=4.69 $Y2=2.63
r140 33 35 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=8.73 $Y=2.38
+ $X2=8.73 $Y2=2.045
r141 31 33 6.82051 $w=2.3e-07 $l=1.67929e-07 $layer=LI1_cond $X=8.61 $Y=2.495
+ $X2=8.73 $Y2=2.38
r142 31 32 50.6073 $w=2.28e-07 $l=1.01e-06 $layer=LI1_cond $X=8.61 $Y=2.495
+ $X2=7.6 $Y2=2.495
r143 30 32 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.515 $Y=2.38
+ $X2=7.6 $Y2=2.495
r144 29 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=2.205
+ $X2=7.515 $Y2=2.12
r145 29 30 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.515 $Y=2.205
+ $X2=7.515 $Y2=2.38
r146 28 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=2.035
+ $X2=7.515 $Y2=2.12
r147 27 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.515 $Y=1.12
+ $X2=7.515 $Y2=0.955
r148 27 28 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.515 $Y=1.12
+ $X2=7.515 $Y2=2.035
r149 26 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.615 $Y=2.12
+ $X2=6.53 $Y2=2.12
r150 25 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=2.12
+ $X2=7.515 $Y2=2.12
r151 25 26 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=7.43 $Y=2.12
+ $X2=6.615 $Y2=2.12
r152 24 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.775 $Y=2.02
+ $X2=4.69 $Y2=2.02
r153 23 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.445 $Y=2.02
+ $X2=6.53 $Y2=2.02
r154 23 24 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=6.445 $Y=2.02
+ $X2=4.775 $Y2=2.02
r155 22 40 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.69 $Y=2.525
+ $X2=4.69 $Y2=2.63
r156 21 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=2.105
+ $X2=4.69 $Y2=2.02
r157 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.69 $Y=2.105
+ $X2=4.69 $Y2=2.525
r158 20 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=1.935
+ $X2=4.69 $Y2=2.02
r159 19 20 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.69 $Y=1.185
+ $X2=4.69 $Y2=1.935
r160 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.605 $Y=1.1
+ $X2=4.69 $Y2=1.185
r161 17 18 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.605 $Y=1.1
+ $X2=4.2 $Y2=1.1
r162 13 18 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=4.087 $Y=1.015
+ $X2=4.2 $Y2=1.1
r163 13 15 11.5244 $w=2.23e-07 $l=2.25e-07 $layer=LI1_cond $X=4.087 $Y=1.015
+ $X2=4.087 $Y2=0.79
r164 4 35 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.605
+ $Y=1.835 $X2=8.745 $Y2=2.045
r165 3 38 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=2.505 $X2=4.55 $Y2=2.63
r166 2 50 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=7.49
+ $Y=0.745 $X2=7.615 $Y2=0.955
r167 1 15 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.585 $X2=4.105 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%X 1 2 7 8 9 10 11 12 13
r10 13 39 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.86 $Y=2.775
+ $X2=9.86 $Y2=2.91
r11 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.86 $Y=2.405
+ $X2=9.86 $Y2=2.775
r12 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.86 $Y=1.98
+ $X2=9.86 $Y2=2.405
r13 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.86 $Y=1.665
+ $X2=9.86 $Y2=1.98
r14 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.86 $Y=1.295
+ $X2=9.86 $Y2=1.665
r15 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.86 $Y=0.925 $X2=9.86
+ $Y2=1.295
r16 7 8 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.86 $Y=0.54 $X2=9.86
+ $Y2=0.925
r17 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=2.91
r18 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=1.98
r19 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.68
+ $Y=0.395 $X2=9.82 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_33_81# 1 2 9 11 12 14 15 16 17
c44 16 0 9.426e-20 $X=1.225 $Y=0.35
r45 17 20 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.06 $Y=0.35
+ $X2=2.06 $Y2=0.555
r46 15 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0.35
+ $X2=2.06 $Y2=0.35
r47 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.895 $Y=0.35
+ $X2=1.225 $Y2=0.35
r48 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.14 $Y=0.435
+ $X2=1.225 $Y2=0.35
r49 13 14 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.14 $Y=0.435
+ $X2=1.14 $Y2=0.815
r50 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.055 $Y=0.9
+ $X2=1.14 $Y2=0.815
r51 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.055 $Y=0.9
+ $X2=0.385 $Y2=0.9
r52 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.255 $Y=0.815
+ $X2=0.385 $Y2=0.9
r53 7 9 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=0.255 $Y=0.815 $X2=0.255
+ $Y2=0.615
r54 2 20 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=1.85
+ $Y=0.405 $X2=2.06 $Y2=0.555
r55 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.405 $X2=0.29 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 39 41 46
+ 54 66 75 76 79 82 85 88
r104 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r105 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r106 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r107 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r108 76 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r109 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r110 73 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.555 $Y=0 $X2=9.39
+ $Y2=0
r111 73 75 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.555 $Y=0
+ $X2=9.84 $Y2=0
r112 72 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r113 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r114 69 72 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r115 68 71 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.88
+ $Y2=0
r116 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r117 66 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=0 $X2=9.39
+ $Y2=0
r118 66 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.225 $Y=0 $X2=8.88
+ $Y2=0
r119 65 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r120 65 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=5.52
+ $Y2=0
r121 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r122 62 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.72 $Y=0 $X2=5.555
+ $Y2=0
r123 62 64 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.72 $Y=0 $X2=6.48
+ $Y2=0
r124 58 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r125 57 60 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r126 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r127 55 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=3.155
+ $Y2=0
r128 55 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=3.6
+ $Y2=0
r129 54 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.39 $Y=0 $X2=5.555
+ $Y2=0
r130 54 60 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.39 $Y=0 $X2=5.04
+ $Y2=0
r131 53 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r132 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r133 50 53 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r134 50 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r135 49 52 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r136 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r137 47 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.72
+ $Y2=0
r138 47 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.2
+ $Y2=0
r139 46 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.155
+ $Y2=0
r140 46 52 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.64
+ $Y2=0
r141 44 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r142 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r143 41 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.72
+ $Y2=0
r144 41 43 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0
+ $X2=0.24 $Y2=0
r145 39 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r146 39 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r147 39 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r148 37 64 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.49 $Y=0 $X2=6.48
+ $Y2=0
r149 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.49 $Y=0 $X2=6.655
+ $Y2=0
r150 36 68 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.96
+ $Y2=0
r151 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.655
+ $Y2=0
r152 32 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=0.085
+ $X2=9.39 $Y2=0
r153 32 34 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=9.39 $Y=0.085
+ $X2=9.39 $Y2=0.54
r154 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.655 $Y=0.085
+ $X2=6.655 $Y2=0
r155 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.655 $Y=0.085
+ $X2=6.655 $Y2=0.76
r156 24 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.555 $Y=0.085
+ $X2=5.555 $Y2=0
r157 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.555 $Y=0.085
+ $X2=5.555 $Y2=0.36
r158 20 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=0.085
+ $X2=3.155 $Y2=0
r159 20 22 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=3.155 $Y=0.085
+ $X2=3.155 $Y2=0.805
r160 16 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r161 16 18 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.53
r162 5 34 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=9.265
+ $Y=0.395 $X2=9.39 $Y2=0.54
r163 4 30 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=6.53
+ $Y=0.595 $X2=6.655 $Y2=0.76
r164 3 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.235 $X2=5.555 $Y2=0.36
r165 2 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.595 $X2=3.155 $Y2=0.805
r166 1 18 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.405 $X2=0.72 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_710_117# 1 2 9 12 14 15
r26 14 15 8.88925 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=0.365
+ $X2=4.89 $Y2=0.365
r27 12 15 63.3349 $w=1.88e-07 $l=1.085e-06 $layer=LI1_cond $X=3.805 $Y=0.35
+ $X2=4.89 $Y2=0.35
r28 7 12 7.24045 $w=1.9e-07 $l=1.89642e-07 $layer=LI1_cond $X=3.657 $Y=0.445
+ $X2=3.805 $Y2=0.35
r29 7 9 13.4777 $w=2.93e-07 $l=3.45e-07 $layer=LI1_cond $X=3.657 $Y=0.445
+ $X2=3.657 $Y2=0.79
r30 2 14 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.235 $X2=5.055 $Y2=0.38
r31 1 9 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.585 $X2=3.675 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_1%A_879_117# 1 2 7 11 16
r30 14 16 8.49442 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=0.73
+ $X2=4.7 $Y2=0.73
r31 9 11 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.025 $Y=0.645
+ $X2=6.025 $Y2=0.44
r32 7 9 7.01501 $w=2e-07 $l=1.78115e-07 $layer=LI1_cond $X=5.89 $Y=0.745
+ $X2=6.025 $Y2=0.645
r33 7 16 65.9909 $w=1.98e-07 $l=1.19e-06 $layer=LI1_cond $X=5.89 $Y=0.745
+ $X2=4.7 $Y2=0.745
r34 2 11 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.855
+ $Y=0.235 $X2=5.995 $Y2=0.44
r35 1 14 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.395
+ $Y=0.585 $X2=4.535 $Y2=0.745
.ends

