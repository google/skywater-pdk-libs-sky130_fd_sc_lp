* File: sky130_fd_sc_lp__nor2b_4.spice
* Created: Wed Sep  2 10:08:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor2b_4.pex.spice"
.subckt sky130_fd_sc_lp__nor2b_4  VNB VPB B_N A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_B_N_M1012_g N_A_60_47#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.2226 PD=1.2 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75003.7
+ A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1012_d N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84 AD=0.1512
+ AS=0.1176 PD=1.2 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.7 SB=75003.2
+ A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1001_s N_A_60_47#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1006 N_Y_M1006_d N_A_60_47#_M1006_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75001.9 A=0.126
+ P=1.98 MULT=1
MM1009 N_VGND_M1002_d N_A_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4 SB=75001.5 A=0.126
+ P=1.98 MULT=1
MM1010 N_Y_M1009_s N_A_60_47#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1017 N_Y_M1017_d N_A_60_47#_M1017_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_A_M1016_g N_Y_M1017_d VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_B_N_M1013_g N_A_60_47#_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.3339 PD=1.62 PS=3.05 NRD=9.3772 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1000 N_A_245_367#_M1000_d N_A_M1000_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75000.7
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1003 N_A_245_367#_M1000_d N_A_60_47#_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1007 N_A_245_367#_M1007_d N_A_60_47#_M1007_g N_Y_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1005 N_A_245_367#_M1007_d N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75001.9
+ A=0.189 P=2.82 MULT=1
MM1014 N_A_245_367#_M1014_d N_A_M1014_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_A_245_367#_M1014_d N_A_60_47#_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_A_245_367#_M1011_d N_A_60_47#_M1011_g N_Y_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_245_367#_M1011_d N_A_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__nor2b_4.pxi.spice"
*
.ends
*
*
