* File: sky130_fd_sc_lp__sdfstp_2.spice
* Created: Wed Sep  2 10:35:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfstp_2.pex.spice"
.subckt sky130_fd_sc_lp__sdfstp_2  VNB VPB SCD D SCE CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1022 A_172_121# N_SCD_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1011 N_A_244_121#_M1011_d N_SCE_M1011_g A_172_121# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 A_330_121# N_D_M1015_g N_A_244_121#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_358_429#_M1009_g A_330_121# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0441 PD=1.04 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1026 N_A_358_429#_M1026_d N_SCE_M1026_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1302 PD=1.37 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_CLK_M1010_g N_A_794_47#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1023 N_A_963_47#_M1023_d N_A_794_47#_M1023_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1034 N_A_1237_55#_M1034_d N_A_794_47#_M1034_g N_A_244_121#_M1034_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.3174 PD=0.7 PS=2.37 NRD=0 NRS=101.424 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1035 A_1323_55# N_A_963_47#_M1035_g N_A_1237_55#_M1034_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1038 N_VGND_M1038_d N_A_1365_29#_M1038_g A_1323_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 A_1608_125# N_A_1237_55#_M1024_g N_A_1365_29#_M1024_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1281 PD=0.63 PS=1.45 NRD=14.28 NRS=11.424 M=1 R=2.8
+ SA=75000.2 SB=75004.6 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_SET_B_M1027_g A_1608_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.207345 AS=0.0441 PD=1.39075 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75004.2 A=0.063 P=1.14 MULT=1
MM1013 A_1933_125# N_A_1237_55#_M1013_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.315955 PD=0.85 PS=2.11925 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_1998_463#_M1008_d N_A_963_47#_M1008_g A_1933_125# VNB NSHORT L=0.15
+ W=0.64 AD=0.224966 AS=0.0672 PD=1.52151 PS=0.85 NRD=33.276 NRS=9.372 M=1
+ R=4.26667 SA=75001.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1002 A_2159_125# N_A_794_47#_M1002_g N_A_1998_463#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.05775 AS=0.147634 PD=0.695 PS=0.998491 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75003 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1016 A_2244_125# N_A_2214_99#_M1016_g A_2159_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.05775 PD=0.96 PS=0.695 NRD=61.428 NRS=23.568 M=1 R=2.8
+ SA=75003.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_SET_B_M1019_g A_2244_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1134 PD=0.81 PS=0.96 NRD=0 NRS=61.428 M=1 R=2.8 SA=75004.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1031 N_A_2214_99#_M1031_d N_A_1998_463#_M1031_g N_VGND_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=31.428 M=1 R=2.8
+ SA=75004.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_1998_463#_M1006_g N_A_2686_131#_M1006_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0875 AS=0.1113 PD=0.8 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1006_d N_A_2686_131#_M1021_g N_Q_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.175 AS=0.1176 PD=1.6 PS=1.12 NRD=4.284 NRS=0 M=1 R=5.6 SA=75000.4
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1036 N_VGND_M1036_d N_A_2686_131#_M1036_g N_Q_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1037 N_VPWR_M1037_d N_SCD_M1037_g N_A_39_481#_M1037_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1017 A_208_481# N_SCE_M1017_g N_VPWR_M1037_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1018 N_A_244_121#_M1018_d N_D_M1018_g A_208_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=16.9223 NRS=15.3857 M=1 R=4.26667
+ SA=75001 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1033 N_A_39_481#_M1033_d N_A_358_429#_M1033_g N_A_244_121#_M1018_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=16.9223 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_A_358_429#_M1014_d N_SCE_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.3424 PD=1.81 PS=2.35 NRD=0 NRS=80.0214 M=1 R=4.26667
+ SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_VPWR_M1020_d N_CLK_M1020_g N_A_794_47#_M1020_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.3129 PD=0.92 PS=2.66 NRD=0 NRS=133.546 M=1 R=4.26667
+ SA=75000.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_963_47#_M1000_d N_A_794_47#_M1000_g N_VPWR_M1020_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_1237_55#_M1029_d N_A_963_47#_M1029_g N_A_244_121#_M1029_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.2247 PD=0.7 PS=1.91 NRD=0 NRS=126.632 M=1 R=2.8
+ SA=75000.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1001 A_1327_415# N_A_794_47#_M1001_g N_A_1237_55#_M1029_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75002 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_1365_29#_M1005_g A_1327_415# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1323 AS=0.0441 PD=1.05 PS=0.63 NRD=4.6886 NRS=23.443 M=1 R=2.8 SA=75001.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1040 N_A_1365_29#_M1040_d N_A_1237_55#_M1040_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.09135 AS=0.1323 PD=0.975 PS=1.05 NRD=0 NRS=159.471 M=1
+ R=2.8 SA=75002 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_SET_B_M1004_g N_A_1365_29#_M1040_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1008 AS=0.09135 PD=0.863333 PS=0.975 NRD=84.4145 NRS=44.5417 M=1
+ R=2.8 SA=75001.5 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_1781_379#_M1007_d N_A_1237_55#_M1007_g N_VPWR_M1004_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2016 PD=2.21 PS=1.72667 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.2 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1032 N_A_1998_463#_M1032_d N_A_963_47#_M1032_g N_A_1888_463#_M1032_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0952 AS=0.1999 PD=0.823333 PS=1.86 NRD=80.5139
+ NRS=56.2829 M=1 R=2.8 SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_A_1781_379#_M1030_d N_A_794_47#_M1030_g N_A_1998_463#_M1032_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.221775 AS=0.1904 PD=2.21 PS=1.64667 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1025 N_VPWR_M1025_d N_A_2214_99#_M1025_g N_A_1888_463#_M1025_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_1998_463#_M1012_d N_SET_B_M1012_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_2214_99#_M1003_d N_A_1998_463#_M1003_g N_VPWR_M1003_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1041 N_VPWR_M1041_d N_A_1998_463#_M1041_g N_A_2686_131#_M1041_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.132952 AS=0.1696 PD=1.09137 PS=1.81 NRD=13.0808 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1028 N_VPWR_M1041_d N_A_2686_131#_M1028_g N_Q_M1028_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.261748 AS=0.1764 PD=2.14863 PS=1.54 NRD=4.1567 NRS=0 M=1 R=8.4
+ SA=75000.4 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1039 N_VPWR_M1039_d N_A_2686_131#_M1039_g N_Q_M1028_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX42_noxref VNB VPB NWDIODE A=29.3551 P=35.21
c_265 VPB 0 2.80948e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfstp_2.pxi.spice"
*
.ends
*
*
