* File: sky130_fd_sc_lp__conb_0.pex.spice
* Created: Wed Sep  2 09:41:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CONB_0%HI 1 6 10 14 15 16 17 18 24 35
r40 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.445
+ $Y=1.375 $X2=0.445 $Y2=1.375
r41 18 26 4.23228 $w=5.83e-07 $l=2.07e-07 $layer=LI1_cond $X=0.572 $Y=2.035
+ $X2=0.572 $Y2=1.828
r42 18 35 10.745 $w=4.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.73 $Y=2.12
+ $X2=0.73 $Y2=2.465
r43 17 26 3.33266 $w=5.83e-07 $l=1.63e-07 $layer=LI1_cond $X=0.572 $Y=1.665
+ $X2=0.572 $Y2=1.828
r44 17 25 5.92928 $w=5.83e-07 $l=2.9e-07 $layer=LI1_cond $X=0.572 $Y=1.665
+ $X2=0.572 $Y2=1.375
r45 16 25 1.63566 $w=5.83e-07 $l=8e-08 $layer=LI1_cond $X=0.572 $Y=1.295
+ $X2=0.572 $Y2=1.375
r46 14 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.445 $Y=1.715
+ $X2=0.445 $Y2=1.375
r47 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.445 $Y=1.715
+ $X2=0.445 $Y2=1.88
r48 13 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.445 $Y=1.21
+ $X2=0.445 $Y2=1.375
r49 10 15 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.535 $Y=2.63
+ $X2=0.535 $Y2=1.88
r50 6 13 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.535 $Y=0.56
+ $X2=0.535 $Y2=1.21
r51 1 35 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=2.31 $X2=0.75 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__CONB_0%LO 1 6 8 11 13 16 18 19 20 21 22 23 30 31 32
r40 30 32 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.087 $Y=1.045
+ $X2=1.087 $Y2=0.88
r41 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.12
+ $Y=1.045 $X2=1.12 $Y2=1.045
r42 22 23 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.665
+ $X2=1.195 $Y2=2.035
r43 21 22 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.665
r44 21 31 9.00346 $w=3.18e-07 $l=2.5e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.045
r45 20 31 2.2929 $w=4.88e-07 $l=3.5e-08 $layer=LI1_cond $X=1.195 $Y=1.01
+ $X2=1.195 $Y2=1.045
r46 18 20 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.035 $Y=0.925
+ $X2=1.195 $Y2=0.925
r47 18 19 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.035 $Y=0.925
+ $X2=0.845 $Y2=0.925
r48 14 19 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.732 $Y=0.84
+ $X2=0.845 $Y2=0.925
r49 14 16 11.0122 $w=2.23e-07 $l=2.15e-07 $layer=LI1_cond $X=0.732 $Y=0.84
+ $X2=0.732 $Y2=0.625
r50 11 13 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=0.965 $Y=2.63
+ $X2=0.965 $Y2=1.55
r51 8 13 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=1.087 $Y=1.353
+ $X2=1.087 $Y2=1.55
r52 7 30 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=1.087 $Y=1.077
+ $X2=1.087 $Y2=1.045
r53 7 8 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=1.087 $Y=1.077
+ $X2=1.087 $Y2=1.353
r54 6 32 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.965 $Y=0.56
+ $X2=0.965 $Y2=0.88
r55 1 16 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.35 $X2=0.75 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LP__CONB_0%VPWR 1 2 7 9 11 13 15 17 27
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 18 23 4.1267 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r24 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 17 26 4.59592 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.237 $Y2=3.33
r26 17 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 11 26 3.00327 $w=3.1e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.237 $Y2=3.33
r31 11 13 29.3687 $w=3.08e-07 $l=7.9e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.455
r32 7 23 3.15799 $w=2.7e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.212 $Y2=3.33
r33 7 9 33.2928 $w=2.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.29 $Y=3.245 $X2=0.29
+ $Y2=2.465
r34 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.31 $X2=1.18 $Y2=2.455
r35 1 9 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=2.31 $X2=0.32 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__CONB_0%VGND 1 2 7 9 11 13 15 17 27
r22 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r23 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 18 23 4.3474 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.225
+ $Y2=0
r25 18 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.72
+ $Y2=0
r26 17 26 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.227
+ $Y2=0
r27 17 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.72
+ $Y2=0
r28 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r29 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r30 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 11 26 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.227 $Y2=0
r32 11 13 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.56
r33 7 23 3.13013 $w=2.95e-07 $l=1.17346e-07 $layer=LI1_cond $X=0.302 $Y=0.085
+ $X2=0.225 $Y2=0
r34 7 9 18.5563 $w=2.93e-07 $l=4.75e-07 $layer=LI1_cond $X=0.302 $Y=0.085
+ $X2=0.302 $Y2=0.56
r35 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.35 $X2=1.18 $Y2=0.56
r36 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.35 $X2=0.32 $Y2=0.56
.ends

