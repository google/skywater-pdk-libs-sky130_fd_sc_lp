* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__einvn_2 A TE_B VGND VNB VPB VPWR Z
M1000 a_220_367# A Z VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=6.678e+11p ps=6.1e+06u
M1001 Z A a_251_47# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=6.804e+11p ps=6.66e+06u
M1002 VGND TE_B a_28_62# VNB nshort w=420000u l=150000u
+  ad=3.465e+11p pd=3.61e+06u as=1.197e+11p ps=1.41e+06u
M1003 a_251_47# A Z VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_28_62# a_251_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_251_47# a_28_62# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR TE_B a_28_62# VPB phighvt w=640000u l=150000u
+  ad=7.382e+11p pd=6.32e+06u as=1.696e+11p ps=1.81e+06u
M1007 VPWR TE_B a_220_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_220_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_220_367# TE_B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
