* File: sky130_fd_sc_lp__nor2_8.pxi.spice
* Created: Fri Aug 28 10:53:45 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_8%A N_A_M1006_g N_A_M1000_g N_A_M1008_g N_A_M1004_g
+ N_A_M1011_g N_A_M1005_g N_A_M1017_g N_A_M1010_g N_A_M1020_g N_A_M1012_g
+ N_A_M1025_g N_A_M1019_g N_A_M1028_g N_A_M1022_g N_A_M1031_g N_A_M1029_g A A A
+ A N_A_c_123_n PM_SKY130_FD_SC_LP__NOR2_8%A
x_PM_SKY130_FD_SC_LP__NOR2_8%B N_B_M1003_g N_B_M1001_g N_B_M1013_g N_B_M1002_g
+ N_B_M1016_g N_B_M1007_g N_B_M1018_g N_B_M1009_g N_B_M1023_g N_B_M1014_g
+ N_B_M1026_g N_B_M1015_g N_B_M1027_g N_B_M1021_g N_B_M1030_g N_B_M1024_g B B B
+ B N_B_c_265_n PM_SKY130_FD_SC_LP__NOR2_8%B
x_PM_SKY130_FD_SC_LP__NOR2_8%A_47_367# N_A_47_367#_M1000_s N_A_47_367#_M1004_s
+ N_A_47_367#_M1010_s N_A_47_367#_M1019_s N_A_47_367#_M1029_s
+ N_A_47_367#_M1002_d N_A_47_367#_M1009_d N_A_47_367#_M1015_d
+ N_A_47_367#_M1024_d N_A_47_367#_c_407_n N_A_47_367#_c_408_n
+ N_A_47_367#_c_413_n N_A_47_367#_c_457_p N_A_47_367#_c_417_n
+ N_A_47_367#_c_454_p N_A_47_367#_c_421_n N_A_47_367#_c_455_p
+ N_A_47_367#_c_409_n N_A_47_367#_c_458_p N_A_47_367#_c_437_n
+ N_A_47_367#_c_439_n N_A_47_367#_c_440_n N_A_47_367#_c_495_p
+ N_A_47_367#_c_442_n N_A_47_367#_c_497_p N_A_47_367#_c_410_n
+ N_A_47_367#_c_411_n N_A_47_367#_c_428_n N_A_47_367#_c_430_n
+ N_A_47_367#_c_412_n N_A_47_367#_c_463_p N_A_47_367#_c_464_p
+ N_A_47_367#_c_465_p PM_SKY130_FD_SC_LP__NOR2_8%A_47_367#
x_PM_SKY130_FD_SC_LP__NOR2_8%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_M1012_d
+ N_VPWR_M1022_d N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n
+ N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n VPWR
+ N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_510_n N_VPWR_c_523_n
+ N_VPWR_c_524_n PM_SKY130_FD_SC_LP__NOR2_8%VPWR
x_PM_SKY130_FD_SC_LP__NOR2_8%Y N_Y_M1006_s N_Y_M1011_s N_Y_M1020_s N_Y_M1028_s
+ N_Y_M1003_d N_Y_M1016_d N_Y_M1023_d N_Y_M1027_d N_Y_M1001_s N_Y_M1007_s
+ N_Y_M1014_s N_Y_M1021_s N_Y_c_617_n N_Y_c_618_n N_Y_c_619_n N_Y_c_620_n
+ N_Y_c_621_n N_Y_c_622_n N_Y_c_623_n N_Y_c_624_n N_Y_c_625_n N_Y_c_626_n
+ N_Y_c_691_n N_Y_c_627_n N_Y_c_628_n N_Y_c_701_n N_Y_c_629_n N_Y_c_630_n
+ N_Y_c_639_n N_Y_c_631_n N_Y_c_632_n N_Y_c_633_n N_Y_c_634_n N_Y_c_670_n
+ N_Y_c_715_n N_Y_c_635_n N_Y_c_723_n N_Y_c_636_n Y Y Y N_Y_c_637_n N_Y_c_638_n
+ Y N_Y_c_737_n PM_SKY130_FD_SC_LP__NOR2_8%Y
x_PM_SKY130_FD_SC_LP__NOR2_8%VGND N_VGND_M1006_d N_VGND_M1008_d N_VGND_M1017_d
+ N_VGND_M1025_d N_VGND_M1031_d N_VGND_M1013_s N_VGND_M1018_s N_VGND_M1026_s
+ N_VGND_M1030_s N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n
+ N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n
+ N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n N_VGND_c_827_n
+ N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n
+ N_VGND_c_833_n VGND N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n
+ N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ PM_SKY130_FD_SC_LP__NOR2_8%VGND
cc_1 VNB N_A_M1006_g 0.0268227f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.745
cc_2 VNB N_A_M1008_g 0.019179f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.745
cc_3 VNB N_A_M1011_g 0.0191786f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.745
cc_4 VNB N_A_M1017_g 0.0191568f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=0.745
cc_5 VNB N_A_M1020_g 0.0191273f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=0.745
cc_6 VNB N_A_M1025_g 0.0187156f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.745
cc_7 VNB N_A_M1028_g 0.0187156f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=0.745
cc_8 VNB N_A_M1031_g 0.018811f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=0.745
cc_9 VNB A 0.00973387f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_10 VNB N_A_c_123_n 0.137876f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.51
cc_11 VNB N_B_M1003_g 0.0188243f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.745
cc_12 VNB N_B_M1013_g 0.0196943f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.745
cc_13 VNB N_B_M1016_g 0.0196942f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.745
cc_14 VNB N_B_M1018_g 0.0187162f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=0.745
cc_15 VNB N_B_M1023_g 0.0190688f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=0.745
cc_16 VNB N_B_M1026_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.745
cc_17 VNB N_B_M1027_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=0.745
cc_18 VNB N_B_M1030_g 0.0230591f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=0.745
cc_19 VNB B 0.00277815f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_20 VNB N_B_c_265_n 0.135562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_510_n 0.322901f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.675
cc_22 VNB N_Y_c_617_n 0.00181291f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=2.465
cc_23 VNB N_Y_c_618_n 0.00304705f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.345
cc_24 VNB N_Y_c_619_n 0.00249829f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.745
cc_25 VNB N_Y_c_620_n 0.00168668f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.675
cc_26 VNB N_Y_c_621_n 0.0041544f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=2.465
cc_27 VNB N_Y_c_622_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=0.745
cc_28 VNB N_Y_c_623_n 0.00257839f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=2.465
cc_29 VNB N_Y_c_624_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=2.465
cc_30 VNB N_Y_c_625_n 0.00284925f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_31 VNB N_Y_c_626_n 0.0044608f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_32 VNB N_Y_c_627_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.51
cc_33 VNB N_Y_c_628_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.51
cc_34 VNB N_Y_c_629_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=1.51
cc_35 VNB N_Y_c_630_n 0.0219142f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.51
cc_36 VNB N_Y_c_631_n 0.019905f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.51
cc_37 VNB N_Y_c_632_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=1.51
cc_38 VNB N_Y_c_633_n 0.00186118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_634_n 0.00579579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_635_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_636_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_637_n 0.0081949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_638_n 0.00251142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_814_n 0.0138616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_815_n 0.0531992f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=2.465
cc_46 VNB N_VGND_c_816_n 0.00178862f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=0.745
cc_47 VNB N_VGND_c_817_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=2.465
cc_48 VNB N_VGND_c_818_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.745
cc_49 VNB N_VGND_c_819_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=2.465
cc_50 VNB N_VGND_c_820_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_821_n 0.00406919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_822_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_823_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_824_n 0.0302167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_825_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_56 VNB N_VGND_c_826_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_57 VNB N_VGND_c_827_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_828_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_829_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_830_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.51
cc_61 VNB N_VGND_c_831_n 0.0108943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_832_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.51
cc_63 VNB N_VGND_c_833_n 0.00581671f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.51
cc_64 VNB N_VGND_c_834_n 0.0146725f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.51
cc_65 VNB N_VGND_c_835_n 0.0143206f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=1.51
cc_66 VNB N_VGND_c_836_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_837_n 0.417829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_838_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_839_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_840_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_841_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_A_M1000_g 0.0238016f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_73 VPB N_A_M1004_g 0.0177715f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.465
cc_74 VPB N_A_M1005_g 0.0177715f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=2.465
cc_75 VPB N_A_M1010_g 0.0177715f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=2.465
cc_76 VPB N_A_M1012_g 0.018136f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.465
cc_77 VPB N_A_M1019_g 0.0184815f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.465
cc_78 VPB N_A_M1022_g 0.0173862f $X=-0.19 $Y=1.655 $X2=3.155 $Y2=2.465
cc_79 VPB N_A_M1029_g 0.0174893f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=2.465
cc_80 VPB A 0.0150158f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_81 VPB N_A_c_123_n 0.0262743f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.51
cc_82 VPB N_B_M1001_g 0.0183435f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_83 VPB N_B_M1002_g 0.0173762f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.465
cc_84 VPB N_B_M1007_g 0.0173762f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=2.465
cc_85 VPB N_B_M1009_g 0.018045f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=2.465
cc_86 VPB N_B_M1014_g 0.0181319f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.465
cc_87 VPB N_B_M1015_g 0.0181378f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.465
cc_88 VPB N_B_M1021_g 0.0181378f $X=-0.19 $Y=1.655 $X2=3.155 $Y2=2.465
cc_89 VPB N_B_M1024_g 0.0225369f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=2.465
cc_90 VPB B 0.0116335f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_91 VPB N_B_c_265_n 0.0276913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_47_367#_c_407_n 0.00927443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_47_367#_c_408_n 0.0371579f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=2.465
cc_94 VPB N_A_47_367#_c_409_n 0.00654072f $X=-0.19 $Y=1.655 $X2=3.155 $Y2=0.745
cc_95 VPB N_A_47_367#_c_410_n 0.00788844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_47_367#_c_411_n 0.0242286f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.51
cc_97 VPB N_A_47_367#_c_412_n 0.00331358f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=1.51
cc_98 VPB N_VPWR_c_511_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.465
cc_99 VPB N_VPWR_c_512_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.435 $Y2=0.745
cc_100 VPB N_VPWR_c_513_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.435 $Y2=2.465
cc_101 VPB N_VPWR_c_514_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.865 $Y2=0.745
cc_102 VPB N_VPWR_c_515_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_516_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.345
cc_104 VPB N_VPWR_c_517_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=0.745
cc_105 VPB N_VPWR_c_518_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_519_n 0.018464f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.465
cc_107 VPB N_VPWR_c_520_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_521_n 0.0971986f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_510_n 0.0565986f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.675
cc_110 VPB N_VPWR_c_523_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_524_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_112 VPB N_Y_c_639_n 0.0171388f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=1.51
cc_113 VPB N_Y_c_631_n 0.0133295f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=1.51
cc_114 N_A_M1031_g N_B_M1003_g 0.0181144f $X=3.585 $Y=0.745 $X2=0 $Y2=0
cc_115 N_A_M1029_g N_B_M1001_g 0.0181144f $X=3.585 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_c_123_n N_B_c_265_n 0.0181144f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_117 N_A_M1000_g N_A_47_367#_c_413_n 0.0122595f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_M1004_g N_A_47_367#_c_413_n 0.0122595f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_119 A N_A_47_367#_c_413_n 0.0411927f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_120 N_A_c_123_n N_A_47_367#_c_413_n 5.51615e-19 $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_121 N_A_M1005_g N_A_47_367#_c_417_n 0.0122595f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_M1010_g N_A_47_367#_c_417_n 0.0122595f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_123 A N_A_47_367#_c_417_n 0.043087f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A_c_123_n N_A_47_367#_c_417_n 5.51615e-19 $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A_M1012_g N_A_47_367#_c_421_n 0.0160306f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_M1019_g N_A_47_367#_c_421_n 0.0137237f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_127 A N_A_47_367#_c_421_n 0.00365635f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A_c_123_n N_A_47_367#_c_421_n 0.002265f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A_M1022_g N_A_47_367#_c_409_n 0.0147238f $X=3.155 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_M1029_g N_A_47_367#_c_409_n 0.0153703f $X=3.585 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_c_123_n N_A_47_367#_c_409_n 0.0027593f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_132 A N_A_47_367#_c_428_n 0.0154822f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A_c_123_n N_A_47_367#_c_428_n 6.23431e-19 $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_134 A N_A_47_367#_c_430_n 0.0154822f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A_c_123_n N_A_47_367#_c_430_n 6.23431e-19 $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_136 N_A_M1019_g N_A_47_367#_c_412_n 0.00257213f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_M1022_g N_A_47_367#_c_412_n 2.94561e-19 $X=3.155 $Y=2.465 $X2=0 $Y2=0
cc_138 A N_A_47_367#_c_412_n 0.00216068f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A_c_123_n N_A_47_367#_c_412_n 0.00288231f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_140 N_A_M1000_g N_VPWR_c_511_n 0.0165759f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_M1004_g N_VPWR_c_511_n 0.014697f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_M1005_g N_VPWR_c_511_n 6.74833e-19 $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_M1004_g N_VPWR_c_512_n 6.74833e-19 $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1005_g N_VPWR_c_512_n 0.014697f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1010_g N_VPWR_c_512_n 0.014697f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1012_g N_VPWR_c_512_n 6.74833e-19 $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1010_g N_VPWR_c_513_n 6.74833e-19 $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_M1012_g N_VPWR_c_513_n 0.014697f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_M1019_g N_VPWR_c_513_n 0.014697f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_M1022_g N_VPWR_c_513_n 6.74833e-19 $X=3.155 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_M1019_g N_VPWR_c_514_n 7.2321e-19 $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_M1022_g N_VPWR_c_514_n 0.0142189f $X=3.155 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_M1029_g N_VPWR_c_514_n 0.0153918f $X=3.585 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_M1010_g N_VPWR_c_515_n 0.00486043f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_M1012_g N_VPWR_c_515_n 0.00486043f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_M1019_g N_VPWR_c_517_n 0.00486043f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_M1022_g N_VPWR_c_517_n 0.00486043f $X=3.155 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_M1000_g N_VPWR_c_519_n 0.00486043f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_M1004_g N_VPWR_c_520_n 0.00486043f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A_M1005_g N_VPWR_c_520_n 0.00486043f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A_M1029_g N_VPWR_c_521_n 0.00486043f $X=3.585 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_M1000_g N_VPWR_c_510_n 0.00926166f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_M1004_g N_VPWR_c_510_n 0.00824727f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A_M1005_g N_VPWR_c_510_n 0.00824727f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_M1010_g N_VPWR_c_510_n 0.00824727f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A_M1012_g N_VPWR_c_510_n 0.00824727f $X=2.295 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_M1019_g N_VPWR_c_510_n 0.00824727f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_M1022_g N_VPWR_c_510_n 0.00824727f $X=3.155 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_M1029_g N_VPWR_c_510_n 0.0082726f $X=3.585 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_M1006_g N_Y_c_617_n 7.36945e-19 $X=0.575 $Y=0.745 $X2=0 $Y2=0
cc_171 N_A_M1008_g N_Y_c_617_n 7.14179e-19 $X=1.005 $Y=0.745 $X2=0 $Y2=0
cc_172 N_A_M1008_g N_Y_c_618_n 0.0130254f $X=1.005 $Y=0.745 $X2=0 $Y2=0
cc_173 N_A_M1011_g N_Y_c_618_n 0.0131657f $X=1.435 $Y=0.745 $X2=0 $Y2=0
cc_174 A N_Y_c_618_n 0.0494427f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A_c_123_n N_Y_c_618_n 0.00243542f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A_M1006_g N_Y_c_619_n 0.00212438f $X=0.575 $Y=0.745 $X2=0 $Y2=0
cc_177 A N_Y_c_619_n 0.0173765f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A_c_123_n N_Y_c_619_n 0.00253619f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A_M1011_g N_Y_c_620_n 7.13716e-19 $X=1.435 $Y=0.745 $X2=0 $Y2=0
cc_180 N_A_M1017_g N_Y_c_620_n 7.13716e-19 $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_181 N_A_M1017_g N_Y_c_621_n 0.0131751f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_182 N_A_M1020_g N_Y_c_621_n 0.0168985f $X=2.295 $Y=0.745 $X2=0 $Y2=0
cc_183 A N_Y_c_621_n 0.0370993f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A_c_123_n N_Y_c_621_n 0.00243542f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A_M1020_g N_Y_c_622_n 8.28776e-19 $X=2.295 $Y=0.745 $X2=0 $Y2=0
cc_186 N_A_M1025_g N_Y_c_622_n 8.28776e-19 $X=2.725 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A_M1028_g N_Y_c_623_n 0.0014183f $X=3.155 $Y=0.745 $X2=0 $Y2=0
cc_188 N_A_M1031_g N_Y_c_623_n 0.00141873f $X=3.585 $Y=0.745 $X2=0 $Y2=0
cc_189 N_A_c_123_n N_Y_c_626_n 0.00121348f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_190 A N_Y_c_632_n 0.0161048f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A_c_123_n N_Y_c_632_n 0.00253619f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_192 N_A_M1020_g N_Y_c_633_n 0.00316014f $X=2.295 $Y=0.745 $X2=0 $Y2=0
cc_193 N_A_M1025_g N_Y_c_633_n 7.45492e-19 $X=2.725 $Y=0.745 $X2=0 $Y2=0
cc_194 A N_Y_c_633_n 0.00557615f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A_c_123_n N_Y_c_633_n 0.0132563f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A_M1025_g N_Y_c_634_n 0.0109978f $X=2.725 $Y=0.745 $X2=0 $Y2=0
cc_197 N_A_M1028_g N_Y_c_634_n 0.0112545f $X=3.155 $Y=0.745 $X2=0 $Y2=0
cc_198 N_A_c_123_n N_Y_c_634_n 0.0223513f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A_c_123_n N_Y_c_670_n 0.00755804f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A_M1031_g N_Y_c_637_n 0.0112451f $X=3.585 $Y=0.745 $X2=0 $Y2=0
cc_201 N_A_c_123_n N_Y_c_637_n 0.00727013f $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_202 N_A_M1006_g N_VGND_c_815_n 0.0162817f $X=0.575 $Y=0.745 $X2=0 $Y2=0
cc_203 N_A_M1008_g N_VGND_c_815_n 6.05476e-19 $X=1.005 $Y=0.745 $X2=0 $Y2=0
cc_204 A N_VGND_c_815_n 5.66516e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A_M1006_g N_VGND_c_816_n 5.39497e-19 $X=0.575 $Y=0.745 $X2=0 $Y2=0
cc_206 N_A_M1008_g N_VGND_c_816_n 0.0102233f $X=1.005 $Y=0.745 $X2=0 $Y2=0
cc_207 N_A_M1011_g N_VGND_c_816_n 0.0101946f $X=1.435 $Y=0.745 $X2=0 $Y2=0
cc_208 N_A_M1017_g N_VGND_c_816_n 5.36081e-19 $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_209 N_A_M1011_g N_VGND_c_817_n 5.36081e-19 $X=1.435 $Y=0.745 $X2=0 $Y2=0
cc_210 N_A_M1017_g N_VGND_c_817_n 0.0101946f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_211 N_A_M1020_g N_VGND_c_817_n 0.0101212f $X=2.295 $Y=0.745 $X2=0 $Y2=0
cc_212 N_A_M1025_g N_VGND_c_817_n 5.09471e-19 $X=2.725 $Y=0.745 $X2=0 $Y2=0
cc_213 N_A_M1020_g N_VGND_c_818_n 5.47664e-19 $X=2.295 $Y=0.745 $X2=0 $Y2=0
cc_214 N_A_M1025_g N_VGND_c_818_n 0.012629f $X=2.725 $Y=0.745 $X2=0 $Y2=0
cc_215 N_A_M1028_g N_VGND_c_818_n 0.012629f $X=3.155 $Y=0.745 $X2=0 $Y2=0
cc_216 N_A_M1031_g N_VGND_c_818_n 5.47664e-19 $X=3.585 $Y=0.745 $X2=0 $Y2=0
cc_217 N_A_c_123_n N_VGND_c_818_n 5.70981e-19 $X=3.585 $Y=1.51 $X2=0 $Y2=0
cc_218 N_A_M1028_g N_VGND_c_819_n 5.47664e-19 $X=3.155 $Y=0.745 $X2=0 $Y2=0
cc_219 N_A_M1031_g N_VGND_c_819_n 0.0125669f $X=3.585 $Y=0.745 $X2=0 $Y2=0
cc_220 N_A_M1020_g N_VGND_c_825_n 0.00414769f $X=2.295 $Y=0.745 $X2=0 $Y2=0
cc_221 N_A_M1025_g N_VGND_c_825_n 0.00414769f $X=2.725 $Y=0.745 $X2=0 $Y2=0
cc_222 N_A_M1028_g N_VGND_c_827_n 0.00414769f $X=3.155 $Y=0.745 $X2=0 $Y2=0
cc_223 N_A_M1031_g N_VGND_c_827_n 0.00414769f $X=3.585 $Y=0.745 $X2=0 $Y2=0
cc_224 N_A_M1006_g N_VGND_c_834_n 0.00464723f $X=0.575 $Y=0.745 $X2=0 $Y2=0
cc_225 N_A_M1008_g N_VGND_c_834_n 0.00414769f $X=1.005 $Y=0.745 $X2=0 $Y2=0
cc_226 N_A_M1011_g N_VGND_c_835_n 0.00414769f $X=1.435 $Y=0.745 $X2=0 $Y2=0
cc_227 N_A_M1017_g N_VGND_c_835_n 0.00414769f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_228 N_A_M1006_g N_VGND_c_837_n 0.00880442f $X=0.575 $Y=0.745 $X2=0 $Y2=0
cc_229 N_A_M1008_g N_VGND_c_837_n 0.00787505f $X=1.005 $Y=0.745 $X2=0 $Y2=0
cc_230 N_A_M1011_g N_VGND_c_837_n 0.00787505f $X=1.435 $Y=0.745 $X2=0 $Y2=0
cc_231 N_A_M1017_g N_VGND_c_837_n 0.00787505f $X=1.865 $Y=0.745 $X2=0 $Y2=0
cc_232 N_A_M1020_g N_VGND_c_837_n 0.00787505f $X=2.295 $Y=0.745 $X2=0 $Y2=0
cc_233 N_A_M1025_g N_VGND_c_837_n 0.00787505f $X=2.725 $Y=0.745 $X2=0 $Y2=0
cc_234 N_A_M1028_g N_VGND_c_837_n 0.00787505f $X=3.155 $Y=0.745 $X2=0 $Y2=0
cc_235 N_A_M1031_g N_VGND_c_837_n 0.00787505f $X=3.585 $Y=0.745 $X2=0 $Y2=0
cc_236 N_B_M1001_g N_A_47_367#_c_409_n 0.00110679f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B_M1001_g N_A_47_367#_c_437_n 0.0114588f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B_M1002_g N_A_47_367#_c_437_n 0.0114565f $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B_c_265_n N_A_47_367#_c_439_n 3.40512e-19 $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_240 N_B_M1007_g N_A_47_367#_c_440_n 0.0115031f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B_M1009_g N_A_47_367#_c_440_n 0.0115031f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B_M1014_g N_A_47_367#_c_442_n 0.0118004f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B_M1015_g N_A_47_367#_c_442_n 0.0117979f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B_M1021_g N_A_47_367#_c_410_n 0.0118004f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B_M1024_g N_A_47_367#_c_410_n 0.0118004f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B_M1001_g N_VPWR_c_514_n 0.00109252f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B_M1001_g N_VPWR_c_521_n 0.00357877f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B_M1002_g N_VPWR_c_521_n 0.00357877f $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_249 N_B_M1007_g N_VPWR_c_521_n 0.00357877f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_250 N_B_M1009_g N_VPWR_c_521_n 0.00357877f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B_M1014_g N_VPWR_c_521_n 0.00357877f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_252 N_B_M1015_g N_VPWR_c_521_n 0.00357877f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_253 N_B_M1021_g N_VPWR_c_521_n 0.00357877f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_254 N_B_M1024_g N_VPWR_c_521_n 0.00357877f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B_M1001_g N_VPWR_c_510_n 0.00537654f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B_M1002_g N_VPWR_c_510_n 0.0053512f $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_257 N_B_M1007_g N_VPWR_c_510_n 0.0053512f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_258 N_B_M1009_g N_VPWR_c_510_n 0.0053512f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B_M1014_g N_VPWR_c_510_n 0.0053512f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B_M1015_g N_VPWR_c_510_n 0.0053512f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_261 N_B_M1021_g N_VPWR_c_510_n 0.0053512f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_262 N_B_M1024_g N_VPWR_c_510_n 0.00641531f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_263 N_B_M1016_g N_Y_c_624_n 8.28776e-19 $X=4.875 $Y=0.745 $X2=0 $Y2=0
cc_264 N_B_M1018_g N_Y_c_624_n 8.28776e-19 $X=5.305 $Y=0.745 $X2=0 $Y2=0
cc_265 N_B_M1018_g N_Y_c_625_n 0.0131128f $X=5.305 $Y=0.745 $X2=0 $Y2=0
cc_266 N_B_M1023_g N_Y_c_625_n 0.013286f $X=5.735 $Y=0.745 $X2=0 $Y2=0
cc_267 B N_Y_c_625_n 0.0324334f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_268 N_B_c_265_n N_Y_c_625_n 0.00246472f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_269 N_B_M1003_g N_Y_c_626_n 0.00285524f $X=4.015 $Y=0.745 $X2=0 $Y2=0
cc_270 N_B_M1001_g N_Y_c_626_n 0.0063144f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_271 N_B_M1013_g N_Y_c_626_n 0.00226795f $X=4.445 $Y=0.745 $X2=0 $Y2=0
cc_272 N_B_M1002_g N_Y_c_626_n 0.0166011f $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_273 N_B_M1016_g N_Y_c_626_n 0.00256544f $X=4.875 $Y=0.745 $X2=0 $Y2=0
cc_274 N_B_M1007_g N_Y_c_626_n 0.0166011f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_275 N_B_M1018_g N_Y_c_626_n 0.00413878f $X=5.305 $Y=0.745 $X2=0 $Y2=0
cc_276 N_B_M1009_g N_Y_c_626_n 0.00651444f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_277 N_B_M1023_g N_Y_c_626_n 4.28404e-19 $X=5.735 $Y=0.745 $X2=0 $Y2=0
cc_278 N_B_M1014_g N_Y_c_626_n 8.63016e-19 $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_279 B N_Y_c_626_n 0.0276322f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_280 N_B_c_265_n N_Y_c_626_n 0.0760078f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_281 N_B_M1009_g N_Y_c_691_n 0.0129633f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_282 N_B_M1014_g N_Y_c_691_n 0.01115f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_283 B N_Y_c_691_n 0.0250873f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_284 N_B_c_265_n N_Y_c_691_n 5.78305e-19 $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_285 N_B_M1023_g N_Y_c_627_n 8.28776e-19 $X=5.735 $Y=0.745 $X2=0 $Y2=0
cc_286 N_B_M1026_g N_Y_c_627_n 8.28776e-19 $X=6.165 $Y=0.745 $X2=0 $Y2=0
cc_287 N_B_M1026_g N_Y_c_628_n 0.0133326f $X=6.165 $Y=0.745 $X2=0 $Y2=0
cc_288 N_B_M1027_g N_Y_c_628_n 0.0133326f $X=6.595 $Y=0.745 $X2=0 $Y2=0
cc_289 B N_Y_c_628_n 0.0491013f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_290 N_B_c_265_n N_Y_c_628_n 0.00246472f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_291 N_B_M1015_g N_Y_c_701_n 0.01115f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_292 N_B_M1021_g N_Y_c_701_n 0.01115f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_293 B N_Y_c_701_n 0.0354228f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_294 N_B_c_265_n N_Y_c_701_n 5.78305e-19 $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_295 N_B_M1027_g N_Y_c_629_n 8.28776e-19 $X=6.595 $Y=0.745 $X2=0 $Y2=0
cc_296 N_B_M1030_g N_Y_c_629_n 8.28776e-19 $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_297 N_B_M1030_g N_Y_c_630_n 0.0151021f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_298 B N_Y_c_630_n 0.0140399f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_299 N_B_M1024_g N_Y_c_639_n 0.0129195f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_300 B N_Y_c_639_n 0.00888173f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_301 N_B_M1030_g N_Y_c_631_n 0.00543294f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_302 N_B_M1024_g N_Y_c_631_n 0.00494811f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_303 B N_Y_c_631_n 0.0158301f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_304 N_B_c_265_n N_Y_c_631_n 0.00196917f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_305 N_B_M1009_g N_Y_c_715_n 5.66402e-19 $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_306 N_B_M1014_g N_Y_c_715_n 0.0112362f $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_307 N_B_M1015_g N_Y_c_715_n 0.0112362f $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_308 N_B_M1021_g N_Y_c_715_n 5.66402e-19 $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_309 B N_Y_c_715_n 0.0230324f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_310 N_B_c_265_n N_Y_c_715_n 6.52992e-19 $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_311 B N_Y_c_635_n 0.0160075f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_312 N_B_c_265_n N_Y_c_635_n 0.00256759f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_313 N_B_M1015_g N_Y_c_723_n 5.66402e-19 $X=6.165 $Y=2.465 $X2=0 $Y2=0
cc_314 N_B_M1021_g N_Y_c_723_n 0.0112362f $X=6.595 $Y=2.465 $X2=0 $Y2=0
cc_315 N_B_M1024_g N_Y_c_723_n 0.0158667f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_316 B N_Y_c_723_n 0.0230324f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_317 N_B_c_265_n N_Y_c_723_n 6.52992e-19 $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_318 B N_Y_c_636_n 0.0160075f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_319 N_B_c_265_n N_Y_c_636_n 0.00256759f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_320 N_B_M1001_g Y 0.0101747f $X=4.015 $Y=2.465 $X2=0 $Y2=0
cc_321 N_B_M1002_g Y 0.0114475f $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_322 N_B_M1007_g Y 5.69231e-19 $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_323 N_B_M1003_g N_Y_c_637_n 0.00811512f $X=4.015 $Y=0.745 $X2=0 $Y2=0
cc_324 N_B_c_265_n N_Y_c_637_n 0.00908345f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_325 N_B_M1003_g N_Y_c_638_n 0.00141873f $X=4.015 $Y=0.745 $X2=0 $Y2=0
cc_326 N_B_M1013_g N_Y_c_638_n 0.00126708f $X=4.445 $Y=0.745 $X2=0 $Y2=0
cc_327 N_B_M1002_g N_Y_c_737_n 5.69231e-19 $X=4.445 $Y=2.465 $X2=0 $Y2=0
cc_328 N_B_M1007_g N_Y_c_737_n 0.0114475f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_329 N_B_M1009_g N_Y_c_737_n 0.0114475f $X=5.305 $Y=2.465 $X2=0 $Y2=0
cc_330 N_B_M1014_g N_Y_c_737_n 5.69231e-19 $X=5.735 $Y=2.465 $X2=0 $Y2=0
cc_331 N_B_M1003_g N_VGND_c_819_n 0.0125669f $X=4.015 $Y=0.745 $X2=0 $Y2=0
cc_332 N_B_M1013_g N_VGND_c_819_n 5.47664e-19 $X=4.445 $Y=0.745 $X2=0 $Y2=0
cc_333 N_B_M1003_g N_VGND_c_820_n 0.00414769f $X=4.015 $Y=0.745 $X2=0 $Y2=0
cc_334 N_B_M1013_g N_VGND_c_820_n 0.00414769f $X=4.445 $Y=0.745 $X2=0 $Y2=0
cc_335 N_B_M1003_g N_VGND_c_821_n 5.901e-19 $X=4.015 $Y=0.745 $X2=0 $Y2=0
cc_336 N_B_M1013_g N_VGND_c_821_n 0.0152898f $X=4.445 $Y=0.745 $X2=0 $Y2=0
cc_337 N_B_M1016_g N_VGND_c_821_n 0.0152795f $X=4.875 $Y=0.745 $X2=0 $Y2=0
cc_338 N_B_M1018_g N_VGND_c_821_n 6.01289e-19 $X=5.305 $Y=0.745 $X2=0 $Y2=0
cc_339 N_B_c_265_n N_VGND_c_821_n 0.00237027f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_340 N_B_M1016_g N_VGND_c_822_n 5.123e-19 $X=4.875 $Y=0.745 $X2=0 $Y2=0
cc_341 N_B_M1018_g N_VGND_c_822_n 0.0102222f $X=5.305 $Y=0.745 $X2=0 $Y2=0
cc_342 N_B_M1023_g N_VGND_c_822_n 0.0102222f $X=5.735 $Y=0.745 $X2=0 $Y2=0
cc_343 N_B_M1026_g N_VGND_c_822_n 5.123e-19 $X=6.165 $Y=0.745 $X2=0 $Y2=0
cc_344 N_B_M1023_g N_VGND_c_823_n 5.123e-19 $X=5.735 $Y=0.745 $X2=0 $Y2=0
cc_345 N_B_M1026_g N_VGND_c_823_n 0.0102222f $X=6.165 $Y=0.745 $X2=0 $Y2=0
cc_346 N_B_M1027_g N_VGND_c_823_n 0.0102222f $X=6.595 $Y=0.745 $X2=0 $Y2=0
cc_347 N_B_M1030_g N_VGND_c_823_n 5.123e-19 $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_348 N_B_M1027_g N_VGND_c_824_n 5.123e-19 $X=6.595 $Y=0.745 $X2=0 $Y2=0
cc_349 N_B_M1030_g N_VGND_c_824_n 0.0112857f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_350 N_B_M1023_g N_VGND_c_829_n 0.00414769f $X=5.735 $Y=0.745 $X2=0 $Y2=0
cc_351 N_B_M1026_g N_VGND_c_829_n 0.00414769f $X=6.165 $Y=0.745 $X2=0 $Y2=0
cc_352 N_B_M1027_g N_VGND_c_832_n 0.00414769f $X=6.595 $Y=0.745 $X2=0 $Y2=0
cc_353 N_B_M1030_g N_VGND_c_832_n 0.00414769f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_354 N_B_M1016_g N_VGND_c_836_n 0.00414769f $X=4.875 $Y=0.745 $X2=0 $Y2=0
cc_355 N_B_M1018_g N_VGND_c_836_n 0.00414769f $X=5.305 $Y=0.745 $X2=0 $Y2=0
cc_356 N_B_M1003_g N_VGND_c_837_n 0.00787505f $X=4.015 $Y=0.745 $X2=0 $Y2=0
cc_357 N_B_M1013_g N_VGND_c_837_n 0.00787505f $X=4.445 $Y=0.745 $X2=0 $Y2=0
cc_358 N_B_M1016_g N_VGND_c_837_n 0.00787505f $X=4.875 $Y=0.745 $X2=0 $Y2=0
cc_359 N_B_M1018_g N_VGND_c_837_n 0.00787505f $X=5.305 $Y=0.745 $X2=0 $Y2=0
cc_360 N_B_M1023_g N_VGND_c_837_n 0.00787505f $X=5.735 $Y=0.745 $X2=0 $Y2=0
cc_361 N_B_M1026_g N_VGND_c_837_n 0.00787505f $X=6.165 $Y=0.745 $X2=0 $Y2=0
cc_362 N_B_M1027_g N_VGND_c_837_n 0.00787505f $X=6.595 $Y=0.745 $X2=0 $Y2=0
cc_363 N_B_M1030_g N_VGND_c_837_n 0.00787505f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_364 N_A_47_367#_c_413_n N_VPWR_M1000_d 0.00333523f $X=1.125 $Y=2.025
+ $X2=-0.19 $Y2=1.655
cc_365 N_A_47_367#_c_417_n N_VPWR_M1005_d 0.00333523f $X=1.985 $Y=2.025 $X2=0
+ $Y2=0
cc_366 N_A_47_367#_c_421_n N_VPWR_M1012_d 0.00421083f $X=2.83 $Y=2.025 $X2=0
+ $Y2=0
cc_367 N_A_47_367#_c_409_n N_VPWR_M1022_d 0.00177993f $X=3.705 $Y=1.812 $X2=0
+ $Y2=0
cc_368 N_A_47_367#_c_413_n N_VPWR_c_511_n 0.0170777f $X=1.125 $Y=2.025 $X2=0
+ $Y2=0
cc_369 N_A_47_367#_c_417_n N_VPWR_c_512_n 0.0170777f $X=1.985 $Y=2.025 $X2=0
+ $Y2=0
cc_370 N_A_47_367#_c_421_n N_VPWR_c_513_n 0.0170777f $X=2.83 $Y=2.025 $X2=0
+ $Y2=0
cc_371 N_A_47_367#_c_409_n N_VPWR_c_514_n 0.0174094f $X=3.705 $Y=1.812 $X2=0
+ $Y2=0
cc_372 N_A_47_367#_c_454_p N_VPWR_c_515_n 0.0124525f $X=2.08 $Y=2.91 $X2=0 $Y2=0
cc_373 N_A_47_367#_c_455_p N_VPWR_c_517_n 0.0124525f $X=2.94 $Y=2.45 $X2=0 $Y2=0
cc_374 N_A_47_367#_c_408_n N_VPWR_c_519_n 0.018528f $X=0.36 $Y=2.91 $X2=0 $Y2=0
cc_375 N_A_47_367#_c_457_p N_VPWR_c_520_n 0.0124525f $X=1.22 $Y=2.91 $X2=0 $Y2=0
cc_376 N_A_47_367#_c_458_p N_VPWR_c_521_n 0.0125234f $X=3.8 $Y=2.905 $X2=0 $Y2=0
cc_377 N_A_47_367#_c_437_n N_VPWR_c_521_n 0.0361172f $X=4.565 $Y=2.99 $X2=0
+ $Y2=0
cc_378 N_A_47_367#_c_440_n N_VPWR_c_521_n 0.0361172f $X=5.425 $Y=2.99 $X2=0
+ $Y2=0
cc_379 N_A_47_367#_c_442_n N_VPWR_c_521_n 0.0362264f $X=6.285 $Y=2.985 $X2=0
+ $Y2=0
cc_380 N_A_47_367#_c_410_n N_VPWR_c_521_n 0.0541447f $X=7.145 $Y=2.985 $X2=0
+ $Y2=0
cc_381 N_A_47_367#_c_463_p N_VPWR_c_521_n 0.0125234f $X=4.66 $Y=2.99 $X2=0 $Y2=0
cc_382 N_A_47_367#_c_464_p N_VPWR_c_521_n 0.0125234f $X=5.52 $Y=2.985 $X2=0
+ $Y2=0
cc_383 N_A_47_367#_c_465_p N_VPWR_c_521_n 0.0125234f $X=6.38 $Y=2.985 $X2=0
+ $Y2=0
cc_384 N_A_47_367#_M1000_s N_VPWR_c_510_n 0.00371702f $X=0.235 $Y=1.835 $X2=0
+ $Y2=0
cc_385 N_A_47_367#_M1004_s N_VPWR_c_510_n 0.00536646f $X=1.08 $Y=1.835 $X2=0
+ $Y2=0
cc_386 N_A_47_367#_M1010_s N_VPWR_c_510_n 0.00536646f $X=1.94 $Y=1.835 $X2=0
+ $Y2=0
cc_387 N_A_47_367#_M1019_s N_VPWR_c_510_n 0.00536646f $X=2.8 $Y=1.835 $X2=0
+ $Y2=0
cc_388 N_A_47_367#_M1029_s N_VPWR_c_510_n 0.00376627f $X=3.66 $Y=1.835 $X2=0
+ $Y2=0
cc_389 N_A_47_367#_M1002_d N_VPWR_c_510_n 0.00223565f $X=4.52 $Y=1.835 $X2=0
+ $Y2=0
cc_390 N_A_47_367#_M1009_d N_VPWR_c_510_n 0.00223565f $X=5.38 $Y=1.835 $X2=0
+ $Y2=0
cc_391 N_A_47_367#_M1015_d N_VPWR_c_510_n 0.00223565f $X=6.24 $Y=1.835 $X2=0
+ $Y2=0
cc_392 N_A_47_367#_M1024_d N_VPWR_c_510_n 0.00215161f $X=7.1 $Y=1.835 $X2=0
+ $Y2=0
cc_393 N_A_47_367#_c_408_n N_VPWR_c_510_n 0.0104192f $X=0.36 $Y=2.91 $X2=0 $Y2=0
cc_394 N_A_47_367#_c_457_p N_VPWR_c_510_n 0.00730901f $X=1.22 $Y=2.91 $X2=0
+ $Y2=0
cc_395 N_A_47_367#_c_454_p N_VPWR_c_510_n 0.00730901f $X=2.08 $Y=2.91 $X2=0
+ $Y2=0
cc_396 N_A_47_367#_c_455_p N_VPWR_c_510_n 0.00730901f $X=2.94 $Y=2.45 $X2=0
+ $Y2=0
cc_397 N_A_47_367#_c_458_p N_VPWR_c_510_n 0.00738676f $X=3.8 $Y=2.905 $X2=0
+ $Y2=0
cc_398 N_A_47_367#_c_437_n N_VPWR_c_510_n 0.023676f $X=4.565 $Y=2.99 $X2=0 $Y2=0
cc_399 N_A_47_367#_c_440_n N_VPWR_c_510_n 0.023676f $X=5.425 $Y=2.99 $X2=0 $Y2=0
cc_400 N_A_47_367#_c_442_n N_VPWR_c_510_n 0.0237058f $X=6.285 $Y=2.985 $X2=0
+ $Y2=0
cc_401 N_A_47_367#_c_410_n N_VPWR_c_510_n 0.033814f $X=7.145 $Y=2.985 $X2=0
+ $Y2=0
cc_402 N_A_47_367#_c_463_p N_VPWR_c_510_n 0.00738676f $X=4.66 $Y=2.99 $X2=0
+ $Y2=0
cc_403 N_A_47_367#_c_464_p N_VPWR_c_510_n 0.00738676f $X=5.52 $Y=2.985 $X2=0
+ $Y2=0
cc_404 N_A_47_367#_c_465_p N_VPWR_c_510_n 0.00738676f $X=6.38 $Y=2.985 $X2=0
+ $Y2=0
cc_405 N_A_47_367#_c_437_n N_Y_M1001_s 0.00332344f $X=4.565 $Y=2.99 $X2=0 $Y2=0
cc_406 N_A_47_367#_c_440_n N_Y_M1007_s 0.00332344f $X=5.425 $Y=2.99 $X2=0 $Y2=0
cc_407 N_A_47_367#_c_442_n N_Y_M1014_s 0.00332931f $X=6.285 $Y=2.985 $X2=0 $Y2=0
cc_408 N_A_47_367#_c_410_n N_Y_M1021_s 0.00332931f $X=7.145 $Y=2.985 $X2=0 $Y2=0
cc_409 N_A_47_367#_M1002_d N_Y_c_626_n 0.001837f $X=4.52 $Y=1.835 $X2=0 $Y2=0
cc_410 N_A_47_367#_c_409_n N_Y_c_626_n 0.0157966f $X=3.705 $Y=1.812 $X2=0 $Y2=0
cc_411 N_A_47_367#_c_439_n N_Y_c_626_n 0.0149669f $X=4.66 $Y=2.425 $X2=0 $Y2=0
cc_412 N_A_47_367#_M1009_d N_Y_c_691_n 0.00332836f $X=5.38 $Y=1.835 $X2=0 $Y2=0
cc_413 N_A_47_367#_c_495_p N_Y_c_691_n 0.0135055f $X=5.52 $Y=2.425 $X2=0 $Y2=0
cc_414 N_A_47_367#_M1015_d N_Y_c_701_n 0.00332836f $X=6.24 $Y=1.835 $X2=0 $Y2=0
cc_415 N_A_47_367#_c_497_p N_Y_c_701_n 0.0135055f $X=6.38 $Y=2.425 $X2=0 $Y2=0
cc_416 N_A_47_367#_M1024_d N_Y_c_639_n 0.00715023f $X=7.1 $Y=1.835 $X2=0 $Y2=0
cc_417 N_A_47_367#_c_411_n N_Y_c_639_n 0.0202165f $X=7.24 $Y=2.425 $X2=0 $Y2=0
cc_418 N_A_47_367#_c_421_n N_Y_c_633_n 0.0063209f $X=2.83 $Y=2.025 $X2=0 $Y2=0
cc_419 N_A_47_367#_c_421_n N_Y_c_634_n 0.0059527f $X=2.83 $Y=2.025 $X2=0 $Y2=0
cc_420 N_A_47_367#_c_409_n N_Y_c_634_n 0.0146262f $X=3.705 $Y=1.812 $X2=0 $Y2=0
cc_421 N_A_47_367#_c_412_n N_Y_c_634_n 0.0141436f $X=2.932 $Y=1.812 $X2=0 $Y2=0
cc_422 N_A_47_367#_c_409_n N_Y_c_670_n 0.0129759f $X=3.705 $Y=1.812 $X2=0 $Y2=0
cc_423 N_A_47_367#_c_442_n N_Y_c_715_n 0.0160814f $X=6.285 $Y=2.985 $X2=0 $Y2=0
cc_424 N_A_47_367#_c_410_n N_Y_c_723_n 0.0160814f $X=7.145 $Y=2.985 $X2=0 $Y2=0
cc_425 N_A_47_367#_c_437_n Y 0.0159805f $X=4.565 $Y=2.99 $X2=0 $Y2=0
cc_426 N_A_47_367#_c_409_n N_Y_c_637_n 0.0288412f $X=3.705 $Y=1.812 $X2=0 $Y2=0
cc_427 N_A_47_367#_c_440_n N_Y_c_737_n 0.0159805f $X=5.425 $Y=2.99 $X2=0 $Y2=0
cc_428 N_VPWR_c_510_n N_Y_M1001_s 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_429 N_VPWR_c_510_n N_Y_M1007_s 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_430 N_VPWR_c_510_n N_Y_M1014_s 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_431 N_VPWR_c_510_n N_Y_M1021_s 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_432 N_Y_c_618_n N_VGND_M1008_d 0.00176461f $X=1.555 $Y=1.16 $X2=0 $Y2=0
cc_433 N_Y_c_621_n N_VGND_M1017_d 0.00176461f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_434 N_Y_c_625_n N_VGND_M1018_s 0.00176461f $X=5.855 $Y=1.17 $X2=0 $Y2=0
cc_435 N_Y_c_628_n N_VGND_M1026_s 0.00176461f $X=6.715 $Y=1.17 $X2=0 $Y2=0
cc_436 N_Y_c_630_n N_VGND_M1030_s 0.00258276f $X=7.425 $Y=1.17 $X2=0 $Y2=0
cc_437 N_Y_c_617_n N_VGND_c_815_n 0.0287988f $X=0.79 $Y=0.48 $X2=0 $Y2=0
cc_438 N_Y_c_619_n N_VGND_c_815_n 0.00502314f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_439 N_Y_c_617_n N_VGND_c_816_n 0.0224866f $X=0.79 $Y=0.48 $X2=0 $Y2=0
cc_440 N_Y_c_618_n N_VGND_c_816_n 0.0170777f $X=1.555 $Y=1.16 $X2=0 $Y2=0
cc_441 N_Y_c_620_n N_VGND_c_816_n 0.0224826f $X=1.65 $Y=0.48 $X2=0 $Y2=0
cc_442 N_Y_c_620_n N_VGND_c_817_n 0.0224826f $X=1.65 $Y=0.48 $X2=0 $Y2=0
cc_443 N_Y_c_621_n N_VGND_c_817_n 0.0170777f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_444 N_Y_c_622_n N_VGND_c_817_n 0.0232405f $X=2.51 $Y=0.47 $X2=0 $Y2=0
cc_445 N_Y_c_622_n N_VGND_c_818_n 0.028306f $X=2.51 $Y=0.47 $X2=0 $Y2=0
cc_446 N_Y_c_623_n N_VGND_c_818_n 0.028306f $X=3.37 $Y=0.47 $X2=0 $Y2=0
cc_447 N_Y_c_634_n N_VGND_c_818_n 0.0225357f $X=3.275 $Y=1.347 $X2=0 $Y2=0
cc_448 N_Y_c_623_n N_VGND_c_819_n 0.028306f $X=3.37 $Y=0.47 $X2=0 $Y2=0
cc_449 N_Y_c_637_n N_VGND_c_819_n 0.0225357f $X=4.065 $Y=1.347 $X2=0 $Y2=0
cc_450 N_Y_c_638_n N_VGND_c_819_n 0.028306f $X=4.23 $Y=0.47 $X2=0 $Y2=0
cc_451 N_Y_c_638_n N_VGND_c_820_n 0.0102275f $X=4.23 $Y=0.47 $X2=0 $Y2=0
cc_452 N_Y_c_624_n N_VGND_c_821_n 0.0299945f $X=5.09 $Y=0.47 $X2=0 $Y2=0
cc_453 N_Y_c_626_n N_VGND_c_821_n 0.0341073f $X=5.245 $Y=1.17 $X2=0 $Y2=0
cc_454 N_Y_c_638_n N_VGND_c_821_n 0.0348527f $X=4.23 $Y=0.47 $X2=0 $Y2=0
cc_455 N_Y_c_624_n N_VGND_c_822_n 0.0236157f $X=5.09 $Y=0.47 $X2=0 $Y2=0
cc_456 N_Y_c_625_n N_VGND_c_822_n 0.0170777f $X=5.855 $Y=1.17 $X2=0 $Y2=0
cc_457 N_Y_c_627_n N_VGND_c_822_n 0.0236157f $X=5.95 $Y=0.47 $X2=0 $Y2=0
cc_458 N_Y_c_627_n N_VGND_c_823_n 0.0236157f $X=5.95 $Y=0.47 $X2=0 $Y2=0
cc_459 N_Y_c_628_n N_VGND_c_823_n 0.0170777f $X=6.715 $Y=1.17 $X2=0 $Y2=0
cc_460 N_Y_c_629_n N_VGND_c_823_n 0.0236157f $X=6.81 $Y=0.47 $X2=0 $Y2=0
cc_461 N_Y_c_629_n N_VGND_c_824_n 0.0236157f $X=6.81 $Y=0.47 $X2=0 $Y2=0
cc_462 N_Y_c_630_n N_VGND_c_824_n 0.0220026f $X=7.425 $Y=1.17 $X2=0 $Y2=0
cc_463 N_Y_c_622_n N_VGND_c_825_n 0.0102275f $X=2.51 $Y=0.47 $X2=0 $Y2=0
cc_464 N_Y_c_623_n N_VGND_c_827_n 0.0102275f $X=3.37 $Y=0.47 $X2=0 $Y2=0
cc_465 N_Y_c_627_n N_VGND_c_829_n 0.0102275f $X=5.95 $Y=0.47 $X2=0 $Y2=0
cc_466 N_Y_c_629_n N_VGND_c_832_n 0.0102275f $X=6.81 $Y=0.47 $X2=0 $Y2=0
cc_467 N_Y_c_617_n N_VGND_c_834_n 0.0105322f $X=0.79 $Y=0.48 $X2=0 $Y2=0
cc_468 N_Y_c_620_n N_VGND_c_835_n 0.00975394f $X=1.65 $Y=0.48 $X2=0 $Y2=0
cc_469 N_Y_c_624_n N_VGND_c_836_n 0.0102275f $X=5.09 $Y=0.47 $X2=0 $Y2=0
cc_470 N_Y_c_617_n N_VGND_c_837_n 0.00765148f $X=0.79 $Y=0.48 $X2=0 $Y2=0
cc_471 N_Y_c_620_n N_VGND_c_837_n 0.0070861f $X=1.65 $Y=0.48 $X2=0 $Y2=0
cc_472 N_Y_c_622_n N_VGND_c_837_n 0.00712543f $X=2.51 $Y=0.47 $X2=0 $Y2=0
cc_473 N_Y_c_623_n N_VGND_c_837_n 0.00712543f $X=3.37 $Y=0.47 $X2=0 $Y2=0
cc_474 N_Y_c_624_n N_VGND_c_837_n 0.00712543f $X=5.09 $Y=0.47 $X2=0 $Y2=0
cc_475 N_Y_c_627_n N_VGND_c_837_n 0.00712543f $X=5.95 $Y=0.47 $X2=0 $Y2=0
cc_476 N_Y_c_629_n N_VGND_c_837_n 0.00712543f $X=6.81 $Y=0.47 $X2=0 $Y2=0
cc_477 N_Y_c_638_n N_VGND_c_837_n 0.00712543f $X=4.23 $Y=0.47 $X2=0 $Y2=0
