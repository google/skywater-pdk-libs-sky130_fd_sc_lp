# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__bufkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__bufkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.775000 0.805000 1.105000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.940800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 0.275000 1.305000 0.775000 ;
        RECT 1.045000 0.775000 2.765000 1.025000 ;
        RECT 1.045000 1.725000 2.765000 1.895000 ;
        RECT 1.045000 1.895000 1.305000 3.060000 ;
        RECT 1.905000 0.275000 2.165000 0.775000 ;
        RECT 1.905000 1.895000 2.165000 3.060000 ;
        RECT 2.255000 1.025000 2.765000 1.725000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.690000 2.810000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.085000  0.275000 0.385000 0.605000 ;
      RECT 0.085000  0.605000 0.255000 1.275000 ;
      RECT 0.085000  1.275000 2.085000 1.535000 ;
      RECT 0.085000  1.535000 0.395000 3.060000 ;
      RECT 0.555000  0.085000 0.830000 0.605000 ;
      RECT 0.565000  1.875000 0.875000 3.060000 ;
      RECT 1.075000  1.205000 2.085000 1.275000 ;
      RECT 1.475000  0.085000 1.730000 0.605000 ;
      RECT 1.475000  2.065000 1.730000 3.075000 ;
      RECT 2.335000  0.085000 2.615000 0.605000 ;
      RECT 2.335000  2.065000 2.620000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.630000  2.725000 0.800000 2.895000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.520000  2.725000 1.690000 2.895000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.390000  2.725000 2.560000 2.895000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_lp__bufkapwr_4
END LIBRARY
