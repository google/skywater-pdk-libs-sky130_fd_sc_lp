* File: sky130_fd_sc_lp__o221a_2.pex.spice
* Created: Wed Sep  2 10:18:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221A_2%C1 1 3 6 8 9 15
c28 6 0 1.27304e-19 $X=0.56 $Y=2.465
c29 1 0 6.95413e-20 $X=0.52 $Y=1.285
r30 15 16 6.10127 $w=3.16e-07 $l=4e-08 $layer=POLY_cond $X=0.52 $Y=1.45 $X2=0.56
+ $Y2=1.45
r31 13 15 36.6076 $w=3.16e-07 $l=2.4e-07 $layer=POLY_cond $X=0.28 $Y=1.45
+ $X2=0.52 $Y2=1.45
r32 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.45 $X2=0.28 $Y2=1.45
r33 9 14 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=0.23 $Y=1.665
+ $X2=0.23 $Y2=1.45
r34 8 14 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.45
r35 4 16 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.615
+ $X2=0.56 $Y2=1.45
r36 4 6 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=0.56 $Y=1.615 $X2=0.56
+ $Y2=2.465
r37 1 15 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.285
+ $X2=0.52 $Y2=1.45
r38 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.52 $Y=1.285 $X2=0.52
+ $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%B1 3 7 8 11 14
c36 8 0 1.27304e-19 $X=1.2 $Y=1.665
c37 3 0 4.83405e-20 $X=0.95 $Y=0.755
r38 11 14 54.0802 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.01 $Y=1.51
+ $X2=1.01 $Y2=1.72
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.51
+ $X2=1.01 $Y2=1.345
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=1.51 $X2=1.01 $Y2=1.51
r41 8 12 5.27625 $w=4.13e-07 $l=1.9e-07 $layer=LI1_cond $X=1.2 $Y=1.552 $X2=1.01
+ $Y2=1.552
r42 7 14 239.393 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.1 $Y=2.465 $X2=1.1
+ $Y2=1.72
r43 3 13 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.95 $Y=0.755
+ $X2=0.95 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%B2 3 7 9 12 13
c39 13 0 4.83405e-20 $X=1.55 $Y=1.5
r40 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.5
+ $X2=1.55 $Y2=1.665
r41 12 14 47.0858 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.55 $Y=1.5 $X2=1.55
+ $Y2=1.33
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.5 $X2=1.55 $Y2=1.5
r43 9 13 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=1.665
+ $X2=1.635 $Y2=1.5
r44 7 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.46 $Y=2.465 $X2=1.46
+ $Y2=1.665
r45 3 14 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=0.755
+ $X2=1.46 $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%A2 3 5 7 8 12 13
c37 13 0 1.60256e-19 $X=2.23 $Y=1.385
c38 12 0 1.85838e-19 $X=2.14 $Y=1.42
r39 11 13 13.9486 $w=3.11e-07 $l=9e-08 $layer=POLY_cond $X=2.14 $Y=1.385
+ $X2=2.23 $Y2=1.385
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.42 $X2=2.14 $Y2=1.42
r41 8 12 7.05871 $w=3.98e-07 $l=2.45e-07 $layer=LI1_cond $X=2.175 $Y=1.665
+ $X2=2.175 $Y2=1.42
r42 5 13 27.8971 $w=3.11e-07 $l=2.75681e-07 $layer=POLY_cond $X=2.41 $Y=1.185
+ $X2=2.23 $Y2=1.385
r43 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.41 $Y=1.185 $X2=2.41
+ $Y2=0.655
r44 1 13 19.8172 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.23 $Y=1.585 $X2=2.23
+ $Y2=1.385
r45 1 3 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.23 $Y=1.585 $X2=2.23
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%A1 1 3 6 8 12 13
c37 13 0 1.48085e-19 $X=2.86 $Y=1.51
c38 6 0 3.46094e-19 $X=2.915 $Y=0.655
r39 12 14 8.89597 $w=2.98e-07 $l=5.5e-08 $layer=POLY_cond $X=2.86 $Y=1.535
+ $X2=2.915 $Y2=1.535
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.86
+ $Y=1.51 $X2=2.86 $Y2=1.51
r41 8 13 6.10934 $w=4.13e-07 $l=2.2e-07 $layer=LI1_cond $X=2.64 $Y=1.552
+ $X2=2.86 $Y2=1.552
r42 4 14 18.8112 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.915 $Y=1.345
+ $X2=2.915 $Y2=1.535
r43 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.915 $Y=1.345
+ $X2=2.915 $Y2=0.655
r44 1 12 43.6711 $w=2.98e-07 $l=3.5242e-07 $layer=POLY_cond $X=2.59 $Y=1.725
+ $X2=2.86 $Y2=1.535
r45 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.59 $Y=1.725 $X2=2.59
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%A_36_67# 1 2 3 12 16 20 24 28 32 35 36 37 40
+ 42 45 49 56 60 66
c119 16 0 3.06591e-19 $X=3.36 $Y=2.465
r120 66 67 2.21101 $w=3.27e-07 $l=1.5e-08 $layer=POLY_cond $X=3.775 $Y=1.51
+ $X2=3.79 $Y2=1.51
r121 63 64 2.21101 $w=3.27e-07 $l=1.5e-08 $layer=POLY_cond $X=3.345 $Y=1.51
+ $X2=3.36 $Y2=1.51
r122 61 66 50.1162 $w=3.27e-07 $l=3.4e-07 $layer=POLY_cond $X=3.435 $Y=1.51
+ $X2=3.775 $Y2=1.51
r123 61 64 11.055 $w=3.27e-07 $l=7.5e-08 $layer=POLY_cond $X=3.435 $Y=1.51
+ $X2=3.36 $Y2=1.51
r124 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.435
+ $Y=1.51 $X2=3.435 $Y2=1.51
r125 57 60 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=3.21 $Y=1.525
+ $X2=3.435 $Y2=1.525
r126 44 57 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.21 $Y=1.645
+ $X2=3.21 $Y2=1.525
r127 44 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.21 $Y=1.645
+ $X2=3.21 $Y2=1.93
r128 43 56 13.5049 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=2.195 $Y=2.015
+ $X2=1.852 $Y2=2.015
r129 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.125 $Y=2.015
+ $X2=3.21 $Y2=1.93
r130 42 43 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.125 $Y=2.015
+ $X2=2.195 $Y2=2.015
r131 38 56 2.81621 $w=6.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.852 $Y=2.1
+ $X2=1.852 $Y2=2.015
r132 38 40 14.1434 $w=6.83e-07 $l=8.1e-07 $layer=LI1_cond $X=1.852 $Y=2.1
+ $X2=1.852 $Y2=2.91
r133 37 54 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.015
+ $X2=0.63 $Y2=2.015
r134 36 56 13.5049 $w=1.7e-07 $l=3.42e-07 $layer=LI1_cond $X=1.51 $Y=2.015
+ $X2=1.852 $Y2=2.015
r135 36 37 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.51 $Y=2.015
+ $X2=0.715 $Y2=2.015
r136 35 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=1.93
+ $X2=0.63 $Y2=2.015
r137 34 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=1.03
+ $X2=0.63 $Y2=0.945
r138 34 35 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=0.63 $Y=1.03 $X2=0.63
+ $Y2=1.93
r139 30 54 19.1155 $w=1.68e-07 $l=2.93e-07 $layer=LI1_cond $X=0.337 $Y=2.015
+ $X2=0.63 $Y2=2.015
r140 30 32 29.6342 $w=3.13e-07 $l=8.1e-07 $layer=LI1_cond $X=0.337 $Y=2.1
+ $X2=0.337 $Y2=2.91
r141 26 49 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.27 $Y=0.945
+ $X2=0.63 $Y2=0.945
r142 26 28 16.8434 $w=2.58e-07 $l=3.8e-07 $layer=LI1_cond $X=0.27 $Y=0.86
+ $X2=0.27 $Y2=0.48
r143 22 67 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=1.675
+ $X2=3.79 $Y2=1.51
r144 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.79 $Y=1.675
+ $X2=3.79 $Y2=2.465
r145 18 66 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.775 $Y=1.345
+ $X2=3.775 $Y2=1.51
r146 18 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.775 $Y=1.345
+ $X2=3.775 $Y2=0.655
r147 14 64 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=1.675
+ $X2=3.36 $Y2=1.51
r148 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.36 $Y=1.675
+ $X2=3.36 $Y2=2.465
r149 10 63 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.345
+ $X2=3.345 $Y2=1.51
r150 10 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.345 $Y=1.345
+ $X2=3.345 $Y2=0.655
r151 3 56 200 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=3 $X=1.535
+ $Y=1.835 $X2=1.675 $Y2=2.015
r152 3 40 200 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=3 $X=1.535
+ $Y=1.835 $X2=1.675 $Y2=2.91
r153 2 30 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.835 $X2=0.345 $Y2=2.015
r154 2 32 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.835 $X2=0.345 $Y2=2.91
r155 1 26 182 $w=1.7e-07 $l=6.69589e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.335 $X2=0.305 $Y2=0.945
r156 1 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.335 $X2=0.305 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%VPWR 1 2 3 14 18 20 22 26 28 33 39 42 48
r54 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 43 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 42 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 37 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 34 42 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.31 $Y=3.33
+ $X2=2.975 $Y2=3.33
r63 34 36 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.31 $Y=3.33 $X2=3.6
+ $Y2=3.33
r64 33 47 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.84 $Y=3.33 $X2=4.08
+ $Y2=3.33
r65 33 36 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.84 $Y=3.33 $X2=3.6
+ $Y2=3.33
r66 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r68 29 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.83 $Y2=3.33
r69 29 31 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 28 42 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=2.975 $Y2=3.33
r71 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r72 26 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 26 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r74 22 25 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.005 $Y=2.25
+ $X2=4.005 $Y2=2.95
r75 20 47 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=4.005 $Y=3.245
+ $X2=4.08 $Y2=3.33
r76 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.005 $Y=3.245
+ $X2=4.005 $Y2=2.95
r77 16 42 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=3.245
+ $X2=2.975 $Y2=3.33
r78 16 18 15.5312 $w=6.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.975 $Y=3.245
+ $X2=2.975 $Y2=2.375
r79 12 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=3.245
+ $X2=0.83 $Y2=3.33
r80 12 14 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.83 $Y=3.245
+ $X2=0.83 $Y2=2.375
r81 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.835 $X2=4.005 $Y2=2.95
r82 3 22 400 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.835 $X2=4.005 $Y2=2.25
r83 2 18 150 $w=1.7e-07 $l=7.42159e-07 $layer=licon1_PDIFF $count=4 $X=2.665
+ $Y=1.835 $X2=3.145 $Y2=2.375
r84 1 14 300 $w=1.7e-07 $l=6.3e-07 $layer=licon1_PDIFF $count=2 $X=0.635
+ $Y=1.835 $X2=0.83 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%X 1 2 9 15 17 18 19 20 28 36
c31 15 0 1.58506e-19 $X=3.995 $Y=1.815
r32 34 36 1.59477 $w=4.48e-07 $l=6e-08 $layer=LI1_cond $X=3.995 $Y=1.235
+ $X2=3.995 $Y2=1.295
r33 26 34 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.555 $Y=1.15
+ $X2=3.995 $Y2=1.15
r34 19 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=1.15
+ $X2=3.995 $Y2=1.15
r35 19 20 9.51547 $w=4.48e-07 $l=3.58e-07 $layer=LI1_cond $X=3.995 $Y=1.307
+ $X2=3.995 $Y2=1.665
r36 19 36 0.318954 $w=4.48e-07 $l=1.2e-08 $layer=LI1_cond $X=3.995 $Y=1.307
+ $X2=3.995 $Y2=1.295
r37 18 26 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=3.555 $Y=0.925
+ $X2=3.555 $Y2=1.065
r38 17 18 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.555 $Y=0.555
+ $X2=3.555 $Y2=0.925
r39 17 28 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=3.555 $Y=0.555
+ $X2=3.555 $Y2=0.42
r40 15 20 3.98693 $w=4.48e-07 $l=1.5e-07 $layer=LI1_cond $X=3.995 $Y=1.815
+ $X2=3.995 $Y2=1.665
r41 12 15 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.575 $Y=1.9
+ $X2=3.995 $Y2=1.9
r42 7 12 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=1.985
+ $X2=3.575 $Y2=1.9
r43 7 9 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=3.575 $Y=1.985
+ $X2=3.575 $Y2=2.91
r44 2 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.835 $X2=3.575 $Y2=1.98
r45 2 9 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.835 $X2=3.575 $Y2=2.91
r46 1 28 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.235 $X2=3.56 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%A_119_67# 1 2 7 11 13
c24 7 0 6.95413e-20 $X=1.57 $Y=0.34
r25 13 16 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.735 $Y=0.34
+ $X2=0.735 $Y2=0.565
r26 9 11 10.0305 $w=2.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.705 $Y=0.425
+ $X2=1.705 $Y2=0.66
r27 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=0.34 $X2=0.735
+ $Y2=0.34
r28 7 9 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.57 $Y=0.34
+ $X2=1.705 $Y2=0.425
r29 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.57 $Y=0.34 $X2=0.9
+ $Y2=0.34
r30 2 11 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.335 $X2=1.675 $Y2=0.66
r31 1 16 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.335 $X2=0.735 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%A_205_67# 1 2 9 11 12 15
r27 13 15 21.376 $w=3.08e-07 $l=5.75e-07 $layer=LI1_cond $X=2.685 $Y=0.995
+ $X2=2.685 $Y2=0.42
r28 11 13 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.53 $Y=1.08
+ $X2=2.685 $Y2=0.995
r29 11 12 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.53 $Y=1.08
+ $X2=1.4 $Y2=1.08
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.235 $Y=0.995
+ $X2=1.4 $Y2=1.08
r31 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.235 $Y=0.995
+ $X2=1.235 $Y2=0.68
r32 2 15 91 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.235 $X2=2.68 $Y2=0.42
r33 1 9 91 $w=1.7e-07 $l=4.37579e-07 $layer=licon1_NDIFF $count=2 $X=1.025
+ $Y=0.335 $X2=1.235 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_2%VGND 1 2 3 12 16 18 20 22 24 32 37 43 46 50
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r55 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r56 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r57 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 38 46 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.132
+ $Y2=0
r59 38 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.6
+ $Y2=0
r60 37 49 4.37118 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=4.087
+ $Y2=0
r61 37 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.6
+ $Y2=0
r62 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r63 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r64 33 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.195
+ $Y2=0
r65 33 35 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.64
+ $Y2=0
r66 32 46 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=3.132
+ $Y2=0
r67 32 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.64
+ $Y2=0
r68 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 27 31 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r70 26 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r71 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r72 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.195
+ $Y2=0
r73 24 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.68
+ $Y2=0
r74 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r75 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r76 22 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r77 18 49 3.14649 $w=3e-07 $l=1.19143e-07 $layer=LI1_cond $X=4.005 $Y=0.085
+ $X2=4.087 $Y2=0
r78 18 20 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=4.005 $Y=0.085
+ $X2=4.005 $Y2=0.38
r79 14 46 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.132 $Y=0.085
+ $X2=3.132 $Y2=0
r80 14 16 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=3.132 $Y=0.085
+ $X2=3.132 $Y2=0.38
r81 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r82 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.38
r83 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.85
+ $Y=0.235 $X2=3.99 $Y2=0.38
r84 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.99
+ $Y=0.235 $X2=3.13 $Y2=0.38
r85 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.07
+ $Y=0.235 $X2=2.195 $Y2=0.38
.ends

