# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__busdriver2_20
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__busdriver2_20 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  24.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.016000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.830000 1.180000 24.835000 1.515000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.180000 0.445000 1.515000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  5.250200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.750000 0.645000 15.400000 0.895000 ;
        RECT 11.305000 0.895000 12.235000 1.505000 ;
        RECT 11.305000 1.505000 20.820000 1.725000 ;
        RECT 11.305000 1.725000 13.010000 1.780000 ;
        RECT 12.820000 1.780000 13.010000 2.715000 ;
        RECT 13.680000 1.725000 13.870000 2.715000 ;
        RECT 14.540000 1.725000 14.730000 2.715000 ;
        RECT 15.400000 1.725000 15.590000 2.715000 ;
        RECT 16.260000 1.725000 16.450000 2.715000 ;
        RECT 16.270000 1.495000 20.820000 1.505000 ;
        RECT 17.120000 1.725000 17.310000 2.715000 ;
        RECT 17.980000 1.725000 18.170000 2.715000 ;
        RECT 18.840000 1.725000 19.030000 2.715000 ;
        RECT 19.700000 1.725000 19.890000 2.715000 ;
        RECT 20.570000 1.725000 20.820000 2.805000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 24.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 24.960000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 25.150000 3.520000 ;
        RECT 11.730000 1.345000 20.980000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 24.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 24.960000 0.085000 ;
      RECT  0.000000  3.245000 24.960000 3.415000 ;
      RECT  0.115000  0.085000  0.445000 1.000000 ;
      RECT  0.115000  1.815000  0.445000 3.245000 ;
      RECT  0.625000  0.265000  0.795000 0.625000 ;
      RECT  0.625000  0.625000  2.360000 0.795000 ;
      RECT  0.625000  0.795000  0.795000 3.065000 ;
      RECT  0.975000  1.815000  1.225000 3.245000 ;
      RECT  1.055000  0.085000  1.385000 0.445000 ;
      RECT  1.405000  1.815000  2.595000 1.985000 ;
      RECT  1.405000  1.985000  1.735000 3.065000 ;
      RECT  1.680000  0.975000  2.010000 1.815000 ;
      RECT  1.915000  2.165000  2.085000 3.245000 ;
      RECT  2.190000  0.795000  2.360000 1.005000 ;
      RECT  2.190000  1.005000  6.150000 1.335000 ;
      RECT  2.265000  1.515000  9.780000 1.685000 ;
      RECT  2.265000  1.685000  2.595000 1.815000 ;
      RECT  2.265000  1.985000  2.595000 3.065000 ;
      RECT  2.340000  0.085000  2.670000 0.445000 ;
      RECT  2.775000  1.855000  2.945000 3.245000 ;
      RECT  2.900000  0.265000  3.230000 0.655000 ;
      RECT  2.900000  0.655000  6.990000 0.825000 ;
      RECT  3.125000  1.865000 10.355000 2.035000 ;
      RECT  3.125000  2.035000  3.455000 2.765000 ;
      RECT  3.410000  0.085000  3.740000 0.475000 ;
      RECT  3.625000  2.205000  3.815000 3.245000 ;
      RECT  3.920000  0.265000  4.090000 0.655000 ;
      RECT  3.985000  2.035000  4.315000 2.765000 ;
      RECT  4.270000  0.085000  4.600000 0.475000 ;
      RECT  4.485000  2.205000  4.675000 3.245000 ;
      RECT  4.780000  0.265000  4.950000 0.655000 ;
      RECT  4.845000  2.035000  5.175000 2.765000 ;
      RECT  5.130000  0.085000  5.460000 0.475000 ;
      RECT  5.345000  2.205000  5.535000 3.245000 ;
      RECT  5.640000  0.265000  5.970000 0.655000 ;
      RECT  5.705000  2.035000  6.035000 2.765000 ;
      RECT  6.150000  0.085000  6.480000 0.475000 ;
      RECT  6.205000  2.205000  6.395000 3.245000 ;
      RECT  6.390000  1.345000  9.780000 1.515000 ;
      RECT  6.565000  2.035000  6.895000 2.765000 ;
      RECT  6.660000  0.265000  6.990000 0.655000 ;
      RECT  6.660000  0.825000  6.990000 0.995000 ;
      RECT  6.660000  0.995000  9.570000 1.165000 ;
      RECT  7.065000  2.205000  7.255000 3.245000 ;
      RECT  7.170000  0.085000  7.340000 0.815000 ;
      RECT  7.425000  2.035000  7.755000 2.765000 ;
      RECT  7.520000  0.265000  7.850000 0.995000 ;
      RECT  7.925000  2.205000  8.115000 3.245000 ;
      RECT  8.030000  0.085000  8.200000 0.815000 ;
      RECT  8.305000  2.035000  8.635000 2.765000 ;
      RECT  8.380000  0.265000  8.710000 0.995000 ;
      RECT  8.805000  2.205000  8.995000 3.245000 ;
      RECT  8.890000  0.085000  9.060000 0.815000 ;
      RECT  9.165000  2.035000  9.495000 2.765000 ;
      RECT  9.240000  0.265000 15.910000 0.475000 ;
      RECT  9.240000  0.475000  9.570000 0.995000 ;
      RECT  9.665000  2.205000  9.855000 3.245000 ;
      RECT 10.025000  1.465000 11.135000 1.635000 ;
      RECT 10.025000  1.635000 10.355000 1.865000 ;
      RECT 10.025000  2.035000 10.355000 3.065000 ;
      RECT 10.535000  1.815000 10.705000 3.245000 ;
      RECT 10.885000  1.635000 11.135000 1.960000 ;
      RECT 10.885000  1.960000 12.650000 2.185000 ;
      RECT 10.885000  2.185000 11.135000 3.065000 ;
      RECT 11.315000  2.365000 11.645000 3.245000 ;
      RECT 12.320000  2.185000 12.650000 2.885000 ;
      RECT 12.320000  2.885000 20.390000 3.065000 ;
      RECT 12.405000  1.075000 21.650000 1.315000 ;
      RECT 12.405000  1.315000 15.455000 1.325000 ;
      RECT 13.180000  1.895000 13.510000 2.885000 ;
      RECT 14.040000  1.895000 14.370000 2.885000 ;
      RECT 14.900000  1.895000 15.230000 2.885000 ;
      RECT 15.580000  0.475000 15.910000 0.805000 ;
      RECT 15.660000  0.985000 23.380000 1.000000 ;
      RECT 15.660000  1.000000 21.650000 1.075000 ;
      RECT 15.760000  1.895000 16.090000 2.885000 ;
      RECT 16.620000  1.895000 16.950000 2.885000 ;
      RECT 17.480000  1.895000 17.810000 2.885000 ;
      RECT 18.340000  1.895000 18.670000 2.885000 ;
      RECT 19.200000  1.895000 19.530000 2.885000 ;
      RECT 20.060000  1.895000 20.390000 2.885000 ;
      RECT 21.050000  1.815000 21.300000 3.245000 ;
      RECT 21.480000  0.830000 23.380000 0.985000 ;
      RECT 21.480000  1.315000 21.650000 1.695000 ;
      RECT 21.480000  1.695000 24.415000 1.865000 ;
      RECT 21.480000  1.865000 21.810000 3.065000 ;
      RECT 21.520000  0.085000 21.850000 0.650000 ;
      RECT 21.990000  2.165000 22.160000 3.245000 ;
      RECT 22.030000  0.295000 22.360000 0.830000 ;
      RECT 22.340000  1.865000 22.670000 3.065000 ;
      RECT 22.540000  0.085000 22.870000 0.650000 ;
      RECT 22.850000  2.045000 23.020000 3.245000 ;
      RECT 23.050000  0.265000 23.380000 0.830000 ;
      RECT 23.200000  1.865000 23.530000 3.065000 ;
      RECT 23.560000  0.085000 23.890000 1.000000 ;
      RECT 23.710000  2.045000 23.880000 3.245000 ;
      RECT 24.085000  1.865000 24.415000 3.065000 ;
      RECT 24.595000  1.815000 24.845000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.245000 18.565000 3.415000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.245000 19.045000 3.415000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.245000 19.525000 3.415000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.245000 20.005000 3.415000 ;
      RECT 20.315000 -0.085000 20.485000 0.085000 ;
      RECT 20.315000  3.245000 20.485000 3.415000 ;
      RECT 20.795000 -0.085000 20.965000 0.085000 ;
      RECT 20.795000  3.245000 20.965000 3.415000 ;
      RECT 21.275000 -0.085000 21.445000 0.085000 ;
      RECT 21.275000  3.245000 21.445000 3.415000 ;
      RECT 21.755000 -0.085000 21.925000 0.085000 ;
      RECT 21.755000  3.245000 21.925000 3.415000 ;
      RECT 22.235000 -0.085000 22.405000 0.085000 ;
      RECT 22.235000  3.245000 22.405000 3.415000 ;
      RECT 22.715000 -0.085000 22.885000 0.085000 ;
      RECT 22.715000  3.245000 22.885000 3.415000 ;
      RECT 23.195000 -0.085000 23.365000 0.085000 ;
      RECT 23.195000  3.245000 23.365000 3.415000 ;
      RECT 23.675000 -0.085000 23.845000 0.085000 ;
      RECT 23.675000  3.245000 23.845000 3.415000 ;
      RECT 24.155000 -0.085000 24.325000 0.085000 ;
      RECT 24.155000  3.245000 24.325000 3.415000 ;
      RECT 24.635000 -0.085000 24.805000 0.085000 ;
      RECT 24.635000  3.245000 24.805000 3.415000 ;
  END
END sky130_fd_sc_lp__busdriver2_20
END LIBRARY
