* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1960_125# a_773_409# a_1751_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 VPWR SET_B a_1960_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_1858_463# a_2205_231# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 Q a_2638_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_2638_53# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR a_2638_53# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_1960_125# a_2205_231# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_218_119# D a_304_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1888_125# a_961_491# a_1960_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_1598_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND SCE a_346_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_2638_53# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_1858_463# a_961_491# a_1960_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 Q a_2638_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_2638_53# a_1960_125# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_1211_463# a_773_409# a_1297_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_1297_463# a_1339_331# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_1315_81# a_1339_331# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_218_119# a_961_491# a_1211_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VGND SCD a_146_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1211_463# a_1751_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 Q a_2638_53# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_773_409# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_218_119# a_346_93# a_27_479# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 VPWR SCE a_346_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_2163_125# a_2205_231# a_2248_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1339_331# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 VGND a_2638_53# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 VPWR SCE a_196_479# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_1960_125# a_773_409# a_2163_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_196_479# D a_218_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 VPWR a_1211_463# a_1339_331# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 a_773_409# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_218_119# a_773_409# a_1211_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND a_1211_463# a_1888_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 Q a_2638_53# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 a_2638_53# a_1960_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 a_1211_463# a_961_491# a_1315_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_1339_331# a_1211_463# a_1598_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_146_119# SCE a_218_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VGND a_773_409# a_961_491# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_2248_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 VPWR a_773_409# a_961_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_27_479# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X44 a_304_119# a_346_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 VPWR a_1960_125# a_2205_231# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
