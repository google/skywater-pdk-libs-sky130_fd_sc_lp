* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_271_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR B1 a_505_529# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_505_529# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_571_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_271_47# a_91_269# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A1_N a_271_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_91_269# B2 a_571_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR A1_N a_271_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 X a_91_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 X a_91_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_91_269# a_271_47# a_505_529# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_271_367# A2_N a_271_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
