* File: sky130_fd_sc_lp__a41oi_0.spice
* Created: Fri Aug 28 10:03:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a41oi_0  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_B1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1007 A_230_47# N_A1_M1007_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.063
+ AS=0.0756 PD=0.72 PS=0.78 NRD=27.132 NRS=17.136 M=1 R=2.8 SA=75000.7
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1005 A_320_47# N_A2_M1005_g A_230_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.063 PD=0.84 PS=0.72 NRD=44.28 NRS=27.132 M=1 R=2.8 SA=75001.1 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1003 A_434_47# N_A3_M1003_g A_320_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0882 PD=0.84 PS=0.84 NRD=44.28 NRS=44.28 M=1 R=2.8 SA=75001.7 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A4_M1008_g A_434_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0882 PD=1.37 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75002.3 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_176_479#_M1001_d N_B1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_176_479#_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1004 N_A_176_479#_M1004_d N_A2_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A3_M1000_g N_A_176_479#_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_176_479#_M1002_d N_A4_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_70 VPB 0 1.83885e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a41oi_0.pxi.spice"
*
.ends
*
*
