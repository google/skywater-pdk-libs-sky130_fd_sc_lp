# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o311ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o311ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.180000 1.860000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.180000 3.795000 1.435000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.465000 1.425000 6.095000 1.750000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.265000 1.425000 7.615000 1.750000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.785000 1.425000 9.995000 1.750000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  3.061800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.080000 1.085000 9.430000 1.255000 ;
        RECT 4.080000 1.255000 4.295000 1.920000 ;
        RECT 4.080000 1.920000 9.570000 2.090000 ;
        RECT 4.080000 2.090000 6.920000 2.120000 ;
        RECT 4.080000 2.120000 4.340000 2.735000 ;
        RECT 5.010000 2.120000 5.200000 2.735000 ;
        RECT 5.870000 2.120000 6.060000 3.075000 ;
        RECT 6.730000 2.120000 6.920000 3.075000 ;
        RECT 7.590000 2.090000 7.780000 3.075000 ;
        RECT 8.100000 0.595000 8.430000 1.085000 ;
        RECT 8.450000 2.090000 8.640000 3.075000 ;
        RECT 9.100000 0.595000 9.430000 1.085000 ;
        RECT 9.310000 2.090000 9.570000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.110000  0.085000  0.440000 1.010000 ;
      RECT 0.110000  1.605000  3.880000 1.775000 ;
      RECT 0.110000  1.775000  0.370000 3.075000 ;
      RECT 0.540000  1.945000  0.870000 3.245000 ;
      RECT 0.610000  0.255000  0.800000 0.840000 ;
      RECT 0.610000  0.840000  7.430000 0.915000 ;
      RECT 0.610000  0.915000  3.910000 1.010000 ;
      RECT 0.970000  0.085000  1.300000 0.670000 ;
      RECT 1.040000  1.775000  1.230000 3.075000 ;
      RECT 1.400000  1.945000  1.730000 3.245000 ;
      RECT 1.470000  0.255000  1.660000 0.840000 ;
      RECT 1.830000  0.085000  2.160000 0.670000 ;
      RECT 1.900000  1.775000  2.090000 3.075000 ;
      RECT 2.260000  1.945000  2.590000 2.905000 ;
      RECT 2.260000  2.905000  5.700000 3.075000 ;
      RECT 2.330000  0.255000  2.520000 0.840000 ;
      RECT 2.690000  0.085000  3.020000 0.670000 ;
      RECT 2.760000  1.775000  2.950000 2.735000 ;
      RECT 3.120000  1.945000  3.450000 2.905000 ;
      RECT 3.190000  0.255000  3.380000 0.745000 ;
      RECT 3.190000  0.745000  7.430000 0.840000 ;
      RECT 3.550000  0.085000  3.880000 0.575000 ;
      RECT 3.620000  1.775000  3.880000 2.735000 ;
      RECT 4.050000  0.255000  4.240000 0.745000 ;
      RECT 4.410000  0.085000  4.740000 0.575000 ;
      RECT 4.510000  2.290000  4.840000 2.905000 ;
      RECT 4.910000  0.255000  5.100000 0.725000 ;
      RECT 4.910000  0.725000  7.430000 0.745000 ;
      RECT 5.270000  0.085000  5.600000 0.555000 ;
      RECT 5.370000  2.290000  5.700000 2.905000 ;
      RECT 5.810000  0.255000  9.860000 0.425000 ;
      RECT 5.810000  0.425000  7.930000 0.555000 ;
      RECT 6.230000  2.290000  6.560000 3.245000 ;
      RECT 7.090000  2.260000  7.420000 3.245000 ;
      RECT 7.600000  0.555000  7.930000 0.915000 ;
      RECT 7.950000  2.260000  8.280000 3.245000 ;
      RECT 8.600000  0.425000  8.930000 0.915000 ;
      RECT 8.810000  2.260000  9.140000 3.245000 ;
      RECT 9.600000  0.425000  9.860000 1.190000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__o311ai_4
END LIBRARY
