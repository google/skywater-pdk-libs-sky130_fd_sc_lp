* File: sky130_fd_sc_lp__o31ai_0.pex.spice
* Created: Wed Sep  2 10:25:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31AI_0%A1 2 3 5 6 8 12 15 18 20 21 22 23 29
r40 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.02 $X2=0.27 $Y2=1.02
r41 22 23 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.247 $Y=1.665
+ $X2=0.247 $Y2=2.035
r42 21 22 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.247 $Y=1.295
+ $X2=0.247 $Y2=1.665
r43 21 30 9.75144 $w=3.23e-07 $l=2.75e-07 $layer=LI1_cond $X=0.247 $Y=1.295
+ $X2=0.247 $Y2=1.02
r44 20 30 3.36868 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=0.247 $Y=0.925
+ $X2=0.247 $Y2=1.02
r45 16 18 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.36 $Y=2.23
+ $X2=0.655 $Y2=2.23
r46 14 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.36
+ $X2=0.27 $Y2=1.02
r47 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.36
+ $X2=0.27 $Y2=1.525
r48 10 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.005
+ $X2=0.27 $Y2=1.02
r49 10 12 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.27 $Y=0.93
+ $X2=0.615 $Y2=0.93
r50 6 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.655 $Y=2.305
+ $X2=0.655 $Y2=2.23
r51 6 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.655 $Y=2.305
+ $X2=0.655 $Y2=2.735
r52 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=0.855
+ $X2=0.615 $Y2=0.93
r53 3 5 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.615 $Y=0.855
+ $X2=0.615 $Y2=0.535
r54 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.155
+ $X2=0.36 $Y2=2.23
r55 2 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.155
+ $X2=0.36 $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_0%A2 2 5 9 11 12 13 14 19
r50 19 21 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.897 $Y=1.41
+ $X2=0.897 $Y2=1.245
r51 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.41 $X2=0.84 $Y2=1.41
r52 13 14 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.792 $Y=1.665
+ $X2=0.792 $Y2=2.035
r53 13 20 6.91466 $w=4.23e-07 $l=2.55e-07 $layer=LI1_cond $X=0.792 $Y=1.665
+ $X2=0.792 $Y2=1.41
r54 12 20 3.11838 $w=4.23e-07 $l=1.15e-07 $layer=LI1_cond $X=0.792 $Y=1.295
+ $X2=0.792 $Y2=1.41
r55 9 11 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.045 $Y=2.735
+ $X2=1.045 $Y2=1.915
r56 5 21 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.045 $Y=0.535
+ $X2=1.045 $Y2=1.245
r57 2 11 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=0.897 $Y=1.693
+ $X2=0.897 $Y2=1.915
r58 1 19 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.897 $Y=1.467
+ $X2=0.897 $Y2=1.41
r59 1 2 28.2451 $w=4.45e-07 $l=2.26e-07 $layer=POLY_cond $X=0.897 $Y=1.467
+ $X2=0.897 $Y2=1.693
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_0%A3 3 7 11 12 13 14 18 19
c42 3 0 2.2249e-20 $X=1.435 $Y=2.735
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.525
+ $Y=1.27 $X2=1.525 $Y2=1.27
r44 13 14 8.27194 $w=5.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.627 $Y=1.295
+ $X2=1.627 $Y2=1.665
r45 13 19 0.558915 $w=5.33e-07 $l=2.5e-08 $layer=LI1_cond $X=1.627 $Y=1.295
+ $X2=1.627 $Y2=1.27
r46 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.525 $Y=1.61
+ $X2=1.525 $Y2=1.27
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.61
+ $X2=1.525 $Y2=1.775
r48 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.105
+ $X2=1.525 $Y2=1.27
r49 7 10 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.575 $Y=0.535
+ $X2=1.575 $Y2=1.105
r50 3 12 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.435 $Y=2.735
+ $X2=1.435 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_0%B1 3 7 9 11 14 16 17 18 19 24 26
c45 17 0 2.2249e-20 $X=2.16 $Y=0.925
r46 24 26 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.127 $Y=1.02
+ $X2=2.127 $Y2=0.855
r47 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.02 $X2=2.16 $Y2=1.02
r48 18 19 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r49 18 25 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.02
r50 17 25 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=1.02
r51 12 14 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.865 $Y=2.09
+ $X2=2.005 $Y2=2.09
r52 11 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.005 $Y=2.015
+ $X2=2.005 $Y2=2.09
r53 11 16 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.005 $Y=2.015
+ $X2=2.005 $Y2=1.525
r54 9 16 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=2.127 $Y=1.328
+ $X2=2.127 $Y2=1.525
r55 8 24 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=2.127 $Y=1.052
+ $X2=2.127 $Y2=1.02
r56 8 9 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=2.127 $Y=1.052
+ $X2=2.127 $Y2=1.328
r57 7 26 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.005 $Y=0.535
+ $X2=2.005 $Y2=0.855
r58 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.865 $Y=2.165
+ $X2=1.865 $Y2=2.09
r59 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.865 $Y=2.165
+ $X2=1.865 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_0%VPWR 1 2 9 13 16 17 18 23 32 33 36
r28 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 33 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 30 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.115 $Y2=3.33
r32 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r36 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 23 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.115 $Y2=3.33
r38 23 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 22 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 18 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 18 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 16 21 2.51176 $w=1.7e-07 $l=3.5e-08 $layer=LI1_cond $X=0.275 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=3.33
+ $X2=0.44 $Y2=3.33
r45 15 25 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.44 $Y2=3.33
r47 11 36 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=3.245
+ $X2=2.115 $Y2=3.33
r48 11 13 30.3624 $w=2.58e-07 $l=6.85e-07 $layer=LI1_cond $X=2.115 $Y=3.245
+ $X2=2.115 $Y2=2.56
r49 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.44 $Y=3.245 $X2=0.44
+ $Y2=3.33
r50 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.44 $Y=3.245
+ $X2=0.44 $Y2=2.56
r51 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=2.415 $X2=2.08 $Y2=2.56
r52 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.315
+ $Y=2.415 $X2=0.44 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_0%Y 1 2 7 8 9 14 15 16 17 18 19 20 36 37
r40 20 37 2.87555 $w=3.65e-07 $l=1.22e-07 $layer=LI1_cond $X=2.607 $Y=2.102
+ $X2=2.607 $Y2=1.98
r41 20 37 0.473607 $w=3.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.607 $Y=1.965
+ $X2=2.607 $Y2=1.98
r42 19 20 9.47213 $w=3.63e-07 $l=3e-07 $layer=LI1_cond $X=2.607 $Y=1.665
+ $X2=2.607 $Y2=1.965
r43 18 19 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.607 $Y=1.295
+ $X2=2.607 $Y2=1.665
r44 17 18 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.607 $Y=0.925
+ $X2=2.607 $Y2=1.295
r45 17 36 8.05131 $w=3.63e-07 $l=2.55e-07 $layer=LI1_cond $X=2.607 $Y=0.925
+ $X2=2.607 $Y2=0.67
r46 16 36 3.25197 $w=3.65e-07 $l=1.65e-07 $layer=LI1_cond $X=2.607 $Y=0.505
+ $X2=2.607 $Y2=0.67
r47 15 32 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.65 $Y=2.775
+ $X2=1.65 $Y2=2.56
r48 14 32 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.65 $Y=2.405
+ $X2=1.65 $Y2=2.56
r49 13 14 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.65 $Y=2.225
+ $X2=1.65 $Y2=2.405
r50 9 16 3.58703 $w=3.3e-07 $l=1.82e-07 $layer=LI1_cond $X=2.425 $Y=0.505
+ $X2=2.607 $Y2=0.505
r51 9 11 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.425 $Y=0.505
+ $X2=2.22 $Y2=0.505
r52 8 13 7.01204 $w=2.45e-07 $l=2.17991e-07 $layer=LI1_cond $X=1.815 $Y=2.102
+ $X2=1.65 $Y2=2.225
r53 7 20 4.28975 $w=2.45e-07 $l=1.82e-07 $layer=LI1_cond $X=2.425 $Y=2.102
+ $X2=2.607 $Y2=2.102
r54 7 8 28.6935 $w=2.43e-07 $l=6.1e-07 $layer=LI1_cond $X=2.425 $Y=2.102
+ $X2=1.815 $Y2=2.102
r55 2 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=2.415 $X2=1.65 $Y2=2.56
r56 1 16 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.325 $X2=2.56 $Y2=0.505
r57 1 11 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.08 $Y=0.325
+ $X2=2.22 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_0%VGND 1 2 7 9 11 15 17 24 25 31
r32 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r34 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r36 22 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r37 21 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r38 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r39 19 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.31
+ $Y2=0
r40 19 21 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.68
+ $Y2=0
r41 17 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r42 17 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r43 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0
r44 13 15 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0.49
r45 12 28 4.52228 $w=1.7e-07 $l=2.83e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.282
+ $Y2=0
r46 11 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=1.31
+ $Y2=0
r47 11 12 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=0.565
+ $Y2=0
r48 7 28 3.2439 $w=3.3e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.4 $Y=0.085
+ $X2=0.282 $Y2=0
r49 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.4 $Y=0.085 $X2=0.4
+ $Y2=0.535
r50 2 15 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.325 $X2=1.31 $Y2=0.49
r51 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.325 $X2=0.4 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_0%A_138_65# 1 2 9 11 12 15
c29 15 0 1.95508e-19 $X=1.79 $Y=0.535
r30 13 15 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.77 $Y=0.765
+ $X2=1.77 $Y2=0.535
r31 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.645 $Y=0.85
+ $X2=1.77 $Y2=0.765
r32 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.645 $Y=0.85
+ $X2=0.975 $Y2=0.85
r33 7 12 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.855 $Y=0.765
+ $X2=0.975 $Y2=0.85
r34 7 9 11.0442 $w=2.38e-07 $l=2.3e-07 $layer=LI1_cond $X=0.855 $Y=0.765
+ $X2=0.855 $Y2=0.535
r35 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.325 $X2=1.79 $Y2=0.535
r36 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.325 $X2=0.83 $Y2=0.535
.ends

