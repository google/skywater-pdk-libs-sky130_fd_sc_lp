* File: sky130_fd_sc_lp__o41a_2.pex.spice
* Created: Wed Sep  2 10:27:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41A_2%A_102_53# 1 2 7 9 12 14 16 19 21 25 28 31 33
+ 34 37 40 47 48
c87 40 0 1.52271e-19 $X=1.757 $Y=1.51
r88 47 48 7.73305 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=2.495
+ $X2=2.405 $Y2=2.33
r89 37 39 16.7296 $w=5.78e-07 $l=6.5e-07 $layer=LI1_cond $X=1.91 $Y=0.39
+ $X2=1.91 $Y2=1.04
r90 34 48 8.58683 $w=2.53e-07 $l=1.9e-07 $layer=LI1_cond $X=2.197 $Y=2.14
+ $X2=2.197 $Y2=2.33
r91 33 34 27.1111 $w=1.78e-07 $l=4.4e-07 $layer=LI1_cond $X=1.757 $Y=2.05
+ $X2=2.197 $Y2=2.05
r92 32 40 5.99569 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=1.757 $Y=1.675
+ $X2=1.757 $Y2=1.51
r93 32 33 11.9435 $w=2.73e-07 $l=2.85e-07 $layer=LI1_cond $X=1.757 $Y=1.675
+ $X2=1.757 $Y2=1.96
r94 31 40 5.99569 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=1.757 $Y=1.345
+ $X2=1.757 $Y2=1.51
r95 31 39 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=1.757 $Y=1.345
+ $X2=1.757 $Y2=1.04
r96 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.495
+ $Y=1.51 $X2=1.495 $Y2=1.51
r97 25 40 0.695019 $w=3.3e-07 $l=1.37e-07 $layer=LI1_cond $X=1.62 $Y=1.51
+ $X2=1.757 $Y2=1.51
r98 25 27 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.62 $Y=1.51
+ $X2=1.495 $Y2=1.51
r99 22 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.585 $Y=1.51
+ $X2=1.015 $Y2=1.51
r100 21 28 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.09 $Y=1.51
+ $X2=1.495 $Y2=1.51
r101 21 24 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.09 $Y=1.51
+ $X2=1.015 $Y2=1.51
r102 17 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=1.51
r103 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=2.465
r104 14 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.345
+ $X2=1.015 $Y2=1.51
r105 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.015 $Y=1.345
+ $X2=1.015 $Y2=0.815
r106 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=1.51
r107 10 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=2.465
r108 7 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.345
+ $X2=0.585 $Y2=1.51
r109 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.585 $Y=1.345
+ $X2=0.585 $Y2=0.815
r110 2 47 150 $w=1.7e-07 $l=8.6741e-07 $layer=licon1_PDIFF $count=4 $X=2.095
+ $Y=1.835 $X2=2.575 $Y2=2.495
r111 2 34 600 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.835 $X2=2.235 $Y2=2.125
r112 1 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.91
+ $Y=0.245 $X2=2.035 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%B1 3 5 7 8 9 17
c40 8 0 1.93916e-19 $X=2.16 $Y=1.295
r41 15 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.16 $Y=1.375 $X2=2.25
+ $Y2=1.375
r42 12 15 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.02 $Y=1.375
+ $X2=2.16 $Y2=1.375
r43 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295 $X2=2.16
+ $Y2=1.665
r44 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.375 $X2=2.16 $Y2=1.375
r45 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.21
+ $X2=2.25 $Y2=1.375
r46 5 7 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.25 $Y=1.21 $X2=2.25
+ $Y2=0.665
r47 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.02 $Y=1.54
+ $X2=2.02 $Y2=1.375
r48 1 3 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.02 $Y=1.54 $X2=2.02
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%A4 3 7 9 10 14 15
c44 7 0 1.93916e-19 $X=2.79 $Y=2.465
r45 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.51 $X2=2.7
+ $Y2=1.675
r46 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.51 $X2=2.7
+ $Y2=1.345
r47 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.51 $X2=2.7 $Y2=1.51
r48 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.655 $Y=1.665
+ $X2=2.655 $Y2=2.035
r49 9 15 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=2.655 $Y=1.665
+ $X2=2.655 $Y2=1.51
r50 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.79 $Y=2.465
+ $X2=2.79 $Y2=1.675
r51 3 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.725 $Y=0.665
+ $X2=2.725 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%A3 3 7 9 10 11 12 18 19
r39 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.51
+ $X2=3.24 $Y2=1.675
r40 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.51
+ $X2=3.24 $Y2=1.345
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.51 $X2=3.24 $Y2=1.51
r42 11 12 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.155 $Y=2.405
+ $X2=3.155 $Y2=2.775
r43 10 11 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.155 $Y=2.035
+ $X2=3.155 $Y2=2.405
r44 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.155 $Y=1.665
+ $X2=3.155 $Y2=2.035
r45 9 19 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.155 $Y=1.665
+ $X2=3.155 $Y2=1.51
r46 7 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.26 $Y=0.665
+ $X2=3.26 $Y2=1.345
r47 3 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.15 $Y=2.465
+ $X2=3.15 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%A2 3 7 9 10 11 12 26 27
c36 26 0 1.77152e-19 $X=3.78 $Y=1.51
r37 26 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.51
+ $X2=3.78 $Y2=1.675
r38 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.51
+ $X2=3.78 $Y2=1.345
r39 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.51 $X2=3.78 $Y2=1.51
r40 11 12 6.50807 $w=6.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.835 $Y=2.405
+ $X2=3.835 $Y2=2.775
r41 10 11 6.50807 $w=6.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.835 $Y=2.035
+ $X2=3.835 $Y2=2.405
r42 9 10 6.50807 $w=6.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.835 $Y=1.665
+ $X2=3.835 $Y2=2.035
r43 9 27 2.72636 $w=6.78e-07 $l=1.55e-07 $layer=LI1_cond $X=3.835 $Y=1.665
+ $X2=3.835 $Y2=1.51
r44 7 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.69 $Y=2.465
+ $X2=3.69 $Y2=1.675
r45 3 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.69 $Y=0.665
+ $X2=3.69 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%A1 3 7 9 14 15
c25 15 0 1.77152e-19 $X=4.51 $Y=1.46
r26 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.46 $X2=4.51 $Y2=1.46
r27 11 14 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=4.23 $Y=1.46
+ $X2=4.51 $Y2=1.46
r28 9 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.51 $Y=1.665
+ $X2=4.51 $Y2=1.46
r29 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.625
+ $X2=4.23 $Y2=1.46
r30 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.23 $Y=1.625 $X2=4.23
+ $Y2=2.465
r31 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.295
+ $X2=4.23 $Y2=1.46
r32 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.23 $Y=1.295 $X2=4.23
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%VPWR 1 2 3 10 12 18 21 22 24 29 31 33 38 50
+ 54
r60 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 42 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 41 44 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r68 39 50 14.9498 $w=1.7e-07 $l=4.18e-07 $layer=LI1_cond $X=1.9 $Y=3.33
+ $X2=1.482 $Y2=3.33
r69 39 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.9 $Y=3.33 $X2=2.16
+ $Y2=3.33
r70 38 53 4.09313 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.572 $Y2=3.33
r71 38 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.08 $Y2=3.33
r72 37 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 34 47 3.99156 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r76 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 33 50 14.9498 $w=1.7e-07 $l=4.17e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.482 $Y2=3.33
r78 33 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 31 45 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=4.08 $Y2=3.33
r80 31 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r81 29 30 5.86895 $w=8.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.482 $Y=2.475
+ $X2=1.482 $Y2=2.31
r82 24 27 36.7074 $w=2.68e-07 $l=8.6e-07 $layer=LI1_cond $X=4.48 $Y=2.09
+ $X2=4.48 $Y2=2.95
r83 22 53 3.19156 $w=2.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.572 $Y2=3.33
r84 22 27 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.95
r85 21 50 3.21326 $w=8.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.482 $Y=3.245
+ $X2=1.482 $Y2=3.33
r86 20 29 3.60972 $w=8.33e-07 $l=2.52e-07 $layer=LI1_cond $X=1.482 $Y=2.727
+ $X2=1.482 $Y2=2.475
r87 20 21 7.41998 $w=8.33e-07 $l=5.18e-07 $layer=LI1_cond $X=1.482 $Y=2.727
+ $X2=1.482 $Y2=3.245
r88 18 30 9.87808 $w=3.83e-07 $l=3.3e-07 $layer=LI1_cond $X=1.257 $Y=1.98
+ $X2=1.257 $Y2=2.31
r89 12 15 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=0.335 $Y=1.98
+ $X2=0.335 $Y2=2.95
r90 10 47 3.22066 $w=2.6e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.232 $Y2=3.33
r91 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.335 $Y2=2.95
r92 3 27 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.835 $X2=4.45 $Y2=2.95
r93 3 24 400 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.835 $X2=4.45 $Y2=2.09
r94 2 29 150 $w=1.7e-07 $l=9.84289e-07 $layer=licon1_PDIFF $count=4 $X=1.09
+ $Y=1.835 $X2=1.805 $Y2=2.475
r95 2 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.835 $X2=1.23 $Y2=1.98
r96 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.95
r97 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%X 1 2 7 8 9 10 11 12 13
r16 13 39 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.765 $Y=2.775
+ $X2=0.765 $Y2=2.91
r17 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.405
+ $X2=0.765 $Y2=2.775
r18 11 12 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=0.765 $Y=1.98
+ $X2=0.765 $Y2=2.405
r19 10 11 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.765 $Y=1.665
+ $X2=0.765 $Y2=1.98
r20 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=1.295
+ $X2=0.765 $Y2=1.665
r21 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=0.925
+ $X2=0.765 $Y2=1.295
r22 7 8 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0.54
+ $X2=0.765 $Y2=0.925
r23 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.91
r24 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=1.98
r25 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.395 $X2=0.8 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%VGND 1 2 3 4 13 15 19 23 27 30 31 33 34 35 37
+ 53 54 60
r58 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r61 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r62 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r63 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r64 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r65 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r66 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r67 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 42 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.23
+ $Y2=0
r69 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.68
+ $Y2=0
r70 41 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r71 41 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r72 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r73 38 57 3.99156 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.232
+ $Y2=0
r74 38 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.72
+ $Y2=0
r75 37 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.23
+ $Y2=0
r76 37 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r77 35 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r78 35 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r79 33 50 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.6 $Y2=0
r80 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.965
+ $Y2=0
r81 32 53 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.13 $Y=0 $X2=4.56
+ $Y2=0
r82 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.13 $Y=0 $X2=3.965
+ $Y2=0
r83 30 47 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=0 $X2=2.64
+ $Y2=0
r84 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=0 $X2=2.995
+ $Y2=0
r85 29 50 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.16 $Y=0 $X2=3.6
+ $Y2=0
r86 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=0 $X2=2.995
+ $Y2=0
r87 25 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=0.085
+ $X2=3.965 $Y2=0
r88 25 27 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.965 $Y=0.085
+ $X2=3.965 $Y2=0.37
r89 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0
r90 21 23 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0.37
r91 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r92 17 19 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.54
r93 13 57 3.22066 $w=2.6e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.232 $Y2=0
r94 13 15 20.1678 $w=2.58e-07 $l=4.55e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.54
r95 4 27 91 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=2 $X=3.765
+ $Y=0.245 $X2=3.965 $Y2=0.37
r96 3 23 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=2.8 $Y=0.245
+ $X2=2.995 $Y2=0.37
r97 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.395 $X2=1.23 $Y2=0.54
r98 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.395 $X2=0.37 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_2%A_465_49# 1 2 3 12 14 15 18 20 24 26
r50 22 24 21.7477 $w=3.08e-07 $l=5.85e-07 $layer=LI1_cond $X=4.455 $Y=1.005
+ $X2=4.455 $Y2=0.42
r51 21 26 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.63 $Y=1.09 $X2=3.48
+ $Y2=1.09
r52 20 22 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=4.3 $Y=1.09
+ $X2=4.455 $Y2=1.005
r53 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.3 $Y=1.09 $X2=3.63
+ $Y2=1.09
r54 16 26 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=1.005 $X2=3.48
+ $Y2=1.09
r55 16 18 22.4726 $w=2.98e-07 $l=5.85e-07 $layer=LI1_cond $X=3.48 $Y=1.005
+ $X2=3.48 $Y2=0.42
r56 14 26 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.33 $Y=1.09 $X2=3.48
+ $Y2=1.09
r57 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.33 $Y=1.09
+ $X2=2.66 $Y2=1.09
r58 10 15 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=2.542 $Y=1.005
+ $X2=2.66 $Y2=1.09
r59 10 12 28.6885 $w=2.33e-07 $l=5.85e-07 $layer=LI1_cond $X=2.542 $Y=1.005
+ $X2=2.542 $Y2=0.42
r60 3 24 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.245 $X2=4.445 $Y2=0.42
r61 2 18 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.335
+ $Y=0.245 $X2=3.475 $Y2=0.42
r62 1 12 91 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.245 $X2=2.51 $Y2=0.42
.ends

