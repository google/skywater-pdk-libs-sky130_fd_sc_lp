* File: sky130_fd_sc_lp__or3_2.pex.spice
* Created: Wed Sep  2 10:30:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3_2%C 3 7 9 10 11 16
c31 16 0 8.25848e-20 $X=0.51 $Y=1.415
r32 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.415
+ $X2=0.51 $Y2=1.58
r33 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.415
+ $X2=0.51 $Y2=1.25
r34 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.415 $X2=0.51 $Y2=1.415
r35 11 30 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=0.75 $Y=2.035
+ $X2=0.75 $Y2=1.775
r36 10 30 5.26802 $w=4.48e-07 $l=1.1e-07 $layer=LI1_cond $X=0.65 $Y=1.665
+ $X2=0.65 $Y2=1.775
r37 10 17 6.64488 $w=4.48e-07 $l=2.5e-07 $layer=LI1_cond $X=0.65 $Y=1.665
+ $X2=0.65 $Y2=1.415
r38 9 17 3.18954 $w=4.48e-07 $l=1.2e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.415
r39 7 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.585 $Y=2.045
+ $X2=0.585 $Y2=1.58
r40 3 18 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.515 $Y=0.51
+ $X2=0.515 $Y2=1.25
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_2%B 3 5 7 9 10 11 19
c33 19 0 8.25848e-20 $X=1.195 $Y=1.205
c34 7 0 1.45091e-19 $X=1.285 $Y=0.51
r35 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.205 $X2=1.195 $Y2=1.205
r36 15 18 38.1986 $w=3.55e-07 $l=2.35e-07 $layer=POLY_cond $X=0.96 $Y=1.192
+ $X2=1.195 $Y2=1.192
r37 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.665
+ $X2=1.195 $Y2=2.035
r38 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.665
r39 9 19 3.45733 $w=2.98e-07 $l=9e-08 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.205
r40 5 18 14.6292 $w=3.55e-07 $l=9e-08 $layer=POLY_cond $X=1.285 $Y=1.192
+ $X2=1.195 $Y2=1.192
r41 5 7 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.285 $Y=1.015
+ $X2=1.285 $Y2=0.51
r42 1 15 22.9692 $w=1.5e-07 $l=1.78e-07 $layer=POLY_cond $X=0.96 $Y=1.37
+ $X2=0.96 $Y2=1.192
r43 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.96 $Y=1.37 $X2=0.96
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_2%A 1 3 4 5 8 10 11 15
c45 15 0 2.86103e-20 $X=1.8 $Y=1.415
r46 15 18 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.8 $Y=1.415 $X2=1.8
+ $Y2=1.655
r47 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.415
+ $X2=1.8 $Y2=1.25
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.8
+ $Y=1.415 $X2=1.8 $Y2=1.415
r49 11 16 6.64488 $w=4.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.74 $Y=1.665
+ $X2=1.74 $Y2=1.415
r50 10 16 3.18954 $w=4.48e-07 $l=1.2e-07 $layer=LI1_cond $X=1.74 $Y=1.295
+ $X2=1.74 $Y2=1.415
r51 8 17 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.715 $Y=0.51
+ $X2=1.715 $Y2=1.25
r52 4 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.655
+ $X2=1.8 $Y2=1.655
r53 4 5 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.635 $Y=1.655
+ $X2=1.395 $Y2=1.655
r54 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.32 $Y=1.73
+ $X2=1.395 $Y2=1.655
r55 1 3 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.32 $Y=1.73 $X2=1.32
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_2%A_35_60# 1 2 3 10 12 15 17 19 22 26 29 30 34
+ 36 38 42 46 48 49 51 52 53
c96 48 0 2.86103e-20 $X=1.535 $Y=0.72
c97 34 0 1.45091e-19 $X=1.5 $Y=0.445
r98 58 59 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=2.735 $Y=1.415
+ $X2=2.765 $Y2=1.415
r99 57 58 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=2.335 $Y=1.415
+ $X2=2.735 $Y2=1.415
r100 55 57 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=2.305 $Y=1.415
+ $X2=2.335 $Y2=1.415
r101 52 59 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.975 $Y=1.415
+ $X2=2.765 $Y2=1.415
r102 51 53 2.34452 $w=4.43e-07 $l=8.5e-08 $layer=LI1_cond $X=3.032 $Y=1.415
+ $X2=3.032 $Y2=1.33
r103 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.415 $X2=2.975 $Y2=1.415
r104 43 46 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.17 $Y=2.11 $X2=0.37
+ $Y2=2.11
r105 40 53 16.9985 $w=3.98e-07 $l=5.9e-07 $layer=LI1_cond $X=3.055 $Y=0.74
+ $X2=3.055 $Y2=1.33
r106 38 40 8.37092 $w=1.7e-07 $l=2.38747e-07 $layer=LI1_cond $X=2.855 $Y=0.655
+ $X2=3.055 $Y2=0.74
r107 38 49 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.855 $Y=0.655
+ $X2=2.08 $Y2=0.655
r108 37 48 5.61476 $w=2.35e-07 $l=1.3e-07 $layer=LI1_cond $X=1.665 $Y=0.72
+ $X2=1.535 $Y2=0.72
r109 36 49 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.93 $Y=0.72
+ $X2=2.08 $Y2=0.72
r110 36 37 10.1799 $w=2.98e-07 $l=2.65e-07 $layer=LI1_cond $X=1.93 $Y=0.72
+ $X2=1.665 $Y2=0.72
r111 32 48 0.981169 $w=2.6e-07 $l=1.5e-07 $layer=LI1_cond $X=1.535 $Y=0.57
+ $X2=1.535 $Y2=0.72
r112 32 34 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=1.535 $Y=0.57
+ $X2=1.535 $Y2=0.445
r113 31 42 2.60907 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=0.785
+ $X2=0.24 $Y2=0.785
r114 30 48 5.61476 $w=2.35e-07 $l=1.59217e-07 $layer=LI1_cond $X=1.405 $Y=0.785
+ $X2=1.535 $Y2=0.72
r115 30 31 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.405 $Y=0.785
+ $X2=0.395 $Y2=0.785
r116 29 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=1.945
+ $X2=0.17 $Y2=2.11
r117 28 42 3.84343 $w=2.4e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.17 $Y=0.87
+ $X2=0.24 $Y2=0.785
r118 28 29 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=0.17 $Y=0.87
+ $X2=0.17 $Y2=1.945
r119 24 42 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=0.7 $X2=0.24
+ $Y2=0.785
r120 24 26 7.06336 $w=3.08e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=0.7
+ $X2=0.24 $Y2=0.51
r121 20 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.58
+ $X2=2.765 $Y2=1.415
r122 20 22 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=2.765 $Y=1.58
+ $X2=2.765 $Y2=2.465
r123 17 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.25
+ $X2=2.735 $Y2=1.415
r124 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.735 $Y=1.25
+ $X2=2.735 $Y2=0.72
r125 13 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.58
+ $X2=2.335 $Y2=1.415
r126 13 15 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=2.335 $Y=1.58
+ $X2=2.335 $Y2=2.465
r127 10 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.25
+ $X2=2.305 $Y2=1.415
r128 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.305 $Y=1.25
+ $X2=2.305 $Y2=0.72
r129 3 46 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.11
r130 2 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.3 $X2=1.5 $Y2=0.445
r131 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.3 $X2=0.3 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_2%VPWR 1 2 9 14 16 20 22 30 36 40
r24 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r25 34 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r26 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r27 31 36 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=1.865 $Y2=3.33
r28 31 33 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.64 $Y2=3.33
r29 30 39 3.90852 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.127 $Y2=3.33
r30 30 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 22 36 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.865 $Y2=3.33
r36 22 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 20 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 20 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 16 19 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=3.02 $Y=1.98
+ $X2=3.02 $Y2=2.95
r41 14 39 3.23464 $w=2.5e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.127 $Y2=3.33
r42 14 19 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=2.95
r43 9 13 7.77451 $w=6.98e-07 $l=4.55e-07 $layer=LI1_cond $X=1.865 $Y=2.085
+ $X2=1.865 $Y2=2.54
r44 7 36 2.86223 $w=7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.865 $Y=3.245 $X2=1.865
+ $Y2=3.33
r45 7 13 12.0462 $w=6.98e-07 $l=7.05e-07 $layer=LI1_cond $X=1.865 $Y=3.245
+ $X2=1.865 $Y2=2.54
r46 2 19 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.835 $X2=2.98 $Y2=2.95
r47 2 16 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.835 $X2=2.98 $Y2=1.98
r48 1 13 300 $w=1.7e-07 $l=1.01821e-06 $layer=licon1_PDIFF $count=2 $X=1.395
+ $Y=1.835 $X2=2.12 $Y2=2.54
r49 1 9 600 $w=1.7e-07 $l=8.40759e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.835 $X2=2.12 $Y2=2.085
r50 1 9 600 $w=1.7e-07 $l=3.37268e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.835 $X2=1.6 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_2%X 1 2 10 13 14 15 30 33
r25 20 33 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.555 $Y=2.04
+ $X2=2.555 $Y2=2.035
r26 15 27 5.93169 $w=3.38e-07 $l=1.75e-07 $layer=LI1_cond $X=2.555 $Y=2.775
+ $X2=2.555 $Y2=2.95
r27 14 15 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.555 $Y=2.405
+ $X2=2.555 $Y2=2.775
r28 13 33 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=2.555 $Y=1.995
+ $X2=2.555 $Y2=2.035
r29 13 30 4.98306 $w=3.38e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=1.995
+ $X2=2.555 $Y2=1.87
r30 13 14 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=2.555 $Y=2.08
+ $X2=2.555 $Y2=2.405
r31 13 20 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=2.555 $Y=2.08
+ $X2=2.555 $Y2=2.04
r32 12 30 32.0876 $w=2.53e-07 $l=7.1e-07 $layer=LI1_cond $X=2.512 $Y=1.16
+ $X2=2.512 $Y2=1.87
r33 10 12 6.3875 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=1.16
r34 2 33 400 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.835 $X2=2.55 $Y2=2.035
r35 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.835 $X2=2.55 $Y2=2.95
r36 1 10 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.3 $X2=2.52 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_2%VGND 1 2 3 10 11 17 28 35 38 40 41
r46 40 43 10.248 $w=3.75e-07 $l=3.15e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.13
+ $Y2=0.315
r47 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 37 38 10.2539 $w=6.13e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0.222
+ $X2=1.235 $Y2=0.222
r49 33 37 6.80695 $w=6.13e-07 $l=3.5e-07 $layer=LI1_cond $X=0.72 $Y=0.222
+ $X2=1.07 $Y2=0.222
r50 33 35 10.0594 $w=6.13e-07 $l=1.55e-07 $layer=LI1_cond $X=0.72 $Y=0.222
+ $X2=0.565 $Y2=0.222
r51 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 31 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r53 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 28 40 5.38787 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.13
+ $Y2=0
r55 28 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.64
+ $Y2=0
r56 26 38 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.235
+ $Y2=0
r57 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r58 21 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.565
+ $Y2=0
r59 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 17 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r61 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r62 17 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r63 13 30 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.64
+ $Y2=0
r64 11 26 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.68
+ $Y2=0
r65 10 15 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.01
+ $Y2=0.315
r66 10 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.175
+ $Y2=0
r67 10 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.845
+ $Y2=0
r68 3 43 182 $w=1.7e-07 $l=2.62393e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.3 $X2=3.065 $Y2=0.315
r69 2 15 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.3 $X2=2.01 $Y2=0.315
r70 1 37 91 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.3 $X2=1.07 $Y2=0.445
.ends

