* File: sky130_fd_sc_lp__nand4b_2.pxi.spice
* Created: Fri Aug 28 10:51:41 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4B_2%A_N N_A_N_c_89_n N_A_N_M1013_g N_A_N_c_91_n
+ N_A_N_c_92_n N_A_N_M1010_g A_N N_A_N_c_94_n N_A_N_c_95_n
+ PM_SKY130_FD_SC_LP__NAND4B_2%A_N
x_PM_SKY130_FD_SC_LP__NAND4B_2%A_27_51# N_A_27_51#_M1013_s N_A_27_51#_M1010_s
+ N_A_27_51#_M1002_g N_A_27_51#_M1003_g N_A_27_51#_M1009_g N_A_27_51#_M1015_g
+ N_A_27_51#_c_127_n N_A_27_51#_c_128_n N_A_27_51#_c_129_n N_A_27_51#_c_130_n
+ N_A_27_51#_c_131_n N_A_27_51#_c_132_n N_A_27_51#_c_138_n N_A_27_51#_c_133_n
+ N_A_27_51#_c_134_n PM_SKY130_FD_SC_LP__NAND4B_2%A_27_51#
x_PM_SKY130_FD_SC_LP__NAND4B_2%B N_B_M1000_g N_B_M1001_g N_B_M1008_g N_B_M1016_g
+ B B N_B_c_210_n PM_SKY130_FD_SC_LP__NAND4B_2%B
x_PM_SKY130_FD_SC_LP__NAND4B_2%C N_C_M1006_g N_C_M1004_g N_C_M1012_g N_C_M1011_g
+ C C C N_C_c_263_n PM_SKY130_FD_SC_LP__NAND4B_2%C
x_PM_SKY130_FD_SC_LP__NAND4B_2%D N_D_M1005_g N_D_M1007_g N_D_M1017_g N_D_M1014_g
+ D D N_D_c_316_n PM_SKY130_FD_SC_LP__NAND4B_2%D
x_PM_SKY130_FD_SC_LP__NAND4B_2%VPWR N_VPWR_M1010_d N_VPWR_M1015_s N_VPWR_M1008_s
+ N_VPWR_M1011_d N_VPWR_M1017_d N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n
+ N_VPWR_c_356_n N_VPWR_c_357_n VPWR N_VPWR_c_358_n N_VPWR_c_359_n
+ N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n
+ N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_352_n PM_SKY130_FD_SC_LP__NAND4B_2%VPWR
x_PM_SKY130_FD_SC_LP__NAND4B_2%Y N_Y_M1002_s N_Y_M1003_d N_Y_M1001_d N_Y_M1004_s
+ N_Y_M1007_s N_Y_c_429_n N_Y_c_431_n N_Y_c_473_n N_Y_c_433_n N_Y_c_425_n
+ N_Y_c_426_n N_Y_c_427_n N_Y_c_459_n N_Y_c_467_n N_Y_c_480_n Y Y Y Y
+ N_Y_c_452_n N_Y_c_463_n N_Y_c_487_n N_Y_c_489_n PM_SKY130_FD_SC_LP__NAND4B_2%Y
x_PM_SKY130_FD_SC_LP__NAND4B_2%VGND N_VGND_M1013_d N_VGND_M1005_d N_VGND_c_504_n
+ N_VGND_c_505_n VGND N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n
+ N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n PM_SKY130_FD_SC_LP__NAND4B_2%VGND
x_PM_SKY130_FD_SC_LP__NAND4B_2%A_217_65# N_A_217_65#_M1002_d N_A_217_65#_M1009_d
+ N_A_217_65#_M1016_s N_A_217_65#_c_561_n N_A_217_65#_c_562_n
+ N_A_217_65#_c_563_n N_A_217_65#_c_574_n N_A_217_65#_c_576_n
+ N_A_217_65#_c_564_n N_A_217_65#_c_577_n PM_SKY130_FD_SC_LP__NAND4B_2%A_217_65#
x_PM_SKY130_FD_SC_LP__NAND4B_2%A_486_65# N_A_486_65#_M1000_d N_A_486_65#_M1006_d
+ N_A_486_65#_c_602_n N_A_486_65#_c_609_n N_A_486_65#_c_603_n
+ PM_SKY130_FD_SC_LP__NAND4B_2%A_486_65#
x_PM_SKY130_FD_SC_LP__NAND4B_2%A_697_69# N_A_697_69#_M1006_s N_A_697_69#_M1012_s
+ N_A_697_69#_M1014_s N_A_697_69#_c_630_n N_A_697_69#_c_631_n
+ N_A_697_69#_c_632_n N_A_697_69#_c_633_n N_A_697_69#_c_634_n
+ N_A_697_69#_c_635_n N_A_697_69#_c_636_n PM_SKY130_FD_SC_LP__NAND4B_2%A_697_69#
cc_1 VNB N_A_N_c_89_n 0.0299002f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.475
cc_2 VNB N_A_N_M1013_g 0.0364358f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.465
cc_3 VNB N_A_N_c_91_n 0.0206306f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.55
cc_4 VNB N_A_N_c_92_n 0.0322613f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.55
cc_5 VNB N_A_N_M1010_g 0.00162716f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=2.045
cc_6 VNB N_A_N_c_94_n 0.0329282f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_7 VNB N_A_N_c_95_n 0.0218556f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_8 VNB N_A_27_51#_M1002_g 0.0236126f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.625
cc_9 VNB N_A_27_51#_M1009_g 0.0201042f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_10 VNB N_A_27_51#_c_127_n 8.72418e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_51#_c_128_n 0.00564986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_51#_c_129_n 0.00836417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_51#_c_130_n 0.0113195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_51#_c_131_n 3.11366e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_51#_c_132_n 0.0137481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_51#_c_133_n 0.00116895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_51#_c_134_n 0.0482443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_M1000_g 0.021176f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.955
cc_19 VNB N_B_M1016_g 0.0245929f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.12
cc_20 VNB B 0.00325317f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=0.955
cc_21 VNB N_B_c_210_n 0.0398398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C_M1006_g 0.0226489f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.955
cc_23 VNB N_C_M1012_g 0.0188729f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=2.045
cc_24 VNB C 0.0107209f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.33
cc_25 VNB N_C_c_263_n 0.0403828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_D_M1005_g 0.0188362f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.955
cc_27 VNB N_D_M1014_g 0.025218f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.12
cc_28 VNB D 0.013634f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=0.955
cc_29 VNB N_D_c_316_n 0.0375798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_352_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_425_n 0.00814296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_426_n 0.00243326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_427_n 0.00676451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_504_n 0.00742391f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.625
cc_35 VNB N_VGND_c_505_n 0.00332106f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_VGND_c_506_n 0.0155965f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_37 VNB N_VGND_c_507_n 0.0940105f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.33
cc_38 VNB N_VGND_c_508_n 0.0187923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_509_n 0.329517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_510_n 0.0052564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_511_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_217_65#_c_561_n 0.0103234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_217_65#_c_562_n 0.00483879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_217_65#_c_563_n 0.0036506f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.12
cc_45 VNB N_A_217_65#_c_564_n 0.00375694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_486_65#_c_602_n 0.0190164f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.55
cc_47 VNB N_A_486_65#_c_603_n 0.00287674f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_48 VNB N_A_697_69#_c_630_n 0.00624587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_697_69#_c_631_n 0.0029562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_697_69#_c_632_n 0.00499518f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.12
cc_51 VNB N_A_697_69#_c_633_n 0.00198077f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=0.955
cc_52 VNB N_A_697_69#_c_634_n 0.0135017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_697_69#_c_635_n 0.0319312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_697_69#_c_636_n 0.0018781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_A_N_M1010_g 0.0321181f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.045
cc_56 VPB N_A_27_51#_M1003_g 0.022671f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_57 VPB N_A_27_51#_M1015_g 0.019398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_27_51#_c_131_n 0.00622732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_27_51#_c_138_n 0.0147537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_27_51#_c_134_n 0.0117219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_B_M1001_g 0.0192086f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.55
cc_62 VPB N_B_M1008_g 0.0209365f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.045
cc_63 VPB B 0.00594436f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=0.955
cc_64 VPB N_B_c_210_n 0.00520336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_C_M1004_g 0.0221579f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.55
cc_66 VPB N_C_M1011_g 0.0180996f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.12
cc_67 VPB C 0.0106347f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.33
cc_68 VPB N_C_c_263_n 0.00769096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_D_M1007_g 0.0183815f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.55
cc_70 VPB N_D_M1017_g 0.0235869f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.045
cc_71 VPB D 0.0122034f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=0.955
cc_72 VPB N_D_c_316_n 0.00523381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_353_n 0.039802f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=0.955
cc_74 VPB N_VPWR_c_354_n 0.00437047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_355_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_356_n 0.0132106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_357_n 0.0483636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_358_n 0.0325333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_359_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_360_n 0.0150212f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_361_n 0.0129657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_362_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_363_n 0.00728331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_364_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_365_n 0.0206365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_366_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_352_n 0.0833059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_Y_c_427_n 0.00477356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 N_A_N_M1010_g N_A_27_51#_M1003_g 0.00904884f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_90 N_A_N_M1013_g N_A_27_51#_c_127_n 0.00103344f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_91 N_A_N_M1013_g N_A_27_51#_c_128_n 0.0177406f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_92 N_A_N_c_91_n N_A_27_51#_c_128_n 0.00117147f $X=0.725 $Y=1.55 $X2=0 $Y2=0
cc_93 N_A_N_c_94_n N_A_27_51#_c_128_n 0.0015658f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_94 N_A_N_c_95_n N_A_27_51#_c_128_n 0.0069087f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_95 N_A_N_c_94_n N_A_27_51#_c_129_n 0.00557802f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_96 N_A_N_c_95_n N_A_27_51#_c_129_n 0.0164461f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_97 N_A_N_M1013_g N_A_27_51#_c_130_n 0.0163472f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_98 N_A_N_c_95_n N_A_27_51#_c_130_n 0.0286701f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_99 N_A_N_M1010_g N_A_27_51#_c_131_n 0.00874929f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_100 N_A_N_c_91_n N_A_27_51#_c_132_n 0.00399141f $X=0.725 $Y=1.55 $X2=0 $Y2=0
cc_101 N_A_N_M1010_g N_A_27_51#_c_132_n 0.00438871f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_102 N_A_N_c_91_n N_A_27_51#_c_138_n 4.61577e-19 $X=0.725 $Y=1.55 $X2=0 $Y2=0
cc_103 N_A_N_c_92_n N_A_27_51#_c_138_n 0.00677539f $X=0.55 $Y=1.55 $X2=0 $Y2=0
cc_104 N_A_N_M1010_g N_A_27_51#_c_138_n 0.00682939f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_105 N_A_N_c_95_n N_A_27_51#_c_138_n 8.77496e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_106 N_A_N_c_89_n N_A_27_51#_c_133_n 7.78185e-19 $X=0.327 $Y=1.475 $X2=0 $Y2=0
cc_107 N_A_N_c_91_n N_A_27_51#_c_133_n 0.0113747f $X=0.725 $Y=1.55 $X2=0 $Y2=0
cc_108 N_A_N_M1010_g N_A_27_51#_c_133_n 4.247e-19 $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_109 N_A_N_c_95_n N_A_27_51#_c_133_n 0.017002f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_110 N_A_N_c_89_n N_A_27_51#_c_134_n 0.00214754f $X=0.327 $Y=1.475 $X2=0 $Y2=0
cc_111 N_A_N_c_91_n N_A_27_51#_c_134_n 0.0131389f $X=0.725 $Y=1.55 $X2=0 $Y2=0
cc_112 N_A_N_M1010_g N_VPWR_c_353_n 0.00645675f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_113 N_A_N_M1013_g N_VGND_c_504_n 0.0108071f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_114 N_A_N_M1013_g N_VGND_c_506_n 0.00346638f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_115 N_A_N_M1013_g N_VGND_c_509_n 0.00507428f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_116 N_A_N_M1013_g N_A_217_65#_c_561_n 0.00465426f $X=0.475 $Y=0.465 $X2=0
+ $Y2=0
cc_117 N_A_27_51#_M1009_g N_B_M1000_g 0.0223864f $X=1.855 $Y=0.745 $X2=0 $Y2=0
cc_118 N_A_27_51#_M1015_g N_B_M1001_g 0.0223864f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_27_51#_M1003_g B 3.3994e-19 $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_27_51#_M1015_g B 0.00243063f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_27_51#_c_132_n B 0.0193004f $X=1.59 $Y=1.51 $X2=0 $Y2=0
cc_122 N_A_27_51#_c_134_n B 0.00879411f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_123 N_A_27_51#_c_134_n N_B_c_210_n 0.0223864f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_124 N_A_27_51#_M1003_g N_VPWR_c_353_n 0.00939649f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_27_51#_c_131_n N_VPWR_c_353_n 0.00604258f $X=0.695 $Y=1.895 $X2=0
+ $Y2=0
cc_126 N_A_27_51#_c_132_n N_VPWR_c_353_n 0.0316172f $X=1.59 $Y=1.51 $X2=0 $Y2=0
cc_127 N_A_27_51#_c_138_n N_VPWR_c_353_n 0.026061f $X=0.695 $Y=2.06 $X2=0 $Y2=0
cc_128 N_A_27_51#_c_134_n N_VPWR_c_353_n 0.00601434f $X=1.855 $Y=1.51 $X2=0
+ $Y2=0
cc_129 N_A_27_51#_M1015_g N_VPWR_c_354_n 0.0027678f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_27_51#_M1003_g N_VPWR_c_359_n 0.00585385f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_27_51#_M1015_g N_VPWR_c_359_n 0.00585385f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_27_51#_M1003_g N_VPWR_c_352_n 0.0118358f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_27_51#_M1015_g N_VPWR_c_352_n 0.0107074f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_27_51#_M1002_g N_Y_c_429_n 0.0054303f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_135 N_A_27_51#_M1009_g N_Y_c_429_n 0.00675298f $X=1.855 $Y=0.745 $X2=0 $Y2=0
cc_136 N_A_27_51#_c_132_n N_Y_c_431_n 0.0112811f $X=1.59 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A_27_51#_c_134_n N_Y_c_431_n 0.00227722f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_138 N_A_27_51#_M1015_g N_Y_c_433_n 0.0154651f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_27_51#_M1009_g N_Y_c_425_n 0.0112929f $X=1.855 $Y=0.745 $X2=0 $Y2=0
cc_140 N_A_27_51#_M1002_g N_Y_c_426_n 0.00529936f $X=1.425 $Y=0.745 $X2=0 $Y2=0
cc_141 N_A_27_51#_M1009_g N_Y_c_426_n 0.00201986f $X=1.855 $Y=0.745 $X2=0 $Y2=0
cc_142 N_A_27_51#_c_132_n N_Y_c_426_n 0.0228472f $X=1.59 $Y=1.51 $X2=0 $Y2=0
cc_143 N_A_27_51#_c_134_n N_Y_c_426_n 0.00252809f $X=1.855 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A_27_51#_M1002_g N_VGND_c_504_n 0.00149641f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_145 N_A_27_51#_c_128_n N_VGND_c_504_n 0.0192074f $X=0.605 $Y=0.78 $X2=0 $Y2=0
cc_146 N_A_27_51#_c_127_n N_VGND_c_506_n 0.0100784f $X=0.26 $Y=0.465 $X2=0 $Y2=0
cc_147 N_A_27_51#_c_128_n N_VGND_c_506_n 0.00265317f $X=0.605 $Y=0.78 $X2=0
+ $Y2=0
cc_148 N_A_27_51#_M1002_g N_VGND_c_507_n 0.00302501f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_149 N_A_27_51#_M1009_g N_VGND_c_507_n 0.00302501f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_150 N_A_27_51#_M1002_g N_VGND_c_509_n 0.0048466f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_151 N_A_27_51#_M1009_g N_VGND_c_509_n 0.00441786f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_152 N_A_27_51#_c_127_n N_VGND_c_509_n 0.00709944f $X=0.26 $Y=0.465 $X2=0
+ $Y2=0
cc_153 N_A_27_51#_c_128_n N_VGND_c_509_n 0.00544199f $X=0.605 $Y=0.78 $X2=0
+ $Y2=0
cc_154 N_A_27_51#_M1002_g N_A_217_65#_c_561_n 0.00354524f $X=1.425 $Y=0.745
+ $X2=0 $Y2=0
cc_155 N_A_27_51#_c_128_n N_A_217_65#_c_561_n 0.0109173f $X=0.605 $Y=0.78 $X2=0
+ $Y2=0
cc_156 N_A_27_51#_c_130_n N_A_217_65#_c_561_n 0.0185751f $X=0.695 $Y=1.415 $X2=0
+ $Y2=0
cc_157 N_A_27_51#_c_132_n N_A_217_65#_c_561_n 0.0171024f $X=1.59 $Y=1.51 $X2=0
+ $Y2=0
cc_158 N_A_27_51#_c_134_n N_A_217_65#_c_561_n 0.00538122f $X=1.855 $Y=1.51 $X2=0
+ $Y2=0
cc_159 N_A_27_51#_M1002_g N_A_217_65#_c_562_n 0.0125492f $X=1.425 $Y=0.745 $X2=0
+ $Y2=0
cc_160 N_A_27_51#_M1009_g N_A_217_65#_c_562_n 0.0115502f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_161 N_B_c_210_n C 2.91423e-19 $X=2.795 $Y=1.51 $X2=0 $Y2=0
cc_162 N_B_M1001_g N_VPWR_c_354_n 0.00272526f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B_M1001_g N_VPWR_c_360_n 0.00585385f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_164 N_B_M1008_g N_VPWR_c_360_n 0.00487821f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B_M1001_g N_VPWR_c_365_n 6.94391e-19 $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_166 N_B_M1008_g N_VPWR_c_365_n 0.0184066f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_167 N_B_M1001_g N_VPWR_c_352_n 0.0107333f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_168 N_B_M1008_g N_VPWR_c_352_n 0.00827319f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_169 N_B_M1000_g N_Y_c_429_n 5.43231e-19 $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_170 N_B_M1001_g N_Y_c_433_n 0.013326f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_171 B N_Y_c_433_n 0.0346419f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_172 N_B_M1000_g N_Y_c_425_n 0.0112174f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_173 N_B_M1016_g N_Y_c_425_n 0.0135334f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_174 B N_Y_c_425_n 0.0618156f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_175 N_B_c_210_n N_Y_c_425_n 0.0043953f $X=2.795 $Y=1.51 $X2=0 $Y2=0
cc_176 N_B_M1000_g N_Y_c_427_n 4.65827e-19 $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_177 N_B_M1016_g N_Y_c_427_n 0.00383612f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_178 B N_Y_c_427_n 0.0274471f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B_c_210_n N_Y_c_427_n 0.0206198f $X=2.795 $Y=1.51 $X2=0 $Y2=0
cc_180 B Y 0.0177466f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_181 N_B_c_210_n Y 7.18291e-19 $X=2.795 $Y=1.51 $X2=0 $Y2=0
cc_182 N_B_M1008_g N_Y_c_452_n 0.0175583f $X=2.795 $Y=2.465 $X2=0 $Y2=0
cc_183 B N_Y_c_452_n 0.00292845f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_184 N_B_M1000_g N_VGND_c_507_n 0.00355797f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_185 N_B_M1016_g N_VGND_c_507_n 0.00302901f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_186 N_B_M1000_g N_VGND_c_509_n 0.00517046f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_187 N_B_M1016_g N_VGND_c_509_n 0.0049033f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_188 N_B_M1000_g N_A_217_65#_c_562_n 0.00285294f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_189 N_B_M1000_g N_A_217_65#_c_574_n 0.00463146f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_190 N_B_M1016_g N_A_217_65#_c_574_n 4.19477e-19 $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_191 N_B_M1000_g N_A_217_65#_c_576_n 7.54017e-19 $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_192 N_B_M1000_g N_A_217_65#_c_577_n 0.00938505f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_193 N_B_M1016_g N_A_217_65#_c_577_n 0.00968245f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_194 N_B_M1016_g N_A_486_65#_c_602_n 0.009647f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_195 N_B_M1000_g N_A_486_65#_c_603_n 0.00179081f $X=2.355 $Y=0.745 $X2=0 $Y2=0
cc_196 N_B_M1016_g N_A_486_65#_c_603_n 0.00788052f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_197 N_B_M1016_g N_A_697_69#_c_630_n 0.00435451f $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_198 N_B_M1016_g N_A_697_69#_c_632_n 7.58088e-19 $X=2.855 $Y=0.745 $X2=0 $Y2=0
cc_199 N_C_M1012_g N_D_M1005_g 0.0242574f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_200 N_C_M1011_g N_D_M1007_g 0.0242574f $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_201 C N_D_M1007_g 0.00193578f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_202 C D 0.0277542f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_203 C N_D_c_316_n 0.007505f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_204 N_C_c_263_n N_D_c_316_n 0.0242574f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_205 N_C_M1004_g N_VPWR_c_355_n 6.80491e-19 $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_206 N_C_M1011_g N_VPWR_c_355_n 0.0145152f $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_207 N_C_M1004_g N_VPWR_c_361_n 0.00487821f $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_208 N_C_M1011_g N_VPWR_c_361_n 0.00486043f $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_209 N_C_M1004_g N_VPWR_c_365_n 0.0182894f $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_210 N_C_M1011_g N_VPWR_c_365_n 6.86512e-19 $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_211 N_C_M1004_g N_VPWR_c_352_n 0.00824731f $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_212 N_C_M1011_g N_VPWR_c_352_n 0.00824727f $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_213 N_C_M1006_g N_Y_c_425_n 6.23791e-19 $X=3.905 $Y=0.765 $X2=0 $Y2=0
cc_214 N_C_M1006_g N_Y_c_427_n 0.00211945f $X=3.905 $Y=0.765 $X2=0 $Y2=0
cc_215 N_C_M1004_g N_Y_c_427_n 0.00417931f $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_216 C N_Y_c_427_n 0.0284456f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_217 N_C_c_263_n N_Y_c_427_n 0.00329977f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_218 N_C_M1011_g N_Y_c_459_n 0.0122129f $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_219 C N_Y_c_459_n 0.0319767f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_220 C Y 0.0153757f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_221 N_C_c_263_n Y 6.52992e-19 $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_222 N_C_M1004_g N_Y_c_463_n 0.0155656f $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_223 C N_Y_c_463_n 0.0455852f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_224 N_C_c_263_n N_Y_c_463_n 4.14878e-19 $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_225 N_C_M1012_g N_VGND_c_505_n 6.40069e-19 $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_226 N_C_M1006_g N_VGND_c_507_n 0.00291444f $X=3.905 $Y=0.765 $X2=0 $Y2=0
cc_227 N_C_M1012_g N_VGND_c_507_n 0.00450424f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_228 N_C_M1006_g N_VGND_c_509_n 0.00428623f $X=3.905 $Y=0.765 $X2=0 $Y2=0
cc_229 N_C_M1012_g N_VGND_c_509_n 0.00862457f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_230 N_C_M1006_g N_A_486_65#_c_602_n 0.0118679f $X=3.905 $Y=0.765 $X2=0 $Y2=0
cc_231 N_C_M1012_g N_A_486_65#_c_602_n 0.00345965f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_232 N_C_M1006_g N_A_486_65#_c_609_n 0.0111491f $X=3.905 $Y=0.765 $X2=0 $Y2=0
cc_233 N_C_M1012_g N_A_486_65#_c_609_n 0.00527422f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_234 N_C_M1006_g N_A_697_69#_c_631_n 0.0139229f $X=3.905 $Y=0.765 $X2=0 $Y2=0
cc_235 N_C_M1012_g N_A_697_69#_c_631_n 0.013073f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_236 C N_A_697_69#_c_631_n 0.0500356f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_237 N_C_c_263_n N_A_697_69#_c_631_n 0.00381774f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_238 C N_A_697_69#_c_632_n 0.0289474f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_239 N_C_c_263_n N_A_697_69#_c_632_n 8.9626e-19 $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_240 N_C_M1012_g N_A_697_69#_c_633_n 8.29132e-19 $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_241 C N_A_697_69#_c_634_n 0.0045171f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_242 C N_A_697_69#_c_636_n 0.017673f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_243 N_D_M1007_g N_VPWR_c_355_n 0.0145152f $X=4.765 $Y=2.465 $X2=0 $Y2=0
cc_244 N_D_M1017_g N_VPWR_c_355_n 6.80491e-19 $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_245 N_D_M1007_g N_VPWR_c_357_n 7.28867e-19 $X=4.765 $Y=2.465 $X2=0 $Y2=0
cc_246 N_D_M1017_g N_VPWR_c_357_n 0.0203776f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_247 D N_VPWR_c_357_n 0.025707f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_248 N_D_M1007_g N_VPWR_c_362_n 0.00486043f $X=4.765 $Y=2.465 $X2=0 $Y2=0
cc_249 N_D_M1017_g N_VPWR_c_362_n 0.00486043f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_250 N_D_M1007_g N_VPWR_c_352_n 0.00824727f $X=4.765 $Y=2.465 $X2=0 $Y2=0
cc_251 N_D_M1017_g N_VPWR_c_352_n 0.00824727f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_252 N_D_M1007_g N_Y_c_459_n 0.0140388f $X=4.765 $Y=2.465 $X2=0 $Y2=0
cc_253 D N_Y_c_467_n 0.0153757f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_254 N_D_c_316_n N_Y_c_467_n 6.52992e-19 $X=5.205 $Y=1.51 $X2=0 $Y2=0
cc_255 N_D_M1005_g N_VGND_c_505_n 0.00960578f $X=4.765 $Y=0.765 $X2=0 $Y2=0
cc_256 N_D_M1014_g N_VGND_c_505_n 0.012812f $X=5.205 $Y=0.765 $X2=0 $Y2=0
cc_257 N_D_M1005_g N_VGND_c_507_n 0.00432557f $X=4.765 $Y=0.765 $X2=0 $Y2=0
cc_258 N_D_M1014_g N_VGND_c_508_n 0.00400407f $X=5.205 $Y=0.765 $X2=0 $Y2=0
cc_259 N_D_M1005_g N_VGND_c_509_n 0.00836275f $X=4.765 $Y=0.765 $X2=0 $Y2=0
cc_260 N_D_M1014_g N_VGND_c_509_n 0.0079758f $X=5.205 $Y=0.765 $X2=0 $Y2=0
cc_261 N_D_M1005_g N_A_486_65#_c_602_n 2.33832e-19 $X=4.765 $Y=0.765 $X2=0 $Y2=0
cc_262 N_D_M1005_g N_A_697_69#_c_633_n 8.46957e-19 $X=4.765 $Y=0.765 $X2=0 $Y2=0
cc_263 N_D_M1005_g N_A_697_69#_c_634_n 0.0153249f $X=4.765 $Y=0.765 $X2=0 $Y2=0
cc_264 N_D_M1014_g N_A_697_69#_c_634_n 0.0137346f $X=5.205 $Y=0.765 $X2=0 $Y2=0
cc_265 D N_A_697_69#_c_634_n 0.0573601f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_266 N_D_c_316_n N_A_697_69#_c_634_n 0.00275417f $X=5.205 $Y=1.51 $X2=0 $Y2=0
cc_267 N_D_M1014_g N_A_697_69#_c_635_n 0.00354659f $X=5.205 $Y=0.765 $X2=0 $Y2=0
cc_268 N_VPWR_c_352_n N_Y_M1003_d 0.0027574f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_c_352_n N_Y_M1001_d 0.00422932f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_270 N_VPWR_c_352_n N_Y_M1004_s 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_271 N_VPWR_c_352_n N_Y_M1007_s 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_359_n N_Y_c_473_n 0.0151136f $X=1.94 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_c_352_n N_Y_c_473_n 0.0102248f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_274 N_VPWR_M1015_s N_Y_c_433_n 0.00502357f $X=1.93 $Y=1.835 $X2=0 $Y2=0
cc_275 N_VPWR_c_354_n N_Y_c_433_n 0.0192006f $X=2.105 $Y=2.385 $X2=0 $Y2=0
cc_276 N_VPWR_M1008_s N_Y_c_427_n 0.0022953f $X=2.87 $Y=1.835 $X2=0 $Y2=0
cc_277 N_VPWR_M1011_d N_Y_c_459_n 0.00353353f $X=4.41 $Y=1.835 $X2=0 $Y2=0
cc_278 N_VPWR_c_355_n N_Y_c_459_n 0.0170777f $X=4.55 $Y=2.39 $X2=0 $Y2=0
cc_279 N_VPWR_c_362_n N_Y_c_480_n 0.0124525f $X=5.245 $Y=3.33 $X2=0 $Y2=0
cc_280 N_VPWR_c_352_n N_Y_c_480_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_281 N_VPWR_M1008_s Y 0.00500257f $X=2.87 $Y=1.835 $X2=0 $Y2=0
cc_282 N_VPWR_c_365_n Y 0.0259215f $X=3.01 $Y=2.375 $X2=0 $Y2=0
cc_283 N_VPWR_c_365_n N_Y_c_452_n 0.00180677f $X=3.01 $Y=2.375 $X2=0 $Y2=0
cc_284 N_VPWR_M1008_s N_Y_c_463_n 0.0213709f $X=2.87 $Y=1.835 $X2=0 $Y2=0
cc_285 N_VPWR_c_365_n N_Y_c_463_n 0.0476696f $X=3.01 $Y=2.375 $X2=0 $Y2=0
cc_286 N_VPWR_c_360_n N_Y_c_487_n 0.0143974f $X=2.845 $Y=3.33 $X2=0 $Y2=0
cc_287 N_VPWR_c_352_n N_Y_c_487_n 0.0090585f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_288 N_VPWR_c_361_n N_Y_c_489_n 0.0124525f $X=4.385 $Y=3.33 $X2=0 $Y2=0
cc_289 N_VPWR_c_352_n N_Y_c_489_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_290 N_Y_c_425_n N_A_217_65#_M1009_d 0.00250873f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_291 N_Y_c_425_n N_A_217_65#_M1016_s 0.00273087f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_292 N_Y_c_426_n N_A_217_65#_c_561_n 0.00539933f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_293 N_Y_M1002_s N_A_217_65#_c_562_n 0.00176461f $X=1.5 $Y=0.325 $X2=0 $Y2=0
cc_294 N_Y_c_429_n N_A_217_65#_c_562_n 0.0159249f $X=1.64 $Y=0.68 $X2=0 $Y2=0
cc_295 N_Y_c_425_n N_A_217_65#_c_562_n 0.00275981f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_296 N_Y_c_425_n N_A_217_65#_c_576_n 0.0209853f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_297 N_Y_c_425_n N_A_217_65#_c_577_n 0.0552053f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_298 N_Y_c_425_n N_A_486_65#_M1000_d 0.00251484f $X=2.905 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_299 N_Y_c_425_n N_A_697_69#_c_630_n 6.81585e-19 $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_300 N_Y_c_425_n N_A_697_69#_c_632_n 0.0121097f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_301 N_Y_c_427_n N_A_697_69#_c_632_n 6.78718e-19 $X=3.06 $Y=1.92 $X2=0 $Y2=0
cc_302 N_Y_c_459_n N_A_697_69#_c_634_n 0.00335436f $X=4.885 $Y=2.005 $X2=0 $Y2=0
cc_303 N_VGND_c_504_n N_A_217_65#_c_561_n 0.00752662f $X=0.69 $Y=0.42 $X2=0
+ $Y2=0
cc_304 N_VGND_c_507_n N_A_217_65#_c_562_n 0.0657172f $X=4.825 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_509_n N_A_217_65#_c_562_n 0.0365173f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_504_n N_A_217_65#_c_563_n 0.0139f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_307 N_VGND_c_507_n N_A_217_65#_c_563_n 0.0186386f $X=4.825 $Y=0 $X2=0 $Y2=0
cc_308 N_VGND_c_509_n N_A_217_65#_c_563_n 0.0101082f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_507_n N_A_217_65#_c_577_n 0.00204091f $X=4.825 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_509_n N_A_217_65#_c_577_n 0.00491956f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_505_n N_A_486_65#_c_602_n 0.00215867f $X=4.99 $Y=0.47 $X2=0
+ $Y2=0
cc_312 N_VGND_c_507_n N_A_486_65#_c_602_n 0.0967555f $X=4.825 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_509_n N_A_486_65#_c_602_n 0.0546872f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_507_n N_A_486_65#_c_603_n 0.0220628f $X=4.825 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_509_n N_A_486_65#_c_603_n 0.0123875f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_505_n N_A_697_69#_c_633_n 0.0228709f $X=4.99 $Y=0.47 $X2=0 $Y2=0
cc_317 N_VGND_c_507_n N_A_697_69#_c_633_n 0.00981731f $X=4.825 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_c_509_n N_A_697_69#_c_633_n 0.00742088f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_M1005_d N_A_697_69#_c_634_n 0.00187091f $X=4.84 $Y=0.345 $X2=0
+ $Y2=0
cc_320 N_VGND_c_505_n N_A_697_69#_c_634_n 0.0171295f $X=4.99 $Y=0.47 $X2=0 $Y2=0
cc_321 N_VGND_c_505_n N_A_697_69#_c_635_n 0.0229093f $X=4.99 $Y=0.47 $X2=0 $Y2=0
cc_322 N_VGND_c_508_n N_A_697_69#_c_635_n 0.0137839f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_509_n N_A_697_69#_c_635_n 0.0104192f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_324 N_A_217_65#_c_577_n N_A_486_65#_M1000_d 0.00473585f $X=2.975 $Y=0.775
+ $X2=-0.19 $Y2=-0.245
cc_325 N_A_217_65#_M1016_s N_A_486_65#_c_602_n 0.00294574f $X=2.93 $Y=0.325
+ $X2=0 $Y2=0
cc_326 N_A_217_65#_c_564_n N_A_486_65#_c_602_n 0.0141492f $X=3.07 $Y=0.81 $X2=0
+ $Y2=0
cc_327 N_A_217_65#_c_577_n N_A_486_65#_c_602_n 0.00476109f $X=2.975 $Y=0.775
+ $X2=0 $Y2=0
cc_328 N_A_217_65#_c_562_n N_A_486_65#_c_603_n 0.0100439f $X=1.975 $Y=0.34 $X2=0
+ $Y2=0
cc_329 N_A_217_65#_c_577_n N_A_486_65#_c_603_n 0.0190318f $X=2.975 $Y=0.775
+ $X2=0 $Y2=0
cc_330 N_A_217_65#_c_564_n N_A_697_69#_c_630_n 0.0192376f $X=3.07 $Y=0.81 $X2=0
+ $Y2=0
cc_331 N_A_486_65#_c_602_n N_A_697_69#_M1006_s 0.00378299f $X=3.955 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_332 N_A_486_65#_c_602_n N_A_697_69#_c_630_n 0.0249442f $X=3.955 $Y=0.34 $X2=0
+ $Y2=0
cc_333 N_A_486_65#_M1006_d N_A_697_69#_c_631_n 0.00176461f $X=3.98 $Y=0.345
+ $X2=0 $Y2=0
cc_334 N_A_486_65#_c_602_n N_A_697_69#_c_631_n 0.00272017f $X=3.955 $Y=0.34
+ $X2=0 $Y2=0
cc_335 N_A_486_65#_c_609_n N_A_697_69#_c_631_n 0.017036f $X=4.12 $Y=0.47 $X2=0
+ $Y2=0
cc_336 N_A_486_65#_c_602_n N_A_697_69#_c_633_n 0.00494821f $X=3.955 $Y=0.34
+ $X2=0 $Y2=0
