* File: sky130_fd_sc_lp__a31oi_0.pex.spice
* Created: Fri Aug 28 09:59:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31OI_0%A3 2 5 7 9 13 14 17 19 20 21 26
c41 26 0 3.46425e-19 $X=0.27 $Y=1.12
c42 5 0 1.56626e-19 $X=0.475 $Y=2.685
c43 2 0 1.10673e-19 $X=0.36 $Y=2.065
r44 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r45 20 21 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r46 20 27 5.45074 $w=3.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.12
r47 19 27 6.07369 $w=3.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.27 $Y=0.925
+ $X2=0.27 $Y2=1.12
r48 15 17 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=0.36 $Y=2.14
+ $X2=0.475 $Y2=2.14
r49 13 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.12
r50 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.625
r51 7 26 60.5302 $w=2.15e-07 $l=4.71036e-07 $layer=POLY_cond $X=0.54 $Y=0.765
+ $X2=0.27 $Y2=1.12
r52 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.765 $X2=0.54
+ $Y2=0.445
r53 3 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.215
+ $X2=0.475 $Y2=2.14
r54 3 5 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.475 $Y=2.215 $X2=0.475
+ $Y2=2.685
r55 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.065
+ $X2=0.36 $Y2=2.14
r56 2 14 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.36 $Y=2.065
+ $X2=0.36 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_0%A2 3 7 11 12 13 14 15 16 22
c42 13 0 1.10673e-19 $X=0.72 $Y=0.555
c43 11 0 1.4009e-19 $X=0.84 $Y=1.66
c44 3 0 2.97244e-19 $X=0.905 $Y=2.685
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.32 $X2=0.84 $Y2=1.32
r46 16 23 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=0.775 $Y=1.665
+ $X2=0.775 $Y2=1.32
r47 15 23 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=0.775 $Y=1.295
+ $X2=0.775 $Y2=1.32
r48 14 15 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.775 $Y=0.925
+ $X2=0.775 $Y2=1.295
r49 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.775 $Y=0.555
+ $X2=0.775 $Y2=0.925
r50 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.84 $Y=1.66
+ $X2=0.84 $Y2=1.32
r51 11 12 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.66
+ $X2=0.84 $Y2=1.825
r52 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.155
+ $X2=0.84 $Y2=1.32
r53 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.93 $Y=0.445
+ $X2=0.93 $Y2=1.155
r54 3 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.905 $Y=2.685
+ $X2=0.905 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_0%A1 3 7 11 12 13 14 15 20
c40 12 0 1.99439e-20 $X=1.41 $Y=1.51
c41 7 0 1.5634e-19 $X=1.335 $Y=2.685
r42 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.41
+ $Y=1.005 $X2=1.41 $Y2=1.005
r43 14 15 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.3 $Y=1.295 $X2=1.3
+ $Y2=1.665
r44 14 21 8.15143 $w=4.08e-07 $l=2.9e-07 $layer=LI1_cond $X=1.3 $Y=1.295 $X2=1.3
+ $Y2=1.005
r45 13 21 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=1.3 $Y=0.925 $X2=1.3
+ $Y2=1.005
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.41 $Y=1.345
+ $X2=1.41 $Y2=1.005
r47 11 12 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.345
+ $X2=1.41 $Y2=1.51
r48 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.84
+ $X2=1.41 $Y2=1.005
r49 7 12 602.5 $w=1.5e-07 $l=1.175e-06 $layer=POLY_cond $X=1.335 $Y=2.685
+ $X2=1.335 $Y2=1.51
r50 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.32 $Y=0.445
+ $X2=1.32 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_0%B1 1 3 7 9 10 11
c30 3 0 1.54676e-19 $X=1.765 $Y=2.685
r31 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.11
+ $Y=1.12 $X2=2.11 $Y2=1.12
r32 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.165 $Y=1.295
+ $X2=2.165 $Y2=1.665
r33 10 17 6.72258 $w=2.98e-07 $l=1.75e-07 $layer=LI1_cond $X=2.165 $Y=1.295
+ $X2=2.165 $Y2=1.12
r34 9 17 7.49088 $w=2.98e-07 $l=1.95e-07 $layer=LI1_cond $X=2.165 $Y=0.925
+ $X2=2.165 $Y2=1.12
r35 5 16 39.3769 $w=3.89e-07 $l=2.05925e-07 $layer=POLY_cond $X=1.89 $Y=0.955
+ $X2=1.982 $Y2=1.12
r36 5 7 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.89 $Y=0.955 $X2=1.89
+ $Y2=0.445
r37 1 16 115.58 $w=3.89e-07 $l=8.8185e-07 $layer=POLY_cond $X=1.765 $Y=1.9
+ $X2=1.982 $Y2=1.12
r38 1 3 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.765 $Y=1.9
+ $X2=1.765 $Y2=2.685
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_0%VPWR 1 2 8 10 11 12 15 17 24 25
c48 11 0 1.99439e-20 $X=0.99 $Y=2.08
c49 10 0 1.40618e-19 $X=0.26 $Y=2.51
r50 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 22 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 21 24 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 19 28 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r56 19 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 17 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 17 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 13 15 17.9515 $w=2.58e-07 $l=4.05e-07 $layer=LI1_cond $X=1.12 $Y=2.165
+ $X2=1.12 $Y2=2.57
r60 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.99 $Y=2.08
+ $X2=1.12 $Y2=2.165
r61 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.99 $Y=2.08 $X2=0.39
+ $Y2=2.08
r62 8 28 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.195 $Y2=3.33
r63 8 10 28.7134 $w=2.93e-07 $l=7.35e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.242 $Y2=2.51
r64 7 12 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.242 $Y=2.165
+ $X2=0.39 $Y2=2.08
r65 7 10 13.4777 $w=2.93e-07 $l=3.45e-07 $layer=LI1_cond $X=0.242 $Y=2.165
+ $X2=0.242 $Y2=2.51
r66 2 15 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.365 $X2=1.12 $Y2=2.57
r67 1 10 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.365 $X2=0.26 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_0%A_110_473# 1 2 9 11 12 15
c22 15 0 3.11016e-19 $X=1.55 $Y=2.51
c23 9 0 3.13252e-19 $X=0.69 $Y=2.51
r24 13 15 17.8516 $w=2.53e-07 $l=3.95e-07 $layer=LI1_cond $X=1.547 $Y=2.905
+ $X2=1.547 $Y2=2.51
r25 11 13 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.42 $Y=2.99
+ $X2=1.547 $Y2=2.905
r26 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.42 $Y=2.99 $X2=0.82
+ $Y2=2.99
r27 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.69 $Y=2.905
+ $X2=0.82 $Y2=2.99
r28 7 9 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=0.69 $Y=2.905
+ $X2=0.69 $Y2=2.51
r29 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.365 $X2=1.55 $Y2=2.51
r30 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.365 $X2=0.69 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_0%Y 1 2 12 14 15 16 29
r32 16 24 6.74385 $w=4.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.08 $Y=2.775
+ $X2=2.08 $Y2=2.51
r33 15 24 2.67209 $w=4.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.08 $Y=2.405
+ $X2=2.08 $Y2=2.51
r34 15 31 5.85315 $w=4.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.08 $Y=2.405
+ $X2=2.08 $Y2=2.175
r35 14 31 3.48349 $w=6.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.995 $Y=2.035
+ $X2=1.995 $Y2=2.175
r36 14 29 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=2.035
+ $X2=1.995 $Y2=1.95
r37 10 12 5.16019 $w=3.33e-07 $l=1.5e-07 $layer=LI1_cond $X=1.61 $Y=0.447
+ $X2=1.76 $Y2=0.447
r38 7 12 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.76 $Y=0.615
+ $X2=1.76 $Y2=0.447
r39 7 29 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=1.76 $Y=0.615
+ $X2=1.76 $Y2=1.95
r40 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.365 $X2=1.98 $Y2=2.51
r41 1 10 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=1.395
+ $Y=0.235 $X2=1.61 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_0%VGND 1 2 7 9 11 13 15 17 30
c31 30 0 1.96469e-19 $X=2.16 $Y=0
c32 17 0 1.49956e-19 $X=2.015 $Y=0
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r36 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r37 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r38 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r39 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 18 26 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r41 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r42 17 29 4.29523 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=2.207
+ $Y2=0
r43 17 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=1.68
+ $Y2=0
r44 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r45 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r46 11 29 3.06482 $w=2.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.207 $Y2=0
r47 11 13 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0.445
r48 7 26 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r49 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.29 $Y2=0.43
r50 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.235 $X2=2.105 $Y2=0.445
r51 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.2 $Y=0.235
+ $X2=0.325 $Y2=0.43
.ends

