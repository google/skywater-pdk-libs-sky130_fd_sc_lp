* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtn_lp D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 a_744_415# a_264_415# a_901_415# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_114_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_27_47# a_712_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_898_47# a_949_335# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_47# D a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND GATE_N a_272_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1222_57# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_949_335# a_1380_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_949_335# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_399_415# a_264_415# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VPWR a_744_415# a_949_335# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_949_335# a_744_415# a_1222_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_949_335# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_712_47# a_264_415# a_744_415# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_27_47# a_646_415# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_272_47# GATE_N a_264_415# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR GATE_N a_264_415# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_646_415# a_399_415# a_744_415# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X18 a_1380_57# a_949_335# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_901_415# a_949_335# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 a_399_415# a_264_415# a_554_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_27_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_554_47# a_264_415# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_744_415# a_399_415# a_898_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
