* File: sky130_fd_sc_lp__nand4b_m.pex.spice
* Created: Wed Sep  2 10:06:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4B_M%A_N 3 7 11 12 13 14 15 16 17 24
r42 24 26 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.642 $Y=1.005
+ $X2=0.642 $Y2=0.84
r43 16 17 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.685 $Y=2.035
+ $X2=0.685 $Y2=2.405
r44 15 16 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.685 $Y=1.665
+ $X2=0.685 $Y2=2.035
r45 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.685 $Y=1.295
+ $X2=0.685 $Y2=1.665
r46 13 14 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.685 $Y=0.925
+ $X2=0.685 $Y2=1.295
r47 13 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.65
+ $Y=1.005 $X2=0.65 $Y2=1.005
r48 11 12 43.8566 $w=3.45e-07 $l=1.5e-07 $layer=POLY_cond $X=0.627 $Y=1.36
+ $X2=0.627 $Y2=1.51
r49 9 24 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=0.642 $Y=1.012
+ $X2=0.642 $Y2=1.005
r50 9 11 58.206 $w=3.45e-07 $l=3.48e-07 $layer=POLY_cond $X=0.642 $Y=1.012
+ $X2=0.642 $Y2=1.36
r51 7 26 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.545 $Y=0.47
+ $X2=0.545 $Y2=0.84
r52 3 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.515 $Y=2.17
+ $X2=0.515 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_M%D 3 8 10 11 12 13 14 15 16 17 22
c48 22 0 2.60315e-20 $X=1.19 $Y=0.955
r49 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=0.925
+ $X2=1.19 $Y2=1.295
r50 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.19
+ $Y=0.955 $X2=1.19 $Y2=0.955
r51 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=0.555
+ $X2=1.19 $Y2=0.925
r52 13 14 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=1.282 $Y=1.7
+ $X2=1.282 $Y2=1.85
r53 12 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.28 $Y=1.46
+ $X2=1.28 $Y2=1.7
r54 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.19 $Y=1.295
+ $X2=1.19 $Y2=0.955
r55 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.295
+ $X2=1.19 $Y2=1.46
r56 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=0.79
+ $X2=1.19 $Y2=0.955
r57 8 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.285 $Y=2.17
+ $X2=1.285 $Y2=1.85
r58 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.28 $Y=0.47 $X2=1.28
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_M%C 3 6 9 10 11 12 13 14 19
c42 19 0 2.60315e-20 $X=1.73 $Y=0.955
r43 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.73 $Y=0.925
+ $X2=1.73 $Y2=1.295
r44 13 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=0.955 $X2=1.73 $Y2=0.955
r45 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.73 $Y=0.555
+ $X2=1.73 $Y2=0.925
r46 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=0.955
r47 10 11 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.46
r48 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.79
+ $X2=1.73 $Y2=0.955
r49 6 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.715 $Y=2.17
+ $X2=1.715 $Y2=1.46
r50 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.64 $Y=0.47 $X2=1.64
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_M%B 3 6 9 10 12 13 14 15 16 17 22
c44 22 0 2.60315e-20 $X=2.27 $Y=0.955
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27
+ $Y=0.955 $X2=2.27 $Y2=0.955
r46 17 23 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.255 $Y=1.295
+ $X2=2.255 $Y2=0.955
r47 16 23 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=2.255 $Y=0.925
+ $X2=2.255 $Y2=0.955
r48 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.255 $Y=0.555
+ $X2=2.255 $Y2=0.925
r49 13 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.27 $Y=1.295
+ $X2=2.27 $Y2=0.955
r50 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.295
+ $X2=2.27 $Y2=1.46
r51 12 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=0.79
+ $X2=2.27 $Y2=0.955
r52 9 10 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=2.162 $Y=1.7
+ $X2=2.162 $Y2=1.85
r53 9 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.18 $Y=1.7 $X2=2.18
+ $Y2=1.46
r54 6 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.18 $Y=0.47 $X2=2.18
+ $Y2=0.79
r55 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.145 $Y=2.17
+ $X2=2.145 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_M%A_35_392# 1 2 7 12 15 19 24 26 32 33
r55 33 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.72 $Y=2.885 $X2=0.72
+ $Y2=2.975
r56 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=2.885 $X2=0.72 $Y2=2.885
r57 29 32 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.275 $Y=2.885
+ $X2=0.72 $Y2=2.885
r58 26 28 4.95036 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.33 $Y=0.535
+ $X2=0.33 $Y2=0.64
r59 24 28 76.7422 $w=2.18e-07 $l=1.465e-06 $layer=LI1_cond $X=0.275 $Y=2.105
+ $X2=0.275 $Y2=0.64
r60 22 29 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=2.72
+ $X2=0.275 $Y2=2.885
r61 22 24 32.216 $w=2.18e-07 $l=6.15e-07 $layer=LI1_cond $X=0.275 $Y=2.72
+ $X2=0.275 $Y2=2.105
r62 17 19 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.575 $Y=1.775
+ $X2=2.72 $Y2=1.775
r63 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.72 $Y=1.7 $X2=2.72
+ $Y2=1.775
r64 13 15 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=2.72 $Y=1.7
+ $X2=2.72 $Y2=0.47
r65 10 12 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.575 $Y=2.9
+ $X2=2.575 $Y2=2.17
r66 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.575 $Y=1.85
+ $X2=2.575 $Y2=1.775
r67 9 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.575 $Y=1.85
+ $X2=2.575 $Y2=2.17
r68 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.885 $Y=2.975
+ $X2=0.72 $Y2=2.975
r69 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.5 $Y=2.975
+ $X2=2.575 $Y2=2.9
r70 7 8 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=2.5 $Y=2.975
+ $X2=0.885 $Y2=2.975
r71 2 24 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.96 $X2=0.3 $Y2=2.105
r72 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.26 $X2=0.33 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_M%VPWR 1 2 3 12 16 20 23 24 26 27 29 30 31 44
+ 45
r36 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 31 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 31 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 29 41 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 29 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.705 $Y=3.33 $X2=2.8
+ $Y2=3.33
r45 28 44 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 28 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.895 $Y=3.33 $X2=2.8
+ $Y2=3.33
r47 26 38 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.93 $Y2=3.33
r49 25 41 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.93 $Y2=3.33
r51 23 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.07 $Y2=3.33
r53 22 38 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.07 $Y2=3.33
r55 18 30 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=3.245 $X2=2.8
+ $Y2=3.33
r56 18 20 58.9569 $w=1.88e-07 $l=1.01e-06 $layer=LI1_cond $X=2.8 $Y=3.245
+ $X2=2.8 $Y2=2.235
r57 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r58 14 16 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.235
r59 10 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r60 10 12 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.235
r61 3 20 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.96 $X2=2.79 $Y2=2.235
r62 2 16 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.96 $X2=1.93 $Y2=2.235
r63 1 12 600 $w=1.7e-07 $l=6.01997e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.96 $X2=1.07 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_M%Y 1 2 3 13 16 18 19 20 32 35 39 46 51
r49 33 35 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=1.68 $Y2=1.665
r50 32 39 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.16 $Y2=1.665
r51 19 20 16.2679 $w=3.38e-07 $l=3.95e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=3.035 $Y2=1.665
r52 19 41 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.525 $Y2=1.665
r53 18 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.195 $Y2=1.665
r54 18 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.525 $Y2=1.665
r55 18 51 10.9968 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=2.36 $Y=1.75
+ $X2=2.36 $Y2=2.105
r56 18 39 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.135 $Y=1.665
+ $X2=2.16 $Y2=1.665
r57 16 33 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=1.39 $Y=1.665
+ $X2=1.665 $Y2=1.665
r58 16 46 10.615 $w=3.98e-07 $l=3.55e-07 $layer=LI1_cond $X=1.5 $Y=1.75 $X2=1.5
+ $Y2=2.105
r59 16 18 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.715 $Y=1.665
+ $X2=2.135 $Y2=1.665
r60 16 35 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.715 $Y=1.665
+ $X2=1.68 $Y2=1.665
r61 14 20 33.3012 $w=3.38e-07 $l=9.4e-07 $layer=LI1_cond $X=3.12 $Y=0.64
+ $X2=3.12 $Y2=1.58
r62 13 14 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.12 $Y=0.535
+ $X2=3.12 $Y2=0.64
r63 11 13 9.77056 $w=2.08e-07 $l=1.85e-07 $layer=LI1_cond $X=2.935 $Y=0.535
+ $X2=3.12 $Y2=0.535
r64 3 51 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.96 $X2=2.36 $Y2=2.105
r65 2 46 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.96 $X2=1.5 $Y2=2.105
r66 1 11 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.26 $X2=2.935 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_M%VGND 1 8 10 17 18 21
c31 18 0 7.80944e-20 $X=3.12 $Y=0
r32 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r34 15 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r35 14 17 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r36 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r37 12 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.76
+ $Y2=0
r38 12 14 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.2
+ $Y2=0
r39 10 18 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r40 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r41 6 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0
r42 6 8 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0.405
r43 1 8 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.26 $X2=0.76 $Y2=0.405
.ends

