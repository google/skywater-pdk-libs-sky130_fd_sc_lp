* File: sky130_fd_sc_lp__maj3_lp.pxi.spice
* Created: Fri Aug 28 10:43:18 2020
* 
x_PM_SKY130_FD_SC_LP__MAJ3_LP%A N_A_M1013_g N_A_M1010_g N_A_M1012_g N_A_M1014_g
+ A A N_A_c_85_n PM_SKY130_FD_SC_LP__MAJ3_LP%A
x_PM_SKY130_FD_SC_LP__MAJ3_LP%B N_B_M1004_g N_B_M1000_g N_B_c_135_n N_B_c_136_n
+ N_B_M1002_g N_B_c_137_n N_B_M1011_g N_B_c_138_n N_B_c_148_n N_B_c_139_n
+ N_B_c_140_n N_B_c_141_n N_B_c_142_n N_B_c_143_n B N_B_c_144_n N_B_c_145_n
+ PM_SKY130_FD_SC_LP__MAJ3_LP%B
x_PM_SKY130_FD_SC_LP__MAJ3_LP%C N_C_M1008_g N_C_M1006_g N_C_c_234_n N_C_M1001_g
+ N_C_M1005_g N_C_c_236_n N_C_c_237_n N_C_c_241_n C N_C_c_238_n N_C_c_243_n
+ PM_SKY130_FD_SC_LP__MAJ3_LP%C
x_PM_SKY130_FD_SC_LP__MAJ3_LP%A_29_419# N_A_29_419#_M1000_s N_A_29_419#_M1006_d
+ N_A_29_419#_M1004_s N_A_29_419#_M1008_d N_A_29_419#_c_303_n
+ N_A_29_419#_M1009_g N_A_29_419#_M1003_g N_A_29_419#_c_304_n
+ N_A_29_419#_M1007_g N_A_29_419#_c_305_n N_A_29_419#_c_306_n
+ N_A_29_419#_c_318_n N_A_29_419#_c_323_n N_A_29_419#_c_307_n
+ N_A_29_419#_c_308_n N_A_29_419#_c_309_n N_A_29_419#_c_310_n
+ N_A_29_419#_c_311_n N_A_29_419#_c_312_n N_A_29_419#_c_320_n
+ N_A_29_419#_c_313_n N_A_29_419#_c_330_n N_A_29_419#_c_314_n
+ N_A_29_419#_c_322_n N_A_29_419#_c_362_n N_A_29_419#_c_315_n
+ PM_SKY130_FD_SC_LP__MAJ3_LP%A_29_419#
x_PM_SKY130_FD_SC_LP__MAJ3_LP%VPWR N_VPWR_M1013_d N_VPWR_M1005_d N_VPWR_c_441_n
+ N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n VPWR N_VPWR_c_445_n
+ N_VPWR_c_446_n N_VPWR_c_440_n N_VPWR_c_448_n PM_SKY130_FD_SC_LP__MAJ3_LP%VPWR
x_PM_SKY130_FD_SC_LP__MAJ3_LP%X N_X_M1007_d N_X_M1003_d N_X_c_493_n X X X
+ N_X_c_496_n N_X_c_494_n PM_SKY130_FD_SC_LP__MAJ3_LP%X
x_PM_SKY130_FD_SC_LP__MAJ3_LP%VGND N_VGND_M1010_d N_VGND_M1001_d N_VGND_c_518_n
+ N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n VGND N_VGND_c_522_n
+ N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n PM_SKY130_FD_SC_LP__MAJ3_LP%VGND
cc_1 VNB N_A_M1010_g 0.0397043f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.835
cc_2 VNB N_A_M1014_g 0.0392678f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=0.835
cc_3 VNB A 9.25061e-19 $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.95
cc_4 VNB N_A_c_85_n 0.0132081f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.77
cc_5 VNB N_B_M1000_g 0.0432027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B_c_135_n 0.134757f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.935
cc_7 VNB N_B_c_136_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=2.595
cc_8 VNB N_B_c_137_n 0.0164779f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=0.835
cc_9 VNB N_B_c_138_n 0.0164321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_139_n 0.0209475f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.77
cc_11 VNB N_B_c_140_n 0.00293005f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.877
cc_12 VNB N_B_c_141_n 0.00811599f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.877
cc_13 VNB N_B_c_142_n 0.00171029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_143_n 0.0213307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_144_n 0.0101187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_145_n 0.00346345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_M1008_g 0.0181153f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=2.595
cc_18 VNB N_C_M1006_g 0.0238068f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.835
cc_19 VNB N_C_c_234_n 0.0385832f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.935
cc_20 VNB N_C_M1001_g 0.0426967f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.605
cc_21 VNB N_C_c_236_n 0.00641209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C_c_237_n 0.012669f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.77
cc_23 VNB N_C_c_238_n 0.0210869f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.77
cc_24 VNB N_A_29_419#_c_303_n 0.0140634f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.605
cc_25 VNB N_A_29_419#_c_304_n 0.0192954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_29_419#_c_305_n 0.0216946f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.77
cc_27 VNB N_A_29_419#_c_306_n 0.0117033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_29_419#_c_307_n 0.0387914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_29_419#_c_308_n 0.00265501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_29_419#_c_309_n 0.00628188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_29_419#_c_310_n 0.0303304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_29_419#_c_311_n 0.0051256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_29_419#_c_312_n 0.0375605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_29_419#_c_313_n 0.0291088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_29_419#_c_314_n 0.00120759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_29_419#_c_315_n 0.0021627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_440_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_493_n 0.025686f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=2.595
cc_39 VNB N_X_c_494_n 0.040914f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.877
cc_40 VNB N_VGND_c_518_n 0.0117822f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.935
cc_41 VNB N_VGND_c_519_n 0.00319234f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.605
cc_42 VNB N_VGND_c_520_n 0.0382009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_521_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_44 VNB N_VGND_c_522_n 0.0448225f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.77
cc_45 VNB N_VGND_c_523_n 0.0278279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_524_n 0.262995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_525_n 0.00567616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_A_M1013_g 0.0238502f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=2.595
cc_49 VPB N_A_M1012_g 0.0228076f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=2.595
cc_50 VPB A 0.00462222f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.95
cc_51 VPB N_A_c_85_n 0.0336366f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=1.77
cc_52 VPB N_B_M1004_g 0.0324526f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=2.595
cc_53 VPB N_B_M1002_g 0.0268629f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.605
cc_54 VPB N_B_c_148_n 0.0147435f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.77
cc_55 VPB N_B_c_140_n 0.00102516f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.877
cc_56 VPB N_B_c_141_n 0.0200005f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.877
cc_57 VPB N_B_c_142_n 8.8959e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B_c_143_n 0.00561291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_C_M1008_g 0.0418295f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=2.595
cc_60 VPB N_C_M1005_g 0.0266551f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_61 VPB N_C_c_241_n 0.0137134f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=1.77
cc_62 VPB N_C_c_238_n 0.00654426f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.77
cc_63 VPB N_C_c_243_n 0.00164715f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.877
cc_64 VPB N_A_29_419#_M1003_g 0.050586f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.95
cc_65 VPB N_A_29_419#_c_306_n 0.00225458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_29_419#_c_318_n 0.0228071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_29_419#_c_311_n 8.75463e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_29_419#_c_320_n 0.0244238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_29_419#_c_313_n 0.0201036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_29_419#_c_322_n 0.00634721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_441_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=1.625 $Y2=1.935
cc_72 VPB N_VPWR_c_442_n 0.00765718f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.605
cc_73 VPB N_VPWR_c_443_n 0.0485959f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.95
cc_74 VPB N_VPWR_c_444_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_445_n 0.0357749f $X=-0.19 $Y=1.655 $X2=1.095 $Y2=1.77
cc_76 VPB N_VPWR_c_446_n 0.0215793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_440_n 0.0464208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_448_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.018649f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.605
cc_80 VPB N_X_c_496_n 0.0414962f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.77
cc_81 VPB N_X_c_494_n 0.0132352f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.877
cc_82 N_A_M1010_g N_B_M1000_g 0.0479575f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_83 N_A_M1010_g N_B_c_135_n 0.00861299f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_84 N_A_M1014_g N_B_c_135_n 0.00865297f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_85 N_A_M1013_g N_B_c_148_n 0.0533063f $X=1.095 $Y=2.595 $X2=0 $Y2=0
cc_86 N_A_M1014_g N_B_c_139_n 0.0109755f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_87 A N_B_c_140_n 0.00968582f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_88 N_A_M1010_g N_B_c_142_n 0.0012627f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_89 A N_B_c_142_n 0.0136936f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_90 N_A_c_85_n N_B_c_142_n 0.00121431f $X=1.625 $Y=1.77 $X2=0 $Y2=0
cc_91 N_A_M1010_g N_B_c_143_n 0.0127515f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_92 A N_B_c_143_n 0.00203758f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_93 N_A_c_85_n N_B_c_143_n 0.0533063f $X=1.625 $Y=1.77 $X2=0 $Y2=0
cc_94 N_A_M1010_g N_B_c_144_n 0.00773469f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_95 N_A_c_85_n N_B_c_144_n 0.00162488f $X=1.625 $Y=1.77 $X2=0 $Y2=0
cc_96 N_A_M1010_g N_B_c_145_n 0.00794853f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_97 N_A_M1014_g N_B_c_145_n 0.00140944f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_98 A N_B_c_145_n 0.0507271f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_99 N_A_c_85_n N_B_c_145_n 0.00638043f $X=1.625 $Y=1.77 $X2=0 $Y2=0
cc_100 A N_C_M1008_g 0.00885459f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_101 N_A_c_85_n N_C_M1008_g 0.0646455f $X=1.625 $Y=1.77 $X2=0 $Y2=0
cc_102 N_A_M1014_g N_C_M1006_g 0.0391908f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_103 N_A_M1014_g N_C_c_236_n 0.0646455f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_104 N_A_M1013_g N_A_29_419#_c_323_n 0.0201962f $X=1.095 $Y=2.595 $X2=0 $Y2=0
cc_105 N_A_M1012_g N_A_29_419#_c_323_n 0.0167309f $X=1.625 $Y=2.595 $X2=0 $Y2=0
cc_106 A N_A_29_419#_c_323_n 0.0400158f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_107 N_A_c_85_n N_A_29_419#_c_323_n 4.2819e-19 $X=1.625 $Y=1.77 $X2=0 $Y2=0
cc_108 N_A_M1010_g N_A_29_419#_c_307_n 0.00124819f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_109 N_A_M1014_g N_A_29_419#_c_308_n 0.00586359f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_110 A N_A_29_419#_c_320_n 0.00136826f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_111 N_A_M1010_g N_A_29_419#_c_330_n 0.0106187f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_112 N_A_M1010_g N_A_29_419#_c_314_n 0.00153295f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_113 N_A_M1014_g N_A_29_419#_c_314_n 0.00734174f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_114 N_A_M1012_g N_A_29_419#_c_322_n 0.00268335f $X=1.625 $Y=2.595 $X2=0 $Y2=0
cc_115 A N_VPWR_M1013_d 0.001878f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_116 N_A_M1013_g N_VPWR_c_441_n 0.0136445f $X=1.095 $Y=2.595 $X2=0 $Y2=0
cc_117 N_A_M1012_g N_VPWR_c_441_n 0.014498f $X=1.625 $Y=2.595 $X2=0 $Y2=0
cc_118 N_A_M1012_g N_VPWR_c_443_n 0.008763f $X=1.625 $Y=2.595 $X2=0 $Y2=0
cc_119 N_A_M1013_g N_VPWR_c_445_n 0.008763f $X=1.095 $Y=2.595 $X2=0 $Y2=0
cc_120 N_A_M1013_g N_VPWR_c_440_n 0.00763092f $X=1.095 $Y=2.595 $X2=0 $Y2=0
cc_121 N_A_M1012_g N_VPWR_c_440_n 0.00763092f $X=1.625 $Y=2.595 $X2=0 $Y2=0
cc_122 N_A_M1010_g N_VGND_c_518_n 0.00365006f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_123 N_A_M1014_g N_VGND_c_518_n 0.00225474f $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_124 N_A_M1010_g N_VGND_c_524_n 9.49986e-19 $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_125 N_A_M1014_g N_VGND_c_524_n 9.49986e-19 $X=1.675 $Y=0.835 $X2=0 $Y2=0
cc_126 N_B_M1002_g N_C_M1008_g 0.0272214f $X=2.615 $Y=2.595 $X2=0 $Y2=0
cc_127 N_B_c_139_n N_C_M1008_g 0.0131634f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_128 N_B_c_140_n N_C_M1008_g 0.00783312f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_129 N_B_c_141_n N_C_M1008_g 0.0211441f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_130 N_B_c_135_n N_C_M1006_g 0.00868355f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_131 N_B_c_137_n N_C_M1006_g 0.00710069f $X=2.575 $Y=0.255 $X2=0 $Y2=0
cc_132 N_B_c_137_n N_C_c_234_n 0.00465755f $X=2.575 $Y=0.255 $X2=0 $Y2=0
cc_133 N_B_c_139_n N_C_c_234_n 0.0164996f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_134 N_B_c_141_n N_C_c_234_n 0.0214008f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_135 N_B_c_135_n N_C_M1001_g 0.026078f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_136 N_B_M1002_g N_C_M1005_g 0.0705419f $X=2.615 $Y=2.595 $X2=0 $Y2=0
cc_137 N_B_c_139_n N_C_c_236_n 0.00749248f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_138 N_B_c_139_n N_C_c_238_n 8.93328e-19 $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_139 N_B_c_140_n N_C_c_238_n 0.0049248f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_140 N_B_c_141_n N_C_c_238_n 0.0200799f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_141 N_B_c_139_n N_C_c_243_n 0.0116028f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_142 N_B_c_140_n N_C_c_243_n 0.0323329f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_143 N_B_c_141_n N_C_c_243_n 0.00114872f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_144 N_B_M1004_g N_A_29_419#_c_323_n 0.019686f $X=0.635 $Y=2.595 $X2=0 $Y2=0
cc_145 N_B_c_142_n N_A_29_419#_c_323_n 0.00991405f $X=0.595 $Y=1.39 $X2=0 $Y2=0
cc_146 N_B_M1000_g N_A_29_419#_c_307_n 0.00722899f $X=0.695 $Y=0.835 $X2=0 $Y2=0
cc_147 N_B_c_138_n N_A_29_419#_c_307_n 0.00162796f $X=0.6 $Y=1.375 $X2=0 $Y2=0
cc_148 N_B_c_142_n N_A_29_419#_c_307_n 0.0141894f $X=0.595 $Y=1.39 $X2=0 $Y2=0
cc_149 N_B_c_135_n N_A_29_419#_c_308_n 0.00456581f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_150 N_B_c_135_n N_A_29_419#_c_309_n 0.00514449f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_151 N_B_c_137_n N_A_29_419#_c_309_n 0.0134089f $X=2.575 $Y=0.255 $X2=0 $Y2=0
cc_152 N_B_c_137_n N_A_29_419#_c_310_n 0.00355141f $X=2.575 $Y=0.255 $X2=0 $Y2=0
cc_153 N_B_c_139_n N_A_29_419#_c_310_n 0.0171588f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_154 N_B_M1004_g N_A_29_419#_c_320_n 0.00570042f $X=0.635 $Y=2.595 $X2=0 $Y2=0
cc_155 N_B_c_148_n N_A_29_419#_c_320_n 6.23284e-19 $X=0.595 $Y=1.895 $X2=0 $Y2=0
cc_156 N_B_c_142_n N_A_29_419#_c_320_n 0.00110853f $X=0.595 $Y=1.39 $X2=0 $Y2=0
cc_157 N_B_M1004_g N_A_29_419#_c_313_n 0.00431633f $X=0.635 $Y=2.595 $X2=0 $Y2=0
cc_158 N_B_M1000_g N_A_29_419#_c_313_n 0.00362326f $X=0.695 $Y=0.835 $X2=0 $Y2=0
cc_159 N_B_c_138_n N_A_29_419#_c_313_n 0.0150793f $X=0.6 $Y=1.375 $X2=0 $Y2=0
cc_160 N_B_c_142_n N_A_29_419#_c_313_n 0.0488992f $X=0.595 $Y=1.39 $X2=0 $Y2=0
cc_161 N_B_M1000_g N_A_29_419#_c_330_n 0.00859422f $X=0.695 $Y=0.835 $X2=0 $Y2=0
cc_162 N_B_c_135_n N_A_29_419#_c_330_n 0.00427163f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_163 N_B_c_139_n N_A_29_419#_c_330_n 0.010189f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_164 N_B_c_142_n N_A_29_419#_c_330_n 0.00695762f $X=0.595 $Y=1.39 $X2=0 $Y2=0
cc_165 N_B_c_144_n N_A_29_419#_c_330_n 0.0158646f $X=1.085 $Y=1.297 $X2=0 $Y2=0
cc_166 N_B_c_145_n N_A_29_419#_c_330_n 0.0142786f $X=1.315 $Y=1.297 $X2=0 $Y2=0
cc_167 N_B_c_135_n N_A_29_419#_c_314_n 2.22778e-19 $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_168 N_B_c_139_n N_A_29_419#_c_314_n 0.0482616f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_169 N_B_M1002_g N_A_29_419#_c_322_n 0.00888631f $X=2.615 $Y=2.595 $X2=0 $Y2=0
cc_170 N_B_c_140_n N_A_29_419#_c_322_n 0.0051969f $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_171 N_B_c_141_n N_A_29_419#_c_322_n 3.63443e-19 $X=2.585 $Y=1.75 $X2=0 $Y2=0
cc_172 N_B_M1002_g N_A_29_419#_c_362_n 0.0137975f $X=2.615 $Y=2.595 $X2=0 $Y2=0
cc_173 N_B_c_139_n N_A_29_419#_c_315_n 0.02628f $X=2.42 $Y=1.33 $X2=0 $Y2=0
cc_174 N_B_M1004_g N_VPWR_c_441_n 0.0027374f $X=0.635 $Y=2.595 $X2=0 $Y2=0
cc_175 N_B_M1002_g N_VPWR_c_442_n 0.0052133f $X=2.615 $Y=2.595 $X2=0 $Y2=0
cc_176 N_B_M1002_g N_VPWR_c_443_n 0.00939541f $X=2.615 $Y=2.595 $X2=0 $Y2=0
cc_177 N_B_M1004_g N_VPWR_c_445_n 0.00975641f $X=0.635 $Y=2.595 $X2=0 $Y2=0
cc_178 N_B_M1004_g N_VPWR_c_440_n 0.010641f $X=0.635 $Y=2.595 $X2=0 $Y2=0
cc_179 N_B_M1002_g N_VPWR_c_440_n 0.0161801f $X=2.615 $Y=2.595 $X2=0 $Y2=0
cc_180 N_B_M1000_g N_VGND_c_518_n 0.00692076f $X=0.695 $Y=0.835 $X2=0 $Y2=0
cc_181 N_B_c_135_n N_VGND_c_518_n 0.0251785f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_182 N_B_c_135_n N_VGND_c_519_n 0.00387647f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_183 N_B_c_136_n N_VGND_c_520_n 0.0215833f $X=0.77 $Y=0.18 $X2=0 $Y2=0
cc_184 N_B_c_135_n N_VGND_c_522_n 0.0351706f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_185 N_B_c_135_n N_VGND_c_524_n 0.0577927f $X=2.5 $Y=0.18 $X2=0 $Y2=0
cc_186 N_B_c_136_n N_VGND_c_524_n 0.00672709f $X=0.77 $Y=0.18 $X2=0 $Y2=0
cc_187 N_C_M1001_g N_A_29_419#_c_303_n 0.0195942f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_188 N_C_M1005_g N_A_29_419#_M1003_g 0.0143068f $X=3.115 $Y=2.595 $X2=0 $Y2=0
cc_189 N_C_c_241_n N_A_29_419#_M1003_g 0.0127715f $X=3.125 $Y=1.915 $X2=0 $Y2=0
cc_190 N_C_c_243_n N_A_29_419#_M1003_g 0.00175947f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_191 N_C_c_238_n N_A_29_419#_c_306_n 0.0127715f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_192 N_C_M1008_g N_A_29_419#_c_323_n 0.020894f $X=2.085 $Y=2.595 $X2=0 $Y2=0
cc_193 N_C_M1006_g N_A_29_419#_c_308_n 0.0131741f $X=2.065 $Y=0.835 $X2=0 $Y2=0
cc_194 N_C_c_236_n N_A_29_419#_c_308_n 8.03654e-19 $X=2.085 $Y=1.3 $X2=0 $Y2=0
cc_195 N_C_M1006_g N_A_29_419#_c_309_n 0.00345837f $X=2.065 $Y=0.835 $X2=0 $Y2=0
cc_196 N_C_M1001_g N_A_29_419#_c_309_n 0.00215559f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_197 N_C_c_234_n N_A_29_419#_c_310_n 0.00688568f $X=2.96 $Y=1.3 $X2=0 $Y2=0
cc_198 N_C_M1001_g N_A_29_419#_c_310_n 0.0167116f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_199 N_C_c_237_n N_A_29_419#_c_310_n 0.00482313f $X=3.125 $Y=1.3 $X2=0 $Y2=0
cc_200 N_C_c_243_n N_A_29_419#_c_310_n 0.0245048f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_201 N_C_M1001_g N_A_29_419#_c_311_n 0.00297244f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_202 N_C_c_237_n N_A_29_419#_c_311_n 0.0030294f $X=3.125 $Y=1.3 $X2=0 $Y2=0
cc_203 N_C_c_243_n N_A_29_419#_c_311_n 0.0254875f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_204 N_C_M1001_g N_A_29_419#_c_312_n 0.00596958f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_205 N_C_c_237_n N_A_29_419#_c_312_n 0.0127715f $X=3.125 $Y=1.3 $X2=0 $Y2=0
cc_206 N_C_c_243_n N_A_29_419#_c_312_n 5.19096e-19 $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_207 N_C_M1006_g N_A_29_419#_c_314_n 2.00237e-19 $X=2.065 $Y=0.835 $X2=0 $Y2=0
cc_208 N_C_M1008_g N_A_29_419#_c_322_n 0.00701617f $X=2.085 $Y=2.595 $X2=0 $Y2=0
cc_209 N_C_M1005_g N_A_29_419#_c_322_n 0.00418715f $X=3.115 $Y=2.595 $X2=0 $Y2=0
cc_210 N_C_M1008_g N_A_29_419#_c_362_n 0.014306f $X=2.085 $Y=2.595 $X2=0 $Y2=0
cc_211 N_C_c_234_n N_A_29_419#_c_315_n 0.00619687f $X=2.96 $Y=1.3 $X2=0 $Y2=0
cc_212 N_C_M1008_g N_VPWR_c_441_n 0.0020846f $X=2.085 $Y=2.595 $X2=0 $Y2=0
cc_213 N_C_M1005_g N_VPWR_c_442_n 0.0251726f $X=3.115 $Y=2.595 $X2=0 $Y2=0
cc_214 N_C_c_243_n N_VPWR_c_442_n 0.00387242f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_215 N_C_M1008_g N_VPWR_c_443_n 0.00939541f $X=2.085 $Y=2.595 $X2=0 $Y2=0
cc_216 N_C_M1005_g N_VPWR_c_443_n 0.008763f $X=3.115 $Y=2.595 $X2=0 $Y2=0
cc_217 N_C_M1008_g N_VPWR_c_440_n 0.00931035f $X=2.085 $Y=2.595 $X2=0 $Y2=0
cc_218 N_C_M1005_g N_VPWR_c_440_n 0.0144844f $X=3.115 $Y=2.595 $X2=0 $Y2=0
cc_219 N_C_M1005_g X 7.46468e-19 $X=3.115 $Y=2.595 $X2=0 $Y2=0
cc_220 N_C_M1001_g N_VGND_c_519_n 0.0117152f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_221 N_C_M1001_g N_VGND_c_522_n 0.0040395f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_222 N_C_M1006_g N_VGND_c_524_n 9.49986e-19 $X=2.065 $Y=0.835 $X2=0 $Y2=0
cc_223 N_C_M1001_g N_VGND_c_524_n 0.00780354f $X=3.035 $Y=0.55 $X2=0 $Y2=0
cc_224 N_A_29_419#_c_323_n A_152_419# 0.00557654f $X=2.185 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A_29_419#_c_323_n N_VPWR_M1013_d 0.00343453f $X=2.185 $Y=2.415
+ $X2=-0.19 $Y2=-0.245
cc_226 N_A_29_419#_c_323_n N_VPWR_c_441_n 0.0159912f $X=2.185 $Y=2.415 $X2=0
+ $Y2=0
cc_227 N_A_29_419#_c_362_n N_VPWR_c_441_n 0.00930336f $X=2.35 $Y=2.415 $X2=0
+ $Y2=0
cc_228 N_A_29_419#_M1003_g N_VPWR_c_442_n 0.022576f $X=3.655 $Y=2.595 $X2=0
+ $Y2=0
cc_229 N_A_29_419#_c_311_n N_VPWR_c_442_n 6.2302e-19 $X=3.695 $Y=1.15 $X2=0
+ $Y2=0
cc_230 N_A_29_419#_c_362_n N_VPWR_c_443_n 0.0177952f $X=2.35 $Y=2.415 $X2=0
+ $Y2=0
cc_231 N_A_29_419#_c_318_n N_VPWR_c_445_n 0.0240223f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_232 N_A_29_419#_M1003_g N_VPWR_c_446_n 0.00879225f $X=3.655 $Y=2.595 $X2=0
+ $Y2=0
cc_233 N_A_29_419#_M1004_s N_VPWR_c_440_n 0.00334885f $X=0.145 $Y=2.095 $X2=0
+ $Y2=0
cc_234 N_A_29_419#_M1008_d N_VPWR_c_440_n 0.00223819f $X=2.21 $Y=2.095 $X2=0
+ $Y2=0
cc_235 N_A_29_419#_M1003_g N_VPWR_c_440_n 0.015232f $X=3.655 $Y=2.595 $X2=0
+ $Y2=0
cc_236 N_A_29_419#_c_318_n N_VPWR_c_440_n 0.0140402f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_237 N_A_29_419#_c_323_n N_VPWR_c_440_n 0.043277f $X=2.185 $Y=2.415 $X2=0
+ $Y2=0
cc_238 N_A_29_419#_c_362_n N_VPWR_c_440_n 0.0123247f $X=2.35 $Y=2.415 $X2=0
+ $Y2=0
cc_239 N_A_29_419#_c_323_n A_350_419# 0.00557654f $X=2.185 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A_29_419#_c_303_n N_X_c_493_n 0.00140093f $X=3.465 $Y=0.835 $X2=0 $Y2=0
cc_241 N_A_29_419#_c_304_n N_X_c_493_n 0.0101099f $X=3.825 $Y=0.835 $X2=0 $Y2=0
cc_242 N_A_29_419#_M1003_g X 0.00885306f $X=3.655 $Y=2.595 $X2=0 $Y2=0
cc_243 N_A_29_419#_c_306_n X 5.86766e-19 $X=3.695 $Y=1.655 $X2=0 $Y2=0
cc_244 N_A_29_419#_c_311_n X 0.00645791f $X=3.695 $Y=1.15 $X2=0 $Y2=0
cc_245 N_A_29_419#_M1003_g N_X_c_496_n 0.0220366f $X=3.655 $Y=2.595 $X2=0 $Y2=0
cc_246 N_A_29_419#_M1003_g N_X_c_494_n 0.00707421f $X=3.655 $Y=2.595 $X2=0 $Y2=0
cc_247 N_A_29_419#_c_304_n N_X_c_494_n 0.00508967f $X=3.825 $Y=0.835 $X2=0 $Y2=0
cc_248 N_A_29_419#_c_310_n N_X_c_494_n 0.0103001f $X=3.525 $Y=0.98 $X2=0 $Y2=0
cc_249 N_A_29_419#_c_311_n N_X_c_494_n 0.0424501f $X=3.695 $Y=1.15 $X2=0 $Y2=0
cc_250 N_A_29_419#_c_312_n N_X_c_494_n 0.0136754f $X=3.695 $Y=1.15 $X2=0 $Y2=0
cc_251 N_A_29_419#_c_330_n A_154_125# 0.00297367f $X=1.495 $Y=0.947 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_29_419#_c_330_n N_VGND_M1010_d 0.00648334f $X=1.495 $Y=0.947
+ $X2=-0.19 $Y2=-0.245
cc_253 N_A_29_419#_c_314_n N_VGND_M1010_d 0.0011772f $X=1.665 $Y=0.947 $X2=-0.19
+ $Y2=-0.245
cc_254 N_A_29_419#_c_307_n N_VGND_c_518_n 9.61732e-19 $X=0.645 $Y=0.915 $X2=0
+ $Y2=0
cc_255 N_A_29_419#_c_309_n N_VGND_c_518_n 0.00984874f $X=2.36 $Y=0.55 $X2=0
+ $Y2=0
cc_256 N_A_29_419#_c_330_n N_VGND_c_518_n 0.0247764f $X=1.495 $Y=0.947 $X2=0
+ $Y2=0
cc_257 N_A_29_419#_c_303_n N_VGND_c_519_n 0.0107512f $X=3.465 $Y=0.835 $X2=0
+ $Y2=0
cc_258 N_A_29_419#_c_304_n N_VGND_c_519_n 0.00174671f $X=3.825 $Y=0.835 $X2=0
+ $Y2=0
cc_259 N_A_29_419#_c_309_n N_VGND_c_519_n 0.0111185f $X=2.36 $Y=0.55 $X2=0 $Y2=0
cc_260 N_A_29_419#_c_310_n N_VGND_c_519_n 0.0207959f $X=3.525 $Y=0.98 $X2=0
+ $Y2=0
cc_261 N_A_29_419#_c_307_n N_VGND_c_520_n 0.00683664f $X=0.645 $Y=0.915 $X2=0
+ $Y2=0
cc_262 N_A_29_419#_c_309_n N_VGND_c_522_n 0.0165487f $X=2.36 $Y=0.55 $X2=0 $Y2=0
cc_263 N_A_29_419#_c_303_n N_VGND_c_523_n 0.0040395f $X=3.465 $Y=0.835 $X2=0
+ $Y2=0
cc_264 N_A_29_419#_c_304_n N_VGND_c_523_n 0.00457319f $X=3.825 $Y=0.835 $X2=0
+ $Y2=0
cc_265 N_A_29_419#_c_303_n N_VGND_c_524_n 0.00772493f $X=3.465 $Y=0.835 $X2=0
+ $Y2=0
cc_266 N_A_29_419#_c_304_n N_VGND_c_524_n 0.00895391f $X=3.825 $Y=0.835 $X2=0
+ $Y2=0
cc_267 N_A_29_419#_c_305_n N_VGND_c_524_n 7.69802e-19 $X=3.825 $Y=0.91 $X2=0
+ $Y2=0
cc_268 N_A_29_419#_c_307_n N_VGND_c_524_n 0.00991258f $X=0.645 $Y=0.915 $X2=0
+ $Y2=0
cc_269 N_A_29_419#_c_309_n N_VGND_c_524_n 0.0109692f $X=2.36 $Y=0.55 $X2=0 $Y2=0
cc_270 N_A_29_419#_c_330_n N_VGND_c_524_n 0.0178749f $X=1.495 $Y=0.947 $X2=0
+ $Y2=0
cc_271 N_A_29_419#_c_314_n N_VGND_c_524_n 0.00365467f $X=1.665 $Y=0.947 $X2=0
+ $Y2=0
cc_272 N_A_29_419#_c_308_n A_350_125# 0.002181f $X=2.195 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_273 A_152_419# N_VPWR_c_440_n 0.00305025f $X=0.76 $Y=2.095 $X2=0 $Y2=0
cc_274 N_VPWR_c_440_n A_350_419# 0.00305025f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_275 N_VPWR_c_440_n A_548_419# 0.0107073f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_276 N_VPWR_c_440_n N_X_M1003_d 0.0023218f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_277 N_VPWR_c_442_n X 0.0629875f $X=3.38 $Y=2.26 $X2=0 $Y2=0
cc_278 N_VPWR_c_446_n N_X_c_496_n 0.0281861f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_c_440_n N_X_c_496_n 0.0173447f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_280 N_X_c_493_n N_VGND_c_519_n 0.0132309f $X=4.04 $Y=0.55 $X2=0 $Y2=0
cc_281 N_X_c_493_n N_VGND_c_523_n 0.0165806f $X=4.04 $Y=0.55 $X2=0 $Y2=0
cc_282 N_X_c_493_n N_VGND_c_524_n 0.0123279f $X=4.04 $Y=0.55 $X2=0 $Y2=0
