* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__einvp_lp A TE VGND VNB VPB VPWR Z
X0 a_314_101# TE a_182_321# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 Z A a_134_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_134_419# a_182_321# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND TE a_314_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_134_141# TE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Z A a_134_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR TE a_182_321# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
