* NGSPICE file created from sky130_fd_sc_lp__o221a_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o221a_lp A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VPWR a_84_21# X VPB phighvt w=1e+06u l=250000u
+  ad=6.65e+11p pd=5.33e+06u as=2.85e+11p ps=2.57e+06u
M1001 a_84_21# A2 a_270_419# VPB phighvt w=1e+06u l=250000u
+  ad=6.05e+11p pd=5.21e+06u as=2.4e+11p ps=2.48e+06u
M1002 a_114_47# a_84_21# X VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1003 a_272_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=2.85425e+11p pd=3.15e+06u as=2.973e+11p ps=3.16e+06u
M1004 VPWR B1 a_482_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1005 a_270_419# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_272_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_272_47# B2 a_490_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1008 a_482_419# B2 a_84_21# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_84_21# a_114_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_84_21# C1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_490_141# B1 a_272_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_84_21# C1 a_490_141# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

