* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_2067_92# a_1920_119# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1575_119# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1232_463# a_1274_401# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR SET_B a_1920_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_1848_119# a_901_441# a_1920_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 VPWR a_1146_463# a_1274_401# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1274_401# a_1146_463# a_1575_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_640_481# a_901_441# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_1146_463# a_1848_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 VGND CLK a_640_481# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_275_481# a_640_481# a_1146_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 Q a_2582_150# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_275_481# a_901_441# a_1146_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_2097_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_640_481# a_901_441# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_34_481# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_34_481# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_275_481# a_34_481# a_383_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_383_481# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VGND a_34_481# a_252_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1146_463# a_1818_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_2025_488# a_2067_92# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VPWR a_1920_119# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_2025_118# a_2067_92# a_2097_118# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR SCE a_203_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_203_481# D a_275_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_1818_379# a_640_481# a_1920_119# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_252_47# D a_275_481# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_1146_463# a_901_441# a_1245_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1146_463# a_640_481# a_1232_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VGND a_1920_119# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_275_481# SCE a_478_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1920_119# a_901_441# a_2025_488# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_2067_92# a_1920_119# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 Q a_2582_150# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 VPWR a_1920_119# a_2582_150# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 VPWR CLK a_640_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 a_1245_119# a_1274_401# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_1274_401# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X39 a_1920_119# a_640_481# a_2025_118# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VGND a_1920_119# a_2582_150# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_478_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
