* File: sky130_fd_sc_lp__a41oi_1.spice
* Created: Fri Aug 28 10:03:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a41oi_1  VNB VPB B1 A4 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_B1_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3066 AS=0.2226 PD=1.57 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1009 A_304_47# N_A4_M1009_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.3066 PD=1.12 PS=1.57 NRD=12.132 NRS=0 M=1 R=5.6 SA=75001.1 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1002 A_390_47# N_A3_M1002_g A_304_47# VNB NSHORT L=0.15 W=0.84 AD=0.1764
+ AS=0.1176 PD=1.26 PS=1.12 NRD=22.14 NRS=12.132 M=1 R=5.6 SA=75001.5 SB=75001.2
+ A=0.126 P=1.98 MULT=1
MM1006 A_504_47# N_A2_M1006_g A_390_47# VNB NSHORT L=0.15 W=0.84 AD=0.1218
+ AS=0.1764 PD=1.13 PS=1.26 NRD=12.852 NRS=22.14 M=1 R=5.6 SA=75002.1 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g A_504_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1218 PD=2.21 PS=1.13 NRD=0 NRS=12.852 M=1 R=5.6 SA=75002.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1001 N_A_128_367#_M1001_d N_B1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.21105 AS=0.3339 PD=1.595 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A4_M1004_g N_A_128_367#_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.49455 AS=0.21105 PD=2.045 PS=1.595 NRD=0 NRS=8.5892 M=1 R=8.4
+ SA=75000.7 SB=75002 A=0.189 P=2.82 MULT=1
MM1000 N_A_128_367#_M1000_d N_A3_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.49455 PD=1.54 PS=2.045 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_128_367#_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75002
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1005 N_A_128_367#_M1005_d N_A1_M1005_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75002.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a41oi_1.pxi.spice"
*
.ends
*
*
