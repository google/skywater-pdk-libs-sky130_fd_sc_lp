* File: sky130_fd_sc_lp__o21ba_4.pxi.spice
* Created: Wed Sep  2 10:16:57 2020
* 
x_PM_SKY130_FD_SC_LP__O21BA_4%B1_N N_B1_N_M1020_g N_B1_N_M1021_g B1_N B1_N
+ N_B1_N_c_108_n N_B1_N_c_109_n PM_SKY130_FD_SC_LP__O21BA_4%B1_N
x_PM_SKY130_FD_SC_LP__O21BA_4%A_180_23# N_A_180_23#_M1001_s N_A_180_23#_M1006_d
+ N_A_180_23#_M1004_d N_A_180_23#_M1007_g N_A_180_23#_M1000_g
+ N_A_180_23#_M1009_g N_A_180_23#_M1002_g N_A_180_23#_M1016_g
+ N_A_180_23#_M1003_g N_A_180_23#_M1019_g N_A_180_23#_M1018_g
+ N_A_180_23#_c_146_n N_A_180_23#_c_147_n N_A_180_23#_c_148_n
+ N_A_180_23#_c_259_p N_A_180_23#_c_149_n N_A_180_23#_c_170_p
+ N_A_180_23#_c_150_n N_A_180_23#_c_151_n N_A_180_23#_c_199_p
+ N_A_180_23#_c_202_p N_A_180_23#_c_152_n N_A_180_23#_c_153_n
+ PM_SKY130_FD_SC_LP__O21BA_4%A_180_23#
x_PM_SKY130_FD_SC_LP__O21BA_4%A_37_49# N_A_37_49#_M1020_s N_A_37_49#_M1021_s
+ N_A_37_49#_M1006_g N_A_37_49#_M1001_g N_A_37_49#_M1011_g N_A_37_49#_M1013_g
+ N_A_37_49#_c_306_n N_A_37_49#_c_312_n N_A_37_49#_c_313_n N_A_37_49#_c_320_n
+ N_A_37_49#_c_365_p N_A_37_49#_c_314_n N_A_37_49#_c_315_n N_A_37_49#_c_307_n
+ N_A_37_49#_c_316_n N_A_37_49#_c_308_n N_A_37_49#_c_318_n N_A_37_49#_c_309_n
+ PM_SKY130_FD_SC_LP__O21BA_4%A_37_49#
x_PM_SKY130_FD_SC_LP__O21BA_4%A1 N_A1_M1005_g N_A1_M1010_g N_A1_M1008_g
+ N_A1_M1014_g N_A1_c_412_n N_A1_c_406_n N_A1_c_414_n N_A1_c_407_n N_A1_c_455_p
+ N_A1_c_408_n N_A1_c_409_n A1 A1 A1 PM_SKY130_FD_SC_LP__O21BA_4%A1
x_PM_SKY130_FD_SC_LP__O21BA_4%A2 N_A2_M1012_g N_A2_M1004_g N_A2_M1017_g
+ N_A2_M1015_g A2 N_A2_c_496_n N_A2_c_493_n PM_SKY130_FD_SC_LP__O21BA_4%A2
x_PM_SKY130_FD_SC_LP__O21BA_4%VPWR N_VPWR_M1021_d N_VPWR_M1002_d N_VPWR_M1018_d
+ N_VPWR_M1011_s N_VPWR_M1014_d N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_575_n
+ N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n VPWR N_VPWR_c_556_n
+ N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n
+ N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_550_n
+ PM_SKY130_FD_SC_LP__O21BA_4%VPWR
x_PM_SKY130_FD_SC_LP__O21BA_4%X N_X_M1007_s N_X_M1016_s N_X_M1000_s N_X_M1003_s
+ N_X_c_656_n N_X_c_652_n N_X_c_653_n N_X_c_698_p N_X_c_654_n X X X X
+ N_X_c_662_n PM_SKY130_FD_SC_LP__O21BA_4%X
x_PM_SKY130_FD_SC_LP__O21BA_4%A_878_367# N_A_878_367#_M1010_s
+ N_A_878_367#_M1015_s N_A_878_367#_c_705_n
+ PM_SKY130_FD_SC_LP__O21BA_4%A_878_367#
x_PM_SKY130_FD_SC_LP__O21BA_4%VGND N_VGND_M1020_d N_VGND_M1009_d N_VGND_M1019_d
+ N_VGND_M1005_d N_VGND_M1017_s N_VGND_c_717_n N_VGND_c_718_n N_VGND_c_719_n
+ N_VGND_c_720_n N_VGND_c_721_n N_VGND_c_722_n N_VGND_c_723_n VGND
+ N_VGND_c_724_n N_VGND_c_725_n N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n
+ N_VGND_c_729_n N_VGND_c_730_n N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n
+ PM_SKY130_FD_SC_LP__O21BA_4%VGND
x_PM_SKY130_FD_SC_LP__O21BA_4%A_575_65# N_A_575_65#_M1001_d N_A_575_65#_M1013_d
+ N_A_575_65#_M1012_d N_A_575_65#_M1008_s N_A_575_65#_c_810_n
+ N_A_575_65#_c_811_n N_A_575_65#_c_812_n N_A_575_65#_c_831_n
+ N_A_575_65#_c_825_n N_A_575_65#_c_826_n N_A_575_65#_c_813_n
+ N_A_575_65#_c_814_n N_A_575_65#_c_815_n N_A_575_65#_c_816_n
+ PM_SKY130_FD_SC_LP__O21BA_4%A_575_65#
cc_1 VNB N_B1_N_M1021_g 0.00660273f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_2 VNB B1_N 0.00766261f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_B1_N_c_108_n 0.0328405f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_4 VNB N_B1_N_c_109_n 0.0202952f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.21
cc_5 VNB N_A_180_23#_M1007_g 0.0228072f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_6 VNB N_A_180_23#_M1009_g 0.0222179f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.375
cc_7 VNB N_A_180_23#_M1016_g 0.022218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_180_23#_M1019_g 0.0283972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_180_23#_c_146_n 0.00336366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_180_23#_c_147_n 0.00407508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_180_23#_c_148_n 0.0165233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_180_23#_c_149_n 0.0077358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_180_23#_c_150_n 0.0114885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_180_23#_c_151_n 0.00308487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_180_23#_c_152_n 0.00496144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_180_23#_c_153_n 0.0684579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_37_49#_M1001_g 0.0302795f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_18 VNB N_A_37_49#_M1013_g 0.0292372f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.665
cc_19 VNB N_A_37_49#_c_306_n 0.025525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_37_49#_c_307_n 0.00698135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_37_49#_c_308_n 0.0293488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_37_49#_c_309_n 0.0491041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_M1005_g 0.0217089f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.665
cc_24 VNB N_A1_M1008_g 0.0264027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_406_n 3.30444e-19 $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.375
cc_26 VNB N_A1_c_407_n 0.0290269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_c_408_n 0.01135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_c_409_n 0.0303307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A2_M1012_g 0.0200032f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.665
cc_30 VNB N_A2_M1017_g 0.019334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_493_n 0.0316395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_550_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_652_n 9.24575e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_653_n 0.00678648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_654_n 0.00221538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_717_n 0.00207168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_718_n 4.87379e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_719_n 0.00958534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_720_n 0.00457468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_721_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_722_n 0.0136175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_723_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_724_n 0.0169166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_725_n 0.0152764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_726_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_727_n 0.0412821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_728_n 0.0212006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_729_n 0.337667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_730_n 0.00405272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_731_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_732_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_733_n 0.00598106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_575_65#_c_810_n 0.00446679f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.21
cc_54 VNB N_A_575_65#_c_811_n 0.00499546f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.295
cc_55 VNB N_A_575_65#_c_812_n 0.00440562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_575_65#_c_813_n 0.00199404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_575_65#_c_814_n 0.0184343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_575_65#_c_815_n 0.00348245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_575_65#_c_816_n 0.0314832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_B1_N_M1021_g 0.0235919f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_61 VPB B1_N 0.00554383f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_62 VPB N_A_180_23#_M1000_g 0.018119f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.54
cc_63 VPB N_A_180_23#_M1002_g 0.0185698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_180_23#_M1003_g 0.0186308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_180_23#_M1018_g 0.0216707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_180_23#_c_149_n 0.00238441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_180_23#_c_151_n 0.00108414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_180_23#_c_153_n 0.0119819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_37_49#_M1006_g 0.0218637f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_70 VPB N_A_37_49#_M1011_g 0.0214162f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=1.295
cc_71 VPB N_A_37_49#_c_312_n 0.0141071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_37_49#_c_313_n 0.0214801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_37_49#_c_314_n 0.00518283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_37_49#_c_315_n 0.0026966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_37_49#_c_316_n 0.00807991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_37_49#_c_308_n 0.0124997f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_37_49#_c_318_n 0.00839616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_37_49#_c_309_n 0.0209299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A1_M1010_g 0.0208346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A1_M1014_g 0.0249722f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.21
cc_81 VPB N_A1_c_412_n 0.00177491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A1_c_406_n 0.001379f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=1.375
cc_83 VPB N_A1_c_414_n 0.00213753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A1_c_407_n 0.00792334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A1_c_409_n 0.00888411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A2_M1004_g 0.0181061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A2_M1015_g 0.018675f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.21
cc_88 VPB N_A2_c_496_n 0.00221113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A2_c_493_n 0.00471591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_551_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_552_n 3.09829e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_553_n 0.00352082f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_554_n 0.0138419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_555_n 0.0562307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_556_n 0.0171007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_557_n 0.0127282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_558_n 0.0383402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_559_n 0.00436638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_560_n 0.00436638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_561_n 0.0128627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_562_n 0.01576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_563_n 0.0134123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_564_n 0.0123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_550_n 0.0500993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_X_c_652_n 0.00153052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 B1_N N_A_180_23#_M1007_g 0.00228708f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B1_N_c_108_n N_A_180_23#_M1007_g 0.0176567f $X=0.525 $Y=1.375 $X2=0
+ $Y2=0
cc_108 N_B1_N_c_109_n N_A_180_23#_M1007_g 0.0159839f $X=0.525 $Y=1.21 $X2=0
+ $Y2=0
cc_109 N_B1_N_M1021_g N_A_180_23#_c_153_n 0.05791f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_110 B1_N N_A_180_23#_c_153_n 0.00215674f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_N_c_108_n N_A_180_23#_c_153_n 0.00235053f $X=0.525 $Y=1.375 $X2=0
+ $Y2=0
cc_112 N_B1_N_M1021_g N_A_37_49#_c_320_n 0.0135806f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_B1_N_c_108_n N_A_37_49#_c_307_n 0.00255043f $X=0.525 $Y=1.375 $X2=0
+ $Y2=0
cc_114 B1_N N_A_37_49#_c_316_n 0.00203547f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B1_N_c_108_n N_A_37_49#_c_316_n 0.00263571f $X=0.525 $Y=1.375 $X2=0
+ $Y2=0
cc_116 N_B1_N_M1021_g N_A_37_49#_c_308_n 0.00499797f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_117 B1_N N_A_37_49#_c_308_n 0.0432568f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B1_N_c_108_n N_A_37_49#_c_308_n 0.00804249f $X=0.525 $Y=1.375 $X2=0
+ $Y2=0
cc_119 N_B1_N_c_109_n N_A_37_49#_c_308_n 0.00400834f $X=0.525 $Y=1.21 $X2=0
+ $Y2=0
cc_120 N_B1_N_M1021_g N_VPWR_c_551_n 0.00893583f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_121 N_B1_N_M1021_g N_VPWR_c_556_n 0.0036352f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_122 N_B1_N_M1021_g N_VPWR_c_550_n 0.00531256f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B1_N_c_109_n N_X_c_656_n 4.0238e-19 $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B1_N_M1021_g N_X_c_652_n 0.00105114f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_125 B1_N N_X_c_652_n 0.0389198f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B1_N_c_108_n N_X_c_652_n 2.22053e-19 $X=0.525 $Y=1.375 $X2=0 $Y2=0
cc_127 B1_N N_X_c_654_n 0.00385581f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B1_N_c_109_n N_X_c_654_n 5.99596e-19 $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B1_N_M1021_g N_X_c_662_n 0.00880701f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_130 B1_N N_X_c_662_n 0.0179193f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_131 B1_N N_VGND_c_717_n 0.0205126f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_N_c_108_n N_VGND_c_717_n 3.65529e-19 $X=0.525 $Y=1.375 $X2=0 $Y2=0
cc_133 N_B1_N_c_109_n N_VGND_c_717_n 0.0142813f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B1_N_c_109_n N_VGND_c_724_n 0.00477554f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_135 N_B1_N_c_109_n N_VGND_c_729_n 0.00925056f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A_180_23#_M1018_g N_A_37_49#_M1006_g 0.00916149f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_180_23#_c_149_n N_A_37_49#_M1006_g 0.00200976f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_138 N_A_180_23#_c_149_n N_A_37_49#_M1001_g 0.00691205f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_139 N_A_180_23#_c_170_p N_A_37_49#_M1001_g 0.0108489f $X=3.51 $Y=0.69 $X2=0
+ $Y2=0
cc_140 N_A_180_23#_c_152_n N_A_37_49#_M1001_g 0.0111914f $X=3.44 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_180_23#_c_149_n N_A_37_49#_M1011_g 0.00269134f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_142 N_A_180_23#_c_149_n N_A_37_49#_M1013_g 0.00445062f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_143 N_A_180_23#_c_170_p N_A_37_49#_M1013_g 0.00684135f $X=3.51 $Y=0.69 $X2=0
+ $Y2=0
cc_144 N_A_180_23#_c_150_n N_A_37_49#_M1013_g 0.0107395f $X=4.525 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_180_23#_c_152_n N_A_37_49#_M1013_g 0.00189414f $X=3.44 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_180_23#_M1000_g N_A_37_49#_c_320_n 0.0122351f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_180_23#_M1002_g N_A_37_49#_c_320_n 0.0123328f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_180_23#_M1003_g N_A_37_49#_c_320_n 0.0123415f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_180_23#_M1018_g N_A_37_49#_c_320_n 0.0168388f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_180_23#_M1018_g N_A_37_49#_c_314_n 0.00300352f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_180_23#_c_146_n N_A_37_49#_c_314_n 0.00496468f $X=2.315 $Y=1.51 $X2=0
+ $Y2=0
cc_152 N_A_180_23#_c_148_n N_A_37_49#_c_314_n 0.00673108f $X=3.205 $Y=1.16 $X2=0
+ $Y2=0
cc_153 N_A_180_23#_c_149_n N_A_37_49#_c_314_n 0.00446611f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_154 N_A_180_23#_M1018_g N_A_37_49#_c_315_n 0.00230602f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_180_23#_c_146_n N_A_37_49#_c_315_n 0.0144545f $X=2.315 $Y=1.51 $X2=0
+ $Y2=0
cc_156 N_A_180_23#_c_148_n N_A_37_49#_c_315_n 0.0249357f $X=3.205 $Y=1.16 $X2=0
+ $Y2=0
cc_157 N_A_180_23#_c_149_n N_A_37_49#_c_315_n 0.0247179f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_158 N_A_180_23#_c_153_n N_A_37_49#_c_315_n 7.1999e-19 $X=2.265 $Y=1.51 $X2=0
+ $Y2=0
cc_159 N_A_180_23#_c_146_n N_A_37_49#_c_309_n 0.00144751f $X=2.315 $Y=1.51 $X2=0
+ $Y2=0
cc_160 N_A_180_23#_c_147_n N_A_37_49#_c_309_n 0.00144392f $X=2.4 $Y=1.415 $X2=0
+ $Y2=0
cc_161 N_A_180_23#_c_148_n N_A_37_49#_c_309_n 0.0150264f $X=3.205 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A_180_23#_c_149_n N_A_37_49#_c_309_n 0.0133805f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_163 N_A_180_23#_c_152_n N_A_37_49#_c_309_n 0.00424403f $X=3.44 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A_180_23#_c_153_n N_A_37_49#_c_309_n 0.0144662f $X=2.265 $Y=1.51 $X2=0
+ $Y2=0
cc_165 N_A_180_23#_c_170_p N_A1_M1005_g 5.84315e-19 $X=3.51 $Y=0.69 $X2=0 $Y2=0
cc_166 N_A_180_23#_c_150_n N_A1_M1005_g 0.0113093f $X=4.525 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_180_23#_c_151_n N_A1_M1005_g 0.00201402f $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_168 N_A_180_23#_c_199_p N_A1_M1010_g 0.00144758f $X=4.695 $Y=2.035 $X2=0
+ $Y2=0
cc_169 N_A_180_23#_c_149_n N_A1_c_412_n 0.00430271f $X=3.33 $Y=1.98 $X2=0 $Y2=0
cc_170 N_A_180_23#_c_199_p N_A1_c_412_n 0.0161971f $X=4.695 $Y=2.035 $X2=0 $Y2=0
cc_171 N_A_180_23#_c_202_p N_A1_c_406_n 0.0101711f $X=4.96 $Y=2.035 $X2=0 $Y2=0
cc_172 N_A_180_23#_c_149_n N_A1_c_414_n 0.00717088f $X=3.33 $Y=1.98 $X2=0 $Y2=0
cc_173 N_A_180_23#_c_150_n N_A1_c_414_n 0.0253118f $X=4.525 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_180_23#_c_151_n N_A1_c_414_n 0.0365981f $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_175 N_A_180_23#_c_149_n N_A1_c_407_n 3.11596e-19 $X=3.33 $Y=1.98 $X2=0 $Y2=0
cc_176 N_A_180_23#_c_150_n N_A1_c_407_n 0.00657789f $X=4.525 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_180_23#_c_151_n N_A1_c_407_n 0.00490004f $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_178 N_A_180_23#_M1004_d A1 0.0034413f $X=4.82 $Y=1.835 $X2=0 $Y2=0
cc_179 N_A_180_23#_c_199_p A1 0.00904562f $X=4.695 $Y=2.035 $X2=0 $Y2=0
cc_180 N_A_180_23#_c_202_p A1 0.0226703f $X=4.96 $Y=2.035 $X2=0 $Y2=0
cc_181 N_A_180_23#_c_150_n N_A2_M1012_g 0.00449664f $X=4.525 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_180_23#_c_151_n N_A2_M1012_g 0.00256346f $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_183 N_A_180_23#_c_151_n N_A2_M1004_g 0.00570342f $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_184 N_A_180_23#_c_199_p N_A2_M1004_g 0.00237488f $X=4.695 $Y=2.035 $X2=0
+ $Y2=0
cc_185 N_A_180_23#_c_202_p N_A2_M1004_g 0.00968336f $X=4.96 $Y=2.035 $X2=0 $Y2=0
cc_186 N_A_180_23#_c_151_n N_A2_M1017_g 4.8453e-19 $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_187 N_A_180_23#_c_151_n N_A2_M1015_g 7.09042e-19 $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_188 N_A_180_23#_c_202_p N_A2_M1015_g 0.00342994f $X=4.96 $Y=2.035 $X2=0 $Y2=0
cc_189 N_A_180_23#_c_151_n N_A2_c_496_n 0.0200214f $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_190 N_A_180_23#_c_202_p N_A2_c_496_n 0.0139282f $X=4.96 $Y=2.035 $X2=0 $Y2=0
cc_191 N_A_180_23#_c_151_n N_A2_c_493_n 0.0102247f $X=4.61 $Y=1.93 $X2=0 $Y2=0
cc_192 N_A_180_23#_c_202_p N_A2_c_493_n 8.95773e-19 $X=4.96 $Y=2.035 $X2=0 $Y2=0
cc_193 N_A_180_23#_M1000_g N_VPWR_c_551_n 0.00949711f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A_180_23#_M1002_g N_VPWR_c_551_n 0.00135454f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_180_23#_M1000_g N_VPWR_c_552_n 0.00135454f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A_180_23#_M1002_g N_VPWR_c_552_n 0.00955913f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A_180_23#_M1003_g N_VPWR_c_552_n 0.00925656f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_180_23#_M1018_g N_VPWR_c_552_n 0.00134502f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_180_23#_M1018_g N_VPWR_c_575_n 0.00428213f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_180_23#_c_149_n N_VPWR_c_553_n 0.0367933f $X=3.33 $Y=1.98 $X2=0 $Y2=0
cc_201 N_A_180_23#_c_150_n N_VPWR_c_553_n 0.00781783f $X=4.525 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_180_23#_c_152_n N_VPWR_c_553_n 0.00292707f $X=3.44 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_A_180_23#_M1000_g N_VPWR_c_557_n 0.0036352f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_180_23#_M1002_g N_VPWR_c_557_n 0.0036352f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_A_180_23#_M1003_g N_VPWR_c_561_n 0.00378092f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_206 N_A_180_23#_M1018_g N_VPWR_c_561_n 0.0036352f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_207 N_A_180_23#_M1003_g N_VPWR_c_562_n 0.00137082f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_208 N_A_180_23#_M1018_g N_VPWR_c_562_n 0.0105717f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_A_180_23#_c_149_n N_VPWR_c_563_n 0.0135169f $X=3.33 $Y=1.98 $X2=0 $Y2=0
cc_210 N_A_180_23#_M1006_d N_VPWR_c_550_n 0.00432284f $X=3.19 $Y=1.835 $X2=0
+ $Y2=0
cc_211 N_A_180_23#_M1004_d N_VPWR_c_550_n 0.00231436f $X=4.82 $Y=1.835 $X2=0
+ $Y2=0
cc_212 N_A_180_23#_M1000_g N_VPWR_c_550_n 0.00436741f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_213 N_A_180_23#_M1002_g N_VPWR_c_550_n 0.00436741f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_214 N_A_180_23#_M1003_g N_VPWR_c_550_n 0.00451808f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_A_180_23#_M1018_g N_VPWR_c_550_n 0.00435022f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_A_180_23#_c_149_n N_VPWR_c_550_n 0.00847534f $X=3.33 $Y=1.98 $X2=0
+ $Y2=0
cc_217 N_A_180_23#_M1007_g N_X_c_656_n 0.00936928f $X=0.975 $Y=0.665 $X2=0 $Y2=0
cc_218 N_A_180_23#_M1007_g N_X_c_652_n 0.00165615f $X=0.975 $Y=0.665 $X2=0 $Y2=0
cc_219 N_A_180_23#_M1000_g N_X_c_652_n 0.00564371f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A_180_23#_M1009_g N_X_c_652_n 0.00216385f $X=1.405 $Y=0.665 $X2=0 $Y2=0
cc_221 N_A_180_23#_M1002_g N_X_c_652_n 0.00500925f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A_180_23#_c_146_n N_X_c_652_n 0.014321f $X=2.315 $Y=1.51 $X2=0 $Y2=0
cc_223 N_A_180_23#_c_153_n N_X_c_652_n 0.0187124f $X=2.265 $Y=1.51 $X2=0 $Y2=0
cc_224 N_A_180_23#_M1009_g N_X_c_653_n 0.0155031f $X=1.405 $Y=0.665 $X2=0 $Y2=0
cc_225 N_A_180_23#_M1016_g N_X_c_653_n 0.0137525f $X=1.835 $Y=0.665 $X2=0 $Y2=0
cc_226 N_A_180_23#_M1019_g N_X_c_653_n 0.00131247f $X=2.265 $Y=0.665 $X2=0 $Y2=0
cc_227 N_A_180_23#_c_146_n N_X_c_653_n 0.0562767f $X=2.315 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_180_23#_c_259_p N_X_c_653_n 0.0146391f $X=2.485 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_180_23#_c_153_n N_X_c_653_n 0.00533319f $X=2.265 $Y=1.51 $X2=0 $Y2=0
cc_230 N_A_180_23#_M1007_g N_X_c_654_n 0.00471564f $X=0.975 $Y=0.665 $X2=0 $Y2=0
cc_231 N_A_180_23#_c_153_n N_X_c_654_n 0.00167841f $X=2.265 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A_180_23#_M1000_g X 0.00249715f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A_180_23#_M1002_g X 0.0135872f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A_180_23#_M1003_g X 0.0136674f $X=1.88 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A_180_23#_M1018_g X 0.00403534f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_180_23#_c_146_n X 0.0334397f $X=2.315 $Y=1.51 $X2=0 $Y2=0
cc_237 N_A_180_23#_c_153_n X 0.00780087f $X=2.265 $Y=1.51 $X2=0 $Y2=0
cc_238 N_A_180_23#_M1000_g N_X_c_662_n 0.0127656f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A_180_23#_c_151_n N_A_878_367#_M1010_s 7.95042e-19 $X=4.61 $Y=1.93
+ $X2=-0.19 $Y2=-0.245
cc_240 N_A_180_23#_c_199_p N_A_878_367#_M1010_s 0.0027899f $X=4.695 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_241 N_A_180_23#_M1004_d N_A_878_367#_c_705_n 0.00366227f $X=4.82 $Y=1.835
+ $X2=0 $Y2=0
cc_242 N_A_180_23#_c_148_n N_VGND_M1019_d 0.00130734f $X=3.205 $Y=1.16 $X2=0
+ $Y2=0
cc_243 N_A_180_23#_c_259_p N_VGND_M1019_d 9.66455e-19 $X=2.485 $Y=1.16 $X2=0
+ $Y2=0
cc_244 N_A_180_23#_c_150_n N_VGND_M1005_d 0.00271357f $X=4.525 $Y=1.16 $X2=0
+ $Y2=0
cc_245 N_A_180_23#_M1007_g N_VGND_c_717_n 0.0018556f $X=0.975 $Y=0.665 $X2=0
+ $Y2=0
cc_246 N_A_180_23#_M1007_g N_VGND_c_718_n 6.97314e-19 $X=0.975 $Y=0.665 $X2=0
+ $Y2=0
cc_247 N_A_180_23#_M1009_g N_VGND_c_718_n 0.0113679f $X=1.405 $Y=0.665 $X2=0
+ $Y2=0
cc_248 N_A_180_23#_M1016_g N_VGND_c_718_n 0.0112407f $X=1.835 $Y=0.665 $X2=0
+ $Y2=0
cc_249 N_A_180_23#_M1019_g N_VGND_c_718_n 6.15775e-19 $X=2.265 $Y=0.665 $X2=0
+ $Y2=0
cc_250 N_A_180_23#_M1016_g N_VGND_c_719_n 6.15775e-19 $X=1.835 $Y=0.665 $X2=0
+ $Y2=0
cc_251 N_A_180_23#_M1019_g N_VGND_c_719_n 0.0126329f $X=2.265 $Y=0.665 $X2=0
+ $Y2=0
cc_252 N_A_180_23#_c_148_n N_VGND_c_719_n 0.0130205f $X=3.205 $Y=1.16 $X2=0
+ $Y2=0
cc_253 N_A_180_23#_c_259_p N_VGND_c_719_n 0.00974177f $X=2.485 $Y=1.16 $X2=0
+ $Y2=0
cc_254 N_A_180_23#_M1007_g N_VGND_c_725_n 0.00554241f $X=0.975 $Y=0.665 $X2=0
+ $Y2=0
cc_255 N_A_180_23#_M1009_g N_VGND_c_725_n 0.00477554f $X=1.405 $Y=0.665 $X2=0
+ $Y2=0
cc_256 N_A_180_23#_M1016_g N_VGND_c_726_n 0.00477554f $X=1.835 $Y=0.665 $X2=0
+ $Y2=0
cc_257 N_A_180_23#_M1019_g N_VGND_c_726_n 0.00477554f $X=2.265 $Y=0.665 $X2=0
+ $Y2=0
cc_258 N_A_180_23#_M1007_g N_VGND_c_729_n 0.0101473f $X=0.975 $Y=0.665 $X2=0
+ $Y2=0
cc_259 N_A_180_23#_M1009_g N_VGND_c_729_n 0.00825815f $X=1.405 $Y=0.665 $X2=0
+ $Y2=0
cc_260 N_A_180_23#_M1016_g N_VGND_c_729_n 0.00825815f $X=1.835 $Y=0.665 $X2=0
+ $Y2=0
cc_261 N_A_180_23#_M1019_g N_VGND_c_729_n 0.00825815f $X=2.265 $Y=0.665 $X2=0
+ $Y2=0
cc_262 N_A_180_23#_c_148_n N_A_575_65#_M1001_d 0.00387431f $X=3.205 $Y=1.16
+ $X2=-0.19 $Y2=-0.245
cc_263 N_A_180_23#_c_150_n N_A_575_65#_M1013_d 0.00267852f $X=4.525 $Y=1.16
+ $X2=0 $Y2=0
cc_264 N_A_180_23#_M1019_g N_A_575_65#_c_810_n 8.28231e-19 $X=2.265 $Y=0.665
+ $X2=0 $Y2=0
cc_265 N_A_180_23#_c_148_n N_A_575_65#_c_810_n 0.0265929f $X=3.205 $Y=1.16 $X2=0
+ $Y2=0
cc_266 N_A_180_23#_M1001_s N_A_575_65#_c_811_n 0.00176461f $X=3.37 $Y=0.325
+ $X2=0 $Y2=0
cc_267 N_A_180_23#_c_170_p N_A_575_65#_c_811_n 0.0159477f $X=3.51 $Y=0.69 $X2=0
+ $Y2=0
cc_268 N_A_180_23#_c_150_n N_A_575_65#_c_811_n 0.00280043f $X=4.525 $Y=1.16
+ $X2=0 $Y2=0
cc_269 N_A_180_23#_c_152_n N_A_575_65#_c_811_n 0.00314961f $X=3.44 $Y=1.16 $X2=0
+ $Y2=0
cc_270 N_A_180_23#_c_150_n N_A_575_65#_c_825_n 0.0276627f $X=4.525 $Y=1.16 $X2=0
+ $Y2=0
cc_271 N_A_180_23#_c_150_n N_A_575_65#_c_826_n 0.0208246f $X=4.525 $Y=1.16 $X2=0
+ $Y2=0
cc_272 N_A_180_23#_c_150_n N_A_575_65#_c_815_n 0.0108938f $X=4.525 $Y=1.16 $X2=0
+ $Y2=0
cc_273 N_A_37_49#_M1013_g N_A1_M1005_g 0.0260861f $X=3.725 $Y=0.745 $X2=0 $Y2=0
cc_274 N_A_37_49#_M1011_g N_A1_M1010_g 0.0105981f $X=3.545 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A_37_49#_M1011_g N_A1_c_412_n 0.00199233f $X=3.545 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A_37_49#_M1013_g N_A1_c_414_n 0.00117416f $X=3.725 $Y=0.745 $X2=0 $Y2=0
cc_277 N_A_37_49#_M1013_g N_A1_c_407_n 0.0214077f $X=3.725 $Y=0.745 $X2=0 $Y2=0
cc_278 N_A_37_49#_c_320_n N_VPWR_M1021_d 0.00349458f $X=2.425 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_279 N_A_37_49#_c_320_n N_VPWR_M1002_d 0.00359984f $X=2.425 $Y=2.52 $X2=0
+ $Y2=0
cc_280 N_A_37_49#_c_320_n N_VPWR_M1018_d 0.00368278f $X=2.425 $Y=2.52 $X2=0
+ $Y2=0
cc_281 N_A_37_49#_c_365_p N_VPWR_M1018_d 0.00899101f $X=2.51 $Y=2.43 $X2=0 $Y2=0
cc_282 N_A_37_49#_c_314_n N_VPWR_M1018_d 0.0120493f $X=2.845 $Y=1.775 $X2=0
+ $Y2=0
cc_283 N_A_37_49#_c_320_n N_VPWR_c_551_n 0.0164573f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_284 N_A_37_49#_c_320_n N_VPWR_c_552_n 0.0164823f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_285 N_A_37_49#_c_320_n N_VPWR_c_575_n 0.0151154f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_286 N_A_37_49#_c_365_p N_VPWR_c_575_n 0.0236636f $X=2.51 $Y=2.43 $X2=0 $Y2=0
cc_287 N_A_37_49#_c_314_n N_VPWR_c_575_n 0.0176226f $X=2.845 $Y=1.775 $X2=0
+ $Y2=0
cc_288 N_A_37_49#_M1011_g N_VPWR_c_553_n 0.0138771f $X=3.545 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_37_49#_c_309_n N_VPWR_c_553_n 0.00616535f $X=3.545 $Y=1.525 $X2=0
+ $Y2=0
cc_290 N_A_37_49#_c_313_n N_VPWR_c_556_n 0.0264135f $X=0.37 $Y=2.91 $X2=0 $Y2=0
cc_291 N_A_37_49#_c_320_n N_VPWR_c_556_n 0.0020344f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_292 N_A_37_49#_c_320_n N_VPWR_c_557_n 0.00670101f $X=2.425 $Y=2.52 $X2=0
+ $Y2=0
cc_293 N_A_37_49#_c_320_n N_VPWR_c_561_n 0.00676879f $X=2.425 $Y=2.52 $X2=0
+ $Y2=0
cc_294 N_A_37_49#_M1006_g N_VPWR_c_562_n 0.00226909f $X=3.115 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_37_49#_c_320_n N_VPWR_c_562_n 0.0148987f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_296 N_A_37_49#_M1006_g N_VPWR_c_563_n 0.00409769f $X=3.115 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A_37_49#_M1011_g N_VPWR_c_563_n 0.00292692f $X=3.545 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A_37_49#_M1006_g N_VPWR_c_564_n 5.6037e-19 $X=3.115 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_A_37_49#_M1011_g N_VPWR_c_564_n 0.00807111f $X=3.545 $Y=2.465 $X2=0
+ $Y2=0
cc_300 N_A_37_49#_M1021_s N_VPWR_c_550_n 0.00235632f $X=0.245 $Y=1.835 $X2=0
+ $Y2=0
cc_301 N_A_37_49#_M1006_g N_VPWR_c_550_n 0.0111916f $X=3.115 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_37_49#_M1011_g N_VPWR_c_550_n 0.00819843f $X=3.545 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_37_49#_c_313_n N_VPWR_c_550_n 0.0146953f $X=0.37 $Y=2.91 $X2=0 $Y2=0
cc_304 N_A_37_49#_c_320_n N_VPWR_c_550_n 0.0335359f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_305 N_A_37_49#_c_320_n N_X_M1000_s 0.00493329f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_306 N_A_37_49#_c_320_n N_X_M1003_s 0.00494544f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_307 N_A_37_49#_c_320_n X 0.00881408f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_308 N_A_37_49#_c_320_n X 0.0569421f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_309 N_A_37_49#_c_320_n N_X_c_662_n 0.0220749f $X=2.425 $Y=2.52 $X2=0 $Y2=0
cc_310 N_A_37_49#_M1001_g N_VGND_c_719_n 0.00241388f $X=3.295 $Y=0.745 $X2=0
+ $Y2=0
cc_311 N_A_37_49#_c_306_n N_VGND_c_724_n 0.0235185f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_312 N_A_37_49#_M1001_g N_VGND_c_727_n 0.0030414f $X=3.295 $Y=0.745 $X2=0
+ $Y2=0
cc_313 N_A_37_49#_M1013_g N_VGND_c_727_n 0.0030414f $X=3.725 $Y=0.745 $X2=0
+ $Y2=0
cc_314 N_A_37_49#_M1020_s N_VGND_c_729_n 0.00384928f $X=0.185 $Y=0.245 $X2=0
+ $Y2=0
cc_315 N_A_37_49#_M1001_g N_VGND_c_729_n 0.00484828f $X=3.295 $Y=0.745 $X2=0
+ $Y2=0
cc_316 N_A_37_49#_M1013_g N_VGND_c_729_n 0.0044277f $X=3.725 $Y=0.745 $X2=0
+ $Y2=0
cc_317 N_A_37_49#_c_306_n N_VGND_c_729_n 0.0131407f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_318 N_A_37_49#_M1001_g N_A_575_65#_c_811_n 0.012837f $X=3.295 $Y=0.745 $X2=0
+ $Y2=0
cc_319 N_A_37_49#_M1013_g N_A_575_65#_c_811_n 0.0116477f $X=3.725 $Y=0.745 $X2=0
+ $Y2=0
cc_320 N_A1_M1005_g N_A2_M1012_g 0.0309308f $X=4.235 $Y=0.745 $X2=0 $Y2=0
cc_321 N_A1_M1010_g N_A2_M1004_g 0.0329315f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A1_c_412_n N_A2_M1004_g 0.00130889f $X=4.21 $Y=2.31 $X2=0 $Y2=0
cc_323 A1 N_A2_M1004_g 0.0111997f $X=5.435 $Y=2.32 $X2=0 $Y2=0
cc_324 N_A1_M1008_g N_A2_M1017_g 0.0291586f $X=5.605 $Y=0.745 $X2=0 $Y2=0
cc_325 N_A1_M1014_g N_A2_M1015_g 0.0291586f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_326 A1 N_A2_M1015_g 0.0127275f $X=5.435 $Y=2.32 $X2=0 $Y2=0
cc_327 N_A1_c_406_n N_A2_c_496_n 0.00807486f $X=5.52 $Y=2.31 $X2=0 $Y2=0
cc_328 N_A1_c_408_n N_A2_c_496_n 0.0173597f $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_329 N_A1_c_409_n N_A2_c_496_n 3.71357e-19 $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_330 A1 N_A2_c_496_n 0.00342405f $X=5.435 $Y=2.32 $X2=0 $Y2=0
cc_331 N_A1_c_406_n N_A2_c_493_n 0.00903169f $X=5.52 $Y=2.31 $X2=0 $Y2=0
cc_332 N_A1_c_414_n N_A2_c_493_n 3.40434e-19 $X=4.18 $Y=1.51 $X2=0 $Y2=0
cc_333 N_A1_c_407_n N_A2_c_493_n 0.0329315f $X=4.18 $Y=1.51 $X2=0 $Y2=0
cc_334 N_A1_c_408_n N_A2_c_493_n 0.00165546f $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_335 N_A1_c_409_n N_A2_c_493_n 0.0291586f $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_336 N_A1_c_412_n N_VPWR_M1011_s 0.00448632f $X=4.21 $Y=2.31 $X2=0 $Y2=0
cc_337 N_A1_c_455_p N_VPWR_M1011_s 0.00332013f $X=4.345 $Y=2.405 $X2=0 $Y2=0
cc_338 N_A1_M1010_g N_VPWR_c_553_n 0.00668172f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A1_c_412_n N_VPWR_c_553_n 0.0389542f $X=4.21 $Y=2.31 $X2=0 $Y2=0
cc_340 N_A1_c_455_p N_VPWR_c_553_n 0.01611f $X=4.345 $Y=2.405 $X2=0 $Y2=0
cc_341 N_A1_M1014_g N_VPWR_c_555_n 0.0167582f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_342 N_A1_c_406_n N_VPWR_c_555_n 0.0511604f $X=5.52 $Y=2.31 $X2=0 $Y2=0
cc_343 N_A1_c_408_n N_VPWR_c_555_n 0.00691319f $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_344 N_A1_c_409_n N_VPWR_c_555_n 0.00202893f $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_345 N_A1_M1010_g N_VPWR_c_558_n 0.00486043f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_346 N_A1_M1014_g N_VPWR_c_558_n 0.00585385f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A1_M1010_g N_VPWR_c_564_n 0.010327f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_348 N_A1_c_455_p N_VPWR_c_564_n 0.00723265f $X=4.345 $Y=2.405 $X2=0 $Y2=0
cc_349 N_A1_M1010_g N_VPWR_c_550_n 0.00460532f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_350 N_A1_M1014_g N_VPWR_c_550_n 0.00970523f $X=5.605 $Y=2.465 $X2=0 $Y2=0
cc_351 N_A1_c_406_n N_VPWR_c_550_n 0.00389047f $X=5.52 $Y=2.31 $X2=0 $Y2=0
cc_352 N_A1_c_455_p N_VPWR_c_550_n 0.00345527f $X=4.345 $Y=2.405 $X2=0 $Y2=0
cc_353 A1 N_VPWR_c_550_n 0.00419895f $X=5.435 $Y=2.32 $X2=0 $Y2=0
cc_354 A1 N_A_878_367#_M1010_s 0.00569401f $X=5.435 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_355 N_A1_c_406_n N_A_878_367#_M1015_s 0.00575453f $X=5.52 $Y=2.31 $X2=0 $Y2=0
cc_356 A1 N_A_878_367#_M1015_s 0.00624995f $X=5.435 $Y=2.32 $X2=0 $Y2=0
cc_357 N_A1_c_406_n N_A_878_367#_c_705_n 0.00310671f $X=5.52 $Y=2.31 $X2=0 $Y2=0
cc_358 A1 N_A_878_367#_c_705_n 0.0554799f $X=5.435 $Y=2.32 $X2=0 $Y2=0
cc_359 N_A1_M1005_g N_VGND_c_720_n 0.00347453f $X=4.235 $Y=0.745 $X2=0 $Y2=0
cc_360 N_A1_M1008_g N_VGND_c_721_n 0.0125458f $X=5.605 $Y=0.745 $X2=0 $Y2=0
cc_361 N_A1_M1005_g N_VGND_c_727_n 0.00356071f $X=4.235 $Y=0.745 $X2=0 $Y2=0
cc_362 N_A1_M1008_g N_VGND_c_728_n 0.00414769f $X=5.605 $Y=0.745 $X2=0 $Y2=0
cc_363 N_A1_M1005_g N_VGND_c_729_n 0.00507138f $X=4.235 $Y=0.745 $X2=0 $Y2=0
cc_364 N_A1_M1008_g N_VGND_c_729_n 0.00827997f $X=5.605 $Y=0.745 $X2=0 $Y2=0
cc_365 N_A1_M1005_g N_A_575_65#_c_811_n 0.00276118f $X=4.235 $Y=0.745 $X2=0
+ $Y2=0
cc_366 N_A1_M1005_g N_A_575_65#_c_831_n 0.00450492f $X=4.235 $Y=0.745 $X2=0
+ $Y2=0
cc_367 N_A1_M1005_g N_A_575_65#_c_825_n 0.00915996f $X=4.235 $Y=0.745 $X2=0
+ $Y2=0
cc_368 N_A1_M1005_g N_A_575_65#_c_826_n 7.41384e-19 $X=4.235 $Y=0.745 $X2=0
+ $Y2=0
cc_369 N_A1_M1008_g N_A_575_65#_c_814_n 0.0138332f $X=5.605 $Y=0.745 $X2=0 $Y2=0
cc_370 N_A1_c_408_n N_A_575_65#_c_814_n 0.0320019f $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_371 N_A1_c_409_n N_A_575_65#_c_814_n 0.0045072f $X=5.695 $Y=1.51 $X2=0 $Y2=0
cc_372 N_A1_M1008_g N_A_575_65#_c_816_n 0.00350978f $X=5.605 $Y=0.745 $X2=0
+ $Y2=0
cc_373 N_A2_M1004_g N_VPWR_c_558_n 0.00373071f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A2_M1015_g N_VPWR_c_558_n 0.00373071f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_375 N_A2_M1004_g N_VPWR_c_564_n 0.00149029f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A2_M1004_g N_VPWR_c_550_n 0.00548684f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_377 N_A2_M1015_g N_VPWR_c_550_n 0.00548684f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_378 N_A2_M1004_g N_A_878_367#_c_705_n 0.0122888f $X=4.745 $Y=2.465 $X2=0
+ $Y2=0
cc_379 N_A2_M1015_g N_A_878_367#_c_705_n 0.0123029f $X=5.175 $Y=2.465 $X2=0
+ $Y2=0
cc_380 N_A2_M1012_g N_VGND_c_720_n 0.00656395f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_381 N_A2_M1017_g N_VGND_c_720_n 3.84006e-19 $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_382 N_A2_M1012_g N_VGND_c_721_n 5.26603e-19 $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_383 N_A2_M1017_g N_VGND_c_721_n 0.00999226f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_384 N_A2_M1012_g N_VGND_c_722_n 0.00304778f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_385 N_A2_M1017_g N_VGND_c_722_n 0.00414769f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_386 N_A2_M1012_g N_VGND_c_729_n 0.00389787f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_387 N_A2_M1017_g N_VGND_c_729_n 0.00787505f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_388 N_A2_M1012_g N_A_575_65#_c_831_n 5.8454e-19 $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_389 N_A2_M1012_g N_A_575_65#_c_825_n 0.0149062f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_390 N_A2_M1012_g N_A_575_65#_c_813_n 5.14142e-19 $X=4.745 $Y=0.745 $X2=0
+ $Y2=0
cc_391 N_A2_M1017_g N_A_575_65#_c_813_n 5.14142e-19 $X=5.175 $Y=0.745 $X2=0
+ $Y2=0
cc_392 N_A2_M1017_g N_A_575_65#_c_814_n 0.0129371f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_393 N_A2_c_496_n N_A_575_65#_c_814_n 0.0141075f $X=5.085 $Y=1.51 $X2=0 $Y2=0
cc_394 N_A2_M1012_g N_A_575_65#_c_815_n 6.54275e-19 $X=4.745 $Y=0.745 $X2=0
+ $Y2=0
cc_395 N_A2_c_496_n N_A_575_65#_c_815_n 0.0113904f $X=5.085 $Y=1.51 $X2=0 $Y2=0
cc_396 N_A2_c_493_n N_A_575_65#_c_815_n 0.00278301f $X=5.175 $Y=1.51 $X2=0 $Y2=0
cc_397 N_VPWR_c_550_n N_X_M1000_s 0.00360572f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_398 N_VPWR_c_550_n N_X_M1003_s 0.00360572f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_399 N_VPWR_M1002_d X 0.00404285f $X=1.52 $Y=1.835 $X2=0 $Y2=0
cc_400 N_VPWR_M1021_d N_X_c_662_n 0.00419166f $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_401 N_VPWR_c_550_n N_A_878_367#_M1010_s 0.00259604f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_402 N_VPWR_c_550_n N_A_878_367#_M1015_s 0.00253292f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_403 N_VPWR_c_558_n N_A_878_367#_c_705_n 0.041633f $X=5.775 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_550_n N_A_878_367#_c_705_n 0.0372579f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_405 N_VPWR_c_555_n N_A_575_65#_c_814_n 0.0058332f $X=5.86 $Y=1.98 $X2=0 $Y2=0
cc_406 N_X_c_653_n N_VGND_M1009_d 0.00176461f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_407 N_X_c_653_n N_VGND_c_718_n 0.0170777f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_408 N_X_c_656_n N_VGND_c_725_n 0.0150063f $X=1.19 $Y=0.42 $X2=0 $Y2=0
cc_409 N_X_c_698_p N_VGND_c_726_n 0.0124525f $X=2.05 $Y=0.42 $X2=0 $Y2=0
cc_410 N_X_M1007_s N_VGND_c_729_n 0.00380103f $X=1.05 $Y=0.245 $X2=0 $Y2=0
cc_411 N_X_M1016_s N_VGND_c_729_n 0.00536646f $X=1.91 $Y=0.245 $X2=0 $Y2=0
cc_412 N_X_c_656_n N_VGND_c_729_n 0.00950443f $X=1.19 $Y=0.42 $X2=0 $Y2=0
cc_413 N_X_c_698_p N_VGND_c_729_n 0.00730901f $X=2.05 $Y=0.42 $X2=0 $Y2=0
cc_414 N_VGND_c_719_n N_A_575_65#_c_810_n 0.0362346f $X=2.48 $Y=0.39 $X2=0 $Y2=0
cc_415 N_VGND_c_720_n N_A_575_65#_c_811_n 0.00963725f $X=4.52 $Y=0.45 $X2=0
+ $Y2=0
cc_416 N_VGND_c_727_n N_A_575_65#_c_811_n 0.0623542f $X=4.355 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_729_n N_A_575_65#_c_811_n 0.0366591f $X=6 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_719_n N_A_575_65#_c_812_n 0.0139001f $X=2.48 $Y=0.39 $X2=0 $Y2=0
cc_419 N_VGND_c_727_n N_A_575_65#_c_812_n 0.0228203f $X=4.355 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_729_n N_A_575_65#_c_812_n 0.0131341f $X=6 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_M1005_d N_A_575_65#_c_825_n 0.00520049f $X=4.31 $Y=0.325 $X2=0
+ $Y2=0
cc_422 N_VGND_c_720_n N_A_575_65#_c_825_n 0.0209591f $X=4.52 $Y=0.45 $X2=0 $Y2=0
cc_423 N_VGND_c_722_n N_A_575_65#_c_825_n 0.00201146f $X=5.225 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_727_n N_A_575_65#_c_825_n 0.00200585f $X=4.355 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_729_n N_A_575_65#_c_825_n 0.00915698f $X=6 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_720_n N_A_575_65#_c_813_n 0.0109102f $X=4.52 $Y=0.45 $X2=0 $Y2=0
cc_427 N_VGND_c_721_n N_A_575_65#_c_813_n 0.0172443f $X=5.39 $Y=0.45 $X2=0 $Y2=0
cc_428 N_VGND_c_722_n N_A_575_65#_c_813_n 0.0107483f $X=5.225 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_729_n N_A_575_65#_c_813_n 0.00716399f $X=6 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_M1017_s N_A_575_65#_c_814_n 0.00176461f $X=5.25 $Y=0.325 $X2=0
+ $Y2=0
cc_431 N_VGND_c_721_n N_A_575_65#_c_814_n 0.0170777f $X=5.39 $Y=0.45 $X2=0 $Y2=0
cc_432 N_VGND_c_721_n N_A_575_65#_c_816_n 0.0222413f $X=5.39 $Y=0.45 $X2=0 $Y2=0
cc_433 N_VGND_c_728_n N_A_575_65#_c_816_n 0.0145797f $X=6 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_729_n N_A_575_65#_c_816_n 0.0101575f $X=6 $Y=0 $X2=0 $Y2=0
