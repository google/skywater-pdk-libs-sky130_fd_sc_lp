* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
X0 a_270_367# B a_360_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND D_N a_528_27# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_79_137# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_450_367# a_528_27# a_270_53# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 X a_270_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND a_79_137# a_270_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR D_N a_528_27# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_270_53# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND A a_270_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 X a_270_53# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_270_53# a_528_27# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_360_367# a_79_137# a_450_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR A a_270_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_79_137# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 X a_270_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR a_270_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VPWR a_270_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_270_53# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VGND a_270_53# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 X a_270_53# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
