* File: sky130_fd_sc_lp__sdfxtp_2.pex.spice
* Created: Wed Sep  2 10:36:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_55_119# 1 2 9 13 16 19 21 22 25 26 30 31
+ 36 41
c86 26 0 1.70252e-19 $X=1.085 $Y=1.8
c87 25 0 5.53709e-20 $X=1.085 $Y=1.8
c88 21 0 2.14447e-20 $X=1 $Y=2.385
r89 33 36 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.195 $Y=0.805
+ $X2=0.42 $Y2=0.805
r90 31 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=2.11
+ $X2=2.015 $Y2=2.275
r91 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=2.11 $X2=2.015 $Y2=2.11
r92 28 41 5.16603 $w=2.5e-07 $l=3.22102e-07 $layer=LI1_cond $X=1.25 $Y=2.11
+ $X2=1 $Y2=1.945
r93 28 30 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.25 $Y=2.11
+ $X2=2.015 $Y2=2.11
r94 26 43 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=1.085 $Y=1.8
+ $X2=1.205 $Y2=1.8
r95 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.8 $X2=1.085 $Y2=1.8
r96 23 41 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=1.945 $X2=1
+ $Y2=1.945
r97 23 25 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=1.125 $Y=1.945
+ $X2=1.125 $Y2=1.8
r98 21 41 5.16603 $w=2.5e-07 $l=4.4e-07 $layer=LI1_cond $X=1 $Y=2.385 $X2=1
+ $Y2=1.945
r99 21 22 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1 $Y=2.385 $X2=0.61
+ $Y2=2.385
r100 17 22 9.65561 $w=1.68e-07 $l=1.48e-07 $layer=LI1_cond $X=0.462 $Y=2.385
+ $X2=0.61 $Y2=2.385
r101 17 38 17.4193 $w=1.68e-07 $l=2.67e-07 $layer=LI1_cond $X=0.462 $Y=2.385
+ $X2=0.195 $Y2=2.385
r102 17 19 3.51593 $w=2.93e-07 $l=9e-08 $layer=LI1_cond $X=0.462 $Y=2.47
+ $X2=0.462 $Y2=2.56
r103 16 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.195 $Y=2.3
+ $X2=0.195 $Y2=2.385
r104 15 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.195 $Y=0.97
+ $X2=0.195 $Y2=0.805
r105 15 16 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=0.195 $Y=0.97
+ $X2=0.195 $Y2=2.3
r106 13 46 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.995 $Y=2.755
+ $X2=1.995 $Y2=2.275
r107 7 43 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.635
+ $X2=1.205 $Y2=1.8
r108 7 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.205 $Y=1.635
+ $X2=1.205 $Y2=0.805
r109 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.335
+ $Y=2.435 $X2=0.48 $Y2=2.56
r110 1 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.595 $X2=0.42 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%D 3 6 8 9 10 21 23
c42 23 0 3.37333e-20 $X=1.655 $Y=1.125
c43 8 0 1.09982e-19 $X=1.68 $Y=0.555
r44 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.655 $Y=1.29
+ $X2=1.655 $Y2=1.455
r45 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.655 $Y=1.29
+ $X2=1.655 $Y2=1.125
r46 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.29 $X2=1.655 $Y2=1.29
r47 10 22 0.092006 $w=6.48e-07 $l=5e-09 $layer=LI1_cond $X=1.44 $Y=1.295
+ $X2=1.44 $Y2=1.29
r48 9 22 6.71644 $w=6.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.44 $Y=0.925
+ $X2=1.44 $Y2=1.29
r49 8 9 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.44 $Y=0.555 $X2=1.44
+ $Y2=0.925
r50 6 24 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=1.565 $Y=2.755
+ $X2=1.565 $Y2=1.455
r51 3 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.565 $Y=0.805
+ $X2=1.565 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%SCE 2 6 7 9 10 11 12 14 16 19 23 24 25 26
+ 27 28 33
c72 24 0 2.14447e-20 $X=0.545 $Y=1.88
c73 2 0 5.53709e-20 $X=0.605 $Y=2.175
r74 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.545
+ $Y=1.375 $X2=0.545 $Y2=1.375
r75 27 28 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=2.035
r76 27 34 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.375
r77 26 34 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=0.64 $Y=1.295 $X2=0.64
+ $Y2=1.375
r78 23 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.545 $Y=1.715
+ $X2=0.545 $Y2=1.375
r79 23 24 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.715
+ $X2=0.545 $Y2=1.88
r80 22 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.21
+ $X2=0.545 $Y2=1.375
r81 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.245 $Y=0.255
+ $X2=2.245 $Y2=0.805
r82 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.205 $Y=2.325
+ $X2=1.205 $Y2=2.755
r83 13 25 5.30422 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=0.77 $Y=2.25
+ $X2=0.65 $Y2=2.25
r84 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.13 $Y=2.25
+ $X2=1.205 $Y2=2.325
r85 12 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.13 $Y=2.25
+ $X2=0.77 $Y2=2.25
r86 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.17 $Y=0.18
+ $X2=2.245 $Y2=0.255
r87 10 11 748.638 $w=1.5e-07 $l=1.46e-06 $layer=POLY_cond $X=2.17 $Y=0.18
+ $X2=0.71 $Y2=0.18
r88 7 25 20.4101 $w=1.5e-07 $l=9.48683e-08 $layer=POLY_cond $X=0.695 $Y=2.325
+ $X2=0.65 $Y2=2.25
r89 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.695 $Y=2.325
+ $X2=0.695 $Y2=2.755
r90 6 22 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.635 $Y=0.805
+ $X2=0.635 $Y2=1.21
r91 3 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.635 $Y=0.255
+ $X2=0.71 $Y2=0.18
r92 3 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.635 $Y=0.255
+ $X2=0.635 $Y2=0.805
r93 2 25 20.4101 $w=1.5e-07 $l=9.48683e-08 $layer=POLY_cond $X=0.605 $Y=2.175
+ $X2=0.65 $Y2=2.25
r94 2 24 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.605 $Y=2.175
+ $X2=0.605 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%SCD 3 7 9 10 14
r48 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.54
+ $X2=2.515 $Y2=1.705
r49 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.54
+ $X2=2.515 $Y2=1.375
r50 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.54 $X2=2.515 $Y2=1.54
r51 10 15 4.50173 $w=3.18e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=2.515 $Y2=1.615
r52 9 15 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=2.515 $Y2=1.615
r53 7 16 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.605 $Y=0.805
+ $X2=2.605 $Y2=1.375
r54 3 17 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.465 $Y=2.755
+ $X2=2.465 $Y2=1.705
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%CLK 3 7 11 12 13 14 15 20
c50 13 0 1.59499e-19 $X=3.6 $Y=1.295
c51 12 0 8.53846e-20 $X=3.202 $Y=2.095
c52 11 0 9.65774e-20 $X=3.202 $Y=1.945
r53 20 22 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.277 $Y=1.59
+ $X2=3.277 $Y2=1.425
r54 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.34
+ $Y=1.59 $X2=3.34 $Y2=1.59
r55 14 15 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.495 $Y=1.665
+ $X2=3.495 $Y2=2.035
r56 14 21 1.86887 $w=4.78e-07 $l=7.5e-08 $layer=LI1_cond $X=3.495 $Y=1.665
+ $X2=3.495 $Y2=1.59
r57 13 21 7.3509 $w=4.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.495 $Y=1.295
+ $X2=3.495 $Y2=1.59
r58 11 12 45.2433 $w=4.55e-07 $l=1.5e-07 $layer=POLY_cond $X=3.202 $Y=1.945
+ $X2=3.202 $Y2=2.095
r59 9 20 7.57836 $w=4.55e-07 $l=6.2e-08 $layer=POLY_cond $X=3.277 $Y=1.652
+ $X2=3.277 $Y2=1.59
r60 9 11 35.8139 $w=4.55e-07 $l=2.93e-07 $layer=POLY_cond $X=3.277 $Y=1.652
+ $X2=3.277 $Y2=1.945
r61 7 22 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.125 $Y=0.805
+ $X2=3.125 $Y2=1.425
r62 3 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.975 $Y=2.755
+ $X2=2.975 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_610_487# 1 2 9 11 13 16 20 24 28 31 34 36
+ 40 41 45 46 48 49 50 52 54 55 58 59 60 62 64 65 66 69 70 73 78 80 85 86 92 98
c236 92 0 1.98119e-19 $X=5.605 $Y=1.59
c237 85 0 2.24563e-19 $X=7.465 $Y=1.93
c238 78 0 1.65685e-19 $X=5.76 $Y=1.59
c239 59 0 1.16002e-19 $X=7.295 $Y=2.83
c240 52 0 8.45676e-20 $X=5.76 $Y=2.115
c241 31 0 1.59499e-19 $X=3.99 $Y=2.085
c242 20 0 3.65866e-19 $X=5.605 $Y=2.465
r243 85 96 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.465 $Y=1.93
+ $X2=7.465 $Y2=2.095
r244 84 86 4.25903 $w=2.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.465 $Y=1.95
+ $X2=7.55 $Y2=1.95
r245 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.465
+ $Y=1.93 $X2=7.465 $Y2=1.93
r246 81 84 4.25903 $w=2.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=1.95
+ $X2=7.465 $Y2=1.95
r247 76 92 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.58 $Y=1.59
+ $X2=5.605 $Y2=1.59
r248 76 89 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.58 $Y=1.59
+ $X2=5.16 $Y2=1.59
r249 75 78 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.58 $Y=1.59
+ $X2=5.76 $Y2=1.59
r250 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.58
+ $Y=1.59 $X2=5.58 $Y2=1.59
r251 70 98 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.185 $Y=1.01
+ $X2=8.185 $Y2=0.845
r252 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.185
+ $Y=1.01 $X2=8.185 $Y2=1.01
r253 67 69 10.1799 $w=2.98e-07 $l=2.65e-07 $layer=LI1_cond $X=8.17 $Y=1.275
+ $X2=8.17 $Y2=1.01
r254 65 67 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=8.02 $Y=1.36
+ $X2=8.17 $Y2=1.275
r255 65 66 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.02 $Y=1.36
+ $X2=7.635 $Y2=1.36
r256 64 86 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.55 $Y=1.835
+ $X2=7.55 $Y2=1.95
r257 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.55 $Y=1.445
+ $X2=7.635 $Y2=1.36
r258 63 64 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.55 $Y=1.445
+ $X2=7.55 $Y2=1.835
r259 61 81 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.38 $Y=2.065
+ $X2=7.38 $Y2=1.95
r260 61 62 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.38 $Y=2.065
+ $X2=7.38 $Y2=2.745
r261 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.295 $Y=2.83
+ $X2=7.38 $Y2=2.745
r262 59 60 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.295 $Y=2.83
+ $X2=6.715 $Y2=2.83
r263 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.63 $Y=2.745
+ $X2=6.715 $Y2=2.83
r264 57 58 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.63 $Y=2.285
+ $X2=6.63 $Y2=2.745
r265 56 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.2
+ $X2=5.76 $Y2=2.2
r266 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.545 $Y=2.2
+ $X2=6.63 $Y2=2.285
r267 55 56 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.545 $Y=2.2
+ $X2=5.845 $Y2=2.2
r268 53 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.285
+ $X2=5.76 $Y2=2.2
r269 53 54 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.76 $Y=2.285
+ $X2=5.76 $Y2=2.835
r270 52 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.115
+ $X2=5.76 $Y2=2.2
r271 51 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=1.755
+ $X2=5.76 $Y2=1.59
r272 51 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.76 $Y=1.755
+ $X2=5.76 $Y2=2.115
r273 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.675 $Y=2.92
+ $X2=5.76 $Y2=2.835
r274 49 50 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=5.675 $Y=2.92
+ $X2=4.145 $Y2=2.92
r275 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=2.835
+ $X2=4.145 $Y2=2.92
r276 47 73 4.40882 $w=2.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.06 $Y=2.47
+ $X2=4.025 $Y2=2.385
r277 47 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.06 $Y=2.47
+ $X2=4.06 $Y2=2.835
r278 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.99
+ $Y=1.59 $X2=3.99 $Y2=1.59
r279 43 73 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=2.3
+ $X2=4.025 $Y2=2.385
r280 43 45 34.0931 $w=2.38e-07 $l=7.1e-07 $layer=LI1_cond $X=4.025 $Y=2.3
+ $X2=4.025 $Y2=1.59
r281 42 72 0.587687 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=1.03
+ $X2=4.025 $Y2=0.865
r282 42 45 26.8903 $w=2.38e-07 $l=5.6e-07 $layer=LI1_cond $X=4.025 $Y=1.03
+ $X2=4.025 $Y2=1.59
r283 40 73 2.0246 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.905 $Y=2.385
+ $X2=4.025 $Y2=2.385
r284 40 41 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.905 $Y=2.385
+ $X2=3.355 $Y2=2.385
r285 36 72 11.5649 $w=3.3e-07 $l=2.85e-07 $layer=LI1_cond $X=3.74 $Y=0.865
+ $X2=4.025 $Y2=0.865
r286 36 38 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.74 $Y=0.865 $X2=3.34
+ $Y2=0.865
r287 32 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.19 $Y=2.47
+ $X2=3.355 $Y2=2.385
r288 32 34 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.19 $Y=2.47
+ $X2=3.19 $Y2=2.58
r289 31 46 86.5563 $w=3.3e-07 $l=4.95e-07 $layer=POLY_cond $X=3.99 $Y=2.085
+ $X2=3.99 $Y2=1.59
r290 30 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=1.425
+ $X2=3.99 $Y2=1.59
r291 28 98 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.275 $Y=0.525
+ $X2=8.275 $Y2=0.845
r292 24 96 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.515 $Y=2.675
+ $X2=7.515 $Y2=2.095
r293 18 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.605 $Y=1.755
+ $X2=5.605 $Y2=1.59
r294 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.605 $Y=1.755
+ $X2=5.605 $Y2=2.465
r295 14 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.16 $Y=1.425
+ $X2=5.16 $Y2=1.59
r296 14 16 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.16 $Y=1.425
+ $X2=5.16 $Y2=0.835
r297 11 31 23.7049 $w=3.05e-07 $l=2.69768e-07 $layer=POLY_cond $X=4.195 $Y=2.235
+ $X2=3.99 $Y2=2.085
r298 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.195 $Y=2.235
+ $X2=4.195 $Y2=2.665
r299 9 30 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.08 $Y=0.445
+ $X2=4.08 $Y2=1.425
r300 2 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.05
+ $Y=2.435 $X2=3.19 $Y2=2.58
r301 1 38 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.595 $X2=3.34 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_831_47# 1 2 8 9 10 11 13 16 19 21 22 23
+ 26 29 32 34 35 39 43 45 46 47 49 50 51 54 55 57 62 67 69
c172 67 0 2.63883e-19 $X=5.61 $Y=0.515
c173 54 0 5.72802e-20 $X=7.63 $Y=1.01
c174 26 0 1.16002e-19 $X=8.04 $Y=2.675
c175 9 0 2.51969e-19 $X=5.1 $Y=2.07
r176 61 62 29.5968 $w=2.18e-07 $l=5.65e-07 $layer=LI1_cond $X=4.425 $Y=0.61
+ $X2=4.425 $Y2=1.175
r177 60 61 7.02548 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=0.445
+ $X2=4.365 $Y2=0.61
r178 57 60 2.37268 $w=3.38e-07 $l=7e-08 $layer=LI1_cond $X=4.365 $Y=0.375
+ $X2=4.365 $Y2=0.445
r179 55 69 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.01
+ $X2=7.615 $Y2=0.845
r180 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.63
+ $Y=1.01 $X2=7.63 $Y2=1.01
r181 52 54 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=7.63 $Y=0.425
+ $X2=7.63 $Y2=1.01
r182 50 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.465 $Y=0.34
+ $X2=7.63 $Y2=0.425
r183 50 51 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.465 $Y=0.34
+ $X2=6.935 $Y2=0.34
r184 48 51 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.825 $Y=0.425
+ $X2=6.935 $Y2=0.34
r185 48 49 15.7151 $w=2.18e-07 $l=3e-07 $layer=LI1_cond $X=6.825 $Y=0.425
+ $X2=6.825 $Y2=0.725
r186 46 49 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.715 $Y=0.81
+ $X2=6.825 $Y2=0.725
r187 46 47 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.715 $Y=0.81
+ $X2=5.965 $Y2=0.81
r188 45 47 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=5.812 $Y=0.725
+ $X2=5.965 $Y2=0.81
r189 44 45 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=5.812 $Y=0.485
+ $X2=5.812 $Y2=0.725
r190 43 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.35
+ $X2=5.61 $Y2=0.515
r191 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.61
+ $Y=0.35 $X2=5.61 $Y2=0.35
r192 40 57 3.28461 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=4.535 $Y=0.375
+ $X2=4.365 $Y2=0.375
r193 40 42 56.3126 $w=2.18e-07 $l=1.075e-06 $layer=LI1_cond $X=4.535 $Y=0.375
+ $X2=5.61 $Y2=0.375
r194 39 44 7.05149 $w=2.2e-07 $l=1.9956e-07 $layer=LI1_cond $X=5.66 $Y=0.375
+ $X2=5.812 $Y2=0.485
r195 39 42 2.61919 $w=2.18e-07 $l=5e-08 $layer=LI1_cond $X=5.66 $Y=0.375
+ $X2=5.61 $Y2=0.375
r196 34 37 42.7519 $w=3.08e-07 $l=1.15e-06 $layer=LI1_cond $X=4.47 $Y=1.34
+ $X2=4.47 $Y2=2.49
r197 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.53
+ $Y=1.34 $X2=4.53 $Y2=1.34
r198 32 62 6.74938 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=4.47 $Y=1.33
+ $X2=4.47 $Y2=1.175
r199 32 34 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=4.47 $Y=1.33
+ $X2=4.47 $Y2=1.34
r200 28 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.53 $Y=1.68
+ $X2=4.53 $Y2=1.34
r201 28 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.53 $Y=1.68
+ $X2=4.53 $Y2=1.845
r202 24 26 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=8.04 $Y=1.535
+ $X2=8.04 $Y2=2.675
r203 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.965 $Y=1.46
+ $X2=8.04 $Y2=1.535
r204 22 23 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.965 $Y=1.46
+ $X2=7.795 $Y2=1.46
r205 21 23 33.3473 $w=1.5e-07 $l=2.14243e-07 $layer=POLY_cond $X=7.615 $Y=1.385
+ $X2=7.795 $Y2=1.46
r206 20 55 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=7.615 $Y=1.025
+ $X2=7.615 $Y2=1.01
r207 20 21 57.7042 $w=3.6e-07 $l=3.6e-07 $layer=POLY_cond $X=7.615 $Y=1.025
+ $X2=7.615 $Y2=1.385
r208 19 69 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.51 $Y=0.525
+ $X2=7.51 $Y2=0.845
r209 16 67 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.67 $Y=0.835
+ $X2=5.67 $Y2=0.515
r210 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.175 $Y=2.145
+ $X2=5.175 $Y2=2.465
r211 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.1 $Y=2.07
+ $X2=5.175 $Y2=2.145
r212 9 10 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=5.1 $Y=2.07
+ $X2=4.695 $Y2=2.07
r213 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.62 $Y=1.995
+ $X2=4.695 $Y2=2.07
r214 8 29 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.62 $Y=1.995
+ $X2=4.62 $Y2=1.845
r215 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=2.345 $X2=4.41 $Y2=2.49
r216 1 60 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.235 $X2=4.295 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_1178_399# 1 2 9 12 16 17 18 20 22 26 30
+ 32
c77 32 0 1.74622e-19 $X=6.355 $Y=1.685
c78 30 0 5.62581e-20 $X=6.19 $Y=1.51
r79 30 35 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.51
+ $X2=6.17 $Y2=1.345
r80 29 32 4.04459 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=1.685
+ $X2=6.355 $Y2=1.685
r81 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.19
+ $Y=1.51 $X2=6.19 $Y2=1.51
r82 24 26 42.9043 $w=1.88e-07 $l=7.35e-07 $layer=LI1_cond $X=7.2 $Y=1.495
+ $X2=7.2 $Y2=0.76
r83 20 22 22.3286 $w=2.38e-07 $l=4.65e-07 $layer=LI1_cond $X=7.005 $Y=1.945
+ $X2=7.005 $Y2=2.41
r84 18 20 9.60442 $w=3.04e-07 $l=2.64102e-07 $layer=LI1_cond $X=7.09 $Y=1.72
+ $X2=7.005 $Y2=1.945
r85 18 24 10.7359 $w=3.04e-07 $l=2.74545e-07 $layer=LI1_cond $X=7.09 $Y=1.72
+ $X2=7.2 $Y2=1.495
r86 18 32 14.0871 $w=4.48e-07 $l=5.3e-07 $layer=LI1_cond $X=6.885 $Y=1.72
+ $X2=6.355 $Y2=1.72
r87 16 17 44.4176 $w=3.7e-07 $l=1.5e-07 $layer=POLY_cond $X=6.122 $Y=1.995
+ $X2=6.122 $Y2=2.145
r88 14 30 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=6.17 $Y=1.53 $X2=6.17
+ $Y2=1.51
r89 14 16 72.5202 $w=3.7e-07 $l=4.65e-07 $layer=POLY_cond $X=6.17 $Y=1.53
+ $X2=6.17 $Y2=1.995
r90 12 35 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.06 $Y=0.835
+ $X2=6.06 $Y2=1.345
r91 9 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.965 $Y=2.465
+ $X2=5.965 $Y2=2.145
r92 2 22 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=2.255 $X2=7.03 $Y2=2.41
r93 1 26 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=7.06
+ $Y=0.315 $X2=7.2 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_1047_125# 1 2 9 11 13 15 18 22 26 29 32
+ 34 39
c95 15 0 2.23659e-19 $X=5.23 $Y=1.935
r96 38 39 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=6.815 $Y=1.23
+ $X2=6.985 $Y2=1.23
r97 33 38 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.77 $Y=1.23
+ $X2=6.815 $Y2=1.23
r98 32 34 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.77 $Y=1.2
+ $X2=6.605 $Y2=1.2
r99 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.23 $X2=6.77 $Y2=1.23
r100 27 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.23 $Y=2.02
+ $X2=5.4 $Y2=2.02
r101 25 26 1.84097 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.49 $Y=1.16
+ $X2=5.317 $Y2=1.16
r102 25 34 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.49 $Y=1.16
+ $X2=6.605 $Y2=1.16
r103 20 29 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=2.105
+ $X2=5.4 $Y2=2.02
r104 20 22 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=5.4 $Y=2.105
+ $X2=5.4 $Y2=2.465
r105 16 26 4.60183 $w=1.95e-07 $l=1.12161e-07 $layer=LI1_cond $X=5.38 $Y=1.075
+ $X2=5.317 $Y2=1.16
r106 16 18 12.5721 $w=2.18e-07 $l=2.4e-07 $layer=LI1_cond $X=5.38 $Y=1.075
+ $X2=5.38 $Y2=0.835
r107 15 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.23 $Y=1.935
+ $X2=5.23 $Y2=2.02
r108 14 26 4.60183 $w=1.95e-07 $l=1.22327e-07 $layer=LI1_cond $X=5.23 $Y=1.245
+ $X2=5.317 $Y2=1.16
r109 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.23 $Y=1.245
+ $X2=5.23 $Y2=1.935
r110 11 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.985 $Y=1.065
+ $X2=6.985 $Y2=1.23
r111 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.985 $Y=1.065
+ $X2=6.985 $Y2=0.635
r112 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.395
+ $X2=6.815 $Y2=1.23
r113 7 9 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=6.815 $Y=1.395
+ $X2=6.815 $Y2=2.675
r114 2 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=2.255 $X2=5.39 $Y2=2.465
r115 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.235
+ $Y=0.625 $X2=5.375 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_1665_381# 1 2 9 13 15 17 20 22 24 27 29
+ 36 40 43 45 48 51 52 53 57 62
r103 61 62 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=10.125 $Y=1.51
+ $X2=10.555 $Y2=1.51
r104 49 61 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=9.97 $Y=1.51
+ $X2=10.125 $Y2=1.51
r105 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.97
+ $Y=1.51 $X2=9.97 $Y2=1.51
r106 46 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.55 $Y=1.51
+ $X2=9.465 $Y2=1.51
r107 46 48 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.55 $Y=1.51
+ $X2=9.97 $Y2=1.51
r108 45 52 4.48993 $w=2.12e-07 $l=1.09407e-07 $layer=LI1_cond $X=9.465 $Y=1.975
+ $X2=9.422 $Y2=2.065
r109 44 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.465 $Y=1.675
+ $X2=9.465 $Y2=1.51
r110 44 45 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.465 $Y=1.675
+ $X2=9.465 $Y2=1.975
r111 43 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.465 $Y=1.345
+ $X2=9.465 $Y2=1.51
r112 43 51 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.465 $Y=1.345
+ $X2=9.465 $Y2=0.895
r113 38 52 4.48993 $w=2.12e-07 $l=9e-08 $layer=LI1_cond $X=9.422 $Y=2.155
+ $X2=9.422 $Y2=2.065
r114 38 40 1.58178 $w=2.53e-07 $l=3.5e-08 $layer=LI1_cond $X=9.422 $Y=2.155
+ $X2=9.422 $Y2=2.19
r115 34 51 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=9.38 $Y=0.725
+ $X2=9.38 $Y2=0.895
r116 34 36 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=9.38 $Y=0.725
+ $X2=9.38 $Y2=0.39
r117 32 57 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=8.49 $Y=2.07
+ $X2=8.635 $Y2=2.07
r118 32 54 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.49 $Y=2.07 $X2=8.4
+ $Y2=2.07
r119 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.49
+ $Y=2.07 $X2=8.49 $Y2=2.07
r120 29 52 1.94654 $w=1.8e-07 $l=1.27e-07 $layer=LI1_cond $X=9.295 $Y=2.065
+ $X2=9.422 $Y2=2.065
r121 29 31 49.601 $w=1.78e-07 $l=8.05e-07 $layer=LI1_cond $X=9.295 $Y=2.065
+ $X2=8.49 $Y2=2.065
r122 25 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.555 $Y=1.675
+ $X2=10.555 $Y2=1.51
r123 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.555 $Y=1.675
+ $X2=10.555 $Y2=2.465
r124 22 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.555 $Y=1.345
+ $X2=10.555 $Y2=1.51
r125 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.555 $Y=1.345
+ $X2=10.555 $Y2=0.815
r126 18 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.125 $Y=1.675
+ $X2=10.125 $Y2=1.51
r127 18 20 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.125 $Y=1.675
+ $X2=10.125 $Y2=2.465
r128 15 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.125 $Y=1.345
+ $X2=10.125 $Y2=1.51
r129 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.125 $Y=1.345
+ $X2=10.125 $Y2=0.815
r130 11 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.635 $Y=1.905
+ $X2=8.635 $Y2=2.07
r131 11 13 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=8.635 $Y=1.905
+ $X2=8.635 $Y2=0.525
r132 7 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.4 $Y=2.235
+ $X2=8.4 $Y2=2.07
r133 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.4 $Y=2.235 $X2=8.4
+ $Y2=2.675
r134 2 40 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.25
+ $Y=2.045 $X2=9.39 $Y2=2.19
r135 1 36 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=9.235
+ $Y=0.235 $X2=9.375 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_1517_63# 1 2 9 13 17 18 23 28 30 32 33 35
+ 37 38
c98 28 0 1.67283e-19 $X=7.985 $Y=1.72
r99 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.115
+ $Y=1.3 $X2=9.115 $Y2=1.3
r100 34 37 9.64003 $w=6.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.575 $Y=1.47
+ $X2=9.115 $Y2=1.47
r101 34 35 9.18355 $w=6.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=1.47
+ $X2=8.49 $Y2=1.47
r102 32 33 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.81 $Y=2.4
+ $X2=7.81 $Y2=2.235
r103 30 34 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.575 $Y=1.135
+ $X2=8.575 $Y2=1.47
r104 29 30 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=8.575 $Y=0.665
+ $X2=8.575 $Y2=1.135
r105 28 35 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=7.985 $Y=1.72
+ $X2=8.49 $Y2=1.72
r106 23 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.49 $Y=0.5
+ $X2=8.575 $Y2=0.665
r107 23 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.49 $Y=0.5
+ $X2=8.06 $Y2=0.5
r108 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.9 $Y=1.805
+ $X2=7.985 $Y2=1.72
r109 21 33 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.9 $Y=1.805
+ $X2=7.9 $Y2=2.235
r110 17 38 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.115 $Y=1.64
+ $X2=9.115 $Y2=1.3
r111 17 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=1.64
+ $X2=9.115 $Y2=1.805
r112 16 38 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=1.135
+ $X2=9.115 $Y2=1.3
r113 13 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.175 $Y=2.465
+ $X2=9.175 $Y2=1.805
r114 9 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.16 $Y=0.555
+ $X2=9.16 $Y2=1.135
r115 2 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.59
+ $Y=2.255 $X2=7.73 $Y2=2.4
r116 1 25 182 $w=1.7e-07 $l=5.59911e-07 $layer=licon1_NDIFF $count=1 $X=7.585
+ $Y=0.315 $X2=8.06 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%VPWR 1 2 3 4 5 6 7 24 28 30 34 38 42 48 52
+ 54 59 60 62 63 64 70 81 88 93 99 102 105 108 112
c140 62 0 1.91244e-19 $X=6.095 $Y=3.33
c141 24 0 6.027e-20 $X=0.945 $Y=2.77
c142 2 0 7.12511e-20 $X=2.54 $Y=2.435
r143 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r144 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r146 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r148 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r149 97 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r150 97 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r151 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r152 94 108 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=10.055 $Y=3.33
+ $X2=9.9 $Y2=3.33
r153 94 96 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.055 $Y=3.33
+ $X2=10.32 $Y2=3.33
r154 93 111 4.47956 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.837 $Y2=3.33
r155 93 96 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.32 $Y2=3.33
r156 92 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r157 92 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r159 89 105 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=8.787 $Y2=3.33
r160 89 91 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 88 108 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.745 $Y=3.33
+ $X2=9.9 $Y2=3.33
r162 88 91 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.745 $Y=3.33
+ $X2=9.36 $Y2=3.33
r163 87 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r164 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r165 84 87 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r166 83 86 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r167 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 81 105 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=8.45 $Y=3.33
+ $X2=8.787 $Y2=3.33
r169 81 86 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=8.45 $Y=3.33 $X2=8.4
+ $Y2=3.33
r170 80 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r171 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r172 77 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r173 76 79 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r174 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 74 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.805 $Y=3.33
+ $X2=3.68 $Y2=3.33
r176 74 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.805 $Y=3.33
+ $X2=4.08 $Y2=3.33
r177 73 100 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r178 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r179 70 99 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.735 $Y2=3.33
r180 70 72 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=1.2 $Y2=3.33
r181 68 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r182 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r183 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r184 64 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.08 $Y2=3.33
r185 62 79 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.095 $Y=3.33 $X2=6
+ $Y2=3.33
r186 62 63 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6.235 $Y2=3.33
r187 61 83 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.375 $Y=3.33
+ $X2=6.48 $Y2=3.33
r188 61 63 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.375 $Y=3.33
+ $X2=6.235 $Y2=3.33
r189 59 67 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.78 $Y=3.33 $X2=0.72
+ $Y2=3.33
r190 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=3.33
+ $X2=0.945 $Y2=3.33
r191 58 72 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.11 $Y=3.33 $X2=1.2
+ $Y2=3.33
r192 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=3.33
+ $X2=0.945 $Y2=3.33
r193 54 57 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=10.785 $Y=1.98
+ $X2=10.785 $Y2=2.95
r194 52 111 3.03811 $w=3e-07 $l=1.07912e-07 $layer=LI1_cond $X=10.785 $Y=3.245
+ $X2=10.837 $Y2=3.33
r195 52 57 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=10.785 $Y=3.245
+ $X2=10.785 $Y2=2.95
r196 48 51 34.945 $w=3.08e-07 $l=9.4e-07 $layer=LI1_cond $X=9.9 $Y=2.01 $X2=9.9
+ $Y2=2.95
r197 46 108 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.9 $Y=3.245
+ $X2=9.9 $Y2=3.33
r198 46 51 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=9.9 $Y=3.245
+ $X2=9.9 $Y2=2.95
r199 42 45 6.20189 $w=6.73e-07 $l=3.5e-07 $layer=LI1_cond $X=8.787 $Y=2.41
+ $X2=8.787 $Y2=2.76
r200 40 105 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=8.787 $Y=3.245
+ $X2=8.787 $Y2=3.33
r201 40 45 8.59404 $w=6.73e-07 $l=4.85e-07 $layer=LI1_cond $X=8.787 $Y=3.245
+ $X2=8.787 $Y2=2.76
r202 36 63 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=3.245
+ $X2=6.235 $Y2=3.33
r203 36 38 25.7242 $w=2.78e-07 $l=6.25e-07 $layer=LI1_cond $X=6.235 $Y=3.245
+ $X2=6.235 $Y2=2.62
r204 32 102 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=3.245
+ $X2=3.68 $Y2=3.33
r205 32 34 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=3.68 $Y=3.245
+ $X2=3.68 $Y2=2.805
r206 31 99 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.735 $Y2=3.33
r207 30 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.555 $Y=3.33
+ $X2=3.68 $Y2=3.33
r208 30 31 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.555 $Y=3.33
+ $X2=2.845 $Y2=3.33
r209 26 99 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=3.245
+ $X2=2.735 $Y2=3.33
r210 26 28 20.4297 $w=2.18e-07 $l=3.9e-07 $layer=LI1_cond $X=2.735 $Y=3.245
+ $X2=2.735 $Y2=2.855
r211 22 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=3.245
+ $X2=0.945 $Y2=3.33
r212 22 24 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.945 $Y=3.245
+ $X2=0.945 $Y2=2.77
r213 7 57 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.835 $X2=10.77 $Y2=2.95
r214 7 54 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.835 $X2=10.77 $Y2=1.98
r215 6 51 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=9.785
+ $Y=1.835 $X2=9.91 $Y2=2.95
r216 6 48 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=9.785
+ $Y=1.835 $X2=9.91 $Y2=2.01
r217 5 45 400 $w=1.7e-07 $l=6.15061e-07 $layer=licon1_PDIFF $count=1 $X=8.475
+ $Y=2.465 $X2=8.96 $Y2=2.76
r218 5 42 400 $w=1.7e-07 $l=5.11762e-07 $layer=licon1_PDIFF $count=1 $X=8.475
+ $Y=2.465 $X2=8.96 $Y2=2.41
r219 4 38 300 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_PDIFF $count=2 $X=6.04
+ $Y=2.255 $X2=6.26 $Y2=2.62
r220 3 34 600 $w=1.7e-07 $l=5.23163e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=2.345 $X2=3.72 $Y2=2.805
r221 2 28 600 $w=1.7e-07 $l=5.10294e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=2.435 $X2=2.74 $Y2=2.855
r222 1 24 600 $w=1.7e-07 $l=4.1334e-07 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=2.435 $X2=0.945 $Y2=2.77
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%A_328_119# 1 2 3 4 17 19 21 22 23 24 26 27
+ 28 30 35 36 39 42 49
c129 49 0 1.51886e-19 $X=4.96 $Y=2.4
c130 42 0 4.62334e-20 $X=5.04 $Y=2.405
c131 39 0 1.92177e-19 $X=2.64 $Y=2.405
c132 27 0 9.81978e-20 $X=4.88 $Y=0.955
c133 22 0 3.37333e-20 $X=2.135 $Y=1.2
c134 21 0 8.53846e-20 $X=2.905 $Y=1.2
r135 42 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.405
+ $X2=5.04 $Y2=2.405
r136 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=2.405
+ $X2=2.64 $Y2=2.405
r137 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=2.405
+ $X2=2.64 $Y2=2.405
r138 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.405
+ $X2=5.04 $Y2=2.405
r139 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.895 $Y=2.405
+ $X2=2.785 $Y2=2.405
r140 32 39 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=2.505 $Y=2.445
+ $X2=2.505 $Y2=2.405
r141 31 39 7.46469 $w=4.38e-07 $l=2.85e-07 $layer=LI1_cond $X=2.505 $Y=2.12
+ $X2=2.505 $Y2=2.405
r142 28 49 2.92684 $w=3.13e-07 $l=8e-08 $layer=LI1_cond $X=4.88 $Y=2.432
+ $X2=4.96 $Y2=2.432
r143 27 34 8.96496 $w=3.09e-07 $l=1.86145e-07 $layer=LI1_cond $X=4.88 $Y=0.955
+ $X2=4.925 $Y2=0.79
r144 27 28 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=4.88 $Y=0.955
+ $X2=4.88 $Y2=2.275
r145 25 26 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.99 $Y=1.285
+ $X2=2.99 $Y2=1.95
r146 24 31 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=2.725 $Y=2.035
+ $X2=2.505 $Y2=2.12
r147 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=2.035
+ $X2=2.99 $Y2=1.95
r148 23 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.905 $Y=2.035
+ $X2=2.725 $Y2=2.035
r149 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=1.2
+ $X2=2.99 $Y2=1.285
r150 21 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.905 $Y=1.2
+ $X2=2.135 $Y2=1.2
r151 20 30 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=2.545
+ $X2=1.78 $Y2=2.545
r152 19 32 29.065 $w=8.9e-08 $l=2.6533e-07 $layer=LI1_cond $X=2.285 $Y=2.545
+ $X2=2.505 $Y2=2.445
r153 19 20 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.285 $Y=2.545
+ $X2=1.945 $Y2=2.545
r154 15 22 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.035 $Y=1.115
+ $X2=2.135 $Y2=1.2
r155 15 17 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=2.035 $Y=1.115
+ $X2=2.035 $Y2=0.805
r156 4 49 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.835
+ $Y=2.255 $X2=4.96 $Y2=2.4
r157 3 30 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.64
+ $Y=2.435 $X2=1.78 $Y2=2.58
r158 2 34 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.8
+ $Y=0.625 $X2=4.925 $Y2=0.79
r159 1 17 182 $w=1.7e-07 $l=4.73498e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.595 $X2=2.02 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%Q 1 2 7 8 9 10 11 12 13
r18 13 39 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=10.345 $Y=2.775
+ $X2=10.345 $Y2=2.91
r19 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=2.405
+ $X2=10.345 $Y2=2.775
r20 11 12 20.4078 $w=2.38e-07 $l=4.25e-07 $layer=LI1_cond $X=10.345 $Y=1.98
+ $X2=10.345 $Y2=2.405
r21 10 11 15.1258 $w=2.38e-07 $l=3.15e-07 $layer=LI1_cond $X=10.345 $Y=1.665
+ $X2=10.345 $Y2=1.98
r22 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=1.295
+ $X2=10.345 $Y2=1.665
r23 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.345 $Y=0.925
+ $X2=10.345 $Y2=1.295
r24 7 8 18.4871 $w=2.38e-07 $l=3.85e-07 $layer=LI1_cond $X=10.345 $Y=0.54
+ $X2=10.345 $Y2=0.925
r25 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.2
+ $Y=1.835 $X2=10.34 $Y2=2.91
r26 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.2
+ $Y=1.835 $X2=10.34 $Y2=1.98
r27 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.2
+ $Y=0.395 $X2=10.34 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 38 42 46 48
+ 50 53 54 56 57 59 60 61 76 83 88 94 97 100 104
r118 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r119 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r120 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r121 95 98 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.88
+ $Y2=0
r122 94 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r123 92 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r124 92 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r125 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r126 89 100 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=10.055 $Y=0
+ $X2=9.9 $Y2=0
r127 89 91 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.055 $Y=0
+ $X2=10.32 $Y2=0
r128 88 103 4.47956 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.837 $Y2=0
r129 88 91 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.32 $Y2=0
r130 87 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r131 87 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r132 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r133 84 97 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=9.04 $Y=0 $X2=8.935
+ $Y2=0
r134 84 86 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.04 $Y=0 $X2=9.36
+ $Y2=0
r135 83 100 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.745 $Y=0 $X2=9.9
+ $Y2=0
r136 83 86 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.745 $Y=0
+ $X2=9.36 $Y2=0
r137 82 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r138 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r139 78 81 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r140 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r141 76 94 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.375
+ $Y2=0
r142 76 81 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6
+ $Y2=0
r143 75 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r144 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r145 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r146 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r147 69 72 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r148 68 71 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r149 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r150 65 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r151 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r152 61 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r153 61 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=4.08 $Y2=0
r154 59 74 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.6
+ $Y2=0
r155 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.86
+ $Y2=0
r156 58 78 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.025 $Y=0 $X2=4.08
+ $Y2=0
r157 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=3.86
+ $Y2=0
r158 56 71 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.64
+ $Y2=0
r159 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.86
+ $Y2=0
r160 55 74 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=3.6
+ $Y2=0
r161 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.86
+ $Y2=0
r162 53 64 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.72
+ $Y2=0
r163 53 54 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.835
+ $Y2=0
r164 52 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r165 52 54 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.835
+ $Y2=0
r166 48 103 3.03811 $w=3e-07 $l=1.07912e-07 $layer=LI1_cond $X=10.785 $Y=0.085
+ $X2=10.837 $Y2=0
r167 48 50 17.4787 $w=2.98e-07 $l=4.55e-07 $layer=LI1_cond $X=10.785 $Y=0.085
+ $X2=10.785 $Y2=0.54
r168 44 100 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.9 $Y=0.085
+ $X2=9.9 $Y2=0
r169 44 46 16.9149 $w=3.08e-07 $l=4.55e-07 $layer=LI1_cond $X=9.9 $Y=0.085
+ $X2=9.9 $Y2=0.54
r170 40 97 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=0.085
+ $X2=8.935 $Y2=0
r171 40 42 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=8.935 $Y=0.085
+ $X2=8.935 $Y2=0.38
r172 39 94 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.545 $Y=0 $X2=6.375
+ $Y2=0
r173 38 97 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.83 $Y=0 $X2=8.935
+ $Y2=0
r174 38 39 149.075 $w=1.68e-07 $l=2.285e-06 $layer=LI1_cond $X=8.83 $Y=0
+ $X2=6.545 $Y2=0
r175 34 94 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0
r176 34 36 12.7108 $w=3.38e-07 $l=3.75e-07 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0.46
r177 30 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0
r178 30 32 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0.41
r179 26 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r180 26 28 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.805
r181 22 54 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.085
+ $X2=0.835 $Y2=0
r182 22 24 37.7163 $w=2.18e-07 $l=7.2e-07 $layer=LI1_cond $X=0.835 $Y=0.085
+ $X2=0.835 $Y2=0.805
r183 7 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.63
+ $Y=0.395 $X2=10.77 $Y2=0.54
r184 6 46 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=9.785
+ $Y=0.395 $X2=9.91 $Y2=0.54
r185 5 42 91 $w=1.7e-07 $l=2.65518e-07 $layer=licon1_NDIFF $count=2 $X=8.71
+ $Y=0.315 $X2=8.945 $Y2=0.38
r186 4 36 182 $w=1.7e-07 $l=3.16938e-07 $layer=licon1_NDIFF $count=1 $X=6.135
+ $Y=0.625 $X2=6.38 $Y2=0.46
r187 3 32 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=0.235 $X2=3.86 $Y2=0.41
r188 2 28 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.68
+ $Y=0.595 $X2=2.86 $Y2=0.805
r189 1 24 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=0.71
+ $Y=0.595 $X2=0.86 $Y2=0.805
.ends

