* File: sky130_fd_sc_lp__a2111o_4.pex.spice
* Created: Fri Aug 28 09:46:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111O_4%D1 3 7 9 13 17 19 20 21 22 26
c47 21 0 8.30185e-20 $X=1.12 $Y=1.42
c48 20 0 1.47171e-19 $X=0.69 $Y=1.51
c49 3 0 7.42059e-20 $X=0.655 $Y=2.465
r50 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.51 $X2=0.37 $Y2=1.51
r51 22 26 4.11983 $w=4.48e-07 $l=1.55e-07 $layer=LI1_cond $X=0.31 $Y=1.665
+ $X2=0.31 $Y2=1.51
r52 19 25 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.58 $Y=1.51
+ $X2=0.37 $Y2=1.51
r53 19 20 6.91837 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.58 $Y=1.51
+ $X2=0.69 $Y2=1.51
r54 15 21 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.155 $Y=1.345
+ $X2=1.12 $Y2=1.42
r55 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.155 $Y=1.345
+ $X2=1.155 $Y2=0.655
r56 11 21 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.085 $Y=1.495
+ $X2=1.12 $Y2=1.42
r57 11 13 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.085 $Y=1.495
+ $X2=1.085 $Y2=2.465
r58 10 20 6.91837 $w=1.5e-07 $l=1.48324e-07 $layer=POLY_cond $X=0.8 $Y=1.42
+ $X2=0.69 $Y2=1.51
r59 9 21 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.01 $Y=1.42 $X2=1.12
+ $Y2=1.42
r60 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.01 $Y=1.42 $X2=0.8
+ $Y2=1.42
r61 5 20 18.1359 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.725 $Y=1.345
+ $X2=0.69 $Y2=1.51
r62 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.725 $Y=1.345
+ $X2=0.725 $Y2=0.655
r63 1 20 18.1359 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.655 $Y=1.675
+ $X2=0.69 $Y2=1.51
r64 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.655 $Y=1.675
+ $X2=0.655 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%C1 3 7 11 15 17 18 19 20 35
c56 20 0 2.21377e-19 $X=2.64 $Y=1.665
r57 33 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.005 $Y=1.51
+ $X2=2.095 $Y2=1.51
r58 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=1.51 $X2=2.005 $Y2=1.51
r59 31 33 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.945 $Y=1.51
+ $X2=2.005 $Y2=1.51
r60 29 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.605 $Y=1.51
+ $X2=1.945 $Y2=1.51
r61 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.605
+ $Y=1.51 $X2=1.605 $Y2=1.51
r62 27 29 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.585 $Y=1.51
+ $X2=1.605 $Y2=1.51
r63 25 27 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.515 $Y=1.51
+ $X2=1.585 $Y2=1.51
r64 19 20 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.597
+ $X2=2.64 $Y2=1.597
r65 19 34 5.17764 $w=3.43e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.597
+ $X2=2.005 $Y2=1.597
r66 18 34 10.8563 $w=3.43e-07 $l=3.25e-07 $layer=LI1_cond $X=1.68 $Y=1.597
+ $X2=2.005 $Y2=1.597
r67 18 30 2.50531 $w=3.43e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=1.597
+ $X2=1.605 $Y2=1.597
r68 17 30 13.5287 $w=3.43e-07 $l=4.05e-07 $layer=LI1_cond $X=1.2 $Y=1.597
+ $X2=1.605 $Y2=1.597
r69 13 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.345
+ $X2=2.095 $Y2=1.51
r70 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.095 $Y=1.345
+ $X2=2.095 $Y2=0.655
r71 9 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=1.675
+ $X2=1.945 $Y2=1.51
r72 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.945 $Y=1.675
+ $X2=1.945 $Y2=2.465
r73 5 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.345
+ $X2=1.585 $Y2=1.51
r74 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.585 $Y=1.345
+ $X2=1.585 $Y2=0.655
r75 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.675
+ $X2=1.515 $Y2=1.51
r76 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.515 $Y=1.675
+ $X2=1.515 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%B1 3 6 9 13 17 24 25 29 35 38
r67 34 38 8.13088 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=1.56
+ $X2=3.375 $Y2=1.56
r68 33 35 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.54 $Y=1.42 $X2=3.56
+ $Y2=1.42
r69 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.54
+ $Y=1.42 $X2=3.54 $Y2=1.42
r70 31 33 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.325 $Y=1.42
+ $X2=3.54 $Y2=1.42
r71 28 29 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.895 $Y=1.42
+ $X2=2.82 $Y2=1.42
r72 24 25 12.7582 $w=4.48e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.56 $X2=4.08
+ $Y2=1.56
r73 24 34 1.59477 $w=4.48e-07 $l=6e-08 $layer=LI1_cond $X=3.6 $Y=1.56 $X2=3.54
+ $Y2=1.56
r74 22 31 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.13 $Y=1.42
+ $X2=3.325 $Y2=1.42
r75 22 28 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.13 $Y=1.42
+ $X2=2.895 $Y2=1.42
r76 21 38 13.5864 $w=1.98e-07 $l=2.45e-07 $layer=LI1_cond $X=3.13 $Y=1.435
+ $X2=3.375 $Y2=1.435
r77 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.13
+ $Y=1.42 $X2=3.13 $Y2=1.42
r78 15 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.255
+ $X2=3.56 $Y2=1.42
r79 15 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.56 $Y=1.255 $X2=3.56
+ $Y2=0.655
r80 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.325 $Y=1.585
+ $X2=3.325 $Y2=1.42
r81 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.325 $Y=1.585
+ $X2=3.325 $Y2=2.375
r82 7 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.895 $Y=1.585
+ $X2=2.895 $Y2=1.42
r83 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.895 $Y=1.585
+ $X2=2.895 $Y2=2.375
r84 6 29 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.6 $Y=1.33 $X2=2.82
+ $Y2=1.33
r85 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.525 $Y=1.255
+ $X2=2.6 $Y2=1.33
r86 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.525 $Y=1.255 $X2=2.525
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%A1 1 3 6 8 10 12 15 17 19 20 23
c61 6 0 1.81945e-19 $X=3.99 $Y=2.375
c62 1 0 1.79874e-19 $X=3.99 $Y=1.185
r63 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.86
+ $Y=1.35 $X2=4.86 $Y2=1.35
r64 20 24 8.82722 $w=2.33e-07 $l=1.8e-07 $layer=LI1_cond $X=5.04 $Y=1.327
+ $X2=4.86 $Y2=1.327
r65 18 23 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=4.495 $Y=1.35
+ $X2=4.86 $Y2=1.35
r66 18 19 6.91837 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.495 $Y=1.35
+ $X2=4.42 $Y2=1.35
r67 13 19 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.42 $Y=1.515
+ $X2=4.42 $Y2=1.35
r68 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.42 $Y=1.515
+ $X2=4.42 $Y2=2.375
r69 10 19 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.42 $Y=1.185
+ $X2=4.42 $Y2=1.35
r70 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.42 $Y=1.185
+ $X2=4.42 $Y2=0.655
r71 9 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.065 $Y=1.26
+ $X2=3.99 $Y2=1.26
r72 8 19 6.91837 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.345 $Y=1.26
+ $X2=4.42 $Y2=1.35
r73 8 9 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.345 $Y=1.26
+ $X2=4.065 $Y2=1.26
r74 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.335
+ $X2=3.99 $Y2=1.26
r75 4 6 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=3.99 $Y=1.335
+ $X2=3.99 $Y2=2.375
r76 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.185
+ $X2=3.99 $Y2=1.26
r77 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.99 $Y=1.185 $X2=3.99
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%A2 1 3 6 8 10 13 15 21 22
c47 21 0 3.30641e-20 $X=5.685 $Y=1.35
r48 20 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.685 $Y=1.35
+ $X2=5.84 $Y2=1.35
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.685
+ $Y=1.35 $X2=5.685 $Y2=1.35
r50 17 20 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=5.41 $Y=1.35
+ $X2=5.685 $Y2=1.35
r51 15 21 8.09162 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=1.327
+ $X2=5.685 $Y2=1.327
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=1.515
+ $X2=5.84 $Y2=1.35
r53 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.84 $Y=1.515
+ $X2=5.84 $Y2=2.465
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=1.185
+ $X2=5.84 $Y2=1.35
r55 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.84 $Y=1.185
+ $X2=5.84 $Y2=0.655
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.41 $Y=1.515
+ $X2=5.41 $Y2=1.35
r57 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.41 $Y=1.515 $X2=5.41
+ $Y2=2.465
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.41 $Y=1.185
+ $X2=5.41 $Y2=1.35
r59 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.41 $Y=1.185 $X2=5.41
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%A_77_47# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 53 59 60 63 65 69 71 73 77 79 82 83 84 90 97 98 99 100 103 104 114
c193 114 0 3.30641e-20 $X=7.56 $Y=1.49
c194 84 0 1.81945e-19 $X=4.515 $Y=1.7
c195 82 0 1.79874e-19 $X=4.43 $Y=1.615
r196 111 112 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.7 $Y=1.49
+ $X2=7.13 $Y2=1.49
r197 104 106 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=6.11 $Y=1.49
+ $X2=6.11 $Y2=1.7
r198 97 98 4.56265 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.87 $Y=2.03 $X2=0.87
+ $Y2=1.93
r199 91 114 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.38 $Y=1.49
+ $X2=7.56 $Y2=1.49
r200 91 112 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.38 $Y=1.49
+ $X2=7.13 $Y2=1.49
r201 90 91 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.38
+ $Y=1.49 $X2=7.38 $Y2=1.49
r202 88 111 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.36 $Y=1.49
+ $X2=6.7 $Y2=1.49
r203 88 108 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.36 $Y=1.49
+ $X2=6.27 $Y2=1.49
r204 87 90 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.36 $Y=1.49
+ $X2=7.38 $Y2=1.49
r205 87 88 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.36
+ $Y=1.49 $X2=6.36 $Y2=1.49
r206 85 104 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.2 $Y=1.49 $X2=6.11
+ $Y2=1.49
r207 85 87 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.2 $Y=1.49
+ $X2=6.36 $Y2=1.49
r208 83 106 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.02 $Y=1.7 $X2=6.11
+ $Y2=1.7
r209 83 84 98.1872 $w=1.68e-07 $l=1.505e-06 $layer=LI1_cond $X=6.02 $Y=1.7
+ $X2=4.515 $Y2=1.7
r210 82 84 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.43 $Y=1.615
+ $X2=4.515 $Y2=1.7
r211 81 82 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.43 $Y=1.155
+ $X2=4.43 $Y2=1.615
r212 80 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.87 $Y=1.07
+ $X2=3.775 $Y2=1.07
r213 79 81 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.345 $Y=1.07
+ $X2=4.43 $Y2=1.155
r214 79 80 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.345 $Y=1.07
+ $X2=3.87 $Y2=1.07
r215 75 102 3.24837 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=3.87 $Y=0.36
+ $X2=3.775 $Y2=0.36
r216 75 77 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=3.87 $Y=0.36
+ $X2=4.635 $Y2=0.36
r217 74 103 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=0.985
+ $X2=3.775 $Y2=1.07
r218 73 102 3.59031 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=3.775 $Y=0.465
+ $X2=3.775 $Y2=0.36
r219 73 74 30.3541 $w=1.88e-07 $l=5.2e-07 $layer=LI1_cond $X=3.775 $Y=0.465
+ $X2=3.775 $Y2=0.985
r220 72 100 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.405 $Y=1.07
+ $X2=2.29 $Y2=1.07
r221 71 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.68 $Y=1.07
+ $X2=3.775 $Y2=1.07
r222 71 72 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.68 $Y=1.07
+ $X2=2.405 $Y2=1.07
r223 67 100 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.985
+ $X2=2.29 $Y2=1.07
r224 67 69 28.31 $w=2.28e-07 $l=5.65e-07 $layer=LI1_cond $X=2.29 $Y=0.985
+ $X2=2.29 $Y2=0.42
r225 66 99 6.59134 $w=1.7e-07 $l=2.69165e-07 $layer=LI1_cond $X=1.505 $Y=1.07
+ $X2=1.275 $Y2=0.985
r226 65 100 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.175 $Y=1.07
+ $X2=2.29 $Y2=1.07
r227 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.175 $Y=1.07
+ $X2=1.505 $Y2=1.07
r228 61 99 0.280307 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.39 $Y=0.985
+ $X2=1.275 $Y2=0.985
r229 61 63 28.31 $w=2.28e-07 $l=5.65e-07 $layer=LI1_cond $X=1.39 $Y=0.985
+ $X2=1.39 $Y2=0.42
r230 59 99 6.59134 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=1.15
+ $X2=1.275 $Y2=0.985
r231 59 60 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.275 $Y=1.15
+ $X2=0.935 $Y2=1.15
r232 55 60 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.82 $Y=1.15
+ $X2=0.935 $Y2=1.15
r233 55 98 34.8238 $w=2.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.82 $Y=1.235
+ $X2=0.82 $Y2=1.93
r234 51 55 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.475 $Y=1.15
+ $X2=0.82 $Y2=1.15
r235 51 53 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=0.475 $Y=1.065
+ $X2=0.475 $Y2=0.42
r236 47 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.56 $Y=1.655
+ $X2=7.56 $Y2=1.49
r237 47 49 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.56 $Y=1.655
+ $X2=7.56 $Y2=2.465
r238 43 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.56 $Y=1.325
+ $X2=7.56 $Y2=1.49
r239 43 45 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.56 $Y=1.325
+ $X2=7.56 $Y2=0.655
r240 39 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.13 $Y=1.655
+ $X2=7.13 $Y2=1.49
r241 39 41 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.13 $Y=1.655
+ $X2=7.13 $Y2=2.465
r242 35 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.13 $Y=1.325
+ $X2=7.13 $Y2=1.49
r243 35 37 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.13 $Y=1.325
+ $X2=7.13 $Y2=0.655
r244 31 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=1.655
+ $X2=6.7 $Y2=1.49
r245 31 33 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.7 $Y=1.655 $X2=6.7
+ $Y2=2.465
r246 27 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=1.325
+ $X2=6.7 $Y2=1.49
r247 27 29 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.7 $Y=1.325
+ $X2=6.7 $Y2=0.655
r248 23 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.27 $Y=1.655
+ $X2=6.27 $Y2=1.49
r249 23 25 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.27 $Y=1.655
+ $X2=6.27 $Y2=2.465
r250 19 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.27 $Y=1.325
+ $X2=6.27 $Y2=1.49
r251 19 21 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.27 $Y=1.325
+ $X2=6.27 $Y2=0.655
r252 6 97 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.835 $X2=0.87 $Y2=2.03
r253 5 77 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=4.495
+ $Y=0.235 $X2=4.635 $Y2=0.37
r254 4 102 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.635
+ $Y=0.235 $X2=3.775 $Y2=0.42
r255 3 69 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.17
+ $Y=0.235 $X2=2.31 $Y2=0.42
r256 2 63 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.23
+ $Y=0.235 $X2=1.37 $Y2=0.42
r257 1 53 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.385
+ $Y=0.235 $X2=0.51 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%A_63_367# 1 2 3 10 12 14 18 20 24 29
c32 18 0 8.30185e-20 $X=1.3 $Y=2.105
r33 22 24 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=2.195 $Y=2.905
+ $X2=2.195 $Y2=2.445
r34 21 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.395 $Y=2.99 $X2=1.3
+ $Y2=2.99
r35 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.065 $Y=2.99
+ $X2=2.195 $Y2=2.905
r36 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.065 $Y=2.99
+ $X2=1.395 $Y2=2.99
r37 16 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.905 $X2=1.3
+ $Y2=2.99
r38 16 18 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=1.3 $Y=2.905 $X2=1.3
+ $Y2=2.105
r39 15 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.535 $Y=2.99
+ $X2=0.405 $Y2=2.99
r40 14 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.205 $Y=2.99 $X2=1.3
+ $Y2=2.99
r41 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.205 $Y=2.99
+ $X2=0.535 $Y2=2.99
r42 10 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.405 $Y=2.905
+ $X2=0.405 $Y2=2.99
r43 10 12 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.405 $Y=2.905
+ $X2=0.405 $Y2=2.085
r44 3 24 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=2.02
+ $Y=1.835 $X2=2.16 $Y2=2.445
r45 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.835 $X2=1.3 $Y2=2.91
r46 2 18 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.835 $X2=1.3 $Y2=2.105
r47 1 27 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=1.835 $X2=0.44 $Y2=2.91
r48 1 12 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=1.835 $X2=0.44 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%A_318_367# 1 2 9 13 16 18
r26 20 21 4.6142 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=2.025
+ $X2=3.085 $Y2=2.11
r27 18 20 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.085 $Y=1.87
+ $X2=3.085 $Y2=2.025
r28 13 21 5.83732 $w=1.88e-07 $l=1e-07 $layer=LI1_cond $X=3.11 $Y=2.21 $X2=3.11
+ $Y2=2.11
r29 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=2.025
+ $X2=1.73 $Y2=2.025
r30 9 20 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.965 $Y=2.025
+ $X2=3.085 $Y2=2.025
r31 9 10 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=2.965 $Y=2.025
+ $X2=1.895 $Y2=2.025
r32 2 18 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.745 $X2=3.11 $Y2=1.87
r33 2 13 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=2.97
+ $Y=1.745 $X2=3.11 $Y2=2.21
r34 1 16 300 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.835 $X2=1.73 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%A_511_349# 1 2 3 4 15 17 18 19 22 23 27 29
+ 33 40
r53 33 35 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=5.625 $Y=2.17
+ $X2=5.625 $Y2=2.85
r54 31 33 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=5.625 $Y=2.125
+ $X2=5.625 $Y2=2.17
r55 30 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.8 $Y=2.04 $X2=4.67
+ $Y2=2.04
r56 29 31 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.53 $Y=2.04
+ $X2=5.625 $Y2=2.125
r57 29 30 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.53 $Y=2.04 $X2=4.8
+ $Y2=2.04
r58 25 40 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.67 $Y=2.125
+ $X2=4.67 $Y2=2.04
r59 25 27 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=4.67 $Y=2.125
+ $X2=4.67 $Y2=2.46
r60 24 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=2.04
+ $X2=3.66 $Y2=2.04
r61 23 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.54 $Y=2.04 $X2=4.67
+ $Y2=2.04
r62 23 24 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=4.54 $Y=2.04
+ $X2=3.825 $Y2=2.04
r63 20 22 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=3.66 $Y=2.905
+ $X2=3.66 $Y2=2.445
r64 19 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=2.125 $X2=3.66
+ $Y2=2.04
r65 19 22 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.66 $Y=2.125
+ $X2=3.66 $Y2=2.445
r66 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.495 $Y=2.99
+ $X2=3.66 $Y2=2.905
r67 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.495 $Y=2.99
+ $X2=2.845 $Y2=2.99
r68 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.68 $Y=2.905
+ $X2=2.845 $Y2=2.99
r69 13 15 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=2.68 $Y=2.905
+ $X2=2.68 $Y2=2.385
r70 4 35 400 $w=1.7e-07 $l=1.08274e-06 $layer=licon1_PDIFF $count=1 $X=5.485
+ $Y=1.835 $X2=5.625 $Y2=2.85
r71 4 33 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=5.485
+ $Y=1.835 $X2=5.625 $Y2=2.17
r72 3 40 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.745 $X2=4.635 $Y2=2.04
r73 3 27 300 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=2 $X=4.495
+ $Y=1.745 $X2=4.635 $Y2=2.46
r74 2 38 600 $w=1.7e-07 $l=4.04629e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.745 $X2=3.66 $Y2=2.04
r75 2 22 300 $w=1.7e-07 $l=8.19756e-07 $layer=licon1_PDIFF $count=2 $X=3.4
+ $Y=1.745 $X2=3.66 $Y2=2.445
r76 1 15 300 $w=1.7e-07 $l=6.99714e-07 $layer=licon1_PDIFF $count=2 $X=2.555
+ $Y=1.745 $X2=2.68 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%VPWR 1 2 3 4 5 18 20 24 28 34 38 40 44 46
+ 51 56 61 67 70 73 76 80
r107 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r110 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r112 65 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r113 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.08 $Y=3.33
+ $X2=6.915 $Y2=3.33
r115 62 64 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.08 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 61 79 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.885 $Y2=3.33
r117 61 64 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r120 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.22 $Y=3.33
+ $X2=6.055 $Y2=3.33
r122 57 59 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.22 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.75 $Y=3.33
+ $X2=6.915 $Y2=3.33
r124 56 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.75 $Y=3.33
+ $X2=6.48 $Y2=3.33
r125 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r126 55 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r127 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 52 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.195 $Y2=3.33
r129 52 54 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.52 $Y2=3.33
r130 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=6.055 $Y2=3.33
r131 51 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=5.52 $Y2=3.33
r132 48 49 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 46 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=3.33
+ $X2=4.205 $Y2=3.33
r134 46 48 247.914 $w=1.68e-07 $l=3.8e-06 $layer=LI1_cond $X=4.04 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 44 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r136 44 49 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 44 67 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 40 43 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=7.775 $Y=2.19
+ $X2=7.775 $Y2=2.95
r139 38 79 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.775 $Y=3.245
+ $X2=7.885 $Y2=3.33
r140 38 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.775 $Y=3.245
+ $X2=7.775 $Y2=2.95
r141 34 37 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.915 $Y=2.18
+ $X2=6.915 $Y2=2.95
r142 32 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=3.245
+ $X2=6.915 $Y2=3.33
r143 32 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.915 $Y=3.245
+ $X2=6.915 $Y2=2.95
r144 28 31 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=6.055 $Y=2.04
+ $X2=6.055 $Y2=2.95
r145 26 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=3.245
+ $X2=6.055 $Y2=3.33
r146 26 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.055 $Y=3.245
+ $X2=6.055 $Y2=2.95
r147 22 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.195 $Y=3.245
+ $X2=5.195 $Y2=3.33
r148 22 24 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=5.195 $Y=3.245
+ $X2=5.195 $Y2=2.42
r149 21 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.205 $Y2=3.33
r150 20 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.03 $Y=3.33
+ $X2=5.195 $Y2=3.33
r151 20 21 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.03 $Y=3.33
+ $X2=4.37 $Y2=3.33
r152 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=3.245
+ $X2=4.205 $Y2=3.33
r153 16 18 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.205 $Y=3.245
+ $X2=4.205 $Y2=2.42
r154 5 43 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.835 $X2=7.775 $Y2=2.95
r155 5 40 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.835 $X2=7.775 $Y2=2.19
r156 4 37 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.835 $X2=6.915 $Y2=2.95
r157 4 34 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.835 $X2=6.915 $Y2=2.18
r158 3 31 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.915
+ $Y=1.835 $X2=6.055 $Y2=2.95
r159 3 28 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.915
+ $Y=1.835 $X2=6.055 $Y2=2.04
r160 2 24 300 $w=1.7e-07 $l=6.44477e-07 $layer=licon1_PDIFF $count=2 $X=5.07
+ $Y=1.835 $X2=5.195 $Y2=2.42
r161 1 18 300 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_PDIFF $count=2 $X=4.065
+ $Y=1.745 $X2=4.205 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41
+ 42 43 44 49 50 52 56
r62 50 56 2.56098 $w=3.58e-07 $l=8e-08 $layer=LI1_cond $X=7.895 $Y=1.745
+ $X2=7.895 $Y2=1.665
r63 49 52 1.92074 $w=3.58e-07 $l=6e-08 $layer=LI1_cond $X=7.895 $Y=1.235
+ $X2=7.895 $Y2=1.295
r64 44 50 2.61705 $w=3.6e-07 $l=9e-08 $layer=LI1_cond $X=7.895 $Y=1.835
+ $X2=7.895 $Y2=1.745
r65 44 56 0.0960369 $w=3.58e-07 $l=3e-09 $layer=LI1_cond $X=7.895 $Y=1.662
+ $X2=7.895 $Y2=1.665
r66 43 49 2.57345 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.895 $Y=1.15
+ $X2=7.895 $Y2=1.235
r67 43 44 11.3644 $w=3.58e-07 $l=3.55e-07 $layer=LI1_cond $X=7.895 $Y=1.307
+ $X2=7.895 $Y2=1.662
r68 43 52 0.384148 $w=3.58e-07 $l=1.2e-08 $layer=LI1_cond $X=7.895 $Y=1.307
+ $X2=7.895 $Y2=1.295
r69 40 42 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.44 $Y=1.835
+ $X2=7.345 $Y2=1.835
r70 39 44 5.2341 $w=1.8e-07 $l=1.8e-07 $layer=LI1_cond $X=7.715 $Y=1.835
+ $X2=7.895 $Y2=1.835
r71 39 40 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=1.835
+ $X2=7.44 $Y2=1.835
r72 38 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.44 $Y=1.15
+ $X2=7.345 $Y2=1.15
r73 37 43 5.44966 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=7.715 $Y=1.15
+ $X2=7.895 $Y2=1.15
r74 37 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=1.15
+ $X2=7.44 $Y2=1.15
r75 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=7.345 $Y=1.98
+ $X2=7.345 $Y2=2.91
r76 31 42 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=7.345 $Y=1.925
+ $X2=7.345 $Y2=1.835
r77 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=7.345 $Y=1.925
+ $X2=7.345 $Y2=1.98
r78 27 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=1.065
+ $X2=7.345 $Y2=1.15
r79 27 29 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=7.345 $Y=1.065
+ $X2=7.345 $Y2=0.42
r80 25 42 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.25 $Y=1.835
+ $X2=7.345 $Y2=1.835
r81 25 26 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.25 $Y=1.835
+ $X2=6.58 $Y2=1.835
r82 23 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.25 $Y=1.15
+ $X2=7.345 $Y2=1.15
r83 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.25 $Y=1.15
+ $X2=6.58 $Y2=1.15
r84 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.485 $Y=1.98
+ $X2=6.485 $Y2=2.91
r85 17 26 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=6.485 $Y=1.925
+ $X2=6.58 $Y2=1.835
r86 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.485 $Y=1.925
+ $X2=6.485 $Y2=1.98
r87 13 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.485 $Y=1.065
+ $X2=6.58 $Y2=1.15
r88 13 15 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=6.485 $Y=1.065
+ $X2=6.485 $Y2=0.42
r89 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.205
+ $Y=1.835 $X2=7.345 $Y2=2.91
r90 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.205
+ $Y=1.835 $X2=7.345 $Y2=1.98
r91 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=1.835 $X2=6.485 $Y2=2.91
r92 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=1.835 $X2=6.485 $Y2=1.98
r93 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.205
+ $Y=0.235 $X2=7.345 $Y2=0.42
r94 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.345
+ $Y=0.235 $X2=6.485 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%VGND 1 2 3 4 5 6 7 24 26 30 36 40 44 46 48
+ 50 51 52 58 63 68 73 79 84 90 92 95 98 102
r120 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r121 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r122 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r123 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r124 89 90 12.2732 $w=8.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=0.365
+ $X2=3.51 $Y2=0.365
r125 86 89 3.05 $w=8.98e-07 $l=2.25e-07 $layer=LI1_cond $X=3.12 $Y=0.365
+ $X2=3.345 $Y2=0.365
r126 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r127 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r128 82 86 6.50667 $w=8.98e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0.365
+ $X2=3.12 $Y2=0.365
r129 82 84 10.9176 $w=8.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.64 $Y=0.365
+ $X2=2.575 $Y2=0.365
r130 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r131 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r132 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r133 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r134 77 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r135 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r136 74 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=6.915
+ $Y2=0
r137 74 76 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=7.44
+ $Y2=0
r138 73 101 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=7.61 $Y=0
+ $X2=7.885 $Y2=0
r139 73 76 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.61 $Y=0 $X2=7.44
+ $Y2=0
r140 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r141 72 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r142 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r143 69 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.22 $Y=0 $X2=6.055
+ $Y2=0
r144 69 71 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.22 $Y=0 $X2=6.48
+ $Y2=0
r145 68 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.75 $Y=0 $X2=6.915
+ $Y2=0
r146 68 71 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.75 $Y=0 $X2=6.48
+ $Y2=0
r147 67 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r148 67 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r149 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r150 64 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.195
+ $Y2=0
r151 64 66 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.52
+ $Y2=0
r152 63 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=0 $X2=6.055
+ $Y2=0
r153 63 66 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.89 $Y=0 $X2=5.52
+ $Y2=0
r154 62 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r155 61 90 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.51
+ $Y2=0
r156 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r157 58 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.03 $Y=0 $X2=5.195
+ $Y2=0
r158 58 61 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=5.03 $Y=0 $X2=3.6
+ $Y2=0
r159 56 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r160 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r161 52 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r162 52 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r163 50 55 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.72
+ $Y2=0
r164 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.94
+ $Y2=0
r165 46 101 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.775 $Y=0.085
+ $X2=7.885 $Y2=0
r166 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.775 $Y=0.085
+ $X2=7.775 $Y2=0.38
r167 42 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0
r168 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0.36
r169 38 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=0.085
+ $X2=6.055 $Y2=0
r170 38 40 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.055 $Y=0.085
+ $X2=6.055 $Y2=0.36
r171 34 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.195 $Y=0.085
+ $X2=5.195 $Y2=0
r172 34 36 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=5.195 $Y=0.085
+ $X2=5.195 $Y2=0.465
r173 33 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.84
+ $Y2=0
r174 33 84 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.575 $Y2=0
r175 28 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r176 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.36
r177 27 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=0.94
+ $Y2=0
r178 26 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.84
+ $Y2=0
r179 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.675 $Y=0
+ $X2=1.105 $Y2=0
r180 22 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=0.085
+ $X2=0.94 $Y2=0
r181 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.94 $Y=0.085
+ $X2=0.94 $Y2=0.38
r182 7 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.635
+ $Y=0.235 $X2=7.775 $Y2=0.38
r183 6 44 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.775
+ $Y=0.235 $X2=6.915 $Y2=0.36
r184 5 40 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.915
+ $Y=0.235 $X2=6.055 $Y2=0.36
r185 4 36 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.235 $X2=5.195 $Y2=0.465
r186 3 89 45.5 $w=1.7e-07 $l=8.05078e-07 $layer=licon1_NDIFF $count=4 $X=2.6
+ $Y=0.235 $X2=3.345 $Y2=0.36
r187 2 30 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=1.66
+ $Y=0.235 $X2=1.84 $Y2=0.36
r188 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.8
+ $Y=0.235 $X2=0.94 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_4%A_813_47# 1 2 11 13 15 17 18
r31 17 18 8.66869 $w=2.78e-07 $l=1.75e-07 $layer=LI1_cond $X=4.685 $Y=0.837
+ $X2=4.86 $Y2=0.837
r32 13 20 4.25761 $w=1.9e-07 $l=1.4e-07 $layer=LI1_cond $X=5.625 $Y=0.76
+ $X2=5.625 $Y2=0.9
r33 13 15 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=5.625 $Y=0.76
+ $X2=5.625 $Y2=0.42
r34 11 20 2.88909 $w=2.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.53 $Y=0.9 $X2=5.625
+ $Y2=0.9
r35 11 18 27.5763 $w=2.78e-07 $l=6.7e-07 $layer=LI1_cond $X=5.53 $Y=0.9 $X2=4.86
+ $Y2=0.9
r36 9 17 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=4.205 $Y=0.725
+ $X2=4.685 $Y2=0.725
r37 2 20 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=5.485
+ $Y=0.235 $X2=5.625 $Y2=0.875
r38 2 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.485
+ $Y=0.235 $X2=5.625 $Y2=0.42
r39 1 9 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=4.065
+ $Y=0.235 $X2=4.205 $Y2=0.72
.ends

