* File: sky130_fd_sc_lp__o22a_0.spice
* Created: Wed Sep  2 10:19:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22a_0.pex.spice"
.subckt sky130_fd_sc_lp__o22a_0  VNB VPB A1 B1 B2 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* B2	B2
* B1	B1
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_80_313#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1323 AS=0.1113 PD=1.05 PS=1.37 NRD=9.996 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1002 N_A_286_125#_M1002_d N_A1_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1323 PD=0.7 PS=1.05 NRD=0 NRS=89.988 M=1 R=2.8 SA=75001
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_80_313#_M1003_d N_B1_M1003_g N_A_286_125#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.0588 PD=0.72 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_286_125#_M1004_d N_B2_M1004_g N_A_80_313#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.063 PD=0.78 PS=0.72 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.8 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_286_125#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1533 AS=0.0756 PD=1.57 PS=0.78 NRD=22.848 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_80_313#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.3712 AS=0.1696 PD=1.8 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1007 A_372_489# N_B1_M1007_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.3712 PD=0.88 PS=1.8 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1001 N_A_80_313#_M1001_d N_B2_M1001_g A_372_489# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.9
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 A_536_489# N_A2_M1009_g N_A_80_313#_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1216 AS=0.0896 PD=1.02 PS=0.92 NRD=41.5473 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_536_489# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1216 PD=1.81 PS=1.02 NRD=0 NRS=41.5473 M=1 R=4.26667 SA=75002.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_82 VPB 0 1.12607e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o22a_0.pxi.spice"
*
.ends
*
*
