* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_85_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 X a_85_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_342_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR A1 a_342_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND A3 a_355_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_355_49# A2 a_427_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 X a_85_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_342_367# B1 a_85_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR A3 a_342_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND a_85_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_427_49# A1 a_85_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_85_23# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
