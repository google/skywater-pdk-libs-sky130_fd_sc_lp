* File: sky130_fd_sc_lp__o2111ai_0.pxi.spice
* Created: Wed Sep  2 10:12:52 2020
* 
x_PM_SKY130_FD_SC_LP__O2111AI_0%D1 N_D1_M1003_g N_D1_M1006_g N_D1_c_74_n
+ N_D1_c_75_n N_D1_c_76_n D1 D1 D1 N_D1_c_78_n PM_SKY130_FD_SC_LP__O2111AI_0%D1
x_PM_SKY130_FD_SC_LP__O2111AI_0%C1 N_C1_M1000_g N_C1_M1007_g N_C1_c_112_n C1 C1
+ C1 C1 N_C1_c_114_n PM_SKY130_FD_SC_LP__O2111AI_0%C1
x_PM_SKY130_FD_SC_LP__O2111AI_0%B1 N_B1_M1009_g N_B1_c_159_n N_B1_c_160_n
+ N_B1_c_166_n N_B1_c_167_n N_B1_M1002_g B1 B1 B1 N_B1_c_162_n N_B1_c_163_n
+ N_B1_c_164_n PM_SKY130_FD_SC_LP__O2111AI_0%B1
x_PM_SKY130_FD_SC_LP__O2111AI_0%A2 N_A2_M1001_g N_A2_c_218_n N_A2_M1005_g
+ N_A2_c_219_n A2 A2 A2 A2 A2 N_A2_c_221_n A2 PM_SKY130_FD_SC_LP__O2111AI_0%A2
x_PM_SKY130_FD_SC_LP__O2111AI_0%A1 N_A1_c_272_n N_A1_M1004_g N_A1_M1008_g
+ N_A1_c_273_n N_A1_c_274_n N_A1_c_279_n N_A1_c_275_n A1 A1 A1 N_A1_c_277_n
+ PM_SKY130_FD_SC_LP__O2111AI_0%A1
x_PM_SKY130_FD_SC_LP__O2111AI_0%VPWR N_VPWR_M1003_s N_VPWR_M1000_d
+ N_VPWR_M1008_d N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n
+ N_VPWR_c_315_n VPWR N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n
+ N_VPWR_c_310_n PM_SKY130_FD_SC_LP__O2111AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O2111AI_0%Y N_Y_M1006_s N_Y_M1003_d N_Y_M1002_d
+ N_Y_c_351_n N_Y_c_352_n N_Y_c_363_n N_Y_c_354_n N_Y_c_355_n N_Y_c_356_n
+ N_Y_c_357_n Y Y Y Y Y PM_SKY130_FD_SC_LP__O2111AI_0%Y
x_PM_SKY130_FD_SC_LP__O2111AI_0%A_339_47# N_A_339_47#_M1009_d
+ N_A_339_47#_M1004_d N_A_339_47#_c_416_n N_A_339_47#_c_437_p
+ N_A_339_47#_c_412_n N_A_339_47#_c_413_n N_A_339_47#_c_414_n
+ N_A_339_47#_c_415_n PM_SKY130_FD_SC_LP__O2111AI_0%A_339_47#
x_PM_SKY130_FD_SC_LP__O2111AI_0%VGND N_VGND_M1001_d N_VGND_c_445_n VGND
+ N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n
+ PM_SKY130_FD_SC_LP__O2111AI_0%VGND
cc_1 VNB N_D1_M1003_g 0.012287f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.645
cc_2 VNB N_D1_c_74_n 0.0194614f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=0.765
cc_3 VNB N_D1_c_75_n 0.0339492f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=0.915
cc_4 VNB N_D1_c_76_n 0.0195476f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.435
cc_5 VNB D1 0.00700254f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_D1_c_78_n 0.0261094f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_7 VNB N_C1_M1007_g 0.0299323f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=0.445
cc_8 VNB N_C1_c_112_n 0.0340284f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.435
cc_9 VNB C1 0.00694535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_C1_c_114_n 0.0165311f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.93
cc_11 VNB N_B1_c_159_n 0.0154273f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=0.765
cc_12 VNB N_B1_c_160_n 0.0117757f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=0.445
cc_13 VNB B1 0.00940018f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_14 VNB N_B1_c_162_n 0.0280014f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_15 VNB N_B1_c_163_n 0.0183174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_164_n 0.0165735f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.295
cc_17 VNB N_A2_M1001_g 0.0409153f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.645
cc_18 VNB N_A2_c_218_n 0.0211702f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=0.445
cc_19 VNB N_A2_c_219_n 0.00241f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.253
cc_20 VNB A2 0.00587781f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.435
cc_21 VNB N_A2_c_221_n 0.0223185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A2 4.40518e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_272_n 0.0194865f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.435
cc_24 VNB N_A1_c_273_n 0.0221147f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.253
cc_25 VNB N_A1_c_274_n 0.00192438f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_A1_c_275_n 0.0393825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A1 0.0224645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_c_277_n 0.0182244f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.93
cc_29 VNB N_VPWR_c_310_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_351_n 0.0517457f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.253
cc_31 VNB N_Y_c_352_n 0.0140333f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.435
cc_32 VNB N_A_339_47#_c_412_n 0.00275974f $X=-0.19 $Y=-0.245 $X2=0.612 $Y2=1.435
cc_33 VNB N_A_339_47#_c_413_n 0.0187111f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_34 VNB N_A_339_47#_c_414_n 0.0124364f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_35 VNB N_A_339_47#_c_415_n 0.0199312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_445_n 0.00527728f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=0.445
cc_37 VNB N_VGND_c_446_n 0.0662179f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=0.915
cc_38 VNB N_VGND_c_447_n 0.0192415f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_39 VNB N_VGND_c_448_n 0.194638f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.93
cc_40 VNB N_VGND_c_449_n 0.00516809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_D1_M1003_g 0.0532152f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.645
cc_42 VPB D1 0.00262414f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_43 VPB N_C1_M1000_g 0.0427582f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.645
cc_44 VPB N_C1_c_112_n 0.0234864f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.435
cc_45 VPB N_B1_c_160_n 0.0257222f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=0.445
cc_46 VPB N_B1_c_166_n 0.0209301f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=0.915
cc_47 VPB N_B1_c_167_n 0.0126217f $X=-0.19 $Y=1.655 $X2=0.702 $Y2=0.765
cc_48 VPB N_B1_M1002_g 0.0229526f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.435
cc_49 VPB B1 0.00289575f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_50 VPB N_A2_M1005_g 0.0382183f $X=-0.19 $Y=1.655 $X2=0.702 $Y2=0.765
cc_51 VPB N_A2_c_219_n 0.0232162f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.253
cc_52 VPB A2 0.00558807f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_53 VPB A2 8.47151e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A1_c_274_n 0.0338401f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_55 VPB N_A1_c_279_n 0.050794f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_56 VPB A1 0.0176359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_311_n 0.0115481f $X=-0.19 $Y=1.655 $X2=0.702 $Y2=0.915
cc_58 VPB N_VPWR_c_312_n 0.0405493f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.435
cc_59 VPB N_VPWR_c_313_n 0.0218302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_314_n 0.0111988f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=0.93
cc_61 VPB N_VPWR_c_315_n 0.0375567f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_62 VPB N_VPWR_c_316_n 0.0181712f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.93
cc_63 VPB N_VPWR_c_317_n 0.0280092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_318_n 0.0167083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_310_n 0.0596337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_Y_c_351_n 0.0141969f $X=-0.19 $Y=1.655 $X2=0.612 $Y2=1.253
cc_67 VPB N_Y_c_354_n 0.00345041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_Y_c_355_n 0.00952805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_Y_c_356_n 0.00372259f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.93
cc_70 VPB N_Y_c_357_n 0.0337564f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.925
cc_71 VPB Y 0.00219217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB Y 0.00238156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 N_D1_c_74_n N_C1_M1007_g 0.0498894f $X=0.702 $Y=0.765 $X2=0 $Y2=0
cc_74 D1 N_C1_M1007_g 7.62652e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_75 N_D1_c_78_n N_C1_M1007_g 0.00689633f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_76 N_D1_M1003_g N_C1_c_112_n 0.0410448f $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_77 N_D1_c_76_n N_C1_c_112_n 0.00735404f $X=0.612 $Y=1.435 $X2=0 $Y2=0
cc_78 D1 N_C1_c_112_n 0.00355573f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_79 N_D1_M1003_g C1 2.67696e-19 $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_80 N_D1_c_74_n C1 0.00488693f $X=0.702 $Y=0.765 $X2=0 $Y2=0
cc_81 D1 C1 0.0804931f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_82 N_D1_c_78_n C1 0.00107759f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_83 D1 N_C1_c_114_n 0.00348581f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_D1_c_78_n N_C1_c_114_n 0.00735404f $X=0.63 $Y=0.93 $X2=0 $Y2=0
cc_85 N_D1_M1003_g N_VPWR_c_312_n 0.00418138f $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_86 N_D1_M1003_g N_VPWR_c_316_n 0.00460962f $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_87 N_D1_M1003_g N_VPWR_c_310_n 0.00904175f $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_88 N_D1_c_74_n N_Y_c_351_n 0.00230936f $X=0.702 $Y=0.765 $X2=0 $Y2=0
cc_89 N_D1_c_75_n N_Y_c_351_n 0.0320775f $X=0.702 $Y=0.915 $X2=0 $Y2=0
cc_90 D1 N_Y_c_351_n 0.0739756f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_91 N_D1_c_74_n N_Y_c_363_n 0.004601f $X=0.702 $Y=0.765 $X2=0 $Y2=0
cc_92 N_D1_c_75_n N_Y_c_363_n 0.00701911f $X=0.702 $Y=0.915 $X2=0 $Y2=0
cc_93 D1 N_Y_c_363_n 0.021752f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_94 N_D1_M1003_g N_Y_c_354_n 0.017474f $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_95 D1 N_Y_c_354_n 0.00217503f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_96 N_D1_M1003_g Y 0.00213566f $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_97 N_D1_c_76_n Y 8.14888e-19 $X=0.612 $Y=1.435 $X2=0 $Y2=0
cc_98 D1 Y 0.0269971f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_99 N_D1_M1003_g Y 0.0165333f $X=0.505 $Y=2.645 $X2=0 $Y2=0
cc_100 N_D1_c_74_n N_VGND_c_446_n 0.0054833f $X=0.702 $Y=0.765 $X2=0 $Y2=0
cc_101 N_D1_c_74_n N_VGND_c_448_n 0.0108543f $X=0.702 $Y=0.765 $X2=0 $Y2=0
cc_102 D1 N_VGND_c_448_n 9.96193e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_103 N_C1_M1007_g N_B1_c_159_n 0.00624792f $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_104 C1 N_B1_c_159_n 0.00107324f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_105 N_C1_c_114_n N_B1_c_159_n 0.0141749f $X=1.2 $Y=1.32 $X2=0 $Y2=0
cc_106 N_C1_M1000_g N_B1_c_160_n 0.0076134f $X=0.935 $Y=2.645 $X2=0 $Y2=0
cc_107 N_C1_c_112_n N_B1_c_160_n 0.0141749f $X=1.2 $Y=1.645 $X2=0 $Y2=0
cc_108 N_C1_M1007_g B1 0.00120242f $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_109 C1 B1 0.0816542f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_110 N_C1_c_114_n B1 0.00354682f $X=1.2 $Y=1.32 $X2=0 $Y2=0
cc_111 C1 N_B1_c_162_n 8.83444e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_112 N_C1_M1007_g N_B1_c_163_n 0.0583926f $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_113 C1 N_B1_c_163_n 0.00186865f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_114 N_C1_c_112_n N_B1_c_164_n 0.0141749f $X=1.2 $Y=1.645 $X2=0 $Y2=0
cc_115 N_C1_M1000_g N_VPWR_c_313_n 0.00434487f $X=0.935 $Y=2.645 $X2=0 $Y2=0
cc_116 N_C1_M1000_g N_VPWR_c_316_n 0.00438034f $X=0.935 $Y=2.645 $X2=0 $Y2=0
cc_117 N_C1_M1000_g N_VPWR_c_310_n 0.00838015f $X=0.935 $Y=2.645 $X2=0 $Y2=0
cc_118 C1 N_Y_c_351_n 0.00498556f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_119 N_C1_M1007_g N_Y_c_363_n 6.401e-19 $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_120 C1 N_Y_c_363_n 0.0169266f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_121 N_C1_M1000_g N_Y_c_357_n 0.0155689f $X=0.935 $Y=2.645 $X2=0 $Y2=0
cc_122 N_C1_c_112_n N_Y_c_357_n 0.0100371f $X=1.2 $Y=1.645 $X2=0 $Y2=0
cc_123 C1 N_Y_c_357_n 0.0262109f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_124 N_C1_M1000_g Y 0.00337072f $X=0.935 $Y=2.645 $X2=0 $Y2=0
cc_125 N_C1_M1000_g Y 0.0166864f $X=0.935 $Y=2.645 $X2=0 $Y2=0
cc_126 C1 A_195_47# 0.0038957f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_127 N_C1_M1007_g N_A_339_47#_c_416_n 7.12782e-19 $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_128 C1 N_A_339_47#_c_412_n 0.00421139f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_129 N_C1_M1007_g N_VGND_c_446_n 0.00381508f $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_130 C1 N_VGND_c_446_n 0.011075f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_131 N_C1_M1007_g N_VGND_c_448_n 0.0051708f $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_132 C1 N_VGND_c_448_n 0.0111988f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_133 B1 N_A2_M1001_g 0.00226025f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_134 N_B1_c_162_n N_A2_M1001_g 0.00706928f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_135 N_B1_c_163_n N_A2_M1001_g 0.00403848f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_136 N_B1_c_160_n N_A2_c_218_n 0.00785911f $X=1.682 $Y=2.035 $X2=0 $Y2=0
cc_137 B1 N_A2_c_218_n 0.00289248f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_138 N_B1_c_164_n N_A2_c_218_n 0.00706928f $X=1.77 $Y=1.27 $X2=0 $Y2=0
cc_139 N_B1_c_160_n N_A2_M1005_g 0.0037997f $X=1.682 $Y=2.035 $X2=0 $Y2=0
cc_140 N_B1_c_166_n N_A2_M1005_g 0.0142871f $X=1.97 $Y=2.11 $X2=0 $Y2=0
cc_141 N_B1_c_159_n A2 0.00109048f $X=1.755 $Y=1.255 $X2=0 $Y2=0
cc_142 N_B1_c_160_n A2 3.41018e-19 $X=1.682 $Y=2.035 $X2=0 $Y2=0
cc_143 B1 A2 0.0199993f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_144 N_B1_c_166_n A2 4.25848e-19 $X=1.97 $Y=2.11 $X2=0 $Y2=0
cc_145 N_B1_c_159_n N_A2_c_221_n 0.00706928f $X=1.755 $Y=1.255 $X2=0 $Y2=0
cc_146 N_B1_c_167_n N_VPWR_c_313_n 0.00913859f $X=1.79 $Y=2.11 $X2=0 $Y2=0
cc_147 N_B1_M1002_g N_VPWR_c_313_n 0.00600275f $X=2.045 $Y=2.645 $X2=0 $Y2=0
cc_148 N_B1_M1002_g N_VPWR_c_317_n 0.00438034f $X=2.045 $Y=2.645 $X2=0 $Y2=0
cc_149 N_B1_M1002_g N_VPWR_c_310_n 0.00838908f $X=2.045 $Y=2.645 $X2=0 $Y2=0
cc_150 N_B1_c_166_n N_Y_c_356_n 0.0036208f $X=1.97 $Y=2.11 $X2=0 $Y2=0
cc_151 N_B1_M1002_g N_Y_c_356_n 0.0141426f $X=2.045 $Y=2.645 $X2=0 $Y2=0
cc_152 N_B1_c_160_n N_Y_c_357_n 0.00779323f $X=1.682 $Y=2.035 $X2=0 $Y2=0
cc_153 N_B1_c_166_n N_Y_c_357_n 0.0161058f $X=1.97 $Y=2.11 $X2=0 $Y2=0
cc_154 N_B1_c_167_n N_Y_c_357_n 0.00485781f $X=1.79 $Y=2.11 $X2=0 $Y2=0
cc_155 B1 N_Y_c_357_n 0.0250764f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_156 N_B1_c_164_n N_Y_c_357_n 0.00149321f $X=1.77 $Y=1.27 $X2=0 $Y2=0
cc_157 N_B1_c_167_n Y 3.27852e-19 $X=1.79 $Y=2.11 $X2=0 $Y2=0
cc_158 B1 N_A_339_47#_c_416_n 0.0137619f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_159 N_B1_c_162_n N_A_339_47#_c_416_n 0.00456035f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_160 N_B1_c_163_n N_A_339_47#_c_416_n 0.005985f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_161 B1 N_A_339_47#_c_412_n 0.0010763f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_162 N_B1_c_163_n N_A_339_47#_c_412_n 0.00158452f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_163 B1 N_A_339_47#_c_414_n 0.0137021f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_164 N_B1_c_162_n N_A_339_47#_c_414_n 0.00168937f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_165 N_B1_c_163_n N_VGND_c_446_n 0.00518687f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_166 B1 N_VGND_c_448_n 0.00432965f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_167 N_B1_c_163_n N_VGND_c_448_n 0.00659148f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_168 N_A2_M1001_g N_A1_c_272_n 0.0191155f $X=2.39 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A2_M1005_g N_A1_c_274_n 0.00834547f $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_170 N_A2_c_219_n N_A1_c_274_n 0.0135799f $X=2.515 $Y=1.825 $X2=0 $Y2=0
cc_171 A2 N_A1_c_274_n 0.00209999f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_172 N_A2_M1005_g N_A1_c_279_n 0.0609861f $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_173 A2 N_A1_c_279_n 0.0073817f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_174 N_A2_M1001_g N_A1_c_275_n 0.00740398f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_175 A2 N_A1_c_275_n 0.00209999f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A2_c_221_n N_A1_c_275_n 0.0135799f $X=2.55 $Y=1.32 $X2=0 $Y2=0
cc_177 N_A2_M1005_g A1 2.69535e-19 $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_178 A2 A1 0.058861f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A2_c_221_n A1 6.86848e-19 $X=2.55 $Y=1.32 $X2=0 $Y2=0
cc_180 N_A2_c_218_n N_A1_c_277_n 0.0135799f $X=2.515 $Y=1.625 $X2=0 $Y2=0
cc_181 A2 N_A1_c_277_n 0.00209999f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_182 N_A2_M1005_g N_VPWR_c_315_n 0.00112226f $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_183 A2 N_VPWR_c_315_n 0.0255918f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_184 N_A2_M1005_g N_VPWR_c_317_n 0.00381391f $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_185 A2 N_VPWR_c_317_n 0.0101914f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_186 N_A2_M1005_g N_VPWR_c_310_n 0.00647042f $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_187 A2 N_VPWR_c_310_n 0.00840595f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_188 N_A2_M1005_g N_Y_c_356_n 0.00349483f $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_189 A2 N_Y_c_356_n 0.0639099f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_190 N_A2_M1005_g N_Y_c_357_n 0.00165431f $X=2.525 $Y=2.645 $X2=0 $Y2=0
cc_191 N_A2_c_219_n N_Y_c_357_n 0.00203223f $X=2.515 $Y=1.825 $X2=0 $Y2=0
cc_192 A2 N_Y_c_357_n 0.0140298f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_193 N_A2_M1001_g N_A_339_47#_c_412_n 0.00239469f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A2_M1001_g N_A_339_47#_c_413_n 0.0142086f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_195 A2 N_A_339_47#_c_413_n 0.026075f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A2_c_221_n N_A_339_47#_c_413_n 0.00167312f $X=2.55 $Y=1.32 $X2=0 $Y2=0
cc_197 N_A2_M1001_g N_VGND_c_445_n 0.00320453f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_198 N_A2_M1001_g N_VGND_c_446_n 0.00585385f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A2_M1001_g N_VGND_c_448_n 0.00684443f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_200 N_A1_c_279_n N_VPWR_c_315_n 0.0230866f $X=3.032 $Y=2.215 $X2=0 $Y2=0
cc_201 A1 N_VPWR_c_315_n 0.0229619f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_202 N_A1_c_279_n N_VPWR_c_317_n 0.00386543f $X=3.032 $Y=2.215 $X2=0 $Y2=0
cc_203 N_A1_c_279_n N_VPWR_c_310_n 0.0076021f $X=3.032 $Y=2.215 $X2=0 $Y2=0
cc_204 N_A1_c_273_n N_A_339_47#_c_413_n 0.0142746f $X=3.002 $Y=0.84 $X2=0 $Y2=0
cc_205 N_A1_c_275_n N_A_339_47#_c_413_n 0.00701143f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_206 A1 N_A_339_47#_c_413_n 0.0152118f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_207 N_A1_c_277_n N_A_339_47#_c_413_n 4.87955e-19 $X=3.09 $Y=1.63 $X2=0 $Y2=0
cc_208 N_A1_c_272_n N_A_339_47#_c_415_n 0.00357871f $X=2.82 $Y=0.765 $X2=0 $Y2=0
cc_209 N_A1_c_273_n N_A_339_47#_c_415_n 0.00448539f $X=3.002 $Y=0.84 $X2=0 $Y2=0
cc_210 N_A1_c_272_n N_VGND_c_445_n 0.00320453f $X=2.82 $Y=0.765 $X2=0 $Y2=0
cc_211 N_A1_c_272_n N_VGND_c_447_n 0.00585385f $X=2.82 $Y=0.765 $X2=0 $Y2=0
cc_212 N_A1_c_273_n N_VGND_c_447_n 6.23557e-19 $X=3.002 $Y=0.84 $X2=0 $Y2=0
cc_213 N_A1_c_272_n N_VGND_c_448_n 0.00721851f $X=2.82 $Y=0.765 $X2=0 $Y2=0
cc_214 N_A1_c_273_n N_VGND_c_448_n 3.40618e-19 $X=3.002 $Y=0.84 $X2=0 $Y2=0
cc_215 N_VPWR_c_312_n N_Y_c_354_n 0.00306684f $X=0.29 $Y=2.47 $X2=0 $Y2=0
cc_216 N_VPWR_c_312_n N_Y_c_355_n 0.0184375f $X=0.29 $Y=2.47 $X2=0 $Y2=0
cc_217 N_VPWR_c_313_n N_Y_c_356_n 0.0263641f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_218 N_VPWR_c_315_n N_Y_c_356_n 3.05712e-19 $X=3.1 $Y=2.48 $X2=0 $Y2=0
cc_219 N_VPWR_c_317_n N_Y_c_356_n 0.0116754f $X=2.935 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_c_310_n N_Y_c_356_n 0.00944183f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_313_n N_Y_c_357_n 0.0676798f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_222 N_VPWR_c_312_n Y 0.0268142f $X=0.29 $Y=2.47 $X2=0 $Y2=0
cc_223 N_VPWR_c_313_n Y 0.0270363f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_224 N_VPWR_c_316_n Y 0.01394f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_225 N_VPWR_c_310_n Y 0.0112748f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_226 N_Y_c_352_n N_VGND_c_446_n 0.0128027f $X=0.365 $Y=0.437 $X2=0 $Y2=0
cc_227 N_Y_c_363_n N_VGND_c_446_n 0.026061f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_228 N_Y_M1006_s N_VGND_c_448_n 0.00503034f $X=0.22 $Y=0.235 $X2=0 $Y2=0
cc_229 N_Y_c_352_n N_VGND_c_448_n 0.00806516f $X=0.365 $Y=0.437 $X2=0 $Y2=0
cc_230 N_Y_c_363_n N_VGND_c_448_n 0.0181003f $X=0.685 $Y=0.445 $X2=0 $Y2=0
cc_231 A_195_47# N_VGND_c_448_n 0.00388585f $X=0.975 $Y=0.235 $X2=0 $Y2=0
cc_232 A_267_47# N_VGND_c_448_n 0.00773626f $X=1.335 $Y=0.235 $X2=3.12 $Y2=0
cc_233 N_A_339_47#_c_413_n N_VGND_c_445_n 0.0169862f $X=2.91 $Y=0.865 $X2=0
+ $Y2=0
cc_234 N_A_339_47#_c_416_n N_VGND_c_446_n 0.0203214f $X=2.035 $Y=0.437 $X2=0
+ $Y2=0
cc_235 N_A_339_47#_c_437_p N_VGND_c_446_n 0.0147885f $X=2.167 $Y=0.595 $X2=0
+ $Y2=0
cc_236 N_A_339_47#_c_415_n N_VGND_c_447_n 0.0162611f $X=3.035 $Y=0.445 $X2=0
+ $Y2=0
cc_237 N_A_339_47#_M1009_d N_VGND_c_448_n 0.00518123f $X=1.695 $Y=0.235 $X2=0
+ $Y2=0
cc_238 N_A_339_47#_M1004_d N_VGND_c_448_n 0.00224632f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_239 N_A_339_47#_c_416_n N_VGND_c_448_n 0.0142487f $X=2.035 $Y=0.437 $X2=0
+ $Y2=0
cc_240 N_A_339_47#_c_437_p N_VGND_c_448_n 0.0101731f $X=2.167 $Y=0.595 $X2=0
+ $Y2=0
cc_241 N_A_339_47#_c_413_n N_VGND_c_448_n 0.0110603f $X=2.91 $Y=0.865 $X2=0
+ $Y2=0
cc_242 N_A_339_47#_c_415_n N_VGND_c_448_n 0.0110561f $X=3.035 $Y=0.445 $X2=0
+ $Y2=0
