* File: sky130_fd_sc_lp__nand4bb_1.spice
* Created: Fri Aug 28 10:52:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4bb_1.pex.spice"
.subckt sky130_fd_sc_lp__nand4bb_1  VNB VPB B_N D C A_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A_N	A_N
* C	C
* D	D
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_B_N_M1006_g N_A_49_367#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.098 AS=0.1197 PD=0.85 PS=1.41 NRD=50.952 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 A_294_47# N_D_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.196 PD=1.05 PS=1.7 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.5 SB=75001.6 A=0.126
+ P=1.98 MULT=1
MM1003 A_366_47# N_C_M1003_g A_294_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75000.9 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1005 A_474_47# N_A_49_367#_M1005_g A_366_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=19.992 M=1 R=5.6 SA=75001.4
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1009_d N_A_552_21#_M1009_g A_474_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_552_21#_M1001_d N_A_N_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_B_N_M1007_g N_A_49_367#_M1007_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.12285 AS=0.1197 PD=0.95 PS=1.41 NRD=121.943 NRS=9.3772 M=1 R=2.8
+ SA=75000.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1011 N_Y_M1011_d N_D_M1011_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.36855 PD=1.54 PS=2.85 NRD=0 NRS=5.2008 M=1 R=8.4 SA=75000.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_C_M1004_g N_Y_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2709 AS=0.1764 PD=1.69 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1000_d N_A_49_367#_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2709 PD=1.54 PS=1.69 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75001.5
+ SB=75000.9 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_552_21#_M1008_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.37485 AS=0.1764 PD=2.715 PS=1.54 NRD=16.154 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.5 A=0.189 P=2.82 MULT=1
MM1010 N_A_552_21#_M1010_d N_A_N_M1010_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.12495 PD=1.37 PS=0.905 NRD=0 NRS=4.6886 M=1 R=2.8
+ SA=75003.1 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__nand4bb_1.pxi.spice"
*
.ends
*
*
