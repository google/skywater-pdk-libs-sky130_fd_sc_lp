* File: sky130_fd_sc_lp__a311oi_4.spice
* Created: Wed Sep  2 09:25:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311oi_4.pex.spice"
.subckt sky130_fd_sc_lp__a311oi_4  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A3_M1012_g N_A_27_47#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1012_d N_A3_M1022_g N_A_27_47#_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_A3_M1024_g N_A_27_47#_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1039 N_VGND_M1024_d N_A3_M1039_g N_A_27_47#_M1039_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1009 N_A_27_47#_M1039_s N_A2_M1009_g N_A_454_47#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1018 N_A_27_47#_M1018_d N_A2_M1018_g N_A_454_47#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1032 N_A_27_47#_M1018_d N_A2_M1032_g N_A_454_47#_M1032_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1033 N_A_27_47#_M1033_d N_A2_M1033_g N_A_454_47#_M1032_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g N_A_454_47#_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75005
+ A=0.126 P=1.98 MULT=1
MM1021 N_Y_M1021_d N_A1_M1021_g N_A_454_47#_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.6 A=0.126 P=1.98 MULT=1
MM1028 N_Y_M1021_d N_A1_M1028_g N_A_454_47#_M1028_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.2 A=0.126 P=1.98 MULT=1
MM1037 N_Y_M1037_d N_A1_M1037_g N_A_454_47#_M1028_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1218 AS=0.1176 PD=1.13 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_B1_M1001_g N_Y_M1037_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1218 PD=1.12 PS=1.13 NRD=0 NRS=1.428 M=1 R=5.6 SA=75001.9
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1001_d N_B1_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_B1_M1015_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.1176 PD=1.22 PS=1.12 NRD=6.42 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1015_d N_B1_M1019_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.1176 PD=1.22 PS=1.12 NRD=7.848 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1019_s N_C1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1016 N_Y_M1016_d N_C1_M1016_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1030 N_Y_M1016_d N_C1_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1031 N_Y_M1031_d N_C1_M1031_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A3_M1008_g N_A_124_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1023_d N_A3_M1023_g N_A_124_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.6 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1023_d N_A3_M1026_g N_A_124_367#_M1026_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.2 A=0.189 P=2.82 MULT=1
MM1034 N_VPWR_M1034_d N_A3_M1034_g N_A_124_367#_M1026_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1004 N_A_124_367#_M1004_d N_A2_M1004_g N_VPWR_M1034_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1014 N_A_124_367#_M1004_d N_A2_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1020 N_A_124_367#_M1020_d N_A2_M1020_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1035 N_A_124_367#_M1020_d N_A2_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2457 PD=1.54 PS=1.65 NRD=0 NRS=8.5892 M=1 R=8.4
+ SA=75003.2 SB=75002 A=0.189 P=2.82 MULT=1
MM1002 N_A_124_367#_M1002_d N_A1_M1002_g N_VPWR_M1035_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2457 PD=1.54 PS=1.65 NRD=0 NRS=8.5892 M=1 R=8.4
+ SA=75003.7 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_A_124_367#_M1002_d N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1010 N_A_124_367#_M1010_d N_A1_M1010_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_A_124_367#_M1010_d N_A1_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_A_124_367#_M1007_d N_B1_M1007_g N_A_1199_367#_M1007_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1025 N_A_124_367#_M1007_d N_B1_M1025_g N_A_1199_367#_M1025_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1029 N_A_124_367#_M1029_d N_B1_M1029_g N_A_1199_367#_M1025_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1036 N_A_124_367#_M1029_d N_B1_M1036_g N_A_1199_367#_M1036_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_A_1199_367#_M1036_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1003_d N_C1_M1011_g N_A_1199_367#_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1027 N_Y_M1027_d N_C1_M1027_g N_A_1199_367#_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1038 N_Y_M1027_d N_C1_M1038_g N_A_1199_367#_M1038_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.5079 P=24.65
*
.include "sky130_fd_sc_lp__a311oi_4.pxi.spice"
*
.ends
*
*
