# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__ebufn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.270000 3.415000 1.940000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.348000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 1.270000 2.780000 1.940000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.345000 0.730000 1.145000 ;
        RECT 0.125000 1.145000 0.355000 1.815000 ;
        RECT 0.125000 1.815000 0.700000 3.075000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.525000  1.315000 0.855000 1.455000 ;
      RECT 0.525000  1.455000 1.860000 1.625000 ;
      RECT 0.525000  1.625000 0.855000 1.645000 ;
      RECT 1.190000  1.795000 1.520000 3.245000 ;
      RECT 1.220000  0.085000 1.550000 1.225000 ;
      RECT 1.690000  1.625000 1.860000 2.905000 ;
      RECT 1.690000  2.905000 2.620000 3.075000 ;
      RECT 1.820000  0.255000 2.200000 0.585000 ;
      RECT 2.030000  0.585000 2.200000 0.640000 ;
      RECT 2.030000  0.640000 2.570000 1.100000 ;
      RECT 2.030000  1.100000 2.280000 2.735000 ;
      RECT 2.450000  2.110000 3.755000 2.280000 ;
      RECT 2.450000  2.280000 2.620000 2.905000 ;
      RECT 2.740000  0.085000 3.070000 1.100000 ;
      RECT 2.790000  2.450000 3.120000 3.245000 ;
      RECT 3.240000  0.640000 3.570000 0.930000 ;
      RECT 3.240000  0.930000 3.755000 1.100000 ;
      RECT 3.290000  2.280000 3.755000 2.790000 ;
      RECT 3.585000  1.100000 3.755000 2.110000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__ebufn_1
END LIBRARY
