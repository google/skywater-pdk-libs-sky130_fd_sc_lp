* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srsdfrtp_1 CLK D RESET_B SCD SCE SLEEP_B KAPWR VGND VNB VPB
+ VPWR Q
M1000 a_999_424# a_969_318# a_332_136# VPB phighvt w=420000u l=150000u
+  ad=4.252e+11p pd=3.81e+06u as=6.772e+11p ps=5.08e+06u
M1001 VPWR a_999_424# a_1176_349# VPB phighvt w=840000u l=150000u
+  ad=2.596e+12p pd=1.588e+07u as=4.788e+11p ps=4.5e+06u
M1002 VGND a_2176_99# a_2206_125# VNB nshort w=420000u l=150000u
+  ad=1.38275e+12p pd=1.474e+07u as=8.82e+10p ps=1.26e+06u
M1003 VGND SCE a_27_110# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1004 a_1128_424# a_1098_271# a_999_424# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1005 a_2836_390# a_969_318# a_1982_397# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=5.244e+11p ps=4.82e+06u
M1006 a_2472_119# a_1982_397# a_2176_99# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.155e+11p ps=1.39e+06u
M1007 a_2544_119# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1008 a_552_466# a_27_110# a_332_136# VPB phighvt w=640000u l=150000u
+  ad=2.304e+11p pd=2e+06u as=0p ps=0u
M1009 VPWR SCD a_552_466# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_534_136# a_27_110# a_462_136# VNB nshort w=420000u l=150000u
+  ad=2.331e+11p pd=2.79e+06u as=8.82e+10p ps=1.26e+06u
M1011 a_2206_125# a_2176_99# a_2134_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 a_3694_73# SLEEP_B a_2586_249# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.155e+11p ps=1.39e+06u
M1013 a_969_318# a_1098_271# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1014 VGND SLEEP_B a_3694_73# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 KAPWR a_1982_397# a_2176_99# VPB phighvt w=1e+06u l=250000u
+  ad=1.23675e+12p pd=8.71e+06u as=2.8e+11p ps=2.56e+06u
M1016 Q a_3751_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1017 a_313_466# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1018 a_2134_125# a_1098_271# a_1982_397# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.99e+11p ps=2.29e+06u
M1019 a_220_136# SCD a_534_136# VNB nshort w=420000u l=150000u
+  ad=2.877e+11p pd=3.05e+06u as=0p ps=0u
M1020 VPWR a_1176_349# a_1128_424# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_462_136# D a_332_136# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.64e+11p ps=3.51e+06u
M1022 KAPWR a_2176_99# a_2836_390# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_534_136# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1098_271# CLK KAPWR VPB phighvt w=640000u l=150000u
+  ad=1.984e+11p pd=1.9e+06u as=0p ps=0u
M1025 a_2586_249# SLEEP_B KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=4.232e+11p pd=2.96e+06u as=0p ps=0u
M1026 a_1982_397# a_969_318# a_1931_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1027 KAPWR SLEEP_B a_1098_271# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_3407_97# SLEEP_B a_3335_97# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1029 a_969_318# a_1098_271# VGND VNB nshort w=420000u l=150000u
+  ad=2.703e+11p pd=2.42e+06u as=0p ps=0u
M1030 VGND SLEEP_B a_3407_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_3751_367# a_1982_397# VGND VNB nshort w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
M1032 a_332_136# a_1098_271# a_999_424# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1033 a_999_424# a_969_318# a_929_152# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.248e+11p ps=3.27e+06u
M1034 VPWR SCE a_27_110# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1035 a_1931_125# a_969_318# a_1176_349# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.52e+11p ps=3.66e+06u
M1036 a_3063_390# a_2586_249# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1037 a_2069_397# a_1098_271# a_1982_397# VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1038 a_1176_349# a_1098_271# a_2069_397# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_332_136# D a_313_466# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_332_136# SCE a_220_136# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_2176_99# RESET_B a_3063_390# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND RESET_B a_1343_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1043 a_999_424# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_2544_119# a_1982_397# a_2472_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_332_136# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VGND a_999_424# a_1176_349# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_2586_249# a_2544_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_3335_97# CLK a_1098_271# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.68e+11p ps=1.64e+06u
M1049 Q a_3751_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.31e+11p pd=2.23e+06u as=0p ps=0u
M1050 a_1343_119# a_1176_349# a_929_152# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VPWR a_1982_397# a_3751_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
.ends
