* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and3b_m A_N B C VGND VNB VPB VPWR X
X0 a_220_53# a_110_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND A_N a_110_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_220_53# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_304_53# B a_376_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A_N a_110_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_376_53# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_220_53# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_220_53# a_110_53# a_304_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_220_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR B a_220_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
