* File: sky130_fd_sc_lp__ebufn_lp2.spice
* Created: Fri Aug 28 10:32:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ebufn_lp2.pex.spice"
.subckt sky130_fd_sc_lp__ebufn_lp2  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_114_47# N_A_M1001_g N_A_27_47#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g A_114_47# VNB NSHORT L=0.15 W=0.42 AD=0.1701
+ AS=0.0504 PD=1.65 PS=0.66 NRD=34.284 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1003 A_425_193# N_A_27_47#_M1003_g N_Z_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.08575 AS=0.1197 PD=0.945 PS=1.41 NRD=42.612 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_232_231#_M1008_g A_425_193# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.08575 PD=0.7 PS=0.945 NRD=0 NRS=42.612 M=1 R=2.8 SA=75000.4
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1006 A_606_153# N_TE_B_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_232_231#_M1002_d N_TE_B_M1002_g A_606_153# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1004 A_475_419# N_A_27_47#_M1004_g N_Z_M1004_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_TE_B_M1009_g A_475_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1005 N_A_232_231#_M1005_d N_TE_B_M1005_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.5154 P=12.69
*
.include "sky130_fd_sc_lp__ebufn_lp2.pxi.spice"
*
.ends
*
*
