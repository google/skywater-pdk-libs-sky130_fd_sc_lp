* File: sky130_fd_sc_lp__clkbuf_lp.pex.spice
* Created: Fri Aug 28 10:15:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUF_LP%A_94_31# 1 2 9 11 13 17 21 24 25 28 32 34
r55 32 34 53.9343 $w=2.48e-07 $l=1.17e-06 $layer=LI1_cond $X=2.1 $Y=1.665
+ $X2=2.1 $Y2=0.495
r56 28 30 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.7 $Y=2.18 $X2=1.7
+ $Y2=2.89
r57 26 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.7 $Y=1.75 $X2=2.1
+ $Y2=1.75
r58 26 28 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.7 $Y=1.835
+ $X2=1.7 $Y2=2.18
r59 24 26 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=1.75
+ $X2=1.7 $Y2=1.75
r60 24 25 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.535 $Y=1.75
+ $X2=1.07 $Y2=1.75
r61 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.905
+ $Y=1.33 $X2=0.905 $Y2=1.33
r62 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.905 $Y=1.665
+ $X2=1.07 $Y2=1.75
r63 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.905 $Y=1.665
+ $X2=0.905 $Y2=1.33
r64 15 22 31.1986 $w=2.74e-07 $l=2.22486e-07 $layer=POLY_cond $X=0.905 $Y=1.165
+ $X2=0.77 $Y2=1.33
r65 15 17 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.905 $Y=1.165
+ $X2=0.905 $Y2=0.495
r66 11 22 58.7894 $w=5.49e-07 $l=5.57293e-07 $layer=POLY_cond $X=0.66 $Y=1.835
+ $X2=0.77 $Y2=1.33
r67 11 13 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.66 $Y=1.835 $X2=0.66
+ $Y2=2.535
r68 7 22 31.1986 $w=2.74e-07 $l=2.96226e-07 $layer=POLY_cond $X=0.545 $Y=1.165
+ $X2=0.77 $Y2=1.33
r69 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.545 $Y=1.165
+ $X2=0.545 $Y2=0.495
r70 2 30 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=2.035 $X2=1.7 $Y2=2.89
r71 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=2.035 $X2=1.7 $Y2=2.18
r72 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.285 $X2=2.06 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_LP%A 1 3 5 7 8 10 11 12 13
r34 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=0.925
+ $X2=1.63 $Y2=1.295
r35 12 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=0.98 $X2=1.63 $Y2=0.98
r36 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=0.555
+ $X2=1.63 $Y2=0.925
r37 8 18 36.9986 $w=2.21e-07 $l=3.01413e-07 $layer=POLY_cond $X=1.845 $Y=0.815
+ $X2=1.615 $Y2=0.98
r38 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.845 $Y=0.815
+ $X2=1.845 $Y2=0.495
r39 5 18 36.9986 $w=2.21e-07 $l=2.20624e-07 $layer=POLY_cond $X=1.485 $Y=0.815
+ $X2=1.615 $Y2=0.98
r40 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.815
+ $X2=1.485 $Y2=0.495
r41 1 18 85.2364 $w=4.43e-07 $l=7.84857e-07 $layer=POLY_cond $X=1.435 $Y=1.68
+ $X2=1.615 $Y2=0.98
r42 1 3 212.428 $w=2.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.435 $Y=1.68
+ $X2=1.435 $Y2=2.535
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_LP%X 1 2 7 8 9 10 11 12 13 24 44
r19 34 44 0.45038 $w=4.33e-07 $l=1.7e-08 $layer=LI1_cond $X=0.342 $Y=2.052
+ $X2=0.342 $Y2=2.035
r20 13 48 3.60668 $w=3.89e-07 $l=1.15e-07 $layer=LI1_cond $X=0.342 $Y=2.775
+ $X2=0.342 $Y2=2.89
r21 13 35 3.02506 $w=4.35e-07 $l=1.02e-07 $layer=LI1_cond $X=0.342 $Y=2.775
+ $X2=0.342 $Y2=2.673
r22 12 35 7.10011 $w=4.33e-07 $l=2.68e-07 $layer=LI1_cond $X=0.342 $Y=2.405
+ $X2=0.342 $Y2=2.673
r23 12 38 5.96091 $w=4.33e-07 $l=2.25e-07 $layer=LI1_cond $X=0.342 $Y=2.405
+ $X2=0.342 $Y2=2.18
r24 11 44 0.90076 $w=4.33e-07 $l=3.4e-08 $layer=LI1_cond $X=0.342 $Y=2.001
+ $X2=0.342 $Y2=2.035
r25 11 42 4.68814 $w=4.33e-07 $l=1.66e-07 $layer=LI1_cond $X=0.342 $Y=2.001
+ $X2=0.342 $Y2=1.835
r26 11 38 2.49034 $w=4.33e-07 $l=9.4e-08 $layer=LI1_cond $X=0.342 $Y=2.086
+ $X2=0.342 $Y2=2.18
r27 11 34 0.90076 $w=4.33e-07 $l=3.4e-08 $layer=LI1_cond $X=0.342 $Y=2.086
+ $X2=0.342 $Y2=2.052
r28 10 42 5.29501 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.31 $Y=1.665
+ $X2=0.31 $Y2=1.835
r29 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.665
r30 8 9 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=0.925 $X2=0.31
+ $Y2=1.295
r31 7 8 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=0.555 $X2=0.31
+ $Y2=0.925
r32 7 24 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=0.31 $Y=0.555 $X2=0.31
+ $Y2=0.495
r33 2 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.25
+ $Y=2.035 $X2=0.395 $Y2=2.89
r34 2 38 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.25
+ $Y=2.035 $X2=0.395 $Y2=2.18
r35 1 24 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.285 $X2=0.33 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_LP%VPWR 1 6 11 12 13 23 24
r22 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r23 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r24 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 13 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 13 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 13 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r28 11 16 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=3.33 $X2=0.72
+ $Y2=3.33
r29 11 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=3.33
+ $X2=0.925 $Y2=3.33
r30 10 20 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 10 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.925 $Y2=3.33
r32 6 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.925 $Y=2.18 $X2=0.925
+ $Y2=2.89
r33 4 12 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=3.33
r34 4 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=2.89
r35 1 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.785
+ $Y=2.035 $X2=0.925 $Y2=2.89
r36 1 6 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.785
+ $Y=2.035 $X2=0.925 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_LP%VGND 1 6 8 10 17 18 21
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r28 15 17 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=2.16
+ $Y2=0
r29 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r31 10 12 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.72
+ $Y2=0
r32 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r33 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r34 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085 $X2=1.12
+ $Y2=0
r36 4 6 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.12 $Y=0.085 $X2=1.12
+ $Y2=0.495
r37 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.285 $X2=1.12 $Y2=0.495
.ends

