* File: sky130_fd_sc_lp__dfrtn_1.spice
* Created: Wed Sep  2 09:43:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfrtn_1.pex.spice"
.subckt sky130_fd_sc_lp__dfrtn_1  VNB VPB D RESET_B CLK_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK_N	CLK_N
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1023 A_142_121# N_RESET_B_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1020 N_A_27_463#_M1020_d N_D_M1020_g A_142_121# VNB NSHORT L=0.15 W=0.42
+ AD=0.1118 AS=0.0441 PD=0.96 PS=0.63 NRD=30 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1001 N_A_336_463#_M1001_d N_A_294_35#_M1001_g N_A_27_463#_M1020_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0609 AS=0.1118 PD=0.71 PS=0.96 NRD=0 NRS=41.424 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1011 A_438_123# N_A_306_277#_M1011_g N_A_336_463#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0609 PD=0.78 PS=0.71 NRD=35.712 NRS=2.856 M=1 R=2.8
+ SA=75001.6 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1006 A_540_123# N_A_501_229#_M1006_g A_438_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.07245 AS=0.0756 PD=0.765 PS=0.78 NRD=33.564 NRS=35.712 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_RESET_B_M1031_g A_540_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.23595 AS=0.07245 PD=2.14 PS=0.765 NRD=144.792 NRS=33.564 M=1 R=2.8
+ SA=75002.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_306_277#_M1016_g N_A_294_35#_M1016_s VNB NSHORT L=0.15
+ W=0.42 AD=0.148308 AS=0.126 PD=1.05396 PS=1.44 NRD=85.164 NRS=4.284 M=1 R=2.8
+ SA=75000.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1028 N_A_501_229#_M1028_d N_A_336_463#_M1028_g N_VGND_M1016_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1408 AS=0.225992 PD=1.08 PS=1.60604 NRD=29.988 NRS=32.808
+ M=1 R=4.26667 SA=75000.7 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1007 N_A_1099_447#_M1007_d N_A_306_277#_M1007_g N_A_501_229#_M1028_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.176423 AS=0.1408 PD=1.52151 PS=1.08 NRD=48.744 NRS=0
+ M=1 R=4.26667 SA=75001.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 A_1275_125# N_A_294_35#_M1018_g N_A_1099_447#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.115777 PD=0.63 PS=0.998491 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1287_276#_M1013_g A_1275_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.111975 AS=0.0441 PD=0.995 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8
+ SA=75002.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1019 A_1465_125# N_RESET_B_M1019_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.111975 PD=0.63 PS=0.995 NRD=14.28 NRS=24.276 M=1 R=2.8
+ SA=75002.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_1287_276#_M1014_d N_A_1099_447#_M1014_g A_1465_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_CLK_N_M1025_g N_A_306_277#_M1025_s VNB NSHORT L=0.15
+ W=0.42 AD=0.204125 AS=0.1113 PD=1.95 PS=1.37 NRD=82.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_1099_447#_M1026_g N_A_1832_367#_M1026_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1010 N_Q_M1010_d N_A_1832_367#_M1010_g N_VGND_M1026_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=2.496 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1029 N_VPWR_M1029_d N_RESET_B_M1029_g N_A_27_463#_M1029_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.135 AS=0.1113 PD=1.085 PS=1.37 NRD=56.2829 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1004 N_A_27_463#_M1004_d N_D_M1004_g N_VPWR_M1029_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.135 PD=0.74 PS=1.085 NRD=0 NRS=56.2829 M=1 R=2.8 SA=75000.8
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1030 N_A_336_463#_M1030_d N_A_306_277#_M1030_g N_A_27_463#_M1004_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.08505 AS=0.0672 PD=0.825 PS=0.74 NRD=37.5088 NRS=18.7544
+ M=1 R=2.8 SA=75001.3 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 A_447_463# N_A_294_35#_M1002_g N_A_336_463#_M1030_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.08505 PD=0.81 PS=0.825 NRD=65.6601 NRS=21.0987 M=1 R=2.8
+ SA=75001.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_501_229#_M1015_g A_447_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.111975 AS=0.0819 PD=0.995 PS=0.81 NRD=39.8531 NRS=65.6601 M=1 R=2.8
+ SA=75002.4 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1022 N_A_336_463#_M1022_d N_RESET_B_M1022_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.111975 PD=1.37 PS=0.995 NRD=0 NRS=39.8531 M=1 R=2.8
+ SA=75003 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_306_277#_M1008_g N_A_294_35#_M1008_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.22907 AS=0.23925 PD=1.52649 PS=2.18 NRD=93.2401 NRS=19.9955
+ M=1 R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1017 N_A_501_229#_M1017_d N_A_336_463#_M1017_g N_VPWR_M1008_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.300655 PD=1.12 PS=2.00351 NRD=0 NRS=21.0987 M=1
+ R=5.6 SA=75000.6 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1003 N_A_1099_447#_M1003_d N_A_294_35#_M1003_g N_A_501_229#_M1017_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2142 AS=0.1176 PD=1.78667 PS=1.12 NRD=0 NRS=0 M=1
+ R=5.6 SA=75001 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1005 A_1229_531# N_A_306_277#_M1005_g N_A_1099_447#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.1071 PD=0.81 PS=0.893333 NRD=65.6601 NRS=93.7917 M=1
+ R=2.8 SA=75001.4 SB=75002 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_A_1287_276#_M1027_g A_1229_531# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0945 AS=0.0819 PD=0.87 PS=0.81 NRD=0 NRS=65.6601 M=1 R=2.8
+ SA=75001.9 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_1287_276#_M1000_d N_RESET_B_M1000_g N_VPWR_M1027_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.14045 AS=0.0945 PD=1.16 PS=0.87 NRD=131.044 NRS=79.7259 M=1 R=2.8
+ SA=75002.5 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_1099_447#_M1021_g N_A_1287_276#_M1000_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0954906 AS=0.14045 PD=0.851887 PS=1.16 NRD=80.8291
+ NRS=11.7215 M=1 R=2.8 SA=75001.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_306_277#_M1009_d N_CLK_N_M1009_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.145509 PD=1.81 PS=1.29811 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_VPWR_M1024_d N_A_1099_447#_M1024_g N_A_1832_367#_M1024_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.14912 AS=0.1696 PD=1.14189 PS=1.81 NRD=33.0763 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 N_Q_M1012_d N_A_1832_367#_M1012_g N_VPWR_M1024_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.29358 PD=3.05 PS=2.24811 NRD=0 NRS=5.2008 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.4031 P=25.61
c_130 VNB 0 1.4009e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfrtn_1.pxi.spice"
*
.ends
*
*
