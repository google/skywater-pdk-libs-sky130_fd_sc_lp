* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VGND a_90_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VPWR B1 a_90_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR a_90_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR A1 a_792_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_792_367# A2 a_90_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A1 a_485_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_90_23# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VPWR a_90_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_792_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X a_90_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 X a_90_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_90_23# A2 a_792_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND a_90_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_485_65# B1 a_90_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_90_23# B1 a_485_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_485_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 X a_90_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VGND A2 a_485_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_485_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 X a_90_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
