# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__maj3_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__maj3_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.605000 1.795000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.225000 1.315000 1.245000 ;
        RECT 0.440000 1.245000 2.750000 1.415000 ;
        RECT 0.440000 1.415000 0.760000 1.895000 ;
        RECT 1.085000 1.180000 1.315000 1.225000 ;
        RECT 2.420000 1.415000 2.750000 1.915000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.960000 1.245000 3.290000 1.915000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.755000 1.920000 4.210000 3.065000 ;
        RECT 3.875000 0.320000 4.210000 0.780000 ;
        RECT 4.040000 0.780000 4.210000 1.920000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.090000  0.875000 1.665000 0.895000 ;
      RECT 0.090000  0.895000 3.695000 0.985000 ;
      RECT 0.090000  0.985000 3.860000 1.000000 ;
      RECT 0.090000  1.000000 0.645000 1.045000 ;
      RECT 0.090000  1.045000 0.260000 2.075000 ;
      RECT 0.090000  2.075000 0.455000 2.330000 ;
      RECT 0.090000  2.330000 2.515000 2.500000 ;
      RECT 0.090000  2.500000 0.455000 3.065000 ;
      RECT 0.315000  0.605000 0.645000 0.830000 ;
      RECT 0.315000  0.830000 1.665000 0.875000 ;
      RECT 1.195000  2.680000 1.525000 3.245000 ;
      RECT 1.215000  0.085000 1.545000 0.650000 ;
      RECT 1.495000  1.000000 3.860000 1.065000 ;
      RECT 2.185000  2.095000 2.515000 2.330000 ;
      RECT 2.185000  2.500000 2.515000 3.065000 ;
      RECT 2.195000  0.320000 2.525000 0.895000 ;
      RECT 3.085000  0.085000 3.415000 0.715000 ;
      RECT 3.215000  2.095000 3.545000 3.245000 ;
      RECT 3.525000  1.065000 3.860000 1.655000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__maj3_lp
END LIBRARY
