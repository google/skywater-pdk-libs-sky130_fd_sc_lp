* File: sky130_fd_sc_lp__xnor3_lp.pex.spice
* Created: Wed Sep  2 10:40:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A 3 7 11 13 19
c40 11 0 1.49436e-20 $X=0.855 $Y=0.755
c41 7 0 2.7607e-19 $X=0.67 $Y=2.545
r42 17 19 6.83688 $w=2.82e-07 $l=4e-08 $layer=POLY_cond $X=0.63 $Y=1.68 $X2=0.67
+ $Y2=1.68
r43 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.68 $X2=0.63 $Y2=1.68
r44 15 17 23.0745 $w=2.82e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=1.68
+ $X2=0.63 $Y2=1.68
r45 13 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.68 $X2=0.63
+ $Y2=1.68
r46 9 19 31.6206 $w=2.82e-07 $l=2.5446e-07 $layer=POLY_cond $X=0.855 $Y=1.515
+ $X2=0.67 $Y2=1.68
r47 9 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.855 $Y=1.515
+ $X2=0.855 $Y2=0.755
r48 5 19 5.69241 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=1.845
+ $X2=0.67 $Y2=1.68
r49 5 7 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.67 $Y=1.845 $X2=0.67
+ $Y2=2.545
r50 1 15 17.5183 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.495 $Y2=1.68
r51 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.495 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A_27_109# 1 2 3 4 13 15 18 22 26 32 34 39
+ 40 41 43 44 45 47 48 49 51 52 53 54 58 62 64 65 67 69
c156 58 0 1.77657e-19 $X=5.96 $Y=0.805
c157 54 0 1.56206e-19 $X=5.795 $Y=0.7
c158 52 0 8.58584e-20 $X=4.425 $Y=0.98
c159 41 0 1.49436e-20 $X=1.505 $Y=0.35
r160 69 71 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.51 $Y=0.7
+ $X2=4.51 $Y2=0.98
r161 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.34
+ $Y=1.33 $X2=1.34 $Y2=1.33
r162 64 65 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.342 $Y=2.19
+ $X2=0.342 $Y2=2.025
r163 58 60 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=5.96 $Y=0.805
+ $X2=5.96 $Y2=1.88
r164 56 58 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=5.96 $Y=0.785
+ $X2=5.96 $Y2=0.805
r165 55 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=0.7
+ $X2=4.51 $Y2=0.7
r166 54 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.795 $Y=0.7
+ $X2=5.96 $Y2=0.785
r167 54 55 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=5.795 $Y=0.7
+ $X2=4.595 $Y2=0.7
r168 52 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=0.98
+ $X2=4.51 $Y2=0.98
r169 52 53 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.425 $Y=0.98
+ $X2=3.895 $Y2=0.98
r170 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=0.895
+ $X2=3.895 $Y2=0.98
r171 50 51 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.81 $Y=0.435
+ $X2=3.81 $Y2=0.895
r172 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=0.35
+ $X2=3.81 $Y2=0.435
r173 48 49 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.725 $Y=0.35
+ $X2=3.075 $Y2=0.35
r174 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.435
+ $X2=3.075 $Y2=0.35
r175 46 47 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.99 $Y=0.435
+ $X2=2.99 $Y2=0.995
r176 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=1.08
+ $X2=2.99 $Y2=0.995
r177 44 45 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.905 $Y=1.08
+ $X2=2.295 $Y2=1.08
r178 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.21 $Y=0.995
+ $X2=2.295 $Y2=1.08
r179 42 43 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.21 $Y=0.435
+ $X2=2.21 $Y2=0.995
r180 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.125 $Y=0.35
+ $X2=2.21 $Y2=0.435
r181 40 41 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.125 $Y=0.35
+ $X2=1.505 $Y2=0.35
r182 39 67 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.42 $Y=1.165
+ $X2=1.34 $Y2=1.25
r183 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.42 $Y=0.435
+ $X2=1.505 $Y2=0.35
r184 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.42 $Y=0.435
+ $X2=1.42 $Y2=1.165
r185 35 62 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.25
+ $X2=0.28 $Y2=1.25
r186 34 67 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=1.25
+ $X2=1.34 $Y2=1.25
r187 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.175 $Y=1.25
+ $X2=0.445 $Y2=1.25
r188 30 64 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=0.342 $Y=2.252
+ $X2=0.342 $Y2=2.19
r189 30 32 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=0.342 $Y=2.252
+ $X2=0.342 $Y2=2.9
r190 28 62 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=1.335
+ $X2=0.28 $Y2=1.25
r191 28 65 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.2 $Y=1.335 $X2=0.2
+ $Y2=2.025
r192 24 62 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=1.165
+ $X2=0.28 $Y2=1.25
r193 24 26 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=1.165
+ $X2=0.28 $Y2=0.755
r194 20 68 35.1394 $w=2.35e-07 $l=3.20038e-07 $layer=POLY_cond $X=1.645 $Y=1.165
+ $X2=1.397 $Y2=1.33
r195 20 22 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.645 $Y=1.165
+ $X2=1.645 $Y2=0.755
r196 16 68 35.1394 $w=2.35e-07 $l=2.13787e-07 $layer=POLY_cond $X=1.285 $Y=1.165
+ $X2=1.397 $Y2=1.33
r197 16 18 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.285 $Y=1.165
+ $X2=1.285 $Y2=0.755
r198 13 68 82.2877 $w=4.7e-07 $l=7.92401e-07 $layer=POLY_cond $X=1.2 $Y=2.03
+ $X2=1.397 $Y2=1.33
r199 13 15 99.292 $w=2.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.2 $Y=2.03 $X2=1.2
+ $Y2=2.545
r200 4 60 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.735 $X2=5.96 $Y2=1.88
r201 3 64 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=2.045 $X2=0.405 $Y2=2.19
r202 3 32 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=2.045 $X2=0.405 $Y2=2.9
r203 2 58 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=5.82
+ $Y=0.555 $X2=5.96 $Y2=0.805
r204 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.545 $X2=0.28 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A_647_367# 1 2 9 10 11 15 17 21 23 25 30 31
+ 35 40 41 47 48 51
c104 51 0 1.01058e-19 $X=3.665 $Y=1.245
c105 48 0 1.58999e-19 $X=3.665 $Y=1.41
c106 31 0 8.58584e-20 $X=4.305 $Y=1.5
c107 23 0 1.56206e-19 $X=5.695 $Y=1.395
r108 48 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.665 $Y=1.41
+ $X2=3.665 $Y2=1.5
r109 48 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.41
+ $X2=3.665 $Y2=1.245
r110 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.665
+ $Y=1.41 $X2=3.665 $Y2=1.41
r111 45 47 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.42 $Y=1.41
+ $X2=3.665 $Y2=1.41
r112 43 45 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=3.417 $Y=1.41
+ $X2=3.42 $Y2=1.41
r113 40 41 6.55101 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=1.98
+ $X2=3.375 $Y2=1.815
r114 37 43 2.50173 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=3.417 $Y=1.575
+ $X2=3.417 $Y2=1.41
r115 37 41 11.2892 $w=2.43e-07 $l=2.4e-07 $layer=LI1_cond $X=3.417 $Y=1.575
+ $X2=3.417 $Y2=1.815
r116 33 45 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=1.245
+ $X2=3.42 $Y2=1.41
r117 33 35 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=3.42 $Y=1.245
+ $X2=3.42 $Y2=0.78
r118 30 32 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.745 $Y=0.765
+ $X2=5.745 $Y2=1.27
r119 27 30 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.745 $Y=0.33
+ $X2=5.745 $Y2=0.765
r120 23 32 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=5.695 $Y=1.395
+ $X2=5.695 $Y2=1.27
r121 23 25 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.695 $Y=1.395
+ $X2=5.695 $Y2=2.235
r122 19 21 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.725 $Y=1.425
+ $X2=4.725 $Y2=0.985
r123 18 31 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.43 $Y=1.5
+ $X2=4.305 $Y2=1.5
r124 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.65 $Y=1.5
+ $X2=4.725 $Y2=1.425
r125 17 18 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.65 $Y=1.5
+ $X2=4.43 $Y2=1.5
r126 13 31 1.63566 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=1.575
+ $X2=4.305 $Y2=1.5
r127 13 15 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.305 $Y=1.575
+ $X2=4.305 $Y2=2.235
r128 12 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.5
+ $X2=3.665 $Y2=1.5
r129 11 31 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.18 $Y=1.5
+ $X2=4.305 $Y2=1.5
r130 11 12 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.18 $Y=1.5
+ $X2=3.83 $Y2=1.5
r131 9 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.67 $Y=0.255
+ $X2=5.745 $Y2=0.33
r132 9 10 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=5.67 $Y=0.255
+ $X2=3.83 $Y2=0.255
r133 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.755 $Y=0.33
+ $X2=3.83 $Y2=0.255
r134 7 51 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.755 $Y=0.33
+ $X2=3.755 $Y2=1.245
r135 2 40 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.235
+ $Y=1.835 $X2=3.375 $Y2=1.98
r136 1 35 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.505 $X2=3.46 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%B 3 8 11 13 14 18 20 23 25 29 31 34 36 37
+ 38 40 41 48 50
c121 48 0 1.58999e-19 $X=2.865 $Y=1.51
c122 34 0 4.30949e-20 $X=6.225 $Y=2.235
c123 31 0 1.27293e-19 $X=6.225 $Y=1.635
c124 29 0 7.10868e-21 $X=6.175 $Y=0.765
c125 18 0 1.77657e-19 $X=5.165 $Y=2.235
c126 11 0 1.75594e-19 $X=3.165 $Y=0.715
r127 49 50 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.11 $Y=1.51
+ $X2=3.165 $Y2=1.51
r128 47 49 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.865 $Y=1.51
+ $X2=3.11 $Y2=1.51
r129 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.51 $X2=2.865 $Y2=1.51
r130 44 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.775 $Y=1.51
+ $X2=2.865 $Y2=1.51
r131 41 48 5.96091 $w=4.33e-07 $l=2.25e-07 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=2.865 $Y2=1.562
r132 40 41 12.7166 $w=4.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=2.64 $Y2=1.562
r133 35 36 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.175 $Y=1.51
+ $X2=5.175 $Y2=1.66
r134 32 34 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.225 $Y=3.075
+ $X2=6.225 $Y2=2.235
r135 31 39 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.225 $Y=1.635
+ $X2=6.225 $Y2=1.51
r136 31 34 149.072 $w=2.5e-07 $l=6e-07 $layer=POLY_cond $X=6.225 $Y=1.635
+ $X2=6.225 $Y2=2.235
r137 29 39 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=6.175 $Y=0.765
+ $X2=6.175 $Y2=1.51
r138 26 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.19 $Y=3.15
+ $X2=5.115 $Y2=3.15
r139 25 32 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=6.1 $Y=3.15
+ $X2=6.225 $Y2=3.075
r140 25 26 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=6.1 $Y=3.15
+ $X2=5.19 $Y2=3.15
r141 23 35 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.235 $Y=0.985
+ $X2=5.235 $Y2=1.51
r142 20 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.115 $Y=3.075
+ $X2=5.115 $Y2=3.15
r143 20 37 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.115 $Y=3.075
+ $X2=5.115 $Y2=2.865
r144 18 36 142.861 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.165 $Y=2.235
+ $X2=5.165 $Y2=1.66
r145 16 37 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=5.165 $Y=2.74
+ $X2=5.165 $Y2=2.865
r146 16 18 125.469 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.165 $Y=2.74
+ $X2=5.165 $Y2=2.235
r147 13 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.04 $Y=3.15
+ $X2=5.115 $Y2=3.15
r148 13 14 925.543 $w=1.5e-07 $l=1.805e-06 $layer=POLY_cond $X=5.04 $Y=3.15
+ $X2=3.235 $Y2=3.15
r149 9 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.345
+ $X2=3.165 $Y2=1.51
r150 9 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.165 $Y=1.345
+ $X2=3.165 $Y2=0.715
r151 6 14 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.11 $Y=3.075
+ $X2=3.235 $Y2=3.15
r152 6 8 183.856 $w=2.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.11 $Y=3.075
+ $X2=3.11 $Y2=2.335
r153 5 49 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.675
+ $X2=3.11 $Y2=1.51
r154 5 8 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.675
+ $X2=3.11 $Y2=2.335
r155 1 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.345
+ $X2=2.775 $Y2=1.51
r156 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.775 $Y=1.345
+ $X2=2.775 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A_1318_85# 1 2 9 14 15 16 18 20 21 27 32 35
c89 35 0 6.27877e-20 $X=8.215 $Y=1.68
c90 14 0 1.07536e-19 $X=6.835 $Y=2.165
c91 9 0 2.18243e-19 $X=6.665 $Y=0.765
r92 35 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.215 $Y=1.68
+ $X2=8.215 $Y2=1.845
r93 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.215
+ $Y=1.68 $X2=8.215 $Y2=1.68
r94 31 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=8.56 $Y=0.795
+ $X2=8.56 $Y2=1.56
r95 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.48 $Y=2.15 $X2=8.48
+ $Y2=2.86
r96 25 32 3.92321 $w=2.33e-07 $l=8e-08 $layer=LI1_cond $X=8.48 $Y=1.677 $X2=8.56
+ $Y2=1.677
r97 25 34 12.9956 $w=2.33e-07 $l=2.65e-07 $layer=LI1_cond $X=8.48 $Y=1.677
+ $X2=8.215 $Y2=1.677
r98 25 27 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=8.48 $Y=1.795
+ $X2=8.48 $Y2=2.15
r99 21 31 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=8.475 $Y=0.705
+ $X2=8.56 $Y2=0.795
r100 21 23 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=8.475 $Y=0.705
+ $X2=7.88 $Y2=0.705
r101 19 20 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.775 $Y=1.44
+ $X2=6.775 $Y2=1.59
r102 18 42 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=8.125 $Y=3.035
+ $X2=8.125 $Y2=1.845
r103 15 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.05 $Y=3.11
+ $X2=8.125 $Y2=3.035
r104 15 16 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=8.05 $Y=3.11
+ $X2=6.96 $Y2=3.11
r105 14 20 142.861 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.835 $Y=2.165
+ $X2=6.835 $Y2=1.59
r106 12 16 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=6.835 $Y=3.035
+ $X2=6.96 $Y2=3.11
r107 12 14 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.835 $Y=3.035
+ $X2=6.835 $Y2=2.165
r108 9 19 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=6.665 $Y=0.765
+ $X2=6.665 $Y2=1.44
r109 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=2.005 $X2=8.48 $Y2=2.86
r110 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=2.005 $X2=8.48 $Y2=2.15
r111 1 23 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=7.735
+ $Y=0.445 $X2=7.88 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%C 1 3 6 9 10 12 13 15 17 20 25 26 30 31 33
c75 33 0 1.94241e-19 $X=8.17 $Y=1.14
c76 30 0 6.27877e-20 $X=7.895 $Y=1.14
c77 25 0 1.92026e-19 $X=8.682 $Y=1.23
c78 20 0 3.34909e-19 $X=8.745 $Y=2.505
c79 15 0 1.26986e-19 $X=8.57 $Y=1.155
c80 6 0 1.56469e-19 $X=7.365 $Y=2.165
r81 32 33 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.095 $Y=1.14
+ $X2=8.17 $Y2=1.14
r82 29 32 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.895 $Y=1.14
+ $X2=8.095 $Y2=1.14
r83 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.895 $Y=1.14
+ $X2=7.73 $Y2=1.14
r84 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.895
+ $Y=1.14 $X2=7.895 $Y2=1.14
r85 26 30 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.895 $Y=1.295
+ $X2=7.895 $Y2=1.14
r86 18 25 15.9654 $w=2e-07 $l=1.01735e-07 $layer=POLY_cond $X=8.745 $Y=1.305
+ $X2=8.682 $Y2=1.23
r87 18 20 298.144 $w=2.5e-07 $l=1.2e-06 $layer=POLY_cond $X=8.745 $Y=1.305
+ $X2=8.745 $Y2=2.505
r88 15 25 15.9654 $w=2e-07 $l=1.4472e-07 $layer=POLY_cond $X=8.57 $Y=1.155
+ $X2=8.682 $Y2=1.23
r89 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.57 $Y=1.155
+ $X2=8.57 $Y2=0.87
r90 13 25 9.46703 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=8.495 $Y=1.23
+ $X2=8.682 $Y2=1.23
r91 13 33 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=8.495 $Y=1.23
+ $X2=8.17 $Y2=1.23
r92 10 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=0.975
+ $X2=8.095 $Y2=1.14
r93 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.095 $Y=0.975
+ $X2=8.095 $Y2=0.655
r94 9 31 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.49 $Y=1.125
+ $X2=7.73 $Y2=1.125
r95 4 9 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.365 $Y=1.125
+ $X2=7.49 $Y2=1.125
r96 4 22 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.365 $Y=1.125
+ $X2=7.095 $Y2=1.125
r97 4 6 239.758 $w=2.5e-07 $l=9.65e-07 $layer=POLY_cond $X=7.365 $Y=1.2
+ $X2=7.365 $Y2=2.165
r98 1 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.095 $Y=1.05
+ $X2=7.095 $Y2=1.125
r99 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.095 $Y=1.05 $X2=7.095
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A_1348_111# 1 2 10 11 13 15 17 19 24 26 30
+ 33 35 40
c82 40 0 1.92026e-19 $X=9.3 $Y=0.385
c83 33 0 1.26986e-19 $X=9.02 $Y=0.385
c84 30 0 1.56469e-19 $X=7.1 $Y=1.81
c85 26 0 7.10868e-21 $X=6.965 $Y=0.35
c86 24 0 1.27293e-19 $X=6.88 $Y=0.765
c87 15 0 1.1992e-19 $X=9.51 $Y=0.475
r88 39 40 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.225 $Y=0.385
+ $X2=9.3 $Y2=0.385
r89 34 39 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=9.02 $Y=0.385
+ $X2=9.225 $Y2=0.385
r90 33 35 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=9.02 $Y=0.407
+ $X2=8.855 $Y2=0.407
r91 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.02
+ $Y=0.385 $X2=9.02 $Y2=0.385
r92 27 30 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=6.84 $Y=1.81 $X2=7.1
+ $Y2=1.81
r93 26 35 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=6.965 $Y=0.35
+ $X2=8.855 $Y2=0.35
r94 22 27 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=6.84 $Y=1.645
+ $X2=6.84 $Y2=1.81
r95 22 24 40.566 $w=2.48e-07 $l=8.8e-07 $layer=LI1_cond $X=6.84 $Y=1.645
+ $X2=6.84 $Y2=0.765
r96 21 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.84 $Y=0.435
+ $X2=6.965 $Y2=0.35
r97 21 24 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=6.84 $Y=0.435
+ $X2=6.84 $Y2=0.765
r98 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.585 $Y=0.55
+ $X2=9.585 $Y2=0.87
r99 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.51 $Y=0.475
+ $X2=9.585 $Y2=0.55
r100 15 40 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.51 $Y=0.475
+ $X2=9.3 $Y2=0.475
r101 11 20 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=9.275 $Y=1.575
+ $X2=9.275 $Y2=1.45
r102 11 13 231.062 $w=2.5e-07 $l=9.3e-07 $layer=POLY_cond $X=9.275 $Y=1.575
+ $X2=9.275 $Y2=2.505
r103 10 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.225 $Y=0.87
+ $X2=9.225 $Y2=1.45
r104 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.225 $Y=0.55
+ $X2=9.225 $Y2=0.385
r105 7 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.225 $Y=0.55
+ $X2=9.225 $Y2=0.87
r106 2 30 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.96
+ $Y=1.665 $X2=7.1 $Y2=1.81
r107 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.74
+ $Y=0.555 $X2=6.88 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%VPWR 1 2 3 12 18 22 27 28 29 35 39 46 47 50
+ 53
r65 53 54 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r66 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 47 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r68 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r69 44 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=3.33
+ $X2=9.01 $Y2=3.33
r70 44 46 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=9.175 $Y=3.33
+ $X2=9.84 $Y2=3.33
r71 43 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 42 43 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 40 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=2.765 $Y2=3.33
r74 40 42 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 39 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=9.01 $Y2=3.33
r76 39 42 373.503 $w=1.68e-07 $l=5.725e-06 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=3.12 $Y2=3.33
r77 38 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r79 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=3.33
+ $X2=2.765 $Y2=3.33
r80 35 37 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.6 $Y=3.33 $X2=1.2
+ $Y2=3.33
r81 33 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r82 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 29 54 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=8.88 $Y2=3.33
r84 29 43 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 27 32 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=3.33 $X2=0.72
+ $Y2=3.33
r86 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=3.33
+ $X2=0.935 $Y2=3.33
r87 26 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r88 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=0.935 $Y2=3.33
r89 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.01 $Y=2.15 $X2=9.01
+ $Y2=2.86
r90 20 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=3.245
+ $X2=9.01 $Y2=3.33
r91 20 25 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.01 $Y=3.245
+ $X2=9.01 $Y2=2.86
r92 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=3.245
+ $X2=2.765 $Y2=3.33
r93 16 18 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.765 $Y=3.245
+ $X2=2.765 $Y2=2.76
r94 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.935 $Y=2.19
+ $X2=0.935 $Y2=2.9
r95 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=3.33
r96 10 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=2.9
r97 3 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.87
+ $Y=2.005 $X2=9.01 $Y2=2.86
r98 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.87
+ $Y=2.005 $X2=9.01 $Y2=2.15
r99 2 18 600 $w=1.7e-07 $l=9.94862e-07 $layer=licon1_PDIFF $count=1 $X=2.62
+ $Y=1.835 $X2=2.765 $Y2=2.76
r100 1 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.795
+ $Y=2.045 $X2=0.935 $Y2=2.9
r101 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.795
+ $Y=2.045 $X2=0.935 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A_265_409# 1 2 3 4 15 18 19 21 24 29 31
c67 29 0 1.0345e-19 $X=1.865 $Y=2.22
c68 24 0 1.41873e-19 $X=4.57 $Y=1.88
c69 15 0 1.7262e-19 $X=1.465 $Y=2.9
r70 31 33 9.71523 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=1.82 $Y=0.8
+ $X2=1.82 $Y2=0.985
r71 28 29 6.24364 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=2.22
+ $X2=1.865 $Y2=2.22
r72 26 28 9.30819 $w=3.88e-07 $l=3.15e-07 $layer=LI1_cond $X=1.465 $Y=2.22
+ $X2=1.78 $Y2=2.22
r73 22 24 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.57 $Y=2.245
+ $X2=4.57 $Y2=1.88
r74 21 36 14.947 $w=3.02e-07 $l=5.01597e-07 $layer=LI1_cond $X=4.57 $Y=1.415
+ $X2=4.94 $Y2=1.105
r75 21 24 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.57 $Y=1.415
+ $X2=4.57 $Y2=1.88
r76 19 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.405 $Y=2.33
+ $X2=4.57 $Y2=2.245
r77 19 29 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=4.405 $Y=2.33
+ $X2=1.865 $Y2=2.33
r78 18 28 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.78 $Y=2.025
+ $X2=1.78 $Y2=2.22
r79 18 33 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.78 $Y=2.025
+ $X2=1.78 $Y2=0.985
r80 13 26 1.7167 $w=3.3e-07 $l=1.95e-07 $layer=LI1_cond $X=1.465 $Y=2.415
+ $X2=1.465 $Y2=2.22
r81 13 15 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.465 $Y=2.415
+ $X2=1.465 $Y2=2.9
r82 4 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.735 $X2=4.57 $Y2=1.88
r83 3 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=2.045 $X2=1.465 $Y2=2.19
r84 3 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=2.045 $X2=1.465 $Y2=2.9
r85 2 36 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.8
+ $Y=0.775 $X2=4.94 $Y2=1.05
r86 1 31 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.545 $X2=1.86 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A_763_347# 1 2 3 4 13 16 17 18 19 23 27 29
+ 32 33 34 36 38 42 43 47
c133 47 0 3.21756e-19 $X=7.45 $Y=0.805
c134 33 0 5.97696e-20 $X=7.895 $Y=2.06
c135 32 0 1.07536e-19 $X=7.45 $Y=1.975
r136 45 47 4.24584 $w=3.78e-07 $l=1.4e-07 $layer=LI1_cond $X=7.31 $Y=0.805
+ $X2=7.45 $Y2=0.805
r137 38 40 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.96 $Y=2.68 $X2=3.96
+ $Y2=2.98
r138 35 36 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.98 $Y=2.145
+ $X2=7.98 $Y2=2.895
r139 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.895 $Y=2.06
+ $X2=7.98 $Y2=2.145
r140 33 34 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.895 $Y=2.06
+ $X2=7.535 $Y2=2.06
r141 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.45 $Y=1.975
+ $X2=7.535 $Y2=2.06
r142 31 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.45 $Y=0.995
+ $X2=7.45 $Y2=0.805
r143 31 32 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=7.45 $Y=0.995
+ $X2=7.45 $Y2=1.975
r144 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.655 $Y=2.98
+ $X2=6.49 $Y2=2.98
r145 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.895 $Y=2.98
+ $X2=7.98 $Y2=2.895
r146 29 30 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.895 $Y=2.98
+ $X2=6.655 $Y2=2.98
r147 25 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=2.895
+ $X2=6.49 $Y2=2.98
r148 25 27 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.49 $Y=2.895
+ $X2=6.49 $Y2=2.59
r149 21 23 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=5.45 $Y=1.795
+ $X2=5.45 $Y2=1.05
r150 20 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=2.98 $X2=5
+ $Y2=2.98
r151 19 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.325 $Y=2.98
+ $X2=6.49 $Y2=2.98
r152 19 20 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=6.325 $Y=2.98
+ $X2=5.085 $Y2=2.98
r153 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.285 $Y=1.88
+ $X2=5.45 $Y2=1.795
r154 17 18 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.285 $Y=1.88
+ $X2=5.085 $Y2=1.88
r155 16 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=2.895 $X2=5
+ $Y2=2.98
r156 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5 $Y=1.965
+ $X2=5.085 $Y2=1.88
r157 15 16 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=5 $Y=1.965 $X2=5
+ $Y2=2.895
r158 14 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=2.98
+ $X2=3.96 $Y2=2.98
r159 13 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=2.98 $X2=5
+ $Y2=2.98
r160 13 14 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.915 $Y=2.98
+ $X2=4.125 $Y2=2.98
r161 4 27 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.735 $X2=6.49 $Y2=2.59
r162 3 38 600 $w=1.7e-07 $l=1.01491e-06 $layer=licon1_PDIFF $count=1 $X=3.815
+ $Y=1.735 $X2=3.96 $Y2=2.68
r163 2 45 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=7.17
+ $Y=0.555 $X2=7.31 $Y2=0.805
r164 1 23 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.31
+ $Y=0.775 $X2=5.45 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%A_803_81# 1 2 3 4 15 17 18 19 22 23 27 28
+ 30 32 33 37
c81 23 0 4.30949e-20 $X=5.595 $Y=2.24
c82 18 0 1.01058e-19 $X=4.245 $Y=0.35
c83 17 0 9.07277e-20 $X=6.305 $Y=0.35
r84 37 40 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=7.59 $Y=2.41
+ $X2=7.59 $Y2=2.505
r85 33 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.92 $Y=2.24
+ $X2=6.92 $Y2=2.41
r86 31 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.005 $Y=2.41
+ $X2=6.92 $Y2=2.41
r87 30 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.465 $Y=2.41
+ $X2=7.59 $Y2=2.41
r88 30 31 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.465 $Y=2.41
+ $X2=7.005 $Y2=2.41
r89 29 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=2.24
+ $X2=6.39 $Y2=2.24
r90 28 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.835 $Y=2.24
+ $X2=6.92 $Y2=2.24
r91 28 29 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.835 $Y=2.24
+ $X2=6.475 $Y2=2.24
r92 25 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=2.155
+ $X2=6.39 $Y2=2.24
r93 25 27 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=6.39 $Y=2.155
+ $X2=6.39 $Y2=0.765
r94 24 27 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.39 $Y=0.435
+ $X2=6.39 $Y2=0.765
r95 22 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=2.24
+ $X2=6.39 $Y2=2.24
r96 22 23 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.305 $Y=2.24
+ $X2=5.595 $Y2=2.24
r97 19 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.43 $Y=2.325
+ $X2=5.595 $Y2=2.24
r98 19 21 3.88182 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=5.43 $Y=2.325
+ $X2=5.43 $Y2=2.43
r99 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.305 $Y=0.35
+ $X2=6.39 $Y2=0.435
r100 17 18 134.396 $w=1.68e-07 $l=2.06e-06 $layer=LI1_cond $X=6.305 $Y=0.35
+ $X2=4.245 $Y2=0.35
r101 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.16 $Y=0.435
+ $X2=4.245 $Y2=0.35
r102 13 15 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.16 $Y=0.435
+ $X2=4.16 $Y2=0.55
r103 4 40 600 $w=1.7e-07 $l=9.07304e-07 $layer=licon1_PDIFF $count=1 $X=7.49
+ $Y=1.665 $X2=7.63 $Y2=2.505
r104 3 21 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=5.29
+ $Y=1.735 $X2=5.43 $Y2=2.43
r105 2 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.25
+ $Y=0.555 $X2=6.39 $Y2=0.765
r106 1 15 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.405 $X2=4.16 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%X 1 2 9 11 12 13 14 15
c22 15 0 1.15221e-19 $X=9.84 $Y=2.775
c23 12 0 1.59919e-19 $X=9.84 $Y=1.665
c24 11 0 1.1992e-19 $X=9.84 $Y=1.295
r25 15 37 2.04134 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=2.775
+ $X2=9.67 $Y2=2.86
r26 15 22 3.99151 $w=5.9e-07 $l=1.8e-07 $layer=LI1_cond $X=9.67 $Y=2.775
+ $X2=9.67 $Y2=2.595
r27 14 22 3.85178 $w=5.88e-07 $l=1.9e-07 $layer=LI1_cond $X=9.67 $Y=2.405
+ $X2=9.67 $Y2=2.595
r28 14 28 5.16949 $w=5.88e-07 $l=2.55e-07 $layer=LI1_cond $X=9.67 $Y=2.405
+ $X2=9.67 $Y2=2.15
r29 13 28 2.33134 $w=5.88e-07 $l=1.15e-07 $layer=LI1_cond $X=9.67 $Y=2.035
+ $X2=9.67 $Y2=2.15
r30 12 13 7.50083 $w=5.88e-07 $l=3.7e-07 $layer=LI1_cond $X=9.67 $Y=1.665
+ $X2=9.67 $Y2=2.035
r31 12 21 3.85178 $w=5.88e-07 $l=1.9e-07 $layer=LI1_cond $X=9.67 $Y=1.665
+ $X2=9.67 $Y2=1.475
r32 11 21 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=9.67 $Y=1.295
+ $X2=9.67 $Y2=1.475
r33 11 32 6.39252 $w=5.88e-07 $l=1.15e-07 $layer=LI1_cond $X=9.67 $Y=1.295
+ $X2=9.67 $Y2=1.18
r34 9 32 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=9.84 $Y=0.87 $X2=9.84
+ $Y2=1.18
r35 2 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.4
+ $Y=2.005 $X2=9.54 $Y2=2.86
r36 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.4
+ $Y=2.005 $X2=9.54 $Y2=2.15
r37 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.66 $X2=9.8 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_LP%VGND 1 2 3 12 16 18 21 23 24 25 31 32 33 39
+ 54 55 58
c91 16 0 1.75594e-19 $X=2.56 $Y=0.65
r92 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r93 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r94 52 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r95 51 52 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r96 49 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r97 48 51 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=9.36
+ $Y2=0
r98 48 49 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r99 46 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.6
+ $Y2=0
r100 46 48 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=3.12 $Y2=0
r101 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r102 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r103 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r104 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r105 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r106 39 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.6
+ $Y2=0
r107 39 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.16 $Y2=0
r108 37 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r109 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r110 33 52 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=9.36
+ $Y2=0
r111 33 49 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=3.12 $Y2=0
r112 31 51 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=9.365 $Y=0 $X2=9.36
+ $Y2=0
r113 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.365 $Y=0 $X2=9.45
+ $Y2=0
r114 30 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.84 $Y2=0
r115 30 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.45
+ $Y2=0
r116 25 28 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=9.01 $Y=0.815
+ $X2=9.01 $Y2=0.915
r117 23 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r118 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.03
+ $Y2=0
r119 22 41 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.2
+ $Y2=0
r120 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.03
+ $Y2=0
r121 20 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.45 $Y=0.085
+ $X2=9.45 $Y2=0
r122 20 21 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=9.45 $Y=0.085
+ $X2=9.45 $Y2=0.73
r123 19 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=0.815
+ $X2=9.01 $Y2=0.815
r124 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.365 $Y=0.815
+ $X2=9.45 $Y2=0.73
r125 18 19 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.365 $Y=0.815
+ $X2=9.175 $Y2=0.815
r126 14 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=0.085
+ $X2=2.6 $Y2=0
r127 14 16 26.0452 $w=2.48e-07 $l=5.65e-07 $layer=LI1_cond $X=2.6 $Y=0.085
+ $X2=2.6 $Y2=0.65
r128 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=0.085
+ $X2=1.03 $Y2=0
r129 10 12 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.03 $Y=0.085
+ $X2=1.03 $Y2=0.755
r130 3 28 182 $w=1.7e-07 $l=4.7571e-07 $layer=licon1_NDIFF $count=1 $X=8.645
+ $Y=0.66 $X2=9.01 $Y2=0.915
r131 2 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.505 $X2=2.56 $Y2=0.65
r132 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.545 $X2=1.07 $Y2=0.755
.ends

