* NGSPICE file created from sky130_fd_sc_lp__a311o_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_85_21# A1 a_427_47# VNB nshort w=840000u l=150000u
+  ad=5.502e+11p pd=4.67e+06u as=3.276e+11p ps=2.46e+06u
M1001 X a_85_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.6506e+12p ps=1.018e+07u
M1002 a_85_21# C1 a_657_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=4.032e+11p ps=3.16e+06u
M1003 VGND B1 a_85_21# VNB nshort w=840000u l=150000u
+  ad=1.0878e+12p pd=7.63e+06u as=0p ps=0u
M1004 VPWR a_85_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_341_367# A3 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1006 a_427_47# A2 a_355_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1007 a_657_367# B1 a_341_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_85_21# C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_341_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_355_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_341_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_85_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 X a_85_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

