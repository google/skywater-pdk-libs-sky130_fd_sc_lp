* File: sky130_fd_sc_lp__or4b_2.pxi.spice
* Created: Fri Aug 28 11:25:51 2020
* 
x_PM_SKY130_FD_SC_LP__OR4B_2%D_N N_D_N_M1012_g N_D_N_M1008_g D_N N_D_N_c_82_n
+ N_D_N_c_83_n PM_SKY130_FD_SC_LP__OR4B_2%D_N
x_PM_SKY130_FD_SC_LP__OR4B_2%A_189_21# N_A_189_21#_M1010_d N_A_189_21#_M1001_d
+ N_A_189_21#_M1006_d N_A_189_21#_M1002_g N_A_189_21#_M1000_g
+ N_A_189_21#_M1007_g N_A_189_21#_M1009_g N_A_189_21#_c_115_n
+ N_A_189_21#_c_105_n N_A_189_21#_c_197_p N_A_189_21#_c_128_p
+ N_A_189_21#_c_177_p N_A_189_21#_c_106_n N_A_189_21#_c_107_n
+ N_A_189_21#_c_108_n N_A_189_21#_c_109_n N_A_189_21#_c_110_n
+ N_A_189_21#_c_111_n N_A_189_21#_c_112_n PM_SKY130_FD_SC_LP__OR4B_2%A_189_21#
x_PM_SKY130_FD_SC_LP__OR4B_2%A N_A_M1010_g N_A_M1003_g A N_A_c_234_n N_A_c_235_n
+ PM_SKY130_FD_SC_LP__OR4B_2%A
x_PM_SKY130_FD_SC_LP__OR4B_2%B N_B_M1005_g N_B_c_271_n N_B_M1013_g B B B
+ PM_SKY130_FD_SC_LP__OR4B_2%B
x_PM_SKY130_FD_SC_LP__OR4B_2%C N_C_M1001_g N_C_M1004_g N_C_c_313_n N_C_c_314_n C
+ C N_C_c_316_n N_C_c_317_n PM_SKY130_FD_SC_LP__OR4B_2%C
x_PM_SKY130_FD_SC_LP__OR4B_2%A_31_131# N_A_31_131#_M1012_s N_A_31_131#_M1008_s
+ N_A_31_131#_c_355_n N_A_31_131#_M1011_g N_A_31_131#_M1006_g
+ N_A_31_131#_c_356_n N_A_31_131#_c_357_n N_A_31_131#_c_363_n
+ N_A_31_131#_c_364_n N_A_31_131#_c_358_n N_A_31_131#_c_359_n
+ N_A_31_131#_c_366_n N_A_31_131#_c_367_n N_A_31_131#_c_360_n
+ N_A_31_131#_c_368_n PM_SKY130_FD_SC_LP__OR4B_2%A_31_131#
x_PM_SKY130_FD_SC_LP__OR4B_2%VPWR N_VPWR_M1008_d N_VPWR_M1009_s N_VPWR_c_436_n
+ N_VPWR_c_437_n VPWR N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_435_n
+ N_VPWR_c_441_n N_VPWR_c_442_n PM_SKY130_FD_SC_LP__OR4B_2%VPWR
x_PM_SKY130_FD_SC_LP__OR4B_2%X N_X_M1002_d N_X_M1000_d N_X_c_467_n N_X_c_493_p
+ N_X_c_468_n X PM_SKY130_FD_SC_LP__OR4B_2%X
x_PM_SKY130_FD_SC_LP__OR4B_2%VGND N_VGND_M1012_d N_VGND_M1007_s N_VGND_M1005_d
+ N_VGND_M1011_d N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ N_VGND_c_503_n VGND N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n
+ N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n
+ PM_SKY130_FD_SC_LP__OR4B_2%VGND
cc_1 VNB N_D_N_M1012_g 0.0324559f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.865
cc_2 VNB N_D_N_M1008_g 0.00192992f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.045
cc_3 VNB N_D_N_c_82_n 0.0121499f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.46
cc_4 VNB N_D_N_c_83_n 0.0476552f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_5 VNB N_A_189_21#_M1002_g 0.0256774f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.46
cc_6 VNB N_A_189_21#_M1007_g 0.0238024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_189_21#_c_105_n 0.0110124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_189_21#_c_106_n 0.0068108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_189_21#_c_107_n 6.0864e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_189_21#_c_108_n 0.0130005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_189_21#_c_109_n 0.0342134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_189_21#_c_110_n 0.00203286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_189_21#_c_111_n 0.0015861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_189_21#_c_112_n 0.0385356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_M1010_g 0.0491142f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.865
cc_16 VNB N_A_c_234_n 0.0246412f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.46
cc_17 VNB N_A_c_235_n 0.00439671f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.46
cc_18 VNB N_B_M1005_g 0.0275629f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.865
cc_19 VNB N_B_c_271_n 0.0481898f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.625
cc_20 VNB N_B_M1013_g 0.00834689f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.045
cc_21 VNB B 0.0088524f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_C_M1004_g 0.0119263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_313_n 0.0168758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C_c_314_n 0.0144152f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.46
cc_25 VNB C 0.0032236f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.46
cc_26 VNB N_C_c_316_n 0.033377f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.46
cc_27 VNB N_C_c_317_n 0.0131197f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.665
cc_28 VNB N_A_31_131#_c_355_n 0.0209562f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.045
cc_29 VNB N_A_31_131#_c_356_n 0.04111f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_30 VNB N_A_31_131#_c_357_n 0.026992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_31_131#_c_358_n 0.00342807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_31_131#_c_359_n 0.00917466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_31_131#_c_360_n 0.0205271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_435_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_467_n 0.00159518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_468_n 0.0035438f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_37 VNB N_VGND_c_499_n 0.015212f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.46
cc_38 VNB N_VGND_c_500_n 0.00494127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_501_n 0.00234082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_502_n 0.0102016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_503_n 0.0168441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_504_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_505_n 0.0149607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_506_n 0.017305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_507_n 0.0263608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_508_n 0.0062884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_509_n 0.00568293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_510_n 0.217335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VPB N_D_N_M1008_g 0.032574f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.045
cc_50 VPB N_D_N_c_82_n 0.00755294f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.46
cc_51 VPB N_A_189_21#_M1000_g 0.0210796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_189_21#_M1009_g 0.0214157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_189_21#_c_115_n 0.00113824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_189_21#_c_109_n 0.0222717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_189_21#_c_112_n 0.00591248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_M1003_g 0.0231059f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.045
cc_57 VPB N_A_c_234_n 0.00640259f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.46
cc_58 VPB N_A_c_235_n 0.00470303f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.46
cc_59 VPB N_B_M1013_g 0.023929f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.045
cc_60 VPB B 0.00341869f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_61 VPB N_C_M1004_g 0.0239785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB C 0.00262668f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.46
cc_63 VPB N_A_31_131#_M1006_g 0.0349222f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.46
cc_64 VPB N_A_31_131#_c_356_n 4.00125e-19 $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.46
cc_65 VPB N_A_31_131#_c_363_n 0.0278694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_31_131#_c_364_n 0.0361619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_31_131#_c_359_n 0.00322958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_31_131#_c_366_n 0.0384401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_31_131#_c_367_n 0.00966343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_31_131#_c_368_n 0.0607537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_436_n 0.0184347f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=1.46
cc_72 VPB N_VPWR_c_437_n 0.0183629f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.46
cc_73 VPB N_VPWR_c_438_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=1.665
cc_74 VPB N_VPWR_c_439_n 0.0631068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_435_n 0.0995378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_441_n 0.0276197f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_442_n 0.00511034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_X_c_467_n 0.00128022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 N_D_N_M1012_g N_A_189_21#_M1002_g 0.0141264f $X=0.495 $Y=0.865 $X2=0 $Y2=0
cc_80 N_D_N_M1008_g N_A_189_21#_M1000_g 0.0141264f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_81 N_D_N_c_83_n N_A_189_21#_c_112_n 0.0141264f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_82 N_D_N_M1008_g N_A_31_131#_c_364_n 0.0236074f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_83 N_D_N_c_82_n N_A_31_131#_c_364_n 0.0275737f $X=0.315 $Y=1.46 $X2=0 $Y2=0
cc_84 N_D_N_c_83_n N_A_31_131#_c_364_n 0.00135495f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_85 N_D_N_M1012_g N_A_31_131#_c_358_n 0.0142219f $X=0.495 $Y=0.865 $X2=0 $Y2=0
cc_86 N_D_N_c_82_n N_A_31_131#_c_358_n 0.00200438f $X=0.315 $Y=1.46 $X2=0 $Y2=0
cc_87 N_D_N_M1012_g N_A_31_131#_c_359_n 0.012899f $X=0.495 $Y=0.865 $X2=0 $Y2=0
cc_88 N_D_N_c_82_n N_A_31_131#_c_359_n 0.0286577f $X=0.315 $Y=1.46 $X2=0 $Y2=0
cc_89 N_D_N_M1012_g N_A_31_131#_c_360_n 0.00825615f $X=0.495 $Y=0.865 $X2=0
+ $Y2=0
cc_90 N_D_N_c_82_n N_A_31_131#_c_360_n 0.0223805f $X=0.315 $Y=1.46 $X2=0 $Y2=0
cc_91 N_D_N_c_83_n N_A_31_131#_c_360_n 0.00664082f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_92 N_D_N_M1008_g X 2.36254e-19 $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_93 N_D_N_M1012_g N_VGND_c_499_n 0.0058738f $X=0.495 $Y=0.865 $X2=0 $Y2=0
cc_94 N_D_N_M1012_g N_VGND_c_507_n 0.00385987f $X=0.495 $Y=0.865 $X2=0 $Y2=0
cc_95 N_D_N_M1012_g N_VGND_c_510_n 0.0046122f $X=0.495 $Y=0.865 $X2=0 $Y2=0
cc_96 N_A_189_21#_M1007_g N_A_M1010_g 0.0250762f $X=1.45 $Y=0.655 $X2=0 $Y2=0
cc_97 N_A_189_21#_c_105_n N_A_M1010_g 0.0151289f $X=2.06 $Y=1.09 $X2=0 $Y2=0
cc_98 N_A_189_21#_c_106_n N_A_M1010_g 0.00595184f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_189_21#_c_111_n N_A_M1010_g 0.0034005f $X=1.51 $Y=1.335 $X2=0 $Y2=0
cc_100 N_A_189_21#_c_112_n N_A_M1010_g 3.77611e-19 $X=1.45 $Y=1.5 $X2=0 $Y2=0
cc_101 N_A_189_21#_M1009_g N_A_M1003_g 0.0167809f $X=1.45 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_189_21#_c_115_n N_A_M1003_g 0.00345788f $X=1.585 $Y=2.005 $X2=0 $Y2=0
cc_103 N_A_189_21#_c_128_p N_A_M1003_g 0.011364f $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_104 N_A_189_21#_M1009_g N_A_c_234_n 3.32099e-19 $X=1.45 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_189_21#_c_105_n N_A_c_234_n 0.00135123f $X=2.06 $Y=1.09 $X2=0 $Y2=0
cc_106 N_A_189_21#_c_128_p N_A_c_234_n 7.58005e-19 $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_107 N_A_189_21#_c_110_n N_A_c_234_n 0.00199598f $X=1.445 $Y=1.5 $X2=0 $Y2=0
cc_108 N_A_189_21#_c_112_n N_A_c_234_n 0.0169532f $X=1.45 $Y=1.5 $X2=0 $Y2=0
cc_109 N_A_189_21#_M1009_g N_A_c_235_n 5.01563e-19 $X=1.45 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_189_21#_c_105_n N_A_c_235_n 0.0347226f $X=2.06 $Y=1.09 $X2=0 $Y2=0
cc_111 N_A_189_21#_c_128_p N_A_c_235_n 0.0291377f $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_112 N_A_189_21#_c_110_n N_A_c_235_n 0.0377843f $X=1.445 $Y=1.5 $X2=0 $Y2=0
cc_113 N_A_189_21#_c_112_n N_A_c_235_n 3.57814e-19 $X=1.45 $Y=1.5 $X2=0 $Y2=0
cc_114 N_A_189_21#_c_106_n N_B_M1005_g 0.00584781f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_189_21#_c_107_n N_B_M1005_g 4.63661e-19 $X=3.15 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_189_21#_c_108_n N_B_M1005_g 5.64462e-19 $X=3.58 $Y=0.895 $X2=0 $Y2=0
cc_117 N_A_189_21#_c_105_n N_B_c_271_n 0.00140691f $X=2.06 $Y=1.09 $X2=0 $Y2=0
cc_118 N_A_189_21#_c_128_p N_B_c_271_n 5.39104e-19 $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_119 N_A_189_21#_c_128_p N_B_M1013_g 0.0126233f $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_120 N_A_189_21#_c_105_n B 0.0143048f $X=2.06 $Y=1.09 $X2=0 $Y2=0
cc_121 N_A_189_21#_c_128_p B 0.023783f $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_122 N_A_189_21#_c_106_n B 0.0125193f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A_189_21#_c_108_n B 0.00372126f $X=3.58 $Y=0.895 $X2=0 $Y2=0
cc_124 N_A_189_21#_c_109_n B 0.00733142f $X=3.58 $Y=2.005 $X2=0 $Y2=0
cc_125 N_A_189_21#_c_128_p N_C_M1004_g 0.0110812f $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_126 N_A_189_21#_c_109_n N_C_M1004_g 0.00175326f $X=3.58 $Y=2.005 $X2=0 $Y2=0
cc_127 N_A_189_21#_c_107_n N_C_c_313_n 0.00718662f $X=3.15 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A_189_21#_c_108_n N_C_c_313_n 0.00139902f $X=3.58 $Y=0.895 $X2=0 $Y2=0
cc_129 N_A_189_21#_c_107_n N_C_c_314_n 7.08121e-19 $X=3.15 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A_189_21#_c_108_n N_C_c_314_n 0.00680419f $X=3.58 $Y=0.895 $X2=0 $Y2=0
cc_131 N_A_189_21#_c_128_p C 0.0222853f $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_132 N_A_189_21#_c_108_n C 0.0161631f $X=3.58 $Y=0.895 $X2=0 $Y2=0
cc_133 N_A_189_21#_c_109_n C 0.0567473f $X=3.58 $Y=2.005 $X2=0 $Y2=0
cc_134 N_A_189_21#_c_128_p N_C_c_316_n 4.49126e-19 $X=3.415 $Y=2.095 $X2=0 $Y2=0
cc_135 N_A_189_21#_c_108_n N_C_c_316_n 0.00164811f $X=3.58 $Y=0.895 $X2=0 $Y2=0
cc_136 N_A_189_21#_c_109_n N_C_c_316_n 0.00205171f $X=3.58 $Y=2.005 $X2=0 $Y2=0
cc_137 N_A_189_21#_c_109_n N_C_c_317_n 0.00294925f $X=3.58 $Y=2.005 $X2=0 $Y2=0
cc_138 N_A_189_21#_c_107_n N_A_31_131#_c_355_n 0.0119063f $X=3.15 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_189_21#_c_108_n N_A_31_131#_c_355_n 0.00507821f $X=3.58 $Y=0.895
+ $X2=0 $Y2=0
cc_140 N_A_189_21#_c_128_p N_A_31_131#_M1006_g 0.0104154f $X=3.415 $Y=2.095
+ $X2=0 $Y2=0
cc_141 N_A_189_21#_c_109_n N_A_31_131#_M1006_g 0.00604126f $X=3.58 $Y=2.005
+ $X2=0 $Y2=0
cc_142 N_A_189_21#_c_109_n N_A_31_131#_c_356_n 0.0261849f $X=3.58 $Y=2.005 $X2=0
+ $Y2=0
cc_143 N_A_189_21#_c_108_n N_A_31_131#_c_357_n 0.0160707f $X=3.58 $Y=0.895 $X2=0
+ $Y2=0
cc_144 N_A_189_21#_c_109_n N_A_31_131#_c_357_n 0.00388225f $X=3.58 $Y=2.005
+ $X2=0 $Y2=0
cc_145 N_A_189_21#_c_109_n N_A_31_131#_c_363_n 0.0133758f $X=3.58 $Y=2.005 $X2=0
+ $Y2=0
cc_146 N_A_189_21#_M1000_g N_A_31_131#_c_364_n 0.00672425f $X=1.02 $Y=2.465
+ $X2=0 $Y2=0
cc_147 N_A_189_21#_M1002_g N_A_31_131#_c_358_n 0.00137503f $X=1.02 $Y=0.655
+ $X2=0 $Y2=0
cc_148 N_A_189_21#_M1002_g N_A_31_131#_c_359_n 0.0063081f $X=1.02 $Y=0.655 $X2=0
+ $Y2=0
cc_149 N_A_189_21#_M1000_g N_A_31_131#_c_366_n 0.014791f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_189_21#_M1009_g N_A_31_131#_c_366_n 0.0167407f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_189_21#_c_128_p N_A_31_131#_c_366_n 0.113976f $X=3.415 $Y=2.095 $X2=0
+ $Y2=0
cc_152 N_A_189_21#_c_177_p N_A_31_131#_c_366_n 0.00897693f $X=1.67 $Y=2.095
+ $X2=0 $Y2=0
cc_153 N_A_189_21#_c_109_n N_A_31_131#_c_366_n 0.00203388f $X=3.58 $Y=2.005
+ $X2=0 $Y2=0
cc_154 N_A_189_21#_M1002_g N_A_31_131#_c_360_n 5.35638e-19 $X=1.02 $Y=0.655
+ $X2=0 $Y2=0
cc_155 N_A_189_21#_c_128_p N_A_31_131#_c_368_n 5.18629e-19 $X=3.415 $Y=2.095
+ $X2=0 $Y2=0
cc_156 N_A_189_21#_c_115_n N_VPWR_M1009_s 0.00229403f $X=1.585 $Y=2.005 $X2=0
+ $Y2=0
cc_157 N_A_189_21#_c_128_p N_VPWR_M1009_s 0.0126538f $X=3.415 $Y=2.095 $X2=0
+ $Y2=0
cc_158 N_A_189_21#_c_177_p N_VPWR_M1009_s 9.65132e-19 $X=1.67 $Y=2.095 $X2=0
+ $Y2=0
cc_159 N_A_189_21#_M1000_g N_VPWR_c_436_n 0.0140592f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_189_21#_M1009_g N_VPWR_c_436_n 0.00160477f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_189_21#_M1000_g N_VPWR_c_437_n 0.00160477f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_189_21#_M1009_g N_VPWR_c_437_n 0.0140592f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_189_21#_M1000_g N_VPWR_c_438_n 0.00486043f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_189_21#_M1009_g N_VPWR_c_438_n 0.00486043f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_189_21#_M1000_g N_VPWR_c_435_n 0.00454594f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_189_21#_M1009_g N_VPWR_c_435_n 0.00454594f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_189_21#_M1002_g N_X_c_467_n 0.00388494f $X=1.02 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A_189_21#_M1000_g N_X_c_467_n 0.00381885f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_189_21#_M1007_g N_X_c_467_n 0.00123469f $X=1.45 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A_189_21#_M1009_g N_X_c_467_n 0.00120307f $X=1.45 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A_189_21#_c_115_n N_X_c_467_n 0.00800676f $X=1.585 $Y=2.005 $X2=0 $Y2=0
cc_172 N_A_189_21#_c_197_p N_X_c_467_n 9.927e-19 $X=1.67 $Y=1.09 $X2=0 $Y2=0
cc_173 N_A_189_21#_c_110_n N_X_c_467_n 0.0235079f $X=1.445 $Y=1.5 $X2=0 $Y2=0
cc_174 N_A_189_21#_c_111_n N_X_c_467_n 0.00710729f $X=1.51 $Y=1.335 $X2=0 $Y2=0
cc_175 N_A_189_21#_c_112_n N_X_c_467_n 0.0118324f $X=1.45 $Y=1.5 $X2=0 $Y2=0
cc_176 N_A_189_21#_M1002_g N_X_c_468_n 0.00714848f $X=1.02 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A_189_21#_M1007_g N_X_c_468_n 5.94388e-19 $X=1.45 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A_189_21#_c_197_p N_X_c_468_n 0.00956688f $X=1.67 $Y=1.09 $X2=0 $Y2=0
cc_179 N_A_189_21#_c_112_n N_X_c_468_n 0.00371629f $X=1.45 $Y=1.5 $X2=0 $Y2=0
cc_180 N_A_189_21#_M1000_g X 0.00633284f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_189_21#_c_112_n X 0.00401286f $X=1.45 $Y=1.5 $X2=0 $Y2=0
cc_182 N_A_189_21#_c_128_p A_436_385# 0.00368563f $X=3.415 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_189_21#_c_128_p A_508_385# 0.00906975f $X=3.415 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_189_21#_c_128_p A_616_385# 0.0018395f $X=3.415 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_189_21#_c_105_n N_VGND_M1007_s 0.00132228f $X=2.06 $Y=1.09 $X2=0
+ $Y2=0
cc_186 N_A_189_21#_c_197_p N_VGND_M1007_s 9.73829e-19 $X=1.67 $Y=1.09 $X2=0
+ $Y2=0
cc_187 N_A_189_21#_M1002_g N_VGND_c_499_n 0.011899f $X=1.02 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A_189_21#_M1007_g N_VGND_c_499_n 6.0835e-19 $X=1.45 $Y=0.655 $X2=0
+ $Y2=0
cc_189 N_A_189_21#_M1002_g N_VGND_c_500_n 6.17181e-19 $X=1.02 $Y=0.655 $X2=0
+ $Y2=0
cc_190 N_A_189_21#_M1007_g N_VGND_c_500_n 0.014682f $X=1.45 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A_189_21#_c_105_n N_VGND_c_500_n 0.0180881f $X=2.06 $Y=1.09 $X2=0 $Y2=0
cc_192 N_A_189_21#_c_197_p N_VGND_c_500_n 0.00992353f $X=1.67 $Y=1.09 $X2=0
+ $Y2=0
cc_193 N_A_189_21#_c_106_n N_VGND_c_500_n 0.0146167f $X=2.19 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A_189_21#_c_112_n N_VGND_c_500_n 2.40159e-19 $X=1.45 $Y=1.5 $X2=0 $Y2=0
cc_195 N_A_189_21#_c_108_n N_VGND_c_503_n 0.0200782f $X=3.58 $Y=0.895 $X2=0
+ $Y2=0
cc_196 N_A_189_21#_M1002_g N_VGND_c_504_n 0.00486043f $X=1.02 $Y=0.655 $X2=0
+ $Y2=0
cc_197 N_A_189_21#_M1007_g N_VGND_c_504_n 0.00486043f $X=1.45 $Y=0.655 $X2=0
+ $Y2=0
cc_198 N_A_189_21#_c_106_n N_VGND_c_505_n 0.0115062f $X=2.19 $Y=0.445 $X2=0
+ $Y2=0
cc_199 N_A_189_21#_c_107_n N_VGND_c_506_n 0.0185332f $X=3.15 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_A_189_21#_c_108_n N_VGND_c_506_n 0.00237343f $X=3.58 $Y=0.895 $X2=0
+ $Y2=0
cc_201 N_A_189_21#_M1010_d N_VGND_c_510_n 0.00458991f $X=2.05 $Y=0.235 $X2=0
+ $Y2=0
cc_202 N_A_189_21#_M1001_d N_VGND_c_510_n 0.00225167f $X=3.01 $Y=0.235 $X2=0
+ $Y2=0
cc_203 N_A_189_21#_M1002_g N_VGND_c_510_n 0.00824727f $X=1.02 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A_189_21#_M1007_g N_VGND_c_510_n 0.00824727f $X=1.45 $Y=0.655 $X2=0
+ $Y2=0
cc_205 N_A_189_21#_c_106_n N_VGND_c_510_n 0.0081747f $X=2.19 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_189_21#_c_107_n N_VGND_c_510_n 0.0123939f $X=3.15 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_189_21#_c_108_n N_VGND_c_510_n 0.0048982f $X=3.58 $Y=0.895 $X2=0
+ $Y2=0
cc_208 N_A_M1010_g N_B_M1005_g 0.0240943f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A_M1010_g N_B_c_271_n 0.0088837f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_210 N_A_c_234_n N_B_c_271_n 0.0354407f $X=2.015 $Y=1.51 $X2=0 $Y2=0
cc_211 N_A_c_235_n N_B_c_271_n 0.00296712f $X=2.015 $Y=1.51 $X2=0 $Y2=0
cc_212 N_A_M1003_g N_B_M1013_g 0.0354407f $X=2.105 $Y=2.135 $X2=0 $Y2=0
cc_213 N_A_M1010_g B 0.00110038f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A_c_234_n B 4.65361e-19 $X=2.015 $Y=1.51 $X2=0 $Y2=0
cc_215 N_A_c_235_n B 0.0394464f $X=2.015 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A_M1003_g N_A_31_131#_c_366_n 0.00915279f $X=2.105 $Y=2.135 $X2=0 $Y2=0
cc_217 N_A_M1010_g N_VGND_c_500_n 0.00399847f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A_M1010_g N_VGND_c_501_n 6.10505e-19 $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A_M1010_g N_VGND_c_505_n 0.00585385f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_M1010_g N_VGND_c_510_n 0.0108947f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_221 N_B_M1013_g N_C_M1004_g 0.0303317f $X=2.465 $Y=2.135 $X2=0 $Y2=0
cc_222 N_B_M1005_g N_C_c_313_n 0.0169653f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_223 B N_C_c_314_n 8.21294e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_224 N_B_c_271_n C 4.00854e-19 $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_225 N_B_M1013_g C 3.21055e-19 $X=2.465 $Y=2.135 $X2=0 $Y2=0
cc_226 B C 0.0557603f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_227 N_B_c_271_n N_C_c_316_n 0.0204862f $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_228 N_B_M1005_g N_C_c_317_n 7.94268e-19 $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_229 N_B_c_271_n N_C_c_317_n 0.0051273f $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_230 B N_C_c_317_n 0.00723226f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_231 N_B_M1013_g N_A_31_131#_c_366_n 0.00884f $X=2.465 $Y=2.135 $X2=0 $Y2=0
cc_232 N_B_M1005_g N_VGND_c_501_n 0.00866798f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_233 N_B_c_271_n N_VGND_c_501_n 9.3227e-19 $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_234 B N_VGND_c_501_n 0.0192745f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_235 N_B_M1005_g N_VGND_c_505_n 0.00486043f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_236 N_B_M1005_g N_VGND_c_510_n 0.00808569f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_237 B N_VGND_c_510_n 0.00161401f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_238 N_C_c_313_n N_A_31_131#_c_355_n 0.0128416f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_239 N_C_M1004_g N_A_31_131#_c_356_n 0.00306742f $X=3.005 $Y=2.135 $X2=0 $Y2=0
cc_240 C N_A_31_131#_c_356_n 7.2892e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_241 N_C_c_316_n N_A_31_131#_c_356_n 0.017271f $X=3.095 $Y=1.29 $X2=0 $Y2=0
cc_242 N_C_c_317_n N_A_31_131#_c_356_n 0.00284552f $X=3.095 $Y=1.125 $X2=0 $Y2=0
cc_243 N_C_c_314_n N_A_31_131#_c_357_n 0.00971271f $X=2.97 $Y=0.915 $X2=0 $Y2=0
cc_244 N_C_M1004_g N_A_31_131#_c_363_n 0.0513544f $X=3.005 $Y=2.135 $X2=0 $Y2=0
cc_245 C N_A_31_131#_c_363_n 0.00122553f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_246 N_C_M1004_g N_A_31_131#_c_366_n 0.00884f $X=3.005 $Y=2.135 $X2=0 $Y2=0
cc_247 N_C_c_313_n N_VGND_c_501_n 0.0038527f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_248 N_C_c_313_n N_VGND_c_506_n 0.00547966f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_249 N_C_c_313_n N_VGND_c_510_n 0.0101914f $X=2.97 $Y=0.765 $X2=0 $Y2=0
cc_250 N_A_31_131#_c_364_n N_VPWR_M1008_d 0.00864985f $X=0.65 $Y=2.09 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_31_131#_c_359_n N_VPWR_M1008_d 0.00200168f $X=0.74 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_31_131#_c_366_n N_VPWR_M1008_d 0.00277086f $X=3.1 $Y=2.44 $X2=-0.19
+ $Y2=-0.245
cc_253 N_A_31_131#_c_366_n N_VPWR_M1009_s 0.005149f $X=3.1 $Y=2.44 $X2=0 $Y2=0
cc_254 N_A_31_131#_c_364_n N_VPWR_c_436_n 0.0158579f $X=0.65 $Y=2.09 $X2=0 $Y2=0
cc_255 N_A_31_131#_c_366_n N_VPWR_c_436_n 0.00633739f $X=3.1 $Y=2.44 $X2=0 $Y2=0
cc_256 N_A_31_131#_c_366_n N_VPWR_c_437_n 0.021555f $X=3.1 $Y=2.44 $X2=0 $Y2=0
cc_257 N_A_31_131#_c_367_n N_VPWR_c_439_n 0.0192467f $X=3.265 $Y=2.88 $X2=0
+ $Y2=0
cc_258 N_A_31_131#_c_368_n N_VPWR_c_439_n 0.00210337f $X=3.365 $Y=2.88 $X2=0
+ $Y2=0
cc_259 N_A_31_131#_c_364_n N_VPWR_c_435_n 6.50158e-19 $X=0.65 $Y=2.09 $X2=0
+ $Y2=0
cc_260 N_A_31_131#_c_366_n N_VPWR_c_435_n 0.0639779f $X=3.1 $Y=2.44 $X2=0 $Y2=0
cc_261 N_A_31_131#_c_367_n N_VPWR_c_435_n 0.0127274f $X=3.265 $Y=2.88 $X2=0
+ $Y2=0
cc_262 N_A_31_131#_c_366_n N_X_M1000_d 0.00493494f $X=3.1 $Y=2.44 $X2=0 $Y2=0
cc_263 N_A_31_131#_c_359_n N_X_c_467_n 0.0473763f $X=0.74 $Y=1.92 $X2=0 $Y2=0
cc_264 N_A_31_131#_c_358_n N_X_c_468_n 0.0128445f $X=0.65 $Y=1.07 $X2=0 $Y2=0
cc_265 N_A_31_131#_c_364_n X 0.0209498f $X=0.65 $Y=2.09 $X2=0 $Y2=0
cc_266 N_A_31_131#_c_359_n X 0.00521446f $X=0.74 $Y=1.92 $X2=0 $Y2=0
cc_267 N_A_31_131#_c_366_n X 0.018725f $X=3.1 $Y=2.44 $X2=0 $Y2=0
cc_268 N_A_31_131#_c_358_n N_VGND_M1012_d 0.00373869f $X=0.65 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_31_131#_c_358_n N_VGND_c_499_n 0.0169249f $X=0.65 $Y=1.07 $X2=0 $Y2=0
cc_270 N_A_31_131#_c_360_n N_VGND_c_499_n 0.00803151f $X=0.28 $Y=0.865 $X2=0
+ $Y2=0
cc_271 N_A_31_131#_c_355_n N_VGND_c_503_n 0.00327088f $X=3.365 $Y=0.765 $X2=0
+ $Y2=0
cc_272 N_A_31_131#_c_357_n N_VGND_c_503_n 0.00111336f $X=3.575 $Y=0.84 $X2=0
+ $Y2=0
cc_273 N_A_31_131#_c_355_n N_VGND_c_506_n 0.00425023f $X=3.365 $Y=0.765 $X2=0
+ $Y2=0
cc_274 N_A_31_131#_c_360_n N_VGND_c_507_n 0.00489913f $X=0.28 $Y=0.865 $X2=0
+ $Y2=0
cc_275 N_A_31_131#_c_355_n N_VGND_c_510_n 0.00685068f $X=3.365 $Y=0.765 $X2=0
+ $Y2=0
cc_276 N_A_31_131#_c_360_n N_VGND_c_510_n 0.00926534f $X=0.28 $Y=0.865 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_435_n N_X_M1000_d 0.00396212f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_278 N_X_c_493_p N_VGND_c_504_n 0.0124525f $X=1.235 $Y=0.42 $X2=0 $Y2=0
cc_279 N_X_M1002_d N_VGND_c_510_n 0.00536646f $X=1.095 $Y=0.235 $X2=0 $Y2=0
cc_280 N_X_c_493_p N_VGND_c_510_n 0.00730901f $X=1.235 $Y=0.42 $X2=0 $Y2=0
