* File: sky130_fd_sc_lp__o211a_m.spice
* Created: Wed Sep  2 10:14:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211a_m.pex.spice"
.subckt sky130_fd_sc_lp__o211a_m  VNB VPB A1 A2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_80_60#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_217_49#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_A_217_49#_M1005_d N_A2_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_488_49# N_B1_M1008_g N_A_217_49#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_80_60#_M1006_d N_C1_M1006_g A_488_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_60#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09975 AS=0.1113 PD=0.895 PS=1.37 NRD=44.5417 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1007 A_300_371# N_A1_M1007_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.09975 PD=0.63 PS=0.895 NRD=23.443 NRS=46.886 M=1 R=2.8
+ SA=75000.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_80_60#_M1009_d N_A2_M1009_g A_300_371# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_A_80_60#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06825 AS=0.0819 PD=0.745 PS=0.81 NRD=21.0987 NRS=51.5943 M=1 R=2.8
+ SA=75001.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_80_60#_M1001_d N_C1_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.06825 PD=1.37 PS=0.745 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o211a_m.pxi.spice"
*
.ends
*
*
