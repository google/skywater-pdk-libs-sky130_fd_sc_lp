* File: sky130_fd_sc_lp__iso1n_lp.pxi.spice
* Created: Wed Sep  2 09:58:08 2020
* 
x_PM_SKY130_FD_SC_LP__ISO1N_LP%SLEEP_B N_SLEEP_B_M1006_g N_SLEEP_B_M1004_g
+ N_SLEEP_B_M1001_g N_SLEEP_B_M1009_g SLEEP_B SLEEP_B N_SLEEP_B_c_62_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP%SLEEP_B
x_PM_SKY130_FD_SC_LP__ISO1N_LP%A_27_93# N_A_27_93#_M1006_s N_A_27_93#_M1004_s
+ N_A_27_93#_c_101_n N_A_27_93#_M1011_g N_A_27_93#_c_102_n N_A_27_93#_M1007_g
+ N_A_27_93#_M1000_g N_A_27_93#_c_103_n N_A_27_93#_c_108_n N_A_27_93#_c_104_n
+ N_A_27_93#_c_105_n N_A_27_93#_c_110_n N_A_27_93#_c_111_n N_A_27_93#_c_112_n
+ N_A_27_93#_c_113_n N_A_27_93#_c_106_n PM_SKY130_FD_SC_LP__ISO1N_LP%A_27_93#
x_PM_SKY130_FD_SC_LP__ISO1N_LP%A N_A_M1013_g N_A_M1002_g N_A_M1012_g A
+ N_A_c_172_n N_A_c_170_n PM_SKY130_FD_SC_LP__ISO1N_LP%A
x_PM_SKY130_FD_SC_LP__ISO1N_LP%A_340_93# N_A_340_93#_M1007_d N_A_340_93#_M1013_d
+ N_A_340_93#_c_213_n N_A_340_93#_M1003_g N_A_340_93#_M1008_g
+ N_A_340_93#_c_214_n N_A_340_93#_M1005_g N_A_340_93#_M1010_g
+ N_A_340_93#_c_215_n N_A_340_93#_c_216_n N_A_340_93#_c_217_n
+ N_A_340_93#_c_222_n N_A_340_93#_c_223_n N_A_340_93#_c_224_n
+ N_A_340_93#_c_268_p N_A_340_93#_c_247_n N_A_340_93#_c_218_n
+ N_A_340_93#_c_219_n PM_SKY130_FD_SC_LP__ISO1N_LP%A_340_93#
x_PM_SKY130_FD_SC_LP__ISO1N_LP%VPWR N_VPWR_M1009_d N_VPWR_M1008_s N_VPWR_c_289_n
+ N_VPWR_c_290_n VPWR N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n
+ N_VPWR_c_288_n N_VPWR_c_295_n N_VPWR_c_296_n PM_SKY130_FD_SC_LP__ISO1N_LP%VPWR
x_PM_SKY130_FD_SC_LP__ISO1N_LP%X N_X_M1005_d N_X_M1010_d X X X X X N_X_c_330_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP%X
x_PM_SKY130_FD_SC_LP__ISO1N_LP%KAGND N_KAGND_M1001_d N_KAGND_M1012_d KAGND
+ N_KAGND_c_344_n N_KAGND_c_345_n N_KAGND_c_346_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP%KAGND
x_PM_SKY130_FD_SC_LP__ISO1N_LP%VGND VGND N_VGND_c_398_n N_VGND_c_399_n VGND
+ PM_SKY130_FD_SC_LP__ISO1N_LP%VGND
cc_1 VNB N_SLEEP_B_M1006_g 0.0351755f $X=-0.22 $Y=-0.245 $X2=0.475 $Y2=0.675
cc_2 VNB N_SLEEP_B_M1001_g 0.0312541f $X=-0.22 $Y=-0.245 $X2=0.835 $Y2=0.675
cc_3 VNB SLEEP_B 0.00827905f $X=-0.22 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_SLEEP_B_c_62_n 0.0506752f $X=-0.22 $Y=-0.245 $X2=0.995 $Y2=1.485
cc_5 VNB N_A_27_93#_c_101_n 0.0137894f $X=-0.22 $Y=-0.245 $X2=0.695 $Y2=2.655
cc_6 VNB N_A_27_93#_c_102_n 0.0144144f $X=-0.22 $Y=-0.245 $X2=0.835 $Y2=0.675
cc_7 VNB N_A_27_93#_c_103_n 0.0250605f $X=-0.22 $Y=-0.245 $X2=0.475 $Y2=1.32
cc_8 VNB N_A_27_93#_c_104_n 0.0210476f $X=-0.22 $Y=-0.245 $X2=0.995 $Y2=1.485
cc_9 VNB N_A_27_93#_c_105_n 0.0332044f $X=-0.22 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_93#_c_106_n 0.0399924f $X=-0.22 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_M1013_g 5.47154e-19 $X=-0.22 $Y=-0.245 $X2=0.475 $Y2=0.675
cc_12 VNB N_A_M1002_g 0.0300075f $X=-0.22 $Y=-0.245 $X2=0.695 $Y2=2.655
cc_13 VNB N_A_M1012_g 0.0303404f $X=-0.22 $Y=-0.245 $X2=0.835 $Y2=0.675
cc_14 VNB N_A_c_170_n 0.055099f $X=-0.22 $Y=-0.245 $X2=0.475 $Y2=1.32
cc_15 VNB N_A_340_93#_c_213_n 0.016294f $X=-0.22 $Y=-0.245 $X2=0.695 $Y2=2.655
cc_16 VNB N_A_340_93#_c_214_n 0.0198943f $X=-0.22 $Y=-0.245 $X2=1.085 $Y2=2.655
cc_17 VNB N_A_340_93#_c_215_n 0.00163989f $X=-0.22 $Y=-0.245 $X2=0.695 $Y2=1.655
cc_18 VNB N_A_340_93#_c_216_n 0.0170924f $X=-0.22 $Y=-0.245 $X2=0.835 $Y2=1.655
cc_19 VNB N_A_340_93#_c_217_n 0.00433003f $X=-0.22 $Y=-0.245 $X2=0.995 $Y2=1.655
cc_20 VNB N_A_340_93#_c_218_n 0.00767951f $X=-0.22 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_340_93#_c_219_n 0.0637404f $X=-0.22 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_288_n 0.163682f $X=-0.22 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_330_n 0.0588801f $X=-0.22 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_KAGND_c_344_n 0.00710967f $X=-0.22 $Y=-0.245 $X2=0.835 $Y2=0.675
cc_25 VNB N_KAGND_c_345_n 0.00738504f $X=-0.22 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_KAGND_c_346_n 0.0258545f $X=-0.22 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB N_VGND_c_398_n 0.230446f $X=-0.22 $Y=-0.245 $X2=0.695 $Y2=1.99
cc_28 VNB N_VGND_c_399_n 0.112118f $X=-0.22 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_SLEEP_B_M1004_g 0.0392373f $X=-0.22 $Y=1.655 $X2=0.695 $Y2=2.655
cc_30 VPB N_SLEEP_B_M1009_g 0.0342064f $X=-0.22 $Y=1.655 $X2=1.085 $Y2=2.655
cc_31 VPB SLEEP_B 0.00130528f $X=-0.22 $Y=1.655 $X2=0.635 $Y2=1.21
cc_32 VPB N_SLEEP_B_c_62_n 0.0433147f $X=-0.22 $Y=1.655 $X2=0.995 $Y2=1.485
cc_33 VPB N_A_27_93#_M1000_g 0.0335159f $X=-0.22 $Y=1.655 $X2=1.085 $Y2=2.655
cc_34 VPB N_A_27_93#_c_108_n 0.0163859f $X=-0.22 $Y=1.655 $X2=0.995 $Y2=1.655
cc_35 VPB N_A_27_93#_c_105_n 0.027029f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_27_93#_c_110_n 0.0199287f $X=-0.22 $Y=1.655 $X2=0.85 $Y2=1.665
cc_37 VPB N_A_27_93#_c_111_n 0.0255732f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_27_93#_c_112_n 0.0209213f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_93#_c_113_n 0.00184461f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_93#_c_106_n 0.0111978f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_M1013_g 0.0599872f $X=-0.22 $Y=1.655 $X2=0.475 $Y2=0.675
cc_42 VPB N_A_c_172_n 0.00687916f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_340_93#_M1008_g 0.0210318f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_340_93#_M1010_g 0.0196807f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_340_93#_c_222_n 0.0111024f $X=-0.22 $Y=1.655 $X2=1.085 $Y2=1.655
cc_46 VPB N_A_340_93#_c_223_n 0.0124046f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_340_93#_c_224_n 0.00414064f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_340_93#_c_219_n 0.00454175f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_289_n 0.0179168f $X=-0.22 $Y=1.655 $X2=0.835 $Y2=1.32
cc_50 VPB N_VPWR_c_290_n 0.0152895f $X=-0.22 $Y=1.655 $X2=1.085 $Y2=1.99
cc_51 VPB N_VPWR_c_291_n 0.0386257f $X=-0.22 $Y=1.655 $X2=0.635 $Y2=1.21
cc_52 VPB N_VPWR_c_292_n 0.0305824f $X=-0.22 $Y=1.655 $X2=0.695 $Y2=1.655
cc_53 VPB N_VPWR_c_293_n 0.027323f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_288_n 0.102625f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_295_n 0.00632158f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_296_n 0.00601838f $X=-0.22 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_X_c_330_n 0.0631849f $X=-0.22 $Y=1.655 $X2=0.635 $Y2=1.58
cc_58 N_SLEEP_B_M1001_g N_A_27_93#_c_101_n 0.0207816f $X=0.835 $Y=0.675 $X2=0
+ $Y2=0
cc_59 N_SLEEP_B_c_62_n N_A_27_93#_M1000_g 0.0173581f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_60 N_SLEEP_B_M1006_g N_A_27_93#_c_104_n 0.00769044f $X=0.475 $Y=0.675 $X2=0
+ $Y2=0
cc_61 N_SLEEP_B_M1006_g N_A_27_93#_c_105_n 0.0146972f $X=0.475 $Y=0.675 $X2=0
+ $Y2=0
cc_62 N_SLEEP_B_M1004_g N_A_27_93#_c_105_n 0.00556354f $X=0.695 $Y=2.655 $X2=0
+ $Y2=0
cc_63 SLEEP_B N_A_27_93#_c_105_n 0.0672664f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_SLEEP_B_c_62_n N_A_27_93#_c_105_n 0.014424f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_65 N_SLEEP_B_M1004_g N_A_27_93#_c_110_n 0.0050656f $X=0.695 $Y=2.655 $X2=0
+ $Y2=0
cc_66 N_SLEEP_B_M1004_g N_A_27_93#_c_111_n 0.0163715f $X=0.695 $Y=2.655 $X2=0
+ $Y2=0
cc_67 N_SLEEP_B_M1009_g N_A_27_93#_c_111_n 0.0151084f $X=1.085 $Y=2.655 $X2=0
+ $Y2=0
cc_68 N_SLEEP_B_c_62_n N_A_27_93#_c_111_n 4.17406e-19 $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_69 SLEEP_B N_A_27_93#_c_112_n 0.0482347f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_SLEEP_B_c_62_n N_A_27_93#_c_112_n 0.00485258f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_71 SLEEP_B N_A_27_93#_c_113_n 0.0449538f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_SLEEP_B_c_62_n N_A_27_93#_c_113_n 0.00666802f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_73 N_SLEEP_B_M1001_g N_A_27_93#_c_106_n 0.00504883f $X=0.835 $Y=0.675 $X2=0
+ $Y2=0
cc_74 SLEEP_B N_A_27_93#_c_106_n 0.00669964f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_SLEEP_B_c_62_n N_A_27_93#_c_106_n 0.042841f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_76 N_SLEEP_B_M1009_g N_VPWR_c_289_n 0.00389024f $X=1.085 $Y=2.655 $X2=0 $Y2=0
cc_77 N_SLEEP_B_M1004_g N_VPWR_c_291_n 0.00510437f $X=0.695 $Y=2.655 $X2=0 $Y2=0
cc_78 N_SLEEP_B_M1009_g N_VPWR_c_291_n 0.00510437f $X=1.085 $Y=2.655 $X2=0 $Y2=0
cc_79 N_SLEEP_B_M1004_g N_VPWR_c_288_n 0.00515964f $X=0.695 $Y=2.655 $X2=0 $Y2=0
cc_80 N_SLEEP_B_M1009_g N_VPWR_c_288_n 0.00515964f $X=1.085 $Y=2.655 $X2=0 $Y2=0
cc_81 N_SLEEP_B_M1006_g N_KAGND_c_344_n 0.00145275f $X=0.475 $Y=0.675 $X2=0
+ $Y2=0
cc_82 N_SLEEP_B_M1001_g N_KAGND_c_344_n 0.00845552f $X=0.835 $Y=0.675 $X2=0
+ $Y2=0
cc_83 SLEEP_B N_KAGND_c_344_n 0.0128024f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_SLEEP_B_c_62_n N_KAGND_c_344_n 0.00105915f $X=0.995 $Y=1.485 $X2=0 $Y2=0
cc_85 N_SLEEP_B_M1006_g N_KAGND_c_346_n 0.00973274f $X=0.475 $Y=0.675 $X2=0
+ $Y2=0
cc_86 N_SLEEP_B_M1001_g N_KAGND_c_346_n 0.00359794f $X=0.835 $Y=0.675 $X2=0
+ $Y2=0
cc_87 SLEEP_B N_KAGND_c_346_n 0.0144484f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_SLEEP_B_M1006_g N_VGND_c_398_n 0.00310524f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_89 N_SLEEP_B_M1001_g N_VGND_c_398_n 0.00310524f $X=0.835 $Y=0.675 $X2=0 $Y2=0
cc_90 N_SLEEP_B_M1006_g N_VGND_c_399_n 0.00510437f $X=0.475 $Y=0.675 $X2=0 $Y2=0
cc_91 N_SLEEP_B_M1001_g N_VGND_c_399_n 0.0048834f $X=0.835 $Y=0.675 $X2=0 $Y2=0
cc_92 N_A_27_93#_c_108_n N_A_M1013_g 0.0510623f $X=1.535 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_27_93#_c_111_n N_A_M1013_g 5.90946e-19 $X=1.37 $Y=2.245 $X2=0 $Y2=0
cc_94 N_A_27_93#_c_102_n N_A_M1002_g 0.0284349f $X=1.625 $Y=0.96 $X2=0 $Y2=0
cc_95 N_A_27_93#_c_113_n N_A_c_172_n 0.0237482f $X=1.535 $Y=1.48 $X2=0 $Y2=0
cc_96 N_A_27_93#_c_106_n N_A_c_172_n 0.00123182f $X=1.535 $Y=1.48 $X2=0 $Y2=0
cc_97 N_A_27_93#_c_113_n N_A_c_170_n 0.00399595f $X=1.535 $Y=1.48 $X2=0 $Y2=0
cc_98 N_A_27_93#_c_106_n N_A_c_170_n 0.0510623f $X=1.535 $Y=1.48 $X2=0 $Y2=0
cc_99 N_A_27_93#_c_102_n N_A_340_93#_c_215_n 0.00379803f $X=1.625 $Y=0.96 $X2=0
+ $Y2=0
cc_100 N_A_27_93#_c_103_n N_A_340_93#_c_217_n 0.00494368f $X=1.625 $Y=1.035
+ $X2=0 $Y2=0
cc_101 N_A_27_93#_c_111_n N_A_340_93#_c_222_n 0.00729784f $X=1.37 $Y=2.245 $X2=0
+ $Y2=0
cc_102 N_A_27_93#_c_113_n N_A_340_93#_c_222_n 0.00138084f $X=1.535 $Y=1.48 $X2=0
+ $Y2=0
cc_103 N_A_27_93#_c_113_n N_A_340_93#_c_224_n 0.00761536f $X=1.535 $Y=1.48 $X2=0
+ $Y2=0
cc_104 N_A_27_93#_c_102_n N_A_340_93#_c_218_n 0.00268639f $X=1.625 $Y=0.96 $X2=0
+ $Y2=0
cc_105 N_A_27_93#_M1000_g N_VPWR_c_289_n 0.00369545f $X=1.625 $Y=2.655 $X2=0
+ $Y2=0
cc_106 N_A_27_93#_c_108_n N_VPWR_c_289_n 5.1863e-19 $X=1.535 $Y=1.985 $X2=0
+ $Y2=0
cc_107 N_A_27_93#_c_111_n N_VPWR_c_289_n 0.0261221f $X=1.37 $Y=2.245 $X2=0 $Y2=0
cc_108 N_A_27_93#_c_110_n N_VPWR_c_291_n 0.00586831f $X=0.48 $Y=2.655 $X2=0
+ $Y2=0
cc_109 N_A_27_93#_M1000_g N_VPWR_c_292_n 0.00510437f $X=1.625 $Y=2.655 $X2=0
+ $Y2=0
cc_110 N_A_27_93#_M1000_g N_VPWR_c_288_n 0.00515964f $X=1.625 $Y=2.655 $X2=0
+ $Y2=0
cc_111 N_A_27_93#_c_110_n N_VPWR_c_288_n 0.00796314f $X=0.48 $Y=2.655 $X2=0
+ $Y2=0
cc_112 N_A_27_93#_c_101_n N_KAGND_c_344_n 0.018482f $X=1.265 $Y=0.96 $X2=0 $Y2=0
cc_113 N_A_27_93#_c_102_n N_KAGND_c_344_n 0.00196398f $X=1.625 $Y=0.96 $X2=0
+ $Y2=0
cc_114 N_A_27_93#_c_103_n N_KAGND_c_344_n 0.00103068f $X=1.625 $Y=1.035 $X2=0
+ $Y2=0
cc_115 N_A_27_93#_c_104_n N_KAGND_c_344_n 0.00492012f $X=0.242 $Y=0.763 $X2=0
+ $Y2=0
cc_116 N_A_27_93#_c_113_n N_KAGND_c_344_n 0.00488772f $X=1.535 $Y=1.48 $X2=0
+ $Y2=0
cc_117 N_A_27_93#_M1006_s N_KAGND_c_346_n 0.00115614f $X=0.135 $Y=0.465 $X2=0
+ $Y2=0
cc_118 N_A_27_93#_c_102_n N_KAGND_c_346_n 0.00999476f $X=1.625 $Y=0.96 $X2=0
+ $Y2=0
cc_119 N_A_27_93#_c_104_n N_KAGND_c_346_n 0.0314646f $X=0.242 $Y=0.763 $X2=0
+ $Y2=0
cc_120 N_A_27_93#_c_101_n N_VGND_c_398_n 0.00310524f $X=1.265 $Y=0.96 $X2=0
+ $Y2=0
cc_121 N_A_27_93#_c_102_n N_VGND_c_398_n 0.00310524f $X=1.625 $Y=0.96 $X2=0
+ $Y2=0
cc_122 N_A_27_93#_c_104_n N_VGND_c_398_n 0.00266832f $X=0.242 $Y=0.763 $X2=0
+ $Y2=0
cc_123 N_A_27_93#_c_101_n N_VGND_c_399_n 0.00372327f $X=1.265 $Y=0.96 $X2=0
+ $Y2=0
cc_124 N_A_27_93#_c_102_n N_VGND_c_399_n 0.00510437f $X=1.625 $Y=0.96 $X2=0
+ $Y2=0
cc_125 N_A_27_93#_c_104_n N_VGND_c_399_n 0.0081917f $X=0.242 $Y=0.763 $X2=0
+ $Y2=0
cc_126 N_A_M1012_g N_A_340_93#_c_213_n 0.0270073f $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_127 N_A_M1002_g N_A_340_93#_c_215_n 0.00431365f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_128 N_A_M1002_g N_A_340_93#_c_216_n 0.00762601f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_129 N_A_M1012_g N_A_340_93#_c_216_n 0.0108589f $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_130 N_A_c_172_n N_A_340_93#_c_216_n 0.0379774f $X=2.415 $Y=1.48 $X2=0 $Y2=0
cc_131 N_A_c_170_n N_A_340_93#_c_216_n 0.00149434f $X=2.475 $Y=1.48 $X2=0 $Y2=0
cc_132 N_A_M1002_g N_A_340_93#_c_217_n 0.00232854f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_133 N_A_c_172_n N_A_340_93#_c_217_n 0.0130022f $X=2.415 $Y=1.48 $X2=0 $Y2=0
cc_134 N_A_c_170_n N_A_340_93#_c_217_n 0.00391752f $X=2.475 $Y=1.48 $X2=0 $Y2=0
cc_135 N_A_M1013_g N_A_340_93#_c_222_n 0.0114604f $X=1.985 $Y=2.655 $X2=0 $Y2=0
cc_136 N_A_c_172_n N_A_340_93#_c_223_n 0.0192012f $X=2.415 $Y=1.48 $X2=0 $Y2=0
cc_137 N_A_c_170_n N_A_340_93#_c_223_n 0.00143458f $X=2.475 $Y=1.48 $X2=0 $Y2=0
cc_138 N_A_M1013_g N_A_340_93#_c_224_n 0.00477088f $X=1.985 $Y=2.655 $X2=0 $Y2=0
cc_139 N_A_c_172_n N_A_340_93#_c_224_n 0.0164251f $X=2.415 $Y=1.48 $X2=0 $Y2=0
cc_140 N_A_c_170_n N_A_340_93#_c_224_n 0.00126496f $X=2.475 $Y=1.48 $X2=0 $Y2=0
cc_141 N_A_M1012_g N_A_340_93#_c_247_n 5.07822e-19 $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_142 N_A_c_172_n N_A_340_93#_c_247_n 0.0176589f $X=2.415 $Y=1.48 $X2=0 $Y2=0
cc_143 N_A_c_170_n N_A_340_93#_c_247_n 0.00160203f $X=2.475 $Y=1.48 $X2=0 $Y2=0
cc_144 N_A_M1002_g N_A_340_93#_c_218_n 0.0076551f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_145 N_A_M1012_g N_A_340_93#_c_218_n 0.00221179f $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_146 N_A_c_172_n N_A_340_93#_c_219_n 0.00329809f $X=2.415 $Y=1.48 $X2=0 $Y2=0
cc_147 N_A_c_170_n N_A_340_93#_c_219_n 0.0161683f $X=2.475 $Y=1.48 $X2=0 $Y2=0
cc_148 N_A_M1013_g N_VPWR_c_290_n 0.00432655f $X=1.985 $Y=2.655 $X2=0 $Y2=0
cc_149 N_A_M1013_g N_VPWR_c_292_n 0.00510437f $X=1.985 $Y=2.655 $X2=0 $Y2=0
cc_150 N_A_M1013_g N_VPWR_c_288_n 0.00515964f $X=1.985 $Y=2.655 $X2=0 $Y2=0
cc_151 N_A_M1002_g N_KAGND_c_345_n 0.00138219f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_152 N_A_M1012_g N_KAGND_c_345_n 0.00812645f $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_KAGND_c_346_n 0.00331496f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_154 N_A_M1012_g N_KAGND_c_346_n 0.0033271f $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_VGND_c_398_n 0.00310524f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_156 N_A_M1012_g N_VGND_c_398_n 0.00310524f $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_157 N_A_M1002_g N_VGND_c_399_n 0.0048834f $X=2.115 $Y=0.675 $X2=0 $Y2=0
cc_158 N_A_M1012_g N_VGND_c_399_n 0.0048834f $X=2.475 $Y=0.675 $X2=0 $Y2=0
cc_159 N_A_340_93#_c_223_n N_VPWR_M1008_s 0.0109378f $X=2.895 $Y=2.04 $X2=0
+ $Y2=0
cc_160 N_A_340_93#_c_222_n N_VPWR_c_289_n 4.76441e-19 $X=2.2 $Y=2.695 $X2=0
+ $Y2=0
cc_161 N_A_340_93#_M1008_g N_VPWR_c_290_n 0.0255081f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_340_93#_M1010_g N_VPWR_c_290_n 0.00358067f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_340_93#_c_222_n N_VPWR_c_290_n 0.0391837f $X=2.2 $Y=2.695 $X2=0 $Y2=0
cc_164 N_A_340_93#_c_223_n N_VPWR_c_290_n 0.0264831f $X=2.895 $Y=2.04 $X2=0
+ $Y2=0
cc_165 N_A_340_93#_c_222_n N_VPWR_c_292_n 0.00660276f $X=2.2 $Y=2.695 $X2=0
+ $Y2=0
cc_166 N_A_340_93#_M1008_g N_VPWR_c_293_n 0.00388479f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_340_93#_M1010_g N_VPWR_c_293_n 0.00585385f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_340_93#_M1008_g N_VPWR_c_288_n 0.006597f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_340_93#_M1010_g N_VPWR_c_288_n 0.0116546f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_340_93#_c_222_n N_VPWR_c_288_n 0.00720343f $X=2.2 $Y=2.695 $X2=0
+ $Y2=0
cc_171 N_A_340_93#_c_223_n A_602_367# 0.00433061f $X=2.895 $Y=2.04 $X2=-0.22
+ $Y2=-0.245
cc_172 N_A_340_93#_c_214_n N_X_c_330_n 0.0343639f $X=3.295 $Y=1.005 $X2=0 $Y2=0
cc_173 N_A_340_93#_c_268_p N_X_c_330_n 0.0143575f $X=3.06 $Y=1.225 $X2=0 $Y2=0
cc_174 N_A_340_93#_c_247_n N_X_c_330_n 0.0529514f $X=3.06 $Y=1.955 $X2=0 $Y2=0
cc_175 N_A_340_93#_c_218_n N_KAGND_c_344_n 0.00790417f $X=1.9 $Y=0.715 $X2=0
+ $Y2=0
cc_176 N_A_340_93#_c_213_n N_KAGND_c_345_n 0.0139281f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_177 N_A_340_93#_c_214_n N_KAGND_c_345_n 0.00392337f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_178 N_A_340_93#_c_216_n N_KAGND_c_345_n 0.0228171f $X=2.895 $Y=1.14 $X2=0
+ $Y2=0
cc_179 N_A_340_93#_c_268_p N_KAGND_c_345_n 0.0181069f $X=3.06 $Y=1.225 $X2=0
+ $Y2=0
cc_180 N_A_340_93#_c_218_n N_KAGND_c_345_n 0.0120821f $X=1.9 $Y=0.715 $X2=0
+ $Y2=0
cc_181 N_A_340_93#_c_219_n N_KAGND_c_345_n 8.4817e-19 $X=3.06 $Y=1.17 $X2=0
+ $Y2=0
cc_182 N_A_340_93#_M1007_d N_KAGND_c_346_n 0.00135548f $X=1.7 $Y=0.465 $X2=0
+ $Y2=0
cc_183 N_A_340_93#_c_214_n N_KAGND_c_346_n 0.00943673f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_184 N_A_340_93#_c_216_n N_KAGND_c_346_n 0.0176818f $X=2.895 $Y=1.14 $X2=0
+ $Y2=0
cc_185 N_A_340_93#_c_268_p N_KAGND_c_346_n 0.00411381f $X=3.06 $Y=1.225 $X2=0
+ $Y2=0
cc_186 N_A_340_93#_c_218_n N_KAGND_c_346_n 0.0342136f $X=1.9 $Y=0.715 $X2=0
+ $Y2=0
cc_187 N_A_340_93#_c_213_n N_VGND_c_398_n 0.00310524f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_188 N_A_340_93#_c_214_n N_VGND_c_398_n 0.00310524f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_189 N_A_340_93#_c_218_n N_VGND_c_398_n 0.00350771f $X=1.9 $Y=0.715 $X2=0
+ $Y2=0
cc_190 N_A_340_93#_c_213_n N_VGND_c_399_n 0.00372327f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_191 N_A_340_93#_c_214_n N_VGND_c_399_n 0.00510437f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_192 N_A_340_93#_c_218_n N_VGND_c_399_n 0.0108653f $X=1.9 $Y=0.715 $X2=0 $Y2=0
cc_193 N_VPWR_c_288_n A_602_367# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.22 $Y2=-0.245
cc_194 N_VPWR_c_288_n N_X_M1010_d 0.00302127f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_293_n N_X_c_330_n 0.0242556f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_288_n N_X_c_330_n 0.0139182f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_X_c_330_n N_KAGND_c_345_n 0.0150658f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_198 N_X_M1005_d N_KAGND_c_346_n 9.16941e-19 $X=3.37 $Y=0.465 $X2=0 $Y2=0
cc_199 N_X_c_330_n N_KAGND_c_346_n 0.0370046f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_200 N_X_c_330_n N_VGND_c_398_n 0.00165179f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_201 N_X_c_330_n N_VGND_c_399_n 0.0109076f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_202 A_110_93# N_KAGND_c_346_n 0.00255809f $X=0.55 $Y=0.465 $X2=3.02 $Y2=0.555
cc_203 N_KAGND_c_344_n A_268_93# 0.00150499f $X=1.38 $Y=0.555 $X2=-0.22
+ $Y2=-0.245
cc_204 N_KAGND_c_346_n A_268_93# 0.00135548f $X=3.02 $Y=0.555 $X2=-0.22
+ $Y2=-0.245
cc_205 N_KAGND_c_346_n A_438_93# 0.00225912f $X=3.02 $Y=0.555 $X2=-0.22
+ $Y2=-0.245
cc_206 N_KAGND_c_345_n A_602_93# 0.00431788f $X=3.02 $Y=0.555 $X2=-0.22
+ $Y2=-0.245
cc_207 N_KAGND_c_346_n A_602_93# 7.09126e-19 $X=3.02 $Y=0.555 $X2=-0.22
+ $Y2=-0.245
cc_208 N_KAGND_c_344_n N_VGND_c_398_n 0.00640001f $X=1.38 $Y=0.555 $X2=0 $Y2=0
cc_209 N_KAGND_c_345_n N_VGND_c_398_n 0.00640001f $X=3.02 $Y=0.555 $X2=0 $Y2=0
cc_210 N_KAGND_c_346_n N_VGND_c_398_n 0.337693f $X=3.02 $Y=0.555 $X2=0 $Y2=0
cc_211 N_KAGND_c_344_n N_VGND_c_399_n 0.0201323f $X=1.38 $Y=0.555 $X2=0 $Y2=0
cc_212 N_KAGND_c_345_n N_VGND_c_399_n 0.0201323f $X=3.02 $Y=0.555 $X2=0 $Y2=0
cc_213 N_KAGND_c_346_n N_VGND_c_399_n 0.0106921f $X=3.02 $Y=0.555 $X2=0 $Y2=0
