# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.500000 1.175000 1.775000 1.505000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.345000 0.285000 6.635000 3.075000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.295000 2.285000 0.640000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.720000  0.085000 0.945000 1.005000 ;
        RECT 2.825000  0.085000 3.155000 0.485000 ;
        RECT 4.800000  0.085000 5.110000 1.085000 ;
        RECT 5.865000  0.085000 6.175000 1.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.720000 3.415000 ;
        RECT 0.720000 2.385000 0.980000 3.245000 ;
        RECT 2.440000 2.715000 2.700000 3.245000 ;
        RECT 4.450000 2.450000 5.190000 3.245000 ;
        RECT 4.950000 2.305000 5.190000 2.450000 ;
        RECT 5.865000 1.815000 6.175000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.150000 0.675000 0.550000 1.005000 ;
      RECT 0.150000 1.005000 0.330000 1.675000 ;
      RECT 0.150000 1.675000 2.890000 1.865000 ;
      RECT 0.150000 1.865000 0.550000 3.065000 ;
      RECT 1.115000 0.810000 2.275000 0.995000 ;
      RECT 1.115000 0.995000 3.920000 1.005000 ;
      RECT 1.150000 2.385000 1.445000 2.905000 ;
      RECT 1.150000 2.905000 2.270000 3.075000 ;
      RECT 1.730000 2.035000 3.460000 2.205000 ;
      RECT 1.730000 2.205000 1.930000 2.735000 ;
      RECT 1.945000 1.005000 3.920000 1.165000 ;
      RECT 1.945000 1.165000 2.275000 1.505000 ;
      RECT 2.100000 2.375000 3.920000 2.545000 ;
      RECT 2.100000 2.545000 2.270000 2.905000 ;
      RECT 2.455000 0.295000 2.645000 0.655000 ;
      RECT 2.455000 0.655000 4.290000 0.825000 ;
      RECT 2.560000 1.335000 2.890000 1.675000 ;
      RECT 3.130000 1.535000 3.460000 2.035000 ;
      RECT 3.255000 2.715000 4.280000 3.065000 ;
      RECT 3.490000 1.165000 3.920000 1.245000 ;
      RECT 3.670000 1.245000 3.920000 2.375000 ;
      RECT 3.725000 0.275000 4.630000 0.465000 ;
      RECT 4.090000 0.825000 4.290000 1.435000 ;
      RECT 4.090000 1.615000 5.210000 1.785000 ;
      RECT 4.090000 1.785000 4.280000 2.715000 ;
      RECT 4.450000 1.955000 4.780000 1.965000 ;
      RECT 4.450000 1.965000 5.660000 2.135000 ;
      RECT 4.450000 2.135000 4.780000 2.215000 ;
      RECT 4.460000 0.465000 4.630000 1.255000 ;
      RECT 4.460000 1.255000 5.210000 1.615000 ;
      RECT 5.280000 0.255000 5.560000 1.075000 ;
      RECT 5.360000 2.135000 5.660000 3.025000 ;
      RECT 5.390000 1.075000 5.560000 1.255000 ;
      RECT 5.390000 1.255000 6.175000 1.585000 ;
      RECT 5.390000 1.585000 5.660000 1.965000 ;
  END
END sky130_fd_sc_lp__dlxtn_1
