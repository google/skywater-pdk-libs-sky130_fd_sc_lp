* File: sky130_fd_sc_lp__mux2i_lp.pex.spice
* Created: Fri Aug 28 10:45:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2I_LP%S 2 3 4 7 11 13 15 18 22 24 26 29 32 33 34
+ 36 38 39 40 41 50 51
r114 51 52 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=2.835 $Y=0.94
+ $X2=2.86 $Y2=0.94
r115 49 51 41.2928 $w=3.21e-07 $l=2.75e-07 $layer=POLY_cond $X=2.56 $Y=0.94
+ $X2=2.835 $Y2=0.94
r116 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=0.94 $X2=2.56 $Y2=0.94
r117 47 49 12.7632 $w=3.21e-07 $l=8.5e-08 $layer=POLY_cond $X=2.475 $Y=0.94
+ $X2=2.56 $Y2=0.94
r118 46 47 0.750779 $w=3.21e-07 $l=5e-09 $layer=POLY_cond $X=2.47 $Y=0.94
+ $X2=2.475 $Y2=0.94
r119 41 50 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.16 $Y=0.94 $X2=2.56
+ $Y2=0.94
r120 40 41 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.89 $Y=0.94
+ $X2=2.16 $Y2=0.94
r121 39 45 88.0219 $w=4.65e-07 $l=5.05e-07 $layer=POLY_cond $X=0.337 $Y=0.98
+ $X2=0.337 $Y2=1.485
r122 39 44 47.3569 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.337 $Y=0.98
+ $X2=0.337 $Y2=0.815
r123 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=0.98 $X2=0.27 $Y2=0.98
r124 36 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.805 $Y=0.775
+ $X2=1.89 $Y2=0.94
r125 35 36 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.805 $Y=0.425
+ $X2=1.805 $Y2=0.775
r126 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=0.34
+ $X2=1.805 $Y2=0.425
r127 33 34 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.72 $Y=0.34 $X2=0.785
+ $Y2=0.34
r128 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=0.425
+ $X2=0.785 $Y2=0.34
r129 31 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.7 $Y=0.425
+ $X2=0.7 $Y2=0.815
r130 30 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=0.9
+ $X2=0.27 $Y2=0.9
r131 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.615 $Y=0.9
+ $X2=0.7 $Y2=0.815
r132 29 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.615 $Y=0.9
+ $X2=0.435 $Y2=0.9
r133 24 52 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.86 $Y=0.775
+ $X2=2.86 $Y2=0.94
r134 24 26 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.86 $Y=0.775
+ $X2=2.86 $Y2=0.455
r135 20 51 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.105
+ $X2=2.835 $Y2=0.94
r136 20 22 892.213 $w=1.5e-07 $l=1.74e-06 $layer=POLY_cond $X=2.835 $Y=1.105
+ $X2=2.835 $Y2=2.845
r137 16 47 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.475 $Y=1.105
+ $X2=2.475 $Y2=0.94
r138 16 18 892.213 $w=1.5e-07 $l=1.74e-06 $layer=POLY_cond $X=2.475 $Y=1.105
+ $X2=2.475 $Y2=2.845
r139 13 46 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=0.775
+ $X2=2.47 $Y2=0.94
r140 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.47 $Y=0.775
+ $X2=2.47 $Y2=0.455
r141 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.55 $Y=2.445 $X2=0.55
+ $Y2=2.845
r142 7 44 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=0.495 $Y=0.455
+ $X2=0.495 $Y2=0.815
r143 3 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=2.37
+ $X2=0.55 $Y2=2.445
r144 3 4 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.475 $Y=2.37
+ $X2=0.255 $Y2=2.37
r145 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=2.295
+ $X2=0.255 $Y2=2.37
r146 2 45 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.18 $Y=2.295
+ $X2=0.18 $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP%A1 3 7 10 11 15 16 18 21
c68 16 0 2.19138e-19 $X=1.42 $Y=2.28
r69 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.32
+ $X2=0.975 $Y2=1.155
r70 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.32 $X2=0.975 $Y2=1.32
r71 18 22 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.72 $Y=1.32
+ $X2=0.975 $Y2=1.32
r72 16 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=2.28
+ $X2=1.42 $Y2=2.445
r73 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=2.28 $X2=1.42 $Y2=2.28
r74 12 15 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.12 $Y=2.28 $X2=1.42
+ $Y2=2.28
r75 11 22 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.035 $Y=1.32
+ $X2=0.975 $Y2=1.32
r76 10 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=2.115
+ $X2=1.12 $Y2=2.28
r77 9 11 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.12 $Y=1.485
+ $X2=1.035 $Y2=1.32
r78 9 10 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.12 $Y=1.485
+ $X2=1.12 $Y2=2.115
r79 7 27 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.37 $Y=2.845 $X2=1.37
+ $Y2=2.445
r80 3 23 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.885 $Y=0.455
+ $X2=0.885 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP%A0 3 5 8 11 14 15 16 24
c58 16 0 2.27745e-20 $X=0.72 $Y=2.035
c59 3 0 2.10122e-20 $X=0.94 $Y=2.845
r60 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.94 $Y=1.89
+ $X2=1.015 $Y2=1.89
r61 20 23 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.7 $Y=1.89 $X2=0.94
+ $Y2=1.89
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.89 $X2=0.7 $Y2=1.89
r63 16 21 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=0.72 $Y=1.937 $X2=0.7
+ $Y2=1.937
r64 15 21 12.4735 $w=4.23e-07 $l=4.6e-07 $layer=LI1_cond $X=0.24 $Y=1.937
+ $X2=0.7 $Y2=1.937
r65 13 14 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.527 $Y=0.885
+ $X2=1.527 $Y2=1.035
r66 11 13 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.545 $Y=0.455
+ $X2=1.545 $Y2=0.885
r67 8 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.51 $Y=1.725
+ $X2=1.51 $Y2=1.035
r68 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.435 $Y=1.8
+ $X2=1.51 $Y2=1.725
r69 5 24 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.435 $Y=1.8
+ $X2=1.015 $Y2=1.8
r70 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=2.055
+ $X2=0.94 $Y2=1.89
r71 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.94 $Y=2.055 $X2=0.94
+ $Y2=2.845
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP%A_365_255# 1 2 9 13 15 18 22 26 28
r65 24 28 5.00808 $w=3.42e-07 $l=1.71377e-07 $layer=LI1_cond $X=3.075 $Y=1.275
+ $X2=3.062 $Y2=1.44
r66 24 26 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=3.075 $Y=1.275
+ $X2=3.075 $Y2=0.47
r67 20 28 5.00808 $w=3.42e-07 $l=1.65e-07 $layer=LI1_cond $X=3.062 $Y=1.605
+ $X2=3.062 $Y2=1.44
r68 20 22 40.2543 $w=3.53e-07 $l=1.24e-06 $layer=LI1_cond $X=3.062 $Y=1.605
+ $X2=3.062 $Y2=2.845
r69 18 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.44
+ $X2=1.99 $Y2=1.605
r70 18 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.44
+ $X2=1.99 $Y2=1.275
r71 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.44 $X2=1.99 $Y2=1.44
r72 15 28 1.47678 $w=3.3e-07 $l=1.77e-07 $layer=LI1_cond $X=2.885 $Y=1.44
+ $X2=3.062 $Y2=1.44
r73 15 17 31.2557 $w=3.28e-07 $l=8.95e-07 $layer=LI1_cond $X=2.885 $Y=1.44
+ $X2=1.99 $Y2=1.44
r74 13 30 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.935 $Y=0.455
+ $X2=1.935 $Y2=1.275
r75 9 31 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=1.9 $Y=2.845 $X2=1.9
+ $Y2=1.605
r76 2 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=2.635 $X2=3.05 $Y2=2.845
r77 1 26 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.935
+ $Y=0.245 $X2=3.075 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP%VPWR 1 2 7 9 13 15 17 24 25 31
r39 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.26 $Y2=3.33
r44 22 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 18 28 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=3.33 $X2=0.25
+ $Y2=3.33
r48 18 20 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=3.33 $X2=0.72
+ $Y2=3.33
r49 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.26 $Y2=3.33
r50 17 20 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 15 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=3.245
+ $X2=2.26 $Y2=3.33
r54 11 13 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.26 $Y=3.245
+ $X2=2.26 $Y2=2.89
r55 7 28 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.25 $Y2=3.33
r56 7 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.335 $Y=3.245 $X2=0.335
+ $Y2=2.845
r57 2 13 600 $w=1.7e-07 $l=3.92301e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=2.635 $X2=2.26 $Y2=2.89
r58 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=2.635 $X2=0.335 $Y2=2.845
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP%Y 1 2 7 10 11 12 13 21 24 25 34
c77 11 0 1.96363e-19 $X=1.755 $Y=1.86
c78 7 0 2.10122e-20 $X=1.755 $Y=2.7
r79 29 34 2.06799 $w=5.2e-07 $l=5e-08 $layer=LI1_cond $X=2.015 $Y=2.355
+ $X2=2.015 $Y2=2.405
r80 25 34 0.544357 $w=3.81e-07 $l=1.7e-08 $layer=LI1_cond $X=2.015 $Y=2.422
+ $X2=2.015 $Y2=2.405
r81 25 29 0.414027 $w=5.18e-07 $l=1.8e-08 $layer=LI1_cond $X=2.015 $Y=2.337
+ $X2=2.015 $Y2=2.355
r82 24 25 6.94646 $w=5.18e-07 $l=3.02e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=2.015 $Y2=2.337
r83 23 24 2.07014 $w=5.18e-07 $l=9e-08 $layer=LI1_cond $X=2.015 $Y=1.945
+ $X2=2.015 $Y2=2.035
r84 19 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.215 $Y=0.76
+ $X2=1.465 $Y2=0.76
r85 13 16 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.155 $Y=2.7
+ $X2=1.155 $Y2=2.845
r86 11 23 9.39785 $w=1.7e-07 $l=2.995e-07 $layer=LI1_cond $X=1.755 $Y=1.86
+ $X2=2.015 $Y2=1.945
r87 11 12 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.755 $Y=1.86
+ $X2=1.55 $Y2=1.86
r88 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.465 $Y=1.775
+ $X2=1.55 $Y2=1.86
r89 9 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0.925
+ $X2=1.465 $Y2=0.76
r90 9 10 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.465 $Y=0.925
+ $X2=1.465 $Y2=1.775
r91 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=2.7 $X2=1.155
+ $Y2=2.7
r92 7 25 8.90184 $w=3.81e-07 $l=3.86735e-07 $layer=LI1_cond $X=1.755 $Y=2.7
+ $X2=2.015 $Y2=2.422
r93 7 8 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.755 $Y=2.7 $X2=1.32
+ $Y2=2.7
r94 2 16 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=2.635 $X2=1.155 $Y2=2.845
r95 1 19 182 $w=1.7e-07 $l=6.29722e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.245 $X2=1.215 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP%VGND 1 2 7 9 13 15 17 27 28 34
r43 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 28 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r46 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.225
+ $Y2=0
r48 25 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=3.12
+ $Y2=0
r49 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r50 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r51 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 18 31 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r53 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r54 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=2.225
+ $Y2=0
r55 17 23 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=1.68
+ $Y2=0
r56 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r57 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r58 15 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0
r60 11 13 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0.415
r61 7 31 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r62 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.435
r63 2 13 182 $w=1.7e-07 $l=2.87706e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.245 $X2=2.225 $Y2=0.415
r64 1 9 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.245 $X2=0.28 $Y2=0.435
.ends

