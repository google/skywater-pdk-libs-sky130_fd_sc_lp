* File: sky130_fd_sc_lp__or4b_m.pxi.spice
* Created: Fri Aug 28 11:26:15 2020
* 
x_PM_SKY130_FD_SC_LP__OR4B_M%D_N N_D_N_c_80_n N_D_N_M1003_g N_D_N_M1004_g
+ N_D_N_c_82_n D_N D_N N_D_N_c_78_n N_D_N_c_79_n PM_SKY130_FD_SC_LP__OR4B_M%D_N
x_PM_SKY130_FD_SC_LP__OR4B_M%A_38_125# N_A_38_125#_M1003_s N_A_38_125#_M1004_s
+ N_A_38_125#_M1005_g N_A_38_125#_c_118_n N_A_38_125#_c_119_n
+ N_A_38_125#_M1000_g N_A_38_125#_c_111_n N_A_38_125#_c_112_n
+ N_A_38_125#_c_113_n N_A_38_125#_c_122_n N_A_38_125#_c_123_n
+ N_A_38_125#_c_124_n N_A_38_125#_c_114_n N_A_38_125#_c_115_n
+ N_A_38_125#_c_116_n N_A_38_125#_c_125_n N_A_38_125#_c_117_n
+ PM_SKY130_FD_SC_LP__OR4B_M%A_38_125#
x_PM_SKY130_FD_SC_LP__OR4B_M%C N_C_c_180_n N_C_M1006_g N_C_c_181_n N_C_c_182_n
+ N_C_M1008_g C C C N_C_c_186_n PM_SKY130_FD_SC_LP__OR4B_M%C
x_PM_SKY130_FD_SC_LP__OR4B_M%B N_B_M1002_g N_B_M1009_g B B N_B_c_226_n
+ PM_SKY130_FD_SC_LP__OR4B_M%B
x_PM_SKY130_FD_SC_LP__OR4B_M%A N_A_M1010_g N_A_M1011_g A A A A N_A_c_254_n
+ PM_SKY130_FD_SC_LP__OR4B_M%A
x_PM_SKY130_FD_SC_LP__OR4B_M%A_215_125# N_A_215_125#_M1005_d
+ N_A_215_125#_M1002_d N_A_215_125#_M1000_s N_A_215_125#_c_296_n
+ N_A_215_125#_M1001_g N_A_215_125#_M1007_g N_A_215_125#_c_299_n
+ N_A_215_125#_c_292_n N_A_215_125#_c_293_n N_A_215_125#_c_294_n
+ N_A_215_125#_c_313_n N_A_215_125#_c_332_n N_A_215_125#_c_301_n
+ N_A_215_125#_c_315_n N_A_215_125#_c_295_n N_A_215_125#_c_302_n
+ N_A_215_125#_c_303_n PM_SKY130_FD_SC_LP__OR4B_M%A_215_125#
x_PM_SKY130_FD_SC_LP__OR4B_M%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_c_399_n
+ N_VPWR_c_400_n N_VPWR_c_421_n N_VPWR_c_401_n N_VPWR_c_402_n VPWR
+ N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_398_n N_VPWR_c_406_n
+ PM_SKY130_FD_SC_LP__OR4B_M%VPWR
x_PM_SKY130_FD_SC_LP__OR4B_M%X N_X_M1007_d N_X_M1001_d X X X X X X X X
+ PM_SKY130_FD_SC_LP__OR4B_M%X
x_PM_SKY130_FD_SC_LP__OR4B_M%VGND N_VGND_M1003_d N_VGND_M1006_d N_VGND_M1011_d
+ N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n
+ VGND N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n
+ N_VGND_c_472_n PM_SKY130_FD_SC_LP__OR4B_M%VGND
cc_1 VNB N_D_N_M1003_g 0.045172f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.835
cc_2 VNB N_D_N_c_78_n 0.0209029f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_3 VNB N_D_N_c_79_n 0.00897674f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_4 VNB N_A_38_125#_c_111_n 0.0177845f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_5 VNB N_A_38_125#_c_112_n 0.0228909f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_6 VNB N_A_38_125#_c_113_n 0.0150538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_38_125#_c_114_n 0.018664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_38_125#_c_115_n 0.00304611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_38_125#_c_116_n 0.0152645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_38_125#_c_117_n 2.20898e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_c_180_n 0.0204214f $X=-0.19 $Y=-0.245 $X2=0.412 $Y2=1.682
cc_12 VNB N_C_c_181_n 0.0414698f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.835
cc_13 VNB N_C_c_182_n 0.00637224f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.835
cc_14 VNB N_C_M1008_g 0.020077f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.73
cc_15 VNB N_B_M1002_g 0.0364999f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.49
cc_16 VNB B 0.0085f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.73
cc_17 VNB N_B_c_226_n 0.0469572f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_A_M1011_g 0.0343381f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.16
cc_19 VNB A 0.0114287f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB N_A_c_254_n 0.0166046f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_21 VNB N_A_215_125#_M1007_g 0.0467561f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_22 VNB N_A_215_125#_c_292_n 0.00141675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_215_125#_c_293_n 0.00445248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_215_125#_c_294_n 0.0123635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_215_125#_c_295_n 0.00102738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_398_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0633268f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.16
cc_28 VNB N_VGND_c_463_n 0.0282592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_464_n 0.0212377f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.655
cc_30 VNB N_VGND_c_465_n 0.0200255f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.665
cc_31 VNB N_VGND_c_466_n 0.0289556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_467_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_468_n 0.0217182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_469_n 0.0233753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_470_n 0.264058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_471_n 0.0271851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_472_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_D_N_c_80_n 0.0253966f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=1.968
cc_39 VPB N_D_N_M1004_g 0.044193f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.73
cc_40 VPB N_D_N_c_82_n 0.0245287f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=2.16
cc_41 VPB N_D_N_c_78_n 0.00232285f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.655
cc_42 VPB N_D_N_c_79_n 0.0232509f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.655
cc_43 VPB N_A_38_125#_c_118_n 0.0374002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_38_125#_c_119_n 0.0183314f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=2.16
cc_45 VPB N_A_38_125#_M1000_g 0.0228091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_38_125#_c_112_n 0.00130279f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.655
cc_47 VPB N_A_38_125#_c_122_n 4.08405e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_38_125#_c_123_n 0.0117264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_38_125#_c_124_n 0.00844209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_38_125#_c_125_n 0.0115888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_38_125#_c_117_n 0.0106219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_C_M1008_g 0.0416861f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.73
cc_53 VPB C 0.0316906f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_54 VPB N_C_c_186_n 0.0453368f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.655
cc_55 VPB N_B_M1002_g 0.027495f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.49
cc_56 VPB N_A_M1010_g 0.0176383f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.49
cc_57 VPB A 0.00961775f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_58 VPB N_A_c_254_n 0.0171819f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.655
cc_59 VPB N_A_215_125#_c_296_n 0.0366734f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_215_125#_M1001_g 0.029343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_215_125#_M1007_g 0.00333657f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.655
cc_62 VPB N_A_215_125#_c_299_n 0.0102663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_215_125#_c_293_n 0.00804418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_215_125#_c_301_n 0.00592732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_215_125#_c_302_n 0.00225151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_215_125#_c_303_n 0.0434158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_399_n 0.0135676f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.73
cc_68 VPB N_VPWR_c_400_n 0.0155423f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_69 VPB N_VPWR_c_401_n 0.0538491f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=1.49
cc_70 VPB N_VPWR_c_402_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.655
cc_71 VPB N_VPWR_c_403_n 0.0194802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_404_n 0.0215374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_398_n 0.0866132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_406_n 0.00628367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB X 0.0154271f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.16
cc_76 VPB X 0.0511648f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=2.16
cc_77 N_D_N_c_80_n N_A_38_125#_c_119_n 0.0137845f $X=0.412 $Y=1.968 $X2=0 $Y2=0
cc_78 N_D_N_M1003_g N_A_38_125#_c_111_n 0.0106134f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_79 N_D_N_c_78_n N_A_38_125#_c_112_n 0.0137845f $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_80 N_D_N_c_79_n N_A_38_125#_c_112_n 2.53578e-19 $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_81 N_D_N_M1003_g N_A_38_125#_c_113_n 0.00781288f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_82 N_D_N_M1004_g N_A_38_125#_c_122_n 3.52891e-19 $X=0.53 $Y=2.73 $X2=0 $Y2=0
cc_83 N_D_N_M1004_g N_A_38_125#_c_123_n 0.01813f $X=0.53 $Y=2.73 $X2=0 $Y2=0
cc_84 N_D_N_c_82_n N_A_38_125#_c_123_n 3.7612e-19 $X=0.412 $Y=2.16 $X2=0 $Y2=0
cc_85 N_D_N_c_79_n N_A_38_125#_c_123_n 0.00518419f $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_86 N_D_N_c_82_n N_A_38_125#_c_124_n 0.00135198f $X=0.412 $Y=2.16 $X2=0 $Y2=0
cc_87 N_D_N_c_79_n N_A_38_125#_c_124_n 0.0158411f $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_88 N_D_N_M1003_g N_A_38_125#_c_114_n 0.019066f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_89 N_D_N_c_78_n N_A_38_125#_c_114_n 0.0016167f $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_90 N_D_N_c_79_n N_A_38_125#_c_114_n 0.0241613f $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_91 N_D_N_M1003_g N_A_38_125#_c_115_n 0.00787729f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_92 N_D_N_c_79_n N_A_38_125#_c_115_n 0.0496577f $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_93 N_D_N_M1003_g N_A_38_125#_c_116_n 0.0137845f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_94 N_D_N_c_82_n N_A_38_125#_c_125_n 0.00787729f $X=0.412 $Y=2.16 $X2=0 $Y2=0
cc_95 N_D_N_c_78_n N_A_38_125#_c_117_n 0.00787729f $X=0.385 $Y=1.655 $X2=0 $Y2=0
cc_96 N_D_N_M1004_g C 8.38678e-19 $X=0.53 $Y=2.73 $X2=0 $Y2=0
cc_97 N_D_N_M1004_g N_VPWR_c_399_n 0.015388f $X=0.53 $Y=2.73 $X2=0 $Y2=0
cc_98 N_D_N_M1004_g N_VPWR_c_403_n 0.00468165f $X=0.53 $Y=2.73 $X2=0 $Y2=0
cc_99 N_D_N_M1004_g N_VPWR_c_398_n 0.00453141f $X=0.53 $Y=2.73 $X2=0 $Y2=0
cc_100 N_D_N_M1003_g N_VGND_c_463_n 0.0032771f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_101 N_D_N_M1003_g N_VGND_c_470_n 0.00469432f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_102 N_D_N_M1003_g N_VGND_c_471_n 0.00415323f $X=0.53 $Y=0.835 $X2=0 $Y2=0
cc_103 N_A_38_125#_c_111_n N_C_c_180_n 0.0113899f $X=0.98 $Y=1.155 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_38_125#_c_118_n N_C_c_182_n 0.0101358f $X=1.54 $Y=1.75 $X2=0 $Y2=0
cc_105 N_A_38_125#_c_116_n N_C_c_182_n 0.00933311f $X=0.98 $Y=1.32 $X2=0 $Y2=0
cc_106 N_A_38_125#_c_118_n N_C_M1008_g 0.0559316f $X=1.54 $Y=1.75 $X2=0 $Y2=0
cc_107 N_A_38_125#_M1000_g C 0.00445046f $X=1.615 $Y=2.195 $X2=0 $Y2=0
cc_108 N_A_38_125#_c_118_n A 0.00482268f $X=1.54 $Y=1.75 $X2=0 $Y2=0
cc_109 N_A_38_125#_c_111_n N_A_215_125#_c_292_n 0.00353471f $X=0.98 $Y=1.155
+ $X2=0 $Y2=0
cc_110 N_A_38_125#_c_114_n N_A_215_125#_c_292_n 0.00635016f $X=0.857 $Y=1.31
+ $X2=0 $Y2=0
cc_111 N_A_38_125#_c_116_n N_A_215_125#_c_292_n 4.31144e-19 $X=0.98 $Y=1.32
+ $X2=0 $Y2=0
cc_112 N_A_38_125#_c_118_n N_A_215_125#_c_293_n 0.0139379f $X=1.54 $Y=1.75 $X2=0
+ $Y2=0
cc_113 N_A_38_125#_M1000_g N_A_215_125#_c_293_n 0.00608003f $X=1.615 $Y=2.195
+ $X2=0 $Y2=0
cc_114 N_A_38_125#_c_112_n N_A_215_125#_c_293_n 0.00683278f $X=0.98 $Y=1.675
+ $X2=0 $Y2=0
cc_115 N_A_38_125#_c_115_n N_A_215_125#_c_293_n 0.030826f $X=0.98 $Y=1.32 $X2=0
+ $Y2=0
cc_116 N_A_38_125#_c_125_n N_A_215_125#_c_293_n 0.0219192f $X=0.735 $Y=2.34
+ $X2=0 $Y2=0
cc_117 N_A_38_125#_c_118_n N_A_215_125#_c_294_n 0.00193003f $X=1.54 $Y=1.75
+ $X2=0 $Y2=0
cc_118 N_A_38_125#_c_118_n N_A_215_125#_c_313_n 0.00258034f $X=1.54 $Y=1.75
+ $X2=0 $Y2=0
cc_119 N_A_38_125#_M1000_g N_A_215_125#_c_313_n 0.0126675f $X=1.615 $Y=2.195
+ $X2=0 $Y2=0
cc_120 N_A_38_125#_c_111_n N_A_215_125#_c_315_n 0.00349634f $X=0.98 $Y=1.155
+ $X2=0 $Y2=0
cc_121 N_A_38_125#_c_113_n N_A_215_125#_c_315_n 6.7135e-19 $X=0.315 $Y=0.9 $X2=0
+ $Y2=0
cc_122 N_A_38_125#_c_114_n N_A_215_125#_c_315_n 9.87196e-19 $X=0.857 $Y=1.31
+ $X2=0 $Y2=0
cc_123 N_A_38_125#_c_116_n N_A_215_125#_c_315_n 0.00185023f $X=0.98 $Y=1.32
+ $X2=0 $Y2=0
cc_124 N_A_38_125#_c_114_n N_A_215_125#_c_295_n 0.00716961f $X=0.857 $Y=1.31
+ $X2=0 $Y2=0
cc_125 N_A_38_125#_c_115_n N_A_215_125#_c_295_n 0.00693738f $X=0.98 $Y=1.32
+ $X2=0 $Y2=0
cc_126 N_A_38_125#_c_116_n N_A_215_125#_c_295_n 0.00287912f $X=0.98 $Y=1.32
+ $X2=0 $Y2=0
cc_127 N_A_38_125#_c_123_n N_VPWR_c_399_n 0.0171134f $X=0.65 $Y=2.425 $X2=0
+ $Y2=0
cc_128 N_A_38_125#_c_122_n N_VPWR_c_403_n 0.00488264f $X=0.315 $Y=2.665 $X2=0
+ $Y2=0
cc_129 N_A_38_125#_c_122_n N_VPWR_c_398_n 0.00619834f $X=0.315 $Y=2.665 $X2=0
+ $Y2=0
cc_130 N_A_38_125#_c_123_n N_VPWR_c_398_n 0.00679911f $X=0.65 $Y=2.425 $X2=0
+ $Y2=0
cc_131 N_A_38_125#_c_111_n N_VGND_c_463_n 0.0032771f $X=0.98 $Y=1.155 $X2=0
+ $Y2=0
cc_132 N_A_38_125#_c_114_n N_VGND_c_463_n 0.0149335f $X=0.857 $Y=1.31 $X2=0
+ $Y2=0
cc_133 N_A_38_125#_c_116_n N_VGND_c_463_n 3.95657e-19 $X=0.98 $Y=1.32 $X2=0
+ $Y2=0
cc_134 N_A_38_125#_c_111_n N_VGND_c_468_n 0.00400711f $X=0.98 $Y=1.155 $X2=0
+ $Y2=0
cc_135 N_A_38_125#_c_111_n N_VGND_c_470_n 0.00469432f $X=0.98 $Y=1.155 $X2=0
+ $Y2=0
cc_136 N_A_38_125#_c_113_n N_VGND_c_470_n 0.0124764f $X=0.315 $Y=0.9 $X2=0 $Y2=0
cc_137 N_C_c_181_n N_B_M1002_g 0.0894236f $X=1.9 $Y=1.23 $X2=0 $Y2=0
cc_138 N_C_c_180_n N_B_c_226_n 2.63776e-19 $X=1.43 $Y=1.155 $X2=0 $Y2=0
cc_139 N_C_c_181_n A 0.00144442f $X=1.9 $Y=1.23 $X2=0 $Y2=0
cc_140 N_C_M1008_g A 0.0113271f $X=1.975 $Y=2.195 $X2=0 $Y2=0
cc_141 N_C_c_180_n N_A_215_125#_c_292_n 0.00942018f $X=1.43 $Y=1.155 $X2=0 $Y2=0
cc_142 N_C_c_182_n N_A_215_125#_c_292_n 0.00364557f $X=1.505 $Y=1.23 $X2=0 $Y2=0
cc_143 N_C_M1008_g N_A_215_125#_c_293_n 0.00513201f $X=1.975 $Y=2.195 $X2=0
+ $Y2=0
cc_144 C N_A_215_125#_c_293_n 0.00870619f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_145 N_C_c_181_n N_A_215_125#_c_294_n 0.0241492f $X=1.9 $Y=1.23 $X2=0 $Y2=0
cc_146 N_C_c_182_n N_A_215_125#_c_294_n 0.00528402f $X=1.505 $Y=1.23 $X2=0 $Y2=0
cc_147 N_C_M1008_g N_A_215_125#_c_294_n 0.00622105f $X=1.975 $Y=2.195 $X2=0
+ $Y2=0
cc_148 N_C_M1008_g N_A_215_125#_c_313_n 0.0162978f $X=1.975 $Y=2.195 $X2=0 $Y2=0
cc_149 C N_A_215_125#_c_313_n 0.0324279f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_150 N_C_c_186_n N_A_215_125#_c_313_n 7.47713e-19 $X=1.885 $Y=2.94 $X2=0 $Y2=0
cc_151 N_C_c_181_n N_A_215_125#_c_332_n 4.03038e-19 $X=1.9 $Y=1.23 $X2=0 $Y2=0
cc_152 N_C_M1008_g N_A_215_125#_c_301_n 0.00472319f $X=1.975 $Y=2.195 $X2=0
+ $Y2=0
cc_153 C N_A_215_125#_c_301_n 0.0105642f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_154 N_C_c_180_n N_A_215_125#_c_315_n 0.00504799f $X=1.43 $Y=1.155 $X2=0 $Y2=0
cc_155 N_C_c_182_n N_A_215_125#_c_295_n 0.00171366f $X=1.505 $Y=1.23 $X2=0 $Y2=0
cc_156 C N_A_215_125#_c_302_n 0.0109901f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_157 C N_A_215_125#_c_303_n 0.00160457f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_158 N_C_c_186_n N_A_215_125#_c_303_n 0.0090743f $X=1.885 $Y=2.94 $X2=0 $Y2=0
cc_159 C N_VPWR_c_399_n 0.0258132f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_160 C N_VPWR_c_401_n 0.0571344f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_161 N_C_c_186_n N_VPWR_c_401_n 0.00617531f $X=1.885 $Y=2.94 $X2=0 $Y2=0
cc_162 C N_VPWR_c_398_n 0.0403696f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_163 N_C_c_186_n N_VPWR_c_398_n 0.00817532f $X=1.885 $Y=2.94 $X2=0 $Y2=0
cc_164 N_C_c_180_n N_VGND_c_464_n 0.00777773f $X=1.43 $Y=1.155 $X2=0 $Y2=0
cc_165 N_C_c_181_n N_VGND_c_464_n 0.00426967f $X=1.9 $Y=1.23 $X2=0 $Y2=0
cc_166 N_C_c_180_n N_VGND_c_468_n 0.00380255f $X=1.43 $Y=1.155 $X2=0 $Y2=0
cc_167 N_C_c_180_n N_VGND_c_470_n 0.00469432f $X=1.43 $Y=1.155 $X2=0 $Y2=0
cc_168 B N_A_M1011_g 0.00486092f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_169 N_B_c_226_n N_A_M1011_g 0.0312751f $X=2.245 $Y=0.35 $X2=0 $Y2=0
cc_170 N_B_M1002_g A 0.0102127f $X=2.335 $Y=0.835 $X2=0 $Y2=0
cc_171 N_B_M1002_g N_A_c_254_n 0.0669187f $X=2.335 $Y=0.835 $X2=0 $Y2=0
cc_172 B N_A_215_125#_M1002_d 0.00191751f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_173 N_B_M1002_g N_A_215_125#_c_294_n 0.0112932f $X=2.335 $Y=0.835 $X2=0 $Y2=0
cc_174 B N_A_215_125#_c_294_n 0.00827314f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_175 N_B_M1002_g N_A_215_125#_c_313_n 0.0194505f $X=2.335 $Y=0.835 $X2=0 $Y2=0
cc_176 N_B_M1002_g N_A_215_125#_c_332_n 0.0152299f $X=2.335 $Y=0.835 $X2=0 $Y2=0
cc_177 B N_A_215_125#_c_332_n 0.0154218f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_178 N_B_M1002_g N_A_215_125#_c_301_n 0.00445047f $X=2.335 $Y=0.835 $X2=0
+ $Y2=0
cc_179 N_B_M1002_g N_VPWR_c_398_n 0.00393927f $X=2.335 $Y=0.835 $X2=0 $Y2=0
cc_180 B N_VGND_M1006_d 0.00275636f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_181 N_B_M1002_g N_VGND_c_464_n 0.00732016f $X=2.335 $Y=0.835 $X2=0 $Y2=0
cc_182 B N_VGND_c_464_n 0.0229984f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_183 N_B_c_226_n N_VGND_c_464_n 0.00372015f $X=2.245 $Y=0.35 $X2=0 $Y2=0
cc_184 B N_VGND_c_465_n 0.0299028f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_185 N_B_c_226_n N_VGND_c_465_n 0.0024312f $X=2.245 $Y=0.35 $X2=0 $Y2=0
cc_186 B N_VGND_c_466_n 0.0406224f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_187 N_B_c_226_n N_VGND_c_466_n 0.00651318f $X=2.245 $Y=0.35 $X2=0 $Y2=0
cc_188 B N_VGND_c_470_n 0.0232288f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_189 N_B_c_226_n N_VGND_c_470_n 0.0101042f $X=2.245 $Y=0.35 $X2=0 $Y2=0
cc_190 N_A_M1011_g N_A_215_125#_M1007_g 0.0213173f $X=2.765 $Y=0.835 $X2=0 $Y2=0
cc_191 A N_A_215_125#_M1007_g 0.00419239f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A_c_254_n N_A_215_125#_M1007_g 0.0134293f $X=2.785 $Y=1.66 $X2=0 $Y2=0
cc_193 N_A_M1010_g N_A_215_125#_c_299_n 0.0149381f $X=2.695 $Y=2.195 $X2=0 $Y2=0
cc_194 A N_A_215_125#_c_299_n 0.00264771f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A_c_254_n N_A_215_125#_c_299_n 0.00661485f $X=2.785 $Y=1.66 $X2=0 $Y2=0
cc_196 A N_A_215_125#_c_293_n 0.0134121f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A_M1011_g N_A_215_125#_c_294_n 0.00574949f $X=2.765 $Y=0.835 $X2=0
+ $Y2=0
cc_198 A N_A_215_125#_c_294_n 0.080853f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_199 N_A_c_254_n N_A_215_125#_c_294_n 0.00207212f $X=2.785 $Y=1.66 $X2=0 $Y2=0
cc_200 N_A_M1010_g N_A_215_125#_c_313_n 0.00898785f $X=2.695 $Y=2.195 $X2=0
+ $Y2=0
cc_201 A N_A_215_125#_c_313_n 0.0491611f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_202 N_A_M1011_g N_A_215_125#_c_332_n 0.00927039f $X=2.765 $Y=0.835 $X2=0
+ $Y2=0
cc_203 N_A_M1010_g N_A_215_125#_c_301_n 0.00426762f $X=2.695 $Y=2.195 $X2=0
+ $Y2=0
cc_204 N_A_M1010_g N_A_215_125#_c_302_n 7.61518e-19 $X=2.695 $Y=2.195 $X2=0
+ $Y2=0
cc_205 N_A_M1010_g N_A_215_125#_c_303_n 0.00919007f $X=2.695 $Y=2.195 $X2=0
+ $Y2=0
cc_206 N_A_M1010_g N_VPWR_c_400_n 0.0013097f $X=2.695 $Y=2.195 $X2=0 $Y2=0
cc_207 N_A_M1010_g N_VPWR_c_421_n 0.00183352f $X=2.695 $Y=2.195 $X2=0 $Y2=0
cc_208 A N_VPWR_c_421_n 0.0117596f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A_c_254_n N_VPWR_c_421_n 0.00240497f $X=2.785 $Y=1.66 $X2=0 $Y2=0
cc_210 A X 0.0137596f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_211 N_A_M1011_g N_VGND_c_465_n 0.00538278f $X=2.765 $Y=0.835 $X2=0 $Y2=0
cc_212 A N_VGND_c_465_n 0.00640199f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A_c_254_n N_VGND_c_465_n 8.10212e-19 $X=2.785 $Y=1.66 $X2=0 $Y2=0
cc_214 N_A_M1011_g N_VGND_c_466_n 0.00331069f $X=2.765 $Y=0.835 $X2=0 $Y2=0
cc_215 N_A_M1011_g N_VGND_c_470_n 0.00359898f $X=2.765 $Y=0.835 $X2=0 $Y2=0
cc_216 N_A_215_125#_c_296_n N_VPWR_c_400_n 0.0153837f $X=3.16 $Y=2.85 $X2=0
+ $Y2=0
cc_217 N_A_215_125#_M1001_g N_VPWR_c_400_n 0.00944898f $X=3.235 $Y=2.195 $X2=0
+ $Y2=0
cc_218 N_A_215_125#_c_301_n N_VPWR_c_400_n 0.0215009f $X=2.57 $Y=2.855 $X2=0
+ $Y2=0
cc_219 N_A_215_125#_c_302_n N_VPWR_c_400_n 0.0118902f $X=2.65 $Y=2.94 $X2=0
+ $Y2=0
cc_220 N_A_215_125#_c_303_n N_VPWR_c_400_n 0.00351565f $X=2.65 $Y=2.85 $X2=0
+ $Y2=0
cc_221 N_A_215_125#_c_296_n N_VPWR_c_421_n 0.0048325f $X=3.16 $Y=2.85 $X2=0
+ $Y2=0
cc_222 N_A_215_125#_M1001_g N_VPWR_c_421_n 0.00199068f $X=3.235 $Y=2.195 $X2=0
+ $Y2=0
cc_223 N_A_215_125#_c_313_n N_VPWR_c_421_n 0.0141759f $X=2.485 $Y=2.17 $X2=0
+ $Y2=0
cc_224 N_A_215_125#_c_301_n N_VPWR_c_421_n 0.00203065f $X=2.57 $Y=2.855 $X2=0
+ $Y2=0
cc_225 N_A_215_125#_c_296_n N_VPWR_c_401_n 0.00445258f $X=3.16 $Y=2.85 $X2=0
+ $Y2=0
cc_226 N_A_215_125#_c_302_n N_VPWR_c_401_n 0.0152941f $X=2.65 $Y=2.94 $X2=0
+ $Y2=0
cc_227 N_A_215_125#_c_303_n N_VPWR_c_401_n 0.00593936f $X=2.65 $Y=2.85 $X2=0
+ $Y2=0
cc_228 N_A_215_125#_c_296_n N_VPWR_c_404_n 0.00449461f $X=3.16 $Y=2.85 $X2=0
+ $Y2=0
cc_229 N_A_215_125#_c_296_n N_VPWR_c_398_n 0.009566f $X=3.16 $Y=2.85 $X2=0 $Y2=0
cc_230 N_A_215_125#_c_302_n N_VPWR_c_398_n 0.0104794f $X=2.65 $Y=2.94 $X2=0
+ $Y2=0
cc_231 N_A_215_125#_c_303_n N_VPWR_c_398_n 0.00799516f $X=2.65 $Y=2.85 $X2=0
+ $Y2=0
cc_232 N_A_215_125#_c_313_n A_338_397# 0.00250064f $X=2.485 $Y=2.17 $X2=-0.19
+ $Y2=-0.245
cc_233 N_A_215_125#_c_313_n A_410_397# 0.00273154f $X=2.485 $Y=2.17 $X2=-0.19
+ $Y2=-0.245
cc_234 N_A_215_125#_c_313_n A_482_397# 0.00196393f $X=2.485 $Y=2.17 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_215_125#_c_301_n A_482_397# 7.62448e-19 $X=2.57 $Y=2.855 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_215_125#_M1001_g X 0.00219531f $X=3.235 $Y=2.195 $X2=0 $Y2=0
cc_237 N_A_215_125#_M1007_g X 0.031562f $X=3.255 $Y=0.835 $X2=0 $Y2=0
cc_238 N_A_215_125#_c_294_n X 0.00488805f $X=2.385 $Y=1.31 $X2=0 $Y2=0
cc_239 N_A_215_125#_c_332_n X 0.0062003f $X=2.55 $Y=0.92 $X2=0 $Y2=0
cc_240 N_A_215_125#_c_296_n X 0.00757462f $X=3.16 $Y=2.85 $X2=0 $Y2=0
cc_241 N_A_215_125#_M1001_g X 0.00757462f $X=3.235 $Y=2.195 $X2=0 $Y2=0
cc_242 N_A_215_125#_c_294_n N_VGND_c_464_n 0.010902f $X=2.385 $Y=1.31 $X2=0
+ $Y2=0
cc_243 N_A_215_125#_c_332_n N_VGND_c_464_n 0.00286318f $X=2.55 $Y=0.92 $X2=0
+ $Y2=0
cc_244 N_A_215_125#_c_315_n N_VGND_c_464_n 0.0133701f $X=1.33 $Y=0.855 $X2=0
+ $Y2=0
cc_245 N_A_215_125#_M1007_g N_VGND_c_465_n 0.0025396f $X=3.255 $Y=0.835 $X2=0
+ $Y2=0
cc_246 N_A_215_125#_c_332_n N_VGND_c_465_n 0.0068835f $X=2.55 $Y=0.92 $X2=0
+ $Y2=0
cc_247 N_A_215_125#_c_315_n N_VGND_c_468_n 0.0042271f $X=1.33 $Y=0.855 $X2=0
+ $Y2=0
cc_248 N_A_215_125#_M1007_g N_VGND_c_469_n 0.00415323f $X=3.255 $Y=0.835 $X2=0
+ $Y2=0
cc_249 N_A_215_125#_M1007_g N_VGND_c_470_n 0.00469432f $X=3.255 $Y=0.835 $X2=0
+ $Y2=0
cc_250 N_A_215_125#_c_315_n N_VGND_c_470_n 0.00950543f $X=1.33 $Y=0.855 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_400_n X 0.0342148f $X=3.08 $Y=3.245 $X2=0 $Y2=0
cc_252 N_VPWR_c_404_n X 0.010134f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_253 N_VPWR_c_398_n X 0.0115466f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_254 X N_VGND_c_465_n 0.0171985f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_255 X N_VGND_c_469_n 0.00893474f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_256 X N_VGND_c_470_n 0.0101801f $X=3.515 $Y=0.47 $X2=0 $Y2=0
