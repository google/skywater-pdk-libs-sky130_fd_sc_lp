* File: sky130_fd_sc_lp__xnor2_m.pxi.spice
* Created: Fri Aug 28 11:35:31 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR2_M%A N_A_M1007_g N_A_c_61_n N_A_M1001_g N_A_M1003_g
+ N_A_M1008_g N_A_c_63_n A A A N_A_c_65_n PM_SKY130_FD_SC_LP__XNOR2_M%A
x_PM_SKY130_FD_SC_LP__XNOR2_M%B N_B_M1002_g N_B_M1000_g N_B_c_109_n N_B_c_110_n
+ N_B_M1005_g N_B_M1009_g B B B N_B_c_113_n PM_SKY130_FD_SC_LP__XNOR2_M%B
x_PM_SKY130_FD_SC_LP__XNOR2_M%A_56_90# N_A_56_90#_M1002_s N_A_56_90#_M1000_d
+ N_A_56_90#_c_157_n N_A_56_90#_c_158_n N_A_56_90#_M1004_g N_A_56_90#_M1006_g
+ N_A_56_90#_c_161_n N_A_56_90#_c_162_n N_A_56_90#_c_168_n N_A_56_90#_c_169_n
+ N_A_56_90#_c_187_n N_A_56_90#_c_170_n N_A_56_90#_c_163_n N_A_56_90#_c_164_n
+ N_A_56_90#_c_165_n N_A_56_90#_c_172_n PM_SKY130_FD_SC_LP__XNOR2_M%A_56_90#
x_PM_SKY130_FD_SC_LP__XNOR2_M%VPWR N_VPWR_M1000_s N_VPWR_M1001_d N_VPWR_M1004_d
+ N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ N_VPWR_c_232_n VPWR N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n
+ N_VPWR_c_219_n PM_SKY130_FD_SC_LP__XNOR2_M%VPWR
x_PM_SKY130_FD_SC_LP__XNOR2_M%Y N_Y_M1006_s N_Y_M1009_d N_Y_c_256_n Y Y Y Y Y
+ N_Y_c_262_n PM_SKY130_FD_SC_LP__XNOR2_M%Y
x_PM_SKY130_FD_SC_LP__XNOR2_M%VGND N_VGND_M1007_d N_VGND_M1005_d N_VGND_c_281_n
+ N_VGND_c_282_n N_VGND_c_283_n N_VGND_c_284_n VGND N_VGND_c_285_n
+ N_VGND_c_286_n N_VGND_c_287_n N_VGND_c_288_n PM_SKY130_FD_SC_LP__XNOR2_M%VGND
x_PM_SKY130_FD_SC_LP__XNOR2_M%A_297_90# N_A_297_90#_M1003_d N_A_297_90#_M1006_d
+ N_A_297_90#_c_322_n N_A_297_90#_c_323_n N_A_297_90#_c_324_n
+ PM_SKY130_FD_SC_LP__XNOR2_M%A_297_90#
cc_1 VNB N_A_M1007_g 0.0233457f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.66
cc_2 VNB N_A_c_61_n 0.00242284f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.8
cc_3 VNB N_A_M1003_g 0.0221223f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.66
cc_4 VNB N_A_c_63_n 0.0183641f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.28
cc_5 VNB A 0.0121511f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_6 VNB N_A_c_65_n 0.0297178f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.295
cc_7 VNB N_B_M1002_g 0.0553696f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.66
cc_8 VNB N_B_M1005_g 0.0543604f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.66
cc_9 VNB N_A_56_90#_c_157_n 0.0113895f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=2.32
cc_10 VNB N_A_56_90#_c_158_n 0.0192639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_56_90#_M1004_g 0.0163653f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.66
cc_12 VNB N_A_56_90#_M1006_g 0.0483998f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=2.32
cc_13 VNB N_A_56_90#_c_161_n 0.0238539f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.28
cc_14 VNB N_A_56_90#_c_162_n 0.0392328f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.8
cc_15 VNB N_A_56_90#_c_163_n 0.00406093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_56_90#_c_164_n 0.0147762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_56_90#_c_165_n 0.00868346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_219_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.48
cc_19 VNB N_Y_c_256_n 0.00275203f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.13
cc_20 VNB Y 0.0109558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_281_n 0.0124918f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.66
cc_22 VNB N_VGND_c_282_n 0.0053519f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.66
cc_23 VNB N_VGND_c_283_n 0.00355854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_284_n 0.0129086f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=2.32
cc_25 VNB N_VGND_c_285_n 0.0353187f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.65
cc_26 VNB N_VGND_c_286_n 0.0525549f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_27 VNB N_VGND_c_287_n 0.23258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_288_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_297_90#_c_322_n 0.0360272f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=2.32
cc_30 VNB N_A_297_90#_c_323_n 4.08405e-19 $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.66
cc_31 VNB N_A_297_90#_c_324_n 0.00304379f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.8
cc_32 VPB N_A_c_61_n 0.0155706f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=1.8
cc_33 VPB N_A_M1001_g 0.0233546f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=2.32
cc_34 VPB N_A_M1008_g 0.0227909f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=2.32
cc_35 VPB A 0.00478329f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_36 VPB N_B_M1002_g 0.0509583f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=0.66
cc_37 VPB N_B_c_109_n 0.0662308f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=2.32
cc_38 VPB N_B_c_110_n 0.0106743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_B_M1005_g 0.0375426f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=0.66
cc_40 VPB B 0.0275539f $X=-0.19 $Y=1.655 $X2=1.23 $Y2=1.28
cc_41 VPB N_B_c_113_n 0.0418418f $X=-0.19 $Y=1.655 $X2=1.265 $Y2=1.8
cc_42 VPB N_A_56_90#_M1004_g 0.0518149f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=0.66
cc_43 VPB N_A_56_90#_c_162_n 0.0131231f $X=-0.19 $Y=1.655 $X2=1.265 $Y2=1.8
cc_44 VPB N_A_56_90#_c_168_n 0.00821678f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_45 VPB N_A_56_90#_c_169_n 0.00931523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_56_90#_c_170_n 0.0270883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_56_90#_c_164_n 0.0287748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_56_90#_c_172_n 0.00157719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_220_n 0.0161782f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=0.66
cc_50 VPB N_VPWR_c_221_n 0.0379128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_222_n 0.0107519f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=2.32
cc_52 VPB N_VPWR_c_223_n 0.0142828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_224_n 0.0373033f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=1.13
cc_54 VPB N_VPWR_c_225_n 0.016802f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_55 VPB N_VPWR_c_226_n 0.0433262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_227_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_219_n 0.0857124f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.48
cc_58 VPB Y 0.00304833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 N_A_M1007_g N_B_M1002_g 0.0586995f $X=0.98 $Y=0.66 $X2=0 $Y2=0
cc_60 A N_B_M1002_g 0.0178575f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A_c_65_n N_B_M1002_g 0.0464563f $X=1.29 $Y=1.295 $X2=0 $Y2=0
cc_62 N_A_M1001_g N_B_c_109_n 0.00918879f $X=1.05 $Y=2.32 $X2=0 $Y2=0
cc_63 N_A_M1008_g N_B_c_109_n 0.00925194f $X=1.48 $Y=2.32 $X2=0 $Y2=0
cc_64 N_A_c_61_n N_B_M1005_g 0.0642926f $X=1.05 $Y=1.8 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_B_M1005_g 0.0467659f $X=1.41 $Y=0.66 $X2=0 $Y2=0
cc_66 A N_B_M1005_g 0.00910798f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_67 A N_A_56_90#_c_158_n 0.00141838f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_68 A N_A_56_90#_c_162_n 0.0347785f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_69 A N_A_56_90#_c_168_n 0.00858322f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_c_61_n N_A_56_90#_c_170_n 0.00276204f $X=1.05 $Y=1.8 $X2=0 $Y2=0
cc_71 N_A_M1001_g N_A_56_90#_c_170_n 0.0140674f $X=1.05 $Y=2.32 $X2=0 $Y2=0
cc_72 N_A_M1008_g N_A_56_90#_c_170_n 0.0136263f $X=1.48 $Y=2.32 $X2=0 $Y2=0
cc_73 A N_A_56_90#_c_170_n 0.0632125f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_74 A N_A_56_90#_c_163_n 0.016482f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_M1007_g N_A_56_90#_c_165_n 5.86076e-19 $X=0.98 $Y=0.66 $X2=0 $Y2=0
cc_76 A N_A_56_90#_c_172_n 0.0146064f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_M1001_g N_VPWR_c_221_n 6.85327e-19 $X=1.05 $Y=2.32 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_VPWR_c_222_n 0.00423953f $X=1.05 $Y=2.32 $X2=0 $Y2=0
cc_79 N_A_M1008_g N_VPWR_c_222_n 0.00352685f $X=1.48 $Y=2.32 $X2=0 $Y2=0
cc_80 N_A_M1001_g N_VPWR_c_232_n 0.00306117f $X=1.05 $Y=2.32 $X2=0 $Y2=0
cc_81 N_A_M1008_g N_VPWR_c_232_n 0.00415887f $X=1.48 $Y=2.32 $X2=0 $Y2=0
cc_82 N_A_M1007_g N_VGND_c_281_n 0.00358099f $X=0.98 $Y=0.66 $X2=0 $Y2=0
cc_83 N_A_M1003_g N_VGND_c_281_n 0.00127127f $X=1.41 $Y=0.66 $X2=0 $Y2=0
cc_84 N_A_c_61_n N_VGND_c_282_n 2.00262e-19 $X=1.05 $Y=1.8 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_VGND_c_282_n 0.0111847f $X=1.41 $Y=0.66 $X2=0 $Y2=0
cc_86 A N_VGND_c_282_n 0.036919f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A_M1007_g N_VGND_c_283_n 0.00516145f $X=0.98 $Y=0.66 $X2=0 $Y2=0
cc_88 N_A_c_63_n N_VGND_c_283_n 0.00296805f $X=1.195 $Y=1.28 $X2=0 $Y2=0
cc_89 A N_VGND_c_283_n 0.0158841f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A_M1007_g N_VGND_c_285_n 0.00520566f $X=0.98 $Y=0.66 $X2=0 $Y2=0
cc_91 N_A_M1003_g N_VGND_c_286_n 0.0045043f $X=1.41 $Y=0.66 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_VGND_c_287_n 0.00520574f $X=0.98 $Y=0.66 $X2=0 $Y2=0
cc_93 N_A_M1003_g N_VGND_c_287_n 0.00437282f $X=1.41 $Y=0.66 $X2=0 $Y2=0
cc_94 N_A_M1003_g N_A_297_90#_c_324_n 0.00593437f $X=1.41 $Y=0.66 $X2=0 $Y2=0
cc_95 N_B_M1005_g N_A_56_90#_c_158_n 0.0417769f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_96 B N_A_56_90#_M1004_g 0.00191729f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_97 N_B_M1002_g N_A_56_90#_c_162_n 0.0303355f $X=0.62 $Y=0.66 $X2=0 $Y2=0
cc_98 N_B_M1002_g N_A_56_90#_c_168_n 0.0184639f $X=0.62 $Y=0.66 $X2=0 $Y2=0
cc_99 N_B_c_109_n N_A_56_90#_c_187_n 0.00376433f $X=1.765 $Y=2.975 $X2=0 $Y2=0
cc_100 N_B_M1005_g N_A_56_90#_c_170_n 0.017969f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_101 B N_A_56_90#_c_170_n 0.0196396f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_102 N_B_c_113_n N_A_56_90#_c_170_n 8.77211e-19 $X=1.93 $Y=2.885 $X2=0 $Y2=0
cc_103 N_B_M1005_g N_A_56_90#_c_163_n 0.00240468f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_104 N_B_M1002_g N_A_56_90#_c_165_n 0.00509686f $X=0.62 $Y=0.66 $X2=0 $Y2=0
cc_105 N_B_M1002_g N_VPWR_c_221_n 0.0180733f $X=0.62 $Y=0.66 $X2=0 $Y2=0
cc_106 N_B_c_110_n N_VPWR_c_221_n 0.00759502f $X=0.695 $Y=2.975 $X2=0 $Y2=0
cc_107 N_B_M1002_g N_VPWR_c_222_n 0.00458799f $X=0.62 $Y=0.66 $X2=0 $Y2=0
cc_108 N_B_c_109_n N_VPWR_c_222_n 0.0179126f $X=1.765 $Y=2.975 $X2=0 $Y2=0
cc_109 N_B_M1005_g N_VPWR_c_222_n 0.00193052f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_110 B N_VPWR_c_222_n 0.0143687f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_111 B N_VPWR_c_224_n 0.0227194f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_112 N_B_c_109_n N_VPWR_c_232_n 0.00341545f $X=1.765 $Y=2.975 $X2=0 $Y2=0
cc_113 N_B_M1005_g N_VPWR_c_232_n 0.00104529f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_114 N_B_c_110_n N_VPWR_c_225_n 0.017109f $X=0.695 $Y=2.975 $X2=0 $Y2=0
cc_115 N_B_c_109_n N_VPWR_c_226_n 0.0213085f $X=1.765 $Y=2.975 $X2=0 $Y2=0
cc_116 B N_VPWR_c_226_n 0.0440299f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_117 N_B_c_110_n N_VPWR_c_219_n 0.0422803f $X=0.695 $Y=2.975 $X2=0 $Y2=0
cc_118 B N_VPWR_c_219_n 0.0398621f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_119 N_B_M1005_g Y 0.00949544f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_120 N_B_M1005_g Y 0.00701747f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_121 B Y 0.0220415f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_122 B N_Y_c_262_n 0.0101004f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_123 N_B_M1005_g N_VGND_c_282_n 0.0165917f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_124 N_B_M1005_g N_VGND_c_284_n 0.00150478f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_125 N_B_M1002_g N_VGND_c_285_n 0.00500116f $X=0.62 $Y=0.66 $X2=0 $Y2=0
cc_126 N_B_M1005_g N_VGND_c_286_n 8.17648e-19 $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_127 N_B_M1002_g N_VGND_c_287_n 0.00520574f $X=0.62 $Y=0.66 $X2=0 $Y2=0
cc_128 N_B_M1005_g N_A_297_90#_c_322_n 0.00930696f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_129 N_B_M1005_g N_A_297_90#_c_324_n 0.0113461f $X=1.84 $Y=0.66 $X2=0 $Y2=0
cc_130 N_A_56_90#_c_168_n N_VPWR_c_221_n 0.00992485f $X=0.75 $Y=2.015 $X2=0
+ $Y2=0
cc_131 N_A_56_90#_c_169_n N_VPWR_c_221_n 0.0149239f $X=0.41 $Y=2.015 $X2=0 $Y2=0
cc_132 N_A_56_90#_M1004_g N_VPWR_c_224_n 0.0065579f $X=2.74 $Y=2.32 $X2=0 $Y2=0
cc_133 N_A_56_90#_c_170_n N_VPWR_c_232_n 0.0193134f $X=2.205 $Y=2.015 $X2=0
+ $Y2=0
cc_134 N_A_56_90#_M1004_g N_VPWR_c_226_n 0.00206046f $X=2.74 $Y=2.32 $X2=0 $Y2=0
cc_135 N_A_56_90#_M1004_g N_VPWR_c_219_n 0.00254193f $X=2.74 $Y=2.32 $X2=0 $Y2=0
cc_136 N_A_56_90#_c_157_n N_Y_c_256_n 0.00196876f $X=2.665 $Y=1.355 $X2=0 $Y2=0
cc_137 N_A_56_90#_M1006_g N_Y_c_256_n 0.00592697f $X=2.87 $Y=0.66 $X2=0 $Y2=0
cc_138 N_A_56_90#_c_161_n N_Y_c_256_n 0.00143753f $X=2.87 $Y=1.355 $X2=0 $Y2=0
cc_139 N_A_56_90#_c_157_n Y 0.00658661f $X=2.665 $Y=1.355 $X2=0 $Y2=0
cc_140 N_A_56_90#_M1004_g Y 0.04149f $X=2.74 $Y=2.32 $X2=0 $Y2=0
cc_141 N_A_56_90#_M1006_g Y 0.0163878f $X=2.87 $Y=0.66 $X2=0 $Y2=0
cc_142 N_A_56_90#_c_161_n Y 0.00810804f $X=2.87 $Y=1.355 $X2=0 $Y2=0
cc_143 N_A_56_90#_c_170_n Y 0.0136946f $X=2.205 $Y=2.015 $X2=0 $Y2=0
cc_144 N_A_56_90#_c_163_n Y 0.0439021f $X=2.29 $Y=1.445 $X2=0 $Y2=0
cc_145 N_A_56_90#_c_164_n Y 0.00322571f $X=2.29 $Y=1.445 $X2=0 $Y2=0
cc_146 N_A_56_90#_c_170_n Y 0.0121311f $X=2.205 $Y=2.015 $X2=0 $Y2=0
cc_147 N_A_56_90#_c_164_n Y 0.00356582f $X=2.29 $Y=1.445 $X2=0 $Y2=0
cc_148 N_A_56_90#_M1004_g N_Y_c_262_n 0.00796994f $X=2.74 $Y=2.32 $X2=0 $Y2=0
cc_149 N_A_56_90#_c_158_n N_VGND_c_284_n 0.00400518f $X=2.455 $Y=1.355 $X2=0
+ $Y2=0
cc_150 N_A_56_90#_c_163_n N_VGND_c_284_n 0.00595928f $X=2.29 $Y=1.445 $X2=0
+ $Y2=0
cc_151 N_A_56_90#_c_165_n N_VGND_c_285_n 0.00557519f $X=0.405 $Y=0.725 $X2=0
+ $Y2=0
cc_152 N_A_56_90#_M1006_g N_VGND_c_286_n 8.23325e-19 $X=2.87 $Y=0.66 $X2=0 $Y2=0
cc_153 N_A_56_90#_c_165_n N_VGND_c_287_n 0.00958017f $X=0.405 $Y=0.725 $X2=0
+ $Y2=0
cc_154 N_A_56_90#_M1006_g N_A_297_90#_c_322_n 0.0149949f $X=2.87 $Y=0.66 $X2=0
+ $Y2=0
cc_155 N_A_56_90#_M1006_g N_A_297_90#_c_323_n 3.52891e-19 $X=2.87 $Y=0.66 $X2=0
+ $Y2=0
cc_156 N_VPWR_c_224_n Y 0.00674363f $X=2.99 $Y=2.345 $X2=0 $Y2=0
cc_157 N_VPWR_c_224_n N_Y_c_262_n 0.0155273f $X=2.99 $Y=2.345 $X2=0 $Y2=0
cc_158 N_Y_c_256_n N_VGND_c_284_n 0.0161706f $X=2.655 $Y=0.725 $X2=0 $Y2=0
cc_159 Y N_VGND_c_284_n 0.0118715f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_160 N_Y_c_256_n N_A_297_90#_c_322_n 0.0214064f $X=2.655 $Y=0.725 $X2=0 $Y2=0
cc_161 N_VGND_c_282_n N_A_297_90#_M1003_d 0.0017847f $X=1.97 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_162 N_VGND_c_282_n N_A_297_90#_c_322_n 0.00460834f $X=1.97 $Y=0.945 $X2=0
+ $Y2=0
cc_163 N_VGND_c_284_n N_A_297_90#_c_322_n 0.0234181f $X=2.135 $Y=0.725 $X2=0
+ $Y2=0
cc_164 N_VGND_c_286_n N_A_297_90#_c_322_n 0.083389f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_165 N_VGND_c_287_n N_A_297_90#_c_322_n 0.0523493f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_166 N_VGND_c_281_n N_A_297_90#_c_324_n 0.0214824f $X=1.195 $Y=0.725 $X2=0
+ $Y2=0
cc_167 N_VGND_c_282_n N_A_297_90#_c_324_n 0.0153029f $X=1.97 $Y=0.945 $X2=0
+ $Y2=0
cc_168 N_VGND_c_286_n N_A_297_90#_c_324_n 0.0206856f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_169 N_VGND_c_287_n N_A_297_90#_c_324_n 0.0124904f $X=3.12 $Y=0 $X2=0 $Y2=0
