* File: sky130_fd_sc_lp__or3b_2.pxi.spice
* Created: Wed Sep  2 10:31:12 2020
* 
x_PM_SKY130_FD_SC_LP__OR3B_2%C_N N_C_N_M1004_g N_C_N_c_78_n N_C_N_M1002_g C_N
+ N_C_N_c_76_n N_C_N_c_77_n PM_SKY130_FD_SC_LP__OR3B_2%C_N
x_PM_SKY130_FD_SC_LP__OR3B_2%A_195_21# N_A_195_21#_M1011_d N_A_195_21#_M1005_d
+ N_A_195_21#_M1009_d N_A_195_21#_c_99_n N_A_195_21#_M1001_g N_A_195_21#_M1006_g
+ N_A_195_21#_c_101_n N_A_195_21#_M1007_g N_A_195_21#_M1010_g
+ N_A_195_21#_c_103_n N_A_195_21#_c_104_n N_A_195_21#_c_105_n
+ N_A_195_21#_c_172_p N_A_195_21#_c_106_n N_A_195_21#_c_107_n
+ N_A_195_21#_c_108_n N_A_195_21#_c_109_n N_A_195_21#_c_110_n
+ N_A_195_21#_c_111_n PM_SKY130_FD_SC_LP__OR3B_2%A_195_21#
x_PM_SKY130_FD_SC_LP__OR3B_2%A N_A_M1011_g N_A_M1000_g A A N_A_c_203_n
+ N_A_c_204_n PM_SKY130_FD_SC_LP__OR3B_2%A
x_PM_SKY130_FD_SC_LP__OR3B_2%B N_B_c_245_n N_B_M1003_g N_B_M1008_g N_B_c_247_n B
+ B B N_B_c_249_n N_B_c_250_n PM_SKY130_FD_SC_LP__OR3B_2%B
x_PM_SKY130_FD_SC_LP__OR3B_2%A_33_131# N_A_33_131#_M1004_s N_A_33_131#_M1002_s
+ N_A_33_131#_c_291_n N_A_33_131#_M1005_g N_A_33_131#_M1009_g
+ N_A_33_131#_c_292_n N_A_33_131#_c_293_n N_A_33_131#_c_300_n
+ N_A_33_131#_c_294_n N_A_33_131#_c_295_n N_A_33_131#_c_296_n
+ N_A_33_131#_c_297_n N_A_33_131#_c_302_n N_A_33_131#_c_303_n
+ N_A_33_131#_c_304_n N_A_33_131#_c_305_n PM_SKY130_FD_SC_LP__OR3B_2%A_33_131#
x_PM_SKY130_FD_SC_LP__OR3B_2%VPWR N_VPWR_M1002_d N_VPWR_M1010_d N_VPWR_c_377_n
+ N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n VPWR
+ N_VPWR_c_382_n N_VPWR_c_376_n N_VPWR_c_384_n PM_SKY130_FD_SC_LP__OR3B_2%VPWR
x_PM_SKY130_FD_SC_LP__OR3B_2%X N_X_M1001_d N_X_M1006_s N_X_c_409_n N_X_c_411_n X
+ X N_X_c_424_n X PM_SKY130_FD_SC_LP__OR3B_2%X
x_PM_SKY130_FD_SC_LP__OR3B_2%VGND N_VGND_M1004_d N_VGND_M1007_s N_VGND_M1003_d
+ N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n VGND N_VGND_c_447_n
+ N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n
+ N_VGND_c_453_n N_VGND_c_454_n PM_SKY130_FD_SC_LP__OR3B_2%VGND
cc_1 VNB N_C_N_M1004_g 0.034327f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.865
cc_2 VNB N_C_N_c_76_n 0.0135774f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.51
cc_3 VNB N_C_N_c_77_n 0.0391802f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.535
cc_4 VNB N_A_195_21#_c_99_n 0.0189365f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.535
cc_5 VNB N_A_195_21#_M1006_g 0.00695666f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.577
cc_6 VNB N_A_195_21#_c_101_n 0.0163436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_195_21#_M1010_g 0.00662945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_195_21#_c_103_n 0.00352885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_195_21#_c_104_n 0.0511253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_195_21#_c_105_n 0.00837519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_195_21#_c_106_n 0.00221551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_195_21#_c_107_n 0.0143649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_195_21#_c_108_n 0.0200792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_195_21#_c_109_n 0.0309983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_195_21#_c_110_n 0.00701581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_195_21#_c_111_n 0.00692367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_M1011_g 0.0490811f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.865
cc_18 VNB N_A_c_203_n 0.0241778f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.725
cc_19 VNB N_A_c_204_n 0.00201086f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.577
cc_20 VNB N_B_c_245_n 0.0165803f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.345
cc_21 VNB N_B_M1008_g 0.0108455f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_B_c_247_n 0.012465f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.51
cc_23 VNB B 0.00553531f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.725
cc_24 VNB N_B_c_249_n 0.0325031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_c_250_n 0.0128672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_33_131#_c_291_n 0.0194298f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.045
cc_27 VNB N_A_33_131#_c_292_n 0.0410815f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.577
cc_28 VNB N_A_33_131#_c_293_n 0.0236857f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.577
cc_29 VNB N_A_33_131#_c_294_n 0.0142555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_33_131#_c_295_n 0.00397538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_33_131#_c_296_n 0.00956297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_33_131#_c_297_n 0.00816974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_376_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_409_n 0.00303382f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_VGND_c_444_n 0.0165009f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.51
cc_36 VNB N_VGND_c_445_n 0.00576457f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.577
cc_37 VNB N_VGND_c_446_n 4.03531e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_447_n 0.0187954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_448_n 0.0154314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_449_n 0.0146425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_450_n 0.0159488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_451_n 0.196464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_452_n 0.00720971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_453_n 0.00648074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_454_n 0.00436966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_C_N_c_78_n 0.0208401f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.725
cc_47 VPB N_C_N_c_76_n 0.0142025f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.51
cc_48 VPB N_C_N_c_77_n 0.017394f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.535
cc_49 VPB N_A_195_21#_M1006_g 0.0213356f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.577
cc_50 VPB N_A_195_21#_M1010_g 0.0222614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_195_21#_c_109_n 0.0262894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_M1000_g 0.0229278f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.045
cc_53 VPB N_A_c_203_n 0.00634839f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.725
cc_54 VPB N_A_c_204_n 0.00319652f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.577
cc_55 VPB N_B_M1008_g 0.0191703f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_56 VPB N_A_33_131#_M1009_g 0.0365425f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.535
cc_57 VPB N_A_33_131#_c_292_n 4.00125e-19 $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.577
cc_58 VPB N_A_33_131#_c_300_n 0.0282908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_33_131#_c_297_n 0.00295073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_33_131#_c_302_n 0.0105332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_33_131#_c_303_n 0.00722989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_33_131#_c_304_n 0.0446786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_33_131#_c_305_n 0.0637715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_377_n 0.0204989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_378_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.51
cc_66 VPB N_VPWR_c_379_n 0.010221f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.577
cc_67 VPB N_VPWR_c_380_n 0.0280782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_381_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.577
cc_69 VPB N_VPWR_c_382_n 0.0427613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_376_n 0.107468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_384_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_X_c_409_n 0.00111556f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_73 VPB N_X_c_411_n 0.00558857f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.51
cc_74 N_C_N_M1004_g N_A_195_21#_c_99_n 0.0150661f $X=0.505 $Y=0.865 $X2=0 $Y2=0
cc_75 N_C_N_c_77_n N_A_195_21#_M1006_g 0.0250283f $X=0.505 $Y=1.535 $X2=0 $Y2=0
cc_76 N_C_N_M1004_g N_A_195_21#_c_104_n 0.00197756f $X=0.505 $Y=0.865 $X2=0
+ $Y2=0
cc_77 N_C_N_M1004_g N_A_33_131#_c_295_n 0.0157252f $X=0.505 $Y=0.865 $X2=0 $Y2=0
cc_78 N_C_N_c_76_n N_A_33_131#_c_295_n 0.014106f $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_79 N_C_N_c_77_n N_A_33_131#_c_295_n 0.00673603f $X=0.505 $Y=1.535 $X2=0 $Y2=0
cc_80 N_C_N_c_76_n N_A_33_131#_c_296_n 0.022044f $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_81 N_C_N_c_77_n N_A_33_131#_c_296_n 0.0037027f $X=0.505 $Y=1.535 $X2=0 $Y2=0
cc_82 N_C_N_M1004_g N_A_33_131#_c_297_n 0.00392057f $X=0.505 $Y=0.865 $X2=0
+ $Y2=0
cc_83 N_C_N_c_76_n N_A_33_131#_c_297_n 0.0269441f $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_84 N_C_N_c_77_n N_A_33_131#_c_297_n 0.00534141f $X=0.505 $Y=1.535 $X2=0 $Y2=0
cc_85 N_C_N_c_78_n N_A_33_131#_c_304_n 0.0236486f $X=0.67 $Y=1.725 $X2=0 $Y2=0
cc_86 N_C_N_c_76_n N_A_33_131#_c_304_n 0.0229258f $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_87 N_C_N_c_77_n N_A_33_131#_c_304_n 0.00196114f $X=0.505 $Y=1.535 $X2=0 $Y2=0
cc_88 N_C_N_M1004_g X 5.23494e-19 $X=0.505 $Y=0.865 $X2=0 $Y2=0
cc_89 N_C_N_M1004_g N_VGND_c_444_n 0.012423f $X=0.505 $Y=0.865 $X2=0 $Y2=0
cc_90 N_C_N_M1004_g N_VGND_c_447_n 0.00332367f $X=0.505 $Y=0.865 $X2=0 $Y2=0
cc_91 N_C_N_M1004_g N_VGND_c_451_n 0.00387424f $X=0.505 $Y=0.865 $X2=0 $Y2=0
cc_92 N_A_195_21#_c_101_n N_A_M1011_g 0.0207887f $X=1.48 $Y=1.185 $X2=0 $Y2=0
cc_93 N_A_195_21#_c_103_n N_A_M1011_g 0.00231261f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_94 N_A_195_21#_c_104_n N_A_M1011_g 0.00873853f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_95 N_A_195_21#_c_105_n N_A_M1011_g 0.0152451f $X=2.1 $Y=1.15 $X2=0 $Y2=0
cc_96 N_A_195_21#_c_106_n N_A_M1011_g 0.00106123f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_195_21#_c_110_n N_A_M1011_g 0.00597694f $X=2.207 $Y=0.87 $X2=0 $Y2=0
cc_98 N_A_195_21#_M1010_g N_A_M1000_g 0.0232899f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_195_21#_c_103_n N_A_c_203_n 0.00228987f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_100 N_A_195_21#_c_104_n N_A_c_203_n 0.0205679f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_101 N_A_195_21#_c_105_n N_A_c_203_n 0.00102782f $X=2.1 $Y=1.15 $X2=0 $Y2=0
cc_102 N_A_195_21#_c_110_n N_A_c_203_n 0.00414616f $X=2.207 $Y=0.87 $X2=0 $Y2=0
cc_103 N_A_195_21#_M1010_g N_A_c_204_n 0.00496036f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_195_21#_c_103_n N_A_c_204_n 0.00691778f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_105 N_A_195_21#_c_105_n N_A_c_204_n 0.0133f $X=2.1 $Y=1.15 $X2=0 $Y2=0
cc_106 N_A_195_21#_c_110_n N_A_c_204_n 0.0170371f $X=2.207 $Y=0.87 $X2=0 $Y2=0
cc_107 N_A_195_21#_c_106_n N_B_c_245_n 0.00184315f $X=2.22 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_108 N_A_195_21#_c_109_n N_B_M1008_g 7.85336e-19 $X=3.1 $Y=2.135 $X2=0 $Y2=0
cc_109 N_A_195_21#_c_107_n N_B_c_247_n 0.0103633f $X=2.985 $Y=0.87 $X2=0 $Y2=0
cc_110 N_A_195_21#_c_107_n B 0.0267022f $X=2.985 $Y=0.87 $X2=0 $Y2=0
cc_111 N_A_195_21#_c_109_n B 0.071529f $X=3.1 $Y=2.135 $X2=0 $Y2=0
cc_112 N_A_195_21#_c_110_n B 0.00929532f $X=2.207 $Y=0.87 $X2=0 $Y2=0
cc_113 N_A_195_21#_c_107_n N_B_c_249_n 0.00126891f $X=2.985 $Y=0.87 $X2=0 $Y2=0
cc_114 N_A_195_21#_c_109_n N_B_c_249_n 9.97443e-19 $X=3.1 $Y=2.135 $X2=0 $Y2=0
cc_115 N_A_195_21#_c_107_n N_B_c_250_n 0.00477414f $X=2.985 $Y=0.87 $X2=0 $Y2=0
cc_116 N_A_195_21#_c_109_n N_B_c_250_n 0.00367226f $X=3.1 $Y=2.135 $X2=0 $Y2=0
cc_117 N_A_195_21#_c_110_n N_B_c_250_n 0.00524568f $X=2.207 $Y=0.87 $X2=0 $Y2=0
cc_118 N_A_195_21#_c_108_n N_A_33_131#_c_291_n 0.00359736f $X=3.1 $Y=0.445 $X2=0
+ $Y2=0
cc_119 N_A_195_21#_c_109_n N_A_33_131#_M1009_g 0.00281739f $X=3.1 $Y=2.135 $X2=0
+ $Y2=0
cc_120 N_A_195_21#_c_109_n N_A_33_131#_c_292_n 0.0240653f $X=3.1 $Y=2.135 $X2=0
+ $Y2=0
cc_121 N_A_195_21#_c_111_n N_A_33_131#_c_292_n 0.00117977f $X=3.125 $Y=0.87
+ $X2=0 $Y2=0
cc_122 N_A_195_21#_c_107_n N_A_33_131#_c_293_n 0.00965738f $X=2.985 $Y=0.87
+ $X2=0 $Y2=0
cc_123 N_A_195_21#_c_108_n N_A_33_131#_c_293_n 0.00509979f $X=3.1 $Y=0.445 $X2=0
+ $Y2=0
cc_124 N_A_195_21#_c_111_n N_A_33_131#_c_293_n 0.00520416f $X=3.125 $Y=0.87
+ $X2=0 $Y2=0
cc_125 N_A_195_21#_c_109_n N_A_33_131#_c_300_n 0.0119065f $X=3.1 $Y=2.135 $X2=0
+ $Y2=0
cc_126 N_A_195_21#_c_99_n N_A_33_131#_c_295_n 0.00172885f $X=1.05 $Y=1.185 $X2=0
+ $Y2=0
cc_127 N_A_195_21#_M1006_g N_A_33_131#_c_297_n 3.42426e-19 $X=1.195 $Y=2.465
+ $X2=0 $Y2=0
cc_128 N_A_195_21#_c_104_n N_A_33_131#_c_297_n 0.0027848f $X=1.535 $Y=1.355
+ $X2=0 $Y2=0
cc_129 N_A_195_21#_M1006_g N_A_33_131#_c_302_n 0.0154434f $X=1.195 $Y=2.465
+ $X2=0 $Y2=0
cc_130 N_A_195_21#_M1010_g N_A_33_131#_c_302_n 0.0186874f $X=1.625 $Y=2.465
+ $X2=0 $Y2=0
cc_131 N_A_195_21#_M1006_g N_A_33_131#_c_304_n 0.00544648f $X=1.195 $Y=2.465
+ $X2=0 $Y2=0
cc_132 N_A_195_21#_M1006_g N_VPWR_c_377_n 0.0157379f $X=1.195 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_195_21#_M1010_g N_VPWR_c_377_n 0.00176668f $X=1.625 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_195_21#_M1006_g N_VPWR_c_378_n 0.00486043f $X=1.195 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_195_21#_M1010_g N_VPWR_c_378_n 0.00486043f $X=1.625 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_195_21#_M1006_g N_VPWR_c_379_n 0.00176668f $X=1.195 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_195_21#_M1010_g N_VPWR_c_379_n 0.0157379f $X=1.625 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_A_195_21#_M1006_g N_VPWR_c_376_n 0.00835506f $X=1.195 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_195_21#_M1010_g N_VPWR_c_376_n 0.00835506f $X=1.625 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_195_21#_c_99_n N_X_c_409_n 0.00328059f $X=1.05 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A_195_21#_M1006_g N_X_c_409_n 0.0102891f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_195_21#_c_101_n N_X_c_409_n 0.00192984f $X=1.48 $Y=1.185 $X2=0 $Y2=0
cc_143 N_A_195_21#_M1010_g N_X_c_409_n 0.00118583f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_195_21#_c_103_n N_X_c_409_n 0.0200502f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_145 N_A_195_21#_c_104_n N_X_c_409_n 0.0139562f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_146 N_A_195_21#_c_172_p N_X_c_409_n 0.0102238f $X=1.72 $Y=1.15 $X2=0 $Y2=0
cc_147 N_A_195_21#_M1006_g N_X_c_411_n 0.00870978f $X=1.195 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_195_21#_M1010_g N_X_c_411_n 0.0053094f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_195_21#_c_103_n N_X_c_411_n 0.0069428f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_150 N_A_195_21#_c_104_n N_X_c_411_n 0.00328837f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_151 N_A_195_21#_c_99_n N_X_c_424_n 0.00703996f $X=1.05 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A_195_21#_c_99_n X 0.00239543f $X=1.05 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A_195_21#_c_104_n X 0.00216562f $X=1.535 $Y=1.355 $X2=0 $Y2=0
cc_154 N_A_195_21#_c_105_n N_VGND_M1007_s 0.00105239f $X=2.1 $Y=1.15 $X2=0 $Y2=0
cc_155 N_A_195_21#_c_172_p N_VGND_M1007_s 0.00116967f $X=1.72 $Y=1.15 $X2=0
+ $Y2=0
cc_156 N_A_195_21#_c_99_n N_VGND_c_444_n 0.00507914f $X=1.05 $Y=1.185 $X2=0
+ $Y2=0
cc_157 N_A_195_21#_c_99_n N_VGND_c_445_n 6.79059e-19 $X=1.05 $Y=1.185 $X2=0
+ $Y2=0
cc_158 N_A_195_21#_c_101_n N_VGND_c_445_n 0.0163601f $X=1.48 $Y=1.185 $X2=0
+ $Y2=0
cc_159 N_A_195_21#_c_104_n N_VGND_c_445_n 7.06489e-19 $X=1.535 $Y=1.355 $X2=0
+ $Y2=0
cc_160 N_A_195_21#_c_105_n N_VGND_c_445_n 0.0173055f $X=2.1 $Y=1.15 $X2=0 $Y2=0
cc_161 N_A_195_21#_c_172_p N_VGND_c_445_n 0.010804f $X=1.72 $Y=1.15 $X2=0 $Y2=0
cc_162 N_A_195_21#_c_106_n N_VGND_c_445_n 0.0231513f $X=2.22 $Y=0.445 $X2=0
+ $Y2=0
cc_163 N_A_195_21#_c_110_n N_VGND_c_445_n 0.00985927f $X=2.207 $Y=0.87 $X2=0
+ $Y2=0
cc_164 N_A_195_21#_c_107_n N_VGND_c_446_n 0.0207225f $X=2.985 $Y=0.87 $X2=0
+ $Y2=0
cc_165 N_A_195_21#_c_99_n N_VGND_c_448_n 0.0054895f $X=1.05 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A_195_21#_c_101_n N_VGND_c_448_n 0.00486043f $X=1.48 $Y=1.185 $X2=0
+ $Y2=0
cc_167 N_A_195_21#_c_106_n N_VGND_c_449_n 0.0115062f $X=2.22 $Y=0.445 $X2=0
+ $Y2=0
cc_168 N_A_195_21#_c_108_n N_VGND_c_450_n 0.0159678f $X=3.1 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_195_21#_M1011_d N_VGND_c_451_n 0.00324303f $X=2.08 $Y=0.235 $X2=0
+ $Y2=0
cc_170 N_A_195_21#_M1005_d N_VGND_c_451_n 0.00230518f $X=2.96 $Y=0.235 $X2=0
+ $Y2=0
cc_171 N_A_195_21#_c_99_n N_VGND_c_451_n 0.0110654f $X=1.05 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A_195_21#_c_101_n N_VGND_c_451_n 0.00824727f $X=1.48 $Y=1.185 $X2=0
+ $Y2=0
cc_173 N_A_195_21#_c_106_n N_VGND_c_451_n 0.0081803f $X=2.22 $Y=0.445 $X2=0
+ $Y2=0
cc_174 N_A_195_21#_c_107_n N_VGND_c_451_n 0.0114207f $X=2.985 $Y=0.87 $X2=0
+ $Y2=0
cc_175 N_A_195_21#_c_108_n N_VGND_c_451_n 0.0106767f $X=3.1 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A_M1011_g N_B_c_245_n 0.0175141f $X=2.005 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_177 N_A_M1000_g N_B_M1008_g 0.03469f $X=2.165 $Y=2.135 $X2=0 $Y2=0
cc_178 N_A_M1011_g B 7.12363e-19 $X=2.005 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A_c_203_n B 0.00127117f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_c_204_n B 0.0555729f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A_c_203_n N_B_c_249_n 0.03469f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_c_204_n N_B_c_249_n 0.00383853f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A_M1011_g N_B_c_250_n 0.0124006f $X=2.005 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_M1000_g N_A_33_131#_c_302_n 0.0139483f $X=2.165 $Y=2.135 $X2=0 $Y2=0
cc_185 N_A_c_203_n N_A_33_131#_c_302_n 4.50807e-19 $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A_c_204_n N_A_33_131#_c_302_n 0.0219613f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_187 N_A_c_204_n N_VPWR_M1010_d 0.0046277f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A_M1000_g N_VPWR_c_376_n 0.00380473f $X=2.165 $Y=2.135 $X2=0 $Y2=0
cc_189 N_A_c_203_n N_X_c_409_n 2.34898e-19 $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A_c_204_n N_X_c_409_n 0.00761998f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A_M1000_g N_X_c_411_n 2.60816e-19 $X=2.165 $Y=2.135 $X2=0 $Y2=0
cc_192 N_A_c_204_n N_X_c_411_n 0.0146288f $X=2.075 $Y=1.51 $X2=0 $Y2=0
cc_193 N_A_c_204_n A_448_385# 0.00173922f $X=2.075 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_194 N_A_M1011_g N_VGND_c_445_n 0.00463887f $X=2.005 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A_M1011_g N_VGND_c_446_n 6.00618e-19 $X=2.005 $Y=0.445 $X2=0 $Y2=0
cc_196 N_A_M1011_g N_VGND_c_449_n 0.00583607f $X=2.005 $Y=0.445 $X2=0 $Y2=0
cc_197 N_A_M1011_g N_VGND_c_451_n 0.0108595f $X=2.005 $Y=0.445 $X2=0 $Y2=0
cc_198 N_B_c_245_n N_A_33_131#_c_291_n 0.0107318f $X=2.435 $Y=0.765 $X2=0 $Y2=0
cc_199 B N_A_33_131#_M1009_g 0.00556915f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_200 N_B_M1008_g N_A_33_131#_c_292_n 0.00306742f $X=2.525 $Y=2.135 $X2=0 $Y2=0
cc_201 B N_A_33_131#_c_292_n 0.00147055f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_202 N_B_c_249_n N_A_33_131#_c_292_n 0.018078f $X=2.615 $Y=1.29 $X2=0 $Y2=0
cc_203 N_B_c_250_n N_A_33_131#_c_292_n 0.00288958f $X=2.615 $Y=1.125 $X2=0 $Y2=0
cc_204 N_B_c_247_n N_A_33_131#_c_293_n 0.0097334f $X=2.525 $Y=0.84 $X2=0 $Y2=0
cc_205 N_B_M1008_g N_A_33_131#_c_300_n 0.0517096f $X=2.525 $Y=2.135 $X2=0 $Y2=0
cc_206 B N_A_33_131#_c_300_n 0.00353467f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_207 N_B_M1008_g N_A_33_131#_c_302_n 0.00955848f $X=2.525 $Y=2.135 $X2=0 $Y2=0
cc_208 B N_A_33_131#_c_302_n 0.0193702f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_209 N_B_M1008_g N_A_33_131#_c_303_n 0.00165504f $X=2.525 $Y=2.135 $X2=0 $Y2=0
cc_210 N_B_M1008_g N_A_33_131#_c_305_n 0.00636429f $X=2.525 $Y=2.135 $X2=0 $Y2=0
cc_211 B N_A_33_131#_c_305_n 5.90859e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_212 N_B_M1008_g N_VPWR_c_376_n 8.89433e-19 $X=2.525 $Y=2.135 $X2=0 $Y2=0
cc_213 B A_520_385# 9.70164e-19 $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_214 N_B_c_245_n N_VGND_c_446_n 0.00845795f $X=2.435 $Y=0.765 $X2=0 $Y2=0
cc_215 N_B_c_247_n N_VGND_c_446_n 0.002329f $X=2.525 $Y=0.84 $X2=0 $Y2=0
cc_216 N_B_c_245_n N_VGND_c_449_n 0.00486043f $X=2.435 $Y=0.765 $X2=0 $Y2=0
cc_217 N_B_c_245_n N_VGND_c_451_n 0.00453118f $X=2.435 $Y=0.765 $X2=0 $Y2=0
cc_218 N_A_33_131#_c_297_n N_VPWR_M1002_d 0.00111036f $X=0.84 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A_33_131#_c_302_n N_VPWR_M1002_d 0.00655748f $X=2.485 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_220 N_A_33_131#_c_304_n N_VPWR_M1002_d 0.00544769f $X=0.93 $Y=2.19 $X2=-0.19
+ $Y2=-0.245
cc_221 N_A_33_131#_c_302_n N_VPWR_M1010_d 0.00961011f $X=2.485 $Y=2.375 $X2=0
+ $Y2=0
cc_222 N_A_33_131#_c_304_n N_VPWR_c_377_n 0.0217712f $X=0.93 $Y=2.19 $X2=0 $Y2=0
cc_223 N_A_33_131#_c_302_n N_VPWR_c_379_n 0.021083f $X=2.485 $Y=2.375 $X2=0
+ $Y2=0
cc_224 N_A_33_131#_c_303_n N_VPWR_c_379_n 0.0121534f $X=2.65 $Y=2.88 $X2=0 $Y2=0
cc_225 N_A_33_131#_c_305_n N_VPWR_c_379_n 0.00732408f $X=2.885 $Y=2.88 $X2=0
+ $Y2=0
cc_226 N_A_33_131#_c_303_n N_VPWR_c_382_n 0.01284f $X=2.65 $Y=2.88 $X2=0 $Y2=0
cc_227 N_A_33_131#_c_305_n N_VPWR_c_382_n 0.0125969f $X=2.885 $Y=2.88 $X2=0
+ $Y2=0
cc_228 N_A_33_131#_c_303_n N_VPWR_c_376_n 0.0117243f $X=2.65 $Y=2.88 $X2=0 $Y2=0
cc_229 N_A_33_131#_c_305_n N_VPWR_c_376_n 0.0155249f $X=2.885 $Y=2.88 $X2=0
+ $Y2=0
cc_230 N_A_33_131#_c_302_n N_X_M1006_s 0.00810274f $X=2.485 $Y=2.375 $X2=0 $Y2=0
cc_231 N_A_33_131#_c_295_n N_X_c_409_n 0.0131672f $X=0.75 $Y=1.15 $X2=0 $Y2=0
cc_232 N_A_33_131#_c_297_n N_X_c_409_n 0.0434407f $X=0.84 $Y=1.92 $X2=0 $Y2=0
cc_233 N_A_33_131#_c_297_n N_X_c_411_n 0.00464704f $X=0.84 $Y=1.92 $X2=0 $Y2=0
cc_234 N_A_33_131#_c_302_n N_X_c_411_n 0.0249186f $X=2.485 $Y=2.375 $X2=0 $Y2=0
cc_235 N_A_33_131#_c_302_n A_448_385# 0.00347026f $X=2.485 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_33_131#_c_302_n A_520_385# 0.00106212f $X=2.485 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_237 N_A_33_131#_c_295_n N_VGND_M1004_d 0.00313716f $X=0.75 $Y=1.15 $X2=-0.19
+ $Y2=-0.245
cc_238 N_A_33_131#_c_295_n N_VGND_c_444_n 0.0260903f $X=0.75 $Y=1.15 $X2=0 $Y2=0
cc_239 N_A_33_131#_c_291_n N_VGND_c_446_n 0.00915651f $X=2.885 $Y=0.765 $X2=0
+ $Y2=0
cc_240 N_A_33_131#_c_294_n N_VGND_c_447_n 0.00421179f $X=0.29 $Y=0.865 $X2=0
+ $Y2=0
cc_241 N_A_33_131#_c_291_n N_VGND_c_450_n 0.00564095f $X=2.885 $Y=0.765 $X2=0
+ $Y2=0
cc_242 N_A_33_131#_c_293_n N_VGND_c_450_n 8.13583e-19 $X=3.095 $Y=0.84 $X2=0
+ $Y2=0
cc_243 N_A_33_131#_c_291_n N_VGND_c_451_n 0.0061326f $X=2.885 $Y=0.765 $X2=0
+ $Y2=0
cc_244 N_A_33_131#_c_293_n N_VGND_c_451_n 5.53504e-19 $X=3.095 $Y=0.84 $X2=0
+ $Y2=0
cc_245 N_A_33_131#_c_294_n N_VGND_c_451_n 0.00737625f $X=0.29 $Y=0.865 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_376_n N_X_M1006_s 0.0119922f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_247 N_X_c_424_n N_VGND_c_448_n 0.015688f $X=1.265 $Y=0.42 $X2=0 $Y2=0
cc_248 N_X_M1001_d N_VGND_c_451_n 0.00380103f $X=1.125 $Y=0.235 $X2=0 $Y2=0
cc_249 N_X_c_424_n N_VGND_c_451_n 0.00984745f $X=1.265 $Y=0.42 $X2=0 $Y2=0
