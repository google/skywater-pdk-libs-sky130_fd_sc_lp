* File: sky130_fd_sc_lp__nor3b_2.spice
* Created: Fri Aug 28 10:56:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor3b_2.pex.spice"
.subckt sky130_fd_sc_lp__nor3b_2  VNB VPB C_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_C_N_M1012_g N_A_27_131#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1575 AS=0.1113 PD=1.13333 PS=1.37 NRD=91.428 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1012_d N_A_27_131#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.315 AS=0.1617 PD=2.26667 PS=1.225 NRD=0 NRS=8.568 M=1 R=5.6 SA=75000.7
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_27_131#_M1004_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1554 AS=0.1617 PD=1.21 PS=1.225 NRD=7.14 NRS=6.42 M=1 R=5.6 SA=75001.2
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1004_d N_B_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1554
+ AS=0.1176 PD=1.21 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75001.7 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_B_M1007_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.2 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.6 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1011 N_Y_M1005_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_C_N_M1001_g N_A_27_131#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_217_365#_M1006_d N_A_27_131#_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1009 N_A_217_365#_M1009_d N_A_27_131#_M1009_g N_Y_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1002 N_A_472_365#_M1002_d N_B_M1002_g N_A_217_365#_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_472_365#_M1002_d N_B_M1010_g N_A_217_365#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_A_472_365#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_472_365#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.684 P=14.11
*
.include "sky130_fd_sc_lp__nor3b_2.pxi.spice"
*
.ends
*
*
