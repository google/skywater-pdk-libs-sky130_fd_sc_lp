* File: sky130_fd_sc_lp__nor3_0.pxi.spice
* Created: Fri Aug 28 10:55:07 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3_0%A N_A_c_49_n N_A_M1002_g N_A_c_56_n N_A_M1000_g
+ N_A_c_50_n N_A_c_51_n N_A_c_52_n N_A_c_57_n A A A A N_A_c_54_n
+ PM_SKY130_FD_SC_LP__NOR3_0%A
x_PM_SKY130_FD_SC_LP__NOR3_0%B N_B_M1001_g N_B_M1003_g N_B_c_91_n N_B_c_96_n B B
+ B B B N_B_c_93_n B PM_SKY130_FD_SC_LP__NOR3_0%B
x_PM_SKY130_FD_SC_LP__NOR3_0%C N_C_M1005_g N_C_M1004_g N_C_c_145_n N_C_c_150_n C
+ C C N_C_c_147_n PM_SKY130_FD_SC_LP__NOR3_0%C
x_PM_SKY130_FD_SC_LP__NOR3_0%VPWR N_VPWR_M1000_s N_VPWR_c_180_n N_VPWR_c_181_n
+ VPWR N_VPWR_c_182_n N_VPWR_c_179_n PM_SKY130_FD_SC_LP__NOR3_0%VPWR
x_PM_SKY130_FD_SC_LP__NOR3_0%Y N_Y_M1002_d N_Y_M1004_d N_Y_M1005_d N_Y_c_199_n
+ N_Y_c_200_n N_Y_c_205_n N_Y_c_201_n Y Y Y N_Y_c_203_n N_Y_c_204_n
+ PM_SKY130_FD_SC_LP__NOR3_0%Y
x_PM_SKY130_FD_SC_LP__NOR3_0%VGND N_VGND_M1002_s N_VGND_M1001_d N_VGND_c_241_n
+ N_VGND_c_242_n N_VGND_c_243_n VGND N_VGND_c_244_n N_VGND_c_245_n
+ N_VGND_c_246_n N_VGND_c_247_n PM_SKY130_FD_SC_LP__NOR3_0%VGND
cc_1 VNB N_A_c_49_n 0.00799035f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.155
cc_2 VNB N_A_c_50_n 0.0211236f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.855
cc_3 VNB N_A_c_51_n 0.0305908f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_4 VNB N_A_c_52_n 0.0185667f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_5 VNB A 0.033577f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A_c_54_n 0.0303222f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_7 VNB N_B_M1001_g 0.0364772f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.855
cc_8 VNB N_B_c_91_n 0.0154103f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_9 VNB B 0.00528862f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_10 VNB N_B_c_93_n 0.0155587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_M1004_g 0.0420812f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.735
cc_12 VNB N_C_c_145_n 0.0191071f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_13 VNB C 0.00467826f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_14 VNB N_C_c_147_n 0.016229f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_VPWR_c_179_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.23
cc_16 VNB N_Y_c_199_n 0.00390632f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.855
cc_17 VNB N_Y_c_200_n 8.38975e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.36
cc_18 VNB N_Y_c_201_n 0.0299162f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_19 VNB Y 0.0141514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_203_n 0.00928982f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_21 VNB N_Y_c_204_n 0.0224461f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=1.295
cc_22 VNB N_VGND_c_241_n 0.0118455f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.735
cc_23 VNB N_VGND_c_242_n 0.020607f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_24 VNB N_VGND_c_243_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_25 VNB N_VGND_c_244_n 0.0144674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_245_n 0.0184227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_246_n 0.133181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_247_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_A_c_49_n 0.0323458f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.155
cc_30 VPB N_A_c_56_n 0.0213851f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.305
cc_31 VPB N_A_c_57_n 0.0272706f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.23
cc_32 VPB A 0.0248792f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_33 VPB N_B_M1003_g 0.0346294f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.735
cc_34 VPB N_B_c_91_n 0.00593676f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.005
cc_35 VPB N_B_c_96_n 0.0156011f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.36
cc_36 VPB B 0.00230661f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.525
cc_37 VPB B 0.00150533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB B 0.00190145f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.23
cc_39 VPB N_C_M1005_g 0.0448772f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.855
cc_40 VPB N_C_c_145_n 0.00404058f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.005
cc_41 VPB N_C_c_150_n 0.0168167f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.36
cc_42 VPB C 0.0129487f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.525
cc_43 VPB N_VPWR_c_180_n 0.0131454f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.535
cc_44 VPB N_VPWR_c_181_n 0.0353237f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.305
cc_45 VPB N_VPWR_c_182_n 0.0423956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_179_n 0.0614348f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.23
cc_47 VPB N_Y_c_205_n 0.0391258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_Y_c_201_n 0.0362803f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_49 N_A_c_50_n N_B_M1001_g 0.0178694f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_50 A N_B_M1001_g 0.00107052f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_51 N_A_c_54_n N_B_M1001_g 0.00702299f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_52 N_A_c_49_n N_B_M1003_g 0.00540078f $X=0.36 $Y=2.155 $X2=0 $Y2=0
cc_53 N_A_c_57_n N_B_M1003_g 0.0531007f $X=0.54 $Y=2.23 $X2=0 $Y2=0
cc_54 A N_B_M1003_g 2.28296e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_55 N_A_c_52_n N_B_c_91_n 0.0113126f $X=0.27 $Y=1.525 $X2=0 $Y2=0
cc_56 N_A_c_49_n N_B_c_96_n 0.0113126f $X=0.36 $Y=2.155 $X2=0 $Y2=0
cc_57 A B 0.0781988f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A_c_54_n B 0.00312077f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_59 N_A_c_52_n B 0.00312077f $X=0.27 $Y=1.525 $X2=0 $Y2=0
cc_60 N_A_c_57_n B 0.00513027f $X=0.54 $Y=2.23 $X2=0 $Y2=0
cc_61 N_A_c_57_n B 0.00701126f $X=0.54 $Y=2.23 $X2=0 $Y2=0
cc_62 A N_B_c_93_n 6.67555e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A_c_54_n N_B_c_93_n 0.0113126f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_64 N_A_c_56_n N_VPWR_c_181_n 0.0052936f $X=0.54 $Y=2.305 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_VPWR_c_181_n 0.00650559f $X=0.54 $Y=2.23 $X2=0 $Y2=0
cc_66 A N_VPWR_c_181_n 0.0193792f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A_c_56_n N_VPWR_c_182_n 0.00543892f $X=0.54 $Y=2.305 $X2=0 $Y2=0
cc_68 N_A_c_56_n N_VPWR_c_179_n 0.010971f $X=0.54 $Y=2.305 $X2=0 $Y2=0
cc_69 N_A_c_50_n N_Y_c_199_n 0.00306602f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_70 A N_Y_c_199_n 0.0160684f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_71 N_A_c_54_n N_Y_c_199_n 3.18588e-19 $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_72 N_A_c_50_n N_Y_c_200_n 0.00115611f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_73 N_A_c_50_n N_VGND_c_242_n 0.01027f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_74 N_A_c_51_n N_VGND_c_242_n 0.00201721f $X=0.34 $Y=1.005 $X2=0 $Y2=0
cc_75 A N_VGND_c_242_n 0.0238221f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A_c_50_n N_VGND_c_243_n 5.37826e-19 $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_77 N_A_c_50_n N_VGND_c_244_n 0.00414769f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_78 N_A_c_50_n N_VGND_c_246_n 0.0078848f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_79 A N_VGND_c_246_n 0.00241005f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_B_c_96_n N_C_M1005_g 0.0661145f $X=0.84 $Y=1.915 $X2=0 $Y2=0
cc_81 B N_C_M1005_g 2.7465e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 B N_C_M1005_g 0.00247266f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_83 N_B_M1001_g N_C_M1004_g 0.0283358f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_84 N_B_c_93_n N_C_c_145_n 0.0137354f $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B_c_91_n N_C_c_150_n 0.0137354f $X=0.84 $Y=1.75 $X2=0 $Y2=0
cc_86 N_B_M1001_g C 0.00656284f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_87 B C 0.0792053f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_M1001_g N_C_c_147_n 0.0137354f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_89 B N_C_c_147_n 5.8273e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 B N_VPWR_c_181_n 0.0190316f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_91 N_B_M1003_g N_VPWR_c_182_n 0.00464216f $X=0.93 $Y=2.735 $X2=0 $Y2=0
cc_92 B N_VPWR_c_182_n 0.00697579f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_93 N_B_M1003_g N_VPWR_c_179_n 0.00797501f $X=0.93 $Y=2.735 $X2=0 $Y2=0
cc_94 B N_VPWR_c_179_n 0.00949194f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_95 B A_123_483# 0.0019099f $X=0.635 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_96 N_B_M1001_g N_Y_c_199_n 7.00936e-19 $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_97 B N_Y_c_199_n 0.0216254f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_98 N_B_c_93_n N_Y_c_199_n 9.55128e-19 $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B_M1001_g N_Y_c_200_n 6.75895e-19 $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_100 N_B_M1003_g N_Y_c_205_n 0.00229434f $X=0.93 $Y=2.735 $X2=0 $Y2=0
cc_101 B N_Y_c_205_n 0.0162797f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_102 N_B_M1001_g N_Y_c_203_n 0.0153698f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_103 B N_Y_c_203_n 0.00911953f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B_c_93_n N_Y_c_203_n 2.85404e-19 $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B_M1001_g N_VGND_c_242_n 5.37826e-19 $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_106 N_B_M1001_g N_VGND_c_243_n 0.00828067f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_107 N_B_M1001_g N_VGND_c_244_n 0.00414769f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_108 N_B_M1001_g N_VGND_c_246_n 0.00414907f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_109 N_C_M1005_g N_VPWR_c_182_n 0.00511657f $X=1.32 $Y=2.735 $X2=0 $Y2=0
cc_110 N_C_M1005_g N_VPWR_c_179_n 0.0103852f $X=1.32 $Y=2.735 $X2=0 $Y2=0
cc_111 N_C_M1005_g N_Y_c_205_n 0.0122847f $X=1.32 $Y=2.735 $X2=0 $Y2=0
cc_112 N_C_c_150_n N_Y_c_205_n 0.00296106f $X=1.38 $Y=1.88 $X2=0 $Y2=0
cc_113 C N_Y_c_205_n 0.00767352f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_C_M1005_g N_Y_c_201_n 0.00661148f $X=1.32 $Y=2.735 $X2=0 $Y2=0
cc_115 N_C_M1004_g N_Y_c_201_n 0.00403827f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_116 C N_Y_c_201_n 0.0772501f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_C_c_147_n N_Y_c_201_n 0.0165356f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_118 N_C_c_147_n Y 0.00309682f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_119 N_C_M1004_g N_Y_c_203_n 0.0147349f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_120 C N_Y_c_203_n 0.0297242f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_121 N_C_c_147_n N_Y_c_203_n 0.00134773f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_122 N_C_M1004_g N_Y_c_204_n 0.00321699f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_123 N_C_M1004_g N_VGND_c_243_n 0.0119778f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_124 N_C_M1004_g N_VGND_c_245_n 0.00414769f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_125 N_C_M1004_g N_VGND_c_246_n 0.00452535f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_126 N_VPWR_c_182_n N_Y_c_205_n 0.0311147f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_127 N_VPWR_c_179_n N_Y_c_205_n 0.0178003f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_128 N_Y_c_203_n N_VGND_c_243_n 0.0213027f $X=1.48 $Y=0.94 $X2=0 $Y2=0
cc_129 N_Y_c_200_n N_VGND_c_244_n 0.00726487f $X=0.715 $Y=0.53 $X2=0 $Y2=0
cc_130 N_Y_c_204_n N_VGND_c_245_n 0.0143843f $X=1.575 $Y=0.53 $X2=0 $Y2=0
cc_131 N_Y_c_199_n N_VGND_c_246_n 0.00168524f $X=0.715 $Y=0.79 $X2=0 $Y2=0
cc_132 N_Y_c_200_n N_VGND_c_246_n 0.00687863f $X=0.715 $Y=0.53 $X2=0 $Y2=0
cc_133 N_Y_c_203_n N_VGND_c_246_n 0.0111883f $X=1.48 $Y=0.94 $X2=0 $Y2=0
cc_134 N_Y_c_204_n N_VGND_c_246_n 0.0129176f $X=1.575 $Y=0.53 $X2=0 $Y2=0
