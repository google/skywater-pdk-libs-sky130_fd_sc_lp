* File: sky130_fd_sc_lp__dfrtp_1.spice
* Created: Wed Sep  2 09:43:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfrtp_1.pex.spice"
.subckt sky130_fd_sc_lp__dfrtp_1  VNB VPB CLK D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_CLK_M1013_g N_A_27_114#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.1113 PD=0.97 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1026 N_A_196_462#_M1026_d N_A_27_114#_M1026_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1155 PD=1.37 PS=0.97 NRD=0 NRS=77.136 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 A_492_149# N_RESET_B_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_304_533#_M1002_d N_D_M1002_g A_492_149# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_559_533#_M1004_d N_A_27_114#_M1004_g N_A_304_533#_M1002_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.12915 AS=0.0588 PD=1.035 PS=0.7 NRD=82.848 NRS=0 M=1 R=2.8
+ SA=75001 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1027 A_803_149# N_A_196_462#_M1027_g N_A_559_533#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.12915 PD=0.63 PS=1.035 NRD=14.28 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1018 A_875_149# N_A_695_375#_M1018_g A_803_149# VNB NSHORT L=0.15 W=0.42
+ AD=0.09345 AS=0.0441 PD=1.02 PS=0.63 NRD=47.856 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_RESET_B_M1014_g A_875_149# VNB NSHORT L=0.15 W=0.42
+ AD=0.140423 AS=0.09345 PD=1.05396 PS=1.02 NRD=79.8 NRS=47.856 M=1 R=2.8
+ SA=75001.4 SB=75003 A=0.063 P=1.14 MULT=1
MM1028 N_A_695_375#_M1028_d N_A_559_533#_M1028_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.18205 AS=0.213977 PD=1.28 PS=1.60604 NRD=22.5 NRS=22.5 M=1
+ R=4.26667 SA=75001.5 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1031 N_A_1247_89#_M1031_d N_A_196_462#_M1031_g N_A_695_375#_M1028_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.243925 AS=0.18205 PD=1.61811 PS=1.28 NRD=44.052 NRS=21.552
+ M=1 R=4.26667 SA=75002 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1030 A_1417_133# N_A_27_114#_M1030_g N_A_1247_89#_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.160075 PD=0.72 PS=1.06189 NRD=27.132 NRS=52.848 M=1 R=2.8
+ SA=75003.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_1467_419#_M1000_g A_1417_133# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.063 PD=0.7 PS=0.72 NRD=0 NRS=27.132 M=1 R=2.8 SA=75003.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 A_1593_133# N_RESET_B_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_1467_419#_M1025_d N_A_1247_89#_M1025_g A_1593_133# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_1247_89#_M1017_g N_A_1832_367#_M1017_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0875 AS=0.1113 PD=0.8 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_Q_M1019_d N_A_1832_367#_M1019_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.175 PD=2.21 PS=1.6 NRD=0 NRS=0.708 M=1 R=5.6 SA=75000.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 N_VPWR_M1020_d N_CLK_M1020_g N_A_27_114#_M1020_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_196_462#_M1006_d N_A_27_114#_M1006_g N_VPWR_M1020_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_RESET_B_M1007_g N_A_304_533#_M1007_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1021 N_A_304_533#_M1021_d N_D_M1021_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1015 N_A_559_533#_M1015_d N_A_196_462#_M1015_g N_A_304_533#_M1021_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=18.7544 NRS=0 M=1
+ R=2.8 SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 A_653_533# N_A_27_114#_M1009_g N_A_559_533#_M1015_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1029 N_VPWR_M1029_d N_A_695_375#_M1029_g A_653_533# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.08085 AS=0.0441 PD=0.805 PS=0.63 NRD=37.5088 NRS=23.443 M=1 R=2.8
+ SA=75001.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_A_559_533#_M1022_d N_RESET_B_M1022_g N_VPWR_M1029_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.08085 PD=1.37 PS=0.805 NRD=0 NRS=11.7215 M=1 R=2.8
+ SA=75002.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_695_375#_M1012_d N_A_559_533#_M1012_g N_VPWR_M1012_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1666 AS=0.365 PD=1.245 PS=2.68 NRD=16.4101 NRS=28.1316 M=1
+ R=5.6 SA=75000.3 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1011 N_A_1247_89#_M1011_d N_A_27_114#_M1011_g N_A_695_375#_M1012_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1792 AS=0.1666 PD=1.62 PS=1.245 NRD=0 NRS=10.5395 M=1 R=5.6
+ SA=75000.9 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1005 A_1379_517# N_A_196_462#_M1005_g N_A_1247_89#_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.0896 PD=0.86 PS=0.81 NRD=77.3816 NRS=46.886 M=1 R=2.8
+ SA=75001.4 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_1467_419#_M1016_g A_1379_517# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1155 AS=0.0924 PD=0.97 PS=0.86 NRD=53.9386 NRS=77.3816 M=1 R=2.8
+ SA=75002 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_1467_419#_M1003_d N_RESET_B_M1003_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1155 PD=0.7 PS=0.97 NRD=0 NRS=72.693 M=1 R=2.8
+ SA=75002.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1247_89#_M1008_g N_A_1467_419#_M1003_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_1247_89#_M1023_g N_A_1832_367#_M1023_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.137128 AS=0.1696 PD=1.09137 PS=1.81 NRD=18.4589 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1024 N_Q_M1024_d N_A_1832_367#_M1024_g N_VPWR_M1023_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.269972 PD=3.05 PS=2.14863 NRD=0 NRS=2.3443 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.4031 P=25.61
*
.include "sky130_fd_sc_lp__dfrtp_1.pxi.spice"
*
.ends
*
*
