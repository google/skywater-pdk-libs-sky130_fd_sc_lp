* File: sky130_fd_sc_lp__sdfsbp_2.pxi.spice
* Created: Fri Aug 28 11:29:17 2020
* 
x_PM_SKY130_FD_SC_LP__SDFSBP_2%SCE N_SCE_c_294_n N_SCE_M1029_g N_SCE_M1004_g
+ N_SCE_M1005_g N_SCE_M1011_g N_SCE_c_297_n N_SCE_c_304_n N_SCE_c_298_n
+ N_SCE_c_299_n SCE SCE SCE SCE N_SCE_c_308_n N_SCE_c_309_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%SCE
x_PM_SKY130_FD_SC_LP__SDFSBP_2%D N_D_M1008_g N_D_M1016_g N_D_c_391_n N_D_c_392_n
+ D D D D N_D_c_388_n N_D_c_389_n PM_SKY130_FD_SC_LP__SDFSBP_2%D
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_27_467# N_A_27_467#_M1004_s N_A_27_467#_M1029_s
+ N_A_27_467#_M1027_g N_A_27_467#_c_442_n N_A_27_467#_c_443_n
+ N_A_27_467#_M1020_g N_A_27_467#_c_445_n N_A_27_467#_c_446_n
+ N_A_27_467#_c_447_n N_A_27_467#_c_448_n N_A_27_467#_c_449_n
+ N_A_27_467#_c_450_n PM_SKY130_FD_SC_LP__SDFSBP_2%A_27_467#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%SCD N_SCD_c_511_n N_SCD_M1021_g N_SCD_c_512_n
+ N_SCD_c_513_n N_SCD_M1012_g N_SCD_c_506_n N_SCD_c_507_n N_SCD_c_508_n
+ N_SCD_c_514_n SCD SCD N_SCD_c_510_n PM_SKY130_FD_SC_LP__SDFSBP_2%SCD
x_PM_SKY130_FD_SC_LP__SDFSBP_2%CLK N_CLK_c_562_n N_CLK_M1023_g N_CLK_M1025_g CLK
+ N_CLK_c_565_n PM_SKY130_FD_SC_LP__SDFSBP_2%CLK
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_920_73# N_A_920_73#_M1033_d N_A_920_73#_M1006_d
+ N_A_920_73#_c_617_n N_A_920_73#_M1001_g N_A_920_73#_M1019_g
+ N_A_920_73#_M1041_g N_A_920_73#_c_607_n N_A_920_73#_M1043_g
+ N_A_920_73#_c_608_n N_A_920_73#_c_609_n N_A_920_73#_c_610_n
+ N_A_920_73#_c_623_n N_A_920_73#_c_611_n N_A_920_73#_c_612_n
+ N_A_920_73#_c_613_n N_A_920_73#_c_614_n N_A_920_73#_c_615_n
+ N_A_920_73#_c_616_n PM_SKY130_FD_SC_LP__SDFSBP_2%A_920_73#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_1291_93# N_A_1291_93#_M1036_s
+ N_A_1291_93#_M1003_d N_A_1291_93#_c_762_n N_A_1291_93#_M1035_g
+ N_A_1291_93#_c_769_n N_A_1291_93#_M1034_g N_A_1291_93#_c_763_n
+ N_A_1291_93#_c_764_n N_A_1291_93#_c_771_n N_A_1291_93#_c_820_p
+ N_A_1291_93#_c_772_n N_A_1291_93#_c_765_n N_A_1291_93#_c_773_n
+ N_A_1291_93#_c_766_n N_A_1291_93#_c_767_n N_A_1291_93#_c_775_n
+ N_A_1291_93#_c_776_n N_A_1291_93#_c_812_p N_A_1291_93#_c_768_n
+ N_A_1291_93#_c_777_n N_A_1291_93#_c_804_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%A_1291_93#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_1163_119# N_A_1163_119#_M1039_d
+ N_A_1163_119#_M1001_d N_A_1163_119#_M1003_g N_A_1163_119#_c_914_n
+ N_A_1163_119#_M1036_g N_A_1163_119#_M1013_g N_A_1163_119#_c_915_n
+ N_A_1163_119#_M1017_g N_A_1163_119#_c_916_n N_A_1163_119#_c_926_n
+ N_A_1163_119#_c_917_n N_A_1163_119#_c_927_n N_A_1163_119#_c_918_n
+ N_A_1163_119#_c_919_n N_A_1163_119#_c_920_n N_A_1163_119#_c_930_n
+ N_A_1163_119#_c_921_n N_A_1163_119#_c_922_n N_A_1163_119#_c_923_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%A_1163_119#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%SET_B N_SET_B_M1030_g N_SET_B_M1024_g
+ N_SET_B_c_1043_n N_SET_B_M1045_g N_SET_B_M1000_g N_SET_B_c_1044_n
+ N_SET_B_c_1045_n N_SET_B_c_1052_n N_SET_B_c_1053_n N_SET_B_c_1046_n
+ N_SET_B_c_1054_n N_SET_B_c_1055_n N_SET_B_c_1056_n SET_B N_SET_B_c_1047_n
+ N_SET_B_c_1048_n N_SET_B_c_1059_n N_SET_B_c_1060_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%SET_B
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_629_47# N_A_629_47#_M1023_d N_A_629_47#_M1025_d
+ N_A_629_47#_M1033_g N_A_629_47#_M1006_g N_A_629_47#_c_1173_n
+ N_A_629_47#_c_1174_n N_A_629_47#_c_1185_n N_A_629_47#_c_1186_n
+ N_A_629_47#_M1039_g N_A_629_47#_c_1176_n N_A_629_47#_M1026_g
+ N_A_629_47#_c_1188_n N_A_629_47#_M1031_g N_A_629_47#_M1032_g
+ N_A_629_47#_c_1178_n N_A_629_47#_c_1190_n N_A_629_47#_c_1179_n
+ N_A_629_47#_c_1180_n N_A_629_47#_c_1181_n N_A_629_47#_c_1182_n
+ N_A_629_47#_c_1183_n PM_SKY130_FD_SC_LP__SDFSBP_2%A_629_47#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_1946_369# N_A_1946_369#_M1028_s
+ N_A_1946_369#_M1010_s N_A_1946_369#_M1002_g N_A_1946_369#_M1038_g
+ N_A_1946_369#_c_1303_n N_A_1946_369#_c_1304_n N_A_1946_369#_c_1305_n
+ N_A_1946_369#_c_1306_n N_A_1946_369#_c_1307_n N_A_1946_369#_c_1313_n
+ N_A_1946_369#_c_1308_n N_A_1946_369#_c_1309_n N_A_1946_369#_c_1310_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%A_1946_369#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_1799_408# N_A_1799_408#_M1041_d
+ N_A_1799_408#_M1031_d N_A_1799_408#_M1000_d N_A_1799_408#_M1028_g
+ N_A_1799_408#_M1010_g N_A_1799_408#_c_1395_n N_A_1799_408#_M1018_g
+ N_A_1799_408#_M1022_g N_A_1799_408#_M1037_g N_A_1799_408#_M1040_g
+ N_A_1799_408#_c_1400_n N_A_1799_408#_c_1401_n N_A_1799_408#_M1042_g
+ N_A_1799_408#_M1009_g N_A_1799_408#_c_1404_n N_A_1799_408#_c_1414_n
+ N_A_1799_408#_c_1405_n N_A_1799_408#_c_1406_n N_A_1799_408#_c_1416_n
+ N_A_1799_408#_c_1417_n N_A_1799_408#_c_1418_n N_A_1799_408#_c_1419_n
+ N_A_1799_408#_c_1456_n N_A_1799_408#_c_1420_n N_A_1799_408#_c_1407_n
+ N_A_1799_408#_c_1408_n N_A_1799_408#_c_1421_n N_A_1799_408#_c_1409_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%A_1799_408#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_2624_49# N_A_2624_49#_M1042_d
+ N_A_2624_49#_M1009_d N_A_2624_49#_M1007_g N_A_2624_49#_M1014_g
+ N_A_2624_49#_M1015_g N_A_2624_49#_M1044_g N_A_2624_49#_c_1573_n
+ N_A_2624_49#_c_1574_n N_A_2624_49#_c_1575_n N_A_2624_49#_c_1576_n
+ N_A_2624_49#_c_1577_n N_A_2624_49#_c_1578_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%A_2624_49#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%VPWR N_VPWR_M1029_d N_VPWR_M1021_d N_VPWR_M1006_s
+ N_VPWR_M1034_d N_VPWR_M1030_d N_VPWR_M1002_d N_VPWR_M1010_d N_VPWR_M1040_d
+ N_VPWR_M1014_s N_VPWR_M1044_s N_VPWR_c_1628_n N_VPWR_c_1629_n N_VPWR_c_1630_n
+ N_VPWR_c_1631_n N_VPWR_c_1632_n N_VPWR_c_1633_n N_VPWR_c_1634_n
+ N_VPWR_c_1635_n N_VPWR_c_1636_n N_VPWR_c_1637_n N_VPWR_c_1638_n
+ N_VPWR_c_1639_n N_VPWR_c_1640_n N_VPWR_c_1641_n N_VPWR_c_1642_n
+ N_VPWR_c_1643_n N_VPWR_c_1644_n N_VPWR_c_1645_n N_VPWR_c_1646_n
+ N_VPWR_c_1647_n VPWR N_VPWR_c_1648_n N_VPWR_c_1649_n N_VPWR_c_1650_n
+ N_VPWR_c_1651_n N_VPWR_c_1652_n N_VPWR_c_1653_n N_VPWR_c_1654_n
+ N_VPWR_c_1655_n N_VPWR_c_1656_n N_VPWR_c_1627_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%VPWR
x_PM_SKY130_FD_SC_LP__SDFSBP_2%A_268_467# N_A_268_467#_M1016_d
+ N_A_268_467#_M1039_s N_A_268_467#_M1008_d N_A_268_467#_M1001_s
+ N_A_268_467#_c_1806_n N_A_268_467#_c_1796_n N_A_268_467#_c_1797_n
+ N_A_268_467#_c_1798_n N_A_268_467#_c_1799_n N_A_268_467#_c_1800_n
+ N_A_268_467#_c_1801_n N_A_268_467#_c_1802_n N_A_268_467#_c_1808_n
+ N_A_268_467#_c_1809_n N_A_268_467#_c_1810_n N_A_268_467#_c_1811_n
+ N_A_268_467#_c_1803_n N_A_268_467#_c_1804_n N_A_268_467#_c_1805_n
+ N_A_268_467#_c_1813_n PM_SKY130_FD_SC_LP__SDFSBP_2%A_268_467#
x_PM_SKY130_FD_SC_LP__SDFSBP_2%Q_N N_Q_N_M1018_d N_Q_N_M1022_s Q_N Q_N Q_N Q_N
+ Q_N N_Q_N_c_1930_n N_Q_N_c_1935_n N_Q_N_c_1932_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%Q_N
x_PM_SKY130_FD_SC_LP__SDFSBP_2%Q N_Q_M1007_s N_Q_M1014_d Q Q Q Q Q Q Q
+ N_Q_c_1960_n PM_SKY130_FD_SC_LP__SDFSBP_2%Q
x_PM_SKY130_FD_SC_LP__SDFSBP_2%VGND N_VGND_M1004_d N_VGND_M1012_d N_VGND_M1033_s
+ N_VGND_M1035_d N_VGND_M1024_d N_VGND_M1045_d N_VGND_M1028_d N_VGND_M1037_s
+ N_VGND_M1007_d N_VGND_M1015_d N_VGND_c_1982_n N_VGND_c_1983_n N_VGND_c_1984_n
+ N_VGND_c_1985_n N_VGND_c_1986_n N_VGND_c_1987_n N_VGND_c_1988_n
+ N_VGND_c_1989_n N_VGND_c_1990_n N_VGND_c_1991_n N_VGND_c_1992_n
+ N_VGND_c_1993_n N_VGND_c_1994_n N_VGND_c_1995_n N_VGND_c_1996_n
+ N_VGND_c_1997_n N_VGND_c_1998_n N_VGND_c_1999_n N_VGND_c_2000_n
+ N_VGND_c_2001_n N_VGND_c_2002_n N_VGND_c_2003_n VGND N_VGND_c_2004_n
+ N_VGND_c_2005_n N_VGND_c_2006_n N_VGND_c_2007_n N_VGND_c_2008_n
+ N_VGND_c_2009_n N_VGND_c_2010_n N_VGND_c_2011_n N_VGND_c_2012_n
+ PM_SKY130_FD_SC_LP__SDFSBP_2%VGND
cc_1 VNB N_SCE_c_294_n 0.00200128f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.845
cc_2 VNB N_SCE_M1004_g 0.0599247f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_3 VNB N_SCE_M1011_g 0.0374923f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.445
cc_4 VNB N_SCE_c_297_n 0.0242476f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.53
cc_5 VNB N_SCE_c_298_n 0.00131314f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.33
cc_6 VNB N_SCE_c_299_n 0.039977f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.33
cc_7 VNB SCE 0.0098913f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB D 0.010536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D_c_388_n 0.03185f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.33
cc_10 VNB N_D_c_389_n 0.016341f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.33
cc_11 VNB N_A_27_467#_M1027_g 0.0196595f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_12 VNB N_A_27_467#_c_442_n 0.034101f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.175
cc_13 VNB N_A_27_467#_c_443_n 0.0164235f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.655
cc_14 VNB N_A_27_467#_M1020_g 0.0102743f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.165
cc_15 VNB N_A_27_467#_c_445_n 0.0261111f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.53
cc_16 VNB N_A_27_467#_c_446_n 0.035751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_467#_c_447_n 0.00728713f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.165
cc_18 VNB N_A_27_467#_c_448_n 0.0439039f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.33
cc_19 VNB N_A_27_467#_c_449_n 0.0122561f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_20 VNB N_A_27_467#_c_450_n 0.0141769f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_21 VNB N_SCD_c_506_n 0.0158306f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.175
cc_22 VNB N_SCD_c_507_n 0.0110479f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.655
cc_23 VNB N_SCD_c_508_n 0.0319482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB SCD 0.00310715f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.445
cc_25 VNB N_SCD_c_510_n 0.00973642f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.53
cc_26 VNB N_CLK_c_562_n 0.0198078f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.605
cc_27 VNB N_CLK_M1025_g 0.0350669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB CLK 0.00510864f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_29 VNB N_CLK_c_565_n 0.0365676f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.165
cc_30 VNB N_A_920_73#_M1019_g 0.0375273f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.165
cc_31 VNB N_A_920_73#_M1041_g 0.0178303f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.53
cc_32 VNB N_A_920_73#_c_607_n 0.0139546f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.53
cc_33 VNB N_A_920_73#_c_608_n 0.0254417f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.33
cc_34 VNB N_A_920_73#_c_609_n 0.0102311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_920_73#_c_610_n 0.00203491f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_36 VNB N_A_920_73#_c_611_n 0.00100362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_920_73#_c_612_n 0.0249805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_920_73#_c_613_n 0.00713979f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_39 VNB N_A_920_73#_c_614_n 0.0318021f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_40 VNB N_A_920_73#_c_615_n 0.00247483f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_41 VNB N_A_920_73#_c_616_n 0.0157461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1291_93#_c_762_n 0.0189083f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.455
cc_43 VNB N_A_1291_93#_c_763_n 0.0204908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1291_93#_c_764_n 0.0208244f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.445
cc_45 VNB N_A_1291_93#_c_765_n 0.0013688f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_46 VNB N_A_1291_93#_c_766_n 0.00259013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1291_93#_c_767_n 0.00567093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1291_93#_c_768_n 8.64496e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_49 VNB N_A_1163_119#_M1003_g 0.0116946f $X=-0.19 $Y=-0.245 $X2=0.725
+ $Y2=0.445
cc_50 VNB N_A_1163_119#_c_914_n 0.0192996f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=2.175
cc_51 VNB N_A_1163_119#_c_915_n 0.0165597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1163_119#_c_916_n 0.00112185f $X=-0.19 $Y=-0.245 $X2=2.255
+ $Y2=1.33
cc_53 VNB N_A_1163_119#_c_917_n 0.00894766f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_54 VNB N_A_1163_119#_c_918_n 0.0297801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1163_119#_c_919_n 0.00406213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1163_119#_c_920_n 0.00494961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1163_119#_c_921_n 0.0432415f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_58 VNB N_A_1163_119#_c_922_n 0.0240389f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_59 VNB N_A_1163_119#_c_923_n 3.8708e-19 $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.01
cc_60 VNB N_SET_B_M1024_g 0.0453898f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.455
cc_61 VNB N_SET_B_c_1043_n 0.0200737f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_62 VNB N_SET_B_c_1044_n 0.0348391f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.445
cc_63 VNB N_SET_B_c_1045_n 0.00649978f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.445
cc_64 VNB N_SET_B_c_1046_n 0.021458f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.33
cc_65 VNB N_SET_B_c_1047_n 0.00709537f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_66 VNB N_SET_B_c_1048_n 0.00141224f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_67 VNB N_A_629_47#_M1033_g 0.0132445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_629_47#_M1006_g 0.00728621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_629_47#_c_1173_n 0.0846783f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.165
cc_70 VNB N_A_629_47#_c_1174_n 0.0125025f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.445
cc_71 VNB N_A_629_47#_M1039_g 0.045345f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.53
cc_72 VNB N_A_629_47#_c_1176_n 0.290561f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.33
cc_73 VNB N_A_629_47#_M1032_g 0.0413639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_629_47#_c_1178_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_629_47#_c_1179_n 0.0149126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_629_47#_c_1180_n 0.00420747f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.01
cc_77 VNB N_A_629_47#_c_1181_n 0.00972793f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_78 VNB N_A_629_47#_c_1182_n 0.0614268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_629_47#_c_1183_n 0.0955028f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_80 VNB N_A_1946_369#_M1038_g 0.0400515f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=2.655
cc_81 VNB N_A_1946_369#_c_1303_n 0.00666474f $X=-0.19 $Y=-0.245 $X2=2.28
+ $Y2=0.445
cc_82 VNB N_A_1946_369#_c_1304_n 0.0248955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1946_369#_c_1305_n 0.00928997f $X=-0.19 $Y=-0.245 $X2=0.725
+ $Y2=1.53
cc_84 VNB N_A_1946_369#_c_1306_n 0.0100653f $X=-0.19 $Y=-0.245 $X2=2.255
+ $Y2=1.165
cc_85 VNB N_A_1946_369#_c_1307_n 0.00695336f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=2.33
cc_86 VNB N_A_1946_369#_c_1308_n 0.00252727f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_87 VNB N_A_1946_369#_c_1309_n 0.0026983f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_88 VNB N_A_1946_369#_c_1310_n 0.0211329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1799_408#_M1028_g 0.0313721f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=2.655
cc_90 VNB N_A_1799_408#_c_1395_n 0.0135294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1799_408#_M1018_g 0.026728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1799_408#_M1022_g 0.00731487f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=2.33
cc_93 VNB N_A_1799_408#_M1037_g 0.0241414f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.33
cc_94 VNB N_A_1799_408#_M1040_g 0.00861806f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_95 VNB N_A_1799_408#_c_1400_n 0.0107227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1799_408#_c_1401_n 0.0222774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1799_408#_M1042_g 0.0540006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1799_408#_M1009_g 0.00935016f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_99 VNB N_A_1799_408#_c_1404_n 0.0174907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1799_408#_c_1405_n 0.00569716f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=2.367
cc_101 VNB N_A_1799_408#_c_1406_n 0.012175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1799_408#_c_1407_n 0.00412153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1799_408#_c_1408_n 4.02031e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1799_408#_c_1409_n 0.0344947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2624_49#_M1007_g 0.0290117f $X=-0.19 $Y=-0.245 $X2=0.725
+ $Y2=0.445
cc_106 VNB N_A_2624_49#_M1014_g 0.00392759f $X=-0.19 $Y=-0.245 $X2=0.905
+ $Y2=2.655
cc_107 VNB N_A_2624_49#_M1015_g 0.0312807f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.445
cc_108 VNB N_A_2624_49#_M1044_g 0.00373837f $X=-0.19 $Y=-0.245 $X2=0.725
+ $Y2=1.53
cc_109 VNB N_A_2624_49#_c_1573_n 0.0149126f $X=-0.19 $Y=-0.245 $X2=2.255
+ $Y2=1.165
cc_110 VNB N_A_2624_49#_c_1574_n 0.00196628f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.245
cc_111 VNB N_A_2624_49#_c_1575_n 0.00871972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2624_49#_c_1576_n 0.00443288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2624_49#_c_1577_n 0.00589363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2624_49#_c_1578_n 0.112317f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_115 VNB N_VPWR_c_1627_n 0.641339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_268_467#_c_1796_n 3.9527e-19 $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=1.53
cc_117 VNB N_A_268_467#_c_1797_n 0.00688344f $X=-0.19 $Y=-0.245 $X2=0.725
+ $Y2=1.53
cc_118 VNB N_A_268_467#_c_1798_n 0.00703243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_268_467#_c_1799_n 0.00293709f $X=-0.19 $Y=-0.245 $X2=2.255
+ $Y2=1.165
cc_120 VNB N_A_268_467#_c_1800_n 0.00998033f $X=-0.19 $Y=-0.245 $X2=2.09
+ $Y2=2.33
cc_121 VNB N_A_268_467#_c_1801_n 0.00206549f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=2.33
cc_122 VNB N_A_268_467#_c_1802_n 0.00249515f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=1.33
cc_123 VNB N_A_268_467#_c_1803_n 0.00834486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_268_467#_c_1804_n 0.00961345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_268_467#_c_1805_n 0.00852984f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=2.01
cc_126 VNB N_Q_N_c_1930_n 0.00280345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB Q 0.00270177f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_128 VNB N_Q_c_1960_n 0.00422824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1982_n 0.00557476f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_130 VNB N_VGND_c_1983_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1984_n 0.0141145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1985_n 0.0236139f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.01
cc_133 VNB N_VGND_c_1986_n 0.0192507f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.245
cc_134 VNB N_VGND_c_1987_n 0.0324314f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_135 VNB N_VGND_c_1988_n 0.0177141f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.367
cc_136 VNB N_VGND_c_1989_n 0.0183986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1990_n 0.018857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1991_n 0.0156606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1992_n 0.0120163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1993_n 0.0487156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1994_n 0.023462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1995_n 0.00632207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1996_n 0.0414647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1997_n 0.00436557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1998_n 0.0279103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1999_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2000_n 0.0632418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2001_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2002_n 0.0549943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2003_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2004_n 0.0338825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2005_n 0.0269506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2006_n 0.0176662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2007_n 0.0255466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2008_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2009_n 0.00836712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2010_n 0.00644364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2011_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2012_n 0.757157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VPB N_SCE_c_294_n 0.00876651f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.845
cc_161 VPB N_SCE_M1029_g 0.0229304f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.655
cc_162 VPB N_SCE_M1005_g 0.0173795f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.655
cc_163 VPB N_SCE_c_304_n 0.017226f $X=-0.19 $Y=1.655 $X2=2.09 $Y2=2.33
cc_164 VPB N_SCE_c_298_n 0.00506236f $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.33
cc_165 VPB N_SCE_c_299_n 0.019163f $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.33
cc_166 VPB SCE 0.00573277f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_167 VPB N_SCE_c_308_n 0.0474039f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.01
cc_168 VPB N_SCE_c_309_n 0.00134721f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.367
cc_169 VPB N_D_M1008_g 0.0214103f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.175
cc_170 VPB N_D_c_391_n 0.00405932f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.445
cc_171 VPB N_D_c_392_n 0.030947f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.175
cc_172 VPB D 0.00261969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_27_467#_M1020_g 0.0493687f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=1.165
cc_174 VPB N_A_27_467#_c_446_n 0.0620385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_SCD_c_511_n 0.0196221f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.605
cc_176 VPB N_SCD_c_512_n 0.0358959f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.655
cc_177 VPB N_SCD_c_513_n 0.006911f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.655
cc_178 VPB N_SCD_c_514_n 0.0251124f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=1.165
cc_179 VPB SCD 0.00784991f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=0.445
cc_180 VPB N_SCD_c_510_n 0.00568302f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.53
cc_181 VPB N_CLK_M1025_g 0.051406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_920_73#_c_617_n 0.023067f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.455
cc_183 VPB N_A_920_73#_M1001_g 0.0413716f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.175
cc_184 VPB N_A_920_73#_c_607_n 0.00674565f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.53
cc_185 VPB N_A_920_73#_M1043_g 0.0510453f $X=-0.19 $Y=1.655 $X2=2.09 $Y2=2.33
cc_186 VPB N_A_920_73#_c_609_n 0.0143417f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_920_73#_c_610_n 0.00554911f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_188 VPB N_A_920_73#_c_623_n 0.00980108f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_189 VPB N_A_920_73#_c_611_n 0.00254336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_920_73#_c_612_n 0.0100932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_920_73#_c_613_n 0.00483639f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.01
cc_192 VPB N_A_920_73#_c_614_n 0.0441499f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.01
cc_193 VPB N_A_920_73#_c_615_n 0.00437715f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.295
cc_194 VPB N_A_920_73#_c_616_n 0.0322545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1291_93#_c_769_n 0.059405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1291_93#_c_763_n 0.00855423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_1291_93#_c_771_n 0.00100759f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.53
cc_198 VPB N_A_1291_93#_c_772_n 0.00200767f $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.33
cc_199 VPB N_A_1291_93#_c_773_n 0.0012428f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_200 VPB N_A_1291_93#_c_767_n 0.00458843f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1291_93#_c_775_n 0.00324838f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.01
cc_202 VPB N_A_1291_93#_c_776_n 0.00191573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1291_93#_c_777_n 0.00149069f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.01
cc_204 VPB N_A_1163_119#_M1003_g 0.0438186f $X=-0.19 $Y=1.655 $X2=0.725
+ $Y2=0.445
cc_205 VPB N_A_1163_119#_M1013_g 0.0244519f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=0.445
cc_206 VPB N_A_1163_119#_c_926_n 8.5954e-19 $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.33
cc_207 VPB N_A_1163_119#_c_927_n 7.2632e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1163_119#_c_918_n 0.00635824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_1163_119#_c_920_n 0.0022095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1163_119#_c_930_n 0.00373541f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=2.01
cc_211 VPB N_SET_B_M1030_g 0.0204698f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.175
cc_212 VPB N_SET_B_M1024_g 0.00994982f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.455
cc_213 VPB N_SET_B_M1000_g 0.0260934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_SET_B_c_1052_n 0.0310281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_SET_B_c_1053_n 0.0105484f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.53
cc_216 VPB N_SET_B_c_1054_n 0.0305143f $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.165
cc_217 VPB N_SET_B_c_1055_n 0.0292415f $X=-0.19 $Y=1.655 $X2=2.09 $Y2=2.33
cc_218 VPB N_SET_B_c_1056_n 0.00148081f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.33
cc_219 VPB N_SET_B_c_1047_n 0.0116372f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_220 VPB N_SET_B_c_1048_n 0.00188574f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_221 VPB N_SET_B_c_1059_n 0.00220422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_SET_B_c_1060_n 0.0430219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_629_47#_M1006_g 0.0618206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_629_47#_c_1185_n 0.119996f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=0.445
cc_225 VPB N_A_629_47#_c_1186_n 0.0125055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_629_47#_M1026_g 0.0344598f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.245
cc_227 VPB N_A_629_47#_c_1188_n 0.198179f $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.33
cc_228 VPB N_A_629_47#_M1031_g 0.0232926f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_229 VPB N_A_629_47#_c_1190_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_629_47#_c_1180_n 0.032141f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.01
cc_231 VPB N_A_1946_369#_M1002_g 0.0357328f $X=-0.19 $Y=1.655 $X2=0.725
+ $Y2=0.445
cc_232 VPB N_A_1946_369#_c_1303_n 0.00292636f $X=-0.19 $Y=1.655 $X2=2.28
+ $Y2=0.445
cc_233 VPB N_A_1946_369#_c_1313_n 0.00177205f $X=-0.19 $Y=1.655 $X2=2.215
+ $Y2=1.33
cc_234 VPB N_A_1946_369#_c_1308_n 0.0010891f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.58
cc_235 VPB N_A_1946_369#_c_1310_n 0.0457351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_1799_408#_M1010_g 0.0264706f $X=-0.19 $Y=1.655 $X2=2.28 $Y2=0.445
cc_237 VPB N_A_1799_408#_M1022_g 0.0215146f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.33
cc_238 VPB N_A_1799_408#_M1040_g 0.0230546f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_239 VPB N_A_1799_408#_M1009_g 0.0276976f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.01
cc_240 VPB N_A_1799_408#_c_1414_n 0.00579189f $X=-0.19 $Y=1.655 $X2=0.72
+ $Y2=1.665
cc_241 VPB N_A_1799_408#_c_1406_n 0.00385034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1799_408#_c_1416_n 0.00103228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1799_408#_c_1417_n 0.0136317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1799_408#_c_1418_n 0.00162215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_1799_408#_c_1419_n 0.0214036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1799_408#_c_1420_n 0.0181934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_1799_408#_c_1421_n 0.00110508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_1799_408#_c_1409_n 0.0163349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_2624_49#_M1014_g 0.0265631f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.655
cc_250 VPB N_A_2624_49#_M1044_g 0.0266392f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.53
cc_251 VPB N_A_2624_49#_c_1574_n 0.0233443f $X=-0.19 $Y=1.655 $X2=2.215
+ $Y2=2.245
cc_252 VPB N_VPWR_c_1628_n 0.0035785f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_253 VPB N_VPWR_c_1629_n 0.0144464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1630_n 0.0141605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1631_n 0.0146598f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.01
cc_256 VPB N_VPWR_c_1632_n 0.00976411f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.245
cc_257 VPB N_VPWR_c_1633_n 0.0233031f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_258 VPB N_VPWR_c_1634_n 0.0350539f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.367
cc_259 VPB N_VPWR_c_1635_n 0.0382456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1636_n 0.0119904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1637_n 0.0637164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1638_n 0.0335573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1639_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1640_n 0.0228034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1641_n 0.00435574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1642_n 0.0481716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1643_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1644_n 0.0478018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1645_n 0.00497181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1646_n 0.0172627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1647_n 0.00651392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1648_n 0.0165577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1649_n 0.0446726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1650_n 0.0735102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1651_n 0.0295308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1652_n 0.0152106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1653_n 0.00583335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1654_n 0.0137656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1655_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1656_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1627_n 0.16228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_A_268_467#_c_1806_n 0.00138873f $X=-0.19 $Y=1.655 $X2=0.905
+ $Y2=2.655
cc_283 VPB N_A_268_467#_c_1802_n 0.00478689f $X=-0.19 $Y=1.655 $X2=2.215
+ $Y2=1.33
cc_284 VPB N_A_268_467#_c_1808_n 0.0123576f $X=-0.19 $Y=1.655 $X2=2.255 $Y2=1.33
cc_285 VPB N_A_268_467#_c_1809_n 0.00741151f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.21
cc_286 VPB N_A_268_467#_c_1810_n 0.0214484f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_287 VPB N_A_268_467#_c_1811_n 0.0091522f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_288 VPB N_A_268_467#_c_1804_n 0.0131271f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_A_268_467#_c_1813_n 0.00862067f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.01
cc_290 VPB N_Q_N_c_1930_n 0.00278593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_Q_N_c_1932_n 0.0041135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB Q 0.00173401f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.445
cc_293 N_SCE_M1005_g N_D_M1008_g 0.0398232f $X=0.905 $Y=2.655 $X2=0 $Y2=0
cc_294 N_SCE_c_304_n N_D_M1008_g 0.0150921f $X=2.09 $Y=2.33 $X2=0 $Y2=0
cc_295 N_SCE_c_304_n N_D_c_391_n 0.0468159f $X=2.09 $Y=2.33 $X2=0 $Y2=0
cc_296 N_SCE_c_298_n N_D_c_391_n 0.0141079f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_297 SCE N_D_c_391_n 0.0128874f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_298 N_SCE_c_308_n N_D_c_391_n 9.43609e-19 $X=0.905 $Y=2.01 $X2=0 $Y2=0
cc_299 N_SCE_c_304_n N_D_c_392_n 0.00438369f $X=2.09 $Y=2.33 $X2=0 $Y2=0
cc_300 SCE N_D_c_392_n 0.00138145f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_301 N_SCE_c_308_n N_D_c_392_n 0.0398232f $X=0.905 $Y=2.01 $X2=0 $Y2=0
cc_302 N_SCE_M1011_g D 0.00390812f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_303 N_SCE_c_298_n D 0.0314453f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_304 N_SCE_c_299_n D 0.0050324f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_305 SCE D 0.0108966f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_306 N_SCE_M1011_g N_D_c_388_n 0.0120185f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_307 N_SCE_M1011_g N_D_c_389_n 0.00964823f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_308 N_SCE_M1004_g N_A_27_467#_M1027_g 0.0106876f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_309 N_SCE_c_298_n N_A_27_467#_c_442_n 0.00176846f $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_310 N_SCE_c_299_n N_A_27_467#_c_442_n 0.0302653f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_311 N_SCE_c_304_n N_A_27_467#_M1020_g 0.0138207f $X=2.09 $Y=2.33 $X2=0 $Y2=0
cc_312 N_SCE_c_298_n N_A_27_467#_M1020_g 0.0084694f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_313 N_SCE_c_297_n N_A_27_467#_c_445_n 0.0212475f $X=0.725 $Y=1.53 $X2=0 $Y2=0
cc_314 SCE N_A_27_467#_c_445_n 0.00213052f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_315 N_SCE_M1004_g N_A_27_467#_c_446_n 0.00705019f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_316 N_SCE_c_297_n N_A_27_467#_c_446_n 0.0249343f $X=0.725 $Y=1.53 $X2=0 $Y2=0
cc_317 SCE N_A_27_467#_c_446_n 0.0774898f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_318 N_SCE_c_309_n N_A_27_467#_c_446_n 0.00681727f $X=0.985 $Y=2.367 $X2=0
+ $Y2=0
cc_319 N_SCE_M1004_g N_A_27_467#_c_447_n 0.00945748f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_320 SCE N_A_27_467#_c_447_n 0.0177592f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_321 N_SCE_M1004_g N_A_27_467#_c_448_n 0.0161485f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_322 N_SCE_c_297_n N_A_27_467#_c_448_n 0.0058583f $X=0.725 $Y=1.53 $X2=0 $Y2=0
cc_323 SCE N_A_27_467#_c_448_n 0.00960052f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_324 N_SCE_M1004_g N_A_27_467#_c_449_n 0.00133947f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_325 SCE N_A_27_467#_c_449_n 0.0258349f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_326 N_SCE_M1004_g N_A_27_467#_c_450_n 0.0212475f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_327 N_SCE_c_304_n N_SCD_c_511_n 0.0126988f $X=2.09 $Y=2.33 $X2=-0.19
+ $Y2=-0.245
cc_328 N_SCE_c_298_n N_SCD_c_511_n 4.4694e-19 $X=2.255 $Y=1.33 $X2=-0.19
+ $Y2=-0.245
cc_329 N_SCE_c_298_n N_SCD_c_513_n 0.00588711f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_330 N_SCE_c_299_n N_SCD_c_513_n 0.0111972f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_331 N_SCE_M1011_g N_SCD_c_506_n 0.050605f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_332 N_SCE_M1011_g N_SCD_c_508_n 0.00992485f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_333 N_SCE_c_298_n N_SCD_c_508_n 0.0013866f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_334 N_SCE_c_299_n N_SCD_c_508_n 0.0207245f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_335 N_SCE_c_298_n N_SCD_c_514_n 0.0012864f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_336 N_SCE_c_304_n SCD 4.24054e-19 $X=2.09 $Y=2.33 $X2=0 $Y2=0
cc_337 N_SCE_c_298_n SCD 0.0559694f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_338 N_SCE_c_299_n SCD 0.00201777f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_339 N_SCE_c_299_n N_SCD_c_510_n 0.0207245f $X=2.255 $Y=1.33 $X2=0 $Y2=0
cc_340 N_SCE_c_309_n N_VPWR_M1029_d 0.00205792f $X=0.985 $Y=2.367 $X2=-0.19
+ $Y2=-0.245
cc_341 N_SCE_M1029_g N_VPWR_c_1628_n 0.011459f $X=0.475 $Y=2.655 $X2=0 $Y2=0
cc_342 N_SCE_M1005_g N_VPWR_c_1628_n 0.0102067f $X=0.905 $Y=2.655 $X2=0 $Y2=0
cc_343 N_SCE_c_309_n N_VPWR_c_1628_n 0.0153247f $X=0.985 $Y=2.367 $X2=0 $Y2=0
cc_344 N_SCE_M1029_g N_VPWR_c_1648_n 0.00393414f $X=0.475 $Y=2.655 $X2=0 $Y2=0
cc_345 N_SCE_M1005_g N_VPWR_c_1649_n 0.00393414f $X=0.905 $Y=2.655 $X2=0 $Y2=0
cc_346 N_SCE_M1029_g N_VPWR_c_1627_n 0.00782316f $X=0.475 $Y=2.655 $X2=0 $Y2=0
cc_347 N_SCE_M1005_g N_VPWR_c_1627_n 0.00391996f $X=0.905 $Y=2.655 $X2=0 $Y2=0
cc_348 N_SCE_c_309_n N_VPWR_c_1627_n 0.00473938f $X=0.985 $Y=2.367 $X2=0 $Y2=0
cc_349 N_SCE_c_304_n A_196_467# 0.00366293f $X=2.09 $Y=2.33 $X2=-0.19 $Y2=-0.245
cc_350 N_SCE_c_304_n N_A_268_467#_M1008_d 0.00384225f $X=2.09 $Y=2.33 $X2=0
+ $Y2=0
cc_351 N_SCE_c_304_n N_A_268_467#_c_1806_n 0.0554139f $X=2.09 $Y=2.33 $X2=0
+ $Y2=0
cc_352 N_SCE_M1011_g N_A_268_467#_c_1796_n 0.00763355f $X=2.28 $Y=0.445 $X2=0
+ $Y2=0
cc_353 N_SCE_M1011_g N_A_268_467#_c_1797_n 0.00980763f $X=2.28 $Y=0.445 $X2=0
+ $Y2=0
cc_354 N_SCE_c_298_n N_A_268_467#_c_1797_n 0.0058811f $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_355 N_SCE_c_299_n N_A_268_467#_c_1797_n 0.00235049f $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_356 N_SCE_M1011_g N_A_268_467#_c_1798_n 0.00244801f $X=2.28 $Y=0.445 $X2=0
+ $Y2=0
cc_357 N_SCE_c_298_n N_A_268_467#_c_1798_n 0.00755136f $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_358 N_SCE_c_299_n N_A_268_467#_c_1798_n 8.19163e-19 $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_359 N_SCE_M1011_g N_A_268_467#_c_1799_n 0.00596137f $X=2.28 $Y=0.445 $X2=0
+ $Y2=0
cc_360 N_SCE_c_298_n N_A_268_467#_c_1799_n 0.00207847f $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_361 N_SCE_c_298_n N_A_268_467#_c_1801_n 0.013491f $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_362 N_SCE_c_299_n N_A_268_467#_c_1801_n 0.00122794f $X=2.255 $Y=1.33 $X2=0
+ $Y2=0
cc_363 N_SCE_c_304_n A_376_467# 0.00265142f $X=2.09 $Y=2.33 $X2=-0.19 $Y2=-0.245
cc_364 N_SCE_M1004_g N_VGND_c_1982_n 0.00327093f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_365 N_SCE_M1011_g N_VGND_c_1983_n 0.00205524f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_366 N_SCE_M1004_g N_VGND_c_1994_n 0.00571971f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_367 N_SCE_M1011_g N_VGND_c_1996_n 0.00429366f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_368 N_SCE_M1004_g N_VGND_c_2012_n 0.00764979f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_369 N_SCE_M1011_g N_VGND_c_2012_n 0.00645269f $X=2.28 $Y=0.445 $X2=0 $Y2=0
cc_370 D N_A_27_467#_M1027_g 0.00418128f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_371 N_D_c_389_n N_A_27_467#_M1027_g 0.0307721f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_372 N_D_c_391_n N_A_27_467#_c_442_n 0.00103215f $X=1.515 $Y=1.945 $X2=0 $Y2=0
cc_373 D N_A_27_467#_c_442_n 0.0156817f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_374 N_D_c_388_n N_A_27_467#_c_442_n 0.0193412f $X=1.715 $Y=0.93 $X2=0 $Y2=0
cc_375 N_D_c_392_n N_A_27_467#_c_443_n 0.0129101f $X=1.355 $Y=1.98 $X2=0 $Y2=0
cc_376 N_D_M1008_g N_A_27_467#_M1020_g 0.0254527f $X=1.265 $Y=2.655 $X2=0 $Y2=0
cc_377 N_D_c_391_n N_A_27_467#_M1020_g 0.00769087f $X=1.515 $Y=1.945 $X2=0 $Y2=0
cc_378 N_D_c_392_n N_A_27_467#_M1020_g 0.0215105f $X=1.355 $Y=1.98 $X2=0 $Y2=0
cc_379 D N_A_27_467#_M1020_g 0.0112828f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_380 N_D_c_391_n N_A_27_467#_c_449_n 0.00705441f $X=1.515 $Y=1.945 $X2=0 $Y2=0
cc_381 N_D_c_392_n N_A_27_467#_c_449_n 7.25738e-19 $X=1.355 $Y=1.98 $X2=0 $Y2=0
cc_382 D N_A_27_467#_c_449_n 0.0544013f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_383 N_D_c_388_n N_A_27_467#_c_449_n 9.10603e-19 $X=1.715 $Y=0.93 $X2=0 $Y2=0
cc_384 D N_A_27_467#_c_450_n 0.00261839f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_385 N_D_c_388_n N_A_27_467#_c_450_n 0.0307721f $X=1.715 $Y=0.93 $X2=0 $Y2=0
cc_386 N_D_M1008_g N_VPWR_c_1628_n 0.00199365f $X=1.265 $Y=2.655 $X2=0 $Y2=0
cc_387 N_D_M1008_g N_VPWR_c_1649_n 0.00473823f $X=1.265 $Y=2.655 $X2=0 $Y2=0
cc_388 N_D_M1008_g N_VPWR_c_1627_n 0.00938177f $X=1.265 $Y=2.655 $X2=0 $Y2=0
cc_389 D N_A_268_467#_M1016_d 0.00304546f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_390 N_D_M1008_g N_A_268_467#_c_1806_n 0.00459578f $X=1.265 $Y=2.655 $X2=0
+ $Y2=0
cc_391 D N_A_268_467#_c_1796_n 0.0249741f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_392 N_D_c_389_n N_A_268_467#_c_1796_n 0.00326261f $X=1.715 $Y=0.765 $X2=0
+ $Y2=0
cc_393 D N_A_268_467#_c_1798_n 0.0145039f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_394 N_D_c_388_n N_A_268_467#_c_1798_n 9.83449e-19 $X=1.715 $Y=0.93 $X2=0
+ $Y2=0
cc_395 N_D_c_389_n N_A_268_467#_c_1798_n 2.17334e-19 $X=1.715 $Y=0.765 $X2=0
+ $Y2=0
cc_396 D N_VGND_c_1996_n 0.0088773f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_397 N_D_c_388_n N_VGND_c_1996_n 0.00166803f $X=1.715 $Y=0.93 $X2=0 $Y2=0
cc_398 N_D_c_389_n N_VGND_c_1996_n 0.00383378f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_399 D N_VGND_c_2012_n 0.00949469f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_400 N_D_c_388_n N_VGND_c_2012_n 0.00191911f $X=1.715 $Y=0.93 $X2=0 $Y2=0
cc_401 N_D_c_389_n N_VGND_c_2012_n 0.00586206f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_402 N_A_27_467#_M1020_g N_SCD_c_513_n 0.0360076f $X=1.805 $Y=2.655 $X2=0
+ $Y2=0
cc_403 N_A_27_467#_c_446_n N_VPWR_c_1628_n 0.0125559f $X=0.26 $Y=2.48 $X2=0
+ $Y2=0
cc_404 N_A_27_467#_c_446_n N_VPWR_c_1648_n 0.0117477f $X=0.26 $Y=2.48 $X2=0
+ $Y2=0
cc_405 N_A_27_467#_M1020_g N_VPWR_c_1649_n 0.00322996f $X=1.805 $Y=2.655 $X2=0
+ $Y2=0
cc_406 N_A_27_467#_M1020_g N_VPWR_c_1627_n 0.0042288f $X=1.805 $Y=2.655 $X2=0
+ $Y2=0
cc_407 N_A_27_467#_c_446_n N_VPWR_c_1627_n 0.00955733f $X=0.26 $Y=2.48 $X2=0
+ $Y2=0
cc_408 N_A_27_467#_M1020_g N_A_268_467#_c_1806_n 0.0108572f $X=1.805 $Y=2.655
+ $X2=0 $Y2=0
cc_409 N_A_27_467#_M1027_g N_VGND_c_1982_n 0.00327093f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_27_467#_c_447_n N_VGND_c_1982_n 0.0140415f $X=1.055 $Y=0.9 $X2=0
+ $Y2=0
cc_411 N_A_27_467#_c_449_n N_VGND_c_1982_n 0.00636687f $X=1.175 $Y=0.98 $X2=0
+ $Y2=0
cc_412 N_A_27_467#_c_450_n N_VGND_c_1982_n 0.00188101f $X=1.175 $Y=0.98 $X2=0
+ $Y2=0
cc_413 N_A_27_467#_c_448_n N_VGND_c_1994_n 0.0337169f $X=0.51 $Y=0.44 $X2=0
+ $Y2=0
cc_414 N_A_27_467#_M1027_g N_VGND_c_1996_n 0.00585385f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_A_27_467#_M1004_s N_VGND_c_2012_n 0.00215817f $X=0.385 $Y=0.235 $X2=0
+ $Y2=0
cc_416 N_A_27_467#_M1027_g N_VGND_c_2012_n 0.00638409f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_417 N_A_27_467#_c_447_n N_VGND_c_2012_n 0.00575544f $X=1.055 $Y=0.9 $X2=0
+ $Y2=0
cc_418 N_A_27_467#_c_448_n N_VGND_c_2012_n 0.0215772f $X=0.51 $Y=0.44 $X2=0
+ $Y2=0
cc_419 N_A_27_467#_c_449_n N_VGND_c_2012_n 0.00651975f $X=1.175 $Y=0.98 $X2=0
+ $Y2=0
cc_420 N_SCD_c_506_n N_CLK_c_562_n 0.0140399f $X=2.672 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_421 N_SCD_c_508_n N_CLK_M1025_g 0.0122608f $X=2.795 $Y=1.58 $X2=0 $Y2=0
cc_422 SCD N_CLK_M1025_g 8.31211e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_423 N_SCD_c_510_n N_CLK_M1025_g 0.0330165f $X=2.795 $Y=1.745 $X2=0 $Y2=0
cc_424 N_SCD_c_507_n CLK 8.41963e-19 $X=2.672 $Y=0.925 $X2=0 $Y2=0
cc_425 N_SCD_c_507_n N_CLK_c_565_n 0.0190894f $X=2.672 $Y=0.925 $X2=0 $Y2=0
cc_426 N_SCD_c_511_n N_VPWR_c_1649_n 0.00322996f $X=2.315 $Y=2.225 $X2=0 $Y2=0
cc_427 N_SCD_c_511_n N_VPWR_c_1654_n 0.00531821f $X=2.315 $Y=2.225 $X2=0 $Y2=0
cc_428 N_SCD_c_511_n N_VPWR_c_1627_n 0.00434817f $X=2.315 $Y=2.225 $X2=0 $Y2=0
cc_429 N_SCD_c_511_n N_A_268_467#_c_1806_n 0.0214354f $X=2.315 $Y=2.225 $X2=0
+ $Y2=0
cc_430 N_SCD_c_512_n N_A_268_467#_c_1806_n 0.00730387f $X=2.63 $Y=2.15 $X2=0
+ $Y2=0
cc_431 SCD N_A_268_467#_c_1806_n 0.0197739f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_432 N_SCD_c_506_n N_A_268_467#_c_1796_n 0.0015207f $X=2.672 $Y=0.775 $X2=0
+ $Y2=0
cc_433 N_SCD_c_506_n N_A_268_467#_c_1797_n 0.00560374f $X=2.672 $Y=0.775 $X2=0
+ $Y2=0
cc_434 N_SCD_c_507_n N_A_268_467#_c_1797_n 0.00304675f $X=2.672 $Y=0.925 $X2=0
+ $Y2=0
cc_435 SCD N_A_268_467#_c_1797_n 2.80624e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_436 N_SCD_c_507_n N_A_268_467#_c_1799_n 0.00260884f $X=2.672 $Y=0.925 $X2=0
+ $Y2=0
cc_437 N_SCD_c_508_n N_A_268_467#_c_1799_n 0.00663903f $X=2.795 $Y=1.58 $X2=0
+ $Y2=0
cc_438 N_SCD_c_508_n N_A_268_467#_c_1800_n 0.00760397f $X=2.795 $Y=1.58 $X2=0
+ $Y2=0
cc_439 SCD N_A_268_467#_c_1800_n 0.0160518f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_440 N_SCD_c_510_n N_A_268_467#_c_1800_n 0.00343765f $X=2.795 $Y=1.745 $X2=0
+ $Y2=0
cc_441 N_SCD_c_508_n N_A_268_467#_c_1801_n 0.00259804f $X=2.795 $Y=1.58 $X2=0
+ $Y2=0
cc_442 SCD N_A_268_467#_c_1801_n 0.0153249f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_443 N_SCD_c_511_n N_A_268_467#_c_1802_n 0.00688395f $X=2.315 $Y=2.225 $X2=0
+ $Y2=0
cc_444 N_SCD_c_508_n N_A_268_467#_c_1802_n 0.0033915f $X=2.795 $Y=1.58 $X2=0
+ $Y2=0
cc_445 SCD N_A_268_467#_c_1802_n 0.0545353f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_446 N_SCD_c_510_n N_A_268_467#_c_1802_n 0.00437239f $X=2.795 $Y=1.745 $X2=0
+ $Y2=0
cc_447 N_SCD_c_506_n N_VGND_c_1983_n 0.0103655f $X=2.672 $Y=0.775 $X2=0 $Y2=0
cc_448 N_SCD_c_507_n N_VGND_c_1983_n 0.0015255f $X=2.672 $Y=0.925 $X2=0 $Y2=0
cc_449 N_SCD_c_506_n N_VGND_c_1996_n 0.003617f $X=2.672 $Y=0.775 $X2=0 $Y2=0
cc_450 N_SCD_c_506_n N_VGND_c_2012_n 0.0041518f $X=2.672 $Y=0.775 $X2=0 $Y2=0
cc_451 CLK N_A_629_47#_c_1179_n 0.0136301f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_452 N_CLK_c_565_n N_A_629_47#_c_1179_n 0.00437f $X=3.28 $Y=0.93 $X2=0 $Y2=0
cc_453 N_CLK_M1025_g N_A_629_47#_c_1180_n 0.0171492f $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_454 N_CLK_c_562_n N_A_629_47#_c_1181_n 0.00430217f $X=3.07 $Y=0.765 $X2=0
+ $Y2=0
cc_455 CLK N_A_629_47#_c_1181_n 0.0101544f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_456 N_CLK_c_565_n N_A_629_47#_c_1181_n 0.00127497f $X=3.28 $Y=0.93 $X2=0
+ $Y2=0
cc_457 N_CLK_M1025_g N_A_629_47#_c_1182_n 0.00486814f $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_458 CLK N_A_629_47#_c_1182_n 0.0115894f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_459 N_CLK_c_565_n N_A_629_47#_c_1182_n 0.00594439f $X=3.28 $Y=0.93 $X2=0
+ $Y2=0
cc_460 N_CLK_c_565_n N_A_629_47#_c_1183_n 0.00579939f $X=3.28 $Y=0.93 $X2=0
+ $Y2=0
cc_461 N_CLK_M1025_g N_VPWR_c_1638_n 0.00299045f $X=3.28 $Y=2.655 $X2=0 $Y2=0
cc_462 N_CLK_M1025_g N_VPWR_c_1654_n 0.00299821f $X=3.28 $Y=2.655 $X2=0 $Y2=0
cc_463 N_CLK_M1025_g N_VPWR_c_1627_n 0.0042382f $X=3.28 $Y=2.655 $X2=0 $Y2=0
cc_464 N_CLK_M1025_g N_A_268_467#_c_1806_n 0.0133408f $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_465 N_CLK_c_562_n N_A_268_467#_c_1797_n 4.17749e-19 $X=3.07 $Y=0.765 $X2=0
+ $Y2=0
cc_466 CLK N_A_268_467#_c_1797_n 0.00503449f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_467 N_CLK_M1025_g N_A_268_467#_c_1799_n 4.81379e-19 $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_468 CLK N_A_268_467#_c_1799_n 0.00672812f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_469 N_CLK_c_565_n N_A_268_467#_c_1799_n 5.83394e-19 $X=3.28 $Y=0.93 $X2=0
+ $Y2=0
cc_470 N_CLK_M1025_g N_A_268_467#_c_1800_n 0.00489948f $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_471 CLK N_A_268_467#_c_1800_n 0.0187013f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_472 N_CLK_c_565_n N_A_268_467#_c_1800_n 0.00589607f $X=3.28 $Y=0.93 $X2=0
+ $Y2=0
cc_473 N_CLK_M1025_g N_A_268_467#_c_1802_n 0.0255981f $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_474 N_CLK_M1025_g N_A_268_467#_c_1808_n 0.0139427f $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_475 N_CLK_M1025_g N_A_268_467#_c_1809_n 0.00281736f $X=3.28 $Y=2.655 $X2=0
+ $Y2=0
cc_476 N_CLK_c_562_n N_VGND_c_1983_n 0.00945238f $X=3.07 $Y=0.765 $X2=0 $Y2=0
cc_477 CLK N_VGND_c_1983_n 0.00128977f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_478 N_CLK_c_562_n N_VGND_c_1998_n 0.00486043f $X=3.07 $Y=0.765 $X2=0 $Y2=0
cc_479 N_CLK_c_565_n N_VGND_c_1998_n 8.7631e-19 $X=3.28 $Y=0.93 $X2=0 $Y2=0
cc_480 N_CLK_c_562_n N_VGND_c_2012_n 0.00586712f $X=3.07 $Y=0.765 $X2=0 $Y2=0
cc_481 CLK N_VGND_c_2012_n 0.00570205f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_482 N_CLK_c_565_n N_VGND_c_2012_n 0.0010536f $X=3.28 $Y=0.93 $X2=0 $Y2=0
cc_483 N_A_920_73#_M1019_g N_A_1291_93#_c_762_n 0.0485918f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_484 N_A_920_73#_M1001_g N_A_1291_93#_c_769_n 0.00435398f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_485 N_A_920_73#_c_609_n N_A_1291_93#_c_769_n 0.0059473f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_486 N_A_920_73#_c_616_n N_A_1291_93#_c_769_n 0.00126329f $X=6.17 $Y=1.68
+ $X2=0 $Y2=0
cc_487 N_A_920_73#_M1019_g N_A_1291_93#_c_763_n 0.00724969f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_488 N_A_920_73#_c_609_n N_A_1291_93#_c_763_n 0.0112104f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_489 N_A_920_73#_c_610_n N_A_1291_93#_c_763_n 0.00126511f $X=6.43 $Y=1.635
+ $X2=0 $Y2=0
cc_490 N_A_920_73#_c_616_n N_A_1291_93#_c_763_n 0.0164248f $X=6.17 $Y=1.68 $X2=0
+ $Y2=0
cc_491 N_A_920_73#_c_609_n N_A_1291_93#_c_764_n 0.00113101f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_492 N_A_920_73#_M1001_g N_A_1291_93#_c_771_n 3.09558e-19 $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_493 N_A_920_73#_c_609_n N_A_1291_93#_c_771_n 0.0242623f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_494 N_A_920_73#_M1043_g N_A_1291_93#_c_773_n 0.00696222f $X=9.445 $Y=2.67
+ $X2=0 $Y2=0
cc_495 N_A_920_73#_c_623_n N_A_1291_93#_c_773_n 0.0465451f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_496 N_A_920_73#_c_612_n N_A_1291_93#_c_773_n 0.00475191f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_497 N_A_920_73#_M1041_g N_A_1291_93#_c_766_n 0.0142711f $X=9.045 $Y=0.915
+ $X2=0 $Y2=0
cc_498 N_A_920_73#_c_607_n N_A_1291_93#_c_766_n 0.00279887f $X=9.37 $Y=1.625
+ $X2=0 $Y2=0
cc_499 N_A_920_73#_c_611_n N_A_1291_93#_c_766_n 0.0146993f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_500 N_A_920_73#_c_612_n N_A_1291_93#_c_766_n 0.002095f $X=9.05 $Y=1.535 $X2=0
+ $Y2=0
cc_501 N_A_920_73#_M1041_g N_A_1291_93#_c_767_n 0.00563211f $X=9.045 $Y=0.915
+ $X2=0 $Y2=0
cc_502 N_A_920_73#_c_607_n N_A_1291_93#_c_767_n 0.0102729f $X=9.37 $Y=1.625
+ $X2=0 $Y2=0
cc_503 N_A_920_73#_M1043_g N_A_1291_93#_c_767_n 0.0128303f $X=9.445 $Y=2.67
+ $X2=0 $Y2=0
cc_504 N_A_920_73#_c_623_n N_A_1291_93#_c_767_n 0.0136416f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_505 N_A_920_73#_c_611_n N_A_1291_93#_c_767_n 0.0358132f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_506 N_A_920_73#_c_612_n N_A_1291_93#_c_767_n 0.00209509f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_507 N_A_920_73#_c_609_n N_A_1291_93#_c_775_n 0.0111986f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_508 N_A_920_73#_c_615_n N_A_1291_93#_c_777_n 0.010592f $X=8.13 $Y=1.635 $X2=0
+ $Y2=0
cc_509 N_A_920_73#_c_623_n N_A_1291_93#_c_804_n 0.00406017f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_510 N_A_920_73#_c_611_n N_A_1291_93#_c_804_n 0.00227419f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_511 N_A_920_73#_c_612_n N_A_1291_93#_c_804_n 2.05478e-19 $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_512 N_A_920_73#_c_609_n N_A_1163_119#_M1003_g 0.0135657f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_513 N_A_920_73#_c_623_n N_A_1163_119#_M1013_g 0.0103447f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_514 N_A_920_73#_c_611_n N_A_1163_119#_M1013_g 0.00295826f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_515 N_A_920_73#_c_612_n N_A_1163_119#_M1013_g 7.3937e-19 $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_516 N_A_920_73#_c_615_n N_A_1163_119#_M1013_g 0.00242094f $X=8.13 $Y=1.635
+ $X2=0 $Y2=0
cc_517 N_A_920_73#_M1041_g N_A_1163_119#_c_915_n 0.0363547f $X=9.045 $Y=0.915
+ $X2=0 $Y2=0
cc_518 N_A_920_73#_M1019_g N_A_1163_119#_c_916_n 0.00989281f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_519 N_A_920_73#_M1001_g N_A_1163_119#_c_926_n 0.00136222f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_520 N_A_920_73#_M1041_g N_A_1163_119#_c_917_n 8.25101e-19 $X=9.045 $Y=0.915
+ $X2=0 $Y2=0
cc_521 N_A_920_73#_c_623_n N_A_1163_119#_c_917_n 0.00479203f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_522 N_A_920_73#_c_611_n N_A_1163_119#_c_917_n 2.42097e-19 $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_523 N_A_920_73#_c_615_n N_A_1163_119#_c_917_n 0.0134731f $X=8.13 $Y=1.635
+ $X2=0 $Y2=0
cc_524 N_A_920_73#_c_623_n N_A_1163_119#_c_927_n 0.0124821f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_525 N_A_920_73#_c_611_n N_A_1163_119#_c_927_n 0.0130847f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_526 N_A_920_73#_c_612_n N_A_1163_119#_c_927_n 0.00101117f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_527 N_A_920_73#_c_615_n N_A_1163_119#_c_927_n 0.00937335f $X=8.13 $Y=1.635
+ $X2=0 $Y2=0
cc_528 N_A_920_73#_c_623_n N_A_1163_119#_c_918_n 0.00505558f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_529 N_A_920_73#_c_611_n N_A_1163_119#_c_918_n 0.00116981f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_530 N_A_920_73#_c_612_n N_A_1163_119#_c_918_n 0.017615f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_531 N_A_920_73#_c_615_n N_A_1163_119#_c_918_n 9.72842e-19 $X=8.13 $Y=1.635
+ $X2=0 $Y2=0
cc_532 N_A_920_73#_M1019_g N_A_1163_119#_c_919_n 0.00508391f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_533 N_A_920_73#_c_616_n N_A_1163_119#_c_919_n 2.11952e-19 $X=6.17 $Y=1.68
+ $X2=0 $Y2=0
cc_534 N_A_920_73#_M1001_g N_A_1163_119#_c_920_n 0.00526863f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_535 N_A_920_73#_M1019_g N_A_1163_119#_c_920_n 0.00636908f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_536 N_A_920_73#_c_610_n N_A_1163_119#_c_920_n 0.0249531f $X=6.43 $Y=1.635
+ $X2=0 $Y2=0
cc_537 N_A_920_73#_c_616_n N_A_1163_119#_c_920_n 0.0117572f $X=6.17 $Y=1.68
+ $X2=0 $Y2=0
cc_538 N_A_920_73#_M1001_g N_A_1163_119#_c_930_n 0.0115674f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_539 N_A_920_73#_c_610_n N_A_1163_119#_c_930_n 0.00695518f $X=6.43 $Y=1.635
+ $X2=0 $Y2=0
cc_540 N_A_920_73#_c_616_n N_A_1163_119#_c_930_n 0.00623512f $X=6.17 $Y=1.68
+ $X2=0 $Y2=0
cc_541 N_A_920_73#_c_609_n N_A_1163_119#_c_921_n 0.0049889f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_542 N_A_920_73#_M1019_g N_A_1163_119#_c_922_n 0.0123367f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_543 N_A_920_73#_c_609_n N_A_1163_119#_c_922_n 0.0497508f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_544 N_A_920_73#_c_610_n N_A_1163_119#_c_922_n 0.0200037f $X=6.43 $Y=1.635
+ $X2=0 $Y2=0
cc_545 N_A_920_73#_c_616_n N_A_1163_119#_c_922_n 0.00128623f $X=6.17 $Y=1.68
+ $X2=0 $Y2=0
cc_546 N_A_920_73#_c_609_n N_A_1163_119#_c_923_n 0.0619067f $X=8.045 $Y=1.635
+ $X2=0 $Y2=0
cc_547 N_A_920_73#_c_609_n N_SET_B_M1024_g 0.011839f $X=8.045 $Y=1.635 $X2=0
+ $Y2=0
cc_548 N_A_920_73#_c_615_n N_SET_B_M1024_g 0.0060177f $X=8.13 $Y=1.635 $X2=0
+ $Y2=0
cc_549 N_A_920_73#_M1043_g N_SET_B_c_1055_n 0.00247177f $X=9.445 $Y=2.67 $X2=0
+ $Y2=0
cc_550 N_A_920_73#_c_609_n N_SET_B_c_1055_n 0.00620214f $X=8.045 $Y=1.635 $X2=0
+ $Y2=0
cc_551 N_A_920_73#_c_623_n N_SET_B_c_1055_n 0.0347839f $X=8.885 $Y=1.94 $X2=0
+ $Y2=0
cc_552 N_A_920_73#_c_612_n N_SET_B_c_1055_n 0.00362346f $X=9.05 $Y=1.535 $X2=0
+ $Y2=0
cc_553 N_A_920_73#_c_615_n N_SET_B_c_1055_n 0.00580558f $X=8.13 $Y=1.635 $X2=0
+ $Y2=0
cc_554 N_A_920_73#_c_609_n N_SET_B_c_1056_n 0.00206217f $X=8.045 $Y=1.635 $X2=0
+ $Y2=0
cc_555 N_A_920_73#_c_609_n N_SET_B_c_1059_n 0.0410575f $X=8.045 $Y=1.635 $X2=0
+ $Y2=0
cc_556 N_A_920_73#_c_615_n N_SET_B_c_1059_n 0.008943f $X=8.13 $Y=1.635 $X2=0
+ $Y2=0
cc_557 N_A_920_73#_c_609_n N_SET_B_c_1060_n 0.00686585f $X=8.045 $Y=1.635 $X2=0
+ $Y2=0
cc_558 N_A_920_73#_c_608_n N_A_629_47#_M1033_g 0.0100821f $X=4.74 $Y=0.565 $X2=0
+ $Y2=0
cc_559 N_A_920_73#_c_613_n N_A_629_47#_M1006_g 0.034913f $X=5.21 $Y=1.65 $X2=0
+ $Y2=0
cc_560 N_A_920_73#_c_608_n N_A_629_47#_c_1173_n 0.00488572f $X=4.74 $Y=0.565
+ $X2=0 $Y2=0
cc_561 N_A_920_73#_M1001_g N_A_629_47#_c_1185_n 0.0104164f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_562 N_A_920_73#_c_617_n N_A_629_47#_M1039_g 0.00504415f $X=5.795 $Y=1.77
+ $X2=0 $Y2=0
cc_563 N_A_920_73#_M1019_g N_A_629_47#_M1039_g 0.0131514f $X=6.17 $Y=0.805 $X2=0
+ $Y2=0
cc_564 N_A_920_73#_M1019_g N_A_629_47#_c_1176_n 0.0103162f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_565 N_A_920_73#_M1041_g N_A_629_47#_c_1176_n 0.0104164f $X=9.045 $Y=0.915
+ $X2=0 $Y2=0
cc_566 N_A_920_73#_M1001_g N_A_629_47#_M1026_g 0.0131778f $X=5.87 $Y=2.525 $X2=0
+ $Y2=0
cc_567 N_A_920_73#_c_610_n N_A_629_47#_M1026_g 9.36651e-19 $X=6.43 $Y=1.635
+ $X2=0 $Y2=0
cc_568 N_A_920_73#_c_616_n N_A_629_47#_M1026_g 0.00545952f $X=6.17 $Y=1.68 $X2=0
+ $Y2=0
cc_569 N_A_920_73#_M1043_g N_A_629_47#_M1031_g 0.0299718f $X=9.445 $Y=2.67 $X2=0
+ $Y2=0
cc_570 N_A_920_73#_c_623_n N_A_629_47#_M1031_g 0.00709238f $X=8.885 $Y=1.94
+ $X2=0 $Y2=0
cc_571 N_A_920_73#_c_612_n N_A_629_47#_M1031_g 0.00717607f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_572 N_A_920_73#_M1041_g N_A_629_47#_M1032_g 0.0104325f $X=9.045 $Y=0.915
+ $X2=0 $Y2=0
cc_573 N_A_920_73#_c_607_n N_A_629_47#_M1032_g 0.00102543f $X=9.37 $Y=1.625
+ $X2=0 $Y2=0
cc_574 N_A_920_73#_c_608_n N_A_629_47#_c_1181_n 0.00499444f $X=4.74 $Y=0.565
+ $X2=0 $Y2=0
cc_575 N_A_920_73#_c_608_n N_A_629_47#_c_1182_n 0.0470966f $X=4.74 $Y=0.565
+ $X2=0 $Y2=0
cc_576 N_A_920_73#_c_613_n N_A_629_47#_c_1182_n 0.00671663f $X=5.21 $Y=1.65
+ $X2=0 $Y2=0
cc_577 N_A_920_73#_c_608_n N_A_629_47#_c_1183_n 0.0216077f $X=4.74 $Y=0.565
+ $X2=0 $Y2=0
cc_578 N_A_920_73#_c_613_n N_A_629_47#_c_1183_n 0.00272782f $X=5.21 $Y=1.65
+ $X2=0 $Y2=0
cc_579 N_A_920_73#_c_614_n N_A_629_47#_c_1183_n 0.0133243f $X=5.21 $Y=1.65 $X2=0
+ $Y2=0
cc_580 N_A_920_73#_c_612_n N_A_1946_369#_M1038_g 0.00184666f $X=9.05 $Y=1.535
+ $X2=0 $Y2=0
cc_581 N_A_920_73#_c_607_n N_A_1946_369#_c_1310_n 0.00928678f $X=9.37 $Y=1.625
+ $X2=0 $Y2=0
cc_582 N_A_920_73#_M1043_g N_A_1946_369#_c_1310_n 0.0718584f $X=9.445 $Y=2.67
+ $X2=0 $Y2=0
cc_583 N_A_920_73#_M1043_g N_A_1799_408#_c_1414_n 0.0166143f $X=9.445 $Y=2.67
+ $X2=0 $Y2=0
cc_584 N_A_920_73#_c_607_n N_A_1799_408#_c_1405_n 6.11233e-19 $X=9.37 $Y=1.625
+ $X2=0 $Y2=0
cc_585 N_A_920_73#_M1041_g N_A_1799_408#_c_1406_n 4.37238e-19 $X=9.045 $Y=0.915
+ $X2=0 $Y2=0
cc_586 N_A_920_73#_c_607_n N_A_1799_408#_c_1406_n 0.003615f $X=9.37 $Y=1.625
+ $X2=0 $Y2=0
cc_587 N_A_920_73#_M1043_g N_A_1799_408#_c_1416_n 0.00387812f $X=9.445 $Y=2.67
+ $X2=0 $Y2=0
cc_588 N_A_920_73#_M1043_g N_A_1799_408#_c_1421_n 0.00109343f $X=9.445 $Y=2.67
+ $X2=0 $Y2=0
cc_589 N_A_920_73#_c_623_n N_VPWR_M1030_d 4.84848e-19 $X=8.885 $Y=1.94 $X2=0
+ $Y2=0
cc_590 N_A_920_73#_c_615_n N_VPWR_M1030_d 0.00127784f $X=8.13 $Y=1.635 $X2=0
+ $Y2=0
cc_591 N_A_920_73#_M1043_g N_VPWR_c_1642_n 0.00380912f $X=9.445 $Y=2.67 $X2=0
+ $Y2=0
cc_592 N_A_920_73#_M1001_g N_VPWR_c_1627_n 9.39239e-19 $X=5.87 $Y=2.525 $X2=0
+ $Y2=0
cc_593 N_A_920_73#_M1043_g N_VPWR_c_1627_n 0.00520574f $X=9.445 $Y=2.67 $X2=0
+ $Y2=0
cc_594 N_A_920_73#_M1006_d N_A_268_467#_c_1810_n 0.00572003f $X=4.6 $Y=1.945
+ $X2=0 $Y2=0
cc_595 N_A_920_73#_c_617_n N_A_268_467#_c_1810_n 2.32303e-19 $X=5.795 $Y=1.77
+ $X2=0 $Y2=0
cc_596 N_A_920_73#_c_613_n N_A_268_467#_c_1810_n 0.0547894f $X=5.21 $Y=1.65
+ $X2=0 $Y2=0
cc_597 N_A_920_73#_c_614_n N_A_268_467#_c_1810_n 0.00494739f $X=5.21 $Y=1.65
+ $X2=0 $Y2=0
cc_598 N_A_920_73#_c_608_n N_A_268_467#_c_1803_n 0.0248611f $X=4.74 $Y=0.565
+ $X2=0 $Y2=0
cc_599 N_A_920_73#_c_617_n N_A_268_467#_c_1804_n 0.0152623f $X=5.795 $Y=1.77
+ $X2=0 $Y2=0
cc_600 N_A_920_73#_M1001_g N_A_268_467#_c_1804_n 0.00598396f $X=5.87 $Y=2.525
+ $X2=0 $Y2=0
cc_601 N_A_920_73#_M1019_g N_A_268_467#_c_1804_n 0.00110501f $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_602 N_A_920_73#_c_608_n N_A_268_467#_c_1804_n 0.00857917f $X=4.74 $Y=0.565
+ $X2=0 $Y2=0
cc_603 N_A_920_73#_c_613_n N_A_268_467#_c_1804_n 0.0517973f $X=5.21 $Y=1.65
+ $X2=0 $Y2=0
cc_604 N_A_920_73#_c_614_n N_A_268_467#_c_1804_n 0.00552066f $X=5.21 $Y=1.65
+ $X2=0 $Y2=0
cc_605 N_A_920_73#_c_617_n N_A_268_467#_c_1805_n 2.9533e-19 $X=5.795 $Y=1.77
+ $X2=0 $Y2=0
cc_606 N_A_920_73#_M1019_g N_A_268_467#_c_1805_n 8.59694e-19 $X=6.17 $Y=0.805
+ $X2=0 $Y2=0
cc_607 N_A_920_73#_c_614_n N_A_268_467#_c_1805_n 6.03365e-19 $X=5.21 $Y=1.65
+ $X2=0 $Y2=0
cc_608 N_A_920_73#_c_617_n N_A_268_467#_c_1813_n 0.00130195f $X=5.795 $Y=1.77
+ $X2=0 $Y2=0
cc_609 N_A_920_73#_c_623_n A_1697_379# 9.68801e-19 $X=8.885 $Y=1.94 $X2=-0.19
+ $Y2=-0.245
cc_610 N_A_920_73#_M1019_g N_VGND_c_1985_n 0.00177594f $X=6.17 $Y=0.805 $X2=0
+ $Y2=0
cc_611 N_A_920_73#_c_608_n N_VGND_c_2000_n 0.0104813f $X=4.74 $Y=0.565 $X2=0
+ $Y2=0
cc_612 N_A_920_73#_M1019_g N_VGND_c_2012_n 9.39239e-19 $X=6.17 $Y=0.805 $X2=0
+ $Y2=0
cc_613 N_A_920_73#_M1041_g N_VGND_c_2012_n 9.39239e-19 $X=9.045 $Y=0.915 $X2=0
+ $Y2=0
cc_614 N_A_920_73#_c_608_n N_VGND_c_2012_n 0.0102908f $X=4.74 $Y=0.565 $X2=0
+ $Y2=0
cc_615 N_A_1291_93#_c_769_n N_A_1163_119#_M1003_g 0.0385637f $X=6.66 $Y=2.205
+ $X2=0 $Y2=0
cc_616 N_A_1291_93#_c_763_n N_A_1163_119#_M1003_g 0.0126038f $X=6.74 $Y=1.825
+ $X2=0 $Y2=0
cc_617 N_A_1291_93#_c_771_n N_A_1163_119#_M1003_g 0.0034893f $X=6.8 $Y=1.99
+ $X2=0 $Y2=0
cc_618 N_A_1291_93#_c_775_n N_A_1163_119#_M1003_g 0.00881125f $X=7.3 $Y=2.495
+ $X2=0 $Y2=0
cc_619 N_A_1291_93#_c_776_n N_A_1163_119#_M1003_g 0.00549076f $X=7.63 $Y=2.495
+ $X2=0 $Y2=0
cc_620 N_A_1291_93#_c_812_p N_A_1163_119#_c_914_n 0.0123278f $X=7.79 $Y=0.837
+ $X2=0 $Y2=0
cc_621 N_A_1291_93#_c_768_n N_A_1163_119#_c_914_n 0.00177462f $X=7.96 $Y=0.837
+ $X2=0 $Y2=0
cc_622 N_A_1291_93#_c_773_n N_A_1163_119#_M1013_g 0.0150259f $X=9.315 $Y=2.29
+ $X2=0 $Y2=0
cc_623 N_A_1291_93#_c_777_n N_A_1163_119#_M1013_g 0.00279844f $X=8.13 $Y=2.29
+ $X2=0 $Y2=0
cc_624 N_A_1291_93#_c_765_n N_A_1163_119#_c_915_n 0.0140714f $X=8.745 $Y=0.95
+ $X2=0 $Y2=0
cc_625 N_A_1291_93#_c_768_n N_A_1163_119#_c_915_n 8.34682e-19 $X=7.96 $Y=0.837
+ $X2=0 $Y2=0
cc_626 N_A_1291_93#_c_804_n N_A_1163_119#_c_915_n 0.00422463f $X=8.83 $Y=0.95
+ $X2=0 $Y2=0
cc_627 N_A_1291_93#_c_762_n N_A_1163_119#_c_916_n 0.00175436f $X=6.53 $Y=1.125
+ $X2=0 $Y2=0
cc_628 N_A_1291_93#_c_820_p N_A_1163_119#_c_926_n 0.00696295f $X=6.965 $Y=2.385
+ $X2=0 $Y2=0
cc_629 N_A_1291_93#_c_765_n N_A_1163_119#_c_917_n 0.0102525f $X=8.745 $Y=0.95
+ $X2=0 $Y2=0
cc_630 N_A_1291_93#_c_812_p N_A_1163_119#_c_917_n 0.0147625f $X=7.79 $Y=0.837
+ $X2=0 $Y2=0
cc_631 N_A_1291_93#_c_768_n N_A_1163_119#_c_917_n 0.0438326f $X=7.96 $Y=0.837
+ $X2=0 $Y2=0
cc_632 N_A_1291_93#_c_765_n N_A_1163_119#_c_918_n 9.59778e-19 $X=8.745 $Y=0.95
+ $X2=0 $Y2=0
cc_633 N_A_1291_93#_c_769_n N_A_1163_119#_c_920_n 0.00132584f $X=6.66 $Y=2.205
+ $X2=0 $Y2=0
cc_634 N_A_1291_93#_c_771_n N_A_1163_119#_c_920_n 0.00177981f $X=6.8 $Y=1.99
+ $X2=0 $Y2=0
cc_635 N_A_1291_93#_c_769_n N_A_1163_119#_c_930_n 0.00342005f $X=6.66 $Y=2.205
+ $X2=0 $Y2=0
cc_636 N_A_1291_93#_c_771_n N_A_1163_119#_c_930_n 0.0116451f $X=6.8 $Y=1.99
+ $X2=0 $Y2=0
cc_637 N_A_1291_93#_c_764_n N_A_1163_119#_c_921_n 0.0126038f $X=6.74 $Y=1.2
+ $X2=0 $Y2=0
cc_638 N_A_1291_93#_c_812_p N_A_1163_119#_c_921_n 0.00581201f $X=7.79 $Y=0.837
+ $X2=0 $Y2=0
cc_639 N_A_1291_93#_c_763_n N_A_1163_119#_c_922_n 0.00525495f $X=6.74 $Y=1.825
+ $X2=0 $Y2=0
cc_640 N_A_1291_93#_c_764_n N_A_1163_119#_c_922_n 0.0176879f $X=6.74 $Y=1.2
+ $X2=0 $Y2=0
cc_641 N_A_1291_93#_c_812_p N_A_1163_119#_c_923_n 0.0165944f $X=7.79 $Y=0.837
+ $X2=0 $Y2=0
cc_642 N_A_1291_93#_c_772_n N_SET_B_M1030_g 0.00749562f $X=8.045 $Y=2.385 $X2=0
+ $Y2=0
cc_643 N_A_1291_93#_c_776_n N_SET_B_M1030_g 0.00954683f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_644 N_A_1291_93#_c_777_n N_SET_B_M1030_g 0.00214371f $X=8.13 $Y=2.29 $X2=0
+ $Y2=0
cc_645 N_A_1291_93#_c_765_n N_SET_B_M1024_g 0.0053815f $X=8.745 $Y=0.95 $X2=0
+ $Y2=0
cc_646 N_A_1291_93#_c_768_n N_SET_B_M1024_g 0.0135573f $X=7.96 $Y=0.837 $X2=0
+ $Y2=0
cc_647 N_A_1291_93#_c_772_n N_SET_B_c_1055_n 0.0048351f $X=8.045 $Y=2.385 $X2=0
+ $Y2=0
cc_648 N_A_1291_93#_c_773_n N_SET_B_c_1055_n 0.0325411f $X=9.315 $Y=2.29 $X2=0
+ $Y2=0
cc_649 N_A_1291_93#_c_767_n N_SET_B_c_1055_n 0.0175662f $X=9.4 $Y=2.205 $X2=0
+ $Y2=0
cc_650 N_A_1291_93#_c_776_n N_SET_B_c_1055_n 0.00198458f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_651 N_A_1291_93#_c_777_n N_SET_B_c_1055_n 0.00467138f $X=8.13 $Y=2.29 $X2=0
+ $Y2=0
cc_652 N_A_1291_93#_c_771_n N_SET_B_c_1056_n 0.00208971f $X=6.8 $Y=1.99 $X2=0
+ $Y2=0
cc_653 N_A_1291_93#_c_775_n N_SET_B_c_1056_n 0.00797915f $X=7.3 $Y=2.495 $X2=0
+ $Y2=0
cc_654 N_A_1291_93#_c_769_n N_SET_B_c_1059_n 7.38407e-19 $X=6.66 $Y=2.205 $X2=0
+ $Y2=0
cc_655 N_A_1291_93#_c_771_n N_SET_B_c_1059_n 0.00969171f $X=6.8 $Y=1.99 $X2=0
+ $Y2=0
cc_656 N_A_1291_93#_c_775_n N_SET_B_c_1059_n 0.0402788f $X=7.3 $Y=2.495 $X2=0
+ $Y2=0
cc_657 N_A_1291_93#_c_772_n N_SET_B_c_1060_n 0.00712114f $X=8.045 $Y=2.385 $X2=0
+ $Y2=0
cc_658 N_A_1291_93#_c_776_n N_SET_B_c_1060_n 0.00165016f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_659 N_A_1291_93#_c_762_n N_A_629_47#_c_1176_n 0.0103107f $X=6.53 $Y=1.125
+ $X2=0 $Y2=0
cc_660 N_A_1291_93#_c_765_n N_A_629_47#_c_1176_n 0.00468275f $X=8.745 $Y=0.95
+ $X2=0 $Y2=0
cc_661 N_A_1291_93#_c_812_p N_A_629_47#_c_1176_n 0.0078914f $X=7.79 $Y=0.837
+ $X2=0 $Y2=0
cc_662 N_A_1291_93#_c_768_n N_A_629_47#_c_1176_n 2.57061e-19 $X=7.96 $Y=0.837
+ $X2=0 $Y2=0
cc_663 N_A_1291_93#_c_804_n N_A_629_47#_c_1176_n 0.00395037f $X=8.83 $Y=0.95
+ $X2=0 $Y2=0
cc_664 N_A_1291_93#_c_769_n N_A_629_47#_M1026_g 0.0401248f $X=6.66 $Y=2.205
+ $X2=0 $Y2=0
cc_665 N_A_1291_93#_c_771_n N_A_629_47#_M1026_g 3.51659e-19 $X=6.8 $Y=1.99 $X2=0
+ $Y2=0
cc_666 N_A_1291_93#_c_820_p N_A_629_47#_M1026_g 5.20381e-19 $X=6.965 $Y=2.385
+ $X2=0 $Y2=0
cc_667 N_A_1291_93#_c_769_n N_A_629_47#_c_1188_n 0.0101854f $X=6.66 $Y=2.205
+ $X2=0 $Y2=0
cc_668 N_A_1291_93#_c_820_p N_A_629_47#_c_1188_n 8.71037e-19 $X=6.965 $Y=2.385
+ $X2=0 $Y2=0
cc_669 N_A_1291_93#_c_772_n N_A_629_47#_c_1188_n 0.00430896f $X=8.045 $Y=2.385
+ $X2=0 $Y2=0
cc_670 N_A_1291_93#_c_775_n N_A_629_47#_c_1188_n 8.3992e-19 $X=7.3 $Y=2.495
+ $X2=0 $Y2=0
cc_671 N_A_1291_93#_c_776_n N_A_629_47#_c_1188_n 0.00473617f $X=7.63 $Y=2.495
+ $X2=0 $Y2=0
cc_672 N_A_1291_93#_c_777_n N_A_629_47#_c_1188_n 5.12858e-19 $X=8.13 $Y=2.29
+ $X2=0 $Y2=0
cc_673 N_A_1291_93#_c_773_n N_A_629_47#_M1031_g 0.0150243f $X=9.315 $Y=2.29
+ $X2=0 $Y2=0
cc_674 N_A_1291_93#_c_767_n N_A_629_47#_M1031_g 0.00306066f $X=9.4 $Y=2.205
+ $X2=0 $Y2=0
cc_675 N_A_1291_93#_c_766_n N_A_629_47#_M1032_g 0.00117313f $X=9.315 $Y=1.115
+ $X2=0 $Y2=0
cc_676 N_A_1291_93#_c_767_n N_A_1946_369#_c_1310_n 4.50524e-19 $X=9.4 $Y=2.205
+ $X2=0 $Y2=0
cc_677 N_A_1291_93#_c_766_n N_A_1799_408#_M1041_d 0.00475134f $X=9.315 $Y=1.115
+ $X2=-0.19 $Y2=-0.245
cc_678 N_A_1291_93#_c_767_n N_A_1799_408#_M1041_d 5.16052e-19 $X=9.4 $Y=2.205
+ $X2=-0.19 $Y2=-0.245
cc_679 N_A_1291_93#_c_773_n N_A_1799_408#_M1031_d 0.00377277f $X=9.315 $Y=2.29
+ $X2=0 $Y2=0
cc_680 N_A_1291_93#_c_773_n N_A_1799_408#_c_1414_n 0.030633f $X=9.315 $Y=2.29
+ $X2=0 $Y2=0
cc_681 N_A_1291_93#_c_766_n N_A_1799_408#_c_1405_n 0.0229619f $X=9.315 $Y=1.115
+ $X2=0 $Y2=0
cc_682 N_A_1291_93#_c_766_n N_A_1799_408#_c_1406_n 0.013583f $X=9.315 $Y=1.115
+ $X2=0 $Y2=0
cc_683 N_A_1291_93#_c_767_n N_A_1799_408#_c_1406_n 0.0659953f $X=9.4 $Y=2.205
+ $X2=0 $Y2=0
cc_684 N_A_1291_93#_c_773_n N_A_1799_408#_c_1416_n 0.00302417f $X=9.315 $Y=2.29
+ $X2=0 $Y2=0
cc_685 N_A_1291_93#_c_773_n N_A_1799_408#_c_1421_n 0.0110966f $X=9.315 $Y=2.29
+ $X2=0 $Y2=0
cc_686 N_A_1291_93#_c_767_n N_A_1799_408#_c_1421_n 0.00383202f $X=9.4 $Y=2.205
+ $X2=0 $Y2=0
cc_687 N_A_1291_93#_c_820_p N_VPWR_M1034_d 0.00194695f $X=6.965 $Y=2.385 $X2=0
+ $Y2=0
cc_688 N_A_1291_93#_c_775_n N_VPWR_M1034_d 0.00159635f $X=7.3 $Y=2.495 $X2=0
+ $Y2=0
cc_689 N_A_1291_93#_c_772_n N_VPWR_M1030_d 0.00348296f $X=8.045 $Y=2.385 $X2=0
+ $Y2=0
cc_690 N_A_1291_93#_c_773_n N_VPWR_M1030_d 0.00187785f $X=9.315 $Y=2.29 $X2=0
+ $Y2=0
cc_691 N_A_1291_93#_c_777_n N_VPWR_M1030_d 0.00612902f $X=8.13 $Y=2.29 $X2=0
+ $Y2=0
cc_692 N_A_1291_93#_c_769_n N_VPWR_c_1630_n 0.00510427f $X=6.66 $Y=2.205 $X2=0
+ $Y2=0
cc_693 N_A_1291_93#_c_820_p N_VPWR_c_1630_n 0.0150492f $X=6.965 $Y=2.385 $X2=0
+ $Y2=0
cc_694 N_A_1291_93#_c_775_n N_VPWR_c_1630_n 0.0121604f $X=7.3 $Y=2.495 $X2=0
+ $Y2=0
cc_695 N_A_1291_93#_c_772_n N_VPWR_c_1631_n 0.00723305f $X=8.045 $Y=2.385 $X2=0
+ $Y2=0
cc_696 N_A_1291_93#_c_773_n N_VPWR_c_1631_n 0.0033515f $X=9.315 $Y=2.29 $X2=0
+ $Y2=0
cc_697 N_A_1291_93#_c_776_n N_VPWR_c_1631_n 0.00234875f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_698 N_A_1291_93#_c_777_n N_VPWR_c_1631_n 0.0134073f $X=8.13 $Y=2.29 $X2=0
+ $Y2=0
cc_699 N_A_1291_93#_c_776_n N_VPWR_c_1640_n 0.00496982f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_700 N_A_1291_93#_c_769_n N_VPWR_c_1627_n 9.39239e-19 $X=6.66 $Y=2.205 $X2=0
+ $Y2=0
cc_701 N_A_1291_93#_c_820_p N_VPWR_c_1627_n 0.0055517f $X=6.965 $Y=2.385 $X2=0
+ $Y2=0
cc_702 N_A_1291_93#_c_772_n N_VPWR_c_1627_n 0.00955131f $X=8.045 $Y=2.385 $X2=0
+ $Y2=0
cc_703 N_A_1291_93#_c_775_n N_VPWR_c_1627_n 0.00551049f $X=7.3 $Y=2.495 $X2=0
+ $Y2=0
cc_704 N_A_1291_93#_c_776_n N_VPWR_c_1627_n 0.00834044f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_705 N_A_1291_93#_c_777_n N_VPWR_c_1627_n 5.43685e-19 $X=8.13 $Y=2.29 $X2=0
+ $Y2=0
cc_706 N_A_1291_93#_c_773_n A_1697_379# 0.0116703f $X=9.315 $Y=2.29 $X2=-0.19
+ $Y2=-0.245
cc_707 N_A_1291_93#_c_765_n N_VGND_M1024_d 0.00888018f $X=8.745 $Y=0.95 $X2=0
+ $Y2=0
cc_708 N_A_1291_93#_c_762_n N_VGND_c_1985_n 0.0117736f $X=6.53 $Y=1.125 $X2=0
+ $Y2=0
cc_709 N_A_1291_93#_c_764_n N_VGND_c_1985_n 0.00520024f $X=6.74 $Y=1.2 $X2=0
+ $Y2=0
cc_710 N_A_1291_93#_c_812_p N_VGND_c_1985_n 0.0171493f $X=7.79 $Y=0.837 $X2=0
+ $Y2=0
cc_711 N_A_1291_93#_c_765_n N_VGND_c_1986_n 0.0266042f $X=8.745 $Y=0.95 $X2=0
+ $Y2=0
cc_712 N_A_1291_93#_c_768_n N_VGND_c_1986_n 0.00426821f $X=7.96 $Y=0.837 $X2=0
+ $Y2=0
cc_713 N_A_1291_93#_c_812_p N_VGND_c_2004_n 0.0109953f $X=7.79 $Y=0.837 $X2=0
+ $Y2=0
cc_714 N_A_1291_93#_c_762_n N_VGND_c_2012_n 7.88961e-19 $X=6.53 $Y=1.125 $X2=0
+ $Y2=0
cc_715 N_A_1291_93#_c_812_p N_VGND_c_2012_n 0.0175771f $X=7.79 $Y=0.837 $X2=0
+ $Y2=0
cc_716 N_A_1291_93#_c_804_n N_VGND_c_2012_n 0.005401f $X=8.83 $Y=0.95 $X2=0
+ $Y2=0
cc_717 N_A_1291_93#_c_812_p A_1530_119# 0.00219687f $X=7.79 $Y=0.837 $X2=-0.19
+ $Y2=-0.245
cc_718 N_A_1291_93#_c_768_n A_1530_119# 7.91627e-19 $X=7.96 $Y=0.837 $X2=-0.19
+ $Y2=-0.245
cc_719 N_A_1291_93#_c_765_n A_1735_119# 0.00112168f $X=8.745 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_720 N_A_1291_93#_c_804_n A_1735_119# 0.00707295f $X=8.83 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_721 N_A_1163_119#_M1003_g N_SET_B_M1030_g 0.0144806f $X=7.25 $Y=2.525 $X2=0
+ $Y2=0
cc_722 N_A_1163_119#_M1013_g N_SET_B_M1030_g 0.0119468f $X=8.41 $Y=2.315 $X2=0
+ $Y2=0
cc_723 N_A_1163_119#_M1003_g N_SET_B_M1024_g 0.00839305f $X=7.25 $Y=2.525 $X2=0
+ $Y2=0
cc_724 N_A_1163_119#_c_914_n N_SET_B_M1024_g 0.051977f $X=7.575 $Y=1.125 $X2=0
+ $Y2=0
cc_725 N_A_1163_119#_M1013_g N_SET_B_M1024_g 0.0174681f $X=8.41 $Y=2.315 $X2=0
+ $Y2=0
cc_726 N_A_1163_119#_c_915_n N_SET_B_M1024_g 0.0178805f $X=8.6 $Y=1.345 $X2=0
+ $Y2=0
cc_727 N_A_1163_119#_c_917_n N_SET_B_M1024_g 0.0113302f $X=8.385 $Y=1.29 $X2=0
+ $Y2=0
cc_728 N_A_1163_119#_c_927_n N_SET_B_M1024_g 9.15467e-19 $X=8.48 $Y=1.51 $X2=0
+ $Y2=0
cc_729 N_A_1163_119#_c_918_n N_SET_B_M1024_g 0.0136954f $X=8.48 $Y=1.51 $X2=0
+ $Y2=0
cc_730 N_A_1163_119#_c_921_n N_SET_B_M1024_g 0.00679914f $X=7.34 $Y=1.29 $X2=0
+ $Y2=0
cc_731 N_A_1163_119#_c_923_n N_SET_B_M1024_g 3.05142e-19 $X=7.505 $Y=1.257 $X2=0
+ $Y2=0
cc_732 N_A_1163_119#_M1013_g N_SET_B_c_1055_n 0.00243139f $X=8.41 $Y=2.315 $X2=0
+ $Y2=0
cc_733 N_A_1163_119#_c_917_n N_SET_B_c_1055_n 0.00171411f $X=8.385 $Y=1.29 $X2=0
+ $Y2=0
cc_734 N_A_1163_119#_c_927_n N_SET_B_c_1055_n 0.00112058f $X=8.48 $Y=1.51 $X2=0
+ $Y2=0
cc_735 N_A_1163_119#_M1003_g N_SET_B_c_1056_n 5.88375e-19 $X=7.25 $Y=2.525 $X2=0
+ $Y2=0
cc_736 N_A_1163_119#_M1003_g N_SET_B_c_1059_n 0.00718947f $X=7.25 $Y=2.525 $X2=0
+ $Y2=0
cc_737 N_A_1163_119#_M1013_g N_SET_B_c_1059_n 6.97942e-19 $X=8.41 $Y=2.315 $X2=0
+ $Y2=0
cc_738 N_A_1163_119#_M1003_g N_SET_B_c_1060_n 0.0220402f $X=7.25 $Y=2.525 $X2=0
+ $Y2=0
cc_739 N_A_1163_119#_c_921_n N_SET_B_c_1060_n 0.00178572f $X=7.34 $Y=1.29 $X2=0
+ $Y2=0
cc_740 N_A_1163_119#_c_926_n N_A_629_47#_c_1185_n 0.00324268f $X=6.085 $Y=2.525
+ $X2=0 $Y2=0
cc_741 N_A_1163_119#_c_916_n N_A_629_47#_M1039_g 0.00107485f $X=5.955 $Y=0.805
+ $X2=0 $Y2=0
cc_742 N_A_1163_119#_c_914_n N_A_629_47#_c_1176_n 0.00979198f $X=7.575 $Y=1.125
+ $X2=0 $Y2=0
cc_743 N_A_1163_119#_c_915_n N_A_629_47#_c_1176_n 0.0100759f $X=8.6 $Y=1.345
+ $X2=0 $Y2=0
cc_744 N_A_1163_119#_c_916_n N_A_629_47#_c_1176_n 0.00339559f $X=5.955 $Y=0.805
+ $X2=0 $Y2=0
cc_745 N_A_1163_119#_c_926_n N_A_629_47#_M1026_g 0.00975559f $X=6.085 $Y=2.525
+ $X2=0 $Y2=0
cc_746 N_A_1163_119#_c_930_n N_A_629_47#_M1026_g 3.38663e-19 $X=6.037 $Y=2.19
+ $X2=0 $Y2=0
cc_747 N_A_1163_119#_M1003_g N_A_629_47#_c_1188_n 0.0100244f $X=7.25 $Y=2.525
+ $X2=0 $Y2=0
cc_748 N_A_1163_119#_M1013_g N_A_629_47#_c_1188_n 0.0104164f $X=8.41 $Y=2.315
+ $X2=0 $Y2=0
cc_749 N_A_1163_119#_M1013_g N_A_629_47#_M1031_g 0.0330879f $X=8.41 $Y=2.315
+ $X2=0 $Y2=0
cc_750 N_A_1163_119#_M1013_g N_A_1799_408#_c_1414_n 0.00144167f $X=8.41 $Y=2.315
+ $X2=0 $Y2=0
cc_751 N_A_1163_119#_M1003_g N_VPWR_c_1630_n 0.00434527f $X=7.25 $Y=2.525 $X2=0
+ $Y2=0
cc_752 N_A_1163_119#_M1013_g N_VPWR_c_1631_n 0.00468574f $X=8.41 $Y=2.315 $X2=0
+ $Y2=0
cc_753 N_A_1163_119#_c_926_n N_VPWR_c_1650_n 0.00462306f $X=6.085 $Y=2.525 $X2=0
+ $Y2=0
cc_754 N_A_1163_119#_M1003_g N_VPWR_c_1627_n 9.39239e-19 $X=7.25 $Y=2.525 $X2=0
+ $Y2=0
cc_755 N_A_1163_119#_M1013_g N_VPWR_c_1627_n 9.39239e-19 $X=8.41 $Y=2.315 $X2=0
+ $Y2=0
cc_756 N_A_1163_119#_c_926_n N_VPWR_c_1627_n 0.00777186f $X=6.085 $Y=2.525 $X2=0
+ $Y2=0
cc_757 N_A_1163_119#_c_916_n N_A_268_467#_c_1803_n 0.0100624f $X=5.955 $Y=0.805
+ $X2=0 $Y2=0
cc_758 N_A_1163_119#_c_926_n N_A_268_467#_c_1804_n 0.00713098f $X=6.085 $Y=2.525
+ $X2=0 $Y2=0
cc_759 N_A_1163_119#_c_920_n N_A_268_467#_c_1804_n 0.063059f $X=6.037 $Y=2.02
+ $X2=0 $Y2=0
cc_760 N_A_1163_119#_c_919_n N_A_268_467#_c_1805_n 0.0176253f $X=5.972 $Y=1.242
+ $X2=0 $Y2=0
cc_761 N_A_1163_119#_c_917_n N_VGND_M1024_d 0.00328644f $X=8.385 $Y=1.29 $X2=0
+ $Y2=0
cc_762 N_A_1163_119#_c_914_n N_VGND_c_1985_n 0.00388132f $X=7.575 $Y=1.125 $X2=0
+ $Y2=0
cc_763 N_A_1163_119#_c_916_n N_VGND_c_1985_n 0.0109469f $X=5.955 $Y=0.805 $X2=0
+ $Y2=0
cc_764 N_A_1163_119#_c_922_n N_VGND_c_1985_n 0.0239807f $X=7.175 $Y=1.257 $X2=0
+ $Y2=0
cc_765 N_A_1163_119#_c_915_n N_VGND_c_1986_n 0.00452992f $X=8.6 $Y=1.345 $X2=0
+ $Y2=0
cc_766 N_A_1163_119#_c_916_n N_VGND_c_2000_n 0.00458155f $X=5.955 $Y=0.805 $X2=0
+ $Y2=0
cc_767 N_A_1163_119#_c_914_n N_VGND_c_2012_n 9.39239e-19 $X=7.575 $Y=1.125 $X2=0
+ $Y2=0
cc_768 N_A_1163_119#_c_915_n N_VGND_c_2012_n 9.39239e-19 $X=8.6 $Y=1.345 $X2=0
+ $Y2=0
cc_769 N_A_1163_119#_c_916_n N_VGND_c_2012_n 0.00767083f $X=5.955 $Y=0.805 $X2=0
+ $Y2=0
cc_770 N_SET_B_M1024_g N_A_629_47#_c_1176_n 0.00988663f $X=7.935 $Y=0.805 $X2=0
+ $Y2=0
cc_771 N_SET_B_M1030_g N_A_629_47#_c_1188_n 0.0100244f $X=7.68 $Y=2.525 $X2=0
+ $Y2=0
cc_772 N_SET_B_c_1055_n N_A_629_47#_M1031_g 0.00251975f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_773 N_SET_B_c_1053_n N_A_1946_369#_M1002_g 0.0174351f $X=10.47 $Y=2.225 $X2=0
+ $Y2=0
cc_774 N_SET_B_c_1055_n N_A_1946_369#_M1002_g 0.00212443f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_SET_B_c_1043_n N_A_1946_369#_M1038_g 0.0477771f $X=10.29 $Y=1.125 $X2=0
+ $Y2=0
cc_776 N_SET_B_c_1046_n N_A_1946_369#_M1038_g 0.0015531f $X=10.8 $Y=1.63 $X2=0
+ $Y2=0
cc_777 N_SET_B_c_1045_n N_A_1946_369#_c_1303_n 0.00255064f $X=10.365 $Y=1.2
+ $X2=0 $Y2=0
cc_778 N_SET_B_c_1046_n N_A_1946_369#_c_1303_n 0.00504687f $X=10.8 $Y=1.63 $X2=0
+ $Y2=0
cc_779 N_SET_B_c_1055_n N_A_1946_369#_c_1303_n 0.00977948f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_780 N_SET_B_c_1048_n N_A_1946_369#_c_1303_n 0.00845622f $X=10.8 $Y=1.795
+ $X2=0 $Y2=0
cc_781 N_SET_B_c_1043_n N_A_1946_369#_c_1304_n 0.0012427f $X=10.29 $Y=1.125
+ $X2=0 $Y2=0
cc_782 N_SET_B_c_1044_n N_A_1946_369#_c_1304_n 0.0285112f $X=10.635 $Y=1.2 $X2=0
+ $Y2=0
cc_783 N_SET_B_c_1045_n N_A_1946_369#_c_1304_n 9.28404e-19 $X=10.365 $Y=1.2
+ $X2=0 $Y2=0
cc_784 N_SET_B_c_1047_n N_A_1946_369#_c_1304_n 0.00298905f $X=10.8 $Y=1.795
+ $X2=0 $Y2=0
cc_785 N_SET_B_c_1048_n N_A_1946_369#_c_1304_n 0.00797154f $X=10.8 $Y=1.795
+ $X2=0 $Y2=0
cc_786 N_SET_B_c_1043_n N_A_1946_369#_c_1305_n 0.00700072f $X=10.29 $Y=1.125
+ $X2=0 $Y2=0
cc_787 N_SET_B_c_1045_n N_A_1946_369#_c_1305_n 0.00247347f $X=10.365 $Y=1.2
+ $X2=0 $Y2=0
cc_788 N_SET_B_c_1045_n N_A_1946_369#_c_1310_n 0.007194f $X=10.365 $Y=1.2 $X2=0
+ $Y2=0
cc_789 N_SET_B_c_1053_n N_A_1946_369#_c_1310_n 0.00105822f $X=10.47 $Y=2.225
+ $X2=0 $Y2=0
cc_790 N_SET_B_c_1046_n N_A_1946_369#_c_1310_n 0.0147029f $X=10.8 $Y=1.63 $X2=0
+ $Y2=0
cc_791 N_SET_B_c_1054_n N_A_1946_369#_c_1310_n 0.00375368f $X=10.8 $Y=2.15 $X2=0
+ $Y2=0
cc_792 N_SET_B_c_1055_n N_A_1946_369#_c_1310_n 0.00887519f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_793 N_SET_B_c_1048_n N_A_1946_369#_c_1310_n 8.18306e-19 $X=10.8 $Y=1.795
+ $X2=0 $Y2=0
cc_794 N_SET_B_c_1055_n N_A_1799_408#_M1031_d 0.00196494f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_795 N_SET_B_c_1044_n N_A_1799_408#_M1028_g 0.00394105f $X=10.635 $Y=1.2 $X2=0
+ $Y2=0
cc_796 N_SET_B_c_1047_n N_A_1799_408#_M1010_g 0.00473869f $X=10.8 $Y=1.795 $X2=0
+ $Y2=0
cc_797 N_SET_B_c_1055_n N_A_1799_408#_c_1414_n 0.00789257f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_SET_B_c_1055_n N_A_1799_408#_c_1406_n 0.0257785f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_799 N_SET_B_M1000_g N_A_1799_408#_c_1416_n 6.01315e-19 $X=10.395 $Y=2.67
+ $X2=0 $Y2=0
cc_800 N_SET_B_M1000_g N_A_1799_408#_c_1417_n 0.00343401f $X=10.395 $Y=2.67
+ $X2=0 $Y2=0
cc_801 N_SET_B_c_1052_n N_A_1799_408#_c_1417_n 0.00533095f $X=10.635 $Y=2.225
+ $X2=0 $Y2=0
cc_802 N_SET_B_c_1053_n N_A_1799_408#_c_1417_n 0.0063074f $X=10.47 $Y=2.225
+ $X2=0 $Y2=0
cc_803 N_SET_B_c_1055_n N_A_1799_408#_c_1417_n 0.0297298f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_804 N_SET_B_c_1048_n N_A_1799_408#_c_1417_n 0.0111307f $X=10.8 $Y=1.795 $X2=0
+ $Y2=0
cc_805 N_SET_B_M1000_g N_A_1799_408#_c_1418_n 0.00608752f $X=10.395 $Y=2.67
+ $X2=0 $Y2=0
cc_806 N_SET_B_c_1052_n N_A_1799_408#_c_1419_n 0.0109098f $X=10.635 $Y=2.225
+ $X2=0 $Y2=0
cc_807 N_SET_B_c_1055_n N_A_1799_408#_c_1419_n 0.00456025f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_808 SET_B N_A_1799_408#_c_1419_n 0.00501838f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_809 N_SET_B_c_1048_n N_A_1799_408#_c_1419_n 0.0124755f $X=10.8 $Y=1.795 $X2=0
+ $Y2=0
cc_810 N_SET_B_M1000_g N_A_1799_408#_c_1456_n 0.00670927f $X=10.395 $Y=2.67
+ $X2=0 $Y2=0
cc_811 N_SET_B_M1000_g N_A_1799_408#_c_1420_n 9.35868e-19 $X=10.395 $Y=2.67
+ $X2=0 $Y2=0
cc_812 SET_B N_A_1799_408#_c_1420_n 0.00669814f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_813 N_SET_B_c_1047_n N_A_1799_408#_c_1420_n 0.00809747f $X=10.8 $Y=1.795
+ $X2=0 $Y2=0
cc_814 N_SET_B_c_1048_n N_A_1799_408#_c_1420_n 0.044913f $X=10.8 $Y=1.795 $X2=0
+ $Y2=0
cc_815 N_SET_B_c_1046_n N_A_1799_408#_c_1407_n 0.00493213f $X=10.8 $Y=1.63 $X2=0
+ $Y2=0
cc_816 N_SET_B_c_1048_n N_A_1799_408#_c_1407_n 0.00119132f $X=10.8 $Y=1.795
+ $X2=0 $Y2=0
cc_817 N_SET_B_c_1046_n N_A_1799_408#_c_1409_n 0.00721088f $X=10.8 $Y=1.63 $X2=0
+ $Y2=0
cc_818 N_SET_B_c_1047_n N_A_1799_408#_c_1409_n 0.00187231f $X=10.8 $Y=1.795
+ $X2=0 $Y2=0
cc_819 N_SET_B_c_1055_n N_VPWR_M1030_d 0.00184562f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_820 N_SET_B_M1030_g N_VPWR_c_1631_n 0.00500072f $X=7.68 $Y=2.525 $X2=0 $Y2=0
cc_821 N_SET_B_c_1055_n N_VPWR_c_1631_n 7.53696e-19 $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_822 N_SET_B_M1000_g N_VPWR_c_1632_n 0.006799f $X=10.395 $Y=2.67 $X2=0 $Y2=0
cc_823 N_SET_B_M1000_g N_VPWR_c_1644_n 0.00426287f $X=10.395 $Y=2.67 $X2=0 $Y2=0
cc_824 N_SET_B_M1030_g N_VPWR_c_1627_n 9.39239e-19 $X=7.68 $Y=2.525 $X2=0 $Y2=0
cc_825 N_SET_B_M1000_g N_VPWR_c_1627_n 0.00520574f $X=10.395 $Y=2.67 $X2=0 $Y2=0
cc_826 N_SET_B_c_1055_n A_1697_379# 0.00266935f $X=10.655 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_827 N_SET_B_M1024_g N_VGND_c_1986_n 0.00526528f $X=7.935 $Y=0.805 $X2=0 $Y2=0
cc_828 N_SET_B_c_1043_n N_VGND_c_1987_n 0.0109909f $X=10.29 $Y=1.125 $X2=0 $Y2=0
cc_829 N_SET_B_c_1044_n N_VGND_c_1987_n 0.00201433f $X=10.635 $Y=1.2 $X2=0 $Y2=0
cc_830 N_SET_B_c_1043_n N_VGND_c_2002_n 0.0035863f $X=10.29 $Y=1.125 $X2=0 $Y2=0
cc_831 N_SET_B_M1024_g N_VGND_c_2012_n 9.39239e-19 $X=7.935 $Y=0.805 $X2=0 $Y2=0
cc_832 N_SET_B_c_1043_n N_VGND_c_2012_n 0.00401353f $X=10.29 $Y=1.125 $X2=0
+ $Y2=0
cc_833 N_A_629_47#_M1032_g N_A_1946_369#_M1038_g 0.0384845f $X=9.57 $Y=0.805
+ $X2=0 $Y2=0
cc_834 N_A_629_47#_M1031_g N_A_1799_408#_c_1414_n 0.00815929f $X=8.92 $Y=2.46
+ $X2=0 $Y2=0
cc_835 N_A_629_47#_c_1176_n N_A_1799_408#_c_1405_n 0.00509664f $X=9.495 $Y=0.18
+ $X2=0 $Y2=0
cc_836 N_A_629_47#_M1032_g N_A_1799_408#_c_1405_n 0.0144847f $X=9.57 $Y=0.805
+ $X2=0 $Y2=0
cc_837 N_A_629_47#_M1032_g N_A_1799_408#_c_1406_n 0.00164539f $X=9.57 $Y=0.805
+ $X2=0 $Y2=0
cc_838 N_A_629_47#_M1006_g N_VPWR_c_1629_n 0.0218258f $X=4.525 $Y=2.265 $X2=0
+ $Y2=0
cc_839 N_A_629_47#_M1026_g N_VPWR_c_1630_n 0.00636556f $X=6.3 $Y=2.525 $X2=0
+ $Y2=0
cc_840 N_A_629_47#_c_1188_n N_VPWR_c_1630_n 0.0254367f $X=8.845 $Y=3.15 $X2=0
+ $Y2=0
cc_841 N_A_629_47#_c_1188_n N_VPWR_c_1631_n 0.0254148f $X=8.845 $Y=3.15 $X2=0
+ $Y2=0
cc_842 N_A_629_47#_M1031_g N_VPWR_c_1631_n 0.00561647f $X=8.92 $Y=2.46 $X2=0
+ $Y2=0
cc_843 N_A_629_47#_c_1188_n N_VPWR_c_1640_n 0.0257522f $X=8.845 $Y=3.15 $X2=0
+ $Y2=0
cc_844 N_A_629_47#_c_1188_n N_VPWR_c_1642_n 0.0257758f $X=8.845 $Y=3.15 $X2=0
+ $Y2=0
cc_845 N_A_629_47#_c_1186_n N_VPWR_c_1650_n 0.0781767f $X=4.6 $Y=3.15 $X2=0
+ $Y2=0
cc_846 N_A_629_47#_c_1185_n N_VPWR_c_1627_n 0.0475104f $X=6.225 $Y=3.15 $X2=0
+ $Y2=0
cc_847 N_A_629_47#_c_1186_n N_VPWR_c_1627_n 0.00709472f $X=4.6 $Y=3.15 $X2=0
+ $Y2=0
cc_848 N_A_629_47#_c_1188_n N_VPWR_c_1627_n 0.079907f $X=8.845 $Y=3.15 $X2=0
+ $Y2=0
cc_849 N_A_629_47#_c_1190_n N_VPWR_c_1627_n 0.00847591f $X=6.3 $Y=3.15 $X2=0
+ $Y2=0
cc_850 N_A_629_47#_c_1182_n N_A_268_467#_c_1800_n 0.0152015f $X=3.745 $Y=1.23
+ $X2=0 $Y2=0
cc_851 N_A_629_47#_c_1180_n N_A_268_467#_c_1802_n 0.0656163f $X=3.495 $Y=2.46
+ $X2=0 $Y2=0
cc_852 N_A_629_47#_c_1182_n N_A_268_467#_c_1802_n 0.0161001f $X=3.745 $Y=1.23
+ $X2=0 $Y2=0
cc_853 N_A_629_47#_M1025_d N_A_268_467#_c_1808_n 0.00484253f $X=3.355 $Y=2.335
+ $X2=0 $Y2=0
cc_854 N_A_629_47#_c_1180_n N_A_268_467#_c_1808_n 0.0138446f $X=3.495 $Y=2.46
+ $X2=0 $Y2=0
cc_855 N_A_629_47#_M1006_g N_A_268_467#_c_1809_n 0.00417195f $X=4.525 $Y=2.265
+ $X2=0 $Y2=0
cc_856 N_A_629_47#_c_1180_n N_A_268_467#_c_1809_n 0.00965725f $X=3.495 $Y=2.46
+ $X2=0 $Y2=0
cc_857 N_A_629_47#_M1006_g N_A_268_467#_c_1810_n 0.0198448f $X=4.525 $Y=2.265
+ $X2=0 $Y2=0
cc_858 N_A_629_47#_c_1185_n N_A_268_467#_c_1810_n 0.0177093f $X=6.225 $Y=3.15
+ $X2=0 $Y2=0
cc_859 N_A_629_47#_c_1180_n N_A_268_467#_c_1811_n 0.0142359f $X=3.495 $Y=2.46
+ $X2=0 $Y2=0
cc_860 N_A_629_47#_c_1173_n N_A_268_467#_c_1803_n 0.00410445f $X=5.665 $Y=0.18
+ $X2=0 $Y2=0
cc_861 N_A_629_47#_M1039_g N_A_268_467#_c_1803_n 0.00336364f $X=5.74 $Y=0.805
+ $X2=0 $Y2=0
cc_862 N_A_629_47#_c_1185_n N_A_268_467#_c_1813_n 0.00563294f $X=6.225 $Y=3.15
+ $X2=0 $Y2=0
cc_863 N_A_629_47#_c_1174_n N_VGND_c_1984_n 0.0110948f $X=4.6 $Y=0.18 $X2=0
+ $Y2=0
cc_864 N_A_629_47#_c_1179_n N_VGND_c_1984_n 0.0251521f $X=3.55 $Y=0.44 $X2=0
+ $Y2=0
cc_865 N_A_629_47#_c_1181_n N_VGND_c_1984_n 0.00868213f $X=3.745 $Y=0.895 $X2=0
+ $Y2=0
cc_866 N_A_629_47#_c_1182_n N_VGND_c_1984_n 0.0220981f $X=3.745 $Y=1.23 $X2=0
+ $Y2=0
cc_867 N_A_629_47#_c_1183_n N_VGND_c_1984_n 0.00198652f $X=4.24 $Y=1.06 $X2=0
+ $Y2=0
cc_868 N_A_629_47#_c_1176_n N_VGND_c_1985_n 0.0257254f $X=9.495 $Y=0.18 $X2=0
+ $Y2=0
cc_869 N_A_629_47#_c_1176_n N_VGND_c_1986_n 0.0254542f $X=9.495 $Y=0.18 $X2=0
+ $Y2=0
cc_870 N_A_629_47#_c_1176_n N_VGND_c_1987_n 0.00651874f $X=9.495 $Y=0.18 $X2=0
+ $Y2=0
cc_871 N_A_629_47#_c_1179_n N_VGND_c_1998_n 0.0457994f $X=3.55 $Y=0.44 $X2=0
+ $Y2=0
cc_872 N_A_629_47#_c_1174_n N_VGND_c_2000_n 0.0666735f $X=4.6 $Y=0.18 $X2=0
+ $Y2=0
cc_873 N_A_629_47#_c_1176_n N_VGND_c_2002_n 0.0366508f $X=9.495 $Y=0.18 $X2=0
+ $Y2=0
cc_874 N_A_629_47#_c_1176_n N_VGND_c_2004_n 0.0358829f $X=9.495 $Y=0.18 $X2=0
+ $Y2=0
cc_875 N_A_629_47#_M1023_d N_VGND_c_2012_n 0.00240648f $X=3.145 $Y=0.235 $X2=0
+ $Y2=0
cc_876 N_A_629_47#_c_1173_n N_VGND_c_2012_n 0.0409824f $X=5.665 $Y=0.18 $X2=0
+ $Y2=0
cc_877 N_A_629_47#_c_1174_n N_VGND_c_2012_n 0.0105884f $X=4.6 $Y=0.18 $X2=0
+ $Y2=0
cc_878 N_A_629_47#_c_1176_n N_VGND_c_2012_n 0.115442f $X=9.495 $Y=0.18 $X2=0
+ $Y2=0
cc_879 N_A_629_47#_c_1178_n N_VGND_c_2012_n 0.00926736f $X=5.74 $Y=0.18 $X2=0
+ $Y2=0
cc_880 N_A_629_47#_c_1179_n N_VGND_c_2012_n 0.0285977f $X=3.55 $Y=0.44 $X2=0
+ $Y2=0
cc_881 N_A_1946_369#_c_1307_n N_A_1799_408#_M1028_g 0.0159779f $X=11.755 $Y=1.17
+ $X2=0 $Y2=0
cc_882 N_A_1946_369#_c_1308_n N_A_1799_408#_M1028_g 0.00195831f $X=11.84
+ $Y=1.815 $X2=0 $Y2=0
cc_883 N_A_1946_369#_c_1313_n N_A_1799_408#_M1010_g 0.0169673f $X=11.755 $Y=1.98
+ $X2=0 $Y2=0
cc_884 N_A_1946_369#_c_1308_n N_A_1799_408#_M1010_g 0.00401423f $X=11.84
+ $Y=1.815 $X2=0 $Y2=0
cc_885 N_A_1946_369#_c_1308_n N_A_1799_408#_c_1395_n 0.00791517f $X=11.84
+ $Y=1.815 $X2=0 $Y2=0
cc_886 N_A_1946_369#_c_1307_n N_A_1799_408#_M1018_g 0.00178606f $X=11.755
+ $Y=1.17 $X2=0 $Y2=0
cc_887 N_A_1946_369#_c_1308_n N_A_1799_408#_M1018_g 8.1579e-19 $X=11.84 $Y=1.815
+ $X2=0 $Y2=0
cc_888 N_A_1946_369#_c_1313_n N_A_1799_408#_M1022_g 0.0015048f $X=11.755 $Y=1.98
+ $X2=0 $Y2=0
cc_889 N_A_1946_369#_c_1308_n N_A_1799_408#_M1022_g 0.00111759f $X=11.84
+ $Y=1.815 $X2=0 $Y2=0
cc_890 N_A_1946_369#_M1002_g N_A_1799_408#_c_1414_n 0.00942094f $X=9.805 $Y=2.67
+ $X2=0 $Y2=0
cc_891 N_A_1946_369#_M1038_g N_A_1799_408#_c_1405_n 9.90202e-19 $X=9.93 $Y=0.805
+ $X2=0 $Y2=0
cc_892 N_A_1946_369#_M1002_g N_A_1799_408#_c_1406_n 0.00565709f $X=9.805 $Y=2.67
+ $X2=0 $Y2=0
cc_893 N_A_1946_369#_M1038_g N_A_1799_408#_c_1406_n 0.0130104f $X=9.93 $Y=0.805
+ $X2=0 $Y2=0
cc_894 N_A_1946_369#_c_1303_n N_A_1799_408#_c_1406_n 0.0434954f $X=10.18 $Y=1.68
+ $X2=0 $Y2=0
cc_895 N_A_1946_369#_c_1305_n N_A_1799_408#_c_1406_n 0.0137764f $X=10.345
+ $Y=1.17 $X2=0 $Y2=0
cc_896 N_A_1946_369#_c_1310_n N_A_1799_408#_c_1406_n 0.00981139f $X=9.93
+ $Y=1.755 $X2=0 $Y2=0
cc_897 N_A_1946_369#_M1002_g N_A_1799_408#_c_1416_n 0.00545993f $X=9.805 $Y=2.67
+ $X2=0 $Y2=0
cc_898 N_A_1946_369#_M1002_g N_A_1799_408#_c_1417_n 0.00614731f $X=9.805 $Y=2.67
+ $X2=0 $Y2=0
cc_899 N_A_1946_369#_c_1303_n N_A_1799_408#_c_1417_n 0.00955454f $X=10.18
+ $Y=1.68 $X2=0 $Y2=0
cc_900 N_A_1946_369#_c_1310_n N_A_1799_408#_c_1417_n 0.00658326f $X=9.93
+ $Y=1.755 $X2=0 $Y2=0
cc_901 N_A_1946_369#_M1002_g N_A_1799_408#_c_1418_n 5.89204e-19 $X=9.805 $Y=2.67
+ $X2=0 $Y2=0
cc_902 N_A_1946_369#_c_1313_n N_A_1799_408#_c_1420_n 0.0246275f $X=11.755
+ $Y=1.98 $X2=0 $Y2=0
cc_903 N_A_1946_369#_c_1308_n N_A_1799_408#_c_1420_n 0.00520515f $X=11.84
+ $Y=1.815 $X2=0 $Y2=0
cc_904 N_A_1946_369#_c_1304_n N_A_1799_408#_c_1407_n 0.00460752f $X=11.12
+ $Y=1.17 $X2=0 $Y2=0
cc_905 N_A_1946_369#_c_1309_n N_A_1799_408#_c_1407_n 0.0106004f $X=11.25 $Y=1.17
+ $X2=0 $Y2=0
cc_906 N_A_1946_369#_c_1307_n N_A_1799_408#_c_1408_n 0.0136149f $X=11.755
+ $Y=1.17 $X2=0 $Y2=0
cc_907 N_A_1946_369#_c_1313_n N_A_1799_408#_c_1408_n 0.0122999f $X=11.755
+ $Y=1.98 $X2=0 $Y2=0
cc_908 N_A_1946_369#_c_1308_n N_A_1799_408#_c_1408_n 0.0154823f $X=11.84
+ $Y=1.815 $X2=0 $Y2=0
cc_909 N_A_1946_369#_c_1309_n N_A_1799_408#_c_1408_n 0.0116776f $X=11.25 $Y=1.17
+ $X2=0 $Y2=0
cc_910 N_A_1946_369#_M1002_g N_A_1799_408#_c_1421_n 0.00237435f $X=9.805 $Y=2.67
+ $X2=0 $Y2=0
cc_911 N_A_1946_369#_c_1307_n N_A_1799_408#_c_1409_n 0.00412051f $X=11.755
+ $Y=1.17 $X2=0 $Y2=0
cc_912 N_A_1946_369#_c_1313_n N_A_1799_408#_c_1409_n 0.00650677f $X=11.755
+ $Y=1.98 $X2=0 $Y2=0
cc_913 N_A_1946_369#_c_1308_n N_A_1799_408#_c_1409_n 0.0104928f $X=11.84
+ $Y=1.815 $X2=0 $Y2=0
cc_914 N_A_1946_369#_c_1309_n N_A_1799_408#_c_1409_n 0.00343667f $X=11.25
+ $Y=1.17 $X2=0 $Y2=0
cc_915 N_A_1946_369#_c_1313_n N_VPWR_M1010_d 0.00448227f $X=11.755 $Y=1.98 $X2=0
+ $Y2=0
cc_916 N_A_1946_369#_M1002_g N_VPWR_c_1632_n 0.00598823f $X=9.805 $Y=2.67 $X2=0
+ $Y2=0
cc_917 N_A_1946_369#_c_1313_n N_VPWR_c_1633_n 0.0058393f $X=11.755 $Y=1.98 $X2=0
+ $Y2=0
cc_918 N_A_1946_369#_M1002_g N_VPWR_c_1642_n 0.00422736f $X=9.805 $Y=2.67 $X2=0
+ $Y2=0
cc_919 N_A_1946_369#_M1002_g N_VPWR_c_1627_n 0.00520574f $X=9.805 $Y=2.67 $X2=0
+ $Y2=0
cc_920 N_A_1946_369#_c_1307_n N_Q_N_c_1930_n 0.0113727f $X=11.755 $Y=1.17 $X2=0
+ $Y2=0
cc_921 N_A_1946_369#_c_1308_n N_Q_N_c_1930_n 0.0340037f $X=11.84 $Y=1.815 $X2=0
+ $Y2=0
cc_922 N_A_1946_369#_c_1313_n N_Q_N_c_1935_n 0.00109262f $X=11.755 $Y=1.98 $X2=0
+ $Y2=0
cc_923 N_A_1946_369#_c_1313_n N_Q_N_c_1932_n 0.0111851f $X=11.755 $Y=1.98 $X2=0
+ $Y2=0
cc_924 N_A_1946_369#_c_1307_n N_VGND_M1028_d 0.00188126f $X=11.755 $Y=1.17 $X2=0
+ $Y2=0
cc_925 N_A_1946_369#_M1038_g N_VGND_c_1987_n 0.00153352f $X=9.93 $Y=0.805 $X2=0
+ $Y2=0
cc_926 N_A_1946_369#_c_1304_n N_VGND_c_1987_n 0.0240949f $X=11.12 $Y=1.17 $X2=0
+ $Y2=0
cc_927 N_A_1946_369#_c_1306_n N_VGND_c_1987_n 0.00855781f $X=11.285 $Y=0.875
+ $X2=0 $Y2=0
cc_928 N_A_1946_369#_c_1307_n N_VGND_c_1988_n 0.0294016f $X=11.755 $Y=1.17 $X2=0
+ $Y2=0
cc_929 N_A_1946_369#_M1038_g N_VGND_c_2002_n 0.00431487f $X=9.93 $Y=0.805 $X2=0
+ $Y2=0
cc_930 N_A_1946_369#_c_1306_n N_VGND_c_2005_n 0.00413385f $X=11.285 $Y=0.875
+ $X2=0 $Y2=0
cc_931 N_A_1946_369#_M1038_g N_VGND_c_2012_n 0.00477801f $X=9.93 $Y=0.805 $X2=0
+ $Y2=0
cc_932 N_A_1946_369#_c_1306_n N_VGND_c_2012_n 0.00732771f $X=11.285 $Y=0.875
+ $X2=0 $Y2=0
cc_933 N_A_1799_408#_M1042_g N_A_2624_49#_c_1573_n 0.0159719f $X=13.045 $Y=0.455
+ $X2=0 $Y2=0
cc_934 N_A_1799_408#_M1040_g N_A_2624_49#_c_1574_n 0.00109001f $X=12.67 $Y=2.465
+ $X2=0 $Y2=0
cc_935 N_A_1799_408#_M1009_g N_A_2624_49#_c_1574_n 0.014823f $X=13.195 $Y=2.155
+ $X2=0 $Y2=0
cc_936 N_A_1799_408#_M1040_g N_A_2624_49#_c_1577_n 4.88052e-19 $X=12.67 $Y=2.465
+ $X2=0 $Y2=0
cc_937 N_A_1799_408#_M1042_g N_A_2624_49#_c_1577_n 0.00219723f $X=13.045
+ $Y=0.455 $X2=0 $Y2=0
cc_938 N_A_1799_408#_M1009_g N_A_2624_49#_c_1577_n 0.00396269f $X=13.195
+ $Y=2.155 $X2=0 $Y2=0
cc_939 N_A_1799_408#_c_1404_n N_A_2624_49#_c_1577_n 0.0105059f $X=13.195 $Y=1.42
+ $X2=0 $Y2=0
cc_940 N_A_1799_408#_M1042_g N_A_2624_49#_c_1578_n 8.82307e-19 $X=13.045
+ $Y=0.455 $X2=0 $Y2=0
cc_941 N_A_1799_408#_c_1404_n N_A_2624_49#_c_1578_n 0.00616394f $X=13.195
+ $Y=1.42 $X2=0 $Y2=0
cc_942 N_A_1799_408#_c_1414_n N_VPWR_c_1632_n 0.0261401f $X=9.665 $Y=2.72 $X2=0
+ $Y2=0
cc_943 N_A_1799_408#_c_1416_n N_VPWR_c_1632_n 0.00350689f $X=9.75 $Y=2.555 $X2=0
+ $Y2=0
cc_944 N_A_1799_408#_c_1417_n N_VPWR_c_1632_n 0.0147698f $X=10.365 $Y=2.245
+ $X2=0 $Y2=0
cc_945 N_A_1799_408#_c_1456_n N_VPWR_c_1632_n 0.0261401f $X=10.535 $Y=2.67 $X2=0
+ $Y2=0
cc_946 N_A_1799_408#_M1010_g N_VPWR_c_1633_n 9.96206e-19 $X=11.715 $Y=2.045
+ $X2=0 $Y2=0
cc_947 N_A_1799_408#_M1022_g N_VPWR_c_1633_n 0.00477819f $X=12.24 $Y=2.465 $X2=0
+ $Y2=0
cc_948 N_A_1799_408#_c_1419_n N_VPWR_c_1633_n 0.0115586f $X=11.065 $Y=2.67 $X2=0
+ $Y2=0
cc_949 N_A_1799_408#_c_1420_n N_VPWR_c_1633_n 0.00593128f $X=11.15 $Y=2.505
+ $X2=0 $Y2=0
cc_950 N_A_1799_408#_M1040_g N_VPWR_c_1634_n 0.00645359f $X=12.67 $Y=2.465 $X2=0
+ $Y2=0
cc_951 N_A_1799_408#_c_1400_n N_VPWR_c_1634_n 0.00774041f $X=12.97 $Y=1.42 $X2=0
+ $Y2=0
cc_952 N_A_1799_408#_M1009_g N_VPWR_c_1634_n 0.00534442f $X=13.195 $Y=2.155
+ $X2=0 $Y2=0
cc_953 N_A_1799_408#_c_1414_n N_VPWR_c_1642_n 0.0259479f $X=9.665 $Y=2.72 $X2=0
+ $Y2=0
cc_954 N_A_1799_408#_c_1419_n N_VPWR_c_1644_n 0.018576f $X=11.065 $Y=2.67 $X2=0
+ $Y2=0
cc_955 N_A_1799_408#_c_1456_n N_VPWR_c_1644_n 0.00368997f $X=10.535 $Y=2.67
+ $X2=0 $Y2=0
cc_956 N_A_1799_408#_M1022_g N_VPWR_c_1646_n 0.0054895f $X=12.24 $Y=2.465 $X2=0
+ $Y2=0
cc_957 N_A_1799_408#_M1040_g N_VPWR_c_1646_n 0.00585385f $X=12.67 $Y=2.465 $X2=0
+ $Y2=0
cc_958 N_A_1799_408#_M1009_g N_VPWR_c_1651_n 0.00312414f $X=13.195 $Y=2.155
+ $X2=0 $Y2=0
cc_959 N_A_1799_408#_M1022_g N_VPWR_c_1627_n 0.0110654f $X=12.24 $Y=2.465 $X2=0
+ $Y2=0
cc_960 N_A_1799_408#_M1040_g N_VPWR_c_1627_n 0.0118221f $X=12.67 $Y=2.465 $X2=0
+ $Y2=0
cc_961 N_A_1799_408#_M1009_g N_VPWR_c_1627_n 0.00410284f $X=13.195 $Y=2.155
+ $X2=0 $Y2=0
cc_962 N_A_1799_408#_c_1414_n N_VPWR_c_1627_n 0.0290003f $X=9.665 $Y=2.72 $X2=0
+ $Y2=0
cc_963 N_A_1799_408#_c_1419_n N_VPWR_c_1627_n 0.0229522f $X=11.065 $Y=2.67 $X2=0
+ $Y2=0
cc_964 N_A_1799_408#_c_1456_n N_VPWR_c_1627_n 0.00557571f $X=10.535 $Y=2.67
+ $X2=0 $Y2=0
cc_965 N_A_1799_408#_c_1414_n A_1904_492# 0.00165422f $X=9.665 $Y=2.72 $X2=-0.19
+ $Y2=-0.245
cc_966 N_A_1799_408#_c_1416_n A_1904_492# 0.00107328f $X=9.75 $Y=2.555 $X2=-0.19
+ $Y2=-0.245
cc_967 N_A_1799_408#_M1028_g N_Q_N_c_1930_n 7.54206e-19 $X=11.5 $Y=0.875 $X2=0
+ $Y2=0
cc_968 N_A_1799_408#_M1018_g N_Q_N_c_1930_n 0.0168112f $X=12.09 $Y=0.665 $X2=0
+ $Y2=0
cc_969 N_A_1799_408#_M1022_g N_Q_N_c_1930_n 0.00844614f $X=12.24 $Y=2.465 $X2=0
+ $Y2=0
cc_970 N_A_1799_408#_M1037_g N_Q_N_c_1930_n 0.0171897f $X=12.52 $Y=0.665 $X2=0
+ $Y2=0
cc_971 N_A_1799_408#_M1040_g N_Q_N_c_1930_n 0.00771396f $X=12.67 $Y=2.465 $X2=0
+ $Y2=0
cc_972 N_A_1799_408#_c_1401_n N_Q_N_c_1930_n 0.0177218f $X=12.745 $Y=1.42 $X2=0
+ $Y2=0
cc_973 N_A_1799_408#_M1042_g N_Q_N_c_1930_n 0.0012801f $X=13.045 $Y=0.455 $X2=0
+ $Y2=0
cc_974 N_A_1799_408#_c_1409_n N_Q_N_c_1930_n 5.93685e-19 $X=11.79 $Y=1.51 $X2=0
+ $Y2=0
cc_975 N_A_1799_408#_M1010_g N_Q_N_c_1935_n 8.32713e-19 $X=11.715 $Y=2.045 $X2=0
+ $Y2=0
cc_976 N_A_1799_408#_M1022_g N_Q_N_c_1935_n 0.0134085f $X=12.24 $Y=2.465 $X2=0
+ $Y2=0
cc_977 N_A_1799_408#_M1010_g N_Q_N_c_1932_n 5.93685e-19 $X=11.715 $Y=2.045 $X2=0
+ $Y2=0
cc_978 N_A_1799_408#_M1022_g N_Q_N_c_1932_n 0.0125329f $X=12.24 $Y=2.465 $X2=0
+ $Y2=0
cc_979 N_A_1799_408#_M1040_g N_Q_N_c_1932_n 8.58208e-19 $X=12.67 $Y=2.465 $X2=0
+ $Y2=0
cc_980 N_A_1799_408#_c_1401_n N_Q_N_c_1932_n 0.0018554f $X=12.745 $Y=1.42 $X2=0
+ $Y2=0
cc_981 N_A_1799_408#_c_1405_n N_VGND_c_1987_n 0.00425916f $X=9.665 $Y=0.725
+ $X2=0 $Y2=0
cc_982 N_A_1799_408#_M1028_g N_VGND_c_1988_n 0.0128601f $X=11.5 $Y=0.875 $X2=0
+ $Y2=0
cc_983 N_A_1799_408#_M1018_g N_VGND_c_1988_n 0.00551624f $X=12.09 $Y=0.665 $X2=0
+ $Y2=0
cc_984 N_A_1799_408#_c_1409_n N_VGND_c_1988_n 9.30313e-19 $X=11.79 $Y=1.51 $X2=0
+ $Y2=0
cc_985 N_A_1799_408#_M1037_g N_VGND_c_1989_n 0.00471817f $X=12.52 $Y=0.665 $X2=0
+ $Y2=0
cc_986 N_A_1799_408#_c_1401_n N_VGND_c_1989_n 0.00842547f $X=12.745 $Y=1.42
+ $X2=0 $Y2=0
cc_987 N_A_1799_408#_M1042_g N_VGND_c_1989_n 0.00901344f $X=13.045 $Y=0.455
+ $X2=0 $Y2=0
cc_988 N_A_1799_408#_M1042_g N_VGND_c_1990_n 0.00575161f $X=13.045 $Y=0.455
+ $X2=0 $Y2=0
cc_989 N_A_1799_408#_M1042_g N_VGND_c_1991_n 0.00378367f $X=13.045 $Y=0.455
+ $X2=0 $Y2=0
cc_990 N_A_1799_408#_c_1405_n N_VGND_c_2002_n 0.014476f $X=9.665 $Y=0.725 $X2=0
+ $Y2=0
cc_991 N_A_1799_408#_M1028_g N_VGND_c_2005_n 0.0032821f $X=11.5 $Y=0.875 $X2=0
+ $Y2=0
cc_992 N_A_1799_408#_M1018_g N_VGND_c_2006_n 0.00561834f $X=12.09 $Y=0.665 $X2=0
+ $Y2=0
cc_993 N_A_1799_408#_M1037_g N_VGND_c_2006_n 0.00554431f $X=12.52 $Y=0.665 $X2=0
+ $Y2=0
cc_994 N_A_1799_408#_M1028_g N_VGND_c_2012_n 0.00385154f $X=11.5 $Y=0.875 $X2=0
+ $Y2=0
cc_995 N_A_1799_408#_M1018_g N_VGND_c_2012_n 0.0115933f $X=12.09 $Y=0.665 $X2=0
+ $Y2=0
cc_996 N_A_1799_408#_M1037_g N_VGND_c_2012_n 0.0103951f $X=12.52 $Y=0.665 $X2=0
+ $Y2=0
cc_997 N_A_1799_408#_M1042_g N_VGND_c_2012_n 0.0120944f $X=13.045 $Y=0.455 $X2=0
+ $Y2=0
cc_998 N_A_1799_408#_c_1405_n N_VGND_c_2012_n 0.0190889f $X=9.665 $Y=0.725 $X2=0
+ $Y2=0
cc_999 N_A_2624_49#_c_1574_n N_VPWR_c_1634_n 0.0268602f $X=13.41 $Y=1.98 $X2=0
+ $Y2=0
cc_1000 N_A_2624_49#_M1014_g N_VPWR_c_1635_n 0.0222944f $X=14.405 $Y=2.465 $X2=0
+ $Y2=0
cc_1001 N_A_2624_49#_M1044_g N_VPWR_c_1635_n 9.1316e-19 $X=14.835 $Y=2.465 $X2=0
+ $Y2=0
cc_1002 N_A_2624_49#_c_1574_n N_VPWR_c_1635_n 0.0285516f $X=13.41 $Y=1.98 $X2=0
+ $Y2=0
cc_1003 N_A_2624_49#_c_1575_n N_VPWR_c_1635_n 0.0230893f $X=14.27 $Y=1.44 $X2=0
+ $Y2=0
cc_1004 N_A_2624_49#_c_1578_n N_VPWR_c_1635_n 0.00757143f $X=14.835 $Y=1.44
+ $X2=0 $Y2=0
cc_1005 N_A_2624_49#_M1044_g N_VPWR_c_1637_n 0.00720408f $X=14.835 $Y=2.465
+ $X2=0 $Y2=0
cc_1006 N_A_2624_49#_M1014_g N_VPWR_c_1652_n 0.00486043f $X=14.405 $Y=2.465
+ $X2=0 $Y2=0
cc_1007 N_A_2624_49#_M1044_g N_VPWR_c_1652_n 0.00564131f $X=14.835 $Y=2.465
+ $X2=0 $Y2=0
cc_1008 N_A_2624_49#_M1014_g N_VPWR_c_1627_n 0.00824727f $X=14.405 $Y=2.465
+ $X2=0 $Y2=0
cc_1009 N_A_2624_49#_M1044_g N_VPWR_c_1627_n 0.0110855f $X=14.835 $Y=2.465 $X2=0
+ $Y2=0
cc_1010 N_A_2624_49#_c_1574_n N_VPWR_c_1627_n 0.0121821f $X=13.41 $Y=1.98 $X2=0
+ $Y2=0
cc_1011 N_A_2624_49#_M1007_g Q 0.00340711f $X=14.035 $Y=0.655 $X2=0 $Y2=0
cc_1012 N_A_2624_49#_M1014_g Q 0.0064279f $X=14.405 $Y=2.465 $X2=0 $Y2=0
cc_1013 N_A_2624_49#_M1015_g Q 0.0100708f $X=14.835 $Y=0.655 $X2=0 $Y2=0
cc_1014 N_A_2624_49#_M1044_g Q 0.025153f $X=14.835 $Y=2.465 $X2=0 $Y2=0
cc_1015 N_A_2624_49#_c_1575_n Q 0.0256674f $X=14.27 $Y=1.44 $X2=0 $Y2=0
cc_1016 N_A_2624_49#_c_1578_n Q 0.0314822f $X=14.835 $Y=1.44 $X2=0 $Y2=0
cc_1017 N_A_2624_49#_M1007_g N_Q_c_1960_n 0.00137803f $X=14.035 $Y=0.655 $X2=0
+ $Y2=0
cc_1018 N_A_2624_49#_M1015_g N_Q_c_1960_n 0.011261f $X=14.835 $Y=0.655 $X2=0
+ $Y2=0
cc_1019 N_A_2624_49#_c_1575_n N_Q_c_1960_n 0.0197123f $X=14.27 $Y=1.44 $X2=0
+ $Y2=0
cc_1020 N_A_2624_49#_c_1578_n N_Q_c_1960_n 0.0118278f $X=14.835 $Y=1.44 $X2=0
+ $Y2=0
cc_1021 N_A_2624_49#_c_1573_n N_VGND_c_1989_n 0.0249455f $X=13.37 $Y=1.275 $X2=0
+ $Y2=0
cc_1022 N_A_2624_49#_c_1576_n N_VGND_c_1990_n 0.0174874f $X=13.37 $Y=0.455 $X2=0
+ $Y2=0
cc_1023 N_A_2624_49#_M1007_g N_VGND_c_1991_n 0.00847481f $X=14.035 $Y=0.655
+ $X2=0 $Y2=0
cc_1024 N_A_2624_49#_c_1573_n N_VGND_c_1991_n 0.0363167f $X=13.37 $Y=1.275 $X2=0
+ $Y2=0
cc_1025 N_A_2624_49#_c_1575_n N_VGND_c_1991_n 0.0231067f $X=14.27 $Y=1.44 $X2=0
+ $Y2=0
cc_1026 N_A_2624_49#_c_1576_n N_VGND_c_1991_n 0.026119f $X=13.37 $Y=0.455 $X2=0
+ $Y2=0
cc_1027 N_A_2624_49#_c_1578_n N_VGND_c_1991_n 0.00519251f $X=14.835 $Y=1.44
+ $X2=0 $Y2=0
cc_1028 N_A_2624_49#_M1015_g N_VGND_c_1993_n 0.00827062f $X=14.835 $Y=0.655
+ $X2=0 $Y2=0
cc_1029 N_A_2624_49#_M1007_g N_VGND_c_2007_n 0.00585385f $X=14.035 $Y=0.655
+ $X2=0 $Y2=0
cc_1030 N_A_2624_49#_M1015_g N_VGND_c_2007_n 0.00564131f $X=14.835 $Y=0.655
+ $X2=0 $Y2=0
cc_1031 N_A_2624_49#_M1042_d N_VGND_c_2012_n 0.00266853f $X=13.12 $Y=0.245 $X2=0
+ $Y2=0
cc_1032 N_A_2624_49#_M1007_g N_VGND_c_2012_n 0.0125413f $X=14.035 $Y=0.655 $X2=0
+ $Y2=0
cc_1033 N_A_2624_49#_M1015_g N_VGND_c_2012_n 0.0117775f $X=14.835 $Y=0.655 $X2=0
+ $Y2=0
cc_1034 N_A_2624_49#_c_1576_n N_VGND_c_2012_n 0.0127213f $X=13.37 $Y=0.455 $X2=0
+ $Y2=0
cc_1035 N_VPWR_M1021_d N_A_268_467#_c_1806_n 0.0276724f $X=2.39 $Y=2.335 $X2=0
+ $Y2=0
cc_1036 N_VPWR_c_1628_n N_A_268_467#_c_1806_n 0.00459348f $X=0.69 $Y=2.85 $X2=0
+ $Y2=0
cc_1037 N_VPWR_c_1638_n N_A_268_467#_c_1806_n 0.0144738f $X=4.1 $Y=3.33 $X2=0
+ $Y2=0
cc_1038 N_VPWR_c_1649_n N_A_268_467#_c_1806_n 0.0208997f $X=2.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1039 N_VPWR_c_1654_n N_A_268_467#_c_1806_n 0.0255255f $X=2.61 $Y=3.07 $X2=0
+ $Y2=0
cc_1040 N_VPWR_c_1627_n N_A_268_467#_c_1806_n 0.0475688f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1041 N_VPWR_M1021_d N_A_268_467#_c_1802_n 0.00441108f $X=2.39 $Y=2.335 $X2=0
+ $Y2=0
cc_1042 N_VPWR_c_1629_n N_A_268_467#_c_1808_n 0.0163171f $X=4.195 $Y=2.84 $X2=0
+ $Y2=0
cc_1043 N_VPWR_c_1638_n N_A_268_467#_c_1808_n 0.0306168f $X=4.1 $Y=3.33 $X2=0
+ $Y2=0
cc_1044 N_VPWR_c_1627_n N_A_268_467#_c_1808_n 0.0247217f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1045 N_VPWR_c_1629_n N_A_268_467#_c_1809_n 0.00988817f $X=4.195 $Y=2.84 $X2=0
+ $Y2=0
cc_1046 N_VPWR_M1006_s N_A_268_467#_c_1810_n 0.0195224f $X=4.05 $Y=1.945 $X2=0
+ $Y2=0
cc_1047 N_VPWR_c_1629_n N_A_268_467#_c_1810_n 0.0205372f $X=4.195 $Y=2.84 $X2=0
+ $Y2=0
cc_1048 N_VPWR_c_1627_n N_A_268_467#_c_1810_n 0.0414575f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1049 N_VPWR_c_1650_n N_A_268_467#_c_1813_n 0.00556665f $X=6.79 $Y=3.33 $X2=0
+ $Y2=0
cc_1050 N_VPWR_c_1627_n N_A_268_467#_c_1813_n 0.00800162f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1051 N_VPWR_c_1627_n N_Q_N_M1022_s 0.00258346f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1052 N_VPWR_c_1646_n N_Q_N_c_1935_n 0.0169299f $X=12.755 $Y=3.33 $X2=0 $Y2=0
cc_1053 N_VPWR_c_1627_n N_Q_N_c_1935_n 0.0112082f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1054 N_VPWR_c_1634_n N_Q_N_c_1932_n 0.0016168f $X=12.93 $Y=1.98 $X2=0 $Y2=0
cc_1055 N_VPWR_c_1627_n N_Q_M1014_d 0.00380103f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1635_n Q 0.0476491f $X=14.19 $Y=1.985 $X2=0 $Y2=0
cc_1057 N_VPWR_c_1637_n Q 0.0456941f $X=15.05 $Y=1.985 $X2=0 $Y2=0
cc_1058 N_VPWR_c_1652_n Q 0.0150063f $X=14.945 $Y=3.33 $X2=0 $Y2=0
cc_1059 N_VPWR_c_1627_n Q 0.00950443f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1060 N_A_268_467#_c_1806_n A_376_467# 0.00639212f $X=3.06 $Y=2.695 $X2=-0.19
+ $Y2=-0.245
cc_1061 N_A_268_467#_c_1796_n N_VGND_c_1983_n 0.0082008f $X=2.055 $Y=0.445 $X2=0
+ $Y2=0
cc_1062 N_A_268_467#_c_1800_n N_VGND_c_1983_n 0.00706412f $X=3.06 $Y=1.28 $X2=0
+ $Y2=0
cc_1063 N_A_268_467#_c_1796_n N_VGND_c_1996_n 0.0131634f $X=2.055 $Y=0.445 $X2=0
+ $Y2=0
cc_1064 N_A_268_467#_c_1797_n N_VGND_c_1996_n 0.00717712f $X=2.52 $Y=0.79 $X2=0
+ $Y2=0
cc_1065 N_A_268_467#_c_1803_n N_VGND_c_2000_n 0.00516835f $X=5.525 $Y=0.805
+ $X2=0 $Y2=0
cc_1066 N_A_268_467#_M1016_d N_VGND_c_2012_n 0.00829206f $X=1.7 $Y=0.235 $X2=0
+ $Y2=0
cc_1067 N_A_268_467#_c_1796_n N_VGND_c_2012_n 0.00941296f $X=2.055 $Y=0.445
+ $X2=0 $Y2=0
cc_1068 N_A_268_467#_c_1797_n N_VGND_c_2012_n 0.0116807f $X=2.52 $Y=0.79 $X2=0
+ $Y2=0
cc_1069 N_A_268_467#_c_1803_n N_VGND_c_2012_n 0.00768579f $X=5.525 $Y=0.805
+ $X2=0 $Y2=0
cc_1070 N_Q_N_c_1930_n N_VGND_c_1989_n 0.0319331f $X=12.305 $Y=0.43 $X2=0 $Y2=0
cc_1071 N_Q_N_c_1930_n N_VGND_c_2006_n 0.0161961f $X=12.305 $Y=0.43 $X2=0 $Y2=0
cc_1072 N_Q_N_M1018_d N_VGND_c_2012_n 0.00223819f $X=12.165 $Y=0.245 $X2=0 $Y2=0
cc_1073 N_Q_N_c_1930_n N_VGND_c_2012_n 0.0114725f $X=12.305 $Y=0.43 $X2=0 $Y2=0
cc_1074 N_Q_c_1960_n N_VGND_c_1991_n 0.0340252f $X=14.62 $Y=0.42 $X2=0 $Y2=0
cc_1075 N_Q_c_1960_n N_VGND_c_1993_n 0.0358485f $X=14.62 $Y=0.42 $X2=0 $Y2=0
cc_1076 N_Q_c_1960_n N_VGND_c_2007_n 0.0426186f $X=14.62 $Y=0.42 $X2=0 $Y2=0
cc_1077 N_Q_M1007_s N_VGND_c_2012_n 0.00530851f $X=14.11 $Y=0.235 $X2=0 $Y2=0
cc_1078 N_Q_c_1960_n N_VGND_c_2012_n 0.0256387f $X=14.62 $Y=0.42 $X2=0 $Y2=0
cc_1079 N_VGND_c_2012_n A_268_47# 0.00768839f $X=15.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1080 N_VGND_c_2012_n A_471_47# 0.00265676f $X=15.12 $Y=0 $X2=-0.19 $Y2=-0.245
