* File: sky130_fd_sc_lp__o2111a_m.spice
* Created: Fri Aug 28 11:00:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111a_m.pex.spice"
.subckt sky130_fd_sc_lp__o2111a_m  VNB VPB D1 C1 B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_80_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_348_47# N_D1_M1000_g N_A_80_21#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.21 PD=0.63 PS=1.84 NRD=14.28 NRS=67.14 M=1 R=2.8 SA=75000.4
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 A_420_47# N_C1_M1007_g A_348_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.8 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_492_47#_M1009_d N_B1_M1009_g A_420_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_492_47#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_492_47#_M1006_d N_A1_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_80_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_80_21#_M1011_d N_D1_M1011_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75000.7
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_C1_M1008_g N_A_80_21#_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.11445 AS=0.0588 PD=0.965 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1010 N_A_80_21#_M1010_d N_B1_M1010_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.11445 PD=0.7 PS=0.965 NRD=0 NRS=114.91 M=1 R=2.8 SA=75001.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_564_535# N_A2_M1003_g N_A_80_21#_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_564_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_89 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o2111a_m.pxi.spice"
*
.ends
*
*
