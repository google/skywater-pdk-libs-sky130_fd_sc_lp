* File: sky130_fd_sc_lp__o32a_4.pex.spice
* Created: Fri Aug 28 11:17:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32A_4%A2 3 7 11 14 16 19 23 24 26 27 28 37 40 42 51
c92 40 0 1.55487e-19 $X=2.21 $Y=1.275
c93 16 0 1.53236e-19 $X=2.01 $Y=1.78
r94 36 42 8.90524 $w=4.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.77 $Y=1.645
+ $X2=1.11 $Y2=1.645
r95 35 37 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=0.77 $Y=1.51 $X2=0.9
+ $Y2=1.51
r96 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.51 $X2=0.77 $Y2=1.51
r97 32 35 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.56 $Y=1.51
+ $X2=0.77 $Y2=1.51
r98 28 51 7.9186 $w=4.38e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=1.645 $X2=1.33
+ $Y2=1.645
r99 28 42 2.35727 $w=4.38e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.645 $X2=1.11
+ $Y2=1.645
r100 27 36 1.30959 $w=4.38e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.645
+ $X2=0.77 $Y2=1.645
r101 26 27 12.5721 $w=4.38e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.645
+ $X2=0.72 $Y2=1.645
r102 24 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.44
+ $X2=2.21 $Y2=1.605
r103 24 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.44
+ $X2=2.21 $Y2=1.275
r104 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.44 $X2=2.21 $Y2=1.44
r105 20 23 5.00117 $w=2.63e-07 $l=1.15e-07 $layer=LI1_cond $X=2.095 $Y=1.402
+ $X2=2.21 $Y2=1.402
r106 18 20 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.095 $Y=1.535
+ $X2=2.095 $Y2=1.402
r107 18 19 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.095 $Y=1.535
+ $X2=2.095 $Y2=1.695
r108 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.01 $Y=1.78
+ $X2=2.095 $Y2=1.695
r109 16 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.01 $Y=1.78
+ $X2=1.33 $Y2=1.78
r110 14 41 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.23 $Y=2.465
+ $X2=2.23 $Y2=1.605
r111 11 40 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.19 $Y=0.745
+ $X2=2.19 $Y2=1.275
r112 5 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=1.675
+ $X2=0.9 $Y2=1.51
r113 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.9 $Y=1.675 $X2=0.9
+ $Y2=2.465
r114 1 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.345
+ $X2=0.56 $Y2=1.51
r115 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.56 $Y=1.345 $X2=0.56
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%A1 1 3 6 8 10 13 15 22
r53 20 22 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.665 $Y=1.44
+ $X2=1.76 $Y2=1.44
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.44 $X2=1.665 $Y2=1.44
r55 17 20 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.33 $Y=1.44
+ $X2=1.665 $Y2=1.44
r56 15 21 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.665 $Y=1.295
+ $X2=1.665 $Y2=1.44
r57 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.605
+ $X2=1.76 $Y2=1.44
r58 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.76 $Y=1.605
+ $X2=1.76 $Y2=2.465
r59 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.275
+ $X2=1.76 $Y2=1.44
r60 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.76 $Y=1.275
+ $X2=1.76 $Y2=0.745
r61 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.605
+ $X2=1.33 $Y2=1.44
r62 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.33 $Y=1.605 $X2=1.33
+ $Y2=2.465
r63 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.275
+ $X2=1.33 $Y2=1.44
r64 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.33 $Y=1.275 $X2=1.33
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%A3 1 3 6 10 12 14 15 16 17 26
c53 6 0 1.53236e-19 $X=2.66 $Y=2.465
c54 1 0 1.62159e-19 $X=2.66 $Y=1.275
r55 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.44 $X2=3.18 $Y2=1.44
r56 26 28 9.9528 $w=3.39e-07 $l=7e-08 $layer=POLY_cond $X=3.11 $Y=1.43 $X2=3.18
+ $Y2=1.43
r57 25 26 2.84366 $w=3.39e-07 $l=2e-08 $layer=POLY_cond $X=3.09 $Y=1.43 $X2=3.11
+ $Y2=1.43
r58 23 25 35.5457 $w=3.39e-07 $l=2.5e-07 $layer=POLY_cond $X=2.84 $Y=1.43
+ $X2=3.09 $Y2=1.43
r59 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.44 $X2=2.84 $Y2=1.44
r60 17 29 14.8931 $w=3.23e-07 $l=4.2e-07 $layer=LI1_cond $X=3.6 $Y=1.372
+ $X2=3.18 $Y2=1.372
r61 16 29 2.12759 $w=3.23e-07 $l=6e-08 $layer=LI1_cond $X=3.12 $Y=1.372 $X2=3.18
+ $Y2=1.372
r62 16 24 9.92874 $w=3.23e-07 $l=2.8e-07 $layer=LI1_cond $X=3.12 $Y=1.372
+ $X2=2.84 $Y2=1.372
r63 15 24 7.09196 $w=3.23e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=1.372 $X2=2.84
+ $Y2=1.372
r64 12 26 21.8644 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.11 $Y=1.255
+ $X2=3.11 $Y2=1.43
r65 12 14 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.11 $Y=1.255
+ $X2=3.11 $Y2=0.745
r66 8 25 21.8644 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.09 $Y=1.605
+ $X2=3.09 $Y2=1.43
r67 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.09 $Y=1.605
+ $X2=3.09 $Y2=2.465
r68 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.66 $Y=1.605 $X2=2.66
+ $Y2=2.465
r69 1 23 25.5929 $w=3.39e-07 $l=1.8e-07 $layer=POLY_cond $X=2.66 $Y=1.43
+ $X2=2.84 $Y2=1.43
r70 1 4 21.8644 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.66 $Y=1.43 $X2=2.66
+ $Y2=1.605
r71 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.66 $Y=1.275 $X2=2.66
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%B2 3 5 7 11 15 19 23 24 25 30 34 40
c97 30 0 1.49418e-19 $X=5.46 $Y=1.51
c98 25 0 1.67221e-19 $X=5.52 $Y=1.665
r99 31 34 7.72661 $w=4.38e-07 $l=2.95e-07 $layer=LI1_cond $X=5.46 $Y=1.645
+ $X2=5.165 $Y2=1.645
r100 30 33 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=5.442 $Y=1.51
+ $X2=5.442 $Y2=1.675
r101 30 32 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=5.442 $Y=1.51
+ $X2=5.442 $Y2=1.345
r102 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.46
+ $Y=1.51 $X2=5.46 $Y2=1.51
r103 25 31 1.57151 $w=4.38e-07 $l=6e-08 $layer=LI1_cond $X=5.52 $Y=1.645
+ $X2=5.46 $Y2=1.645
r104 24 34 3.27399 $w=4.38e-07 $l=1.25e-07 $layer=LI1_cond $X=5.04 $Y=1.645
+ $X2=5.165 $Y2=1.645
r105 24 40 7.00188 $w=4.38e-07 $l=9.5e-08 $layer=LI1_cond $X=5.04 $Y=1.645
+ $X2=4.945 $Y2=1.645
r106 23 40 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.195 $Y=1.78
+ $X2=4.945 $Y2=1.78
r107 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.51 $X2=4.025 $Y2=1.51
r108 17 23 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=4.027 $Y=1.695
+ $X2=4.195 $Y2=1.78
r109 17 19 6.36424 $w=3.33e-07 $l=1.85e-07 $layer=LI1_cond $X=4.027 $Y=1.695
+ $X2=4.027 $Y2=1.51
r110 15 32 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.34 $Y=0.745 $X2=5.34
+ $Y2=1.345
r111 11 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.335 $Y=2.465
+ $X2=5.335 $Y2=1.675
r112 5 20 38.5938 $w=3.29e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.04 $Y=1.675
+ $X2=4.025 $Y2=1.51
r113 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.04 $Y=1.675
+ $X2=4.04 $Y2=2.465
r114 1 20 38.5938 $w=3.29e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.975 $Y=1.345
+ $X2=4.025 $Y2=1.51
r115 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.975 $Y=1.345 $X2=3.975
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%B1 1 3 6 8 10 13 15 22
c53 8 0 2.39709e-19 $X=4.905 $Y=1.275
c54 1 0 6.53712e-20 $X=4.475 $Y=1.275
r55 20 22 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=4.61 $Y=1.44
+ $X2=4.905 $Y2=1.44
r56 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.61
+ $Y=1.44 $X2=4.61 $Y2=1.44
r57 17 20 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.475 $Y=1.44
+ $X2=4.61 $Y2=1.44
r58 15 21 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.61 $Y=1.295
+ $X2=4.61 $Y2=1.44
r59 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.605
+ $X2=4.905 $Y2=1.44
r60 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.905 $Y=1.605
+ $X2=4.905 $Y2=2.465
r61 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.275
+ $X2=4.905 $Y2=1.44
r62 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.905 $Y=1.275
+ $X2=4.905 $Y2=0.745
r63 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.475 $Y=1.605
+ $X2=4.475 $Y2=1.44
r64 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.475 $Y=1.605
+ $X2=4.475 $Y2=2.465
r65 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.475 $Y=1.275
+ $X2=4.475 $Y2=1.44
r66 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.475 $Y=1.275
+ $X2=4.475 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%A_547_367# 1 2 3 4 5 18 22 26 30 34 38 42 46
+ 48 50 52 54 57 58 60 62 66 69 75 83 86 104
c159 104 0 1.67221e-19 $X=7.655 $Y=1.49
c160 86 0 1.49418e-19 $X=5.12 $Y=0.7
c161 62 0 5.52737e-20 $X=5.795 $Y=1.165
r162 101 102 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.795 $Y=1.49
+ $X2=7.225 $Y2=1.49
r163 88 89 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.12 $Y=0.955
+ $X2=5.12 $Y2=1.165
r164 86 88 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.12 $Y=0.7
+ $X2=5.12 $Y2=0.955
r165 83 84 10.8226 $w=3.1e-07 $l=2.75e-07 $layer=LI1_cond $X=4.19 $Y=0.68
+ $X2=4.19 $Y2=0.955
r166 76 104 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.475 $Y=1.49
+ $X2=7.655 $Y2=1.49
r167 76 102 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.475 $Y=1.49
+ $X2=7.225 $Y2=1.49
r168 75 76 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.475
+ $Y=1.49 $X2=7.475 $Y2=1.49
r169 73 101 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.455 $Y=1.49
+ $X2=6.795 $Y2=1.49
r170 73 98 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.455 $Y=1.49
+ $X2=6.365 $Y2=1.49
r171 72 75 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=6.455 $Y=1.49
+ $X2=7.475 $Y2=1.49
r172 72 73 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.455
+ $Y=1.49 $X2=6.455 $Y2=1.49
r173 70 97 6.52558 $w=1.9e-07 $l=2.53e-07 $layer=LI1_cond $X=6.3 $Y=1.49
+ $X2=6.047 $Y2=1.49
r174 70 72 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=6.3 $Y=1.49
+ $X2=6.455 $Y2=1.49
r175 69 92 32.4246 $w=1.68e-07 $l=4.97e-07 $layer=LI1_cond $X=6.047 $Y=2.12
+ $X2=5.55 $Y2=2.12
r176 68 97 2.25005 $w=5.03e-07 $l=9.5e-08 $layer=LI1_cond $X=6.047 $Y=1.585
+ $X2=6.047 $Y2=1.49
r177 68 69 10.6581 $w=5.03e-07 $l=4.5e-07 $layer=LI1_cond $X=6.047 $Y=1.585
+ $X2=6.047 $Y2=2.035
r178 66 92 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=5.585 $Y=2.515
+ $X2=5.585 $Y2=2.205
r179 63 89 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=1.165
+ $X2=5.12 $Y2=1.165
r180 62 97 7.69753 $w=5.03e-07 $l=3.25e-07 $layer=LI1_cond $X=6.047 $Y=1.165
+ $X2=6.047 $Y2=1.49
r181 62 63 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.795 $Y=1.165
+ $X2=5.285 $Y2=1.165
r182 61 84 4.25403 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=0.955
+ $X2=4.19 $Y2=0.955
r183 60 88 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.955 $Y=0.955
+ $X2=5.12 $Y2=0.955
r184 60 61 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.955 $Y=0.955
+ $X2=4.355 $Y2=0.955
r185 59 81 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.92 $Y=2.12
+ $X2=3.79 $Y2=2.12
r186 58 92 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.455 $Y=2.12
+ $X2=5.55 $Y2=2.12
r187 58 59 100.144 $w=1.68e-07 $l=1.535e-06 $layer=LI1_cond $X=5.455 $Y=2.12
+ $X2=3.92 $Y2=2.12
r188 55 57 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=3.79 $Y=2.905
+ $X2=3.79 $Y2=2.52
r189 54 81 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=2.205
+ $X2=3.79 $Y2=2.12
r190 54 57 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.79 $Y=2.205
+ $X2=3.79 $Y2=2.52
r191 53 79 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=2.99
+ $X2=2.875 $Y2=2.99
r192 52 55 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.66 $Y=2.99
+ $X2=3.79 $Y2=2.905
r193 52 53 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.66 $Y=2.99
+ $X2=3.04 $Y2=2.99
r194 48 79 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=2.905
+ $X2=2.875 $Y2=2.99
r195 48 50 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=2.875 $Y=2.905
+ $X2=2.875 $Y2=2.13
r196 44 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.655
+ $X2=7.655 $Y2=1.49
r197 44 46 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.655 $Y=1.655
+ $X2=7.655 $Y2=2.465
r198 40 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.325
+ $X2=7.655 $Y2=1.49
r199 40 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.655 $Y=1.325
+ $X2=7.655 $Y2=0.665
r200 36 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.655
+ $X2=7.225 $Y2=1.49
r201 36 38 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.225 $Y=1.655
+ $X2=7.225 $Y2=2.465
r202 32 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.325
+ $X2=7.225 $Y2=1.49
r203 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.225 $Y=1.325
+ $X2=7.225 $Y2=0.665
r204 28 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.655
+ $X2=6.795 $Y2=1.49
r205 28 30 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.795 $Y=1.655
+ $X2=6.795 $Y2=2.465
r206 24 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.325
+ $X2=6.795 $Y2=1.49
r207 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.795 $Y=1.325
+ $X2=6.795 $Y2=0.665
r208 20 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.655
+ $X2=6.365 $Y2=1.49
r209 20 22 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.365 $Y=1.655
+ $X2=6.365 $Y2=2.465
r210 16 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.325
+ $X2=6.365 $Y2=1.49
r211 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.365 $Y=1.325
+ $X2=6.365 $Y2=0.665
r212 5 92 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.835 $X2=5.55 $Y2=2.12
r213 5 66 300 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=2 $X=5.41
+ $Y=1.835 $X2=5.55 $Y2=2.515
r214 4 81 600 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=1.835 $X2=3.825 $Y2=2.12
r215 4 57 300 $w=1.7e-07 $l=7.44883e-07 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=1.835 $X2=3.825 $Y2=2.52
r216 3 79 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.735
+ $Y=1.835 $X2=2.875 $Y2=2.91
r217 3 50 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.735
+ $Y=1.835 $X2=2.875 $Y2=2.13
r218 2 86 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=4.98
+ $Y=0.325 $X2=5.12 $Y2=0.7
r219 1 83 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=4.05
+ $Y=0.325 $X2=4.19 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%A_112_367# 1 2 3 10 12 14 22 24 25 28
r47 26 28 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=3.34 $Y=1.875
+ $X2=3.34 $Y2=1.98
r48 24 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.21 $Y=1.79
+ $X2=3.34 $Y2=1.875
r49 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.21 $Y=1.79
+ $X2=2.54 $Y2=1.79
r50 20 32 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=2.205
+ $X2=2.445 $Y2=2.12
r51 20 22 14.3014 $w=1.88e-07 $l=2.45e-07 $layer=LI1_cond $X=2.445 $Y=2.205
+ $X2=2.445 $Y2=2.45
r52 17 32 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=2.035
+ $X2=2.445 $Y2=2.12
r53 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=2.445 $Y=2.035
+ $X2=2.445 $Y2=1.98
r54 16 25 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.445 $Y=1.875
+ $X2=2.54 $Y2=1.79
r55 16 19 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=2.445 $Y=1.875
+ $X2=2.445 $Y2=1.98
r56 15 31 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.78 $Y=2.12 $X2=0.65
+ $Y2=2.12
r57 14 32 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.35 $Y=2.12
+ $X2=2.445 $Y2=2.12
r58 14 15 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=2.35 $Y=2.12
+ $X2=0.78 $Y2=2.12
r59 10 31 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=2.205
+ $X2=0.65 $Y2=2.12
r60 10 12 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.65 $Y=2.205
+ $X2=0.65 $Y2=2.52
r61 3 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.835 $X2=3.305 $Y2=1.98
r62 2 22 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=2.305
+ $Y=1.835 $X2=2.445 $Y2=2.45
r63 2 19 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=1.835 $X2=2.445 $Y2=1.98
r64 1 31 600 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.685 $Y2=2.12
r65 1 12 300 $w=1.7e-07 $l=7.44883e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=1.835 $X2=0.685 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%A_195_367# 1 2 7 9 11 13 15
r23 13 20 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=2.545 $X2=2.03
+ $Y2=2.46
r24 13 15 14.0214 $w=2.98e-07 $l=3.65e-07 $layer=LI1_cond $X=2.03 $Y=2.545
+ $X2=2.03 $Y2=2.91
r25 12 18 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.21 $Y=2.46 $X2=1.08
+ $Y2=2.46
r26 11 20 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.88 $Y=2.46 $X2=2.03
+ $Y2=2.46
r27 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.88 $Y=2.46
+ $X2=1.21 $Y2=2.46
r28 7 18 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=2.545 $X2=1.08
+ $Y2=2.46
r29 7 9 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=1.08 $Y=2.545
+ $X2=1.08 $Y2=2.91
r30 2 20 600 $w=1.7e-07 $l=7.09313e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.835 $X2=2.015 $Y2=2.46
r31 2 15 600 $w=1.7e-07 $l=1.16152e-06 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.835 $X2=2.015 $Y2=2.91
r32 1 18 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.835 $X2=1.115 $Y2=2.46
r33 1 9 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.835 $X2=1.115 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%VPWR 1 2 3 4 5 18 20 24 28 32 36 38 42 44 52
+ 57 62 68 71 74 77 81 88
r113 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r116 72 88 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.32 $Y2=3.33
r117 71 72 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 68 69 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r119 66 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 66 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 63 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=3.33
+ $X2=7.01 $Y2=3.33
r123 63 65 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.175 $Y=3.33
+ $X2=7.44 $Y2=3.33
r124 62 80 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.932 $Y2=3.33
r125 62 65 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.44 $Y2=3.33
r126 61 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r127 61 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r128 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r129 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.315 $Y=3.33
+ $X2=6.15 $Y2=3.33
r130 58 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.315 $Y=3.33
+ $X2=6.48 $Y2=3.33
r131 57 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=3.33
+ $X2=7.01 $Y2=3.33
r132 57 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.845 $Y=3.33
+ $X2=6.48 $Y2=3.33
r133 56 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r134 56 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r136 53 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.69 $Y2=3.33
r137 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.04 $Y2=3.33
r138 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=3.33
+ $X2=6.15 $Y2=3.33
r139 52 55 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=5.985 $Y=3.33
+ $X2=5.04 $Y2=3.33
r140 51 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r141 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r143 46 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r144 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r145 44 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=3.33
+ $X2=1.545 $Y2=3.33
r146 44 50 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.38 $Y=3.33
+ $X2=1.2 $Y2=3.33
r147 42 88 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.32 $Y2=3.33
r148 42 69 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=1.68 $Y2=3.33
r149 38 41 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=7.87 $Y=2.18
+ $X2=7.87 $Y2=2.95
r150 36 80 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=7.87 $Y=3.245
+ $X2=7.932 $Y2=3.33
r151 36 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.87 $Y=3.245
+ $X2=7.87 $Y2=2.95
r152 32 35 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=7.01 $Y=2.18
+ $X2=7.01 $Y2=2.95
r153 30 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=3.245
+ $X2=7.01 $Y2=3.33
r154 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.01 $Y=3.245
+ $X2=7.01 $Y2=2.95
r155 26 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.15 $Y=3.245
+ $X2=6.15 $Y2=3.33
r156 26 28 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.15 $Y=3.245
+ $X2=6.15 $Y2=2.475
r157 22 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=3.33
r158 22 24 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=2.835
r159 21 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=3.33
+ $X2=1.545 $Y2=3.33
r160 20 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.69 $Y2=3.33
r161 20 21 183.652 $w=1.68e-07 $l=2.815e-06 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=1.71 $Y2=3.33
r162 16 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=3.245
+ $X2=1.545 $Y2=3.33
r163 16 18 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.545 $Y=3.245
+ $X2=1.545 $Y2=2.84
r164 5 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.835 $X2=7.87 $Y2=2.95
r165 5 38 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.835 $X2=7.87 $Y2=2.18
r166 4 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.87
+ $Y=1.835 $X2=7.01 $Y2=2.95
r167 4 32 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=6.87
+ $Y=1.835 $X2=7.01 $Y2=2.18
r168 3 28 300 $w=1.7e-07 $l=6.99714e-07 $layer=licon1_PDIFF $count=2 $X=6.025
+ $Y=1.835 $X2=6.15 $Y2=2.475
r169 2 24 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=4.55
+ $Y=1.835 $X2=4.69 $Y2=2.835
r170 1 18 600 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.835 $X2=1.545 $Y2=2.84
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%A_823_367# 1 2 7 9 11 13 15
r24 13 20 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=2.545
+ $X2=5.155 $Y2=2.46
r25 13 15 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=2.545
+ $X2=5.155 $Y2=2.91
r26 12 18 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.355 $Y=2.46
+ $X2=4.222 $Y2=2.46
r27 11 20 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.025 $Y=2.46
+ $X2=5.155 $Y2=2.46
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.025 $Y=2.46
+ $X2=4.355 $Y2=2.46
r29 7 18 2.82608 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.222 $Y=2.545
+ $X2=4.222 $Y2=2.46
r30 7 9 15.8733 $w=2.63e-07 $l=3.65e-07 $layer=LI1_cond $X=4.222 $Y=2.545
+ $X2=4.222 $Y2=2.91
r31 2 20 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.835 $X2=5.12 $Y2=2.46
r32 2 15 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.835 $X2=5.12 $Y2=2.91
r33 1 18 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.835 $X2=4.255 $Y2=2.46
r34 1 9 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.835 $X2=4.255 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41 42
+ 44 45 49 51
r59 49 51 3.04419 $w=2.63e-07 $l=7e-08 $layer=LI1_cond $X=7.942 $Y=1.225
+ $X2=7.942 $Y2=1.295
r60 44 49 2.8391 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.942 $Y=1.14
+ $X2=7.942 $Y2=1.225
r61 44 45 15.7863 $w=2.63e-07 $l=3.63e-07 $layer=LI1_cond $X=7.942 $Y=1.302
+ $X2=7.942 $Y2=1.665
r62 44 51 0.304419 $w=2.63e-07 $l=7e-09 $layer=LI1_cond $X=7.942 $Y=1.302
+ $X2=7.942 $Y2=1.295
r63 43 45 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=7.942 $Y=1.755
+ $X2=7.942 $Y2=1.665
r64 40 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.535 $Y=1.84
+ $X2=7.44 $Y2=1.84
r65 39 43 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=7.81 $Y=1.84
+ $X2=7.942 $Y2=1.755
r66 39 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.81 $Y=1.84
+ $X2=7.535 $Y2=1.84
r67 38 41 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.525 $Y=1.14 $X2=7.435
+ $Y2=1.14
r68 37 44 4.40896 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.81 $Y=1.14
+ $X2=7.942 $Y2=1.14
r69 37 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.81 $Y=1.14
+ $X2=7.525 $Y2=1.14
r70 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=7.44 $Y=1.98
+ $X2=7.44 $Y2=2.91
r71 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.44 $Y=1.925
+ $X2=7.44 $Y2=1.84
r72 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=7.44 $Y=1.925
+ $X2=7.44 $Y2=1.98
r73 27 41 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=1.055
+ $X2=7.435 $Y2=1.14
r74 27 29 39.1263 $w=1.78e-07 $l=6.35e-07 $layer=LI1_cond $X=7.435 $Y=1.055
+ $X2=7.435 $Y2=0.42
r75 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.345 $Y=1.84
+ $X2=7.44 $Y2=1.84
r76 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.345 $Y=1.84
+ $X2=6.675 $Y2=1.84
r77 23 41 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.345 $Y=1.14 $X2=7.435
+ $Y2=1.14
r78 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.345 $Y=1.14
+ $X2=6.665 $Y2=1.14
r79 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.58 $Y=1.98
+ $X2=6.58 $Y2=2.91
r80 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.58 $Y=1.925
+ $X2=6.675 $Y2=1.84
r81 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.58 $Y=1.925
+ $X2=6.58 $Y2=1.98
r82 13 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.575 $Y=1.055
+ $X2=6.665 $Y2=1.14
r83 13 15 39.1263 $w=1.78e-07 $l=6.35e-07 $layer=LI1_cond $X=6.575 $Y=1.055
+ $X2=6.575 $Y2=0.42
r84 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.835 $X2=7.44 $Y2=2.91
r85 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.835 $X2=7.44 $Y2=1.98
r86 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.835 $X2=6.58 $Y2=2.91
r87 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.835 $X2=6.58 $Y2=1.98
r88 2 29 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=7.3
+ $Y=0.245 $X2=7.44 $Y2=0.42
r89 1 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=6.44
+ $Y=0.245 $X2=6.58 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%A_44_65# 1 2 3 4 5 6 21 23 24 27 29 30 33 35
+ 41 42 43 47 50 51
c87 51 0 1.84435e-19 $X=4.655 $Y=0.34
c88 43 0 6.53712e-20 $X=5.465 $Y=0.345
c89 33 0 3.17646e-19 $X=2.435 $Y=0.47
r90 53 55 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=4.655 $Y=0.345
+ $X2=4.655 $Y2=0.535
r91 51 53 0.221624 $w=2.58e-07 $l=5e-09 $layer=LI1_cond $X=4.655 $Y=0.34
+ $X2=4.655 $Y2=0.345
r92 45 47 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=5.63 $Y=0.435
+ $X2=5.63 $Y2=0.47
r93 44 53 2.89065 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.785 $Y=0.345
+ $X2=4.655 $Y2=0.345
r94 43 45 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.465 $Y=0.345
+ $X2=5.63 $Y2=0.435
r95 43 44 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=5.465 $Y=0.345
+ $X2=4.785 $Y2=0.345
r96 41 51 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.525 $Y=0.34
+ $X2=4.655 $Y2=0.34
r97 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.525 $Y=0.34
+ $X2=3.855 $Y2=0.34
r98 38 40 7.6549 $w=6.23e-07 $l=4e-07 $layer=LI1_cond $X=3.542 $Y=0.87 $X2=3.542
+ $Y2=0.47
r99 37 42 10.24 $w=1.7e-07 $l=3.5295e-07 $layer=LI1_cond $X=3.542 $Y=0.425
+ $X2=3.855 $Y2=0.34
r100 37 40 0.861176 $w=6.23e-07 $l=4.5e-08 $layer=LI1_cond $X=3.542 $Y=0.425
+ $X2=3.542 $Y2=0.47
r101 36 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.56 $Y=0.955
+ $X2=2.435 $Y2=0.955
r102 35 38 10.24 $w=1.7e-07 $l=3.51943e-07 $layer=LI1_cond $X=3.23 $Y=0.955
+ $X2=3.542 $Y2=0.87
r103 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.23 $Y=0.955
+ $X2=2.56 $Y2=0.955
r104 31 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.87
+ $X2=2.435 $Y2=0.955
r105 31 33 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=2.435 $Y=0.87
+ $X2=2.435 $Y2=0.47
r106 30 49 7.02746 $w=2.46e-07 $l=1.54771e-07 $layer=LI1_cond $X=1.64 $Y=0.955
+ $X2=1.522 $Y2=1.04
r107 29 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.31 $Y=0.955
+ $X2=2.435 $Y2=0.955
r108 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.31 $Y=0.955
+ $X2=1.64 $Y2=0.955
r109 25 49 1.01869 $w=2.35e-07 $l=1.7e-07 $layer=LI1_cond $X=1.522 $Y=0.87
+ $X2=1.522 $Y2=1.04
r110 25 27 20.5969 $w=2.33e-07 $l=4.2e-07 $layer=LI1_cond $X=1.522 $Y=0.87
+ $X2=1.522 $Y2=0.45
r111 23 49 19.1283 $w=2.46e-07 $l=4.22024e-07 $layer=LI1_cond $X=1.16 $Y=1.17
+ $X2=1.522 $Y2=1.04
r112 23 24 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.16 $Y=1.17
+ $X2=0.44 $Y2=1.17
r113 19 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.31 $Y=1.085
+ $X2=0.44 $Y2=1.17
r114 19 21 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=0.31 $Y=1.085
+ $X2=0.31 $Y2=0.47
r115 6 47 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=5.415
+ $Y=0.325 $X2=5.63 $Y2=0.47
r116 5 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.55
+ $Y=0.325 $X2=4.69 $Y2=0.535
r117 4 40 45.5 $w=1.7e-07 $l=6.43428e-07 $layer=licon1_NDIFF $count=4 $X=3.185
+ $Y=0.325 $X2=3.76 $Y2=0.47
r118 3 33 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.325 $X2=2.435 $Y2=0.47
r119 2 27 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.325 $X2=1.545 $Y2=0.45
r120 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.325 $X2=0.345 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_4%VGND 1 2 3 4 5 6 21 25 29 33 35 37 40 41 43
+ 44 45 47 59 63 68 77 81 84 88 97
r109 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r110 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r111 82 97 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.32
+ $Y2=0
r112 81 82 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6
+ $Y2=0
r113 77 79 8.26381 $w=5.61e-07 $l=3.8e-07 $layer=LI1_cond $X=0.922 $Y=0.45
+ $X2=0.922 $Y2=0.83
r114 74 77 9.7861 $w=5.61e-07 $l=4.5e-07 $layer=LI1_cond $X=0.922 $Y=0 $X2=0.922
+ $Y2=0.45
r115 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r116 72 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r117 72 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r118 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r119 69 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=0 $X2=7.01
+ $Y2=0
r120 69 71 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.175 $Y=0
+ $X2=7.44 $Y2=0
r121 68 87 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=7.705 $Y=0
+ $X2=7.932 $Y2=0
r122 68 71 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.705 $Y=0
+ $X2=7.44 $Y2=0
r123 67 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r124 67 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r125 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r126 64 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.315 $Y=0 $X2=6.15
+ $Y2=0
r127 64 66 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.315 $Y=0
+ $X2=6.48 $Y2=0
r128 63 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=0 $X2=7.01
+ $Y2=0
r129 63 66 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.845 $Y=0
+ $X2=6.48 $Y2=0
r130 61 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r131 59 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=0 $X2=6.15
+ $Y2=0
r132 59 61 186.914 $w=1.68e-07 $l=2.865e-06 $layer=LI1_cond $X=5.985 $Y=0
+ $X2=3.12 $Y2=0
r133 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r134 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r135 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r136 55 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r137 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r138 52 74 7.88553 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=0.922 $Y2=0
r139 52 54 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=1.68 $Y2=0
r140 50 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r141 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r142 47 74 7.88553 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.922
+ $Y2=0
r143 47 49 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.24
+ $Y2=0
r144 45 97 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.32 $Y2=0
r145 45 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r146 43 57 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.64
+ $Y2=0
r147 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.895
+ $Y2=0
r148 42 61 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.06 $Y=0 $X2=3.12
+ $Y2=0
r149 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=0 $X2=2.895
+ $Y2=0
r150 40 54 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.68
+ $Y2=0
r151 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.975
+ $Y2=0
r152 39 57 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.64
+ $Y2=0
r153 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=1.975
+ $Y2=0
r154 35 87 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.932 $Y2=0
r155 35 37 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0.39
r156 31 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0
r157 31 33 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0.37
r158 27 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0
r159 27 29 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0.39
r160 23 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0
r161 23 25 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0.595
r162 19 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0
r163 19 21 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0.595
r164 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.73
+ $Y=0.245 $X2=7.87 $Y2=0.39
r165 5 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.87
+ $Y=0.245 $X2=7.01 $Y2=0.37
r166 4 29 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.025
+ $Y=0.245 $X2=6.15 $Y2=0.39
r167 3 25 182 $w=1.7e-07 $l=3.40734e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.325 $X2=2.895 $Y2=0.595
r168 2 21 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=1.835
+ $Y=0.325 $X2=1.975 $Y2=0.595
r169 1 79 121.333 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1
+ $X=0.635 $Y=0.325 $X2=0.775 $Y2=0.83
r170 1 77 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1
+ $X=0.635 $Y=0.325 $X2=0.775 $Y2=0.45
.ends

