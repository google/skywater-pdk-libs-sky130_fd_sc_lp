* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__invkapwr_2 A KAPWR VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.226e+11p ps=2.74e+06u
M1001 KAPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=6.867e+11p ps=6.13e+06u
M1002 KAPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A KAPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
