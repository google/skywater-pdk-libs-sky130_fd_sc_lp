* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 VGND a_91_123# a_260_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_483_123# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_359_123# a_91_123# a_454_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_1143_125# a_1203_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1199_449# a_1203_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 Q a_1673_409# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Q a_1673_409# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND a_1475_449# a_1673_409# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND a_1673_409# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_359_123# SCE a_483_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1475_449# a_641_123# a_1670_61# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1203_99# a_850_51# a_1475_449# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND CLK a_641_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_359_123# a_850_51# a_1053_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_1631_507# a_1673_409# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 Q a_1673_409# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VPWR a_1673_409# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR a_1053_125# a_1203_99# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 a_1053_125# a_850_51# a_1143_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR a_1475_449# a_1673_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR CLK a_641_123# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_641_123# a_850_51# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VPWR a_1673_409# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_454_491# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_91_123# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_1203_99# a_641_123# a_1475_449# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X26 a_1670_61# a_1673_409# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VPWR SCE a_296_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_296_491# D a_359_123# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_91_123# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_1053_125# a_641_123# a_1199_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_1475_449# a_850_51# a_1631_507# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 a_260_123# D a_359_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VGND a_1673_409# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 Q a_1673_409# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 VGND a_641_123# a_850_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VGND a_1053_125# a_1203_99# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X37 a_359_123# a_641_123# a_1053_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
