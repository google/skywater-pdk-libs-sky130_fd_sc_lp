* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VGND CLK a_1161_95# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1033_121# a_1075_95# a_722_23# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_2040_125# a_2082_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_196_119# D a_304_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_2409_367# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND a_2409_367# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND a_2082_99# a_2409_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND SCE a_324_431# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_196_119# a_1075_95# a_722_23# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1075_95# a_1161_95# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_2082_99# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR a_767_121# a_974_425# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VGND a_1873_497# a_2082_99# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VPWR CLK a_1161_95# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_1786_497# a_1075_95# a_1873_497# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_722_23# a_1161_95# a_196_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1873_497# a_1161_95# a_767_121# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_722_23# a_1161_95# a_974_425# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 VPWR SCE a_196_483# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_196_483# D a_196_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_767_121# a_722_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1786_497# a_2082_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VPWR a_1873_497# a_2082_99# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 a_27_483# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 VGND a_767_121# a_1033_121# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_767_121# a_1075_95# a_1873_497# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_324_431# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1873_497# a_1161_95# a_2040_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_2409_367# a_2082_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_196_119# a_324_431# a_27_483# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_124_119# SCE a_196_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_767_121# a_722_23# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 a_304_119# a_324_431# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VGND SCD a_124_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1075_95# a_1161_95# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 Q a_2082_99# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
