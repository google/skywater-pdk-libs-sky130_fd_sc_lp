* File: sky130_fd_sc_lp__fa_1.spice
* Created: Fri Aug 28 10:34:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fa_1.pex.spice"
.subckt sky130_fd_sc_lp__fa_1  VNB VPB A B CIN COUT VPWR SUM VGND
* 
* VGND	VGND
* SUM	SUM
* VPWR	VPWR
* COUT	COUT
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_A_80_27#_M1016_g N_COUT_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.252 AS=0.2226 PD=1.96667 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1006 A_267_137# N_A_M1006_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.126 PD=0.66 PS=0.983333 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1026 N_A_80_27#_M1026_d N_B_M1026_g A_267_137# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_A_431_137#_M1001_d N_CIN_M1001_g N_A_80_27#_M1026_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_M1020_g N_A_431_137#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1021 N_A_431_137#_M1021_d N_B_M1021_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1022 N_A_818_83#_M1022_d N_B_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.05985 AS=0.1113 PD=0.705 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_CIN_M1024_g N_A_818_83#_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.05985 PD=0.715 PS=0.705 NRD=4.284 NRS=1.428 M=1 R=2.8
+ SA=75000.6 SB=75002 A=0.063 P=1.14 MULT=1
MM1007 N_A_818_83#_M1007_d N_A_M1007_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.42
+ AD=0.13755 AS=0.06195 PD=1.14 PS=0.715 NRD=32.136 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_1118_411#_M1025_d N_A_80_27#_M1025_g N_A_818_83#_M1007_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.13755 PD=0.7 PS=1.14 NRD=0 NRS=34.992 M=1 R=2.8
+ SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1027 A_1212_125# N_CIN_M1027_g N_A_1118_411#_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1014 A_1290_125# N_B_M1014_g A_1212_125# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8 SA=75001.8 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g A_1290_125# VNB NSHORT L=0.15 W=0.42 AD=0.0966
+ AS=0.0882 PD=0.843333 PS=0.84 NRD=42.852 NRS=44.28 M=1 R=2.8 SA=75002.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1023 N_SUM_M1023_d N_A_1118_411#_M1023_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1932 PD=2.25 PS=1.68667 NRD=2.856 NRS=0 M=1 R=5.6
+ SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_A_80_27#_M1017_g N_COUT_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.319725 AS=0.3339 PD=2.5575 PS=3.05 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 A_231_457# N_A_M1004_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0735
+ AS=0.106575 PD=0.77 PS=0.8525 NRD=56.2829 NRS=70.3487 M=1 R=2.8 SA=75000.8
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1008 N_A_80_27#_M1008_d N_B_M1008_g A_231_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=56.2829 M=1 R=2.8 SA=75001.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_417_457#_M1015_d N_CIN_M1015_g N_A_80_27#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_417_457#_M1015_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.117775 AS=0.0588 PD=1.035 PS=0.7 NRD=105.73 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1012 N_A_417_457#_M1012_d N_B_M1012_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.117775 PD=1.37 PS=1.035 NRD=0 NRS=105.73 M=1 R=2.8 SA=75002.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_854_411#_M1002_d N_B_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0651 AS=0.1113 PD=0.73 PS=1.37 NRD=14.0658 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.7 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_CIN_M1003_g N_A_854_411#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0651 PD=0.7 PS=0.73 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_854_411#_M1010_d N_A_M1010_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1018 N_A_1118_411#_M1018_d N_A_80_27#_M1018_g N_A_854_411#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=18.7544 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1011 A_1212_411# N_CIN_M1011_g N_A_1118_411#_M1018_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0672 PD=0.66 PS=0.74 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75002
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1000 A_1290_411# N_B_M1000_g A_1212_411# VPB PHIGHVT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=72.693 NRS=30.4759 M=1 R=2.8 SA=75002.4
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A_M1019_g A_1290_411# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.120225 AS=0.0882 PD=0.925 PS=0.84 NRD=108.448 NRS=72.693 M=1 R=2.8
+ SA=75002.9 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1013 N_SUM_M1013_d N_A_1118_411#_M1013_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.360675 PD=3.05 PS=2.775 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.4 SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.9271 P=20.81
c_160 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__fa_1.pxi.spice"
*
.ends
*
*
