* File: sky130_fd_sc_lp__dlclkp_4.pex.spice
* Created: Wed Sep  2 09:45:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%A_73_269# 1 2 9 13 15 18 19 21 22 24 26 27
+ 31 35 37
c110 37 0 1.61743e-19 $X=1.675 $Y=2.365
c111 31 0 1.79399e-19 $X=1.12 $Y=1.645
r112 37 40 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.675 $Y=2.365
+ $X2=1.675 $Y2=2.57
r113 32 35 9.3636 $w=2.38e-07 $l=1.95e-07 $layer=LI1_cond $X=1.57 $Y=0.725
+ $X2=1.765 $Y2=0.725
r114 27 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.51
+ $X2=0.53 $Y2=1.675
r115 27 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.51
+ $X2=0.53 $Y2=1.345
r116 26 29 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.56 $Y=1.51
+ $X2=0.56 $Y2=1.645
r117 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.51 $X2=0.53 $Y2=1.51
r118 23 32 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.57 $Y=0.845
+ $X2=1.57 $Y2=0.725
r119 23 24 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.57 $Y=0.845
+ $X2=1.57 $Y2=1.56
r120 21 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=2.365
+ $X2=1.675 $Y2=2.365
r121 21 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.51 $Y=2.365
+ $X2=1.205 $Y2=2.365
r122 20 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.645
+ $X2=1.12 $Y2=1.645
r123 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=1.645
+ $X2=1.57 $Y2=1.56
r124 19 20 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.485 $Y=1.645
+ $X2=1.205 $Y2=1.645
r125 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=2.28
+ $X2=1.205 $Y2=2.365
r126 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.73
+ $X2=1.12 $Y2=1.645
r127 17 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.12 $Y=1.73
+ $X2=1.12 $Y2=2.28
r128 16 29 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.685 $Y=1.645
+ $X2=0.56 $Y2=1.645
r129 15 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=1.645
+ $X2=1.12 $Y2=1.645
r130 15 16 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.035 $Y=1.645
+ $X2=0.685 $Y2=1.645
r131 13 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.5 $Y=0.655
+ $X2=0.5 $Y2=1.345
r132 9 44 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.675
r133 2 40 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=2.325 $X2=1.675 $Y2=2.57
r134 1 35 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.405 $X2=1.765 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%GATE 3 7 9 12
c54 3 0 1.75443e-19 $X=1.1 $Y=2.645
r55 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.295
+ $X2=1.1 $Y2=1.13
r56 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.295 $X2=1.1 $Y2=1.295
r57 9 13 5.23838 $w=2.18e-07 $l=1e-07 $layer=LI1_cond $X=1.2 $Y=1.28 $X2=1.1
+ $Y2=1.28
r58 7 14 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.19 $Y=0.615
+ $X2=1.19 $Y2=1.13
r59 1 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.46 $X2=1.1
+ $Y2=1.295
r60 1 3 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=1.1 $Y=1.46 $X2=1.1
+ $Y2=2.645
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%A_277_367# 1 2 9 13 14 17 21 22 24 26 28 31
+ 32 34 39 46
c129 14 0 1.6638e-19 $X=1.835 $Y=2.005
c130 9 0 8.7847e-20 $X=1.46 $Y=2.645
r131 39 41 4.72258 $w=3.1e-07 $l=1.2e-07 $layer=LI1_cond $X=3.53 $Y=2.25
+ $X2=3.53 $Y2=2.37
r132 38 39 9.05161 $w=3.1e-07 $l=2.3e-07 $layer=LI1_cond $X=3.53 $Y=2.02
+ $X2=3.53 $Y2=2.25
r133 34 36 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=3.245 $Y=0.63
+ $X2=3.245 $Y2=0.71
r134 30 31 41.397 $w=3.78e-07 $l=1.365e-06 $layer=LI1_cond $X=4.89 $Y=0.795
+ $X2=4.89 $Y2=2.16
r135 29 39 3.91789 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=2.25
+ $X2=3.53 $Y2=2.25
r136 28 31 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=4.7 $Y=2.25
+ $X2=4.89 $Y2=2.16
r137 28 29 61.9242 $w=1.78e-07 $l=1.005e-06 $layer=LI1_cond $X=4.7 $Y=2.25
+ $X2=3.695 $Y2=2.25
r138 27 36 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.375 $Y=0.71
+ $X2=3.245 $Y2=0.71
r139 26 30 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=4.7 $Y=0.71
+ $X2=4.89 $Y2=0.795
r140 26 27 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=4.7 $Y=0.71
+ $X2=3.375 $Y2=0.71
r141 25 32 7.80489 $w=1.95e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.165 $Y=2.02
+ $X2=2 $Y2=2.005
r142 24 38 3.91789 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=2.02
+ $X2=3.53 $Y2=2.02
r143 24 25 73.9394 $w=1.78e-07 $l=1.2e-06 $layer=LI1_cond $X=3.365 $Y=2.02
+ $X2=2.165 $Y2=2.02
r144 22 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.1 $X2=2
+ $Y2=0.935
r145 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2 $Y=1.1
+ $X2=2 $Y2=1.1
r146 19 32 0.463323 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=2 $Y=1.9 $X2=2
+ $Y2=2.005
r147 19 21 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=2 $Y=1.9 $X2=2 $Y2=1.1
r148 17 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=2 $X2=1.55
+ $Y2=2.165
r149 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55 $Y=2
+ $X2=1.55 $Y2=2
r150 14 32 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=2.005
+ $X2=2 $Y2=2.005
r151 14 16 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=1.835 $Y=2.005
+ $X2=1.55 $Y2=2.005
r152 13 46 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.98 $Y=0.615
+ $X2=1.98 $Y2=0.935
r153 9 44 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.46 $Y=2.645
+ $X2=1.46 $Y2=2.165
r154 2 41 600 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=2.095 $X2=3.49 $Y2=2.37
r155 1 34 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.405 $X2=3.21 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%A_295_55# 1 2 9 11 12 15 19 22 25 28 29 30
+ 33 35 36 37 43 47
c114 37 0 1.83398e-19 $X=4.2 $Y=1.08
c115 36 0 1.89073e-19 $X=3.075 $Y=1.475
c116 19 0 1.34147e-19 $X=2.995 $Y=0.615
c117 12 0 1.6638e-19 $X=1.625 $Y=1.55
c118 11 0 1.61743e-19 $X=1.925 $Y=1.55
r119 47 51 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.14
+ $X2=3.1 $Y2=0.975
r120 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.085
+ $Y=1.14 $X2=3.085 $Y2=1.14
r121 41 43 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.365 $Y=1.195
+ $X2=4.365 $Y2=1.895
r122 38 46 4.02592 $w=2.3e-07 $l=1.55e-07 $layer=LI1_cond $X=3.23 $Y=1.08
+ $X2=3.075 $Y2=1.08
r123 38 40 47.6009 $w=2.28e-07 $l=9.5e-07 $layer=LI1_cond $X=3.23 $Y=1.08
+ $X2=4.18 $Y2=1.08
r124 37 41 7.10306 $w=2.3e-07 $l=2.14942e-07 $layer=LI1_cond $X=4.2 $Y=1.08
+ $X2=4.365 $Y2=1.195
r125 37 40 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=4.2 $Y=1.08 $X2=4.18
+ $Y2=1.08
r126 35 46 2.98697 $w=3.1e-07 $l=1.15e-07 $layer=LI1_cond $X=3.075 $Y=1.195
+ $X2=3.075 $Y2=1.08
r127 35 36 10.4092 $w=3.08e-07 $l=2.8e-07 $layer=LI1_cond $X=3.075 $Y=1.195
+ $X2=3.075 $Y2=1.475
r128 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.64 $X2=2.51 $Y2=1.64
r129 30 36 6.83216 $w=2.85e-07 $l=2.14558e-07 $layer=LI1_cond $X=2.92 $Y=1.617
+ $X2=3.075 $Y2=1.475
r130 30 32 16.579 $w=2.83e-07 $l=4.1e-07 $layer=LI1_cond $X=2.92 $Y=1.617
+ $X2=2.51 $Y2=1.617
r131 27 33 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=2.075 $Y=1.64
+ $X2=2.51 $Y2=1.64
r132 27 28 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=2.075 $Y=1.64 $X2=2
+ $Y2=1.64
r133 25 29 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.205 $Y=2.415
+ $X2=3.205 $Y2=1.645
r134 22 29 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=3.1 $Y=1.465 $X2=3.1
+ $Y2=1.645
r135 21 47 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=3.1 $Y=1.155
+ $X2=3.1 $Y2=1.14
r136 21 22 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=3.1 $Y=1.155
+ $X2=3.1 $Y2=1.465
r137 19 51 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.995 $Y=0.615
+ $X2=2.995 $Y2=0.975
r138 13 28 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.805 $X2=2
+ $Y2=1.64
r139 13 15 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2 $Y=1.805 $X2=2
+ $Y2=2.535
r140 11 28 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.925 $Y=1.55
+ $X2=2 $Y2=1.64
r141 11 12 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.925 $Y=1.55
+ $X2=1.625 $Y2=1.55
r142 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.55 $Y=1.475
+ $X2=1.625 $Y2=1.55
r143 7 9 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.55 $Y=1.475
+ $X2=1.55 $Y2=0.615
r144 2 43 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=1.77 $X2=4.365 $Y2=1.895
r145 1 40 182 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.655 $X2=4.18 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%A_27_367# 1 2 9 13 14 15 16 18 21 25 31 33
+ 36 37 38 39 42 43 44 46 48 50 51 54 55 61 62 63 64 68 75 76 80 81 82 87 90 97
c246 87 0 1.3918e-19 $X=5.885 $Y=1.535
c247 76 0 8.68225e-20 $X=2.54 $Y=1.1
c248 44 0 8.7847e-20 $X=2.19 $Y=2.365
c249 39 0 1.75443e-19 $X=2.02 $Y=2.99
c250 37 0 1.34147e-19 $X=2.345 $Y=0.35
r251 85 97 2.88623 $w=3.34e-07 $l=2e-08 $layer=POLY_cond $X=5.765 $Y=1.425
+ $X2=5.745 $Y2=1.425
r252 84 87 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=5.765 $Y=1.535
+ $X2=5.885 $Y2=1.535
r253 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.765
+ $Y=1.5 $X2=5.765 $Y2=1.5
r254 80 94 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.98 $Y=2.94
+ $X2=3.98 $Y2=3.15
r255 79 82 18.2906 $w=5.63e-07 $l=5.6e-07 $layer=LI1_cond $X=3.98 $Y=2.792
+ $X2=4.54 $Y2=2.792
r256 79 81 6.12322 $w=5.63e-07 $l=1.75e-07 $layer=LI1_cond $X=3.98 $Y=2.792
+ $X2=3.805 $Y2=2.792
r257 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.98
+ $Y=2.94 $X2=3.98 $Y2=2.94
r258 76 90 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.54 $Y=1.1
+ $X2=2.54 $Y2=0.935
r259 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.1 $X2=2.54 $Y2=1.1
r260 72 75 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=2.43 $Y=1.14
+ $X2=2.54 $Y2=1.14
r261 68 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.2 $Y=2.715
+ $X2=1.2 $Y2=2.99
r262 63 66 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=0.265 $Y=2.715
+ $X2=0.265 $Y2=2.91
r263 63 64 2.88111 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.715
+ $X2=0.265 $Y2=2.63
r264 61 62 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.26 $Y2=1.9
r265 59 62 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.18 $Y=1.095
+ $X2=0.18 $Y2=1.9
r266 58 59 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=0.93
+ $X2=0.272 $Y2=1.095
r267 55 58 0.486948 $w=3.53e-07 $l=1.5e-08 $layer=LI1_cond $X=0.272 $Y=0.915
+ $X2=0.272 $Y2=0.93
r268 55 56 3.24083 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=0.272 $Y=0.915
+ $X2=0.272 $Y2=0.83
r269 53 87 2.89065 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=5.885 $Y=1.665
+ $X2=5.885 $Y2=1.535
r270 53 54 52.0657 $w=1.78e-07 $l=8.45e-07 $layer=LI1_cond $X=5.885 $Y=1.665
+ $X2=5.885 $Y2=2.51
r271 51 54 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.795 $Y=2.595
+ $X2=5.885 $Y2=2.51
r272 51 82 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=5.795 $Y=2.595
+ $X2=4.54 $Y2=2.595
r273 50 81 22.6771 $w=3.08e-07 $l=6.1e-07 $layer=LI1_cond $X=3.195 $Y=2.92
+ $X2=3.805 $Y2=2.92
r274 48 50 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=3.11 $Y=2.765
+ $X2=3.195 $Y2=2.92
r275 47 48 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.11 $Y=2.45
+ $X2=3.11 $Y2=2.765
r276 46 72 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.43 $Y=1.015
+ $X2=2.43 $Y2=1.14
r277 45 46 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.43 $Y=0.435
+ $X2=2.43 $Y2=1.015
r278 43 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=2.365
+ $X2=3.11 $Y2=2.45
r279 43 44 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.025 $Y=2.365
+ $X2=2.19 $Y2=2.365
r280 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.105 $Y=2.45
+ $X2=2.19 $Y2=2.365
r281 41 42 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.105 $Y=2.45
+ $X2=2.105 $Y2=2.905
r282 40 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.99
+ $X2=1.2 $Y2=2.99
r283 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.02 $Y=2.99
+ $X2=2.105 $Y2=2.905
r284 39 40 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.02 $Y=2.99
+ $X2=1.285 $Y2=2.99
r285 37 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.345 $Y=0.35
+ $X2=2.43 $Y2=0.435
r286 37 38 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.345 $Y=0.35
+ $X2=1.23 $Y2=0.35
r287 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=0.435
+ $X2=1.23 $Y2=0.35
r288 35 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.145 $Y=0.435
+ $X2=1.145 $Y2=0.83
r289 34 55 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.45 $Y=0.915
+ $X2=0.272 $Y2=0.915
r290 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=0.915
+ $X2=1.145 $Y2=0.83
r291 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.06 $Y=0.915
+ $X2=0.45 $Y2=0.915
r292 32 63 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.435 $Y=2.715
+ $X2=0.265 $Y2=2.715
r293 31 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.715
+ $X2=1.2 $Y2=2.715
r294 31 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.115 $Y=2.715
+ $X2=0.435 $Y2=2.715
r295 29 61 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.26 $Y=2.065
+ $X2=0.26 $Y2=2.015
r296 29 64 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.26 $Y=2.065
+ $X2=0.26 $Y2=2.63
r297 25 56 16.579 $w=2.83e-07 $l=4.1e-07 $layer=LI1_cond $X=0.237 $Y=0.42
+ $X2=0.237 $Y2=0.83
r298 19 97 21.5099 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.745 $Y=1.665
+ $X2=5.745 $Y2=1.425
r299 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.745 $Y=1.665
+ $X2=5.745 $Y2=2.465
r300 16 97 47.6228 $w=3.34e-07 $l=4.33705e-07 $layer=POLY_cond $X=5.415 $Y=1.185
+ $X2=5.745 $Y2=1.425
r301 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.415 $Y=1.185
+ $X2=5.415 $Y2=0.655
r302 14 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.98 $Y2=3.15
r303 14 15 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=2.435 $Y2=3.15
r304 13 90 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.45 $Y=0.615
+ $X2=2.45 $Y2=0.935
r305 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.36 $Y=3.075
+ $X2=2.435 $Y2=3.15
r306 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.36 $Y=3.075
+ $X2=2.36 $Y2=2.535
r307 2 66 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r308 2 61 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.015
r309 1 58 182 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.93
r310 1 25 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%CLK 1 5 9 11 12 15 19 24 26 29 30
c76 29 0 1.02251e-19 $X=3.685 $Y=1.53
c77 24 0 1.3918e-19 $X=5.315 $Y=1.62
c78 15 0 1.83398e-19 $X=5.055 $Y=0.655
r79 29 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.685 $Y=1.53
+ $X2=3.685 $Y2=1.62
r80 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=1.53 $X2=3.685 $Y2=1.53
r81 26 30 3.58824 $w=4.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.625 $Y=1.665
+ $X2=3.625 $Y2=1.53
r82 23 24 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.055 $Y=1.62
+ $X2=5.315 $Y2=1.62
r83 21 22 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.51 $Y=1.62
+ $X2=4.695 $Y2=1.62
r84 17 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.315 $Y=1.695
+ $X2=5.315 $Y2=1.62
r85 17 19 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.315 $Y=1.695
+ $X2=5.315 $Y2=2.465
r86 13 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.055 $Y=1.545
+ $X2=5.055 $Y2=1.62
r87 13 15 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.055 $Y=1.545
+ $X2=5.055 $Y2=0.655
r88 12 22 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.77 $Y=1.62
+ $X2=4.695 $Y2=1.62
r89 11 23 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.98 $Y=1.62
+ $X2=5.055 $Y2=1.62
r90 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.98 $Y=1.62
+ $X2=4.77 $Y2=1.62
r91 7 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.695 $Y=1.695
+ $X2=4.695 $Y2=1.62
r92 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.695 $Y=1.695
+ $X2=4.695 $Y2=2.155
r93 3 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.51 $Y=1.545
+ $X2=4.51 $Y2=1.62
r94 3 5 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.51 $Y=1.545 $X2=4.51
+ $Y2=0.865
r95 2 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=1.62
+ $X2=3.685 $Y2=1.62
r96 1 21 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.435 $Y=1.62
+ $X2=4.51 $Y2=1.62
r97 1 2 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=4.435 $Y=1.62
+ $X2=3.85 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%A_1078_367# 1 2 9 13 17 21 25 29 33 37 40
+ 43 45 48 51 54 58 71
r119 70 71 43.1182 $w=3.13e-07 $l=2.8e-07 $layer=POLY_cond $X=7.225 $Y=1.5
+ $X2=7.505 $Y2=1.5
r120 69 70 23.099 $w=3.13e-07 $l=1.5e-07 $layer=POLY_cond $X=7.075 $Y=1.5
+ $X2=7.225 $Y2=1.5
r121 66 67 23.099 $w=3.13e-07 $l=1.5e-07 $layer=POLY_cond $X=6.645 $Y=1.5
+ $X2=6.795 $Y2=1.5
r122 65 66 43.1182 $w=3.13e-07 $l=2.8e-07 $layer=POLY_cond $X=6.365 $Y=1.5
+ $X2=6.645 $Y2=1.5
r123 62 65 8.46965 $w=3.13e-07 $l=5.5e-08 $layer=POLY_cond $X=6.31 $Y=1.5
+ $X2=6.365 $Y2=1.5
r124 62 63 14.6294 $w=3.13e-07 $l=9.5e-08 $layer=POLY_cond $X=6.31 $Y=1.5
+ $X2=6.215 $Y2=1.5
r125 61 62 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=1.5 $X2=6.31 $Y2=1.5
r126 55 58 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.335 $Y=2.175
+ $X2=5.53 $Y2=2.175
r127 52 69 13.0895 $w=3.13e-07 $l=8.5e-08 $layer=POLY_cond $X=6.99 $Y=1.5
+ $X2=7.075 $Y2=1.5
r128 52 67 30.0288 $w=3.13e-07 $l=1.95e-07 $layer=POLY_cond $X=6.99 $Y=1.5
+ $X2=6.795 $Y2=1.5
r129 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.99
+ $Y=1.5 $X2=6.99 $Y2=1.5
r130 49 61 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.315 $Y=1.5
+ $X2=6.23 $Y2=1.5
r131 49 51 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.315 $Y=1.5
+ $X2=6.99 $Y2=1.5
r132 48 61 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.23 $Y=1.415
+ $X2=6.23 $Y2=1.5
r133 47 48 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.23 $Y=1.235
+ $X2=6.23 $Y2=1.415
r134 46 54 2.76166 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=5.795 $Y=1.15
+ $X2=5.522 $Y2=1.15
r135 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.145 $Y=1.15
+ $X2=6.23 $Y2=1.235
r136 45 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.145 $Y=1.15
+ $X2=5.795 $Y2=1.15
r137 41 54 3.70735 $w=2.5e-07 $l=1.44375e-07 $layer=LI1_cond $X=5.63 $Y=1.065
+ $X2=5.522 $Y2=1.15
r138 41 43 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=5.63 $Y=1.065
+ $X2=5.63 $Y2=0.42
r139 40 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.01
+ $X2=5.335 $Y2=2.175
r140 39 54 3.70735 $w=2.5e-07 $l=2.2553e-07 $layer=LI1_cond $X=5.335 $Y=1.235
+ $X2=5.522 $Y2=1.15
r141 39 40 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=5.335 $Y=1.235
+ $X2=5.335 $Y2=2.01
r142 35 71 23.099 $w=3.13e-07 $l=2.2798e-07 $layer=POLY_cond $X=7.655 $Y=1.335
+ $X2=7.505 $Y2=1.5
r143 35 37 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.655 $Y=1.335
+ $X2=7.655 $Y2=0.655
r144 31 71 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.505 $Y=1.665
+ $X2=7.505 $Y2=1.5
r145 31 33 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=7.505 $Y=1.665
+ $X2=7.505 $Y2=2.465
r146 27 70 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.335
+ $X2=7.225 $Y2=1.5
r147 27 29 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.225 $Y=1.335
+ $X2=7.225 $Y2=0.655
r148 23 69 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.075 $Y=1.665
+ $X2=7.075 $Y2=1.5
r149 23 25 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=7.075 $Y=1.665
+ $X2=7.075 $Y2=2.465
r150 19 67 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.335
+ $X2=6.795 $Y2=1.5
r151 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.795 $Y=1.335
+ $X2=6.795 $Y2=0.655
r152 15 66 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=1.665
+ $X2=6.645 $Y2=1.5
r153 15 17 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=6.645 $Y=1.665
+ $X2=6.645 $Y2=2.465
r154 11 65 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.365 $Y=1.335
+ $X2=6.365 $Y2=1.5
r155 11 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.365 $Y=1.335
+ $X2=6.365 $Y2=0.655
r156 7 63 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.215 $Y=1.665
+ $X2=6.215 $Y2=1.5
r157 7 9 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=6.215 $Y=1.665
+ $X2=6.215 $Y2=2.465
r158 2 58 600 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.835 $X2=5.53 $Y2=2.175
r159 1 43 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.49
+ $Y=0.235 $X2=5.63 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 44 45 46
+ 48 53 61 69 78 83 90 93 96 100
r108 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r109 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r110 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 83 86 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.77 $Y=3.065
+ $X2=0.77 $Y2=3.33
r114 81 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r115 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 78 99 3.91666 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.932 $Y2=3.33
r117 78 80 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 77 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r119 77 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r120 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 74 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.125 $Y=3.33
+ $X2=5.96 $Y2=3.33
r122 74 76 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.125 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 73 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r124 73 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 70 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.005 $Y2=3.33
r127 70 72 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 69 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=3.33
+ $X2=5.96 $Y2=3.33
r129 69 72 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.795 $Y=3.33
+ $X2=5.52 $Y2=3.33
r130 68 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r132 65 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r134 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r135 62 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.69 $Y2=3.33
r136 62 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r137 61 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=5.005 $Y2=3.33
r138 61 67 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r139 60 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r140 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 57 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r144 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r145 54 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.77 $Y2=3.33
r146 54 56 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.2 $Y2=3.33
r147 53 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.69 $Y2=3.33
r148 53 59 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r149 51 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r150 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r151 48 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.77 $Y2=3.33
r152 48 50 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 46 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 46 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r155 44 76 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.48 $Y2=3.33
r156 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.86 $Y2=3.33
r157 43 80 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=7.44 $Y2=3.33
r158 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=6.86 $Y2=3.33
r159 39 42 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=7.83 $Y=1.98
+ $X2=7.83 $Y2=2.95
r160 37 99 3.2265 $w=2.5e-07 $l=1.38109e-07 $layer=LI1_cond $X=7.83 $Y=3.245
+ $X2=7.932 $Y2=3.33
r161 37 42 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.83 $Y=3.245
+ $X2=7.83 $Y2=2.95
r162 33 36 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.86 $Y=2.27
+ $X2=6.86 $Y2=2.95
r163 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=3.33
r164 31 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=2.95
r165 27 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=3.245
+ $X2=5.96 $Y2=3.33
r166 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.96 $Y=3.245
+ $X2=5.96 $Y2=2.95
r167 23 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=3.33
r168 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=2.95
r169 19 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=3.33
r170 19 21 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=2.745
r171 6 42 400 $w=1.7e-07 $l=1.21547e-06 $layer=licon1_PDIFF $count=1 $X=7.58
+ $Y=1.835 $X2=7.79 $Y2=2.95
r172 6 39 400 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=7.58
+ $Y=1.835 $X2=7.79 $Y2=1.98
r173 5 36 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.72
+ $Y=1.835 $X2=6.86 $Y2=2.95
r174 5 33 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=6.72
+ $Y=1.835 $X2=6.86 $Y2=2.27
r175 4 29 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.835 $X2=5.96 $Y2=2.95
r176 3 25 600 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=4.77
+ $Y=1.835 $X2=5.005 $Y2=2.95
r177 2 21 600 $w=1.7e-07 $l=5.32447e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=2.325 $X2=2.69 $Y2=2.745
r178 1 83 600 $w=1.7e-07 $l=1.33548e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.77 $Y2=3.065
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%GCLK 1 2 3 4 13 15 19 21 23 24 27 28 29 30
+ 31 32 33 45 54 60
r54 58 60 1.69477 $w=3.38e-07 $l=5e-08 $layer=LI1_cond $X=7.365 $Y=1.985
+ $X2=7.365 $Y2=2.035
r55 51 54 3.08081 $w=1.78e-07 $l=5e-08 $layer=LI1_cond $X=7.445 $Y=1.245
+ $X2=7.445 $Y2=1.295
r56 33 67 4.57588 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=7.365 $Y=2.775
+ $X2=7.365 $Y2=2.91
r57 32 33 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=7.365 $Y=2.405
+ $X2=7.365 $Y2=2.775
r58 31 52 3.58051 $w=2.6e-07 $l=1.18427e-07 $layer=LI1_cond $X=7.365 $Y=1.9
+ $X2=7.445 $Y2=1.815
r59 31 58 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.365 $Y=1.9
+ $X2=7.365 $Y2=1.985
r60 31 32 11.9651 $w=3.38e-07 $l=3.53e-07 $layer=LI1_cond $X=7.365 $Y=2.052
+ $X2=7.365 $Y2=2.405
r61 31 60 0.576222 $w=3.38e-07 $l=1.7e-08 $layer=LI1_cond $X=7.365 $Y=2.052
+ $X2=7.365 $Y2=2.035
r62 30 52 9.24242 $w=1.78e-07 $l=1.5e-07 $layer=LI1_cond $X=7.445 $Y=1.665
+ $X2=7.445 $Y2=1.815
r63 29 43 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=7.44 $Y=1.16
+ $X2=7.44 $Y2=1.075
r64 29 51 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=7.44 $Y=1.16
+ $X2=7.445 $Y2=1.245
r65 29 30 21.7505 $w=1.78e-07 $l=3.53e-07 $layer=LI1_cond $X=7.445 $Y=1.312
+ $X2=7.445 $Y2=1.665
r66 29 54 1.04747 $w=1.78e-07 $l=1.7e-08 $layer=LI1_cond $X=7.445 $Y=1.312
+ $X2=7.445 $Y2=1.295
r67 28 43 8.75598 $w=1.88e-07 $l=1.5e-07 $layer=LI1_cond $X=7.44 $Y=0.925
+ $X2=7.44 $Y2=1.075
r68 27 28 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.44 $Y=0.555
+ $X2=7.44 $Y2=0.925
r69 27 45 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=7.44 $Y=0.555
+ $X2=7.44 $Y2=0.42
r70 23 29 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.345 $Y=1.16
+ $X2=7.44 $Y2=1.16
r71 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.345 $Y=1.16
+ $X2=6.675 $Y2=1.16
r72 22 26 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.525 $Y=1.9
+ $X2=6.41 $Y2=1.9
r73 21 31 2.90867 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.195 $Y=1.9
+ $X2=7.365 $Y2=1.9
r74 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.195 $Y=1.9
+ $X2=6.525 $Y2=1.9
r75 17 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.58 $Y=1.075
+ $X2=6.675 $Y2=1.16
r76 17 19 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=6.58 $Y=1.075
+ $X2=6.58 $Y2=0.42
r77 13 26 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=1.985 $X2=6.41
+ $Y2=1.9
r78 13 15 46.3483 $w=2.28e-07 $l=9.25e-07 $layer=LI1_cond $X=6.41 $Y=1.985
+ $X2=6.41 $Y2=2.91
r79 4 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.15
+ $Y=1.835 $X2=7.29 $Y2=1.98
r80 4 67 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.15
+ $Y=1.835 $X2=7.29 $Y2=2.91
r81 3 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.835 $X2=6.43 $Y2=1.98
r82 3 15 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.835 $X2=6.43 $Y2=2.91
r83 2 45 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.3
+ $Y=0.235 $X2=7.44 $Y2=0.42
r84 1 19 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.44
+ $Y=0.235 $X2=6.58 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 47 48 49 51 69 73 78 84 87 90 94
r98 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r99 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r100 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r101 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r102 82 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r103 82 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r104 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r105 79 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=0 $X2=7.01
+ $Y2=0
r106 79 81 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.175 $Y=0
+ $X2=7.44 $Y2=0
r107 78 93 4.38626 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.74 $Y=0 $X2=7.95
+ $Y2=0
r108 78 81 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.74 $Y=0 $X2=7.44
+ $Y2=0
r109 77 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r110 77 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r111 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r112 74 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.315 $Y=0 $X2=6.15
+ $Y2=0
r113 74 76 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.315 $Y=0
+ $X2=6.48 $Y2=0
r114 73 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=0 $X2=7.01
+ $Y2=0
r115 73 76 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.845 $Y=0
+ $X2=6.48 $Y2=0
r116 72 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r117 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r118 69 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=0 $X2=6.15
+ $Y2=0
r119 69 71 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=5.985 $Y=0
+ $X2=5.04 $Y2=0
r120 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r121 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r122 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r123 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r124 62 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r125 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r126 59 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r127 59 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r128 58 61 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r129 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r130 56 84 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.72
+ $Y2=0
r131 56 58 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r132 54 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r133 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r134 51 84 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.72
+ $Y2=0
r135 51 53 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r136 49 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r137 49 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r138 47 67 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.675 $Y=0
+ $X2=4.56 $Y2=0
r139 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=4.84
+ $Y2=0
r140 46 71 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.005 $Y=0 $X2=5.04
+ $Y2=0
r141 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=4.84
+ $Y2=0
r142 44 61 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.64
+ $Y2=0
r143 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.815
+ $Y2=0
r144 43 64 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.945 $Y=0
+ $X2=3.12 $Y2=0
r145 43 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.815
+ $Y2=0
r146 39 93 3.09127 $w=2.95e-07 $l=1.12161e-07 $layer=LI1_cond $X=7.887 $Y=0.085
+ $X2=7.95 $Y2=0
r147 39 41 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=7.887 $Y=0.085
+ $X2=7.887 $Y2=0.38
r148 35 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0
r149 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0.38
r150 31 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0
r151 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0.38
r152 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0
r153 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0.36
r154 23 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=0.085
+ $X2=2.815 $Y2=0
r155 23 25 23.4921 $w=2.58e-07 $l=5.3e-07 $layer=LI1_cond $X=2.815 $Y=0.085
+ $X2=2.815 $Y2=0.615
r156 19 84 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r157 19 21 15.2529 $w=3.38e-07 $l=4.5e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.535
r158 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.73
+ $Y=0.235 $X2=7.87 $Y2=0.38
r159 5 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.87
+ $Y=0.235 $X2=7.01 $Y2=0.38
r160 4 33 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.025
+ $Y=0.235 $X2=6.15 $Y2=0.38
r161 3 29 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.655 $X2=4.84 $Y2=0.36
r162 2 25 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.405 $X2=2.78 $Y2=0.615
r163 1 21 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.535
.ends

