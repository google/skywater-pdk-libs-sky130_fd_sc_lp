* File: sky130_fd_sc_lp__a21bo_2.pxi.spice
* Created: Wed Sep  2 09:18:47 2020
* 
x_PM_SKY130_FD_SC_LP__A21BO_2%A_22_259# N_A_22_259#_M1006_d N_A_22_259#_M1010_s
+ N_A_22_259#_c_73_n N_A_22_259#_M1000_g N_A_22_259#_M1001_g N_A_22_259#_c_75_n
+ N_A_22_259#_c_76_n N_A_22_259#_M1008_g N_A_22_259#_M1007_g N_A_22_259#_c_78_n
+ N_A_22_259#_c_79_n N_A_22_259#_c_85_n N_A_22_259#_c_86_n N_A_22_259#_c_87_n
+ N_A_22_259#_c_88_n N_A_22_259#_c_89_n N_A_22_259#_c_101_p N_A_22_259#_c_104_p
+ N_A_22_259#_c_114_p N_A_22_259#_c_80_n N_A_22_259#_c_91_n N_A_22_259#_c_81_n
+ PM_SKY130_FD_SC_LP__A21BO_2%A_22_259#
x_PM_SKY130_FD_SC_LP__A21BO_2%B1_N N_B1_N_M1002_g N_B1_N_M1004_g B1_N B1_N B1_N
+ N_B1_N_c_166_n N_B1_N_c_167_n PM_SKY130_FD_SC_LP__A21BO_2%B1_N
x_PM_SKY130_FD_SC_LP__A21BO_2%A_304_153# N_A_304_153#_M1002_d
+ N_A_304_153#_M1004_d N_A_304_153#_c_192_n N_A_304_153#_M1006_g
+ N_A_304_153#_M1010_g N_A_304_153#_c_195_n N_A_304_153#_c_196_n
+ N_A_304_153#_c_197_n N_A_304_153#_c_198_n
+ PM_SKY130_FD_SC_LP__A21BO_2%A_304_153#
x_PM_SKY130_FD_SC_LP__A21BO_2%A1 N_A1_M1011_g N_A1_M1005_g A1 A1 N_A1_c_238_n
+ N_A1_c_239_n PM_SKY130_FD_SC_LP__A21BO_2%A1
x_PM_SKY130_FD_SC_LP__A21BO_2%A2 N_A2_M1009_g N_A2_M1003_g A2 N_A2_c_272_n
+ N_A2_c_273_n PM_SKY130_FD_SC_LP__A21BO_2%A2
x_PM_SKY130_FD_SC_LP__A21BO_2%VPWR N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_M1005_d
+ N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n VPWR
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_294_n N_VPWR_c_303_n
+ N_VPWR_c_304_n PM_SKY130_FD_SC_LP__A21BO_2%VPWR
x_PM_SKY130_FD_SC_LP__A21BO_2%X N_X_M1000_s N_X_M1001_s X X X X X
+ PM_SKY130_FD_SC_LP__A21BO_2%X
x_PM_SKY130_FD_SC_LP__A21BO_2%A_508_367# N_A_508_367#_M1010_d
+ N_A_508_367#_M1003_d N_A_508_367#_c_362_n N_A_508_367#_c_358_n
+ N_A_508_367#_c_359_n N_A_508_367#_c_360_n
+ PM_SKY130_FD_SC_LP__A21BO_2%A_508_367#
x_PM_SKY130_FD_SC_LP__A21BO_2%VGND N_VGND_M1000_d N_VGND_M1008_d N_VGND_M1006_s
+ N_VGND_M1009_d N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n
+ N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n VGND N_VGND_c_388_n
+ N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n
+ PM_SKY130_FD_SC_LP__A21BO_2%VGND
cc_1 VNB N_A_22_259#_c_73_n 0.0211732f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.295
cc_2 VNB N_A_22_259#_M1001_g 0.00178952f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_3 VNB N_A_22_259#_c_75_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.37
cc_4 VNB N_A_22_259#_c_76_n 0.0184299f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.295
cc_5 VNB N_A_22_259#_M1007_g 0.0104807f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_6 VNB N_A_22_259#_c_78_n 0.00492193f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.37
cc_7 VNB N_A_22_259#_c_79_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.46
cc_8 VNB N_A_22_259#_c_80_n 0.00657399f $X=-0.19 $Y=-0.245 $X2=2.222 $Y2=1.815
cc_9 VNB N_A_22_259#_c_81_n 0.0525738f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.46
cc_10 VNB N_B1_N_M1004_g 0.00158942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B1_N 0.00802569f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.765
cc_12 VNB N_B1_N_c_166_n 0.0311062f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.37
cc_13 VNB N_B1_N_c_167_n 0.0212912f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.765
cc_14 VNB N_A_304_153#_c_192_n 0.0229486f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.295
cc_15 VNB N_A_304_153#_M1006_g 0.023941f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_16 VNB N_A_304_153#_M1010_g 0.0106133f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.37
cc_17 VNB N_A_304_153#_c_195_n 0.00391059f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.765
cc_18 VNB N_A_304_153#_c_196_n 0.0189899f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.765
cc_19 VNB N_A_304_153#_c_197_n 4.25797e-19 $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_20 VNB N_A_304_153#_c_198_n 0.0399505f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.46
cc_21 VNB N_A1_M1005_g 0.00774116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A1 0.0115786f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.765
cc_23 VNB N_A1_c_238_n 0.0300839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_239_n 0.0170382f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.37
cc_25 VNB N_A2_M1003_g 0.0116295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB A2 0.0130194f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.765
cc_27 VNB N_A2_c_272_n 0.0363285f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_28 VNB N_A2_c_273_n 0.0218156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_294_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=0.945
cc_30 VNB X 0.0066318f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.295
cc_31 VNB N_VGND_c_381_n 0.0116782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_382_n 0.0431588f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.37
cc_33 VNB N_VGND_c_383_n 0.0232831f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.445
cc_34 VNB N_VGND_c_384_n 0.0249166f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.37
cc_35 VNB N_VGND_c_385_n 0.0196257f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.46
cc_36 VNB N_VGND_c_386_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.41
cc_37 VNB N_VGND_c_387_n 0.0334596f $X=-0.19 $Y=-0.245 $X2=2.222 $Y2=1.952
cc_38 VNB N_VGND_c_388_n 0.0155275f $X=-0.19 $Y=-0.245 $X2=2.222 $Y2=2.495
cc_39 VNB N_VGND_c_389_n 0.0271101f $X=-0.19 $Y=-0.245 $X2=2.272 $Y2=1.815
cc_40 VNB N_VGND_c_390_n 0.0058666f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.46
cc_41 VNB N_VGND_c_391_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.46
cc_42 VNB N_VGND_c_392_n 0.229873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A_22_259#_M1001_g 0.0235194f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_44 VPB N_A_22_259#_M1007_g 0.0224586f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_45 VPB N_A_22_259#_c_79_n 0.0257756f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.46
cc_46 VPB N_A_22_259#_c_85_n 0.029535f $X=-0.19 $Y=1.655 $X2=2.085 $Y2=2.41
cc_47 VPB N_A_22_259#_c_86_n 0.0075223f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=2.41
cc_48 VPB N_A_22_259#_c_87_n 0.00287275f $X=-0.19 $Y=1.655 $X2=2.222 $Y2=1.952
cc_49 VPB N_A_22_259#_c_88_n 0.00449971f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=1.98
cc_50 VPB N_A_22_259#_c_89_n 0.0222208f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=2.91
cc_51 VPB N_A_22_259#_c_80_n 0.00340738f $X=-0.19 $Y=1.655 $X2=2.222 $Y2=1.815
cc_52 VPB N_A_22_259#_c_91_n 2.51509e-19 $X=-0.19 $Y=1.655 $X2=2.222 $Y2=2.41
cc_53 VPB N_B1_N_M1004_g 0.0225995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB B1_N 0.00133979f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.765
cc_55 VPB N_A_304_153#_M1010_g 0.022606f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.37
cc_56 VPB N_A_304_153#_c_197_n 0.00616266f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_57 VPB N_A1_M1005_g 0.0189925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A2_M1003_g 0.0247156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_295_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.625
cc_60 VPB N_VPWR_c_296_n 0.0195232f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_61 VPB N_VPWR_c_297_n 0.0195239f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.295
cc_62 VPB N_VPWR_c_298_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_63 VPB N_VPWR_c_299_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.46
cc_64 VPB N_VPWR_c_300_n 0.0467082f $X=-0.19 $Y=1.655 $X2=2.222 $Y2=1.952
cc_65 VPB N_VPWR_c_301_n 0.0158241f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.945
cc_66 VPB N_VPWR_c_294_n 0.0563338f $X=-0.19 $Y=1.655 $X2=2.36 $Y2=0.945
cc_67 VPB N_VPWR_c_303_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.222 $Y2=2.41
cc_68 VPB N_VPWR_c_304_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.46
cc_69 VPB X 0.00355002f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.295
cc_70 VPB N_A_508_367#_c_358_n 0.0151588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_508_367#_c_359_n 0.00224829f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.37
cc_72 VPB N_A_508_367#_c_360_n 0.0465671f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.765
cc_73 N_A_22_259#_M1007_g N_B1_N_M1004_g 0.0211544f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A_22_259#_c_85_n N_B1_N_M1004_g 0.010385f $X=2.085 $Y=2.41 $X2=0 $Y2=0
cc_75 N_A_22_259#_c_87_n N_B1_N_M1004_g 0.0042998f $X=2.222 $Y=1.952 $X2=0 $Y2=0
cc_76 N_A_22_259#_c_76_n B1_N 0.00847135f $X=0.92 $Y=1.295 $X2=0 $Y2=0
cc_77 N_A_22_259#_c_85_n B1_N 0.0254338f $X=2.085 $Y=2.41 $X2=0 $Y2=0
cc_78 N_A_22_259#_c_78_n N_B1_N_c_166_n 0.0203185f $X=0.92 $Y=1.37 $X2=0 $Y2=0
cc_79 N_A_22_259#_c_76_n N_B1_N_c_167_n 0.0114661f $X=0.92 $Y=1.295 $X2=0 $Y2=0
cc_80 N_A_22_259#_c_87_n N_A_304_153#_c_192_n 0.00329104f $X=2.222 $Y=1.952
+ $X2=0 $Y2=0
cc_81 N_A_22_259#_c_80_n N_A_304_153#_c_192_n 0.0143025f $X=2.222 $Y=1.815 $X2=0
+ $Y2=0
cc_82 N_A_22_259#_c_101_p N_A_304_153#_M1006_g 0.0151611f $X=2.585 $Y=0.945
+ $X2=0 $Y2=0
cc_83 N_A_22_259#_c_80_n N_A_304_153#_M1006_g 0.00801685f $X=2.222 $Y=1.815
+ $X2=0 $Y2=0
cc_84 N_A_22_259#_c_80_n N_A_304_153#_M1010_g 0.0106004f $X=2.222 $Y=1.815 $X2=0
+ $Y2=0
cc_85 N_A_22_259#_c_104_p N_A_304_153#_c_196_n 0.0107622f $X=2.36 $Y=0.945 $X2=0
+ $Y2=0
cc_86 N_A_22_259#_c_80_n N_A_304_153#_c_196_n 0.0455045f $X=2.222 $Y=1.815 $X2=0
+ $Y2=0
cc_87 N_A_22_259#_c_85_n N_A_304_153#_c_197_n 0.021403f $X=2.085 $Y=2.41 $X2=0
+ $Y2=0
cc_88 N_A_22_259#_c_87_n N_A_304_153#_c_197_n 0.0244313f $X=2.222 $Y=1.952 $X2=0
+ $Y2=0
cc_89 N_A_22_259#_c_80_n N_A_304_153#_c_197_n 0.00993957f $X=2.222 $Y=1.815
+ $X2=0 $Y2=0
cc_90 N_A_22_259#_c_80_n N_A_304_153#_c_198_n 0.00134666f $X=2.222 $Y=1.815
+ $X2=0 $Y2=0
cc_91 N_A_22_259#_c_101_p A1 0.0214056f $X=2.585 $Y=0.945 $X2=0 $Y2=0
cc_92 N_A_22_259#_c_80_n A1 0.0244019f $X=2.222 $Y=1.815 $X2=0 $Y2=0
cc_93 N_A_22_259#_c_101_p N_A1_c_238_n 0.00148141f $X=2.585 $Y=0.945 $X2=0 $Y2=0
cc_94 N_A_22_259#_c_101_p N_A1_c_239_n 0.00349802f $X=2.585 $Y=0.945 $X2=0 $Y2=0
cc_95 N_A_22_259#_c_114_p N_A1_c_239_n 0.0117658f $X=2.68 $Y=0.42 $X2=0 $Y2=0
cc_96 N_A_22_259#_c_101_p N_A2_c_273_n 5.39154e-19 $X=2.585 $Y=0.945 $X2=0 $Y2=0
cc_97 N_A_22_259#_c_114_p N_A2_c_273_n 0.00183298f $X=2.68 $Y=0.42 $X2=0 $Y2=0
cc_98 N_A_22_259#_c_79_n N_VPWR_M1001_d 0.00230064f $X=0.275 $Y=1.46 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_22_259#_c_86_n N_VPWR_M1001_d 0.00306947f $X=0.44 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_22_259#_c_85_n N_VPWR_M1007_d 0.00514235f $X=2.085 $Y=2.41 $X2=0
+ $Y2=0
cc_101 N_A_22_259#_M1001_g N_VPWR_c_296_n 0.014885f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_22_259#_M1007_g N_VPWR_c_296_n 0.00169308f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_A_22_259#_c_86_n N_VPWR_c_296_n 0.0237968f $X=0.44 $Y=2.41 $X2=0 $Y2=0
cc_104 N_A_22_259#_M1001_g N_VPWR_c_297_n 0.00169308f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_A_22_259#_M1007_g N_VPWR_c_297_n 0.014886f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_22_259#_c_85_n N_VPWR_c_297_n 0.0215105f $X=2.085 $Y=2.41 $X2=0 $Y2=0
cc_107 N_A_22_259#_M1001_g N_VPWR_c_299_n 0.00486043f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_22_259#_M1007_g N_VPWR_c_299_n 0.00486043f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_A_22_259#_c_89_n N_VPWR_c_300_n 0.0183433f $X=2.25 $Y=2.91 $X2=0 $Y2=0
cc_110 N_A_22_259#_M1010_s N_VPWR_c_294_n 0.00319521f $X=2.125 $Y=1.835 $X2=0
+ $Y2=0
cc_111 N_A_22_259#_M1001_g N_VPWR_c_294_n 0.00459245f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_A_22_259#_M1007_g N_VPWR_c_294_n 0.00460886f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_22_259#_c_85_n N_VPWR_c_294_n 0.0449337f $X=2.085 $Y=2.41 $X2=0 $Y2=0
cc_114 N_A_22_259#_c_86_n N_VPWR_c_294_n 0.00119414f $X=0.44 $Y=2.41 $X2=0 $Y2=0
cc_115 N_A_22_259#_c_89_n N_VPWR_c_294_n 0.0106136f $X=2.25 $Y=2.91 $X2=0 $Y2=0
cc_116 N_A_22_259#_c_85_n N_X_M1001_s 0.00508781f $X=2.085 $Y=2.41 $X2=0 $Y2=0
cc_117 N_A_22_259#_c_73_n X 0.00302902f $X=0.49 $Y=1.295 $X2=0 $Y2=0
cc_118 N_A_22_259#_c_75_n X 0.0137561f $X=0.845 $Y=1.37 $X2=0 $Y2=0
cc_119 N_A_22_259#_c_76_n X 0.00201958f $X=0.92 $Y=1.295 $X2=0 $Y2=0
cc_120 N_A_22_259#_M1007_g X 0.00340751f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_22_259#_c_79_n X 0.0468567f $X=0.275 $Y=1.46 $X2=0 $Y2=0
cc_122 N_A_22_259#_c_85_n X 0.0135055f $X=2.085 $Y=2.41 $X2=0 $Y2=0
cc_123 N_A_22_259#_c_81_n X 0.00305982f $X=0.565 $Y=1.46 $X2=0 $Y2=0
cc_124 N_A_22_259#_c_80_n N_A_508_367#_c_359_n 0.0128285f $X=2.222 $Y=1.815
+ $X2=0 $Y2=0
cc_125 N_A_22_259#_c_104_p N_VGND_M1006_s 0.0039849f $X=2.36 $Y=0.945 $X2=0
+ $Y2=0
cc_126 N_A_22_259#_c_80_n N_VGND_M1006_s 5.45101e-19 $X=2.222 $Y=1.815 $X2=0
+ $Y2=0
cc_127 N_A_22_259#_c_73_n N_VGND_c_382_n 0.0177988f $X=0.49 $Y=1.295 $X2=0 $Y2=0
cc_128 N_A_22_259#_c_76_n N_VGND_c_382_n 5.86893e-19 $X=0.92 $Y=1.295 $X2=0
+ $Y2=0
cc_129 N_A_22_259#_c_79_n N_VGND_c_382_n 0.0291318f $X=0.275 $Y=1.46 $X2=0 $Y2=0
cc_130 N_A_22_259#_c_81_n N_VGND_c_382_n 0.00779955f $X=0.565 $Y=1.46 $X2=0
+ $Y2=0
cc_131 N_A_22_259#_c_76_n N_VGND_c_383_n 0.00365171f $X=0.92 $Y=1.295 $X2=0
+ $Y2=0
cc_132 N_A_22_259#_c_101_p N_VGND_c_385_n 0.0017491f $X=2.585 $Y=0.945 $X2=0
+ $Y2=0
cc_133 N_A_22_259#_c_104_p N_VGND_c_385_n 0.0130463f $X=2.36 $Y=0.945 $X2=0
+ $Y2=0
cc_134 N_A_22_259#_c_101_p N_VGND_c_387_n 0.00454195f $X=2.585 $Y=0.945 $X2=0
+ $Y2=0
cc_135 N_A_22_259#_c_114_p N_VGND_c_387_n 0.0164453f $X=2.68 $Y=0.42 $X2=0 $Y2=0
cc_136 N_A_22_259#_c_73_n N_VGND_c_388_n 0.00400407f $X=0.49 $Y=1.295 $X2=0
+ $Y2=0
cc_137 N_A_22_259#_c_76_n N_VGND_c_388_n 0.00480781f $X=0.92 $Y=1.295 $X2=0
+ $Y2=0
cc_138 N_A_22_259#_c_114_p N_VGND_c_389_n 0.015688f $X=2.68 $Y=0.42 $X2=0 $Y2=0
cc_139 N_A_22_259#_M1006_d N_VGND_c_392_n 0.00253254f $X=2.54 $Y=0.235 $X2=0
+ $Y2=0
cc_140 N_A_22_259#_c_73_n N_VGND_c_392_n 0.00774504f $X=0.49 $Y=1.295 $X2=0
+ $Y2=0
cc_141 N_A_22_259#_c_76_n N_VGND_c_392_n 0.00971208f $X=0.92 $Y=1.295 $X2=0
+ $Y2=0
cc_142 N_A_22_259#_c_101_p N_VGND_c_392_n 0.00499226f $X=2.585 $Y=0.945 $X2=0
+ $Y2=0
cc_143 N_A_22_259#_c_104_p N_VGND_c_392_n 6.18499e-19 $X=2.36 $Y=0.945 $X2=0
+ $Y2=0
cc_144 N_A_22_259#_c_114_p N_VGND_c_392_n 0.00984745f $X=2.68 $Y=0.42 $X2=0
+ $Y2=0
cc_145 B1_N N_A_304_153#_c_196_n 0.0338405f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_146 N_B1_N_c_166_n N_A_304_153#_c_196_n 0.00225327f $X=1.37 $Y=1.46 $X2=0
+ $Y2=0
cc_147 N_B1_N_c_167_n N_A_304_153#_c_196_n 0.0115127f $X=1.372 $Y=1.295 $X2=0
+ $Y2=0
cc_148 N_B1_N_M1004_g N_A_304_153#_c_197_n 0.00602905f $X=1.465 $Y=2.045 $X2=0
+ $Y2=0
cc_149 B1_N N_A_304_153#_c_197_n 0.0384703f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_150 B1_N N_A_304_153#_c_198_n 2.81072e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_151 N_B1_N_c_166_n N_A_304_153#_c_198_n 0.0204769f $X=1.37 $Y=1.46 $X2=0
+ $Y2=0
cc_152 B1_N N_VPWR_M1007_d 0.00832999f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_153 B1_N X 0.0493412f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_154 B1_N N_VGND_c_383_n 0.0218792f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B1_N_c_166_n N_VGND_c_383_n 5.98291e-19 $X=1.37 $Y=1.46 $X2=0 $Y2=0
cc_156 N_B1_N_c_167_n N_VGND_c_383_n 0.00651792f $X=1.372 $Y=1.295 $X2=0 $Y2=0
cc_157 N_B1_N_c_167_n N_VGND_c_384_n 0.00348629f $X=1.372 $Y=1.295 $X2=0 $Y2=0
cc_158 N_B1_N_c_167_n N_VGND_c_385_n 0.001352f $X=1.372 $Y=1.295 $X2=0 $Y2=0
cc_159 N_B1_N_c_167_n N_VGND_c_392_n 0.00432409f $X=1.372 $Y=1.295 $X2=0 $Y2=0
cc_160 N_A_304_153#_M1010_g N_A1_M1005_g 0.027103f $X=2.465 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A_304_153#_M1006_g A1 0.0018808f $X=2.465 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A_304_153#_M1010_g A1 0.00137916f $X=2.465 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_304_153#_c_195_n A1 0.00369175f $X=2.465 $Y=1.37 $X2=0 $Y2=0
cc_164 N_A_304_153#_M1006_g N_A1_c_238_n 0.0213596f $X=2.465 $Y=0.655 $X2=0
+ $Y2=0
cc_165 N_A_304_153#_M1006_g N_A1_c_239_n 0.0144853f $X=2.465 $Y=0.655 $X2=0
+ $Y2=0
cc_166 N_A_304_153#_M1010_g N_VPWR_c_298_n 0.0013973f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_304_153#_M1010_g N_VPWR_c_300_n 0.00571722f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_304_153#_M1010_g N_VPWR_c_294_n 0.0117938f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_304_153#_M1010_g N_A_508_367#_c_362_n 0.0132439f $X=2.465 $Y=2.465
+ $X2=0 $Y2=0
cc_170 N_A_304_153#_M1010_g N_A_508_367#_c_359_n 0.00353967f $X=2.465 $Y=2.465
+ $X2=0 $Y2=0
cc_171 N_A_304_153#_c_196_n N_VGND_c_383_n 0.0173913f $X=1.755 $Y=1.625 $X2=0
+ $Y2=0
cc_172 N_A_304_153#_c_192_n N_VGND_c_385_n 0.00314439f $X=2.39 $Y=1.37 $X2=0
+ $Y2=0
cc_173 N_A_304_153#_M1006_g N_VGND_c_385_n 0.0132192f $X=2.465 $Y=0.655 $X2=0
+ $Y2=0
cc_174 N_A_304_153#_M1006_g N_VGND_c_389_n 0.00486043f $X=2.465 $Y=0.655 $X2=0
+ $Y2=0
cc_175 N_A_304_153#_M1006_g N_VGND_c_392_n 0.00460797f $X=2.465 $Y=0.655 $X2=0
+ $Y2=0
cc_176 N_A_304_153#_c_196_n N_VGND_c_392_n 0.0166155f $X=1.755 $Y=1.625 $X2=0
+ $Y2=0
cc_177 N_A1_M1005_g N_A2_M1003_g 0.0233828f $X=2.895 $Y=2.465 $X2=0 $Y2=0
cc_178 A1 A2 0.0252184f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A1_c_238_n A2 3.5333e-19 $X=2.915 $Y=1.35 $X2=0 $Y2=0
cc_180 A1 N_A2_c_272_n 0.00233081f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A1_c_238_n N_A2_c_272_n 0.0206091f $X=2.915 $Y=1.35 $X2=0 $Y2=0
cc_182 N_A1_c_239_n N_A2_c_273_n 0.0402464f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A1_M1005_g N_VPWR_c_298_n 0.0145911f $X=2.895 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A1_M1005_g N_VPWR_c_300_n 0.00564095f $X=2.895 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A1_M1005_g N_VPWR_c_294_n 0.00950825f $X=2.895 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A1_M1005_g N_A_508_367#_c_358_n 0.0147495f $X=2.895 $Y=2.465 $X2=0
+ $Y2=0
cc_187 A1 N_A_508_367#_c_358_n 0.0306187f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A1_c_238_n N_A_508_367#_c_358_n 0.00302458f $X=2.915 $Y=1.35 $X2=0
+ $Y2=0
cc_189 A1 N_A_508_367#_c_359_n 0.0230939f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_c_238_n N_A_508_367#_c_359_n 0.0010483f $X=2.915 $Y=1.35 $X2=0 $Y2=0
cc_191 N_A1_c_239_n N_VGND_c_385_n 0.00124028f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A1_c_239_n N_VGND_c_387_n 0.00337156f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_193 N_A1_c_239_n N_VGND_c_389_n 0.0054895f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_194 N_A1_c_239_n N_VGND_c_392_n 0.0101742f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_195 N_A2_M1003_g N_VPWR_c_298_n 0.0154114f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A2_M1003_g N_VPWR_c_301_n 0.00564095f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A2_M1003_g N_VPWR_c_294_n 0.0104155f $X=3.365 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A2_M1003_g N_A_508_367#_c_358_n 0.0189143f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_199 A2 N_A_508_367#_c_358_n 0.0245287f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A2_c_272_n N_A_508_367#_c_358_n 0.00451858f $X=3.47 $Y=1.35 $X2=0 $Y2=0
cc_201 A2 N_VGND_c_387_n 0.0197533f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_202 N_A2_c_272_n N_VGND_c_387_n 0.00436897f $X=3.47 $Y=1.35 $X2=0 $Y2=0
cc_203 N_A2_c_273_n N_VGND_c_387_n 0.0237311f $X=3.462 $Y=1.185 $X2=0 $Y2=0
cc_204 N_A2_c_273_n N_VGND_c_389_n 0.00486043f $X=3.462 $Y=1.185 $X2=0 $Y2=0
cc_205 N_A2_c_273_n N_VGND_c_392_n 0.00848326f $X=3.462 $Y=1.185 $X2=0 $Y2=0
cc_206 N_VPWR_c_294_n N_X_M1001_s 0.00408795f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_c_294_n N_A_508_367#_M1010_d 0.00310528f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_208 N_VPWR_c_294_n N_A_508_367#_M1003_d 0.00302127f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_300_n N_A_508_367#_c_362_n 0.0153751f $X=2.965 $Y=3.33 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_294_n N_A_508_367#_c_362_n 0.0101105f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_M1005_d N_A_508_367#_c_358_n 0.00218982f $X=2.97 $Y=1.835 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_298_n N_A_508_367#_c_358_n 0.017285f $X=3.13 $Y=2.11 $X2=0 $Y2=0
cc_213 N_VPWR_c_301_n N_A_508_367#_c_360_n 0.0185207f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_294_n N_A_508_367#_c_360_n 0.010808f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_215 X N_VGND_c_382_n 0.0345013f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_216 X N_VGND_c_383_n 0.0300941f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_217 X N_VGND_c_388_n 0.010561f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_218 X N_VGND_c_392_n 0.00798307f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_219 N_A_508_367#_c_358_n N_VGND_c_387_n 0.00206951f $X=3.465 $Y=1.77 $X2=0
+ $Y2=0
cc_220 N_VGND_c_392_n A_594_47# 0.0137053f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
