* File: sky130_fd_sc_lp__o31ai_4.spice
* Created: Fri Aug 28 11:16:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31ai_4.pex.spice"
.subckt sky130_fd_sc_lp__o31ai_4  VNB VPB A2 A1 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_132_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75007.2 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A1_M1010_g N_A_132_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75006.7 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1010_d N_A1_M1016_g N_A_132_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75006.3 A=0.126 P=1.98 MULT=1
MM1027 N_VGND_M1027_d N_A1_M1027_g N_A_132_47#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75005.9 A=0.126 P=1.98 MULT=1
MM1029 N_VGND_M1027_d N_A1_M1029_g N_A_132_47#_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75005.4 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_132_47#_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3 SB=75005
+ A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1007_d N_A2_M1011_g N_A_132_47#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75004.6 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_A2_M1024_g N_A_132_47#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1005 N_A_132_47#_M1005_d N_A3_M1005_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1017 N_A_132_47#_M1005_d N_A3_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=6.42 M=1 R=5.6 SA=75004.1
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1019 N_A_132_47#_M1019_d N_A3_M1019_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=3.564 M=1 R=5.6 SA=75004.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1008 N_A_132_47#_M1019_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005 SB=75002.4
+ A=0.126 P=1.98 MULT=1
MM1014 N_A_132_47#_M1014_d N_B1_M1014_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.4
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1023 N_A_132_47#_M1014_d N_B1_M1023_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.273 PD=1.12 PS=1.49 NRD=0 NRS=0 M=1 R=5.6 SA=75005.8 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1025 N_A_132_47#_M1025_d N_B1_M1025_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.273 PD=1.12 PS=1.49 NRD=0 NRS=0 M=1 R=5.6 SA=75006.6 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1022 N_A_132_47#_M1025_d N_A3_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2898 PD=1.12 PS=2.37 NRD=0 NRS=11.424 M=1 R=5.6 SA=75007.1
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1012 N_A_132_367#_M1012_d N_A2_M1012_g N_A_49_367#_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75007.3 A=0.189 P=2.82 MULT=1
MM1001 N_A_132_367#_M1012_d N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.9 A=0.189 P=2.82 MULT=1
MM1009 N_A_132_367#_M1009_d N_A1_M1009_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75006.4 A=0.189 P=2.82 MULT=1
MM1013 N_A_132_367#_M1009_d N_A1_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75006 A=0.189 P=2.82 MULT=1
MM1026 N_A_132_367#_M1026_d N_A1_M1026_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1020 N_A_132_367#_M1026_d N_A2_M1020_g N_A_49_367#_M1020_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1030 N_A_132_367#_M1030_d N_A2_M1030_g N_A_49_367#_M1020_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1031 N_A_132_367#_M1030_d N_A2_M1031_g N_A_49_367#_M1031_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A3_M1006_g N_A_49_367#_M1031_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75003.8 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1006_d N_A3_M1015_g N_A_49_367#_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1018 N_Y_M1018_d N_A3_M1018_g N_A_49_367#_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5 SB=75003
+ A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_Y_M1018_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3465 AS=0.1764 PD=1.81 PS=1.54 NRD=42.1974 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1000_d N_B1_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3465 AS=0.1764 PD=1.81 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3213 AS=0.1764 PD=1.77 PS=1.54 NRD=9.3772 NRS=0 M=1 R=8.4 SA=75006.1
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1003_d N_B1_M1021_g N_Y_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3213 AS=0.2394 PD=1.77 PS=1.64 NRD=26.5753 NRS=15.6221 M=1 R=8.4
+ SA=75006.7 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1028 N_Y_M1021_s N_A3_M1028_g N_A_49_367#_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2394 AS=0.3906 PD=1.64 PS=3.14 NRD=0 NRS=7.0329 M=1 R=8.4 SA=75007.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.9271 P=20.81
*
.include "sky130_fd_sc_lp__o31ai_4.pxi.spice"
*
.ends
*
*
