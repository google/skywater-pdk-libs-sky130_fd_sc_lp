* File: sky130_fd_sc_lp__o32a_lp.spice
* Created: Fri Aug 28 11:17:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o32a_lp  VNB VPB B1 B2 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_A_134_101#_M1000_d N_B1_M1000_g N_A_31_101#_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.08085 AS=0.1533 PD=0.84 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75000.3 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_31_101#_M1009_d N_B2_M1009_g N_A_134_101#_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.08085 PD=0.7 PS=0.84 NRD=0 NRS=24.276 M=1 R=2.8
+ SA=75000.7 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A3_M1010_g N_A_31_101#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.136625 AS=0.0588 PD=1.165 PS=0.7 NRD=77.22 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1001 N_A_31_101#_M1001_d N_A2_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.136625 PD=0.7 PS=1.165 NRD=0 NRS=77.22 M=1 R=2.8 SA=75001.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A1_M1003_g N_A_31_101#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1008 A_612_89# N_A_134_101#_M1008_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_X_M1011_d N_A_134_101#_M1011_g A_612_89# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_151_419# N_B1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.3 PD=1.24 PS=2.6 NRD=12.7853 NRS=2.9353 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1007 N_A_134_101#_M1007_d N_B2_M1007_g A_151_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.1925 AS=0.12 PD=1.385 PS=1.24 NRD=20.685 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1004 A_376_419# N_A3_M1004_g N_A_134_101#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.1925 PD=1.24 PS=1.385 NRD=12.7853 NRS=0 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1012 A_474_419# N_A2_M1012_g A_376_419# VPB PHIGHVT L=0.25 W=1 AD=0.12 AS=0.12
+ PD=1.24 PS=1.24 NRD=12.7853 NRS=12.7853 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g A_474_419# VPB PHIGHVT L=0.25 W=1 AD=0.145
+ AS=0.12 PD=1.29 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_X_M1006_d N_A_134_101#_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.145 PD=2.57 PS=1.29 NRD=0 NRS=1.9503 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o32a_lp.pxi.spice"
*
.ends
*
*
