* File: sky130_fd_sc_lp__o2111ai_4.pxi.spice
* Created: Fri Aug 28 11:01:11 2020
* 
x_PM_SKY130_FD_SC_LP__O2111AI_4%D1 N_D1_M1010_g N_D1_M1000_g N_D1_M1017_g
+ N_D1_M1011_g N_D1_M1019_g N_D1_M1024_g N_D1_M1037_g N_D1_M1036_g N_D1_c_160_n
+ N_D1_c_175_p N_D1_c_161_n D1 N_D1_c_162_n PM_SKY130_FD_SC_LP__O2111AI_4%D1
x_PM_SKY130_FD_SC_LP__O2111AI_4%C1 N_C1_M1007_g N_C1_M1004_g N_C1_M1013_g
+ N_C1_M1009_g N_C1_M1029_g N_C1_M1025_g N_C1_M1031_g N_C1_M1030_g N_C1_c_236_n
+ N_C1_c_237_n C1 N_C1_c_238_n N_C1_c_239_n PM_SKY130_FD_SC_LP__O2111AI_4%C1
x_PM_SKY130_FD_SC_LP__O2111AI_4%B1 N_B1_c_320_n N_B1_M1002_g N_B1_c_314_n
+ N_B1_M1001_g N_B1_c_321_n N_B1_M1005_g N_B1_c_315_n N_B1_M1016_g N_B1_c_322_n
+ N_B1_M1014_g N_B1_c_316_n N_B1_M1022_g N_B1_c_323_n N_B1_M1032_g N_B1_c_317_n
+ N_B1_M1033_g B1 B1 B1 B1 N_B1_c_319_n PM_SKY130_FD_SC_LP__O2111AI_4%B1
x_PM_SKY130_FD_SC_LP__O2111AI_4%A2 N_A2_c_407_n N_A2_M1003_g N_A2_M1008_g
+ N_A2_c_408_n N_A2_M1015_g N_A2_M1020_g N_A2_c_409_n N_A2_M1026_g N_A2_M1021_g
+ N_A2_c_410_n N_A2_M1027_g N_A2_M1038_g N_A2_c_403_n N_A2_c_404_n A2
+ N_A2_c_406_n PM_SKY130_FD_SC_LP__O2111AI_4%A2
x_PM_SKY130_FD_SC_LP__O2111AI_4%A1 N_A1_M1006_g N_A1_M1018_g N_A1_M1012_g
+ N_A1_M1034_g N_A1_M1023_g N_A1_M1035_g N_A1_M1028_g N_A1_M1039_g A1 A1 A1 A1
+ N_A1_c_507_n N_A1_c_508_n PM_SKY130_FD_SC_LP__O2111AI_4%A1
x_PM_SKY130_FD_SC_LP__O2111AI_4%Y N_Y_M1010_d N_Y_M1019_d N_Y_M1000_s
+ N_Y_M1011_s N_Y_M1036_s N_Y_M1009_s N_Y_M1030_s N_Y_M1005_s N_Y_M1032_s
+ N_Y_M1015_s N_Y_M1027_s N_Y_c_580_n N_Y_c_584_n N_Y_c_602_n N_Y_c_679_p
+ N_Y_c_585_n N_Y_c_680_p N_Y_c_586_n N_Y_c_675_p N_Y_c_587_n N_Y_c_588_n
+ N_Y_c_681_p N_Y_c_636_n N_Y_c_682_p N_Y_c_640_n N_Y_c_684_p N_Y_c_648_n
+ N_Y_c_705_p N_Y_c_589_n N_Y_c_581_n N_Y_c_582_n N_Y_c_590_n N_Y_c_591_n
+ N_Y_c_592_n N_Y_c_644_n N_Y_c_646_n N_Y_c_593_n N_Y_c_594_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__O2111AI_4%Y
x_PM_SKY130_FD_SC_LP__O2111AI_4%VPWR N_VPWR_M1000_d N_VPWR_M1024_d
+ N_VPWR_M1004_d N_VPWR_M1025_d N_VPWR_M1002_d N_VPWR_M1014_d N_VPWR_M1006_s
+ N_VPWR_M1012_s N_VPWR_M1028_s N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_729_n
+ N_VPWR_c_730_n N_VPWR_c_731_n N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n
+ N_VPWR_c_735_n N_VPWR_c_736_n N_VPWR_c_737_n N_VPWR_c_738_n N_VPWR_c_739_n
+ N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_744_n
+ N_VPWR_c_745_n VPWR N_VPWR_c_746_n N_VPWR_c_747_n N_VPWR_c_748_n
+ N_VPWR_c_749_n N_VPWR_c_750_n N_VPWR_c_751_n N_VPWR_c_752_n N_VPWR_c_753_n
+ N_VPWR_c_726_n PM_SKY130_FD_SC_LP__O2111AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O2111AI_4%A_1210_367# N_A_1210_367#_M1003_d
+ N_A_1210_367#_M1026_d N_A_1210_367#_M1006_d N_A_1210_367#_M1023_d
+ N_A_1210_367#_c_883_n N_A_1210_367#_c_886_n N_A_1210_367#_c_889_n
+ N_A_1210_367#_c_891_n N_A_1210_367#_c_893_n N_A_1210_367#_c_882_n
+ N_A_1210_367#_c_901_n N_A_1210_367#_c_904_n N_A_1210_367#_c_937_n
+ N_A_1210_367#_c_905_n N_A_1210_367#_c_909_n N_A_1210_367#_c_941_n
+ N_A_1210_367#_c_897_n N_A_1210_367#_c_911_n
+ PM_SKY130_FD_SC_LP__O2111AI_4%A_1210_367#
x_PM_SKY130_FD_SC_LP__O2111AI_4%A_27_47# N_A_27_47#_M1010_s N_A_27_47#_M1017_s
+ N_A_27_47#_M1037_s N_A_27_47#_M1013_d N_A_27_47#_M1031_d N_A_27_47#_c_948_n
+ N_A_27_47#_c_991_p N_A_27_47#_c_944_n N_A_27_47#_c_945_n N_A_27_47#_c_961_n
+ N_A_27_47#_c_946_n N_A_27_47#_c_947_n PM_SKY130_FD_SC_LP__O2111AI_4%A_27_47#
x_PM_SKY130_FD_SC_LP__O2111AI_4%A_454_47# N_A_454_47#_M1007_s
+ N_A_454_47#_M1029_s N_A_454_47#_M1001_s N_A_454_47#_M1022_s
+ N_A_454_47#_c_1001_n N_A_454_47#_c_1009_n N_A_454_47#_c_1005_n
+ N_A_454_47#_c_1011_n N_A_454_47#_c_1014_n
+ PM_SKY130_FD_SC_LP__O2111AI_4%A_454_47#
x_PM_SKY130_FD_SC_LP__O2111AI_4%A_819_47# N_A_819_47#_M1001_d
+ N_A_819_47#_M1016_d N_A_819_47#_M1033_d N_A_819_47#_M1020_s
+ N_A_819_47#_M1038_s N_A_819_47#_M1034_d N_A_819_47#_M1039_d
+ N_A_819_47#_c_1050_n N_A_819_47#_c_1051_n N_A_819_47#_c_1052_n
+ N_A_819_47#_c_1115_n N_A_819_47#_c_1053_n N_A_819_47#_c_1127_p
+ N_A_819_47#_c_1054_n N_A_819_47#_c_1128_p N_A_819_47#_c_1080_n
+ N_A_819_47#_c_1129_p N_A_819_47#_c_1055_n N_A_819_47#_c_1130_p
+ N_A_819_47#_c_1056_n N_A_819_47#_c_1057_n N_A_819_47#_c_1074_n
+ N_A_819_47#_c_1058_n N_A_819_47#_c_1059_n N_A_819_47#_c_1060_n
+ N_A_819_47#_c_1061_n PM_SKY130_FD_SC_LP__O2111AI_4%A_819_47#
x_PM_SKY130_FD_SC_LP__O2111AI_4%VGND N_VGND_M1008_d N_VGND_M1021_d
+ N_VGND_M1018_s N_VGND_M1035_s N_VGND_c_1145_n N_VGND_c_1146_n N_VGND_c_1147_n
+ N_VGND_c_1148_n N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n
+ N_VGND_c_1152_n VGND N_VGND_c_1153_n N_VGND_c_1154_n N_VGND_c_1155_n
+ N_VGND_c_1156_n N_VGND_c_1157_n N_VGND_c_1158_n
+ PM_SKY130_FD_SC_LP__O2111AI_4%VGND
cc_1 VNB N_D1_M1010_g 0.0232583f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_D1_M1000_g 0.00376879f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_D1_M1017_g 0.0194968f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_4 VNB N_D1_M1011_g 0.0035059f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_5 VNB N_D1_M1019_g 0.0193142f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_6 VNB N_D1_M1024_g 0.00350909f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_7 VNB N_D1_M1037_g 0.0200765f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_8 VNB N_D1_M1036_g 0.00362641f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_9 VNB N_D1_c_160_n 0.00108573f $X=-0.19 $Y=-0.245 $X2=1.097 $Y2=1.352
cc_10 VNB N_D1_c_161_n 0.00576019f $X=-0.19 $Y=-0.245 $X2=1.533 $Y2=1.352
cc_11 VNB N_D1_c_162_n 0.0813648f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.42
cc_12 VNB N_C1_M1007_g 0.0192874f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_13 VNB N_C1_M1004_g 0.00362641f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_14 VNB N_C1_M1013_g 0.0190206f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_15 VNB N_C1_M1009_g 0.00350909f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_16 VNB N_C1_M1029_g 0.0193127f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_17 VNB N_C1_M1025_g 0.00350909f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_18 VNB N_C1_M1031_g 0.0232284f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_19 VNB N_C1_M1030_g 0.00397811f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_20 VNB N_C1_c_236_n 0.00148829f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.42
cc_21 VNB N_C1_c_237_n 0.0012052f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.42
cc_22 VNB N_C1_c_238_n 0.094921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_c_239_n 0.00630066f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.352
cc_24 VNB N_B1_c_314_n 0.0195571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_315_n 0.0152515f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_26 VNB N_B1_c_316_n 0.0152515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_c_317_n 0.0153124f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_28 VNB B1 0.00769054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_c_319_n 0.124321f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.42
cc_30 VNB N_A2_M1008_g 0.0198242f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_31 VNB N_A2_M1020_g 0.0196263f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.585
cc_32 VNB N_A2_M1021_g 0.0200724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_M1038_g 0.0236041f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_34 VNB N_A2_c_403_n 0.00220488f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.42
cc_35 VNB N_A2_c_404_n 0.00140207f $X=-0.19 $Y=-0.245 $X2=1.097 $Y2=1.352
cc_36 VNB A2 0.00734935f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.352
cc_37 VNB N_A2_c_406_n 0.0930819f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.42
cc_38 VNB N_A1_M1006_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_39 VNB N_A1_M1018_g 0.0245523f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_40 VNB N_A1_M1012_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_41 VNB N_A1_M1034_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_42 VNB N_A1_M1023_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_43 VNB N_A1_M1035_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_44 VNB N_A1_M1028_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_45 VNB N_A1_M1039_g 0.0284365f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_46 VNB A1 0.0160169f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.42
cc_47 VNB N_A1_c_507_n 0.0931637f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.42
cc_48 VNB N_A1_c_508_n 0.0438136f $X=-0.19 $Y=-0.245 $X2=1.533 $Y2=1.352
cc_49 VNB N_Y_c_580_n 0.00827133f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.42
cc_50 VNB N_Y_c_581_n 9.80655e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Y_c_582_n 0.00220865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB Y 0.0254479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VPWR_c_726_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_27_47#_c_944_n 0.00314562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_47#_c_945_n 0.00421655f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.255
cc_56 VNB N_A_27_47#_c_946_n 0.0223254f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_57 VNB N_A_27_47#_c_947_n 0.00238485f $X=-0.19 $Y=-0.245 $X2=1.097 $Y2=1.352
cc_58 VNB N_A_454_47#_c_1001_n 0.0128051f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.585
cc_59 VNB N_A_819_47#_c_1050_n 0.00393389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_819_47#_c_1051_n 0.0028872f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_61 VNB N_A_819_47#_c_1052_n 0.00294003f $X=-0.19 $Y=-0.245 $X2=1.765
+ $Y2=0.655
cc_62 VNB N_A_819_47#_c_1053_n 0.00414532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_819_47#_c_1054_n 0.00312279f $X=-0.19 $Y=-0.245 $X2=1.097
+ $Y2=1.352
cc_64 VNB N_A_819_47#_c_1055_n 0.00306842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_819_47#_c_1056_n 0.0122038f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.42
cc_66 VNB N_A_819_47#_c_1057_n 0.0284746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_819_47#_c_1058_n 0.00389908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_819_47#_c_1059_n 0.00204151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_819_47#_c_1060_n 0.0066849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_819_47#_c_1061_n 0.00152782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1145_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_72 VNB N_VGND_c_1146_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_73 VNB N_VGND_c_1147_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_74 VNB N_VGND_c_1148_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_75 VNB N_VGND_c_1149_n 0.144354f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_76 VNB N_VGND_c_1150_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_77 VNB N_VGND_c_1151_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.42
cc_78 VNB N_VGND_c_1152_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.42
cc_79 VNB N_VGND_c_1153_n 0.021009f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_80 VNB N_VGND_c_1154_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.42
cc_81 VNB N_VGND_c_1155_n 0.0179216f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.352
cc_82 VNB N_VGND_c_1156_n 0.474328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1157_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1158_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VPB N_D1_M1000_g 0.0233761f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_86 VPB N_D1_M1011_g 0.0182267f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_87 VPB N_D1_M1024_g 0.0182451f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_88 VPB N_D1_M1036_g 0.0183453f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_89 VPB N_C1_M1004_g 0.0183453f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_90 VPB N_C1_M1009_g 0.0182451f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_91 VPB N_C1_M1025_g 0.0182451f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_92 VPB N_C1_M1030_g 0.0209836f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_93 VPB N_B1_c_320_n 0.0180799f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.255
cc_94 VPB N_B1_c_321_n 0.0157077f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_95 VPB N_B1_c_322_n 0.0157609f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.585
cc_96 VPB N_B1_c_323_n 0.016015f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.655
cc_97 VPB B1 0.0124989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_B1_c_319_n 0.035562f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=1.42
cc_99 VPB N_A2_c_407_n 0.0164331f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.255
cc_100 VPB N_A2_c_408_n 0.0161699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A2_c_409_n 0.0152515f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_102 VPB N_A2_c_410_n 0.0195571f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_103 VPB N_A2_c_406_n 0.0227211f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.42
cc_104 VPB N_A1_M1006_g 0.0231352f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_105 VPB N_A1_M1012_g 0.0187475f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.655
cc_106 VPB N_A1_M1023_g 0.0187475f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.655
cc_107 VPB N_A1_M1028_g 0.0245754f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.655
cc_108 VPB A1 0.0250591f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.42
cc_109 VPB N_Y_c_584_n 0.00320975f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.42
cc_110 VPB N_Y_c_585_n 0.00297559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_Y_c_586_n 0.00297836f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.42
cc_112 VPB N_Y_c_587_n 0.00289786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_Y_c_588_n 0.00288394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_Y_c_589_n 2.17744e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_Y_c_590_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_Y_c_591_n 0.00288887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_Y_c_592_n 0.00143206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_Y_c_593_n 0.00121151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_Y_c_594_n 0.00918573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB Y 9.67293e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB Y 0.00774107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB Y 0.0472745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_727_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_124 VPB N_VPWR_c_728_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.42
cc_125 VPB N_VPWR_c_729_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.352
cc_126 VPB N_VPWR_c_730_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.71 $Y2=1.42
cc_127 VPB N_VPWR_c_731_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_732_n 3.99158e-19 $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.42
cc_129 VPB N_VPWR_c_733_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_734_n 0.00886878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_735_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_736_n 0.0135296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_737_n 0.0478673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_738_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_739_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_740_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_741_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_742_n 0.0204486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_743_n 0.00443527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_744_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_745_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_746_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_747_n 0.0598893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_748_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_749_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_750_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_751_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_752_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_753_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_726_n 0.0524506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_1210_367#_c_882_n 0.0142745f $X=-0.19 $Y=1.655 $X2=1.765
+ $Y2=0.655
cc_152 N_D1_M1037_g N_C1_M1007_g 0.0179875f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_153 N_D1_M1036_g N_C1_M1004_g 0.0235071f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_154 N_D1_c_161_n N_C1_c_237_n 0.0124388f $X=1.533 $Y=1.352 $X2=0 $Y2=0
cc_155 N_D1_c_162_n N_C1_c_237_n 2.50256e-19 $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_156 N_D1_c_161_n N_C1_c_238_n 5.79489e-19 $X=1.533 $Y=1.352 $X2=0 $Y2=0
cc_157 N_D1_c_162_n N_C1_c_238_n 0.0239944f $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_158 N_D1_M1000_g N_Y_c_584_n 0.0168597f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_159 N_D1_M1011_g N_Y_c_584_n 0.0141753f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_160 N_D1_c_175_p N_Y_c_584_n 0.0352929f $X=0.945 $Y=1.352 $X2=0 $Y2=0
cc_161 N_D1_c_162_n N_Y_c_584_n 0.00246472f $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_162 N_D1_M1017_g N_Y_c_602_n 0.0132113f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_163 N_D1_M1019_g N_Y_c_602_n 0.0126234f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_164 N_D1_c_160_n N_Y_c_602_n 0.0395646f $X=1.097 $Y=1.352 $X2=0 $Y2=0
cc_165 N_D1_c_175_p N_Y_c_602_n 0.00626862f $X=0.945 $Y=1.352 $X2=0 $Y2=0
cc_166 N_D1_c_161_n N_Y_c_602_n 0.010314f $X=1.533 $Y=1.352 $X2=0 $Y2=0
cc_167 N_D1_c_162_n N_Y_c_602_n 0.00130915f $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_168 N_D1_M1024_g N_Y_c_585_n 0.0141753f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_169 N_D1_M1036_g N_Y_c_585_n 0.0141253f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_170 N_D1_c_161_n N_Y_c_585_n 0.0476355f $X=1.533 $Y=1.352 $X2=0 $Y2=0
cc_171 N_D1_c_162_n N_Y_c_585_n 0.00332595f $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_172 N_D1_M1010_g N_Y_c_581_n 0.0133008f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_173 N_D1_c_175_p N_Y_c_581_n 0.018047f $X=0.945 $Y=1.352 $X2=0 $Y2=0
cc_174 N_D1_M1017_g N_Y_c_582_n 0.002515f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_175 N_D1_c_162_n N_Y_c_582_n 0.00251669f $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_176 N_D1_c_160_n N_Y_c_590_n 0.015901f $X=1.097 $Y=1.352 $X2=0 $Y2=0
cc_177 N_D1_c_162_n N_Y_c_590_n 0.00256759f $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_178 N_D1_M1010_g Y 0.0193028f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_179 N_D1_c_160_n Y 0.00424439f $X=1.097 $Y=1.352 $X2=0 $Y2=0
cc_180 N_D1_c_175_p Y 0.0138858f $X=0.945 $Y=1.352 $X2=0 $Y2=0
cc_181 N_D1_M1000_g N_VPWR_c_727_n 0.0178941f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_182 N_D1_M1011_g N_VPWR_c_727_n 0.01587f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_183 N_D1_M1024_g N_VPWR_c_727_n 7.49804e-19 $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_184 N_D1_M1011_g N_VPWR_c_728_n 7.49804e-19 $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_185 N_D1_M1024_g N_VPWR_c_728_n 0.01587f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_186 N_D1_M1036_g N_VPWR_c_728_n 0.01587f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_187 N_D1_M1036_g N_VPWR_c_729_n 7.49804e-19 $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_188 N_D1_M1011_g N_VPWR_c_738_n 0.00486043f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_189 N_D1_M1024_g N_VPWR_c_738_n 0.00486043f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_190 N_D1_M1036_g N_VPWR_c_740_n 0.00486043f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_191 N_D1_M1000_g N_VPWR_c_746_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_192 N_D1_M1000_g N_VPWR_c_726_n 0.00917987f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_193 N_D1_M1011_g N_VPWR_c_726_n 0.00824727f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_194 N_D1_M1024_g N_VPWR_c_726_n 0.00824727f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_195 N_D1_M1036_g N_VPWR_c_726_n 0.0082726f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_196 N_D1_M1010_g N_A_27_47#_c_948_n 0.0114156f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_197 N_D1_M1017_g N_A_27_47#_c_948_n 0.0104569f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_198 N_D1_M1019_g N_A_27_47#_c_948_n 0.0103812f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_199 N_D1_M1037_g N_A_27_47#_c_948_n 0.0153414f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_200 N_D1_M1037_g N_A_27_47#_c_945_n 0.00263136f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_201 N_D1_c_161_n N_A_27_47#_c_945_n 0.00155335f $X=1.533 $Y=1.352 $X2=0 $Y2=0
cc_202 N_D1_c_162_n N_A_27_47#_c_945_n 5.10663e-19 $X=1.765 $Y=1.42 $X2=0 $Y2=0
cc_203 N_D1_M1010_g N_A_27_47#_c_946_n 0.00623683f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_204 N_D1_M1017_g N_A_27_47#_c_946_n 8.9618e-19 $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_205 N_D1_M1010_g N_VGND_c_1149_n 0.00359361f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_206 N_D1_M1017_g N_VGND_c_1149_n 0.00357877f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_207 N_D1_M1019_g N_VGND_c_1149_n 0.00357877f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_208 N_D1_M1037_g N_VGND_c_1149_n 0.00357877f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_209 N_D1_M1010_g N_VGND_c_1156_n 0.0062747f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_210 N_D1_M1017_g N_VGND_c_1156_n 0.0053512f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_211 N_D1_M1019_g N_VGND_c_1156_n 0.0053512f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_212 N_D1_M1037_g N_VGND_c_1156_n 0.00537654f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_213 N_C1_M1030_g N_B1_c_320_n 0.00477805f $X=3.485 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_214 N_C1_M1030_g B1 0.002238f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_215 N_C1_c_238_n B1 0.00283248f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_216 N_C1_c_239_n B1 0.0131949f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_217 N_C1_M1031_g N_B1_c_319_n 0.00169371f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_218 N_C1_M1030_g N_B1_c_319_n 0.00341277f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_219 N_C1_c_238_n N_B1_c_319_n 0.0206043f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_220 N_C1_c_239_n N_B1_c_319_n 0.00295192f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_221 N_C1_M1004_g N_Y_c_586_n 0.0141315f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_222 N_C1_M1009_g N_Y_c_586_n 0.0141753f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_223 N_C1_c_237_n N_Y_c_586_n 0.0462455f $X=3.115 $Y=1.33 $X2=0 $Y2=0
cc_224 N_C1_c_238_n N_Y_c_586_n 0.00332737f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_225 N_C1_M1025_g N_Y_c_587_n 0.0141287f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_226 N_C1_M1030_g N_Y_c_587_n 0.0146409f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_227 N_C1_c_237_n N_Y_c_587_n 0.0486534f $X=3.115 $Y=1.33 $X2=0 $Y2=0
cc_228 N_C1_c_238_n N_Y_c_587_n 0.00357126f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_229 N_C1_c_238_n N_Y_c_588_n 0.0043649f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_230 N_C1_c_239_n N_Y_c_588_n 0.014393f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_231 N_C1_c_237_n N_Y_c_592_n 0.015388f $X=3.115 $Y=1.33 $X2=0 $Y2=0
cc_232 N_C1_c_238_n N_Y_c_592_n 0.00256759f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_233 N_C1_M1004_g N_VPWR_c_728_n 7.49804e-19 $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_234 N_C1_M1004_g N_VPWR_c_729_n 0.01587f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_235 N_C1_M1009_g N_VPWR_c_729_n 0.01587f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_236 N_C1_M1025_g N_VPWR_c_729_n 7.49804e-19 $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_237 N_C1_M1009_g N_VPWR_c_730_n 0.00486043f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_238 N_C1_M1025_g N_VPWR_c_730_n 0.00486043f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_239 N_C1_M1009_g N_VPWR_c_731_n 7.49804e-19 $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_240 N_C1_M1025_g N_VPWR_c_731_n 0.01587f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_241 N_C1_M1030_g N_VPWR_c_731_n 0.0178919f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_242 N_C1_M1004_g N_VPWR_c_740_n 0.00486043f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_243 N_C1_M1030_g N_VPWR_c_742_n 0.00486043f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_244 N_C1_M1004_g N_VPWR_c_726_n 0.0082726f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_245 N_C1_M1009_g N_VPWR_c_726_n 0.00824727f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_246 N_C1_M1025_g N_VPWR_c_726_n 0.00824727f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_247 N_C1_M1030_g N_VPWR_c_726_n 0.00888845f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_248 N_C1_M1007_g N_A_27_47#_c_944_n 0.0129997f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_249 N_C1_M1013_g N_A_27_47#_c_944_n 0.0103943f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_250 N_C1_c_237_n N_A_27_47#_c_944_n 0.0462833f $X=3.115 $Y=1.33 $X2=0 $Y2=0
cc_251 N_C1_c_238_n N_A_27_47#_c_944_n 0.00328782f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_252 N_C1_M1029_g N_A_27_47#_c_961_n 0.0134748f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_253 N_C1_M1031_g N_A_27_47#_c_961_n 0.0126055f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_254 N_C1_c_236_n N_A_27_47#_c_961_n 0.0461463f $X=3.29 $Y=1.33 $X2=0 $Y2=0
cc_255 N_C1_c_237_n N_A_27_47#_c_961_n 0.00619999f $X=3.115 $Y=1.33 $X2=0 $Y2=0
cc_256 N_C1_c_238_n N_A_27_47#_c_961_n 0.00170609f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_257 N_C1_M1013_g N_A_27_47#_c_947_n 3.04429e-19 $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_258 N_C1_M1029_g N_A_27_47#_c_947_n 0.00226238f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_259 N_C1_c_237_n N_A_27_47#_c_947_n 0.0156189f $X=3.115 $Y=1.33 $X2=0 $Y2=0
cc_260 N_C1_c_238_n N_A_27_47#_c_947_n 0.00250816f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_261 N_C1_M1013_g N_A_454_47#_c_1001_n 0.0109459f $X=2.625 $Y=0.655 $X2=0
+ $Y2=0
cc_262 N_C1_M1029_g N_A_454_47#_c_1001_n 0.00927192f $X=3.055 $Y=0.655 $X2=0
+ $Y2=0
cc_263 N_C1_M1031_g N_A_454_47#_c_1001_n 0.0120412f $X=3.485 $Y=0.655 $X2=0
+ $Y2=0
cc_264 N_C1_M1007_g N_A_454_47#_c_1005_n 0.00616418f $X=2.195 $Y=0.655 $X2=0
+ $Y2=0
cc_265 N_C1_M1013_g N_A_454_47#_c_1005_n 0.00644475f $X=2.625 $Y=0.655 $X2=0
+ $Y2=0
cc_266 N_C1_M1029_g N_A_454_47#_c_1005_n 8.73235e-19 $X=3.055 $Y=0.655 $X2=0
+ $Y2=0
cc_267 N_C1_M1031_g N_A_819_47#_c_1052_n 0.00426638f $X=3.485 $Y=0.655 $X2=0
+ $Y2=0
cc_268 N_C1_c_239_n N_A_819_47#_c_1052_n 0.00191044f $X=3.61 $Y=1.42 $X2=0 $Y2=0
cc_269 N_C1_M1007_g N_VGND_c_1149_n 0.0054895f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_270 N_C1_M1013_g N_VGND_c_1149_n 0.00359361f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_271 N_C1_M1029_g N_VGND_c_1149_n 0.00357877f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_272 N_C1_M1031_g N_VGND_c_1149_n 0.00357877f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_273 N_C1_M1007_g N_VGND_c_1156_n 0.0099382f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_274 N_C1_M1013_g N_VGND_c_1156_n 0.00534209f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_275 N_C1_M1029_g N_VGND_c_1156_n 0.0053512f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_276 N_C1_M1031_g N_VGND_c_1156_n 0.00675087f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_277 N_B1_c_323_n N_A2_c_407_n 0.00926302f $X=5.545 $Y=1.725 $X2=-0.19
+ $Y2=-0.245
cc_278 N_B1_c_317_n N_A2_M1008_g 0.0208211f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_279 B1 N_A2_c_404_n 0.00842596f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_280 N_B1_c_319_n N_A2_c_404_n 2.10899e-19 $X=5.545 $Y=1.457 $X2=0 $Y2=0
cc_281 B1 N_A2_c_406_n 0.00333597f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_282 N_B1_c_319_n N_A2_c_406_n 0.0302869f $X=5.545 $Y=1.457 $X2=0 $Y2=0
cc_283 N_B1_c_320_n N_Y_c_588_n 0.0034916f $X=4.255 $Y=1.73 $X2=0 $Y2=0
cc_284 B1 N_Y_c_588_n 0.0228692f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_285 N_B1_c_319_n N_Y_c_588_n 0.00119825f $X=5.545 $Y=1.457 $X2=0 $Y2=0
cc_286 N_B1_c_320_n N_Y_c_636_n 0.0124077f $X=4.255 $Y=1.73 $X2=0 $Y2=0
cc_287 N_B1_c_321_n N_Y_c_636_n 0.0125619f $X=4.685 $Y=1.725 $X2=0 $Y2=0
cc_288 B1 N_Y_c_636_n 0.0438829f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_289 N_B1_c_319_n N_Y_c_636_n 0.00147362f $X=5.545 $Y=1.457 $X2=0 $Y2=0
cc_290 N_B1_c_322_n N_Y_c_640_n 0.0125619f $X=5.115 $Y=1.725 $X2=0 $Y2=0
cc_291 N_B1_c_323_n N_Y_c_640_n 0.0125619f $X=5.545 $Y=1.725 $X2=0 $Y2=0
cc_292 B1 N_Y_c_640_n 0.043669f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_293 N_B1_c_319_n N_Y_c_640_n 6.51543e-19 $X=5.545 $Y=1.457 $X2=0 $Y2=0
cc_294 B1 N_Y_c_644_n 0.0156128f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_295 N_B1_c_319_n N_Y_c_644_n 7.31333e-19 $X=5.545 $Y=1.457 $X2=0 $Y2=0
cc_296 B1 N_Y_c_646_n 0.00121827f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_297 N_B1_c_319_n N_Y_c_646_n 0.00371162f $X=5.545 $Y=1.457 $X2=0 $Y2=0
cc_298 N_B1_c_320_n N_VPWR_c_732_n 0.0168789f $X=4.255 $Y=1.73 $X2=0 $Y2=0
cc_299 N_B1_c_321_n N_VPWR_c_732_n 0.0144971f $X=4.685 $Y=1.725 $X2=0 $Y2=0
cc_300 N_B1_c_322_n N_VPWR_c_732_n 6.7792e-19 $X=5.115 $Y=1.725 $X2=0 $Y2=0
cc_301 N_B1_c_321_n N_VPWR_c_733_n 6.77662e-19 $X=4.685 $Y=1.725 $X2=0 $Y2=0
cc_302 N_B1_c_322_n N_VPWR_c_733_n 0.0144971f $X=5.115 $Y=1.725 $X2=0 $Y2=0
cc_303 N_B1_c_323_n N_VPWR_c_733_n 0.0156897f $X=5.545 $Y=1.725 $X2=0 $Y2=0
cc_304 N_B1_c_320_n N_VPWR_c_742_n 0.0046653f $X=4.255 $Y=1.73 $X2=0 $Y2=0
cc_305 N_B1_c_321_n N_VPWR_c_744_n 0.00486043f $X=4.685 $Y=1.725 $X2=0 $Y2=0
cc_306 N_B1_c_322_n N_VPWR_c_744_n 0.00486043f $X=5.115 $Y=1.725 $X2=0 $Y2=0
cc_307 N_B1_c_323_n N_VPWR_c_747_n 0.00486043f $X=5.545 $Y=1.725 $X2=0 $Y2=0
cc_308 N_B1_c_320_n N_VPWR_c_726_n 0.00857954f $X=4.255 $Y=1.73 $X2=0 $Y2=0
cc_309 N_B1_c_321_n N_VPWR_c_726_n 0.00824727f $X=4.685 $Y=1.725 $X2=0 $Y2=0
cc_310 N_B1_c_322_n N_VPWR_c_726_n 0.00824727f $X=5.115 $Y=1.725 $X2=0 $Y2=0
cc_311 N_B1_c_323_n N_VPWR_c_726_n 0.0082726f $X=5.545 $Y=1.725 $X2=0 $Y2=0
cc_312 N_B1_c_314_n N_A_454_47#_c_1001_n 0.012436f $X=4.435 $Y=1.185 $X2=0 $Y2=0
cc_313 N_B1_c_315_n N_A_454_47#_c_1009_n 0.0083908f $X=4.865 $Y=1.185 $X2=0
+ $Y2=0
cc_314 N_B1_c_316_n N_A_454_47#_c_1009_n 0.0083908f $X=5.295 $Y=1.185 $X2=0
+ $Y2=0
cc_315 N_B1_c_314_n N_A_454_47#_c_1011_n 0.0103967f $X=4.435 $Y=1.185 $X2=0
+ $Y2=0
cc_316 N_B1_c_315_n N_A_454_47#_c_1011_n 0.00639056f $X=4.865 $Y=1.185 $X2=0
+ $Y2=0
cc_317 N_B1_c_316_n N_A_454_47#_c_1011_n 3.28947e-19 $X=5.295 $Y=1.185 $X2=0
+ $Y2=0
cc_318 N_B1_c_315_n N_A_454_47#_c_1014_n 5.05504e-19 $X=4.865 $Y=1.185 $X2=0
+ $Y2=0
cc_319 N_B1_c_316_n N_A_454_47#_c_1014_n 0.00638651f $X=5.295 $Y=1.185 $X2=0
+ $Y2=0
cc_320 N_B1_c_317_n N_A_454_47#_c_1014_n 0.00648785f $X=5.725 $Y=1.185 $X2=0
+ $Y2=0
cc_321 N_B1_c_314_n N_A_819_47#_c_1051_n 0.0133491f $X=4.435 $Y=1.185 $X2=0
+ $Y2=0
cc_322 N_B1_c_315_n N_A_819_47#_c_1051_n 0.0121487f $X=4.865 $Y=1.185 $X2=0
+ $Y2=0
cc_323 B1 N_A_819_47#_c_1051_n 0.0498596f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_324 N_B1_c_319_n N_A_819_47#_c_1051_n 0.00459926f $X=5.545 $Y=1.457 $X2=0
+ $Y2=0
cc_325 B1 N_A_819_47#_c_1052_n 0.0206234f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_326 N_B1_c_319_n N_A_819_47#_c_1052_n 0.00840772f $X=5.545 $Y=1.457 $X2=0
+ $Y2=0
cc_327 N_B1_c_316_n N_A_819_47#_c_1053_n 0.0121487f $X=5.295 $Y=1.185 $X2=0
+ $Y2=0
cc_328 N_B1_c_317_n N_A_819_47#_c_1053_n 0.0163862f $X=5.725 $Y=1.185 $X2=0
+ $Y2=0
cc_329 B1 N_A_819_47#_c_1053_n 0.0381358f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_330 N_B1_c_319_n N_A_819_47#_c_1053_n 0.00322408f $X=5.545 $Y=1.457 $X2=0
+ $Y2=0
cc_331 B1 N_A_819_47#_c_1074_n 0.0151973f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_332 N_B1_c_319_n N_A_819_47#_c_1074_n 0.00502918f $X=5.545 $Y=1.457 $X2=0
+ $Y2=0
cc_333 N_B1_c_317_n N_VGND_c_1145_n 0.00125916f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_334 N_B1_c_314_n N_VGND_c_1149_n 0.00357842f $X=4.435 $Y=1.185 $X2=0 $Y2=0
cc_335 N_B1_c_315_n N_VGND_c_1149_n 0.00357842f $X=4.865 $Y=1.185 $X2=0 $Y2=0
cc_336 N_B1_c_316_n N_VGND_c_1149_n 0.00357842f $X=5.295 $Y=1.185 $X2=0 $Y2=0
cc_337 N_B1_c_317_n N_VGND_c_1149_n 0.00547432f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_338 N_B1_c_314_n N_VGND_c_1156_n 0.00675085f $X=4.435 $Y=1.185 $X2=0 $Y2=0
cc_339 N_B1_c_315_n N_VGND_c_1156_n 0.00535118f $X=4.865 $Y=1.185 $X2=0 $Y2=0
cc_340 N_B1_c_316_n N_VGND_c_1156_n 0.00535118f $X=5.295 $Y=1.185 $X2=0 $Y2=0
cc_341 N_B1_c_317_n N_VGND_c_1156_n 0.00990114f $X=5.725 $Y=1.185 $X2=0 $Y2=0
cc_342 N_A2_M1038_g N_A1_M1018_g 0.00644846f $X=7.445 $Y=0.655 $X2=0 $Y2=0
cc_343 A2 N_A1_M1018_g 0.00176393f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_344 A2 A1 0.00958593f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_345 N_A2_c_406_n A1 0.00358544f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_346 A2 N_A1_c_507_n 0.00283805f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_347 N_A2_c_406_n N_A1_c_507_n 0.00903732f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_348 N_A2_c_407_n N_Y_c_648_n 0.0157803f $X=5.975 $Y=1.725 $X2=0 $Y2=0
cc_349 N_A2_c_408_n N_Y_c_648_n 0.0137639f $X=6.405 $Y=1.725 $X2=0 $Y2=0
cc_350 N_A2_c_404_n N_Y_c_648_n 0.0151383f $X=7.135 $Y=1.365 $X2=0 $Y2=0
cc_351 N_A2_c_406_n N_Y_c_648_n 0.0028017f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_352 N_A2_c_409_n N_Y_c_589_n 0.0101867f $X=6.835 $Y=1.725 $X2=0 $Y2=0
cc_353 N_A2_c_410_n N_Y_c_589_n 0.00685606f $X=7.265 $Y=1.725 $X2=0 $Y2=0
cc_354 N_A2_c_404_n N_Y_c_589_n 0.0393724f $X=7.135 $Y=1.365 $X2=0 $Y2=0
cc_355 N_A2_c_406_n N_Y_c_589_n 0.0113715f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_356 N_A2_c_408_n N_Y_c_593_n 0.00278291f $X=6.405 $Y=1.725 $X2=0 $Y2=0
cc_357 N_A2_c_409_n N_Y_c_593_n 2.3962e-19 $X=6.835 $Y=1.725 $X2=0 $Y2=0
cc_358 N_A2_c_404_n N_Y_c_593_n 0.0147221f $X=7.135 $Y=1.365 $X2=0 $Y2=0
cc_359 N_A2_c_406_n N_Y_c_593_n 0.0068357f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_360 N_A2_c_409_n N_Y_c_594_n 5.20508e-19 $X=6.835 $Y=1.725 $X2=0 $Y2=0
cc_361 N_A2_c_410_n N_Y_c_594_n 0.00756873f $X=7.265 $Y=1.725 $X2=0 $Y2=0
cc_362 A2 N_Y_c_594_n 0.0259658f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_363 N_A2_c_406_n N_Y_c_594_n 0.00615858f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_364 N_A2_c_407_n N_VPWR_c_733_n 0.00131998f $X=5.975 $Y=1.725 $X2=0 $Y2=0
cc_365 N_A2_c_410_n N_VPWR_c_734_n 0.00924783f $X=7.265 $Y=1.725 $X2=0 $Y2=0
cc_366 N_A2_c_407_n N_VPWR_c_747_n 0.00547432f $X=5.975 $Y=1.725 $X2=0 $Y2=0
cc_367 N_A2_c_408_n N_VPWR_c_747_n 0.00357842f $X=6.405 $Y=1.725 $X2=0 $Y2=0
cc_368 N_A2_c_409_n N_VPWR_c_747_n 0.00357842f $X=6.835 $Y=1.725 $X2=0 $Y2=0
cc_369 N_A2_c_410_n N_VPWR_c_747_n 0.00547432f $X=7.265 $Y=1.725 $X2=0 $Y2=0
cc_370 N_A2_c_407_n N_VPWR_c_726_n 0.00990114f $X=5.975 $Y=1.725 $X2=0 $Y2=0
cc_371 N_A2_c_408_n N_VPWR_c_726_n 0.00535118f $X=6.405 $Y=1.725 $X2=0 $Y2=0
cc_372 N_A2_c_409_n N_VPWR_c_726_n 0.00535118f $X=6.835 $Y=1.725 $X2=0 $Y2=0
cc_373 N_A2_c_410_n N_VPWR_c_726_n 0.0076668f $X=7.265 $Y=1.725 $X2=0 $Y2=0
cc_374 N_A2_c_407_n N_A_1210_367#_c_883_n 0.00844452f $X=5.975 $Y=1.725 $X2=0
+ $Y2=0
cc_375 N_A2_c_408_n N_A_1210_367#_c_883_n 0.00968553f $X=6.405 $Y=1.725 $X2=0
+ $Y2=0
cc_376 N_A2_c_409_n N_A_1210_367#_c_883_n 5.63573e-19 $X=6.835 $Y=1.725 $X2=0
+ $Y2=0
cc_377 N_A2_c_408_n N_A_1210_367#_c_886_n 0.0107932f $X=6.405 $Y=1.725 $X2=0
+ $Y2=0
cc_378 N_A2_c_409_n N_A_1210_367#_c_886_n 0.0114056f $X=6.835 $Y=1.725 $X2=0
+ $Y2=0
cc_379 N_A2_c_410_n N_A_1210_367#_c_886_n 0.00405982f $X=7.265 $Y=1.725 $X2=0
+ $Y2=0
cc_380 N_A2_c_407_n N_A_1210_367#_c_889_n 0.00203265f $X=5.975 $Y=1.725 $X2=0
+ $Y2=0
cc_381 N_A2_c_408_n N_A_1210_367#_c_889_n 6.12373e-19 $X=6.405 $Y=1.725 $X2=0
+ $Y2=0
cc_382 N_A2_c_409_n N_A_1210_367#_c_891_n 0.00315264f $X=6.835 $Y=1.725 $X2=0
+ $Y2=0
cc_383 N_A2_c_406_n N_A_1210_367#_c_891_n 5.4695e-19 $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_384 N_A2_c_408_n N_A_1210_367#_c_893_n 4.99636e-19 $X=6.405 $Y=1.725 $X2=0
+ $Y2=0
cc_385 N_A2_c_409_n N_A_1210_367#_c_893_n 0.00526271f $X=6.835 $Y=1.725 $X2=0
+ $Y2=0
cc_386 N_A2_c_410_n N_A_1210_367#_c_893_n 0.0122164f $X=7.265 $Y=1.725 $X2=0
+ $Y2=0
cc_387 N_A2_c_410_n N_A_1210_367#_c_882_n 0.0115971f $X=7.265 $Y=1.725 $X2=0
+ $Y2=0
cc_388 N_A2_c_409_n N_A_1210_367#_c_897_n 0.00172556f $X=6.835 $Y=1.725 $X2=0
+ $Y2=0
cc_389 N_A2_c_410_n N_A_1210_367#_c_897_n 9.80814e-19 $X=7.265 $Y=1.725 $X2=0
+ $Y2=0
cc_390 N_A2_M1008_g N_A_819_47#_c_1054_n 0.0134969f $X=6.155 $Y=0.655 $X2=0
+ $Y2=0
cc_391 N_A2_M1020_g N_A_819_47#_c_1054_n 0.0127457f $X=6.585 $Y=0.655 $X2=0
+ $Y2=0
cc_392 N_A2_c_404_n N_A_819_47#_c_1054_n 0.0467631f $X=7.135 $Y=1.365 $X2=0
+ $Y2=0
cc_393 N_A2_c_406_n N_A_819_47#_c_1054_n 0.00419449f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_394 N_A2_M1021_g N_A_819_47#_c_1080_n 0.0121162f $X=7.015 $Y=0.655 $X2=0
+ $Y2=0
cc_395 N_A2_M1038_g N_A_819_47#_c_1080_n 0.0122595f $X=7.445 $Y=0.655 $X2=0
+ $Y2=0
cc_396 N_A2_c_403_n N_A_819_47#_c_1080_n 0.0282422f $X=7.295 $Y=1.365 $X2=0
+ $Y2=0
cc_397 N_A2_c_404_n N_A_819_47#_c_1080_n 0.00600522f $X=7.135 $Y=1.365 $X2=0
+ $Y2=0
cc_398 N_A2_c_406_n N_A_819_47#_c_1080_n 5.77739e-19 $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_399 N_A2_c_404_n N_A_819_47#_c_1058_n 0.00201686f $X=7.135 $Y=1.365 $X2=0
+ $Y2=0
cc_400 N_A2_c_406_n N_A_819_47#_c_1058_n 0.00496491f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_401 N_A2_M1020_g N_A_819_47#_c_1059_n 2.39715e-19 $X=6.585 $Y=0.655 $X2=0
+ $Y2=0
cc_402 N_A2_M1021_g N_A_819_47#_c_1059_n 0.00551859f $X=7.015 $Y=0.655 $X2=0
+ $Y2=0
cc_403 N_A2_M1038_g N_A_819_47#_c_1059_n 8.15368e-19 $X=7.445 $Y=0.655 $X2=0
+ $Y2=0
cc_404 N_A2_c_404_n N_A_819_47#_c_1059_n 0.0203755f $X=7.135 $Y=1.365 $X2=0
+ $Y2=0
cc_405 N_A2_c_406_n N_A_819_47#_c_1059_n 0.00299787f $X=7.265 $Y=1.5 $X2=0 $Y2=0
cc_406 N_A2_M1038_g N_A_819_47#_c_1060_n 0.00341839f $X=7.445 $Y=0.655 $X2=0
+ $Y2=0
cc_407 A2 N_A_819_47#_c_1060_n 0.00811108f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_408 N_A2_M1008_g N_VGND_c_1145_n 0.0114707f $X=6.155 $Y=0.655 $X2=0 $Y2=0
cc_409 N_A2_M1020_g N_VGND_c_1145_n 0.010278f $X=6.585 $Y=0.655 $X2=0 $Y2=0
cc_410 N_A2_M1021_g N_VGND_c_1145_n 6.16837e-19 $X=7.015 $Y=0.655 $X2=0 $Y2=0
cc_411 N_A2_M1020_g N_VGND_c_1146_n 5.74401e-19 $X=6.585 $Y=0.655 $X2=0 $Y2=0
cc_412 N_A2_M1021_g N_VGND_c_1146_n 0.0105198f $X=7.015 $Y=0.655 $X2=0 $Y2=0
cc_413 N_A2_M1038_g N_VGND_c_1146_n 0.0122042f $X=7.445 $Y=0.655 $X2=0 $Y2=0
cc_414 N_A2_M1008_g N_VGND_c_1149_n 0.00486043f $X=6.155 $Y=0.655 $X2=0 $Y2=0
cc_415 N_A2_M1020_g N_VGND_c_1151_n 0.00486043f $X=6.585 $Y=0.655 $X2=0 $Y2=0
cc_416 N_A2_M1021_g N_VGND_c_1151_n 0.00486043f $X=7.015 $Y=0.655 $X2=0 $Y2=0
cc_417 N_A2_M1038_g N_VGND_c_1153_n 0.00486043f $X=7.445 $Y=0.655 $X2=0 $Y2=0
cc_418 N_A2_M1008_g N_VGND_c_1156_n 0.0082726f $X=6.155 $Y=0.655 $X2=0 $Y2=0
cc_419 N_A2_M1020_g N_VGND_c_1156_n 0.00824727f $X=6.585 $Y=0.655 $X2=0 $Y2=0
cc_420 N_A2_M1021_g N_VGND_c_1156_n 0.0075745f $X=7.015 $Y=0.655 $X2=0 $Y2=0
cc_421 N_A2_M1038_g N_VGND_c_1156_n 0.00891413f $X=7.445 $Y=0.655 $X2=0 $Y2=0
cc_422 N_A1_M1006_g N_Y_c_594_n 0.00846192f $X=8.215 $Y=2.465 $X2=0 $Y2=0
cc_423 A1 N_Y_c_594_n 0.00337196f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_424 N_A1_M1006_g N_VPWR_c_734_n 0.0115711f $X=8.215 $Y=2.465 $X2=0 $Y2=0
cc_425 N_A1_M1012_g N_VPWR_c_734_n 5.65914e-19 $X=8.645 $Y=2.465 $X2=0 $Y2=0
cc_426 N_A1_M1006_g N_VPWR_c_735_n 6.14008e-19 $X=8.215 $Y=2.465 $X2=0 $Y2=0
cc_427 N_A1_M1012_g N_VPWR_c_735_n 0.0145375f $X=8.645 $Y=2.465 $X2=0 $Y2=0
cc_428 N_A1_M1023_g N_VPWR_c_735_n 0.0145573f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_429 N_A1_M1028_g N_VPWR_c_735_n 6.77662e-19 $X=9.505 $Y=2.465 $X2=0 $Y2=0
cc_430 N_A1_M1023_g N_VPWR_c_737_n 7.26038e-19 $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A1_M1028_g N_VPWR_c_737_n 0.0200737f $X=9.505 $Y=2.465 $X2=0 $Y2=0
cc_432 A1 N_VPWR_c_737_n 0.0260594f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_433 N_A1_c_507_n N_VPWR_c_737_n 0.00159727f $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_434 N_A1_M1006_g N_VPWR_c_748_n 0.00486043f $X=8.215 $Y=2.465 $X2=0 $Y2=0
cc_435 N_A1_M1012_g N_VPWR_c_748_n 0.00486043f $X=8.645 $Y=2.465 $X2=0 $Y2=0
cc_436 N_A1_M1023_g N_VPWR_c_749_n 0.00486043f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_437 N_A1_M1028_g N_VPWR_c_749_n 0.00486043f $X=9.505 $Y=2.465 $X2=0 $Y2=0
cc_438 N_A1_M1006_g N_VPWR_c_726_n 0.0045304f $X=8.215 $Y=2.465 $X2=0 $Y2=0
cc_439 N_A1_M1012_g N_VPWR_c_726_n 0.00824727f $X=8.645 $Y=2.465 $X2=0 $Y2=0
cc_440 N_A1_M1023_g N_VPWR_c_726_n 0.00824727f $X=9.075 $Y=2.465 $X2=0 $Y2=0
cc_441 N_A1_M1028_g N_VPWR_c_726_n 0.00824727f $X=9.505 $Y=2.465 $X2=0 $Y2=0
cc_442 N_A1_M1006_g N_A_1210_367#_c_882_n 0.0120104f $X=8.215 $Y=2.465 $X2=0
+ $Y2=0
cc_443 A1 N_A_1210_367#_c_882_n 0.00967954f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_444 N_A1_M1006_g N_A_1210_367#_c_901_n 0.00398525f $X=8.215 $Y=2.465 $X2=0
+ $Y2=0
cc_445 A1 N_A_1210_367#_c_901_n 0.019455f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_446 N_A1_c_507_n N_A_1210_367#_c_901_n 5.69681e-19 $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_447 N_A1_M1006_g N_A_1210_367#_c_904_n 0.00856708f $X=8.215 $Y=2.465 $X2=0
+ $Y2=0
cc_448 N_A1_M1012_g N_A_1210_367#_c_905_n 0.0122129f $X=8.645 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A1_M1023_g N_A_1210_367#_c_905_n 0.0122595f $X=9.075 $Y=2.465 $X2=0
+ $Y2=0
cc_450 A1 N_A_1210_367#_c_905_n 0.0434214f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_451 N_A1_c_507_n N_A_1210_367#_c_905_n 5.03185e-19 $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_452 A1 N_A_1210_367#_c_909_n 0.0155814f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_453 N_A1_c_507_n N_A_1210_367#_c_909_n 5.69681e-19 $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_454 N_A1_M1006_g N_A_1210_367#_c_911_n 0.0010444f $X=8.215 $Y=2.465 $X2=0
+ $Y2=0
cc_455 N_A1_M1018_g N_A_819_47#_c_1055_n 0.0140976f $X=8.235 $Y=0.655 $X2=0
+ $Y2=0
cc_456 N_A1_M1034_g N_A_819_47#_c_1055_n 0.0136347f $X=8.665 $Y=0.655 $X2=0
+ $Y2=0
cc_457 A1 N_A_819_47#_c_1055_n 0.0438847f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_458 N_A1_c_507_n N_A_819_47#_c_1055_n 0.00366825f $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_459 N_A1_M1035_g N_A_819_47#_c_1056_n 0.0136347f $X=9.095 $Y=0.655 $X2=0
+ $Y2=0
cc_460 N_A1_M1039_g N_A_819_47#_c_1056_n 0.0144441f $X=9.525 $Y=0.655 $X2=0
+ $Y2=0
cc_461 A1 N_A_819_47#_c_1056_n 0.0634623f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_462 N_A1_c_507_n N_A_819_47#_c_1056_n 0.00250022f $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_463 N_A1_c_508_n N_A_819_47#_c_1056_n 0.0076395f $X=9.79 $Y=1.46 $X2=0 $Y2=0
cc_464 A1 N_A_819_47#_c_1060_n 0.0143313f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_465 N_A1_c_507_n N_A_819_47#_c_1060_n 0.00480554f $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_466 A1 N_A_819_47#_c_1061_n 0.0143344f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_467 N_A1_c_507_n N_A_819_47#_c_1061_n 0.00261251f $X=9.6 $Y=1.46 $X2=0 $Y2=0
cc_468 N_A1_M1018_g N_VGND_c_1147_n 0.0119381f $X=8.235 $Y=0.655 $X2=0 $Y2=0
cc_469 N_A1_M1034_g N_VGND_c_1147_n 0.010177f $X=8.665 $Y=0.655 $X2=0 $Y2=0
cc_470 N_A1_M1035_g N_VGND_c_1147_n 6.14008e-19 $X=9.095 $Y=0.655 $X2=0 $Y2=0
cc_471 N_A1_M1034_g N_VGND_c_1148_n 6.14008e-19 $X=8.665 $Y=0.655 $X2=0 $Y2=0
cc_472 N_A1_M1035_g N_VGND_c_1148_n 0.010177f $X=9.095 $Y=0.655 $X2=0 $Y2=0
cc_473 N_A1_M1039_g N_VGND_c_1148_n 0.0119381f $X=9.525 $Y=0.655 $X2=0 $Y2=0
cc_474 N_A1_M1018_g N_VGND_c_1153_n 0.00486043f $X=8.235 $Y=0.655 $X2=0 $Y2=0
cc_475 N_A1_M1034_g N_VGND_c_1154_n 0.00486043f $X=8.665 $Y=0.655 $X2=0 $Y2=0
cc_476 N_A1_M1035_g N_VGND_c_1154_n 0.00486043f $X=9.095 $Y=0.655 $X2=0 $Y2=0
cc_477 N_A1_M1039_g N_VGND_c_1155_n 0.00486043f $X=9.525 $Y=0.655 $X2=0 $Y2=0
cc_478 N_A1_M1018_g N_VGND_c_1156_n 0.00891413f $X=8.235 $Y=0.655 $X2=0 $Y2=0
cc_479 N_A1_M1034_g N_VGND_c_1156_n 0.00824727f $X=8.665 $Y=0.655 $X2=0 $Y2=0
cc_480 N_A1_M1035_g N_VGND_c_1156_n 0.00824727f $X=9.095 $Y=0.655 $X2=0 $Y2=0
cc_481 N_A1_M1039_g N_VGND_c_1156_n 0.00924722f $X=9.525 $Y=0.655 $X2=0 $Y2=0
cc_482 N_Y_c_584_n N_VPWR_M1000_d 0.00176461f $X=1.025 $Y=1.76 $X2=-0.19
+ $Y2=-0.245
cc_483 N_Y_c_585_n N_VPWR_M1024_d 0.00176461f $X=1.885 $Y=1.76 $X2=0 $Y2=0
cc_484 N_Y_c_586_n N_VPWR_M1004_d 0.00176461f $X=2.745 $Y=1.76 $X2=0 $Y2=0
cc_485 N_Y_c_587_n N_VPWR_M1025_d 0.00176461f $X=3.605 $Y=1.76 $X2=0 $Y2=0
cc_486 N_Y_c_636_n N_VPWR_M1002_d 0.00317167f $X=4.805 $Y=2.01 $X2=0 $Y2=0
cc_487 N_Y_c_640_n N_VPWR_M1014_d 0.00331802f $X=5.665 $Y=2.01 $X2=0 $Y2=0
cc_488 N_Y_c_584_n N_VPWR_c_727_n 0.0170777f $X=1.025 $Y=1.76 $X2=0 $Y2=0
cc_489 N_Y_c_585_n N_VPWR_c_728_n 0.0170777f $X=1.885 $Y=1.76 $X2=0 $Y2=0
cc_490 N_Y_c_586_n N_VPWR_c_729_n 0.0170777f $X=2.745 $Y=1.76 $X2=0 $Y2=0
cc_491 N_Y_c_675_p N_VPWR_c_730_n 0.0124525f $X=2.84 $Y=1.98 $X2=0 $Y2=0
cc_492 N_Y_c_587_n N_VPWR_c_731_n 0.0170777f $X=3.605 $Y=1.76 $X2=0 $Y2=0
cc_493 N_Y_c_636_n N_VPWR_c_732_n 0.0175267f $X=4.805 $Y=2.01 $X2=0 $Y2=0
cc_494 N_Y_c_640_n N_VPWR_c_733_n 0.0171443f $X=5.665 $Y=2.01 $X2=0 $Y2=0
cc_495 N_Y_c_679_p N_VPWR_c_738_n 0.0124525f $X=1.12 $Y=1.98 $X2=0 $Y2=0
cc_496 N_Y_c_680_p N_VPWR_c_740_n 0.0124525f $X=1.98 $Y=1.98 $X2=0 $Y2=0
cc_497 N_Y_c_681_p N_VPWR_c_742_n 0.0361813f $X=3.7 $Y=2.91 $X2=0 $Y2=0
cc_498 N_Y_c_682_p N_VPWR_c_744_n 0.0124525f $X=4.9 $Y=2.505 $X2=0 $Y2=0
cc_499 Y N_VPWR_c_746_n 0.018528f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_500 N_Y_c_684_p N_VPWR_c_747_n 0.0124525f $X=5.76 $Y=2.505 $X2=0 $Y2=0
cc_501 N_Y_M1000_s N_VPWR_c_726_n 0.00371702f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_502 N_Y_M1011_s N_VPWR_c_726_n 0.00536646f $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_503 N_Y_M1036_s N_VPWR_c_726_n 0.00536646f $X=1.84 $Y=1.835 $X2=0 $Y2=0
cc_504 N_Y_M1009_s N_VPWR_c_726_n 0.00536646f $X=2.7 $Y=1.835 $X2=0 $Y2=0
cc_505 N_Y_M1030_s N_VPWR_c_726_n 0.00836199f $X=3.56 $Y=1.835 $X2=0 $Y2=0
cc_506 N_Y_M1005_s N_VPWR_c_726_n 0.00536646f $X=4.76 $Y=1.835 $X2=0 $Y2=0
cc_507 N_Y_M1032_s N_VPWR_c_726_n 0.00536646f $X=5.62 $Y=1.835 $X2=0 $Y2=0
cc_508 N_Y_M1015_s N_VPWR_c_726_n 0.00225186f $X=6.48 $Y=1.835 $X2=0 $Y2=0
cc_509 N_Y_M1027_s N_VPWR_c_726_n 0.00389753f $X=7.34 $Y=1.835 $X2=0 $Y2=0
cc_510 N_Y_c_679_p N_VPWR_c_726_n 0.00730901f $X=1.12 $Y=1.98 $X2=0 $Y2=0
cc_511 N_Y_c_680_p N_VPWR_c_726_n 0.00730901f $X=1.98 $Y=1.98 $X2=0 $Y2=0
cc_512 N_Y_c_675_p N_VPWR_c_726_n 0.00730901f $X=2.84 $Y=1.98 $X2=0 $Y2=0
cc_513 N_Y_c_681_p N_VPWR_c_726_n 0.020333f $X=3.7 $Y=2.91 $X2=0 $Y2=0
cc_514 N_Y_c_682_p N_VPWR_c_726_n 0.00730901f $X=4.9 $Y=2.505 $X2=0 $Y2=0
cc_515 N_Y_c_684_p N_VPWR_c_726_n 0.00730901f $X=5.76 $Y=2.505 $X2=0 $Y2=0
cc_516 Y N_VPWR_c_726_n 0.0104192f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_517 N_Y_c_648_n N_A_1210_367#_M1003_d 0.00402329f $X=6.51 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_518 N_Y_c_589_n N_A_1210_367#_M1026_d 0.00176461f $X=7.315 $Y=1.79 $X2=0
+ $Y2=0
cc_519 N_Y_c_648_n N_A_1210_367#_c_883_n 0.0171443f $X=6.51 $Y=2.01 $X2=0 $Y2=0
cc_520 N_Y_M1015_s N_A_1210_367#_c_886_n 0.00332931f $X=6.48 $Y=1.835 $X2=0
+ $Y2=0
cc_521 N_Y_c_705_p N_A_1210_367#_c_886_n 0.0127141f $X=6.62 $Y=2.56 $X2=0 $Y2=0
cc_522 N_Y_c_589_n N_A_1210_367#_c_891_n 0.0152916f $X=7.315 $Y=1.79 $X2=0 $Y2=0
cc_523 N_Y_M1027_s N_A_1210_367#_c_882_n 0.00716549f $X=7.34 $Y=1.835 $X2=0
+ $Y2=0
cc_524 N_Y_c_589_n N_A_1210_367#_c_882_n 0.00306481f $X=7.315 $Y=1.79 $X2=0
+ $Y2=0
cc_525 N_Y_c_594_n N_A_1210_367#_c_882_n 0.0212796f $X=7.48 $Y=1.79 $X2=0 $Y2=0
cc_526 N_Y_c_594_n N_A_1210_367#_c_901_n 0.00531282f $X=7.48 $Y=1.79 $X2=0 $Y2=0
cc_527 N_Y_c_594_n N_A_1210_367#_c_904_n 0.0015961f $X=7.48 $Y=1.79 $X2=0 $Y2=0
cc_528 N_Y_c_589_n N_A_1210_367#_c_897_n 8.43884e-19 $X=7.315 $Y=1.79 $X2=0
+ $Y2=0
cc_529 N_Y_c_580_n N_A_27_47#_M1010_s 0.00272521f $X=0.355 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_530 N_Y_c_602_n N_A_27_47#_M1017_s 0.00334339f $X=1.55 $Y=0.865 $X2=0 $Y2=0
cc_531 N_Y_M1010_d N_A_27_47#_c_948_n 0.00337742f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_532 N_Y_M1019_d N_A_27_47#_c_948_n 0.00337742f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_533 N_Y_c_581_n N_A_27_47#_c_948_n 0.00394508f $X=0.595 $Y=0.927 $X2=0 $Y2=0
cc_534 N_Y_c_582_n N_A_27_47#_c_948_n 0.0591745f $X=0.775 $Y=0.927 $X2=0 $Y2=0
cc_535 N_Y_c_586_n N_A_27_47#_c_944_n 3.12508e-19 $X=2.745 $Y=1.76 $X2=0 $Y2=0
cc_536 N_Y_c_585_n N_A_27_47#_c_945_n 3.70992e-19 $X=1.885 $Y=1.76 $X2=0 $Y2=0
cc_537 N_Y_c_591_n N_A_27_47#_c_945_n 0.00816307f $X=1.98 $Y=1.76 $X2=0 $Y2=0
cc_538 N_Y_c_580_n N_A_27_47#_c_946_n 0.0220891f $X=0.355 $Y=1.07 $X2=0 $Y2=0
cc_539 N_Y_c_581_n N_A_27_47#_c_946_n 0.00175788f $X=0.595 $Y=0.927 $X2=0 $Y2=0
cc_540 N_Y_M1010_d N_VGND_c_1156_n 0.00225186f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_541 N_Y_M1019_d N_VGND_c_1156_n 0.00225186f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_542 N_VPWR_c_726_n N_A_1210_367#_M1003_d 0.00223559f $X=9.84 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_543 N_VPWR_c_726_n N_A_1210_367#_M1026_d 0.00223559f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_726_n N_A_1210_367#_M1006_d 0.00408089f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_726_n N_A_1210_367#_M1023_d 0.00536646f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_734_n N_A_1210_367#_c_886_n 0.00562533f $X=8 $Y=2.8 $X2=0 $Y2=0
cc_547 N_VPWR_c_747_n N_A_1210_367#_c_886_n 0.049025f $X=7.835 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_726_n N_A_1210_367#_c_886_n 0.0312604f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_747_n N_A_1210_367#_c_889_n 0.01906f $X=7.835 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_726_n N_A_1210_367#_c_889_n 0.0124545f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_734_n N_A_1210_367#_c_893_n 0.00681933f $X=8 $Y=2.8 $X2=0 $Y2=0
cc_552 N_VPWR_M1006_s N_A_1210_367#_c_882_n 0.00792481f $X=7.875 $Y=1.835 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_734_n N_A_1210_367#_c_882_n 0.0215105f $X=8 $Y=2.8 $X2=0 $Y2=0
cc_554 N_VPWR_c_726_n N_A_1210_367#_c_882_n 0.024453f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_748_n N_A_1210_367#_c_937_n 0.0124525f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_726_n N_A_1210_367#_c_937_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_557 N_VPWR_M1012_s N_A_1210_367#_c_905_n 0.00334931f $X=8.72 $Y=1.835 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_735_n N_A_1210_367#_c_905_n 0.0170777f $X=8.86 $Y=2.385 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_749_n N_A_1210_367#_c_941_n 0.0124525f $X=9.555 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_726_n N_A_1210_367#_c_941_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_726_n N_A_1210_367#_c_911_n 0.00246046f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_562 N_A_27_47#_c_944_n N_A_454_47#_M1007_s 0.00176461f $X=2.745 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_563 N_A_27_47#_c_961_n N_A_454_47#_M1029_s 0.00334627f $X=3.7 $Y=0.82 $X2=0
+ $Y2=0
cc_564 N_A_27_47#_M1013_d N_A_454_47#_c_1001_n 0.00335455f $X=2.7 $Y=0.235 $X2=0
+ $Y2=0
cc_565 N_A_27_47#_M1031_d N_A_454_47#_c_1001_n 0.00585785f $X=3.56 $Y=0.235
+ $X2=0 $Y2=0
cc_566 N_A_27_47#_c_944_n N_A_454_47#_c_1001_n 0.00358515f $X=2.745 $Y=1.07
+ $X2=0 $Y2=0
cc_567 N_A_27_47#_c_961_n N_A_454_47#_c_1001_n 0.0469484f $X=3.7 $Y=0.82 $X2=0
+ $Y2=0
cc_568 N_A_27_47#_c_947_n N_A_454_47#_c_1001_n 0.0127705f $X=2.84 $Y=0.82 $X2=0
+ $Y2=0
cc_569 N_A_27_47#_c_944_n N_A_454_47#_c_1005_n 0.0168098f $X=2.745 $Y=1.07 $X2=0
+ $Y2=0
cc_570 N_A_27_47#_c_961_n N_A_819_47#_c_1050_n 0.0211587f $X=3.7 $Y=0.82 $X2=0
+ $Y2=0
cc_571 N_A_27_47#_c_948_n N_VGND_c_1149_n 0.0816421f $X=1.855 $Y=0.392 $X2=0
+ $Y2=0
cc_572 N_A_27_47#_c_991_p N_VGND_c_1149_n 0.0135879f $X=1.965 $Y=0.53 $X2=0
+ $Y2=0
cc_573 N_A_27_47#_c_946_n N_VGND_c_1149_n 0.0207785f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_574 N_A_27_47#_M1010_s N_VGND_c_1156_n 0.00215158f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_575 N_A_27_47#_M1017_s N_VGND_c_1156_n 0.00223577f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_576 N_A_27_47#_M1037_s N_VGND_c_1156_n 0.00376625f $X=1.84 $Y=0.235 $X2=0
+ $Y2=0
cc_577 N_A_27_47#_M1013_d N_VGND_c_1156_n 0.00224381f $X=2.7 $Y=0.235 $X2=0
+ $Y2=0
cc_578 N_A_27_47#_M1031_d N_VGND_c_1156_n 0.0021598f $X=3.56 $Y=0.235 $X2=0
+ $Y2=0
cc_579 N_A_27_47#_c_948_n N_VGND_c_1156_n 0.0514937f $X=1.855 $Y=0.392 $X2=0
+ $Y2=0
cc_580 N_A_27_47#_c_991_p N_VGND_c_1156_n 0.00855309f $X=1.965 $Y=0.53 $X2=0
+ $Y2=0
cc_581 N_A_27_47#_c_946_n N_VGND_c_1156_n 0.0125051f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_582 N_A_454_47#_c_1001_n N_A_819_47#_M1001_d 0.00527599f $X=4.485 $Y=0.37
+ $X2=-0.19 $Y2=-0.245
cc_583 N_A_454_47#_c_1009_n N_A_819_47#_M1016_d 0.00332344f $X=5.345 $Y=0.34
+ $X2=0 $Y2=0
cc_584 N_A_454_47#_c_1001_n N_A_819_47#_c_1050_n 0.0191996f $X=4.485 $Y=0.37
+ $X2=0 $Y2=0
cc_585 N_A_454_47#_M1001_s N_A_819_47#_c_1051_n 0.00176461f $X=4.51 $Y=0.235
+ $X2=0 $Y2=0
cc_586 N_A_454_47#_c_1001_n N_A_819_47#_c_1051_n 0.00340518f $X=4.485 $Y=0.37
+ $X2=0 $Y2=0
cc_587 N_A_454_47#_c_1009_n N_A_819_47#_c_1051_n 0.00301993f $X=5.345 $Y=0.34
+ $X2=0 $Y2=0
cc_588 N_A_454_47#_c_1011_n N_A_819_47#_c_1051_n 0.016881f $X=4.65 $Y=0.38 $X2=0
+ $Y2=0
cc_589 N_A_454_47#_c_1009_n N_A_819_47#_c_1115_n 0.0124977f $X=5.345 $Y=0.34
+ $X2=0 $Y2=0
cc_590 N_A_454_47#_M1022_s N_A_819_47#_c_1053_n 0.00176461f $X=5.37 $Y=0.235
+ $X2=0 $Y2=0
cc_591 N_A_454_47#_c_1009_n N_A_819_47#_c_1053_n 0.00301993f $X=5.345 $Y=0.34
+ $X2=0 $Y2=0
cc_592 N_A_454_47#_c_1014_n N_A_819_47#_c_1053_n 0.016881f $X=5.51 $Y=0.38 $X2=0
+ $Y2=0
cc_593 N_A_454_47#_c_1001_n N_VGND_c_1149_n 0.112645f $X=4.485 $Y=0.37 $X2=0
+ $Y2=0
cc_594 N_A_454_47#_c_1009_n N_VGND_c_1149_n 0.0298674f $X=5.345 $Y=0.34 $X2=0
+ $Y2=0
cc_595 N_A_454_47#_c_1005_n N_VGND_c_1149_n 0.0187157f $X=2.41 $Y=0.37 $X2=0
+ $Y2=0
cc_596 N_A_454_47#_c_1011_n N_VGND_c_1149_n 0.0189074f $X=4.65 $Y=0.38 $X2=0
+ $Y2=0
cc_597 N_A_454_47#_c_1014_n N_VGND_c_1149_n 0.0189074f $X=5.51 $Y=0.38 $X2=0
+ $Y2=0
cc_598 N_A_454_47#_M1007_s N_VGND_c_1156_n 0.00223559f $X=2.27 $Y=0.235 $X2=0
+ $Y2=0
cc_599 N_A_454_47#_M1029_s N_VGND_c_1156_n 0.00223577f $X=3.13 $Y=0.235 $X2=0
+ $Y2=0
cc_600 N_A_454_47#_M1001_s N_VGND_c_1156_n 0.00223559f $X=4.51 $Y=0.235 $X2=0
+ $Y2=0
cc_601 N_A_454_47#_M1022_s N_VGND_c_1156_n 0.00223559f $X=5.37 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_A_454_47#_c_1001_n N_VGND_c_1156_n 0.0696302f $X=4.485 $Y=0.37 $X2=0
+ $Y2=0
cc_603 N_A_454_47#_c_1009_n N_VGND_c_1156_n 0.0187823f $X=5.345 $Y=0.34 $X2=0
+ $Y2=0
cc_604 N_A_454_47#_c_1005_n N_VGND_c_1156_n 0.0123226f $X=2.41 $Y=0.37 $X2=0
+ $Y2=0
cc_605 N_A_454_47#_c_1011_n N_VGND_c_1156_n 0.0124079f $X=4.65 $Y=0.38 $X2=0
+ $Y2=0
cc_606 N_A_454_47#_c_1014_n N_VGND_c_1156_n 0.0124079f $X=5.51 $Y=0.38 $X2=0
+ $Y2=0
cc_607 N_A_819_47#_c_1054_n N_VGND_M1008_d 0.00176461f $X=6.705 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_608 N_A_819_47#_c_1080_n N_VGND_M1021_d 0.00332667f $X=7.565 $Y=0.95 $X2=0
+ $Y2=0
cc_609 N_A_819_47#_c_1055_n N_VGND_M1018_s 0.00176461f $X=8.785 $Y=1.09 $X2=0
+ $Y2=0
cc_610 N_A_819_47#_c_1056_n N_VGND_M1035_s 0.00176461f $X=9.645 $Y=1.09 $X2=0
+ $Y2=0
cc_611 N_A_819_47#_c_1054_n N_VGND_c_1145_n 0.0170777f $X=6.705 $Y=1.1 $X2=0
+ $Y2=0
cc_612 N_A_819_47#_c_1080_n N_VGND_c_1146_n 0.0170777f $X=7.565 $Y=0.95 $X2=0
+ $Y2=0
cc_613 N_A_819_47#_c_1055_n N_VGND_c_1147_n 0.0170777f $X=8.785 $Y=1.09 $X2=0
+ $Y2=0
cc_614 N_A_819_47#_c_1056_n N_VGND_c_1148_n 0.0170777f $X=9.645 $Y=1.09 $X2=0
+ $Y2=0
cc_615 N_A_819_47#_c_1127_p N_VGND_c_1149_n 0.0124525f $X=5.94 $Y=0.42 $X2=0
+ $Y2=0
cc_616 N_A_819_47#_c_1128_p N_VGND_c_1151_n 0.0124525f $X=6.8 $Y=0.42 $X2=0
+ $Y2=0
cc_617 N_A_819_47#_c_1129_p N_VGND_c_1153_n 0.037765f $X=8.02 $Y=0.42 $X2=0
+ $Y2=0
cc_618 N_A_819_47#_c_1130_p N_VGND_c_1154_n 0.0124525f $X=8.88 $Y=0.42 $X2=0
+ $Y2=0
cc_619 N_A_819_47#_c_1057_n N_VGND_c_1155_n 0.0178111f $X=9.74 $Y=0.42 $X2=0
+ $Y2=0
cc_620 N_A_819_47#_M1001_d N_VGND_c_1156_n 0.0021598f $X=4.095 $Y=0.235 $X2=0
+ $Y2=0
cc_621 N_A_819_47#_M1016_d N_VGND_c_1156_n 0.00225186f $X=4.94 $Y=0.235 $X2=0
+ $Y2=0
cc_622 N_A_819_47#_M1033_d N_VGND_c_1156_n 0.00536646f $X=5.8 $Y=0.235 $X2=0
+ $Y2=0
cc_623 N_A_819_47#_M1020_s N_VGND_c_1156_n 0.0041006f $X=6.66 $Y=0.235 $X2=0
+ $Y2=0
cc_624 N_A_819_47#_M1038_s N_VGND_c_1156_n 0.00835561f $X=7.52 $Y=0.235 $X2=0
+ $Y2=0
cc_625 N_A_819_47#_M1034_d N_VGND_c_1156_n 0.00536646f $X=8.74 $Y=0.235 $X2=0
+ $Y2=0
cc_626 N_A_819_47#_M1039_d N_VGND_c_1156_n 0.00371702f $X=9.6 $Y=0.235 $X2=0
+ $Y2=0
cc_627 N_A_819_47#_c_1127_p N_VGND_c_1156_n 0.00730901f $X=5.94 $Y=0.42 $X2=0
+ $Y2=0
cc_628 N_A_819_47#_c_1128_p N_VGND_c_1156_n 0.00730901f $X=6.8 $Y=0.42 $X2=0
+ $Y2=0
cc_629 N_A_819_47#_c_1129_p N_VGND_c_1156_n 0.021305f $X=8.02 $Y=0.42 $X2=0
+ $Y2=0
cc_630 N_A_819_47#_c_1130_p N_VGND_c_1156_n 0.00730901f $X=8.88 $Y=0.42 $X2=0
+ $Y2=0
cc_631 N_A_819_47#_c_1057_n N_VGND_c_1156_n 0.0100304f $X=9.74 $Y=0.42 $X2=0
+ $Y2=0
cc_632 N_A_819_47#_c_1059_n N_VGND_c_1156_n 0.00223353f $X=6.835 $Y=0.95 $X2=0
+ $Y2=0
