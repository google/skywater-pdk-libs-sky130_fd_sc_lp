* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VGND a_22_259# X VNB nshort w=840000u l=150000u
+  ad=9.366e+11p pd=9.06e+06u as=2.352e+11p ps=2.24e+06u
M1001 VPWR a_22_259# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1256e+12p pd=9.52e+06u as=3.528e+11p ps=3.08e+06u
M1002 a_304_153# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.281e+11p pd=1.45e+06u as=0p ps=0u
M1003 a_508_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=0p ps=0u
M1004 a_304_153# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.281e+11p pd=1.45e+06u as=0p ps=0u
M1005 VPWR A1 a_508_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_22_259# a_304_153# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1007 X a_22_259# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_22_259# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_594_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.32e+06u
M1010 a_508_367# a_304_153# a_22_259# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1011 a_594_47# A1 a_22_259# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
