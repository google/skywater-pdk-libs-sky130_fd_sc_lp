* File: sky130_fd_sc_lp__o221a_lp.pex.spice
* Created: Fri Aug 28 11:07:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221A_LP%A_84_21# 1 2 3 10 12 16 19 21 23 25 26 27
+ 28 30 31 33 37 39 44 45 46 53 56
c109 56 0 8.31823e-20 $X=0.6 $Y=1.225
c110 27 0 1.83003e-19 $X=0.6 $Y=1.895
r111 51 53 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.96 $Y=0.85
+ $X2=4.15 $Y2=0.85
r112 45 48 2.66596 $w=8.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.82 $Y=2.055
+ $X2=3.82 $Y2=2.24
r113 45 46 10.4641 $w=8.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=2.055
+ $X2=3.82 $Y2=1.97
r114 41 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.15 $Y=1.015
+ $X2=4.15 $Y2=0.85
r115 41 46 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.15 $Y=1.015
+ $X2=4.15 $Y2=1.97
r116 40 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=2.055
+ $X2=1.98 $Y2=2.055
r117 39 45 10.4562 $w=1.7e-07 $l=4.15e-07 $layer=LI1_cond $X=3.405 $Y=2.055
+ $X2=3.82 $Y2=2.055
r118 39 40 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=3.405 $Y=2.055
+ $X2=2.145 $Y2=2.055
r119 35 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.14
+ $X2=1.98 $Y2=2.055
r120 35 37 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.98 $Y=2.14 $X2=1.98
+ $Y2=2.24
r121 34 43 3.37873 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.84 $Y=2.055
+ $X2=0.67 $Y2=2.055
r122 33 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=2.055
+ $X2=1.98 $Y2=2.055
r123 33 34 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=1.815 $Y=2.055
+ $X2=0.84 $Y2=2.055
r124 31 56 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.39
+ $X2=0.6 $Y2=1.225
r125 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=1.39 $X2=0.615 $Y2=1.39
r126 28 43 12.3276 $w=3.9e-07 $l=3.67287e-07 $layer=LI1_cond $X=0.645 $Y=1.7
+ $X2=0.67 $Y2=2.055
r127 28 30 9.16044 $w=3.88e-07 $l=3.1e-07 $layer=LI1_cond $X=0.645 $Y=1.7
+ $X2=0.645 $Y2=1.39
r128 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=0.855 $Y2=0.445
r129 22 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=0.805
+ $X2=0.495 $Y2=0.805
r130 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.855 $Y2=0.73
r131 21 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.57 $Y2=0.805
r132 19 27 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.59 $Y=2.595
+ $X2=0.59 $Y2=1.895
r133 16 27 31.8466 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.6 $Y=1.715
+ $X2=0.6 $Y2=1.895
r134 15 31 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=0.6 $Y=1.405
+ $X2=0.6 $Y2=1.39
r135 15 16 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=0.6 $Y=1.405
+ $X2=0.6 $Y2=1.715
r136 13 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=0.805
r137 13 56 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=1.225
r138 10 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.805
r139 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.445
r140 3 48 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.43
+ $Y=2.095 $X2=3.57 $Y2=2.24
r141 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.095 $X2=1.98 $Y2=2.24
r142 1 51 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=3.82
+ $Y=0.61 $X2=3.96 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%A1 3 9 11 12 13 14 15 16 17 21
c51 16 0 8.31823e-20 $X=1.2 $Y=1.295
c52 14 0 3.61764e-20 $X=1.28 $Y=0.73
r53 16 17 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.185 $Y=1.285
+ $X2=1.185 $Y2=1.665
r54 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.185
+ $Y=1.285 $X2=1.185 $Y2=1.285
r55 14 15 69.5192 $w=1.6e-07 $l=1.5e-07 $layer=POLY_cond $X=1.28 $Y=0.73
+ $X2=1.28 $Y2=0.88
r56 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.185 $Y=1.625
+ $X2=1.185 $Y2=1.285
r57 12 13 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.625
+ $X2=1.185 $Y2=1.79
r58 11 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.12
+ $X2=1.185 $Y2=1.285
r59 11 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.275 $Y=1.12
+ $X2=1.275 $Y2=0.88
r60 9 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.285 $Y=0.445
+ $X2=1.285 $Y2=0.73
r61 3 13 200.005 $w=2.5e-07 $l=8.05e-07 $layer=POLY_cond $X=1.225 $Y=2.595
+ $X2=1.225 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%A2 3 7 11 12 13 14 18
c44 13 0 6.68456e-20 $X=1.68 $Y=1.295
r45 13 14 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=1.717 $Y=1.285
+ $X2=1.717 $Y2=1.665
r46 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.755
+ $Y=1.285 $X2=1.755 $Y2=1.285
r47 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.755 $Y=1.625
+ $X2=1.755 $Y2=1.285
r48 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.625
+ $X2=1.755 $Y2=1.79
r49 10 18 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.12
+ $X2=1.755 $Y2=1.285
r50 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.715 $Y=0.445
+ $X2=1.715 $Y2=1.12
r51 3 12 200.005 $w=2.5e-07 $l=8.05e-07 $layer=POLY_cond $X=1.715 $Y=2.595
+ $X2=1.715 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%B2 3 7 8 9 11 12 13 17 19
c56 3 0 6.68456e-20 $X=2.285 $Y=2.595
r57 17 20 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.56
+ $X2=2.325 $Y2=1.725
r58 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.56
+ $X2=2.325 $Y2=1.395
r59 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=1.56 $X2=2.325 $Y2=1.56
r60 13 18 9.42908 $w=3.83e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=1.587
+ $X2=2.325 $Y2=1.587
r61 12 18 4.93904 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=1.587
+ $X2=2.325 $Y2=1.587
r62 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.805 $Y=0.63
+ $X2=2.805 $Y2=0.915
r63 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.73 $Y=0.555
+ $X2=2.805 $Y2=0.63
r64 7 8 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=2.73 $Y=0.555
+ $X2=2.375 $Y2=0.555
r65 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.3 $Y=0.63
+ $X2=2.375 $Y2=0.555
r66 5 19 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.3 $Y=0.63 $X2=2.3
+ $Y2=1.395
r67 3 20 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.285 $Y=2.595
+ $X2=2.285 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%B1 1 3 6 7 10 12 13 16 17
c53 10 0 5.08984e-20 $X=3.315 $Y=0.82
c54 7 0 1.41911e-19 $X=2.9 $Y=1.585
r55 16 19 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.245 $Y=1.495
+ $X2=3.245 $Y2=1.585
r56 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.245 $Y=1.495
+ $X2=3.245 $Y2=1.33
r57 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=1.495 $X2=3.245 $Y2=1.495
r58 13 17 6.02816 $w=3.23e-07 $l=1.7e-07 $layer=LI1_cond $X=3.167 $Y=1.665
+ $X2=3.167 $Y2=1.495
r59 10 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.315 $Y=0.82
+ $X2=3.315 $Y2=1.33
r60 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.585
+ $X2=3.245 $Y2=1.585
r61 6 7 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.08 $Y=1.585 $X2=2.9
+ $Y2=1.585
r62 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.825 $Y=1.66
+ $X2=2.9 $Y2=1.585
r63 4 12 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=2.825 $Y=1.66
+ $X2=2.825 $Y2=1.965
r64 1 12 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.775 $Y=2.09
+ $X2=2.775 $Y2=1.965
r65 1 3 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.775 $Y=2.09
+ $X2=2.775 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%C1 1 3 4 5 8 11 12 15 16
r43 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.495
+ $X2=3.785 $Y2=1.66
r44 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.495
+ $X2=3.785 $Y2=1.33
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.785
+ $Y=1.495 $X2=3.785 $Y2=1.495
r46 12 16 4.81032 $w=4.58e-07 $l=1.85e-07 $layer=LI1_cond $X=3.6 $Y=1.56
+ $X2=3.785 $Y2=1.56
r47 11 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.745 $Y=1.87
+ $X2=3.745 $Y2=1.66
r48 8 17 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.745 $Y=0.82
+ $X2=3.745 $Y2=1.33
r49 4 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.67 $Y=1.945
+ $X2=3.745 $Y2=1.87
r50 4 5 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.67 $Y=1.945 $X2=3.43
+ $Y2=1.945
r51 1 5 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.305 $Y=2.02
+ $X2=3.43 $Y2=1.945
r52 1 3 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.305 $Y=2.02
+ $X2=3.305 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%X 1 2 12 13 14 15 26
r26 19 26 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=0.272 $Y=0.868
+ $X2=0.272 $Y2=0.925
r27 15 28 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=0.272 $Y=0.939
+ $X2=0.272 $Y2=1.04
r28 15 26 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=0.272 $Y=0.939
+ $X2=0.272 $Y2=0.925
r29 15 19 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=0.272 $Y=0.854
+ $X2=0.272 $Y2=0.868
r30 14 15 12.8272 $w=3.43e-07 $l=3.84e-07 $layer=LI1_cond $X=0.272 $Y=0.47
+ $X2=0.272 $Y2=0.854
r31 13 28 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=0.185 $Y=2.075
+ $X2=0.185 $Y2=1.04
r32 12 13 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.295 $Y=2.24
+ $X2=0.295 $Y2=2.075
r33 2 12 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.18
+ $Y=2.095 $X2=0.325 $Y2=2.24
r34 1 14 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%VPWR 1 2 11 15 17 19 29 30 33 36
c44 11 0 1.83003e-19 $X=0.855 $Y=2.485
r45 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=3.04 $Y2=3.33
r50 27 29 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=0.855 $Y2=3.33
r57 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.02 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=3.04 $Y2=3.33
r59 19 25 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=3.245
+ $X2=3.04 $Y2=3.33
r63 13 15 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=3.04 $Y=3.245
+ $X2=3.04 $Y2=2.485
r64 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=3.245
+ $X2=0.855 $Y2=3.33
r65 9 11 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.855 $Y=3.245
+ $X2=0.855 $Y2=2.485
r66 2 15 300 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=2.9
+ $Y=2.095 $X2=3.04 $Y2=2.485
r67 1 11 300 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=2 $X=0.715
+ $Y=2.095 $X2=0.855 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%VGND 1 2 9 12 13 14 20 26 27 31
r51 31 34 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.01
+ $Y2=0.28
r52 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r53 24 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.01
+ $Y2=0
r54 24 26 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=2.175 $Y=0
+ $X2=4.08 $Y2=0
r55 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=2.01
+ $Y2=0
r57 20 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.68
+ $Y2=0
r58 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r59 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r60 14 27 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r61 14 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 14 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 12 17 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r64 12 13 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.03
+ $Y2=0
r65 11 22 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.68
+ $Y2=0
r66 11 13 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.03
+ $Y2=0
r67 7 13 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=0.085
+ $X2=1.03 $Y2=0
r68 7 9 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=1.03 $Y=0.085 $X2=1.03
+ $Y2=0.445
r69 2 34 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.235 $X2=2.01 $Y2=0.28
r70 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%A_272_47# 1 2 7 10 14
c37 7 0 8.70748e-20 $X=2.935 $Y=0.63
r38 14 17 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.1 $Y=0.63 $X2=3.1
+ $Y2=0.735
r39 10 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.5 $Y=0.47 $X2=1.5
+ $Y2=0.63
r40 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=0.63 $X2=1.5
+ $Y2=0.63
r41 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0.63 $X2=3.1
+ $Y2=0.63
r42 7 8 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=2.935 $Y=0.63
+ $X2=1.665 $Y2=0.63
r43 2 17 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=2.88
+ $Y=0.705 $X2=3.1 $Y2=0.735
r44 1 10 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.235 $X2=1.5 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_LP%A_490_141# 1 2 7 11 14
r28 14 16 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.59 $Y=0.98
+ $X2=2.59 $Y2=1.075
r29 9 11 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=3.57 $Y=0.99 $X2=3.57
+ $Y2=0.85
r30 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=1.075
+ $X2=2.59 $Y2=1.075
r31 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.445 $Y=1.075
+ $X2=3.57 $Y2=0.99
r32 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.445 $Y=1.075
+ $X2=2.755 $Y2=1.075
r33 2 11 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=3.39
+ $Y=0.61 $X2=3.53 $Y2=0.85
r34 1 14 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.705 $X2=2.59 $Y2=0.98
.ends

