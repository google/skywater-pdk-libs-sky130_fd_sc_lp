* File: sky130_fd_sc_lp__a41o_m.pxi.spice
* Created: Wed Sep  2 09:29:21 2020
* 
x_PM_SKY130_FD_SC_LP__A41O_M%A_80_153# N_A_80_153#_M1004_d N_A_80_153#_M1002_s
+ N_A_80_153#_c_93_n N_A_80_153#_M1009_g N_A_80_153#_c_87_n N_A_80_153#_M1010_g
+ N_A_80_153#_c_88_n N_A_80_153#_c_95_n N_A_80_153#_c_89_n N_A_80_153#_c_97_n
+ N_A_80_153#_c_90_n N_A_80_153#_c_128_p N_A_80_153#_c_98_n N_A_80_153#_c_99_n
+ N_A_80_153#_c_136_p N_A_80_153#_c_91_n N_A_80_153#_c_92_n
+ PM_SKY130_FD_SC_LP__A41O_M%A_80_153#
x_PM_SKY130_FD_SC_LP__A41O_M%B1 N_B1_M1004_g N_B1_M1002_g N_B1_c_160_n
+ N_B1_c_161_n B1 B1 B1 N_B1_c_158_n PM_SKY130_FD_SC_LP__A41O_M%B1
x_PM_SKY130_FD_SC_LP__A41O_M%A1 N_A1_M1001_g N_A1_M1000_g N_A1_c_207_n
+ N_A1_c_212_n A1 A1 A1 A1 A1 N_A1_c_209_n PM_SKY130_FD_SC_LP__A41O_M%A1
x_PM_SKY130_FD_SC_LP__A41O_M%A2 N_A2_M1006_g N_A2_M1007_g N_A2_c_259_n
+ N_A2_c_260_n N_A2_c_261_n A2 A2 A2 A2 A2 N_A2_c_263_n
+ PM_SKY130_FD_SC_LP__A41O_M%A2
x_PM_SKY130_FD_SC_LP__A41O_M%A3 N_A3_M1008_g N_A3_M1003_g N_A3_c_304_n
+ N_A3_c_309_n A3 A3 A3 A3 N_A3_c_306_n PM_SKY130_FD_SC_LP__A41O_M%A3
x_PM_SKY130_FD_SC_LP__A41O_M%A4 N_A4_M1005_g N_A4_M1011_g N_A4_c_350_n
+ N_A4_c_351_n N_A4_c_357_n N_A4_c_352_n A4 A4 A4 A4 N_A4_c_354_n
+ PM_SKY130_FD_SC_LP__A41O_M%A4
x_PM_SKY130_FD_SC_LP__A41O_M%X N_X_M1010_s N_X_M1009_s X X X X X X X N_X_c_387_n
+ PM_SKY130_FD_SC_LP__A41O_M%X
x_PM_SKY130_FD_SC_LP__A41O_M%VPWR N_VPWR_M1009_d N_VPWR_M1000_d N_VPWR_M1003_d
+ N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n
+ N_VPWR_c_408_n N_VPWR_c_409_n VPWR N_VPWR_c_410_n N_VPWR_c_411_n
+ N_VPWR_c_402_n N_VPWR_c_413_n PM_SKY130_FD_SC_LP__A41O_M%VPWR
x_PM_SKY130_FD_SC_LP__A41O_M%A_300_508# N_A_300_508#_M1002_d
+ N_A_300_508#_M1007_d N_A_300_508#_M1011_d N_A_300_508#_c_455_n
+ N_A_300_508#_c_456_n N_A_300_508#_c_457_n N_A_300_508#_c_458_n
+ N_A_300_508#_c_459_n N_A_300_508#_c_460_n N_A_300_508#_c_461_n
+ PM_SKY130_FD_SC_LP__A41O_M%A_300_508#
x_PM_SKY130_FD_SC_LP__A41O_M%VGND N_VGND_M1010_d N_VGND_M1005_d N_VGND_c_494_n
+ N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n VGND N_VGND_c_498_n
+ N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n PM_SKY130_FD_SC_LP__A41O_M%VGND
cc_1 VNB N_A_80_153#_c_87_n 0.0197677f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.765
cc_2 VNB N_A_80_153#_c_88_n 0.0228317f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.84
cc_3 VNB N_A_80_153#_c_89_n 0.00676206f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.01
cc_4 VNB N_A_80_153#_c_90_n 0.0210101f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.86
cc_5 VNB N_A_80_153#_c_91_n 0.00198732f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=0.51
cc_6 VNB N_A_80_153#_c_92_n 0.0406555f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.845
cc_7 VNB N_B1_M1004_g 0.0614417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB B1 0.00360845f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.445
cc_9 VNB N_B1_c_158_n 0.0141057f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.945
cc_10 VNB N_A1_M1001_g 0.0385443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_207_n 0.02506f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_12 VNB A1 0.00387734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_209_n 0.0193653f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.01
cc_14 VNB N_A2_M1007_g 0.0108825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_259_n 0.0178632f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.032
cc_16 VNB N_A2_c_260_n 0.0245543f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.328
cc_17 VNB N_A2_c_261_n 0.0176119f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.515
cc_18 VNB A2 0.00286215f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_19 VNB N_A2_c_263_n 0.018196f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.945
cc_20 VNB N_A3_M1008_g 0.0379042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_c_304_n 0.017609f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.515
cc_22 VNB A3 0.0126846f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_23 VNB N_A3_c_306_n 0.0182566f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.515
cc_24 VNB N_A4_M1005_g 0.0267104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A4_c_350_n 0.00942658f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.328
cc_26 VNB N_A4_c_351_n 0.0453984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A4_c_352_n 0.0191629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB A4 0.0367555f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.515
cc_29 VNB N_A4_c_354_n 0.0289471f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.48
cc_30 VNB X 0.0518257f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.915
cc_31 VNB N_X_c_387_n 0.0168319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_402_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_494_n 0.00494119f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.032
cc_34 VNB N_VGND_c_495_n 0.0126216f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_35 VNB N_VGND_c_496_n 0.023571f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.445
cc_36 VNB N_VGND_c_497_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.445
cc_37 VNB N_VGND_c_498_n 0.0611883f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.395
cc_38 VNB N_VGND_c_499_n 0.0155085f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=2.48
cc_39 VNB N_VGND_c_500_n 0.217959f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.48
cc_40 VNB N_VGND_c_501_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=2.685
cc_41 VPB N_A_80_153#_c_93_n 0.0248979f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.328
cc_42 VPB N_A_80_153#_M1009_g 0.0256331f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_43 VPB N_A_80_153#_c_95_n 0.0227895f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.515
cc_44 VPB N_A_80_153#_c_89_n 0.00159457f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.01
cc_45 VPB N_A_80_153#_c_97_n 0.0234893f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.01
cc_46 VPB N_A_80_153#_c_98_n 0.0179449f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=2.48
cc_47 VPB N_A_80_153#_c_99_n 0.00150838f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.48
cc_48 VPB N_A_80_153#_c_92_n 0.00921799f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.845
cc_49 VPB N_B1_M1002_g 0.0334556f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.915
cc_50 VPB N_B1_c_160_n 0.0274518f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_51 VPB N_B1_c_161_n 0.0344271f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB B1 0.00208417f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.445
cc_53 VPB N_B1_c_158_n 0.00419918f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.945
cc_54 VPB N_A1_M1000_g 0.0490746f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.915
cc_55 VPB N_A1_c_207_n 0.00140001f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_56 VPB N_A1_c_212_n 0.0238258f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_57 VPB A1 0.00677994f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A2_M1007_g 0.0541064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB A2 0.00465125f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_60 VPB N_A3_M1003_g 0.0447179f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.915
cc_61 VPB N_A3_c_304_n 0.00539071f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.515
cc_62 VPB N_A3_c_309_n 0.0165621f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_63 VPB A3 0.00715518f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_64 VPB N_A4_M1011_g 0.0301524f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.915
cc_65 VPB N_A4_c_350_n 0.0310055f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.328
cc_66 VPB N_A4_c_357_n 0.0312125f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.84
cc_67 VPB A4 0.028206f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.515
cc_68 VPB X 0.0489863f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.915
cc_69 VPB N_VPWR_c_403_n 0.00707402f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_70 VPB N_VPWR_c_404_n 0.00331778f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.445
cc_71 VPB N_VPWR_c_405_n 0.00774912f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.84
cc_72 VPB N_VPWR_c_406_n 0.0307955f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.945
cc_73 VPB N_VPWR_c_407_n 0.00601765f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.395
cc_74 VPB N_VPWR_c_408_n 0.0174159f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.01
cc_75 VPB N_VPWR_c_409_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.01
cc_76 VPB N_VPWR_c_410_n 0.0163199f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=2.48
cc_77 VPB N_VPWR_c_411_n 0.0265015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_402_n 0.0734393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_413_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_300_508#_c_455_n 0.00121421f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_81 VPB N_A_300_508#_c_456_n 0.013199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_300_508#_c_457_n 0.00371229f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.765
cc_83 VPB N_A_300_508#_c_458_n 0.0012004f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.84
cc_84 VPB N_A_300_508#_c_459_n 0.0200261f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.84
cc_85 VPB N_A_300_508#_c_460_n 0.00317049f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.395
cc_86 VPB N_A_300_508#_c_461_n 0.00601353f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.01
cc_87 N_A_80_153#_c_87_n N_B1_M1004_g 0.0215275f $X=0.685 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_80_153#_c_89_n N_B1_M1004_g 0.00782749f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_89 N_A_80_153#_c_90_n N_B1_M1004_g 0.0130288f $X=1.225 $Y=0.86 $X2=0 $Y2=0
cc_90 N_A_80_153#_c_91_n N_B1_M1004_g 0.00304795f $X=1.33 $Y=0.51 $X2=0 $Y2=0
cc_91 N_A_80_153#_c_92_n N_B1_M1004_g 0.0100762f $X=0.587 $Y=1.845 $X2=0 $Y2=0
cc_92 N_A_80_153#_c_93_n N_B1_M1002_g 0.00578926f $X=0.587 $Y=2.328 $X2=0 $Y2=0
cc_93 N_A_80_153#_c_89_n N_B1_M1002_g 8.04502e-19 $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_94 N_A_80_153#_c_98_n N_B1_M1002_g 0.0021779f $X=1.105 $Y=2.48 $X2=0 $Y2=0
cc_95 N_A_80_153#_c_89_n N_B1_c_160_n 0.00124165f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_96 N_A_80_153#_c_97_n N_B1_c_160_n 0.0118513f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_97 N_A_80_153#_c_93_n N_B1_c_161_n 0.0118513f $X=0.587 $Y=2.328 $X2=0 $Y2=0
cc_98 N_A_80_153#_c_98_n N_B1_c_161_n 0.00630579f $X=1.105 $Y=2.48 $X2=0 $Y2=0
cc_99 N_A_80_153#_c_89_n B1 0.0395567f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_100 N_A_80_153#_c_97_n B1 0.0012272f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_101 N_A_80_153#_c_90_n B1 0.0127635f $X=1.225 $Y=0.86 $X2=0 $Y2=0
cc_102 N_A_80_153#_c_98_n B1 0.0177586f $X=1.105 $Y=2.48 $X2=0 $Y2=0
cc_103 N_A_80_153#_c_92_n B1 5.36712e-19 $X=0.587 $Y=1.845 $X2=0 $Y2=0
cc_104 N_A_80_153#_c_89_n N_B1_c_158_n 0.00363602f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_105 N_A_80_153#_c_90_n N_B1_c_158_n 0.00272917f $X=1.225 $Y=0.86 $X2=0 $Y2=0
cc_106 N_A_80_153#_c_92_n N_B1_c_158_n 0.00492661f $X=0.587 $Y=1.845 $X2=0 $Y2=0
cc_107 N_A_80_153#_c_90_n N_A1_M1001_g 0.0013666f $X=1.225 $Y=0.86 $X2=0 $Y2=0
cc_108 N_A_80_153#_c_91_n N_A1_M1001_g 0.00371605f $X=1.33 $Y=0.51 $X2=0 $Y2=0
cc_109 N_A_80_153#_c_90_n A1 0.0131875f $X=1.225 $Y=0.86 $X2=0 $Y2=0
cc_110 N_A_80_153#_c_91_n A1 0.0208815f $X=1.33 $Y=0.51 $X2=0 $Y2=0
cc_111 N_A_80_153#_c_87_n X 0.00485291f $X=0.685 $Y=0.765 $X2=0 $Y2=0
cc_112 N_A_80_153#_c_88_n X 0.0493382f $X=0.685 $Y=0.84 $X2=0 $Y2=0
cc_113 N_A_80_153#_c_89_n X 0.100067f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_114 N_A_80_153#_c_128_p X 0.0130705f $X=0.695 $Y=0.86 $X2=0 $Y2=0
cc_115 N_A_80_153#_c_99_n X 0.0130705f $X=0.695 $Y=2.48 $X2=0 $Y2=0
cc_116 N_A_80_153#_c_88_n N_X_c_387_n 0.00664729f $X=0.685 $Y=0.84 $X2=0 $Y2=0
cc_117 N_A_80_153#_c_128_p N_X_c_387_n 0.00294507f $X=0.695 $Y=0.86 $X2=0 $Y2=0
cc_118 N_A_80_153#_M1009_g N_VPWR_c_403_n 0.0123507f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_119 N_A_80_153#_c_95_n N_VPWR_c_403_n 0.00128406f $X=0.587 $Y=2.515 $X2=0
+ $Y2=0
cc_120 N_A_80_153#_c_98_n N_VPWR_c_403_n 0.00829825f $X=1.105 $Y=2.48 $X2=0
+ $Y2=0
cc_121 N_A_80_153#_c_99_n N_VPWR_c_403_n 0.00771077f $X=0.695 $Y=2.48 $X2=0
+ $Y2=0
cc_122 N_A_80_153#_c_136_p N_VPWR_c_403_n 3.00173e-19 $X=1.21 $Y=2.685 $X2=0
+ $Y2=0
cc_123 N_A_80_153#_c_136_p N_VPWR_c_406_n 0.00543295f $X=1.21 $Y=2.685 $X2=0
+ $Y2=0
cc_124 N_A_80_153#_M1009_g N_VPWR_c_410_n 0.00486043f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_125 N_A_80_153#_M1009_g N_VPWR_c_402_n 0.0093594f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_126 N_A_80_153#_c_98_n N_VPWR_c_402_n 0.00997091f $X=1.105 $Y=2.48 $X2=0
+ $Y2=0
cc_127 N_A_80_153#_c_99_n N_VPWR_c_402_n 8.79797e-19 $X=0.695 $Y=2.48 $X2=0
+ $Y2=0
cc_128 N_A_80_153#_c_136_p N_VPWR_c_402_n 0.0069436f $X=1.21 $Y=2.685 $X2=0
+ $Y2=0
cc_129 N_A_80_153#_c_98_n N_A_300_508#_c_455_n 0.00485981f $X=1.105 $Y=2.48
+ $X2=0 $Y2=0
cc_130 N_A_80_153#_c_98_n N_A_300_508#_c_457_n 0.00584815f $X=1.105 $Y=2.48
+ $X2=0 $Y2=0
cc_131 N_A_80_153#_c_87_n N_VGND_c_494_n 0.00288714f $X=0.685 $Y=0.765 $X2=0
+ $Y2=0
cc_132 N_A_80_153#_c_90_n N_VGND_c_494_n 0.0114298f $X=1.225 $Y=0.86 $X2=0 $Y2=0
cc_133 N_A_80_153#_c_87_n N_VGND_c_496_n 0.00585385f $X=0.685 $Y=0.765 $X2=0
+ $Y2=0
cc_134 N_A_80_153#_c_88_n N_VGND_c_496_n 6.32862e-19 $X=0.685 $Y=0.84 $X2=0
+ $Y2=0
cc_135 N_A_80_153#_c_91_n N_VGND_c_498_n 0.00782832f $X=1.33 $Y=0.51 $X2=0 $Y2=0
cc_136 N_A_80_153#_M1004_d N_VGND_c_500_n 0.00680214f $X=1.19 $Y=0.235 $X2=0
+ $Y2=0
cc_137 N_A_80_153#_c_87_n N_VGND_c_500_n 0.00714621f $X=0.685 $Y=0.765 $X2=0
+ $Y2=0
cc_138 N_A_80_153#_c_88_n N_VGND_c_500_n 7.32533e-19 $X=0.685 $Y=0.84 $X2=0
+ $Y2=0
cc_139 N_A_80_153#_c_90_n N_VGND_c_500_n 0.0108793f $X=1.225 $Y=0.86 $X2=0 $Y2=0
cc_140 N_A_80_153#_c_128_p N_VGND_c_500_n 0.00426154f $X=0.695 $Y=0.86 $X2=0
+ $Y2=0
cc_141 N_A_80_153#_c_91_n N_VGND_c_500_n 0.00693508f $X=1.33 $Y=0.51 $X2=0 $Y2=0
cc_142 N_B1_M1004_g N_A1_M1001_g 0.0384935f $X=1.115 $Y=0.445 $X2=0 $Y2=0
cc_143 N_B1_c_160_n N_A1_M1000_g 0.00435287f $X=1.15 $Y=2.065 $X2=0 $Y2=0
cc_144 N_B1_c_161_n N_A1_M1000_g 0.030162f $X=1.425 $Y=2.14 $X2=0 $Y2=0
cc_145 B1 N_A1_M1000_g 5.12415e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_146 B1 N_A1_c_207_n 9.96992e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B1_c_158_n N_A1_c_207_n 0.00872829f $X=1.15 $Y=1.71 $X2=0 $Y2=0
cc_148 N_B1_c_160_n N_A1_c_212_n 0.00872829f $X=1.15 $Y=2.065 $X2=0 $Y2=0
cc_149 N_B1_M1004_g A1 0.00198496f $X=1.115 $Y=0.445 $X2=0 $Y2=0
cc_150 N_B1_c_160_n A1 0.00195346f $X=1.15 $Y=2.065 $X2=0 $Y2=0
cc_151 N_B1_c_161_n A1 5.26462e-19 $X=1.425 $Y=2.14 $X2=0 $Y2=0
cc_152 B1 A1 0.0414717f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B1_c_158_n A1 8.95359e-19 $X=1.15 $Y=1.71 $X2=0 $Y2=0
cc_154 B1 N_A1_c_209_n 0.00254286f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B1_M1002_g N_VPWR_c_403_n 0.00592828f $X=1.425 $Y=2.75 $X2=0 $Y2=0
cc_156 N_B1_M1002_g N_VPWR_c_404_n 0.00116144f $X=1.425 $Y=2.75 $X2=0 $Y2=0
cc_157 N_B1_M1002_g N_VPWR_c_406_n 0.00461464f $X=1.425 $Y=2.75 $X2=0 $Y2=0
cc_158 N_B1_M1002_g N_VPWR_c_402_n 0.00914415f $X=1.425 $Y=2.75 $X2=0 $Y2=0
cc_159 N_B1_M1002_g N_A_300_508#_c_455_n 5.61522e-19 $X=1.425 $Y=2.75 $X2=0
+ $Y2=0
cc_160 N_B1_M1002_g N_A_300_508#_c_457_n 0.00379141f $X=1.425 $Y=2.75 $X2=0
+ $Y2=0
cc_161 N_B1_M1004_g N_VGND_c_494_n 0.00288714f $X=1.115 $Y=0.445 $X2=0 $Y2=0
cc_162 N_B1_M1004_g N_VGND_c_498_n 0.00585385f $X=1.115 $Y=0.445 $X2=0 $Y2=0
cc_163 N_B1_M1004_g N_VGND_c_500_n 0.00630904f $X=1.115 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A1_c_207_n N_A2_M1007_g 0.00746673f $X=1.727 $Y=1.675 $X2=0 $Y2=0
cc_165 N_A1_c_212_n N_A2_M1007_g 0.047348f $X=1.727 $Y=1.825 $X2=0 $Y2=0
cc_166 A1 N_A2_M1007_g 3.61369e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_167 N_A1_M1001_g N_A2_c_259_n 0.0313206f $X=1.6 $Y=0.445 $X2=0 $Y2=0
cc_168 A1 N_A2_c_259_n 0.00473773f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_169 A1 N_A2_c_260_n 8.70585e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_170 N_A1_c_209_n N_A2_c_260_n 0.00864124f $X=1.69 $Y=1.32 $X2=0 $Y2=0
cc_171 N_A1_c_207_n N_A2_c_261_n 0.00864124f $X=1.727 $Y=1.675 $X2=0 $Y2=0
cc_172 N_A1_M1001_g A2 7.56644e-19 $X=1.6 $Y=0.445 $X2=0 $Y2=0
cc_173 N_A1_c_207_n A2 0.00193583f $X=1.727 $Y=1.675 $X2=0 $Y2=0
cc_174 N_A1_c_212_n A2 0.00354618f $X=1.727 $Y=1.825 $X2=0 $Y2=0
cc_175 A1 A2 0.0794202f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_176 N_A1_c_209_n A2 0.00101655f $X=1.69 $Y=1.32 $X2=0 $Y2=0
cc_177 N_A1_M1000_g N_VPWR_c_404_n 0.00825838f $X=1.855 $Y=2.75 $X2=0 $Y2=0
cc_178 N_A1_M1000_g N_VPWR_c_406_n 0.00383152f $X=1.855 $Y=2.75 $X2=0 $Y2=0
cc_179 N_A1_M1000_g N_VPWR_c_402_n 0.00388243f $X=1.855 $Y=2.75 $X2=0 $Y2=0
cc_180 N_A1_M1000_g N_A_300_508#_c_455_n 0.001666f $X=1.855 $Y=2.75 $X2=0 $Y2=0
cc_181 N_A1_M1000_g N_A_300_508#_c_456_n 0.0157953f $X=1.855 $Y=2.75 $X2=0 $Y2=0
cc_182 N_A1_c_212_n N_A_300_508#_c_456_n 3.56428e-19 $X=1.727 $Y=1.825 $X2=0
+ $Y2=0
cc_183 A1 N_A_300_508#_c_456_n 0.00393781f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_184 N_A1_c_212_n N_A_300_508#_c_457_n 0.0026015f $X=1.727 $Y=1.825 $X2=0
+ $Y2=0
cc_185 A1 N_A_300_508#_c_457_n 0.011423f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_186 N_A1_M1001_g N_VGND_c_498_n 0.0048701f $X=1.6 $Y=0.445 $X2=0 $Y2=0
cc_187 A1 N_VGND_c_498_n 0.00426263f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_188 N_A1_M1001_g N_VGND_c_500_n 0.00863017f $X=1.6 $Y=0.445 $X2=0 $Y2=0
cc_189 A1 N_VGND_c_500_n 0.00568396f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_190 A1 A_335_47# 0.00266388f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_191 N_A2_c_259_n N_A3_M1008_g 0.0210363f $X=2.23 $Y=0.765 $X2=0 $Y2=0
cc_192 A2 N_A3_M1008_g 0.00746154f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_193 N_A2_c_263_n N_A3_M1008_g 0.0139295f $X=2.23 $Y=0.93 $X2=0 $Y2=0
cc_194 N_A2_M1007_g N_A3_M1003_g 0.0368547f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_195 A2 N_A3_M1003_g 2.32971e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_196 N_A2_M1007_g N_A3_c_304_n 0.0226224f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_197 N_A2_c_261_n N_A3_c_304_n 0.0139295f $X=2.23 $Y=1.435 $X2=0 $Y2=0
cc_198 N_A2_M1007_g A3 0.00424257f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_199 A2 A3 0.0759025f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_200 N_A2_c_263_n A3 0.00394106f $X=2.23 $Y=0.93 $X2=0 $Y2=0
cc_201 N_A2_c_260_n N_A3_c_306_n 0.0139295f $X=2.23 $Y=1.27 $X2=0 $Y2=0
cc_202 N_A2_M1007_g N_VPWR_c_404_n 0.00825085f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_203 N_A2_M1007_g N_VPWR_c_408_n 0.00383152f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_204 N_A2_M1007_g N_VPWR_c_402_n 0.00388243f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_205 N_A2_M1007_g N_A_300_508#_c_456_n 0.0131492f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_206 A2 N_A_300_508#_c_456_n 0.0184333f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_207 N_A2_M1007_g N_A_300_508#_c_458_n 0.001666f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_208 N_A2_c_259_n N_VGND_c_498_n 0.00412296f $X=2.23 $Y=0.765 $X2=0 $Y2=0
cc_209 A2 N_VGND_c_498_n 0.00590724f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_210 N_A2_c_263_n N_VGND_c_498_n 0.0018659f $X=2.23 $Y=0.93 $X2=0 $Y2=0
cc_211 N_A2_c_259_n N_VGND_c_500_n 0.00662524f $X=2.23 $Y=0.765 $X2=0 $Y2=0
cc_212 A2 N_VGND_c_500_n 0.00743229f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_213 N_A2_c_263_n N_VGND_c_500_n 0.00215369f $X=2.23 $Y=0.93 $X2=0 $Y2=0
cc_214 A2 A_443_47# 0.00307071f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_215 N_A3_M1008_g N_A4_M1005_g 0.0567558f $X=2.68 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A3_M1003_g N_A4_c_350_n 0.00300267f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_217 N_A3_c_309_n N_A4_c_350_n 0.00788767f $X=2.77 $Y=1.9 $X2=0 $Y2=0
cc_218 A3 N_A4_c_350_n 0.0011322f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_219 A3 N_A4_c_351_n 0.00167026f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_220 N_A3_M1003_g N_A4_c_357_n 0.0271213f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_221 N_A3_c_304_n N_A4_c_352_n 0.00788767f $X=2.77 $Y=1.735 $X2=0 $Y2=0
cc_222 N_A3_M1008_g A4 4.6941e-19 $X=2.68 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A3_M1003_g A4 3.34916e-19 $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_224 A3 A4 0.0427562f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_225 N_A3_c_306_n A4 0.0024705f $X=2.77 $Y=1.395 $X2=0 $Y2=0
cc_226 N_A3_M1008_g N_A4_c_354_n 0.00283301f $X=2.68 $Y=0.445 $X2=0 $Y2=0
cc_227 A3 N_A4_c_354_n 0.00355323f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_228 N_A3_c_306_n N_A4_c_354_n 0.00788767f $X=2.77 $Y=1.395 $X2=0 $Y2=0
cc_229 N_A3_M1003_g N_VPWR_c_404_n 7.03005e-19 $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_230 N_A3_M1003_g N_VPWR_c_405_n 0.00169048f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_231 N_A3_M1003_g N_VPWR_c_408_n 0.00461464f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_232 N_A3_M1003_g N_VPWR_c_402_n 0.00468324f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_233 N_A3_M1003_g N_A_300_508#_c_458_n 9.325e-19 $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_234 N_A3_M1003_g N_A_300_508#_c_459_n 0.0119343f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_235 N_A3_c_309_n N_A_300_508#_c_459_n 0.00302311f $X=2.77 $Y=1.9 $X2=0 $Y2=0
cc_236 A3 N_A_300_508#_c_459_n 0.0189043f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_237 A3 N_A_300_508#_c_461_n 0.0043399f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_238 N_A3_M1008_g N_VGND_c_495_n 0.00238543f $X=2.68 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A3_M1008_g N_VGND_c_498_n 0.00585385f $X=2.68 $Y=0.445 $X2=0 $Y2=0
cc_240 N_A3_M1008_g N_VGND_c_500_n 0.00665118f $X=2.68 $Y=0.445 $X2=0 $Y2=0
cc_241 A3 N_VGND_c_500_n 0.0105945f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_242 N_A4_M1011_g N_VPWR_c_405_n 0.00327258f $X=3.145 $Y=2.75 $X2=0 $Y2=0
cc_243 N_A4_M1011_g N_VPWR_c_411_n 0.00461464f $X=3.145 $Y=2.75 $X2=0 $Y2=0
cc_244 N_A4_M1011_g N_VPWR_c_402_n 0.00472399f $X=3.145 $Y=2.75 $X2=0 $Y2=0
cc_245 N_A4_M1011_g N_A_300_508#_c_459_n 0.0168732f $X=3.145 $Y=2.75 $X2=0 $Y2=0
cc_246 N_A4_c_357_n N_A_300_508#_c_459_n 0.00868965f $X=3.34 $Y=2.215 $X2=0
+ $Y2=0
cc_247 A4 N_A_300_508#_c_459_n 0.01022f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_248 N_A4_M1011_g N_A_300_508#_c_460_n 0.0020107f $X=3.145 $Y=2.75 $X2=0 $Y2=0
cc_249 N_A4_M1005_g N_VGND_c_495_n 0.0113072f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A4_c_351_n N_VGND_c_495_n 0.00747768f $X=3.43 $Y=0.99 $X2=0 $Y2=0
cc_251 A4 N_VGND_c_495_n 0.00323297f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_252 N_A4_M1005_g N_VGND_c_498_n 0.00486043f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_253 N_A4_M1005_g N_VGND_c_500_n 0.00818711f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_254 A4 N_VGND_c_500_n 0.0101065f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_255 X N_VPWR_c_410_n 0.00831216f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_256 N_X_M1009_s N_VPWR_c_402_n 0.00489501f $X=0.135 $Y=2.675 $X2=0 $Y2=0
cc_257 X N_VPWR_c_402_n 0.0069578f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_258 N_X_c_387_n N_VGND_c_496_n 0.0257719f $X=0.47 $Y=0.43 $X2=0 $Y2=0
cc_259 N_X_M1010_s N_VGND_c_500_n 0.00234592f $X=0.345 $Y=0.235 $X2=0 $Y2=0
cc_260 N_X_c_387_n N_VGND_c_500_n 0.0159398f $X=0.47 $Y=0.43 $X2=0 $Y2=0
cc_261 N_VPWR_c_406_n N_A_300_508#_c_455_n 0.00493172f $X=1.905 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_402_n N_A_300_508#_c_455_n 0.00631623f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_404_n N_A_300_508#_c_456_n 0.0157665f $X=2.07 $Y=2.815 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_402_n N_A_300_508#_c_456_n 0.0116386f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_c_408_n N_A_300_508#_c_458_n 0.00493172f $X=2.825 $Y=3.33 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_402_n N_A_300_508#_c_458_n 0.00631623f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_405_n N_A_300_508#_c_459_n 0.0142847f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_402_n N_A_300_508#_c_459_n 0.0135041f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_c_411_n N_A_300_508#_c_460_n 0.00549876f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_402_n N_A_300_508#_c_460_n 0.00699584f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_271 N_VGND_c_500_n A_335_47# 0.0134089f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_272 N_VGND_c_500_n A_443_47# 0.0101616f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_273 N_VGND_c_500_n A_551_47# 0.00620535f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
