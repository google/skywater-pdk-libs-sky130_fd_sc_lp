* File: sky130_fd_sc_lp__mux2_lp2.pxi.spice
* Created: Fri Aug 28 10:44:21 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_LP2%A_84_259# N_A_84_259#_M1006_d N_A_84_259#_M1003_d
+ N_A_84_259#_c_76_n N_A_84_259#_M1010_g N_A_84_259#_M1001_g N_A_84_259#_M1007_g
+ N_A_84_259#_c_80_n N_A_84_259#_c_81_n N_A_84_259#_c_82_n N_A_84_259#_c_146_p
+ N_A_84_259#_c_89_p N_A_84_259#_c_112_p N_A_84_259#_c_83_n N_A_84_259#_c_84_n
+ N_A_84_259#_c_96_p PM_SKY130_FD_SC_LP__MUX2_LP2%A_84_259#
x_PM_SKY130_FD_SC_LP__MUX2_LP2%A_182_303# N_A_182_303#_M1009_d
+ N_A_182_303#_M1013_d N_A_182_303#_M1011_g N_A_182_303#_c_163_n
+ N_A_182_303#_c_164_n N_A_182_303#_M1012_g N_A_182_303#_c_165_n
+ N_A_182_303#_c_166_n N_A_182_303#_c_167_n N_A_182_303#_c_168_n
+ N_A_182_303#_c_204_n N_A_182_303#_c_207_n N_A_182_303#_c_175_n
+ N_A_182_303#_c_176_n N_A_182_303#_c_177_n N_A_182_303#_c_178_n
+ N_A_182_303#_c_169_n N_A_182_303#_c_180_n N_A_182_303#_c_170_n
+ PM_SKY130_FD_SC_LP__MUX2_LP2%A_182_303#
x_PM_SKY130_FD_SC_LP__MUX2_LP2%A1 N_A1_M1003_g N_A1_M1004_g N_A1_c_269_n
+ N_A1_c_270_n N_A1_c_271_n N_A1_c_272_n N_A1_c_273_n N_A1_c_274_n A1 A1
+ N_A1_c_276_n PM_SKY130_FD_SC_LP__MUX2_LP2%A1
x_PM_SKY130_FD_SC_LP__MUX2_LP2%A0 N_A0_c_335_n N_A0_M1006_g N_A0_c_336_n
+ N_A0_M1000_g N_A0_c_338_n A0 N_A0_c_340_n PM_SKY130_FD_SC_LP__MUX2_LP2%A0
x_PM_SKY130_FD_SC_LP__MUX2_LP2%S N_S_M1005_g N_S_M1002_g N_S_M1013_g N_S_M1008_g
+ N_S_M1009_g S S S N_S_c_383_n PM_SKY130_FD_SC_LP__MUX2_LP2%S
x_PM_SKY130_FD_SC_LP__MUX2_LP2%X N_X_M1001_s N_X_M1010_s N_X_c_441_n X X X X X X
+ X PM_SKY130_FD_SC_LP__MUX2_LP2%X
x_PM_SKY130_FD_SC_LP__MUX2_LP2%VPWR N_VPWR_M1010_d N_VPWR_M1005_d N_VPWR_c_462_n
+ N_VPWR_c_463_n VPWR N_VPWR_c_464_n N_VPWR_c_465_n N_VPWR_c_461_n
+ N_VPWR_c_467_n N_VPWR_c_468_n PM_SKY130_FD_SC_LP__MUX2_LP2%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_LP2%VGND N_VGND_M1007_d N_VGND_M1002_d N_VGND_c_506_n
+ N_VGND_c_507_n VGND N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n
+ N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n PM_SKY130_FD_SC_LP__MUX2_LP2%VGND
cc_1 VNB N_A_84_259#_c_76_n 0.0657263f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.42
cc_2 VNB N_A_84_259#_M1010_g 0.018416f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_3 VNB N_A_84_259#_M1001_g 0.0249044f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.495
cc_4 VNB N_A_84_259#_M1007_g 0.0226876f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.495
cc_5 VNB N_A_84_259#_c_80_n 0.0123414f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.07
cc_6 VNB N_A_84_259#_c_81_n 0.00150815f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=0.905
cc_7 VNB N_A_84_259#_c_82_n 0.010471f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.065
cc_8 VNB N_A_84_259#_c_83_n 0.0056893f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.07
cc_9 VNB N_A_84_259#_c_84_n 0.00298469f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.495
cc_10 VNB N_A_182_303#_c_163_n 0.0382795f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.495
cc_11 VNB N_A_182_303#_c_164_n 0.0169687f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.495
cc_12 VNB N_A_182_303#_c_165_n 0.0177115f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.495
cc_13 VNB N_A_182_303#_c_166_n 0.00813942f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.495
cc_14 VNB N_A_182_303#_c_167_n 0.0288261f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.07
cc_15 VNB N_A_182_303#_c_168_n 0.00354722f $X=-0.19 $Y=-0.245 $X2=1.505
+ $Y2=0.515
cc_16 VNB N_A_182_303#_c_169_n 0.0455057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_182_303#_c_170_n 0.0251105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1004_g 0.0258607f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.42
cc_19 VNB N_A1_c_269_n 0.0039977f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_20 VNB N_A1_c_270_n 0.0226216f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.495
cc_21 VNB N_A1_c_271_n 0.0059476f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.905
cc_22 VNB N_A1_c_272_n 0.00299153f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.495
cc_23 VNB N_A1_c_273_n 0.00472487f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.495
cc_24 VNB N_A1_c_274_n 0.0348534f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.07
cc_25 VNB A1 0.00378408f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.07
cc_26 VNB N_A1_c_276_n 0.00519794f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=2.15
cc_27 VNB N_A0_c_335_n 0.0192762f $X=-0.19 $Y=-0.245 $X2=2.135 $Y2=0.285
cc_28 VNB N_A0_c_336_n 0.0107181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A0_M1000_g 0.00268641f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_30 VNB N_A0_c_338_n 0.027262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB A0 0.00571694f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.905
cc_32 VNB N_A0_c_340_n 0.0485281f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.905
cc_33 VNB N_S_M1002_g 0.053977f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.42
cc_34 VNB N_S_M1008_g 0.0468596f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.905
cc_35 VNB N_S_M1009_g 0.0534738f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.07
cc_36 VNB N_S_c_383_n 0.0540565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB X 0.0607617f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.905
cc_38 VNB N_VPWR_c_461_n 0.203486f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.15
cc_39 VNB N_VGND_c_506_n 0.00739108f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_40 VNB N_VGND_c_507_n 0.0131801f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.495
cc_41 VNB N_VGND_c_508_n 0.0273115f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.495
cc_42 VNB N_VGND_c_509_n 0.0561827f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.07
cc_43 VNB N_VGND_c_510_n 0.0316536f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.43
cc_44 VNB N_VGND_c_511_n 0.297976f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.15
cc_45 VNB N_VGND_c_512_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_513_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.495
cc_47 VPB N_A_84_259#_M1010_g 0.0471182f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.505
cc_48 VPB N_A_84_259#_c_82_n 0.00271436f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=2.065
cc_49 VPB N_A_182_303#_M1011_g 0.0280101f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.505
cc_50 VPB N_A_182_303#_c_165_n 0.021543f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.495
cc_51 VPB N_A_182_303#_c_166_n 0.00722928f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.495
cc_52 VPB N_A_182_303#_c_168_n 0.00238588f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=0.515
cc_53 VPB N_A_182_303#_c_175_n 0.00211757f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=0.43
cc_54 VPB N_A_182_303#_c_176_n 0.0097966f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.15
cc_55 VPB N_A_182_303#_c_177_n 0.0191615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_182_303#_c_178_n 0.0401659f $X=-0.19 $Y=1.655 $X2=2.66 $Y2=0.535
cc_57 VPB N_A_182_303#_c_169_n 0.0203918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_182_303#_c_180_n 0.00704942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A1_M1003_g 0.0267967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A1_c_269_n 0.00632763f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.505
cc_61 VPB N_A1_c_270_n 0.0130328f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.495
cc_62 VPB N_A0_M1000_g 0.0363301f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.505
cc_63 VPB N_S_M1005_g 0.0278368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_S_M1013_g 0.0368868f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.905
cc_65 VPB N_S_c_383_n 0.0487801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_X_c_441_n 0.0216297f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.505
cc_67 VPB X 0.0278732f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.905
cc_68 VPB X 0.00635268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_462_n 0.00547558f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.905
cc_70 VPB N_VPWR_c_463_n 0.00280617f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=0.905
cc_71 VPB N_VPWR_c_464_n 0.058257f $X=-0.19 $Y=1.655 $X2=1.42 $Y2=1.07
cc_72 VPB N_VPWR_c_465_n 0.0431961f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=0.43
cc_73 VPB N_VPWR_c_461_n 0.095275f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.15
cc_74 VPB N_VPWR_c_467_n 0.0252051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_468_n 0.00546567f $X=-0.19 $Y=1.655 $X2=2.66 $Y2=0.495
cc_76 N_A_84_259#_M1010_g N_A_182_303#_M1011_g 0.0156f $X=0.545 $Y=2.505 $X2=0
+ $Y2=0
cc_77 N_A_84_259#_c_82_n N_A_182_303#_M1011_g 0.00507506f $X=1.505 $Y=2.065
+ $X2=0 $Y2=0
cc_78 N_A_84_259#_c_89_p N_A_182_303#_M1011_g 0.00667497f $X=1.59 $Y=2.15 $X2=0
+ $Y2=0
cc_79 N_A_84_259#_c_76_n N_A_182_303#_c_163_n 0.00615583f $X=0.545 $Y=1.42 $X2=0
+ $Y2=0
cc_80 N_A_84_259#_c_80_n N_A_182_303#_c_163_n 0.00776353f $X=1.42 $Y=1.07 $X2=0
+ $Y2=0
cc_81 N_A_84_259#_c_82_n N_A_182_303#_c_163_n 0.017378f $X=1.505 $Y=2.065 $X2=0
+ $Y2=0
cc_82 N_A_84_259#_c_83_n N_A_182_303#_c_163_n 0.00630992f $X=1.505 $Y=1.07 $X2=0
+ $Y2=0
cc_83 N_A_84_259#_M1007_g N_A_182_303#_c_164_n 0.00472057f $X=0.86 $Y=0.495
+ $X2=0 $Y2=0
cc_84 N_A_84_259#_c_81_n N_A_182_303#_c_164_n 0.0040032f $X=1.505 $Y=0.905 $X2=0
+ $Y2=0
cc_85 N_A_84_259#_c_96_p N_A_182_303#_c_164_n 0.0143678f $X=2.495 $Y=0.535 $X2=0
+ $Y2=0
cc_86 N_A_84_259#_c_76_n N_A_182_303#_c_165_n 0.00228598f $X=0.545 $Y=1.42 $X2=0
+ $Y2=0
cc_87 N_A_84_259#_M1010_g N_A_182_303#_c_165_n 0.0184787f $X=0.545 $Y=2.505
+ $X2=0 $Y2=0
cc_88 N_A_84_259#_c_80_n N_A_182_303#_c_165_n 0.00736108f $X=1.42 $Y=1.07 $X2=0
+ $Y2=0
cc_89 N_A_84_259#_c_82_n N_A_182_303#_c_166_n 0.00931647f $X=1.505 $Y=2.065
+ $X2=0 $Y2=0
cc_90 N_A_84_259#_c_76_n N_A_182_303#_c_167_n 0.00853983f $X=0.545 $Y=1.42 $X2=0
+ $Y2=0
cc_91 N_A_84_259#_M1007_g N_A_182_303#_c_167_n 0.00376291f $X=0.86 $Y=0.495
+ $X2=0 $Y2=0
cc_92 N_A_84_259#_c_80_n N_A_182_303#_c_167_n 0.00207868f $X=1.42 $Y=1.07 $X2=0
+ $Y2=0
cc_93 N_A_84_259#_c_81_n N_A_182_303#_c_167_n 0.00927672f $X=1.505 $Y=0.905
+ $X2=0 $Y2=0
cc_94 N_A_84_259#_c_83_n N_A_182_303#_c_167_n 0.00218092f $X=1.505 $Y=1.07 $X2=0
+ $Y2=0
cc_95 N_A_84_259#_c_76_n N_A_182_303#_c_168_n 2.05376e-19 $X=0.545 $Y=1.42 $X2=0
+ $Y2=0
cc_96 N_A_84_259#_M1010_g N_A_182_303#_c_168_n 0.00802073f $X=0.545 $Y=2.505
+ $X2=0 $Y2=0
cc_97 N_A_84_259#_c_80_n N_A_182_303#_c_168_n 0.0187215f $X=1.42 $Y=1.07 $X2=0
+ $Y2=0
cc_98 N_A_84_259#_c_82_n N_A_182_303#_c_168_n 0.0359208f $X=1.505 $Y=2.065 $X2=0
+ $Y2=0
cc_99 N_A_84_259#_M1003_d N_A_182_303#_c_204_n 0.00625132f $X=2.02 $Y=2.005
+ $X2=0 $Y2=0
cc_100 N_A_84_259#_c_89_p N_A_182_303#_c_204_n 0.00799641f $X=1.59 $Y=2.15 $X2=0
+ $Y2=0
cc_101 N_A_84_259#_c_112_p N_A_182_303#_c_204_n 0.0390209f $X=2.16 $Y=2.15 $X2=0
+ $Y2=0
cc_102 N_A_84_259#_M1010_g N_A_182_303#_c_207_n 0.0021874f $X=0.545 $Y=2.505
+ $X2=0 $Y2=0
cc_103 N_A_84_259#_c_112_p N_A1_M1003_g 0.0130778f $X=2.16 $Y=2.15 $X2=0 $Y2=0
cc_104 N_A_84_259#_c_84_n N_A1_M1004_g 0.00597773f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_105 N_A_84_259#_c_82_n N_A1_c_269_n 0.0250969f $X=1.505 $Y=2.065 $X2=0 $Y2=0
cc_106 N_A_84_259#_c_112_p N_A1_c_269_n 0.0309476f $X=2.16 $Y=2.15 $X2=0 $Y2=0
cc_107 N_A_84_259#_c_82_n N_A1_c_270_n 0.00548145f $X=1.505 $Y=2.065 $X2=0 $Y2=0
cc_108 N_A_84_259#_c_112_p N_A1_c_270_n 0.00159134f $X=2.16 $Y=2.15 $X2=0 $Y2=0
cc_109 N_A_84_259#_c_84_n N_A1_c_272_n 0.0123938f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_110 N_A_84_259#_c_84_n N_A1_c_273_n 0.0145882f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_111 N_A_84_259#_c_84_n N_A1_c_274_n 0.00159161f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_112 N_A_84_259#_c_84_n A1 0.0112319f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_113 N_A_84_259#_c_81_n N_A0_c_335_n 4.148e-19 $X=1.505 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_84_259#_c_84_n N_A0_c_335_n 0.00448919f $X=2.66 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_84_259#_c_96_p N_A0_c_335_n 0.0119615f $X=2.495 $Y=0.535 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_84_259#_c_81_n A0 0.00340374f $X=1.505 $Y=0.905 $X2=0 $Y2=0
cc_117 N_A_84_259#_c_83_n A0 0.0106929f $X=1.505 $Y=1.07 $X2=0 $Y2=0
cc_118 N_A_84_259#_c_96_p A0 0.0133185f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_119 N_A_84_259#_c_83_n N_A0_c_340_n 0.00193138f $X=1.505 $Y=1.07 $X2=0 $Y2=0
cc_120 N_A_84_259#_c_96_p N_A0_c_340_n 0.00606424f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_121 N_A_84_259#_c_84_n N_S_M1002_g 3.579e-19 $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_122 N_A_84_259#_M1010_g N_X_c_441_n 0.0144604f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_123 N_A_84_259#_c_76_n X 0.0217614f $X=0.545 $Y=1.42 $X2=0 $Y2=0
cc_124 N_A_84_259#_M1010_g X 0.0326609f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_125 N_A_84_259#_M1001_g X 0.0156799f $X=0.5 $Y=0.495 $X2=0 $Y2=0
cc_126 N_A_84_259#_M1007_g X 0.00214948f $X=0.86 $Y=0.495 $X2=0 $Y2=0
cc_127 N_A_84_259#_c_80_n X 0.0257681f $X=1.42 $Y=1.07 $X2=0 $Y2=0
cc_128 N_A_84_259#_M1010_g X 0.00341836f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_129 N_A_84_259#_M1010_g N_VPWR_c_462_n 0.0121126f $X=0.545 $Y=2.505 $X2=0
+ $Y2=0
cc_130 N_A_84_259#_M1010_g N_VPWR_c_461_n 0.0135501f $X=0.545 $Y=2.505 $X2=0
+ $Y2=0
cc_131 N_A_84_259#_M1010_g N_VPWR_c_467_n 0.00717535f $X=0.545 $Y=2.505 $X2=0
+ $Y2=0
cc_132 N_A_84_259#_c_82_n A_306_401# 6.88945e-19 $X=1.505 $Y=2.065 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_84_259#_c_112_p A_306_401# 0.00598648f $X=2.16 $Y=2.15 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A_84_259#_c_81_n N_VGND_M1007_d 0.00182157f $X=1.505 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_84_259#_c_146_p N_VGND_M1007_d 0.00309271f $X=1.59 $Y=0.43 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_84_259#_c_76_n N_VGND_c_506_n 5.79521e-19 $X=0.545 $Y=1.42 $X2=0
+ $Y2=0
cc_137 N_A_84_259#_M1001_g N_VGND_c_506_n 0.002112f $X=0.5 $Y=0.495 $X2=0 $Y2=0
cc_138 N_A_84_259#_M1007_g N_VGND_c_506_n 0.0134154f $X=0.86 $Y=0.495 $X2=0
+ $Y2=0
cc_139 N_A_84_259#_c_80_n N_VGND_c_506_n 0.0275493f $X=1.42 $Y=1.07 $X2=0 $Y2=0
cc_140 N_A_84_259#_c_81_n N_VGND_c_506_n 0.0154042f $X=1.505 $Y=0.905 $X2=0
+ $Y2=0
cc_141 N_A_84_259#_c_146_p N_VGND_c_506_n 0.0138719f $X=1.59 $Y=0.43 $X2=0 $Y2=0
cc_142 N_A_84_259#_c_84_n N_VGND_c_507_n 0.00263454f $X=2.66 $Y=0.495 $X2=0
+ $Y2=0
cc_143 N_A_84_259#_M1001_g N_VGND_c_508_n 0.00502664f $X=0.5 $Y=0.495 $X2=0
+ $Y2=0
cc_144 N_A_84_259#_M1007_g N_VGND_c_508_n 0.00445056f $X=0.86 $Y=0.495 $X2=0
+ $Y2=0
cc_145 N_A_84_259#_c_146_p N_VGND_c_509_n 0.00644478f $X=1.59 $Y=0.43 $X2=0
+ $Y2=0
cc_146 N_A_84_259#_c_96_p N_VGND_c_509_n 0.0457842f $X=2.495 $Y=0.535 $X2=0
+ $Y2=0
cc_147 N_A_84_259#_M1001_g N_VGND_c_511_n 0.0100646f $X=0.5 $Y=0.495 $X2=0 $Y2=0
cc_148 N_A_84_259#_M1007_g N_VGND_c_511_n 0.00796275f $X=0.86 $Y=0.495 $X2=0
+ $Y2=0
cc_149 N_A_84_259#_c_146_p N_VGND_c_511_n 0.00629747f $X=1.59 $Y=0.43 $X2=0
+ $Y2=0
cc_150 N_A_84_259#_c_96_p N_VGND_c_511_n 0.042531f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_151 N_A_84_259#_c_96_p A_349_57# 0.0062275f $X=2.495 $Y=0.535 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_182_303#_M1011_g N_A1_M1003_g 0.0467335f $X=1.405 $Y=2.505 $X2=0
+ $Y2=0
cc_153 N_A_182_303#_c_204_n N_A1_M1003_g 0.0177156f $X=3.585 $Y=2.5 $X2=0 $Y2=0
cc_154 N_A_182_303#_c_166_n N_A1_c_269_n 3.65464e-19 $X=1.405 $Y=1.68 $X2=0
+ $Y2=0
cc_155 N_A_182_303#_c_204_n N_A1_c_269_n 0.0087799f $X=3.585 $Y=2.5 $X2=0 $Y2=0
cc_156 N_A_182_303#_c_166_n N_A1_c_270_n 0.0467335f $X=1.405 $Y=1.68 $X2=0 $Y2=0
cc_157 N_A_182_303#_c_164_n N_A0_c_335_n 0.0214344f $X=1.67 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_182_303#_c_204_n N_A0_M1000_g 0.0208309f $X=3.585 $Y=2.5 $X2=0 $Y2=0
cc_159 N_A_182_303#_c_163_n A0 2.46466e-19 $X=1.455 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A_182_303#_c_167_n A0 4.91884e-19 $X=1.67 $Y=0.855 $X2=0 $Y2=0
cc_161 N_A_182_303#_c_163_n N_A0_c_340_n 0.00498062f $X=1.455 $Y=1.515 $X2=0
+ $Y2=0
cc_162 N_A_182_303#_c_167_n N_A0_c_340_n 0.0214344f $X=1.67 $Y=0.855 $X2=0 $Y2=0
cc_163 N_A_182_303#_c_204_n N_S_M1005_g 0.020832f $X=3.585 $Y=2.5 $X2=0 $Y2=0
cc_164 N_A_182_303#_c_175_n N_S_M1005_g 7.25173e-19 $X=3.75 $Y=2.155 $X2=0 $Y2=0
cc_165 N_A_182_303#_c_176_n N_S_M1005_g 0.00111412f $X=3.75 $Y=2.415 $X2=0 $Y2=0
cc_166 N_A_182_303#_c_177_n N_S_M1005_g 6.30887e-19 $X=3.75 $Y=2.86 $X2=0 $Y2=0
cc_167 N_A_182_303#_c_204_n N_S_M1013_g 0.0170744f $X=3.585 $Y=2.5 $X2=0 $Y2=0
cc_168 N_A_182_303#_c_175_n N_S_M1013_g 0.00456803f $X=3.75 $Y=2.155 $X2=0 $Y2=0
cc_169 N_A_182_303#_c_176_n N_S_M1013_g 0.00523018f $X=3.75 $Y=2.415 $X2=0 $Y2=0
cc_170 N_A_182_303#_c_177_n N_S_M1013_g 0.00857868f $X=3.75 $Y=2.86 $X2=0 $Y2=0
cc_171 N_A_182_303#_c_180_n N_S_M1013_g 3.84191e-19 $X=3.75 $Y=2.5 $X2=0 $Y2=0
cc_172 N_A_182_303#_c_170_n N_S_M1008_g 0.00125204f $X=4.38 $Y=0.495 $X2=0 $Y2=0
cc_173 N_A_182_303#_c_169_n N_S_M1009_g 0.0357634f $X=4.46 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_182_303#_c_170_n N_S_M1009_g 0.0101221f $X=4.38 $Y=0.495 $X2=0 $Y2=0
cc_175 N_A_182_303#_c_204_n S 0.0173521f $X=3.585 $Y=2.5 $X2=0 $Y2=0
cc_176 N_A_182_303#_c_175_n S 0.0265437f $X=3.75 $Y=2.155 $X2=0 $Y2=0
cc_177 N_A_182_303#_c_178_n S 0.0201206f $X=4.375 $Y=2.07 $X2=0 $Y2=0
cc_178 N_A_182_303#_c_169_n S 0.0250954f $X=4.46 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_182_303#_c_204_n N_S_c_383_n 0.00159567f $X=3.585 $Y=2.5 $X2=0 $Y2=0
cc_180 N_A_182_303#_c_175_n N_S_c_383_n 0.00814315f $X=3.75 $Y=2.155 $X2=0 $Y2=0
cc_181 N_A_182_303#_c_178_n N_S_c_383_n 0.0090573f $X=4.375 $Y=2.07 $X2=0 $Y2=0
cc_182 N_A_182_303#_c_207_n N_X_c_441_n 0.00244423f $X=1.24 $Y=2.5 $X2=0 $Y2=0
cc_183 N_A_182_303#_c_165_n X 9.75956e-19 $X=1.28 $Y=1.68 $X2=0 $Y2=0
cc_184 N_A_182_303#_c_168_n X 0.0317824f $X=1.075 $Y=1.68 $X2=0 $Y2=0
cc_185 N_A_182_303#_c_207_n X 0.00401418f $X=1.24 $Y=2.5 $X2=0 $Y2=0
cc_186 N_A_182_303#_c_168_n N_VPWR_M1010_d 0.0109704f $X=1.075 $Y=1.68 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_182_303#_c_207_n N_VPWR_M1010_d 0.00990429f $X=1.24 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_182_303#_c_204_n N_VPWR_M1005_d 0.00482647f $X=3.585 $Y=2.5 $X2=0
+ $Y2=0
cc_189 N_A_182_303#_M1011_g N_VPWR_c_462_n 0.00819181f $X=1.405 $Y=2.505 $X2=0
+ $Y2=0
cc_190 N_A_182_303#_c_207_n N_VPWR_c_462_n 0.00524842f $X=1.24 $Y=2.5 $X2=0
+ $Y2=0
cc_191 N_A_182_303#_c_204_n N_VPWR_c_463_n 0.0156967f $X=3.585 $Y=2.5 $X2=0
+ $Y2=0
cc_192 N_A_182_303#_c_177_n N_VPWR_c_463_n 0.0171316f $X=3.75 $Y=2.86 $X2=0
+ $Y2=0
cc_193 N_A_182_303#_M1011_g N_VPWR_c_464_n 0.00614491f $X=1.405 $Y=2.505 $X2=0
+ $Y2=0
cc_194 N_A_182_303#_c_204_n N_VPWR_c_464_n 0.0216386f $X=3.585 $Y=2.5 $X2=0
+ $Y2=0
cc_195 N_A_182_303#_c_207_n N_VPWR_c_464_n 0.00394033f $X=1.24 $Y=2.5 $X2=0
+ $Y2=0
cc_196 N_A_182_303#_c_204_n N_VPWR_c_465_n 0.00254828f $X=3.585 $Y=2.5 $X2=0
+ $Y2=0
cc_197 N_A_182_303#_c_177_n N_VPWR_c_465_n 0.0177662f $X=3.75 $Y=2.86 $X2=0
+ $Y2=0
cc_198 N_A_182_303#_M1011_g N_VPWR_c_461_n 0.00851092f $X=1.405 $Y=2.505 $X2=0
+ $Y2=0
cc_199 N_A_182_303#_c_204_n N_VPWR_c_461_n 0.0482726f $X=3.585 $Y=2.5 $X2=0
+ $Y2=0
cc_200 N_A_182_303#_c_207_n N_VPWR_c_461_n 0.00772312f $X=1.24 $Y=2.5 $X2=0
+ $Y2=0
cc_201 N_A_182_303#_c_177_n N_VPWR_c_461_n 0.0123184f $X=3.75 $Y=2.86 $X2=0
+ $Y2=0
cc_202 N_A_182_303#_c_204_n A_306_401# 0.00376622f $X=3.585 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_182_303#_c_204_n A_518_401# 0.00693206f $X=3.585 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_182_303#_c_164_n N_VGND_c_506_n 0.00433746f $X=1.67 $Y=0.78 $X2=0
+ $Y2=0
cc_205 N_A_182_303#_c_170_n N_VGND_c_507_n 0.0153904f $X=4.38 $Y=0.495 $X2=0
+ $Y2=0
cc_206 N_A_182_303#_c_164_n N_VGND_c_509_n 0.00341756f $X=1.67 $Y=0.78 $X2=0
+ $Y2=0
cc_207 N_A_182_303#_c_167_n N_VGND_c_509_n 0.00120198f $X=1.67 $Y=0.855 $X2=0
+ $Y2=0
cc_208 N_A_182_303#_c_170_n N_VGND_c_510_n 0.0217285f $X=4.38 $Y=0.495 $X2=0
+ $Y2=0
cc_209 N_A_182_303#_c_164_n N_VGND_c_511_n 0.00534735f $X=1.67 $Y=0.78 $X2=0
+ $Y2=0
cc_210 N_A_182_303#_c_167_n N_VGND_c_511_n 0.00108233f $X=1.67 $Y=0.855 $X2=0
+ $Y2=0
cc_211 N_A_182_303#_c_170_n N_VGND_c_511_n 0.0125175f $X=4.38 $Y=0.495 $X2=0
+ $Y2=0
cc_212 N_A1_M1004_g N_A0_c_335_n 0.00748711f $X=2.875 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A1_c_269_n N_A0_c_336_n 0.00998423f $X=2.495 $Y=1.68 $X2=0 $Y2=0
cc_214 N_A1_c_270_n N_A0_c_336_n 0.018117f $X=1.935 $Y=1.68 $X2=0 $Y2=0
cc_215 N_A1_c_271_n N_A0_c_336_n 0.00417995f $X=2.58 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A1_M1003_g N_A0_M1000_g 0.0441834f $X=1.895 $Y=2.505 $X2=0 $Y2=0
cc_217 N_A1_c_269_n N_A0_M1000_g 0.0161793f $X=2.495 $Y=1.68 $X2=0 $Y2=0
cc_218 N_A1_c_271_n N_A0_c_338_n 0.00980278f $X=2.58 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A1_M1004_g A0 5.76477e-19 $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_220 N_A1_c_269_n A0 0.0141301f $X=2.495 $Y=1.68 $X2=0 $Y2=0
cc_221 N_A1_c_270_n A0 4.99128e-19 $X=1.935 $Y=1.68 $X2=0 $Y2=0
cc_222 N_A1_c_273_n A0 0.0193848f $X=2.665 $Y=1.07 $X2=0 $Y2=0
cc_223 N_A1_M1004_g N_A0_c_340_n 0.00198995f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_224 N_A1_c_269_n N_A0_c_340_n 0.00230328f $X=2.495 $Y=1.68 $X2=0 $Y2=0
cc_225 N_A1_c_270_n N_A0_c_340_n 0.00364645f $X=1.935 $Y=1.68 $X2=0 $Y2=0
cc_226 N_A1_c_273_n N_A0_c_340_n 0.00524242f $X=2.665 $Y=1.07 $X2=0 $Y2=0
cc_227 N_A1_c_274_n N_A0_c_340_n 0.0146469f $X=2.895 $Y=1.07 $X2=0 $Y2=0
cc_228 N_A1_M1004_g N_S_M1002_g 0.0218147f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_229 N_A1_c_271_n N_S_M1002_g 0.00505851f $X=2.58 $Y=1.515 $X2=0 $Y2=0
cc_230 N_A1_c_274_n N_S_M1002_g 0.0162467f $X=2.895 $Y=1.07 $X2=0 $Y2=0
cc_231 A1 N_S_M1002_g 0.00697836f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_232 N_A1_c_276_n N_S_M1002_g 0.01014f $X=3.12 $Y=0.905 $X2=0 $Y2=0
cc_233 N_A1_c_269_n S 0.0246693f $X=2.495 $Y=1.68 $X2=0 $Y2=0
cc_234 N_A1_c_271_n S 0.00294774f $X=2.58 $Y=1.515 $X2=0 $Y2=0
cc_235 N_A1_c_272_n S 0.00908682f $X=3.005 $Y=1.07 $X2=0 $Y2=0
cc_236 N_A1_c_274_n S 7.21519e-19 $X=2.895 $Y=1.07 $X2=0 $Y2=0
cc_237 N_A1_c_276_n S 0.0147363f $X=3.12 $Y=0.905 $X2=0 $Y2=0
cc_238 N_A1_c_269_n N_S_c_383_n 0.00327902f $X=2.495 $Y=1.68 $X2=0 $Y2=0
cc_239 N_A1_c_271_n N_S_c_383_n 2.73658e-19 $X=2.58 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A1_c_272_n N_S_c_383_n 7.9666e-19 $X=3.005 $Y=1.07 $X2=0 $Y2=0
cc_241 N_A1_c_274_n N_S_c_383_n 0.0132474f $X=2.895 $Y=1.07 $X2=0 $Y2=0
cc_242 N_A1_c_276_n N_S_c_383_n 0.00456286f $X=3.12 $Y=0.905 $X2=0 $Y2=0
cc_243 N_A1_M1003_g N_VPWR_c_464_n 0.00614491f $X=1.895 $Y=2.505 $X2=0 $Y2=0
cc_244 N_A1_M1003_g N_VPWR_c_461_n 0.00831366f $X=1.895 $Y=2.505 $X2=0 $Y2=0
cc_245 N_A1_M1004_g N_VGND_c_507_n 0.00147238f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_246 A1 N_VGND_c_507_n 0.0197815f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_247 N_A1_M1004_g N_VGND_c_509_n 0.00503642f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_248 A1 N_VGND_c_509_n 0.00719474f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_249 N_A1_M1004_g N_VGND_c_511_n 0.0101211f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_250 A1 N_VGND_c_511_n 0.0079425f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_251 A1 A_590_57# 0.00875576f $X=3.035 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_252 N_A0_M1000_g N_S_M1005_g 0.049115f $X=2.465 $Y=2.505 $X2=0 $Y2=0
cc_253 N_A0_c_336_n S 3.52248e-19 $X=2.465 $Y=1.6 $X2=0 $Y2=0
cc_254 N_A0_c_336_n N_S_c_383_n 0.049115f $X=2.465 $Y=1.6 $X2=0 $Y2=0
cc_255 N_A0_M1000_g N_VPWR_c_463_n 0.00172228f $X=2.465 $Y=2.505 $X2=0 $Y2=0
cc_256 N_A0_M1000_g N_VPWR_c_464_n 0.00614491f $X=2.465 $Y=2.505 $X2=0 $Y2=0
cc_257 N_A0_M1000_g N_VPWR_c_461_n 0.00831366f $X=2.465 $Y=2.505 $X2=0 $Y2=0
cc_258 N_A0_c_335_n N_VGND_c_509_n 0.00341756f $X=2.06 $Y=0.815 $X2=0 $Y2=0
cc_259 N_A0_c_335_n N_VGND_c_511_n 0.0053421f $X=2.06 $Y=0.815 $X2=0 $Y2=0
cc_260 N_S_M1005_g N_VPWR_c_463_n 0.00980665f $X=2.955 $Y=2.505 $X2=0 $Y2=0
cc_261 N_S_M1013_g N_VPWR_c_463_n 0.0107419f $X=3.485 $Y=2.505 $X2=0 $Y2=0
cc_262 N_S_M1005_g N_VPWR_c_464_n 0.00552397f $X=2.955 $Y=2.505 $X2=0 $Y2=0
cc_263 N_S_M1013_g N_VPWR_c_465_n 0.00543943f $X=3.485 $Y=2.505 $X2=0 $Y2=0
cc_264 N_S_M1005_g N_VPWR_c_461_n 0.00698489f $X=2.955 $Y=2.505 $X2=0 $Y2=0
cc_265 N_S_M1013_g N_VPWR_c_461_n 0.00736963f $X=3.485 $Y=2.505 $X2=0 $Y2=0
cc_266 N_S_M1002_g N_VGND_c_507_n 0.0125679f $X=3.375 $Y=0.495 $X2=0 $Y2=0
cc_267 N_S_M1008_g N_VGND_c_507_n 0.0134712f $X=3.805 $Y=0.495 $X2=0 $Y2=0
cc_268 N_S_M1009_g N_VGND_c_507_n 0.002112f $X=4.165 $Y=0.495 $X2=0 $Y2=0
cc_269 N_S_M1002_g N_VGND_c_509_n 0.00445056f $X=3.375 $Y=0.495 $X2=0 $Y2=0
cc_270 N_S_M1008_g N_VGND_c_510_n 0.00445056f $X=3.805 $Y=0.495 $X2=0 $Y2=0
cc_271 N_S_M1009_g N_VGND_c_510_n 0.00502664f $X=4.165 $Y=0.495 $X2=0 $Y2=0
cc_272 N_S_M1002_g N_VGND_c_511_n 0.00822633f $X=3.375 $Y=0.495 $X2=0 $Y2=0
cc_273 N_S_M1008_g N_VGND_c_511_n 0.00796275f $X=3.805 $Y=0.495 $X2=0 $Y2=0
cc_274 N_S_M1009_g N_VGND_c_511_n 0.010132f $X=4.165 $Y=0.495 $X2=0 $Y2=0
cc_275 N_X_c_441_n N_VPWR_c_462_n 0.0171316f $X=0.28 $Y=2.86 $X2=0 $Y2=0
cc_276 N_X_c_441_n N_VPWR_c_461_n 0.0123184f $X=0.28 $Y=2.86 $X2=0 $Y2=0
cc_277 N_X_c_441_n N_VPWR_c_467_n 0.0177662f $X=0.28 $Y=2.86 $X2=0 $Y2=0
cc_278 X N_VGND_c_506_n 0.0154081f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_279 X N_VGND_c_508_n 0.0223692f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_280 X N_VGND_c_511_n 0.0127743f $X=0.155 $Y=0.47 $X2=0 $Y2=0
