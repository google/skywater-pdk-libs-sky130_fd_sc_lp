* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 VGND D a_41_464# VNB nshort w=420000u l=150000u
+  ad=7.791e+11p pd=7.13e+06u as=1.113e+11p ps=1.37e+06u
M1001 VPWR a_249_70# a_371_473# VPB phighvt w=640000u l=150000u
+  ad=1.7295e+12p pd=1.213e+07u as=1.696e+11p ps=1.81e+06u
M1002 a_623_473# a_41_464# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1003 a_587_47# a_41_464# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_809_21# a_659_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1005 a_659_47# a_371_473# a_587_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1006 a_1056_73# a_659_47# a_809_21# VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=2.226e+11p ps=2.21e+06u
M1007 a_659_47# a_249_70# a_623_473# VPB phighvt w=640000u l=150000u
+  ad=2.158e+11p pd=2.03e+06u as=0p ps=0u
M1008 VPWR a_809_21# a_800_473# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 a_767_47# a_249_70# a_659_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VGND a_809_21# a_767_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_809_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1012 VGND a_249_70# a_371_473# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1013 a_249_70# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1014 a_249_70# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=0p ps=0u
M1015 VPWR D a_41_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1016 VPWR RESET_B a_809_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_800_473# a_371_473# a_659_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_809_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1019 VGND RESET_B a_1056_73# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
