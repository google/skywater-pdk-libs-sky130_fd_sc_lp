* File: sky130_fd_sc_lp__a221o_0.spice
* Created: Wed Sep  2 09:21:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221o_0.pex.spice"
.subckt sky130_fd_sc_lp__a221o_0  VNB VPB A2 A1 B1 B2 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_72_312#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1113 PD=0.84 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1009 A_246_47# N_A2_M1009_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=21.42 M=1 R=2.8 SA=75000.8 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_72_312#_M1005_d N_A1_M1005_g A_246_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1323 AS=0.0441 PD=1.05 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 A_474_47# N_B1_M1004_g N_A_72_312#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1323 PD=0.63 PS=1.05 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_B2_M1006_g A_474_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=21.42 NRS=14.28 M=1 R=2.8 SA=75002.3 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_72_312#_M1010_d N_C1_M1010_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=9.996 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_72_312#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.1696 PD=0.94 PS=1.81 NRD=6.1464 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_216_484#_M1001_d N_A2_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.096 PD=0.92 PS=0.94 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_216_484#_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_216_484#_M1002_d N_B1_M1002_g N_A_409_429#_M1002_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=6.1464 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 N_A_409_429#_M1008_d N_B2_M1008_g N_A_216_484#_M1002_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1011 N_A_72_312#_M1011_d N_C1_M1011_g N_A_409_429#_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.112 PD=1.81 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a221o_0.pxi.spice"
*
.ends
*
*
