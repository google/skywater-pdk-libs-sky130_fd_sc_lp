* File: sky130_fd_sc_lp__a211o_lp.pxi.spice
* Created: Fri Aug 28 09:47:55 2020
* 
x_PM_SKY130_FD_SC_LP__A211O_LP%A1 N_A1_c_70_n N_A1_M1000_g N_A1_M1001_g A1 A1
+ N_A1_c_72_n PM_SKY130_FD_SC_LP__A211O_LP%A1
x_PM_SKY130_FD_SC_LP__A211O_LP%A2 N_A2_M1012_g N_A2_c_101_n N_A2_M1009_g
+ N_A2_c_105_n A2 A2 N_A2_c_103_n PM_SKY130_FD_SC_LP__A211O_LP%A2
x_PM_SKY130_FD_SC_LP__A211O_LP%B1 N_B1_c_138_n N_B1_M1002_g N_B1_c_142_n
+ N_B1_M1005_g N_B1_c_139_n N_B1_M1003_g N_B1_c_140_n B1 B1 N_B1_c_141_n
+ PM_SKY130_FD_SC_LP__A211O_LP%B1
x_PM_SKY130_FD_SC_LP__A211O_LP%C1 N_C1_M1011_g N_C1_M1007_g N_C1_M1004_g
+ N_C1_c_188_n N_C1_c_192_n C1 C1 N_C1_c_190_n PM_SKY130_FD_SC_LP__A211O_LP%C1
x_PM_SKY130_FD_SC_LP__A211O_LP%A_43_57# N_A_43_57#_M1001_s N_A_43_57#_M1003_d
+ N_A_43_57#_M1011_d N_A_43_57#_c_236_n N_A_43_57#_M1008_g N_A_43_57#_M1006_g
+ N_A_43_57#_c_238_n N_A_43_57#_M1010_g N_A_43_57#_c_239_n N_A_43_57#_c_240_n
+ N_A_43_57#_c_241_n N_A_43_57#_c_249_n N_A_43_57#_c_250_n N_A_43_57#_c_251_n
+ N_A_43_57#_c_242_n N_A_43_57#_c_283_n N_A_43_57#_c_243_n N_A_43_57#_c_244_n
+ N_A_43_57#_c_245_n N_A_43_57#_c_246_n N_A_43_57#_c_247_n
+ PM_SKY130_FD_SC_LP__A211O_LP%A_43_57#
x_PM_SKY130_FD_SC_LP__A211O_LP%A_29_409# N_A_29_409#_M1000_s N_A_29_409#_M1009_d
+ N_A_29_409#_c_330_n N_A_29_409#_c_331_n N_A_29_409#_c_332_n
+ N_A_29_409#_c_333_n PM_SKY130_FD_SC_LP__A211O_LP%A_29_409#
x_PM_SKY130_FD_SC_LP__A211O_LP%VPWR N_VPWR_M1000_d N_VPWR_M1006_s N_VPWR_c_361_n
+ N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n VPWR N_VPWR_c_365_n
+ N_VPWR_c_360_n N_VPWR_c_367_n PM_SKY130_FD_SC_LP__A211O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A211O_LP%X N_X_M1010_d N_X_M1006_d X X X X X X X
+ PM_SKY130_FD_SC_LP__A211O_LP%X
x_PM_SKY130_FD_SC_LP__A211O_LP%VGND N_VGND_M1012_d N_VGND_M1004_d N_VGND_c_415_n
+ N_VGND_c_416_n VGND N_VGND_c_417_n N_VGND_c_418_n N_VGND_c_419_n
+ N_VGND_c_420_n N_VGND_c_421_n N_VGND_c_422_n PM_SKY130_FD_SC_LP__A211O_LP%VGND
cc_1 VNB N_A1_c_70_n 0.0876617f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.75
cc_2 VNB N_A1_M1001_g 0.032957f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.495
cc_3 VNB N_A1_c_72_n 0.0322022f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.12
cc_4 VNB N_A2_M1012_g 0.0343873f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.545
cc_5 VNB N_A2_c_101_n 0.020484f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.495
cc_6 VNB A2 0.00567617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A2_c_103_n 0.0190177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_138_n 0.0138865f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.75
cc_9 VNB N_B1_c_139_n 0.0137713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_140_n 0.018608f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.12
cc_11 VNB N_B1_c_141_n 0.0527613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C1_M1007_g 0.0310797f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.495
cc_13 VNB N_C1_M1004_g 0.0310567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C1_c_188_n 0.0235666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB C1 0.00414624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_c_190_n 0.0249538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_43_57#_c_236_n 0.0158686f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_A_43_57#_M1006_g 0.0127908f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.12
cc_19 VNB N_A_43_57#_c_238_n 0.0198912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_43_57#_c_239_n 0.0134883f $X=-0.19 $Y=-0.245 $X2=0.305 $Y2=1.665
cc_21 VNB N_A_43_57#_c_240_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_43_57#_c_241_n 0.0181694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_43_57#_c_242_n 8.26572e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_43_57#_c_243_n 0.00291709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_43_57#_c_244_n 0.0330653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_43_57#_c_245_n 0.00927711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_43_57#_c_246_n 0.0796389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_43_57#_c_247_n 0.00467522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_360_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB X 0.0587996f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.495
cc_31 VNB N_VGND_c_415_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_32 VNB N_VGND_c_416_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.12
cc_33 VNB N_VGND_c_417_n 0.0290631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_418_n 0.0352526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_419_n 0.0275168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_420_n 0.231352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_421_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_422_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A1_c_70_n 0.00680514f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.75
cc_40 VPB N_A1_M1000_g 0.0452126f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.545
cc_41 VPB N_A1_c_72_n 0.00794424f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.12
cc_42 VPB N_A2_M1009_g 0.0294655f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_43 VPB N_A2_c_105_n 0.0158437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB A2 0.00243683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B1_c_142_n 0.0138848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B1_M1005_g 0.029037f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.495
cc_47 VPB B1 0.00195814f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=1.295
cc_48 VPB N_B1_c_141_n 0.00134252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_C1_M1011_g 0.0337655f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.545
cc_50 VPB N_C1_c_192_n 0.014908f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=1.665
cc_51 VPB C1 0.00296927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_C1_c_190_n 0.00145704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_43_57#_M1006_g 0.0504419f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.12
cc_54 VPB N_A_43_57#_c_249_n 0.0111748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_43_57#_c_250_n 0.0184783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_43_57#_c_251_n 0.00487352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_43_57#_c_243_n 0.00920236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_29_409#_c_330_n 0.035517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_29_409#_c_331_n 0.0164712f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.12
cc_60 VPB N_A_29_409#_c_332_n 0.0095886f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.12
cc_61 VPB N_A_29_409#_c_333_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_361_n 0.00416786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_362_n 0.0104514f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.12
cc_64 VPB N_VPWR_c_363_n 0.0533915f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=1.295
cc_65 VPB N_VPWR_c_364_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_365_n 0.0192431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_360_n 0.077036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_367_n 0.0247306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB X 0.0573842f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.495
cc_70 N_A1_M1001_g N_A2_M1012_g 0.0388128f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_71 N_A1_c_72_n N_A2_M1012_g 0.00261876f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_72 N_A1_c_70_n N_A2_c_101_n 0.00686598f $X=0.555 $Y=1.75 $X2=0 $Y2=0
cc_73 N_A1_M1000_g N_A2_M1009_g 0.0252746f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_74 N_A1_M1000_g N_A2_c_105_n 0.00686598f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_75 N_A1_c_70_n A2 0.00276674f $X=0.555 $Y=1.75 $X2=0 $Y2=0
cc_76 N_A1_c_72_n A2 0.0213341f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_77 N_A1_c_70_n N_A2_c_103_n 0.0388128f $X=0.555 $Y=1.75 $X2=0 $Y2=0
cc_78 N_A1_c_70_n N_A_43_57#_c_244_n 0.00319779f $X=0.555 $Y=1.75 $X2=0 $Y2=0
cc_79 N_A1_M1001_g N_A_43_57#_c_244_n 0.0263936f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_80 N_A1_c_72_n N_A_43_57#_c_244_n 0.0227324f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_81 N_A1_M1000_g N_A_29_409#_c_330_n 0.0160648f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_82 N_A1_M1000_g N_A_29_409#_c_331_n 0.0240121f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_83 N_A1_c_72_n N_A_29_409#_c_331_n 0.0016489f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_84 N_A1_c_70_n N_A_29_409#_c_332_n 0.00150166f $X=0.555 $Y=1.75 $X2=0 $Y2=0
cc_85 N_A1_M1000_g N_A_29_409#_c_332_n 0.00130637f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_86 N_A1_c_72_n N_A_29_409#_c_332_n 0.0239369f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_87 N_A1_M1000_g N_A_29_409#_c_333_n 8.99696e-19 $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_88 N_A1_M1000_g N_VPWR_c_361_n 0.017429f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_89 N_A1_M1000_g N_VPWR_c_360_n 0.0140911f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_90 N_A1_M1000_g N_VPWR_c_367_n 0.00769046f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_91 N_A1_M1001_g N_VGND_c_415_n 0.00171633f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_92 N_A1_M1001_g N_VGND_c_417_n 0.00366349f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_93 N_A1_M1001_g N_VGND_c_420_n 0.00586405f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_94 N_A2_M1012_g N_B1_c_138_n 0.0191069f $X=0.965 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A2_c_101_n N_B1_c_142_n 0.0176675f $X=1.075 $Y=1.655 $X2=0 $Y2=0
cc_96 N_A2_M1009_g N_B1_M1005_g 0.0174755f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_97 A2 B1 0.0503477f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_98 N_A2_c_103_n B1 7.64192e-19 $X=1.095 $Y=1.335 $X2=0 $Y2=0
cc_99 N_A2_M1012_g N_B1_c_141_n 0.00751394f $X=0.965 $Y=0.495 $X2=0 $Y2=0
cc_100 A2 N_B1_c_141_n 0.0041215f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A2_c_103_n N_B1_c_141_n 0.0176675f $X=1.095 $Y=1.335 $X2=0 $Y2=0
cc_102 N_A2_M1012_g N_A_43_57#_c_239_n 0.0125608f $X=0.965 $Y=0.495 $X2=0 $Y2=0
cc_103 A2 N_A_43_57#_c_239_n 0.0291068f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A2_c_103_n N_A_43_57#_c_239_n 0.00151167f $X=1.095 $Y=1.335 $X2=0 $Y2=0
cc_105 N_A2_M1012_g N_A_43_57#_c_244_n 0.00417832f $X=0.965 $Y=0.495 $X2=0 $Y2=0
cc_106 N_A2_M1009_g N_A_29_409#_c_330_n 8.56315e-19 $X=1.135 $Y=2.545 $X2=0
+ $Y2=0
cc_107 N_A2_M1009_g N_A_29_409#_c_331_n 0.0198967f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_108 N_A2_c_105_n N_A_29_409#_c_331_n 0.00222631f $X=1.075 $Y=1.84 $X2=0 $Y2=0
cc_109 A2 N_A_29_409#_c_331_n 0.0292218f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A2_M1009_g N_A_29_409#_c_333_n 0.0141925f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_111 N_A2_M1009_g N_VPWR_c_361_n 0.0029541f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_112 N_A2_M1009_g N_VPWR_c_363_n 0.0086001f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_113 N_A2_M1009_g N_VPWR_c_360_n 0.0156763f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_114 N_A2_M1012_g N_VGND_c_415_n 0.0102775f $X=0.965 $Y=0.495 $X2=0 $Y2=0
cc_115 N_A2_M1012_g N_VGND_c_417_n 0.00445056f $X=0.965 $Y=0.495 $X2=0 $Y2=0
cc_116 N_A2_M1012_g N_VGND_c_420_n 0.00426841f $X=0.965 $Y=0.495 $X2=0 $Y2=0
cc_117 N_B1_M1005_g N_C1_M1011_g 0.0632364f $X=1.665 $Y=2.545 $X2=0 $Y2=0
cc_118 N_B1_c_139_n N_C1_M1007_g 0.0303431f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_119 B1 N_C1_c_188_n 8.14382e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B1_c_141_n N_C1_c_188_n 0.0177665f $X=1.665 $Y=1.335 $X2=0 $Y2=0
cc_121 B1 C1 0.0447196f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_c_141_n C1 0.00410965f $X=1.665 $Y=1.335 $X2=0 $Y2=0
cc_123 N_B1_c_142_n N_C1_c_190_n 0.0177665f $X=1.665 $Y=1.84 $X2=0 $Y2=0
cc_124 N_B1_c_140_n N_A_43_57#_c_239_n 0.0199287f $X=1.755 $Y=0.855 $X2=0 $Y2=0
cc_125 B1 N_A_43_57#_c_239_n 0.0220537f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B1_c_141_n N_A_43_57#_c_239_n 0.00690231f $X=1.665 $Y=1.335 $X2=0 $Y2=0
cc_127 N_B1_c_138_n N_A_43_57#_c_240_n 0.00171786f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_128 N_B1_c_139_n N_A_43_57#_c_240_n 0.0100195f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_129 N_B1_c_140_n N_A_43_57#_c_240_n 0.00230187f $X=1.755 $Y=0.855 $X2=0 $Y2=0
cc_130 N_B1_M1005_g N_A_43_57#_c_249_n 0.00376238f $X=1.665 $Y=2.545 $X2=0 $Y2=0
cc_131 N_B1_M1005_g N_A_43_57#_c_251_n 7.25172e-19 $X=1.665 $Y=2.545 $X2=0 $Y2=0
cc_132 N_B1_c_140_n N_A_43_57#_c_245_n 0.00156724f $X=1.755 $Y=0.855 $X2=0 $Y2=0
cc_133 B1 N_A_43_57#_c_245_n 0.00193735f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B1_c_141_n N_A_43_57#_c_245_n 0.00119316f $X=1.665 $Y=1.335 $X2=0 $Y2=0
cc_135 N_B1_c_142_n N_A_29_409#_c_331_n 3.02817e-19 $X=1.665 $Y=1.84 $X2=0 $Y2=0
cc_136 N_B1_M1005_g N_A_29_409#_c_331_n 0.00438558f $X=1.665 $Y=2.545 $X2=0
+ $Y2=0
cc_137 B1 N_A_29_409#_c_331_n 0.00534367f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B1_M1005_g N_A_29_409#_c_333_n 0.0181312f $X=1.665 $Y=2.545 $X2=0 $Y2=0
cc_139 N_B1_M1005_g N_VPWR_c_363_n 0.0086001f $X=1.665 $Y=2.545 $X2=0 $Y2=0
cc_140 N_B1_M1005_g N_VPWR_c_360_n 0.0157977f $X=1.665 $Y=2.545 $X2=0 $Y2=0
cc_141 N_B1_c_138_n N_VGND_c_415_n 0.0105659f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_142 N_B1_c_139_n N_VGND_c_415_n 0.00188065f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_143 N_B1_c_138_n N_VGND_c_418_n 0.00445056f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_144 N_B1_c_139_n N_VGND_c_418_n 0.00502664f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_145 N_B1_c_140_n N_VGND_c_418_n 5.84996e-19 $X=1.755 $Y=0.855 $X2=0 $Y2=0
cc_146 N_B1_c_138_n N_VGND_c_420_n 0.00418511f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_147 N_B1_c_139_n N_VGND_c_420_n 0.00562693f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_148 N_B1_c_140_n N_VGND_c_420_n 7.94744e-19 $X=1.755 $Y=0.855 $X2=0 $Y2=0
cc_149 N_C1_M1004_g N_A_43_57#_c_236_n 0.0147173f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_150 N_C1_M1007_g N_A_43_57#_c_240_n 0.0111815f $X=2.185 $Y=0.495 $X2=0 $Y2=0
cc_151 N_C1_M1004_g N_A_43_57#_c_240_n 0.00192036f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_152 N_C1_M1007_g N_A_43_57#_c_241_n 0.00807925f $X=2.185 $Y=0.495 $X2=0 $Y2=0
cc_153 N_C1_M1004_g N_A_43_57#_c_241_n 0.014987f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_154 N_C1_c_188_n N_A_43_57#_c_241_n 2.06387e-19 $X=2.545 $Y=1.245 $X2=0 $Y2=0
cc_155 C1 N_A_43_57#_c_241_n 0.0196738f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_C1_M1011_g N_A_43_57#_c_249_n 0.0182913f $X=2.195 $Y=2.545 $X2=0 $Y2=0
cc_157 N_C1_M1011_g N_A_43_57#_c_251_n 0.00468955f $X=2.195 $Y=2.545 $X2=0 $Y2=0
cc_158 N_C1_c_188_n N_A_43_57#_c_251_n 0.00617539f $X=2.545 $Y=1.245 $X2=0 $Y2=0
cc_159 N_C1_c_192_n N_A_43_57#_c_251_n 6.13648e-19 $X=2.235 $Y=1.84 $X2=0 $Y2=0
cc_160 C1 N_A_43_57#_c_251_n 0.00875454f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_161 N_C1_M1004_g N_A_43_57#_c_283_n 0.0018373f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_162 C1 N_A_43_57#_c_283_n 0.0226385f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_163 N_C1_c_190_n N_A_43_57#_c_283_n 7.21459e-19 $X=2.235 $Y=1.335 $X2=0 $Y2=0
cc_164 N_C1_M1011_g N_A_43_57#_c_243_n 0.00435208f $X=2.195 $Y=2.545 $X2=0 $Y2=0
cc_165 N_C1_c_190_n N_A_43_57#_c_243_n 0.00622524f $X=2.235 $Y=1.335 $X2=0 $Y2=0
cc_166 N_C1_M1007_g N_A_43_57#_c_245_n 0.00275578f $X=2.185 $Y=0.495 $X2=0 $Y2=0
cc_167 N_C1_c_188_n N_A_43_57#_c_245_n 3.10581e-19 $X=2.545 $Y=1.245 $X2=0 $Y2=0
cc_168 C1 N_A_43_57#_c_245_n 0.0075854f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_169 N_C1_M1004_g N_A_43_57#_c_246_n 0.0266754f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_170 C1 N_A_43_57#_c_246_n 0.00123914f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_171 N_C1_c_190_n N_A_43_57#_c_246_n 0.00397189f $X=2.235 $Y=1.335 $X2=0 $Y2=0
cc_172 N_C1_M1011_g N_A_29_409#_c_331_n 7.25172e-19 $X=2.195 $Y=2.545 $X2=0
+ $Y2=0
cc_173 N_C1_M1011_g N_A_29_409#_c_333_n 0.00376238f $X=2.195 $Y=2.545 $X2=0
+ $Y2=0
cc_174 N_C1_M1011_g N_VPWR_c_362_n 0.00316346f $X=2.195 $Y=2.545 $X2=0 $Y2=0
cc_175 N_C1_M1011_g N_VPWR_c_363_n 0.0086001f $X=2.195 $Y=2.545 $X2=0 $Y2=0
cc_176 N_C1_M1011_g N_VPWR_c_360_n 0.0166934f $X=2.195 $Y=2.545 $X2=0 $Y2=0
cc_177 N_C1_M1007_g N_VGND_c_416_n 0.00188065f $X=2.185 $Y=0.495 $X2=0 $Y2=0
cc_178 N_C1_M1004_g N_VGND_c_416_n 0.0105659f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_179 N_C1_M1007_g N_VGND_c_418_n 0.00502664f $X=2.185 $Y=0.495 $X2=0 $Y2=0
cc_180 N_C1_M1004_g N_VGND_c_418_n 0.00445056f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_181 N_C1_M1007_g N_VGND_c_420_n 0.00562693f $X=2.185 $Y=0.495 $X2=0 $Y2=0
cc_182 N_C1_M1004_g N_VGND_c_420_n 0.00418511f $X=2.545 $Y=0.495 $X2=0 $Y2=0
cc_183 N_A_43_57#_c_250_n N_VPWR_M1006_s 0.00494755f $X=2.875 $Y=2.105 $X2=0
+ $Y2=0
cc_184 N_A_43_57#_M1006_g N_VPWR_c_362_n 0.0193891f $X=3.285 $Y=2.545 $X2=0
+ $Y2=0
cc_185 N_A_43_57#_c_249_n N_VPWR_c_362_n 0.0468558f $X=2.46 $Y=2.9 $X2=0 $Y2=0
cc_186 N_A_43_57#_c_250_n N_VPWR_c_362_n 0.0161868f $X=2.875 $Y=2.105 $X2=0
+ $Y2=0
cc_187 N_A_43_57#_c_249_n N_VPWR_c_363_n 0.0220321f $X=2.46 $Y=2.9 $X2=0 $Y2=0
cc_188 N_A_43_57#_M1006_g N_VPWR_c_365_n 0.00769046f $X=3.285 $Y=2.545 $X2=0
+ $Y2=0
cc_189 N_A_43_57#_M1006_g N_VPWR_c_360_n 0.0140911f $X=3.285 $Y=2.545 $X2=0
+ $Y2=0
cc_190 N_A_43_57#_c_249_n N_VPWR_c_360_n 0.0125808f $X=2.46 $Y=2.9 $X2=0 $Y2=0
cc_191 N_A_43_57#_c_236_n X 0.00191848f $X=2.975 $Y=0.82 $X2=0 $Y2=0
cc_192 N_A_43_57#_M1006_g X 0.0440508f $X=3.285 $Y=2.545 $X2=0 $Y2=0
cc_193 N_A_43_57#_c_238_n X 0.012579f $X=3.335 $Y=0.82 $X2=0 $Y2=0
cc_194 N_A_43_57#_c_250_n X 0.00828461f $X=2.875 $Y=2.105 $X2=0 $Y2=0
cc_195 N_A_43_57#_c_242_n X 0.0129587f $X=3.04 $Y=0.99 $X2=0 $Y2=0
cc_196 N_A_43_57#_c_283_n X 0.0357696f $X=3.04 $Y=1.325 $X2=0 $Y2=0
cc_197 N_A_43_57#_c_243_n X 0.0236558f $X=2.96 $Y=2.02 $X2=0 $Y2=0
cc_198 N_A_43_57#_c_246_n X 0.0247553f $X=3.04 $Y=0.985 $X2=0 $Y2=0
cc_199 N_A_43_57#_c_244_n A_130_57# 0.00206159f $X=0.36 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_43_57#_c_239_n N_VGND_c_415_n 0.0199879f $X=1.805 $Y=0.905 $X2=0
+ $Y2=0
cc_201 N_A_43_57#_c_240_n N_VGND_c_415_n 0.0125465f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_202 N_A_43_57#_c_244_n N_VGND_c_415_n 0.00920801f $X=0.36 $Y=0.495 $X2=0
+ $Y2=0
cc_203 N_A_43_57#_c_236_n N_VGND_c_416_n 0.0105649f $X=2.975 $Y=0.82 $X2=0 $Y2=0
cc_204 N_A_43_57#_c_238_n N_VGND_c_416_n 0.00188065f $X=3.335 $Y=0.82 $X2=0
+ $Y2=0
cc_205 N_A_43_57#_c_240_n N_VGND_c_416_n 0.0125465f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_206 N_A_43_57#_c_241_n N_VGND_c_416_n 0.0174453f $X=2.875 $Y=0.905 $X2=0
+ $Y2=0
cc_207 N_A_43_57#_c_242_n N_VGND_c_416_n 0.0027879f $X=3.04 $Y=0.99 $X2=0 $Y2=0
cc_208 N_A_43_57#_c_244_n N_VGND_c_417_n 0.0275623f $X=0.36 $Y=0.495 $X2=0 $Y2=0
cc_209 N_A_43_57#_c_240_n N_VGND_c_418_n 0.021949f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_210 N_A_43_57#_c_236_n N_VGND_c_419_n 0.00445056f $X=2.975 $Y=0.82 $X2=0
+ $Y2=0
cc_211 N_A_43_57#_c_238_n N_VGND_c_419_n 0.00502664f $X=3.335 $Y=0.82 $X2=0
+ $Y2=0
cc_212 N_A_43_57#_c_236_n N_VGND_c_420_n 0.00418302f $X=2.975 $Y=0.82 $X2=0
+ $Y2=0
cc_213 N_A_43_57#_c_238_n N_VGND_c_420_n 0.0100677f $X=3.335 $Y=0.82 $X2=0 $Y2=0
cc_214 N_A_43_57#_c_239_n N_VGND_c_420_n 0.0202154f $X=1.805 $Y=0.905 $X2=0
+ $Y2=0
cc_215 N_A_43_57#_c_240_n N_VGND_c_420_n 0.0124703f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_216 N_A_43_57#_c_241_n N_VGND_c_420_n 0.0153271f $X=2.875 $Y=0.905 $X2=0
+ $Y2=0
cc_217 N_A_43_57#_c_242_n N_VGND_c_420_n 0.00985419f $X=3.04 $Y=0.99 $X2=0 $Y2=0
cc_218 N_A_43_57#_c_244_n N_VGND_c_420_n 0.0215106f $X=0.36 $Y=0.495 $X2=0 $Y2=0
cc_219 N_A_29_409#_c_331_n N_VPWR_M1000_d 0.00235187f $X=1.235 $Y=2.105
+ $X2=-0.19 $Y2=1.655
cc_220 N_A_29_409#_c_330_n N_VPWR_c_361_n 0.045794f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_221 N_A_29_409#_c_331_n N_VPWR_c_361_n 0.0185435f $X=1.235 $Y=2.105 $X2=0
+ $Y2=0
cc_222 N_A_29_409#_c_333_n N_VPWR_c_361_n 0.0197666f $X=1.4 $Y=2.9 $X2=0 $Y2=0
cc_223 N_A_29_409#_c_333_n N_VPWR_c_363_n 0.021949f $X=1.4 $Y=2.9 $X2=0 $Y2=0
cc_224 N_A_29_409#_c_330_n N_VPWR_c_360_n 0.0125808f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_225 N_A_29_409#_c_333_n N_VPWR_c_360_n 0.0124703f $X=1.4 $Y=2.9 $X2=0 $Y2=0
cc_226 N_A_29_409#_c_330_n N_VPWR_c_367_n 0.0220321f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_227 N_VPWR_c_362_n X 0.045794f $X=3.02 $Y=2.535 $X2=0 $Y2=0
cc_228 N_VPWR_c_365_n X 0.0220321f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_c_360_n X 0.0125808f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_230 X N_VGND_c_416_n 0.0125465f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_231 X N_VGND_c_419_n 0.0220321f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_232 X N_VGND_c_420_n 0.0125808f $X=3.515 $Y=0.47 $X2=0 $Y2=0
