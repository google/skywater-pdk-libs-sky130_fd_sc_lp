* File: sky130_fd_sc_lp__nand4_m.pxi.spice
* Created: Fri Aug 28 10:51:21 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4_M%D N_D_M1004_g N_D_M1001_g N_D_c_61_n N_D_c_66_n D
+ D D D N_D_c_63_n PM_SKY130_FD_SC_LP__NAND4_M%D
x_PM_SKY130_FD_SC_LP__NAND4_M%C N_C_M1005_g N_C_M1006_g N_C_c_94_n N_C_c_95_n
+ N_C_c_96_n C C C C N_C_c_98_n PM_SKY130_FD_SC_LP__NAND4_M%C
x_PM_SKY130_FD_SC_LP__NAND4_M%B N_B_M1007_g N_B_M1003_g N_B_c_141_n N_B_c_142_n
+ N_B_c_143_n B B B B N_B_c_145_n PM_SKY130_FD_SC_LP__NAND4_M%B
x_PM_SKY130_FD_SC_LP__NAND4_M%A N_A_M1000_g N_A_M1002_g N_A_c_190_n N_A_c_197_n
+ N_A_c_191_n N_A_c_192_n A A A N_A_c_194_n PM_SKY130_FD_SC_LP__NAND4_M%A
x_PM_SKY130_FD_SC_LP__NAND4_M%VPWR N_VPWR_M1001_s N_VPWR_M1006_d N_VPWR_M1000_d
+ N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n
+ N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_240_n VPWR N_VPWR_c_241_n
+ N_VPWR_c_232_n PM_SKY130_FD_SC_LP__NAND4_M%VPWR
x_PM_SKY130_FD_SC_LP__NAND4_M%Y N_Y_M1002_d N_Y_M1001_d N_Y_M1003_d N_Y_c_266_n
+ N_Y_c_267_n N_Y_c_269_n Y Y Y N_Y_c_272_n Y N_Y_c_273_n N_Y_c_274_n
+ PM_SKY130_FD_SC_LP__NAND4_M%Y
x_PM_SKY130_FD_SC_LP__NAND4_M%VGND N_VGND_M1004_s N_VGND_c_318_n N_VGND_c_319_n
+ N_VGND_c_320_n VGND N_VGND_c_321_n N_VGND_c_322_n
+ PM_SKY130_FD_SC_LP__NAND4_M%VGND
cc_1 VNB N_D_M1004_g 0.0466619f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.445
cc_2 VNB N_D_c_61_n 0.0286295f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_3 VNB D 0.0445505f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_D_c_63_n 0.018587f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_5 VNB N_C_M1006_g 0.0116186f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.52
cc_6 VNB N_C_c_94_n 0.0167966f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_7 VNB N_C_c_95_n 0.0239175f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_8 VNB N_C_c_96_n 0.0172122f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.675
cc_9 VNB C 0.00281609f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_10 VNB N_C_c_98_n 0.0175199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_M1003_g 0.0101297f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.52
cc_12 VNB N_B_c_141_n 0.0176297f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_13 VNB N_B_c_142_n 0.0217661f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_14 VNB N_B_c_143_n 0.0161422f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.675
cc_15 VNB B 0.0105029f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_16 VNB N_B_c_145_n 0.0164565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_M1002_g 0.0251256f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.52
cc_18 VNB N_A_c_190_n 0.00886083f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_19 VNB N_A_c_191_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_20 VNB N_A_c_192_n 0.0173274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A 0.0103336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_194_n 0.0164912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_232_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_266_n 0.0476196f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.675
cc_25 VNB N_Y_c_267_n 0.0212576f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_VGND_c_318_n 0.01277f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.52
cc_27 VNB N_VGND_c_319_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_28 VNB N_VGND_c_320_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.155
cc_29 VNB N_VGND_c_321_n 0.0655869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_322_n 0.17471f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.32
cc_31 VPB N_D_M1001_g 0.0436616f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.52
cc_32 VPB N_D_c_61_n 0.00167004f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_33 VPB N_D_c_66_n 0.032692f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.825
cc_34 VPB D 0.0423187f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_35 VPB N_C_M1006_g 0.044515f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.52
cc_36 VPB C 0.00176994f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_37 VPB N_B_M1003_g 0.0439676f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.52
cc_38 VPB B 0.00244611f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_39 VPB N_A_M1000_g 0.0400602f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.445
cc_40 VPB N_A_c_190_n 0.00116914f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.155
cc_41 VPB N_A_c_197_n 0.0163044f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.825
cc_42 VPB A 0.00202503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_233_n 0.0259256f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_44 VPB N_VPWR_c_234_n 0.0195397f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_45 VPB N_VPWR_c_235_n 0.0140295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_236_n 0.0291792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_237_n 0.0193272f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.32
cc_48 VPB N_VPWR_c_238_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.32
cc_49 VPB N_VPWR_c_239_n 0.0190583f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_240_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_241_n 0.0227638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_232_n 0.0975285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_Y_c_266_n 0.0147507f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.675
cc_54 VPB N_Y_c_269_n 0.028574f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_55 VPB Y 0.00594531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB Y 0.00726222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_272_n 0.0155963f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.295
cc_58 VPB N_Y_c_273_n 0.0110459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_Y_c_274_n 0.0167707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_D_c_61_n N_C_M1006_g 0.00599184f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_61 N_D_c_66_n N_C_M1006_g 0.0319303f $X=0.7 $Y=1.825 $X2=0 $Y2=0
cc_62 D N_C_M1006_g 6.05906e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_63 N_D_M1004_g N_C_c_94_n 0.0236544f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_64 N_D_c_61_n N_C_c_95_n 0.0236544f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_65 N_D_M1004_g C 0.00387617f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_66 N_D_c_61_n C 0.00188577f $X=0.7 $Y=1.675 $X2=0 $Y2=0
cc_67 N_D_c_66_n C 6.64602e-19 $X=0.7 $Y=1.825 $X2=0 $Y2=0
cc_68 D C 0.0351531f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_69 D N_C_c_98_n 0.00200864f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_D_c_63_n N_C_c_98_n 0.0236544f $X=0.63 $Y=1.32 $X2=0 $Y2=0
cc_71 N_D_M1001_g N_VPWR_c_233_n 0.00385941f $X=0.86 $Y=2.52 $X2=0 $Y2=0
cc_72 N_D_c_66_n N_VPWR_c_233_n 0.00194827f $X=0.7 $Y=1.825 $X2=0 $Y2=0
cc_73 D N_VPWR_c_233_n 0.0155616f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_74 N_D_M1001_g N_VPWR_c_239_n 0.00428744f $X=0.86 $Y=2.52 $X2=0 $Y2=0
cc_75 N_D_M1001_g N_VPWR_c_232_n 0.00476395f $X=0.86 $Y=2.52 $X2=0 $Y2=0
cc_76 N_D_M1001_g Y 0.0017351f $X=0.86 $Y=2.52 $X2=0 $Y2=0
cc_77 D Y 0.011747f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_78 N_D_M1001_g N_Y_c_273_n 0.00584267f $X=0.86 $Y=2.52 $X2=0 $Y2=0
cc_79 N_D_M1004_g N_VGND_c_318_n 0.0107712f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_80 D N_VGND_c_318_n 0.013835f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_81 N_D_c_63_n N_VGND_c_318_n 5.94371e-19 $X=0.63 $Y=1.32 $X2=0 $Y2=0
cc_82 N_D_M1004_g N_VGND_c_321_n 0.00486043f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_83 N_D_M1004_g N_VGND_c_322_n 0.00693889f $X=0.72 $Y=0.445 $X2=0 $Y2=0
cc_84 D N_VGND_c_322_n 0.0104926f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_85 N_C_M1006_g N_B_M1003_g 0.0441254f $X=1.29 $Y=2.52 $X2=0 $Y2=0
cc_86 C N_B_M1003_g 3.38916e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_87 N_C_c_94_n N_B_c_141_n 0.0198776f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_88 C N_B_c_141_n 0.0010831f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_89 N_C_c_95_n N_B_c_142_n 0.0118633f $X=1.2 $Y=1.27 $X2=0 $Y2=0
cc_90 N_C_c_96_n N_B_c_143_n 0.0118633f $X=1.2 $Y=1.435 $X2=0 $Y2=0
cc_91 N_C_c_94_n B 4.80776e-19 $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_92 C B 0.0565648f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_93 N_C_c_98_n B 0.00665631f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_94 C N_B_c_145_n 7.52967e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_95 N_C_c_98_n N_B_c_145_n 0.0118633f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_96 N_C_M1006_g N_VPWR_c_234_n 0.00127635f $X=1.29 $Y=2.52 $X2=0 $Y2=0
cc_97 N_C_M1006_g N_VPWR_c_239_n 0.00428744f $X=1.29 $Y=2.52 $X2=0 $Y2=0
cc_98 N_C_M1006_g N_VPWR_c_232_n 0.00476395f $X=1.29 $Y=2.52 $X2=0 $Y2=0
cc_99 N_C_c_96_n Y 0.00299025f $X=1.2 $Y=1.435 $X2=0 $Y2=0
cc_100 C Y 0.00534285f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_101 N_C_M1006_g N_Y_c_272_n 0.017164f $X=1.29 $Y=2.52 $X2=0 $Y2=0
cc_102 C N_Y_c_272_n 0.00721346f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_103 N_C_M1006_g N_Y_c_273_n 0.00375072f $X=1.29 $Y=2.52 $X2=0 $Y2=0
cc_104 N_C_c_94_n N_VGND_c_318_n 0.00229416f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_105 C N_VGND_c_318_n 4.91318e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_106 N_C_c_94_n N_VGND_c_321_n 0.00499463f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_107 C N_VGND_c_321_n 0.00398853f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_C_c_98_n N_VGND_c_321_n 0.00187414f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_109 N_C_c_94_n N_VGND_c_322_n 0.00880207f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_110 C N_VGND_c_322_n 0.00539257f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_111 N_C_c_98_n N_VGND_c_322_n 0.00216458f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_112 C A_237_47# 0.00271716f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_113 N_B_c_141_n N_A_M1002_g 0.0186799f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_114 B N_A_M1002_g 0.00412971f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_115 N_B_c_145_n N_A_M1002_g 0.0117064f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_116 N_B_M1003_g N_A_c_197_n 0.0351133f $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_117 B N_A_c_197_n 4.63942e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_118 N_B_c_143_n N_A_c_191_n 0.0117064f $X=1.77 $Y=1.435 $X2=0 $Y2=0
cc_119 N_B_M1003_g N_A_c_192_n 0.00712579f $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_120 B N_A_c_192_n 7.31847e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_121 N_B_M1003_g A 9.30151e-19 $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_122 B A 0.0595903f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_123 N_B_c_145_n A 0.00426123f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_124 N_B_c_142_n N_A_c_194_n 0.0117064f $X=1.77 $Y=1.27 $X2=0 $Y2=0
cc_125 B N_A_c_194_n 5.64969e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_126 N_B_M1003_g N_VPWR_c_234_n 0.00127635f $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_127 N_B_M1003_g N_VPWR_c_241_n 0.00428744f $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_128 N_B_M1003_g N_VPWR_c_232_n 0.00476395f $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_129 B N_Y_c_267_n 0.00323191f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_130 N_B_c_143_n Y 0.00280598f $X=1.77 $Y=1.435 $X2=0 $Y2=0
cc_131 B Y 0.00200357f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 N_B_M1003_g N_Y_c_272_n 0.0151564f $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_133 N_B_c_143_n N_Y_c_272_n 2.63136e-19 $X=1.77 $Y=1.435 $X2=0 $Y2=0
cc_134 B N_Y_c_272_n 0.0163169f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_135 N_B_M1003_g N_Y_c_274_n 0.0041259f $X=1.72 $Y=2.52 $X2=0 $Y2=0
cc_136 N_B_c_141_n N_VGND_c_321_n 0.00398598f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_137 B N_VGND_c_321_n 0.00634804f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_138 N_B_c_145_n N_VGND_c_321_n 0.00185537f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_139 N_B_c_141_n N_VGND_c_322_n 0.00636002f $X=1.77 $Y=0.765 $X2=0 $Y2=0
cc_140 B N_VGND_c_322_n 0.00806027f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_141 N_B_c_145_n N_VGND_c_322_n 0.00213938f $X=1.77 $Y=0.93 $X2=0 $Y2=0
cc_142 B A_351_47# 0.00330582f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_143 N_A_M1000_g N_VPWR_c_236_n 0.00380493f $X=2.15 $Y=2.52 $X2=0 $Y2=0
cc_144 N_A_M1000_g N_VPWR_c_241_n 6.53249e-19 $X=2.15 $Y=2.52 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_Y_c_266_n 0.00339766f $X=2.15 $Y=2.52 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_Y_c_266_n 0.00546311f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_c_190_n N_Y_c_266_n 0.00130879f $X=2.25 $Y=1.675 $X2=0 $Y2=0
cc_148 N_A_c_197_n N_Y_c_266_n 0.00242178f $X=2.25 $Y=1.75 $X2=0 $Y2=0
cc_149 A N_Y_c_266_n 0.0667326f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_150 N_A_c_194_n N_Y_c_266_n 0.0163648f $X=2.34 $Y=1.005 $X2=0 $Y2=0
cc_151 A N_Y_c_267_n 0.00343308f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_152 N_A_c_194_n N_Y_c_267_n 0.00384253f $X=2.34 $Y=1.005 $X2=0 $Y2=0
cc_153 N_A_c_197_n N_Y_c_269_n 0.00224923f $X=2.25 $Y=1.75 $X2=0 $Y2=0
cc_154 N_A_c_192_n N_Y_c_269_n 0.00290373f $X=2.34 $Y=1.51 $X2=0 $Y2=0
cc_155 A N_Y_c_269_n 0.0130725f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_156 N_A_M1000_g Y 0.0106283f $X=2.15 $Y=2.52 $X2=0 $Y2=0
cc_157 N_A_c_197_n Y 5.85208e-19 $X=2.25 $Y=1.75 $X2=0 $Y2=0
cc_158 A Y 0.0126344f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_159 N_A_M1000_g N_Y_c_274_n 0.0266459f $X=2.15 $Y=2.52 $X2=0 $Y2=0
cc_160 N_A_M1002_g N_VGND_c_321_n 0.00585385f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_M1002_g N_VGND_c_322_n 0.00801226f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_162 A N_VGND_c_322_n 0.010685f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_163 N_VPWR_c_236_n N_Y_c_269_n 0.0170452f $X=2.53 $Y=2.525 $X2=0 $Y2=0
cc_164 N_VPWR_c_234_n N_Y_c_272_n 0.0168699f $X=1.505 $Y=2.525 $X2=0 $Y2=0
cc_165 N_VPWR_c_233_n N_Y_c_273_n 0.0154405f $X=0.645 $Y=2.525 $X2=0 $Y2=0
cc_166 N_VPWR_c_234_n N_Y_c_273_n 0.0154405f $X=1.505 $Y=2.525 $X2=0 $Y2=0
cc_167 N_VPWR_c_239_n N_Y_c_273_n 0.00859063f $X=1.4 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_232_n N_Y_c_273_n 0.0075889f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_169 N_VPWR_c_234_n N_Y_c_274_n 0.0162792f $X=1.505 $Y=2.525 $X2=0 $Y2=0
cc_170 N_VPWR_c_236_n N_Y_c_274_n 0.0339021f $X=2.53 $Y=2.525 $X2=0 $Y2=0
cc_171 N_VPWR_c_241_n N_Y_c_274_n 0.0170574f $X=2.425 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_232_n N_Y_c_274_n 0.0150683f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_173 N_Y_c_267_n N_VGND_c_321_n 0.0178198f $X=2.69 $Y=0.495 $X2=0 $Y2=0
cc_174 N_Y_M1002_d N_VGND_c_322_n 0.0027096f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_175 N_Y_c_267_n N_VGND_c_322_n 0.0144125f $X=2.69 $Y=0.495 $X2=0 $Y2=0
cc_176 N_VGND_c_322_n A_159_47# 0.010279f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_177 N_VGND_c_322_n A_237_47# 0.0125365f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_178 N_VGND_c_322_n A_351_47# 0.0100481f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
