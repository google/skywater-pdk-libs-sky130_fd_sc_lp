* NGSPICE file created from sky130_fd_sc_lp__a2bb2oi_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2bb2oi_m A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A2_N a_202_47# VNB nshort w=420000u l=150000u
+  ad=3.633e+11p pd=4.25e+06u as=1.176e+11p ps=1.4e+06u
M1001 Y a_202_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1002 a_202_47# A2_N a_132_517# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1003 VPWR B2 a_403_387# VPB phighvt w=420000u l=150000u
+  ad=2.625e+11p pd=2.93e+06u as=2.289e+11p ps=2.77e+06u
M1004 VGND B1 a_467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1005 a_202_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_403_387# a_202_47# Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 a_132_517# A1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_467_47# B2 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_403_387# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

