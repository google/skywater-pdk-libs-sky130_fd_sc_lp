* File: sky130_fd_sc_lp__dfstp_2.spice
* Created: Fri Aug 28 10:23:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfstp_2.pex.spice"
.subckt sky130_fd_sc_lp__dfstp_2  VNB VPB CLK D SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_CLK_M1007_g N_A_27_465#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1197 PD=0.74 PS=1.41 NRD=5.712 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_196_465#_M1015_d N_A_27_465#_M1015_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_400_119#_M1006_d N_D_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1029 N_A_486_119#_M1029_d N_A_27_465#_M1029_g N_A_400_119#_M1006_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1031 A_572_119# N_A_196_465#_M1031_g N_A_486_119#_M1029_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_614_93#_M1021_g A_572_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 A_857_47# N_A_486_119#_M1020_g N_A_614_93#_M1020_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_SET_B_M1010_g A_857_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.135747 AS=0.0441 PD=1.01038 PS=0.63 NRD=79.284 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1027 A_1086_47# N_A_486_119#_M1027_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.206853 PD=0.85 PS=1.53962 NRD=9.372 NRS=14.988 M=1 R=4.26667
+ SA=75001 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1030 N_A_1158_47#_M1030_d N_A_196_465#_M1030_g A_1086_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.138023 AS=0.0672 PD=1.24981 PS=0.85 NRD=3.744 NRS=9.372 M=1
+ R=4.26667 SA=75001.3 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1032 A_1267_91# N_A_27_465#_M1032_g N_A_1158_47#_M1030_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0905774 PD=0.63 PS=0.820189 NRD=14.28 NRS=27.852 M=1
+ R=2.8 SA=75001.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 A_1339_91# N_A_1309_65#_M1001_g A_1267_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_SET_B_M1013_g A_1339_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.08925 AS=0.0441 PD=0.845 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1017 N_A_1309_65#_M1017_d N_A_1158_47#_M1017_g N_VGND_M1013_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.08925 PD=1.41 PS=0.845 NRD=5.712 NRS=41.424 M=1
+ R=2.8 SA=75003 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_1158_47#_M1018_g N_A_1855_47#_M1018_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0903 AS=0.1113 PD=0.8 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 N_Q_M1016_d N_A_1855_47#_M1016_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1806 PD=1.12 PS=1.6 NRD=0 NRS=4.284 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1028 N_Q_M1016_d N_A_1855_47#_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_CLK_M1009_g N_A_27_465#_M1009_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1024 N_A_196_465#_M1024_d N_A_27_465#_M1024_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.176 AS=0.0896 PD=1.83 PS=0.92 NRD=3.0732 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_A_400_119#_M1011_d N_D_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.1
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_486_119#_M1002_d N_A_196_465#_M1002_g N_A_400_119#_M1011_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1019 A_572_463# N_A_27_465#_M1019_g N_A_486_119#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_614_93#_M1023_g A_572_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=4.6886 NRS=23.443 M=1 R=2.8 SA=75001.4
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_614_93#_M1003_d N_A_486_119#_M1003_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=46.886 M=1 R=2.8
+ SA=75001.9 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_SET_B_M1025_g N_A_614_93#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1211 AS=0.0588 PD=0.96 PS=0.7 NRD=76.2193 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1000 N_A_988_379#_M1000_d N_A_486_119#_M1000_g N_VPWR_M1025_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2422 PD=2.21 PS=1.92 NRD=0 NRS=37.5088 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1014 N_A_1158_47#_M1014_d N_A_196_465#_M1014_g N_A_1095_425#_M1014_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0952 AS=0.1113 PD=0.823333 PS=1.37 NRD=28.1316
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1026 N_A_988_379#_M1026_d N_A_27_465#_M1026_g N_A_1158_47#_M1014_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.30685 AS=0.1904 PD=2.66 PS=1.64667 NRD=23.443 NRS=12.8838
+ M=1 R=5.6 SA=75000.5 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_1309_65#_M1008_g N_A_1095_425#_M1008_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_1158_47#_M1033_d N_SET_B_M1033_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_1309_65#_M1004_d N_A_1158_47#_M1004_g N_VPWR_M1004_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_1158_47#_M1005_g N_A_1855_47#_M1005_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.129819 AS=0.1696 PD=1.09137 PS=1.81 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 N_Q_M1012_d N_A_1855_47#_M1012_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.255581 PD=1.54 PS=2.14863 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75000.4 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1022 N_Q_M1012_d N_A_1855_47#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=21.5167 P=26.99
c_126 VNB 0 1.77925e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfstp_2.pxi.spice"
*
.ends
*
*
