* File: sky130_fd_sc_lp__sdfrbp_lp.pxi.spice
* Created: Fri Aug 28 11:28:03 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%SCE N_SCE_M1040_g N_SCE_M1024_g N_SCE_M1017_g
+ N_SCE_M1016_g N_SCE_c_382_n N_SCE_c_383_n N_SCE_M1008_g N_SCE_M1013_g
+ N_SCE_c_385_n N_SCE_c_386_n N_SCE_c_387_n SCE SCE SCE N_SCE_c_389_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%SCE
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%D N_D_M1014_g N_D_M1059_g N_D_c_453_n
+ N_D_c_454_n N_D_c_455_n N_D_c_456_n D N_D_c_457_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%D
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_29_47# N_A_29_47#_M1040_s N_A_29_47#_M1024_s
+ N_A_29_47#_M1004_g N_A_29_47#_M1056_g N_A_29_47#_c_502_n N_A_29_47#_c_503_n
+ N_A_29_47#_c_510_n N_A_29_47#_c_504_n N_A_29_47#_c_505_n N_A_29_47#_c_506_n
+ N_A_29_47#_c_507_n N_A_29_47#_c_508_n PM_SKY130_FD_SC_LP__SDFRBP_LP%A_29_47#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%SCD N_SCD_M1023_g N_SCD_c_572_n N_SCD_M1050_g
+ N_SCD_c_573_n N_SCD_c_574_n SCD N_SCD_c_576_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%SCD
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_876_93# N_A_876_93#_M1010_d
+ N_A_876_93#_M1029_d N_A_876_93#_M1032_g N_A_876_93#_M1006_g
+ N_A_876_93#_M1044_g N_A_876_93#_M1051_g N_A_876_93#_c_613_n
+ N_A_876_93#_c_614_n N_A_876_93#_c_615_n N_A_876_93#_c_665_p
+ N_A_876_93#_c_616_n N_A_876_93#_c_617_n N_A_876_93#_c_618_n
+ N_A_876_93#_c_636_p N_A_876_93#_c_637_p N_A_876_93#_c_669_p
+ N_A_876_93#_c_619_n N_A_876_93#_c_620_n N_A_876_93#_c_629_n
+ N_A_876_93#_c_621_n N_A_876_93#_c_622_n N_A_876_93#_c_623_n
+ N_A_876_93#_c_624_n N_A_876_93#_c_625_n N_A_876_93#_c_626_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%A_876_93#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_967_193# N_A_967_193#_M1026_s
+ N_A_967_193#_M1052_s N_A_967_193#_M1015_g N_A_967_193#_M1028_g
+ N_A_967_193#_c_791_n N_A_967_193#_c_792_n N_A_967_193#_M1025_g
+ N_A_967_193#_M1057_g N_A_967_193#_M1029_g N_A_967_193#_M1010_g
+ N_A_967_193#_c_795_n N_A_967_193#_c_796_n N_A_967_193#_c_797_n
+ N_A_967_193#_c_798_n N_A_967_193#_c_799_n N_A_967_193#_c_800_n
+ N_A_967_193#_c_825_n N_A_967_193#_c_826_n N_A_967_193#_M1042_g
+ N_A_967_193#_M1045_g N_A_967_193#_c_802_n N_A_967_193#_c_803_n
+ N_A_967_193#_c_804_n N_A_967_193#_c_805_n N_A_967_193#_c_806_n
+ N_A_967_193#_c_807_n N_A_967_193#_c_828_n N_A_967_193#_c_829_n
+ N_A_967_193#_c_830_n N_A_967_193#_c_831_n N_A_967_193#_c_832_n
+ N_A_967_193#_c_808_n N_A_967_193#_c_809_n N_A_967_193#_c_810_n
+ N_A_967_193#_c_835_n N_A_967_193#_c_836_n N_A_967_193#_c_811_n
+ N_A_967_193#_c_812_n N_A_967_193#_c_813_n N_A_967_193#_c_814_n
+ N_A_967_193#_c_815_n N_A_967_193#_c_816_n N_A_967_193#_c_817_n
+ N_A_967_193#_c_818_n PM_SKY130_FD_SC_LP__SDFRBP_LP%A_967_193#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_1147_490# N_A_1147_490#_M1000_s
+ N_A_1147_490#_M1051_s N_A_1147_490#_M1002_s N_A_1147_490#_M1042_d
+ N_A_1147_490#_c_1103_n N_A_1147_490#_M1003_g N_A_1147_490#_c_1104_n
+ N_A_1147_490#_c_1105_n N_A_1147_490#_M1030_g N_A_1147_490#_c_1091_n
+ N_A_1147_490#_c_1092_n N_A_1147_490#_c_1093_n N_A_1147_490#_c_1094_n
+ N_A_1147_490#_c_1095_n N_A_1147_490#_c_1109_n N_A_1147_490#_c_1184_n
+ N_A_1147_490#_c_1110_n N_A_1147_490#_c_1111_n N_A_1147_490#_c_1112_n
+ N_A_1147_490#_c_1096_n N_A_1147_490#_c_1097_n N_A_1147_490#_c_1098_n
+ N_A_1147_490#_c_1099_n N_A_1147_490#_c_1100_n N_A_1147_490#_c_1101_n
+ N_A_1147_490#_c_1114_n N_A_1147_490#_c_1102_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%A_1147_490#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%RESET_B N_RESET_B_c_1299_n N_RESET_B_M1047_g
+ N_RESET_B_c_1285_n N_RESET_B_c_1286_n N_RESET_B_M1041_g N_RESET_B_c_1288_n
+ N_RESET_B_c_1289_n N_RESET_B_c_1302_n N_RESET_B_M1048_g N_RESET_B_M1043_g
+ N_RESET_B_M1005_g N_RESET_B_M1049_g N_RESET_B_M1054_g N_RESET_B_c_1306_n
+ N_RESET_B_M1038_g N_RESET_B_M1036_g N_RESET_B_c_1292_n N_RESET_B_c_1293_n
+ N_RESET_B_c_1294_n N_RESET_B_c_1295_n N_RESET_B_c_1296_n N_RESET_B_c_1311_n
+ N_RESET_B_c_1312_n N_RESET_B_c_1313_n N_RESET_B_c_1314_n N_RESET_B_c_1315_n
+ N_RESET_B_c_1316_n RESET_B N_RESET_B_c_1297_n N_RESET_B_c_1298_n
+ N_RESET_B_c_1318_n N_RESET_B_c_1319_n N_RESET_B_c_1320_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_911_219# N_A_911_219#_M1032_d
+ N_A_911_219#_M1006_d N_A_911_219#_M1049_d N_A_911_219#_c_1543_n
+ N_A_911_219#_M1000_g N_A_911_219#_M1002_g N_A_911_219#_c_1546_n
+ N_A_911_219#_M1021_g N_A_911_219#_M1009_g N_A_911_219#_c_1549_n
+ N_A_911_219#_c_1550_n N_A_911_219#_c_1560_n N_A_911_219#_c_1551_n
+ N_A_911_219#_c_1561_n N_A_911_219#_c_1562_n N_A_911_219#_c_1552_n
+ N_A_911_219#_c_1553_n N_A_911_219#_c_1554_n N_A_911_219#_c_1565_n
+ N_A_911_219#_c_1566_n N_A_911_219#_c_1619_n N_A_911_219#_c_1653_n
+ N_A_911_219#_c_1555_n N_A_911_219#_c_1556_n N_A_911_219#_c_1567_n
+ N_A_911_219#_c_1622_n N_A_911_219#_c_1568_n N_A_911_219#_c_1557_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%A_911_219#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2388_115# N_A_2388_115#_M1035_d
+ N_A_2388_115#_M1037_d N_A_2388_115#_c_1729_n N_A_2388_115#_M1011_g
+ N_A_2388_115#_M1018_g N_A_2388_115#_c_1730_n N_A_2388_115#_c_1738_n
+ N_A_2388_115#_c_1731_n N_A_2388_115#_c_1732_n N_A_2388_115#_c_1746_n
+ N_A_2388_115#_c_1739_n N_A_2388_115#_c_1740_n N_A_2388_115#_c_1741_n
+ N_A_2388_115#_c_1733_n N_A_2388_115#_c_1734_n N_A_2388_115#_c_1735_n
+ N_A_2388_115#_c_1736_n PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2388_115#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2168_439# N_A_2168_439#_M1051_d
+ N_A_2168_439#_M1044_d N_A_2168_439#_M1037_g N_A_2168_439#_c_1839_n
+ N_A_2168_439#_M1035_g N_A_2168_439#_c_1840_n N_A_2168_439#_c_1841_n
+ N_A_2168_439#_M1019_g N_A_2168_439#_M1046_g N_A_2168_439#_M1033_g
+ N_A_2168_439#_M1031_g N_A_2168_439#_M1007_g N_A_2168_439#_c_1847_n
+ N_A_2168_439#_M1022_g N_A_2168_439#_M1034_g N_A_2168_439#_c_1850_n
+ N_A_2168_439#_M1001_g N_A_2168_439#_M1039_g N_A_2168_439#_c_1853_n
+ N_A_2168_439#_c_1854_n N_A_2168_439#_c_1855_n N_A_2168_439#_c_1874_n
+ N_A_2168_439#_c_1856_n N_A_2168_439#_c_1876_n N_A_2168_439#_c_1877_n
+ N_A_2168_439#_c_1938_n N_A_2168_439#_c_1857_n N_A_2168_439#_c_1858_n
+ N_A_2168_439#_c_1859_n N_A_2168_439#_c_1860_n N_A_2168_439#_c_1861_n
+ N_A_2168_439#_c_1879_n N_A_2168_439#_c_1880_n N_A_2168_439#_c_1862_n
+ N_A_2168_439#_c_1863_n N_A_2168_439#_c_1864_n N_A_2168_439#_c_1865_n
+ N_A_2168_439#_c_1866_n N_A_2168_439#_c_1867_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2168_439#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%CLK N_CLK_M1026_g N_CLK_M1052_g N_CLK_M1027_g
+ N_CLK_M1055_g CLK N_CLK_c_2085_n N_CLK_c_2086_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%CLK
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_3416_137# N_A_3416_137#_M1022_s
+ N_A_3416_137#_M1034_s N_A_3416_137#_M1012_g N_A_3416_137#_M1053_g
+ N_A_3416_137#_M1020_g N_A_3416_137#_M1058_g N_A_3416_137#_c_2133_n
+ N_A_3416_137#_c_2134_n N_A_3416_137#_c_2135_n N_A_3416_137#_c_2136_n
+ N_A_3416_137#_c_2137_n PM_SKY130_FD_SC_LP__SDFRBP_LP%A_3416_137#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%VPWR N_VPWR_M1016_d N_VPWR_M1023_d
+ N_VPWR_M1003_d N_VPWR_M1009_d N_VPWR_M1018_d N_VPWR_M1036_d N_VPWR_M1055_d
+ N_VPWR_M1039_d N_VPWR_c_2192_n N_VPWR_c_2193_n N_VPWR_c_2194_n N_VPWR_c_2195_n
+ N_VPWR_c_2196_n N_VPWR_c_2197_n N_VPWR_c_2198_n N_VPWR_c_2199_n
+ N_VPWR_c_2200_n N_VPWR_c_2201_n N_VPWR_c_2202_n N_VPWR_c_2203_n VPWR
+ N_VPWR_c_2204_n N_VPWR_c_2205_n N_VPWR_c_2206_n N_VPWR_c_2207_n
+ N_VPWR_c_2208_n N_VPWR_c_2209_n N_VPWR_c_2210_n N_VPWR_c_2191_n
+ N_VPWR_c_2212_n N_VPWR_c_2213_n N_VPWR_c_2214_n N_VPWR_c_2215_n
+ N_VPWR_c_2216_n N_VPWR_c_2217_n PM_SKY130_FD_SC_LP__SDFRBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_342_261# N_A_342_261#_M1008_d
+ N_A_342_261#_M1015_d N_A_342_261#_M1014_d N_A_342_261#_M1048_d
+ N_A_342_261#_c_2407_n N_A_342_261#_c_2408_n N_A_342_261#_c_2409_n
+ N_A_342_261#_c_2410_n N_A_342_261#_c_2411_n N_A_342_261#_c_2439_n
+ N_A_342_261#_c_2440_n N_A_342_261#_c_2412_n N_A_342_261#_c_2421_n
+ N_A_342_261#_c_2422_n N_A_342_261#_c_2489_n N_A_342_261#_c_2413_n
+ N_A_342_261#_c_2414_n N_A_342_261#_c_2415_n N_A_342_261#_c_2416_n
+ N_A_342_261#_c_2417_n PM_SKY130_FD_SC_LP__SDFRBP_LP%A_342_261#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2081_439# N_A_2081_439#_M1044_s
+ N_A_2081_439#_M1018_s N_A_2081_439#_c_2552_n N_A_2081_439#_c_2553_n
+ N_A_2081_439#_c_2554_n N_A_2081_439#_c_2555_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2081_439#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2523_397# N_A_2523_397#_M1037_s
+ N_A_2523_397#_M1019_d N_A_2523_397#_c_2582_n N_A_2523_397#_c_2583_n
+ N_A_2523_397#_c_2584_n N_A_2523_397#_c_2585_n N_A_2523_397#_c_2586_n
+ N_A_2523_397#_c_2587_n PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2523_397#
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%Q_N N_Q_N_M1031_d N_Q_N_M1007_d N_Q_N_c_2634_n
+ N_Q_N_c_2635_n N_Q_N_c_2631_n Q_N Q_N N_Q_N_c_2632_n Q_N
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%Q N_Q_M1020_d N_Q_M1058_d Q Q Q Q Q Q Q
+ N_Q_c_2665_n PM_SKY130_FD_SC_LP__SDFRBP_LP%Q
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%VGND N_VGND_M1017_d N_VGND_M1041_s
+ N_VGND_M1005_d N_VGND_M1021_d N_VGND_M1011_d N_VGND_M1027_d N_VGND_M1001_d
+ N_VGND_c_2681_n N_VGND_c_2682_n N_VGND_c_2683_n N_VGND_c_2684_n
+ N_VGND_c_2685_n N_VGND_c_2686_n N_VGND_c_2687_n N_VGND_c_2688_n
+ N_VGND_c_2689_n N_VGND_c_2690_n N_VGND_c_2691_n VGND N_VGND_c_2692_n
+ N_VGND_c_2693_n N_VGND_c_2694_n N_VGND_c_2695_n N_VGND_c_2696_n
+ N_VGND_c_2697_n N_VGND_c_2698_n N_VGND_c_2699_n N_VGND_c_2700_n
+ N_VGND_c_2701_n N_VGND_c_2702_n N_VGND_c_2703_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%VGND
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%noxref_37 N_noxref_37_M1008_s
+ N_noxref_37_M1050_d N_noxref_37_c_2854_n N_noxref_37_c_2855_n
+ N_noxref_37_c_2856_n N_noxref_37_c_2857_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%noxref_37
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%noxref_39 N_noxref_39_M1004_d
+ N_noxref_39_M1041_d N_noxref_39_c_2888_n N_noxref_39_c_2889_n
+ N_noxref_39_c_2890_n N_noxref_39_c_2891_n N_noxref_39_c_2892_n
+ N_noxref_39_c_2893_n N_noxref_39_c_2894_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%noxref_39
x_PM_SKY130_FD_SC_LP__SDFRBP_LP%A_824_219# N_A_824_219#_M1032_s
+ N_A_824_219#_M1030_s N_A_824_219#_c_2941_n N_A_824_219#_c_2942_n
+ N_A_824_219#_c_2943_n N_A_824_219#_c_2944_n
+ PM_SKY130_FD_SC_LP__SDFRBP_LP%A_824_219#
cc_1 VNB N_SCE_M1040_g 0.0498534f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_2 VNB N_SCE_M1017_g 0.0545371f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.445
cc_3 VNB N_SCE_M1016_g 0.00851722f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.775
cc_4 VNB N_SCE_c_382_n 0.0303301f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.91
cc_5 VNB N_SCE_c_383_n 0.0175494f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.835
cc_6 VNB N_SCE_M1013_g 0.0160332f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_7 VNB N_SCE_c_385_n 0.0205046f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.465
cc_8 VNB N_SCE_c_386_n 7.95968e-19 $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.91
cc_9 VNB N_SCE_c_387_n 0.00426715f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.91
cc_10 VNB SCE 0.00340318f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_SCE_c_389_n 0.0251125f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.48
cc_12 VNB N_D_M1014_g 0.0137007f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_13 VNB N_D_M1059_g 0.0537436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_c_453_n 0.00873809f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.445
cc_15 VNB N_D_c_454_n 0.0207365f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.445
cc_16 VNB N_D_c_455_n 0.0522851f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.775
cc_17 VNB N_D_c_456_n 0.00399582f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.91
cc_18 VNB N_D_c_457_n 0.018492f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.985
cc_19 VNB N_A_29_47#_M1004_g 0.0295451f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.445
cc_20 VNB N_A_29_47#_M1056_g 0.0137007f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.985
cc_21 VNB N_A_29_47#_c_502_n 0.00803274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_29_47#_c_503_n 0.017419f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.835
cc_23 VNB N_A_29_47#_c_504_n 0.0131464f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.465
cc_24 VNB N_A_29_47#_c_505_n 0.0364011f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.835
cc_25 VNB N_A_29_47#_c_506_n 0.0127427f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.835
cc_26 VNB N_A_29_47#_c_507_n 0.0378855f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.985
cc_27 VNB N_A_29_47#_c_508_n 0.0376446f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.91
cc_28 VNB N_SCD_M1023_g 0.0196399f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_29 VNB N_SCD_c_572_n 0.018955f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.985
cc_30 VNB N_SCD_c_573_n 0.0219085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_SCD_c_574_n 0.004972f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.445
cc_32 VNB SCD 0.00845378f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.445
cc_33 VNB N_SCD_c_576_n 0.0366643f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.775
cc_34 VNB N_A_876_93#_M1032_g 0.056594f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.315
cc_35 VNB N_A_876_93#_M1051_g 0.0245852f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.835
cc_36 VNB N_A_876_93#_c_613_n 0.0443997f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.515
cc_37 VNB N_A_876_93#_c_614_n 0.0039802f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_38 VNB N_A_876_93#_c_615_n 0.00930618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_876_93#_c_616_n 0.00805422f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.465
cc_40 VNB N_A_876_93#_c_617_n 0.0164389f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.835
cc_41 VNB N_A_876_93#_c_618_n 0.00382049f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.91
cc_42 VNB N_A_876_93#_c_619_n 0.00410127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_876_93#_c_620_n 0.00536567f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.48
cc_44 VNB N_A_876_93#_c_621_n 0.00980626f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_45 VNB N_A_876_93#_c_622_n 0.00480951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_876_93#_c_623_n 0.0443045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_876_93#_c_624_n 0.00165251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_876_93#_c_625_n 9.63216e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_876_93#_c_626_n 0.0412445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_967_193#_M1015_g 0.0423798f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.315
cc_51 VNB N_A_967_193#_M1028_g 0.00222123f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.985
cc_52 VNB N_A_967_193#_c_791_n 0.0461708f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.775
cc_53 VNB N_A_967_193#_c_792_n 0.0142736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_967_193#_M1057_g 0.0280685f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_55 VNB N_A_967_193#_M1010_g 0.0240584f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.835
cc_56 VNB N_A_967_193#_c_795_n 0.0204883f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.91
cc_57 VNB N_A_967_193#_c_796_n 0.0431905f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_58 VNB N_A_967_193#_c_797_n 0.0723197f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_59 VNB N_A_967_193#_c_798_n 0.00748168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_967_193#_c_799_n 0.0907745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_967_193#_c_800_n 0.0101614f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.48
cc_62 VNB N_A_967_193#_M1045_g 0.0466158f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.035
cc_63 VNB N_A_967_193#_c_802_n 0.0721582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_967_193#_c_803_n 0.120142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_967_193#_c_804_n 0.0142074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_967_193#_c_805_n 0.00573649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_967_193#_c_806_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_967_193#_c_807_n 0.0164608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_967_193#_c_808_n 0.00216389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_967_193#_c_809_n 0.00227379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_967_193#_c_810_n 0.00110214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_967_193#_c_811_n 0.00374636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_967_193#_c_812_n 0.0424081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_967_193#_c_813_n 0.0187804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_967_193#_c_814_n 0.0358788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_967_193#_c_815_n 0.0112558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_967_193#_c_816_n 0.0391275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_967_193#_c_817_n 0.0048278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_967_193#_c_818_n 0.0407603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1147_490#_c_1091_n 0.0119755f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=1.985
cc_81 VNB N_A_1147_490#_c_1092_n 0.0295801f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=2.775
cc_82 VNB N_A_1147_490#_c_1093_n 0.00610893f $X=-0.19 $Y=-0.245 $X2=0.7
+ $Y2=1.315
cc_83 VNB N_A_1147_490#_c_1094_n 0.0102175f $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.835
cc_84 VNB N_A_1147_490#_c_1095_n 0.00266884f $X=-0.19 $Y=-0.245 $X2=0.73
+ $Y2=1.985
cc_85 VNB N_A_1147_490#_c_1096_n 0.00837414f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.48
cc_86 VNB N_A_1147_490#_c_1097_n 0.00646202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1147_490#_c_1098_n 0.00392709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1147_490#_c_1099_n 0.0384985f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=2.035
cc_89 VNB N_A_1147_490#_c_1100_n 0.0125507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1147_490#_c_1101_n 0.00513107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1147_490#_c_1102_n 0.0196487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_RESET_B_c_1285_n 0.0112712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_RESET_B_c_1286_n 0.00546427f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.985
cc_94 VNB N_RESET_B_M1041_g 0.009716f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.315
cc_95 VNB N_RESET_B_c_1288_n 0.210326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_RESET_B_c_1289_n 0.0125079f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.985
cc_97 VNB N_RESET_B_M1005_g 0.0611446f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_98 VNB N_RESET_B_M1054_g 0.0477572f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.835
cc_99 VNB N_RESET_B_c_1292_n 0.0196523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_RESET_B_c_1293_n 0.0476797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_RESET_B_c_1294_n 0.0335004f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.035
cc_102 VNB N_RESET_B_c_1295_n 0.00415515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_RESET_B_c_1296_n 0.00698333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_RESET_B_c_1297_n 0.0164615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_RESET_B_c_1298_n 0.0043602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_911_219#_c_1543_n 0.0271963f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=0.445
cc_107 VNB N_A_911_219#_M1000_g 0.0296715f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.775
cc_108 VNB N_A_911_219#_M1002_g 0.00570057f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.91
cc_109 VNB N_A_911_219#_c_1546_n 0.00536358f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=1.515
cc_110 VNB N_A_911_219#_M1021_g 0.0277621f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=2.775
cc_111 VNB N_A_911_219#_M1009_g 0.00430441f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.465
cc_112 VNB N_A_911_219#_c_1549_n 0.0050554f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.91
cc_113 VNB N_A_911_219#_c_1550_n 0.00524433f $X=-0.19 $Y=-0.245 $X2=0.73
+ $Y2=1.835
cc_114 VNB N_A_911_219#_c_1551_n 0.00828387f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_115 VNB N_A_911_219#_c_1552_n 0.00434769f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.48
cc_116 VNB N_A_911_219#_c_1553_n 0.00778581f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.295
cc_117 VNB N_A_911_219#_c_1554_n 0.0221702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_911_219#_c_1555_n 0.00406733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_911_219#_c_1556_n 0.00266631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_911_219#_c_1557_n 0.0271371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_2388_115#_c_1729_n 0.0148867f $X=-0.19 $Y=-0.245 $X2=0.55
+ $Y2=2.775
cc_122 VNB N_A_2388_115#_c_1730_n 0.00229106f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.91
cc_123 VNB N_A_2388_115#_c_1731_n 0.00361641f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=2.775
cc_124 VNB N_A_2388_115#_c_1732_n 5.57369e-19 $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=2.775
cc_125 VNB N_A_2388_115#_c_1733_n 0.0032665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2388_115#_c_1734_n 0.00235012f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.48
cc_127 VNB N_A_2388_115#_c_1735_n 0.00551292f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.665
cc_128 VNB N_A_2388_115#_c_1736_n 0.0579734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_2168_439#_c_1839_n 0.0182525f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=0.445
cc_130 VNB N_A_2168_439#_c_1840_n 0.0166376f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.775
cc_131 VNB N_A_2168_439#_c_1841_n 0.00980698f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.775
cc_132 VNB N_A_2168_439#_M1019_g 0.00721443f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.91
cc_133 VNB N_A_2168_439#_M1046_g 0.0181004f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=1.985
cc_134 VNB N_A_2168_439#_M1033_g 9.19169e-19 $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.465
cc_135 VNB N_A_2168_439#_M1031_g 0.0225459f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.91
cc_136 VNB N_A_2168_439#_M1007_g 9.92454e-19 $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_137 VNB N_A_2168_439#_c_1847_n 0.0592042f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_138 VNB N_A_2168_439#_M1022_g 0.0212901f $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.48
cc_139 VNB N_A_2168_439#_M1034_g 0.0136618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_2168_439#_c_1850_n 0.005583f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.48
cc_141 VNB N_A_2168_439#_M1001_g 0.0197152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_2168_439#_M1039_g 0.010806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_2168_439#_c_1853_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_2168_439#_c_1854_n 0.00524817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_2168_439#_c_1855_n 0.00601219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_A_2168_439#_c_1856_n 0.00857001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_2168_439#_c_1857_n 0.0203296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_A_2168_439#_c_1858_n 0.00493283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_2168_439#_c_1859_n 0.00431825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_A_2168_439#_c_1860_n 0.00970901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_A_2168_439#_c_1861_n 0.00440443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_A_2168_439#_c_1862_n 0.0176661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_2168_439#_c_1863_n 0.00365072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_2168_439#_c_1864_n 0.00223777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_A_2168_439#_c_1865_n 0.00160603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_A_2168_439#_c_1866_n 0.0385654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_A_2168_439#_c_1867_n 0.0302823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_CLK_M1026_g 0.0218178f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_159 VNB N_CLK_M1027_g 0.0208567f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.445
cc_160 VNB N_CLK_c_2085_n 5.67477e-19 $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_161 VNB N_CLK_c_2086_n 0.0287318f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_162 VNB N_A_3416_137#_M1012_g 0.0226389f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=1.315
cc_163 VNB N_A_3416_137#_M1053_g 0.00101744f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=1.985
cc_164 VNB N_A_3416_137#_M1020_g 0.0249073f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=1.91
cc_165 VNB N_A_3416_137#_M1058_g 0.00112085f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=1.515
cc_166 VNB N_A_3416_137#_c_2133_n 0.0093481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_A_3416_137#_c_2134_n 2.41884e-19 $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.835
cc_168 VNB N_A_3416_137#_c_2135_n 0.020007f $X=-0.19 $Y=-0.245 $X2=1.635
+ $Y2=1.91
cc_169 VNB N_A_3416_137#_c_2136_n 0.00212516f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_170 VNB N_A_3416_137#_c_2137_n 0.0378831f $X=-0.19 $Y=-0.245 $X2=0.722
+ $Y2=1.48
cc_171 VNB N_VPWR_c_2191_n 0.800558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_A_342_261#_c_2407_n 0.0134526f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.775
cc_173 VNB N_A_342_261#_c_2408_n 0.0134814f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.775
cc_174 VNB N_A_342_261#_c_2409_n 0.00425636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_A_342_261#_c_2410_n 0.00656037f $X=-0.19 $Y=-0.245 $X2=1.56
+ $Y2=1.91
cc_176 VNB N_A_342_261#_c_2411_n 6.91649e-19 $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.91
cc_177 VNB N_A_342_261#_c_2412_n 0.00843042f $X=-0.19 $Y=-0.245 $X2=0.7
+ $Y2=1.315
cc_178 VNB N_A_342_261#_c_2413_n 4.85034e-19 $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_179 VNB N_A_342_261#_c_2414_n 0.00822935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_A_342_261#_c_2415_n 0.00228872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_A_342_261#_c_2416_n 0.00570885f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.48
cc_182 VNB N_A_342_261#_c_2417_n 0.00244626f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.295
cc_183 VNB N_Q_N_c_2631_n 0.00575777f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.775
cc_184 VNB N_Q_N_c_2632_n 0.01497f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_185 VNB Q_N 0.00356222f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.835
cc_186 VNB N_Q_c_2665_n 0.0567461f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.985
cc_187 VNB N_VGND_c_2681_n 0.00659109f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.775
cc_188 VNB N_VGND_c_2682_n 0.00410504f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.465
cc_189 VNB N_VGND_c_2683_n 0.0075011f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.985
cc_190 VNB N_VGND_c_2684_n 0.00715016f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_191 VNB N_VGND_c_2685_n 0.013655f $X=-0.19 $Y=-0.245 $X2=0.722 $Y2=1.48
cc_192 VNB N_VGND_c_2686_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_193 VNB N_VGND_c_2687_n 0.0197306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_194 VNB N_VGND_c_2688_n 0.0795114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_195 VNB N_VGND_c_2689_n 0.00478044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_196 VNB N_VGND_c_2690_n 0.0761013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_197 VNB N_VGND_c_2691_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_198 VNB N_VGND_c_2692_n 0.0262771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_199 VNB N_VGND_c_2693_n 0.0545609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_200 VNB N_VGND_c_2694_n 0.03929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_201 VNB N_VGND_c_2695_n 0.0825606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_202 VNB N_VGND_c_2696_n 0.0552379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_203 VNB N_VGND_c_2697_n 0.0270669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_204 VNB N_VGND_c_2698_n 0.935355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_205 VNB N_VGND_c_2699_n 0.0051053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_206 VNB N_VGND_c_2700_n 0.00324297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_207 VNB N_VGND_c_2701_n 0.00631443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_208 VNB N_VGND_c_2702_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_209 VNB N_VGND_c_2703_n 0.00536178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_210 VNB N_noxref_37_c_2854_n 0.00108592f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=1.315
cc_211 VNB N_noxref_37_c_2855_n 0.0203054f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=0.445
cc_212 VNB N_noxref_37_c_2856_n 2.77498e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_213 VNB N_noxref_37_c_2857_n 4.24544e-19 $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.775
cc_214 VNB N_noxref_39_c_2888_n 6.47547e-19 $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=1.315
cc_215 VNB N_noxref_39_c_2889_n 0.0274046f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=0.445
cc_216 VNB N_noxref_39_c_2890_n 0.0018464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_217 VNB N_noxref_39_c_2891_n 0.00846169f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.775
cc_218 VNB N_noxref_39_c_2892_n 0.00440851f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.775
cc_219 VNB N_noxref_39_c_2893_n 0.00809854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_220 VNB N_noxref_39_c_2894_n 0.00635915f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.91
cc_221 VNB N_A_824_219#_c_2941_n 0.021156f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.775
cc_222 VNB N_A_824_219#_c_2942_n 0.00991743f $X=-0.19 $Y=-0.245 $X2=0.895
+ $Y2=0.445
cc_223 VNB N_A_824_219#_c_2943_n 0.00992762f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=1.985
cc_224 VNB N_A_824_219#_c_2944_n 0.0190045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_225 VPB N_SCE_M1024_g 0.0382552f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.775
cc_226 VPB N_SCE_M1016_g 0.0285513f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.775
cc_227 VPB N_SCE_M1013_g 0.0222092f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=2.775
cc_228 VPB N_SCE_c_386_n 0.0121278f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.91
cc_229 VPB SCE 0.00826956f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_230 VPB N_SCE_c_389_n 0.0132738f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.48
cc_231 VPB N_D_M1014_g 0.0187279f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.445
cc_232 VPB N_A_29_47#_M1056_g 0.0187279f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.985
cc_233 VPB N_A_29_47#_c_510_n 0.0331156f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=2.775
cc_234 VPB N_A_29_47#_c_505_n 0.0372245f $X=-0.19 $Y=1.655 $X2=0.722 $Y2=1.835
cc_235 VPB N_SCD_M1023_g 0.0221582f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.445
cc_236 VPB N_A_876_93#_M1032_g 0.0201788f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.315
cc_237 VPB N_A_876_93#_M1044_g 0.0338692f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.775
cc_238 VPB N_A_876_93#_c_629_n 0.00153036f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.295
cc_239 VPB N_A_876_93#_c_621_n 0.00411147f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.665
cc_240 VPB N_A_876_93#_c_625_n 0.00463285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_876_93#_c_626_n 0.0126347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_967_193#_M1028_g 0.0245106f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.985
cc_243 VPB N_A_967_193#_c_791_n 0.00625887f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.775
cc_244 VPB N_A_967_193#_M1025_g 0.0209141f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.835
cc_245 VPB N_A_967_193#_M1029_g 0.020201f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.315
cc_246 VPB N_A_967_193#_c_796_n 0.0096014f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_247 VPB N_A_967_193#_c_798_n 0.0721304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_967_193#_c_825_n 0.0760119f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.48
cc_249 VPB N_A_967_193#_c_826_n 0.010539f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.48
cc_250 VPB N_A_967_193#_M1042_g 0.0314211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_967_193#_c_828_n 0.0279518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_967_193#_c_829_n 0.0223695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_967_193#_c_830_n 0.0170956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_967_193#_c_831_n 0.00353434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_967_193#_c_832_n 0.00337873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_967_193#_c_809_n 0.00674171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_967_193#_c_810_n 0.0162832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_967_193#_c_835_n 0.00276398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_967_193#_c_836_n 0.0358979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_1147_490#_c_1103_n 0.0205592f $X=-0.19 $Y=1.655 $X2=0.91
+ $Y2=1.985
cc_261 VPB N_A_1147_490#_c_1104_n 0.0365855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_1147_490#_c_1105_n 0.00773051f $X=-0.19 $Y=1.655 $X2=1.56
+ $Y2=1.91
cc_263 VPB N_A_1147_490#_c_1091_n 0.0428302f $X=-0.19 $Y=1.655 $X2=1.635
+ $Y2=1.985
cc_264 VPB N_A_1147_490#_c_1093_n 0.00780911f $X=-0.19 $Y=1.655 $X2=0.7
+ $Y2=1.315
cc_265 VPB N_A_1147_490#_c_1095_n 0.00145711f $X=-0.19 $Y=1.655 $X2=0.73
+ $Y2=1.985
cc_266 VPB N_A_1147_490#_c_1109_n 0.00310275f $X=-0.19 $Y=1.655 $X2=1.635
+ $Y2=1.91
cc_267 VPB N_A_1147_490#_c_1110_n 0.00531952f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.95
cc_268 VPB N_A_1147_490#_c_1111_n 0.00847087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_1147_490#_c_1112_n 0.00182831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_1147_490#_c_1097_n 0.00443429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_1147_490#_c_1114_n 0.00752496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_RESET_B_c_1299_n 0.0175807f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.315
cc_273 VPB N_RESET_B_c_1285_n 0.00291892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_RESET_B_c_1286_n 0.00265092f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.985
cc_275 VPB N_RESET_B_c_1302_n 0.0177364f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.775
cc_276 VPB N_RESET_B_M1043_g 0.0207205f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.835
cc_277 VPB N_RESET_B_M1005_g 0.0366256f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=2.775
cc_278 VPB N_RESET_B_M1049_g 0.021858f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.315
cc_279 VPB N_RESET_B_c_1306_n 0.02022f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_280 VPB N_RESET_B_M1038_g 0.0208833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_RESET_B_M1036_g 0.0173269f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.48
cc_282 VPB N_RESET_B_c_1295_n 0.00698135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_RESET_B_c_1296_n 0.0148719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_RESET_B_c_1311_n 0.0213405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_RESET_B_c_1312_n 0.00144101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_RESET_B_c_1313_n 0.0347729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_RESET_B_c_1314_n 0.00152042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_RESET_B_c_1315_n 0.00327586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_RESET_B_c_1316_n 0.00697491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_RESET_B_c_1298_n 0.00119617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_RESET_B_c_1318_n 0.0429202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_RESET_B_c_1319_n 7.91879e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_RESET_B_c_1320_n 0.0446132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_A_911_219#_M1002_g 0.0233131f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.91
cc_295 VPB N_A_911_219#_M1009_g 0.0222093f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.465
cc_296 VPB N_A_911_219#_c_1560_n 0.00227434f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.21
cc_297 VPB N_A_911_219#_c_1561_n 0.00365117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_A_911_219#_c_1562_n 0.00106796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_A_911_219#_c_1553_n 0.00286291f $X=-0.19 $Y=1.655 $X2=0.64
+ $Y2=1.295
cc_300 VPB N_A_911_219#_c_1554_n 0.0129652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_A_911_219#_c_1565_n 0.00607507f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.48
cc_302 VPB N_A_911_219#_c_1566_n 0.00210331f $X=-0.19 $Y=1.655 $X2=0.64
+ $Y2=2.035
cc_303 VPB N_A_911_219#_c_1567_n 0.00100726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_A_911_219#_c_1568_n 0.0028892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_A_911_219#_c_1557_n 0.0140647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_A_2388_115#_M1018_g 0.0296496f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.775
cc_307 VPB N_A_2388_115#_c_1738_n 0.0117803f $X=-0.19 $Y=1.655 $X2=1.635
+ $Y2=1.515
cc_308 VPB N_A_2388_115#_c_1739_n 0.00271537f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=1.835
cc_309 VPB N_A_2388_115#_c_1740_n 0.00417204f $X=-0.19 $Y=1.655 $X2=0.73
+ $Y2=1.985
cc_310 VPB N_A_2388_115#_c_1741_n 0.037529f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.91
cc_311 VPB N_A_2388_115#_c_1735_n 0.0350336f $X=-0.19 $Y=1.655 $X2=0.64
+ $Y2=1.665
cc_312 VPB N_A_2168_439#_M1037_g 0.020992f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.315
cc_313 VPB N_A_2168_439#_M1019_g 0.0694152f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.91
cc_314 VPB N_A_2168_439#_M1033_g 0.019089f $X=-0.19 $Y=1.655 $X2=0.722 $Y2=1.465
cc_315 VPB N_A_2168_439#_M1007_g 0.0230552f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_316 VPB N_A_2168_439#_M1034_g 0.0237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_317 VPB N_A_2168_439#_M1039_g 0.0219563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_318 VPB N_A_2168_439#_c_1874_n 0.00733911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_319 VPB N_A_2168_439#_c_1856_n 0.00264111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_320 VPB N_A_2168_439#_c_1876_n 0.0112317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_321 VPB N_A_2168_439#_c_1877_n 0.016437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_A_2168_439#_c_1857_n 0.0176511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_A_2168_439#_c_1879_n 8.16291e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_A_2168_439#_c_1880_n 0.00299687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_CLK_M1052_g 0.0225181f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.775
cc_326 VPB N_CLK_M1055_g 0.0165343f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.775
cc_327 VPB N_CLK_c_2085_n 0.00889399f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=2.775
cc_328 VPB N_CLK_c_2086_n 0.00362791f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=2.775
cc_329 VPB N_A_3416_137#_M1053_g 0.0215386f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.985
cc_330 VPB N_A_3416_137#_M1058_g 0.0234886f $X=-0.19 $Y=1.655 $X2=1.635
+ $Y2=1.515
cc_331 VPB N_A_3416_137#_c_2134_n 0.0143873f $X=-0.19 $Y=1.655 $X2=0.722
+ $Y2=1.835
cc_332 VPB N_VPWR_c_2192_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.315
cc_333 VPB N_VPWR_c_2193_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.835
cc_334 VPB N_VPWR_c_2194_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_335 VPB N_VPWR_c_2195_n 0.00785303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_2196_n 0.00921575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_2197_n 0.00439506f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.035
cc_338 VPB N_VPWR_c_2198_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_2199_n 0.0256831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_2200_n 0.0696723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_2201_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_342 VPB N_VPWR_c_2202_n 0.0420545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_2203_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_2204_n 0.0282044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_2205_n 0.0469379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_346 VPB N_VPWR_c_2206_n 0.072686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_347 VPB N_VPWR_c_2207_n 0.0771899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_348 VPB N_VPWR_c_2208_n 0.0305844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_349 VPB N_VPWR_c_2209_n 0.0574501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_350 VPB N_VPWR_c_2210_n 0.0268694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_351 VPB N_VPWR_c_2191_n 0.170508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_352 VPB N_VPWR_c_2212_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_353 VPB N_VPWR_c_2213_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_354 VPB N_VPWR_c_2214_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_355 VPB N_VPWR_c_2215_n 0.00631846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_356 VPB N_VPWR_c_2216_n 0.00421541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_357 VPB N_VPWR_c_2217_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_358 VPB N_A_342_261#_c_2410_n 0.019121f $X=-0.19 $Y=1.655 $X2=1.56 $Y2=1.91
cc_359 VPB N_A_342_261#_c_2411_n 0.00187622f $X=-0.19 $Y=1.655 $X2=0.985
+ $Y2=1.91
cc_360 VPB N_A_342_261#_c_2412_n 0.0176236f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.315
cc_361 VPB N_A_342_261#_c_2421_n 0.00175918f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.91
cc_362 VPB N_A_342_261#_c_2422_n 6.25841e-19 $X=-0.19 $Y=1.655 $X2=0.73
+ $Y2=1.835
cc_363 VPB N_A_342_261#_c_2413_n 7.4181e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_364 VPB N_A_2081_439#_c_2552_n 0.00404153f $X=-0.19 $Y=1.655 $X2=0.895
+ $Y2=1.315
cc_365 VPB N_A_2081_439#_c_2553_n 8.6014e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_366 VPB N_A_2081_439#_c_2554_n 0.00212228f $X=-0.19 $Y=1.655 $X2=0.91
+ $Y2=2.775
cc_367 VPB N_A_2081_439#_c_2555_n 0.0175054f $X=-0.19 $Y=1.655 $X2=0.91
+ $Y2=2.775
cc_368 VPB N_A_2523_397#_c_2582_n 0.00433473f $X=-0.19 $Y=1.655 $X2=0.55
+ $Y2=2.775
cc_369 VPB N_A_2523_397#_c_2583_n 0.00222373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_370 VPB N_A_2523_397#_c_2584_n 0.026297f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.985
cc_371 VPB N_A_2523_397#_c_2585_n 0.00137688f $X=-0.19 $Y=1.655 $X2=0.91
+ $Y2=2.775
cc_372 VPB N_A_2523_397#_c_2586_n 0.00537743f $X=-0.19 $Y=1.655 $X2=0.985
+ $Y2=1.91
cc_373 VPB N_A_2523_397#_c_2587_n 0.0149405f $X=-0.19 $Y=1.655 $X2=1.635
+ $Y2=1.835
cc_374 VPB N_Q_N_c_2634_n 0.00580357f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.315
cc_375 VPB N_Q_N_c_2635_n 0.0264434f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=0.445
cc_376 VPB N_Q_N_c_2631_n 0.00305138f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.775
cc_377 VPB N_Q_c_2665_n 0.0543794f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.985
cc_378 N_SCE_M1013_g N_D_M1014_g 0.0376119f $X=1.635 $Y=2.775 $X2=0 $Y2=0
cc_379 N_SCE_c_383_n N_D_M1059_g 0.0145734f $X=1.635 $Y=1.835 $X2=0 $Y2=0
cc_380 N_SCE_c_387_n N_D_c_453_n 0.0376119f $X=1.635 $Y=1.91 $X2=0 $Y2=0
cc_381 N_SCE_M1040_g N_A_29_47#_c_503_n 0.00924054f $X=0.505 $Y=0.445 $X2=0
+ $Y2=0
cc_382 N_SCE_M1017_g N_A_29_47#_c_503_n 0.00165355f $X=0.895 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_SCE_M1024_g N_A_29_47#_c_510_n 0.01578f $X=0.55 $Y=2.775 $X2=0 $Y2=0
cc_384 N_SCE_M1016_g N_A_29_47#_c_510_n 0.00184939f $X=0.91 $Y=2.775 $X2=0 $Y2=0
cc_385 SCE N_A_29_47#_c_510_n 0.00127591f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_386 N_SCE_M1040_g N_A_29_47#_c_504_n 0.00500826f $X=0.505 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_SCE_M1040_g N_A_29_47#_c_505_n 0.015297f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_388 SCE N_A_29_47#_c_505_n 0.069684f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_389 N_SCE_c_389_n N_A_29_47#_c_505_n 0.0239167f $X=0.64 $Y=1.48 $X2=0 $Y2=0
cc_390 N_SCE_M1040_g N_A_29_47#_c_508_n 0.00953507f $X=0.505 $Y=0.445 $X2=0
+ $Y2=0
cc_391 N_SCE_M1017_g N_A_29_47#_c_508_n 0.018233f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_392 N_SCE_c_383_n N_A_29_47#_c_508_n 8.03683e-19 $X=1.635 $Y=1.835 $X2=0
+ $Y2=0
cc_393 N_SCE_c_385_n N_A_29_47#_c_508_n 2.86294e-19 $X=0.7 $Y=1.465 $X2=0 $Y2=0
cc_394 SCE N_A_29_47#_c_508_n 0.017973f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_395 N_SCE_M1024_g N_VPWR_c_2192_n 0.00283343f $X=0.55 $Y=2.775 $X2=0 $Y2=0
cc_396 N_SCE_M1016_g N_VPWR_c_2192_n 0.0194416f $X=0.91 $Y=2.775 $X2=0 $Y2=0
cc_397 N_SCE_c_382_n N_VPWR_c_2192_n 5.59578e-19 $X=1.56 $Y=1.91 $X2=0 $Y2=0
cc_398 N_SCE_M1013_g N_VPWR_c_2192_n 0.016003f $X=1.635 $Y=2.775 $X2=0 $Y2=0
cc_399 N_SCE_M1024_g N_VPWR_c_2204_n 0.00549284f $X=0.55 $Y=2.775 $X2=0 $Y2=0
cc_400 N_SCE_M1016_g N_VPWR_c_2204_n 0.00486043f $X=0.91 $Y=2.775 $X2=0 $Y2=0
cc_401 N_SCE_M1013_g N_VPWR_c_2205_n 0.00585385f $X=1.635 $Y=2.775 $X2=0 $Y2=0
cc_402 N_SCE_M1024_g N_VPWR_c_2191_n 0.0109537f $X=0.55 $Y=2.775 $X2=0 $Y2=0
cc_403 N_SCE_M1016_g N_VPWR_c_2191_n 0.00814425f $X=0.91 $Y=2.775 $X2=0 $Y2=0
cc_404 N_SCE_M1013_g N_VPWR_c_2191_n 0.0115332f $X=1.635 $Y=2.775 $X2=0 $Y2=0
cc_405 N_SCE_M1017_g N_A_342_261#_c_2407_n 0.00834554f $X=0.895 $Y=0.445 $X2=0
+ $Y2=0
cc_406 N_SCE_M1016_g N_A_342_261#_c_2407_n 0.00187868f $X=0.91 $Y=2.775 $X2=0
+ $Y2=0
cc_407 N_SCE_c_382_n N_A_342_261#_c_2407_n 0.0110496f $X=1.56 $Y=1.91 $X2=0
+ $Y2=0
cc_408 N_SCE_c_383_n N_A_342_261#_c_2407_n 0.00198037f $X=1.635 $Y=1.835 $X2=0
+ $Y2=0
cc_409 N_SCE_M1013_g N_A_342_261#_c_2407_n 0.00279472f $X=1.635 $Y=2.775 $X2=0
+ $Y2=0
cc_410 SCE N_A_342_261#_c_2407_n 0.0657768f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_411 N_SCE_c_382_n N_A_342_261#_c_2408_n 0.00435107f $X=1.56 $Y=1.91 $X2=0
+ $Y2=0
cc_412 N_SCE_c_383_n N_A_342_261#_c_2408_n 0.00835307f $X=1.635 $Y=1.835 $X2=0
+ $Y2=0
cc_413 N_SCE_M1017_g N_A_342_261#_c_2409_n 0.00625176f $X=0.895 $Y=0.445 $X2=0
+ $Y2=0
cc_414 SCE N_A_342_261#_c_2409_n 0.00466823f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_415 N_SCE_c_382_n N_A_342_261#_c_2410_n 0.00883484f $X=1.56 $Y=1.91 $X2=0
+ $Y2=0
cc_416 N_SCE_M1013_g N_A_342_261#_c_2410_n 0.0160108f $X=1.635 $Y=2.775 $X2=0
+ $Y2=0
cc_417 N_SCE_M1024_g N_A_342_261#_c_2411_n 7.82533e-19 $X=0.55 $Y=2.775 $X2=0
+ $Y2=0
cc_418 N_SCE_M1016_g N_A_342_261#_c_2411_n 0.00628326f $X=0.91 $Y=2.775 $X2=0
+ $Y2=0
cc_419 SCE N_A_342_261#_c_2411_n 4.01705e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_420 N_SCE_c_383_n N_A_342_261#_c_2439_n 0.00680959f $X=1.635 $Y=1.835 $X2=0
+ $Y2=0
cc_421 N_SCE_M1013_g N_A_342_261#_c_2440_n 0.00371475f $X=1.635 $Y=2.775 $X2=0
+ $Y2=0
cc_422 N_SCE_M1040_g N_VGND_c_2681_n 0.00200074f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_423 N_SCE_M1017_g N_VGND_c_2681_n 0.0112286f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_424 N_SCE_M1040_g N_VGND_c_2692_n 0.00425202f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_425 N_SCE_M1017_g N_VGND_c_2692_n 0.00362954f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_426 N_SCE_M1040_g N_VGND_c_2698_n 0.00699576f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_427 N_SCE_M1017_g N_VGND_c_2698_n 0.00423997f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_428 N_SCE_c_383_n N_noxref_37_c_2854_n 0.00188255f $X=1.635 $Y=1.835 $X2=0
+ $Y2=0
cc_429 N_SCE_c_382_n N_noxref_37_c_2855_n 0.00139094f $X=1.56 $Y=1.91 $X2=0
+ $Y2=0
cc_430 N_SCE_c_383_n N_noxref_37_c_2855_n 0.005155f $X=1.635 $Y=1.835 $X2=0
+ $Y2=0
cc_431 N_SCE_c_387_n N_noxref_37_c_2855_n 0.00528237f $X=1.635 $Y=1.91 $X2=0
+ $Y2=0
cc_432 N_SCE_c_382_n N_noxref_37_c_2856_n 0.00819162f $X=1.56 $Y=1.91 $X2=0
+ $Y2=0
cc_433 N_D_c_453_n N_A_29_47#_M1004_g 0.0431201f $X=2.045 $Y=1.985 $X2=0 $Y2=0
cc_434 N_D_M1014_g N_A_29_47#_M1056_g 0.0400038f $X=2.025 $Y=2.775 $X2=0 $Y2=0
cc_435 N_D_M1059_g N_A_29_47#_c_506_n 0.00237323f $X=2.065 $Y=1.515 $X2=0 $Y2=0
cc_436 N_D_c_454_n N_A_29_47#_c_506_n 0.0258204f $X=3.005 $Y=0.35 $X2=0 $Y2=0
cc_437 N_D_c_457_n N_A_29_47#_c_506_n 0.00259977f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_438 N_D_M1059_g N_A_29_47#_c_507_n 0.0431201f $X=2.065 $Y=1.515 $X2=0 $Y2=0
cc_439 N_D_c_454_n N_A_29_47#_c_507_n 0.00821905f $X=3.005 $Y=0.35 $X2=0 $Y2=0
cc_440 N_D_c_457_n N_A_29_47#_c_507_n 0.00136304f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_441 N_D_M1059_g N_A_29_47#_c_508_n 0.0160152f $X=2.065 $Y=1.515 $X2=0 $Y2=0
cc_442 N_D_c_454_n N_A_29_47#_c_508_n 0.00855343f $X=3.005 $Y=0.35 $X2=0 $Y2=0
cc_443 N_D_c_455_n N_A_29_47#_c_508_n 0.00484599f $X=1.945 $Y=0.4 $X2=0 $Y2=0
cc_444 N_D_c_456_n N_A_29_47#_c_508_n 0.0219045f $X=2.11 $Y=0.4 $X2=0 $Y2=0
cc_445 N_D_c_457_n N_RESET_B_M1041_g 0.00225899f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_446 N_D_M1014_g N_VPWR_c_2205_n 0.00549284f $X=2.025 $Y=2.775 $X2=0 $Y2=0
cc_447 N_D_M1014_g N_VPWR_c_2191_n 0.0100377f $X=2.025 $Y=2.775 $X2=0 $Y2=0
cc_448 N_D_M1059_g N_A_342_261#_c_2408_n 0.00643292f $X=2.065 $Y=1.515 $X2=0
+ $Y2=0
cc_449 N_D_M1014_g N_A_342_261#_c_2410_n 0.0109043f $X=2.025 $Y=2.775 $X2=0
+ $Y2=0
cc_450 N_D_M1059_g N_A_342_261#_c_2439_n 0.00717352f $X=2.065 $Y=1.515 $X2=0
+ $Y2=0
cc_451 N_D_M1014_g N_A_342_261#_c_2440_n 0.0176967f $X=2.025 $Y=2.775 $X2=0
+ $Y2=0
cc_452 N_D_M1014_g N_A_342_261#_c_2417_n 0.00275687f $X=2.025 $Y=2.775 $X2=0
+ $Y2=0
cc_453 N_D_c_453_n N_A_342_261#_c_2417_n 0.00110934f $X=2.045 $Y=1.985 $X2=0
+ $Y2=0
cc_454 N_D_c_455_n N_VGND_c_2681_n 0.00235376f $X=1.945 $Y=0.4 $X2=0 $Y2=0
cc_455 N_D_c_456_n N_VGND_c_2681_n 0.00970699f $X=2.11 $Y=0.4 $X2=0 $Y2=0
cc_456 N_D_c_457_n N_VGND_c_2682_n 0.0169046f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_457 N_D_c_455_n N_VGND_c_2693_n 0.00603332f $X=1.945 $Y=0.4 $X2=0 $Y2=0
cc_458 N_D_c_456_n N_VGND_c_2693_n 0.0738992f $X=2.11 $Y=0.4 $X2=0 $Y2=0
cc_459 N_D_c_457_n N_VGND_c_2693_n 0.014793f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_460 N_D_c_455_n N_VGND_c_2698_n 0.00780108f $X=1.945 $Y=0.4 $X2=0 $Y2=0
cc_461 N_D_c_456_n N_VGND_c_2698_n 0.0443932f $X=2.11 $Y=0.4 $X2=0 $Y2=0
cc_462 N_D_c_457_n N_VGND_c_2698_n 0.00870292f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_463 N_D_M1059_g N_noxref_37_c_2855_n 0.00723073f $X=2.065 $Y=1.515 $X2=0
+ $Y2=0
cc_464 N_D_c_453_n N_noxref_37_c_2855_n 0.007716f $X=2.045 $Y=1.985 $X2=0 $Y2=0
cc_465 N_D_M1059_g N_noxref_39_c_2888_n 0.0010357f $X=2.065 $Y=1.515 $X2=0 $Y2=0
cc_466 N_D_c_454_n N_noxref_39_c_2889_n 0.00845112f $X=3.005 $Y=0.35 $X2=0 $Y2=0
cc_467 N_D_c_457_n N_noxref_39_c_2889_n 0.0102857f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_468 N_D_M1059_g N_noxref_39_c_2890_n 4.60392e-19 $X=2.065 $Y=1.515 $X2=0
+ $Y2=0
cc_469 N_D_c_454_n N_noxref_39_c_2890_n 0.00149578f $X=3.005 $Y=0.35 $X2=0 $Y2=0
cc_470 N_D_c_457_n N_noxref_39_c_2894_n 0.00346687f $X=3.12 $Y=0.35 $X2=0 $Y2=0
cc_471 N_A_29_47#_M1056_g N_SCD_M1023_g 0.036868f $X=2.455 $Y=2.775 $X2=0 $Y2=0
cc_472 N_A_29_47#_M1004_g N_SCD_c_572_n 0.0141096f $X=2.425 $Y=1.515 $X2=0 $Y2=0
cc_473 N_A_29_47#_c_502_n N_SCD_c_574_n 0.036868f $X=2.44 $Y=1.985 $X2=0 $Y2=0
cc_474 N_A_29_47#_c_510_n N_VPWR_c_2192_n 0.019242f $X=0.312 $Y=2.622 $X2=0
+ $Y2=0
cc_475 N_A_29_47#_M1056_g N_VPWR_c_2193_n 0.00284989f $X=2.455 $Y=2.775 $X2=0
+ $Y2=0
cc_476 N_A_29_47#_c_510_n N_VPWR_c_2204_n 0.0227389f $X=0.312 $Y=2.622 $X2=0
+ $Y2=0
cc_477 N_A_29_47#_M1056_g N_VPWR_c_2205_n 0.00549284f $X=2.455 $Y=2.775 $X2=0
+ $Y2=0
cc_478 N_A_29_47#_M1024_s N_VPWR_c_2191_n 0.00232985f $X=0.19 $Y=2.455 $X2=0
+ $Y2=0
cc_479 N_A_29_47#_M1056_g N_VPWR_c_2191_n 0.0100377f $X=2.455 $Y=2.775 $X2=0
+ $Y2=0
cc_480 N_A_29_47#_c_510_n N_VPWR_c_2191_n 0.0143009f $X=0.312 $Y=2.622 $X2=0
+ $Y2=0
cc_481 N_A_29_47#_M1004_g N_A_342_261#_c_2408_n 4.60392e-19 $X=2.425 $Y=1.515
+ $X2=0 $Y2=0
cc_482 N_A_29_47#_c_508_n N_A_342_261#_c_2408_n 0.0643575f $X=2.295 $Y=0.75
+ $X2=0 $Y2=0
cc_483 N_A_29_47#_c_508_n N_A_342_261#_c_2409_n 0.0137879f $X=2.295 $Y=0.75
+ $X2=0 $Y2=0
cc_484 N_A_29_47#_M1004_g N_A_342_261#_c_2439_n 0.00103345f $X=2.425 $Y=1.515
+ $X2=0 $Y2=0
cc_485 N_A_29_47#_M1056_g N_A_342_261#_c_2440_n 0.0170571f $X=2.455 $Y=2.775
+ $X2=0 $Y2=0
cc_486 N_A_29_47#_M1056_g N_A_342_261#_c_2412_n 0.0109043f $X=2.455 $Y=2.775
+ $X2=0 $Y2=0
cc_487 N_A_29_47#_M1056_g N_A_342_261#_c_2417_n 0.00275687f $X=2.455 $Y=2.775
+ $X2=0 $Y2=0
cc_488 N_A_29_47#_c_502_n N_A_342_261#_c_2417_n 8.32005e-19 $X=2.44 $Y=1.985
+ $X2=0 $Y2=0
cc_489 N_A_29_47#_c_503_n N_VGND_c_2681_n 0.00855378f $X=0.29 $Y=0.47 $X2=0
+ $Y2=0
cc_490 N_A_29_47#_c_508_n N_VGND_c_2681_n 0.0221837f $X=2.295 $Y=0.75 $X2=0
+ $Y2=0
cc_491 N_A_29_47#_c_503_n N_VGND_c_2692_n 0.0197437f $X=0.29 $Y=0.47 $X2=0 $Y2=0
cc_492 N_A_29_47#_c_508_n N_VGND_c_2692_n 0.00711987f $X=2.295 $Y=0.75 $X2=0
+ $Y2=0
cc_493 N_A_29_47#_c_508_n N_VGND_c_2693_n 0.00782034f $X=2.295 $Y=0.75 $X2=0
+ $Y2=0
cc_494 N_A_29_47#_M1040_s N_VGND_c_2698_n 0.00232985f $X=0.145 $Y=0.235 $X2=0
+ $Y2=0
cc_495 N_A_29_47#_c_503_n N_VGND_c_2698_n 0.0125654f $X=0.29 $Y=0.47 $X2=0 $Y2=0
cc_496 N_A_29_47#_c_508_n N_VGND_c_2698_n 0.0278757f $X=2.295 $Y=0.75 $X2=0
+ $Y2=0
cc_497 N_A_29_47#_M1004_g N_noxref_37_c_2855_n 0.00723073f $X=2.425 $Y=1.515
+ $X2=0 $Y2=0
cc_498 N_A_29_47#_c_502_n N_noxref_37_c_2855_n 0.00738826f $X=2.44 $Y=1.985
+ $X2=0 $Y2=0
cc_499 N_A_29_47#_M1004_g N_noxref_37_c_2857_n 8.13609e-19 $X=2.425 $Y=1.515
+ $X2=0 $Y2=0
cc_500 N_A_29_47#_M1004_g N_noxref_39_c_2888_n 0.00699586f $X=2.425 $Y=1.515
+ $X2=0 $Y2=0
cc_501 N_A_29_47#_M1004_g N_noxref_39_c_2890_n 0.00643292f $X=2.425 $Y=1.515
+ $X2=0 $Y2=0
cc_502 N_A_29_47#_c_506_n N_noxref_39_c_2890_n 0.0159383f $X=2.515 $Y=0.75 $X2=0
+ $Y2=0
cc_503 N_A_29_47#_c_507_n N_noxref_39_c_2890_n 0.00429058f $X=2.515 $Y=0.75
+ $X2=0 $Y2=0
cc_504 N_SCD_M1023_g N_RESET_B_c_1286_n 0.0115185f $X=2.845 $Y=2.775 $X2=0 $Y2=0
cc_505 SCD N_RESET_B_c_1286_n 0.00185458f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_506 N_SCD_c_576_n N_RESET_B_c_1286_n 0.00890713f $X=3.49 $Y=1.8 $X2=0 $Y2=0
cc_507 SCD N_RESET_B_c_1293_n 0.00485946f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_508 N_SCD_c_576_n N_RESET_B_c_1297_n 0.0220935f $X=3.49 $Y=1.8 $X2=0 $Y2=0
cc_509 SCD N_RESET_B_c_1298_n 0.0258623f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_510 N_SCD_c_576_n N_RESET_B_c_1298_n 5.41715e-19 $X=3.49 $Y=1.8 $X2=0 $Y2=0
cc_511 N_SCD_M1023_g N_VPWR_c_2193_n 0.0190607f $X=2.845 $Y=2.775 $X2=0 $Y2=0
cc_512 N_SCD_M1023_g N_VPWR_c_2205_n 0.00486043f $X=2.845 $Y=2.775 $X2=0 $Y2=0
cc_513 N_SCD_M1023_g N_VPWR_c_2191_n 0.00827383f $X=2.845 $Y=2.775 $X2=0 $Y2=0
cc_514 N_SCD_M1023_g N_A_342_261#_c_2440_n 0.0025027f $X=2.845 $Y=2.775 $X2=0
+ $Y2=0
cc_515 N_SCD_M1023_g N_A_342_261#_c_2412_n 0.0155704f $X=2.845 $Y=2.775 $X2=0
+ $Y2=0
cc_516 N_SCD_c_574_n N_A_342_261#_c_2412_n 0.0138067f $X=2.85 $Y=1.91 $X2=0
+ $Y2=0
cc_517 SCD N_A_342_261#_c_2412_n 0.0190561f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_518 N_SCD_c_576_n N_A_342_261#_c_2412_n 0.00320328f $X=3.49 $Y=1.8 $X2=0
+ $Y2=0
cc_519 N_SCD_M1023_g N_A_342_261#_c_2421_n 0.00324315f $X=2.845 $Y=2.775 $X2=0
+ $Y2=0
cc_520 N_SCD_c_572_n N_noxref_37_c_2855_n 0.00468987f $X=2.855 $Y=1.835 $X2=0
+ $Y2=0
cc_521 N_SCD_c_573_n N_noxref_37_c_2855_n 0.00885136f $X=3.325 $Y=1.91 $X2=0
+ $Y2=0
cc_522 N_SCD_c_574_n N_noxref_37_c_2855_n 0.00557949f $X=2.85 $Y=1.91 $X2=0
+ $Y2=0
cc_523 SCD N_noxref_37_c_2855_n 0.0131961f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_524 N_SCD_c_576_n N_noxref_37_c_2855_n 3.44981e-19 $X=3.49 $Y=1.8 $X2=0 $Y2=0
cc_525 N_SCD_c_572_n N_noxref_37_c_2857_n 0.00637046f $X=2.855 $Y=1.835 $X2=0
+ $Y2=0
cc_526 SCD N_noxref_37_c_2857_n 0.0183134f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_527 N_SCD_c_576_n N_noxref_37_c_2857_n 0.00126605f $X=3.49 $Y=1.8 $X2=0 $Y2=0
cc_528 N_SCD_c_572_n N_noxref_39_c_2888_n 0.00175545f $X=2.855 $Y=1.835 $X2=0
+ $Y2=0
cc_529 N_SCD_c_572_n N_noxref_39_c_2889_n 0.00900822f $X=2.855 $Y=1.835 $X2=0
+ $Y2=0
cc_530 N_SCD_c_573_n N_noxref_39_c_2889_n 0.00217117f $X=3.325 $Y=1.91 $X2=0
+ $Y2=0
cc_531 SCD N_noxref_39_c_2889_n 0.0139049f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_532 N_SCD_c_576_n N_noxref_39_c_2889_n 0.00174977f $X=3.49 $Y=1.8 $X2=0 $Y2=0
cc_533 SCD N_noxref_39_c_2892_n 0.00310926f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_534 N_A_876_93#_M1032_g N_A_967_193#_M1015_g 0.0395576f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_535 N_A_876_93#_c_613_n N_A_967_193#_M1015_g 5.20516e-19 $X=6.57 $Y=0.35
+ $X2=0 $Y2=0
cc_536 N_A_876_93#_M1032_g N_A_967_193#_c_792_n 0.0174614f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_537 N_A_876_93#_c_636_p N_A_967_193#_M1057_g 7.95427e-19 $X=8.505 $Y=0.645
+ $X2=0 $Y2=0
cc_538 N_A_876_93#_c_637_p N_A_967_193#_M1057_g 0.0127926f $X=9.765 $Y=0.73
+ $X2=0 $Y2=0
cc_539 N_A_876_93#_c_619_n N_A_967_193#_M1057_g 0.0014773f $X=9.93 $Y=0.43 $X2=0
+ $Y2=0
cc_540 N_A_876_93#_c_620_n N_A_967_193#_M1057_g 0.00108332f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_541 N_A_876_93#_c_629_n N_A_967_193#_M1029_g 0.00198615f $X=9.85 $Y=1.98
+ $X2=0 $Y2=0
cc_542 N_A_876_93#_c_637_p N_A_967_193#_M1010_g 0.0120631f $X=9.765 $Y=0.73
+ $X2=0 $Y2=0
cc_543 N_A_876_93#_c_619_n N_A_967_193#_M1010_g 0.00719413f $X=9.93 $Y=0.43
+ $X2=0 $Y2=0
cc_544 N_A_876_93#_c_620_n N_A_967_193#_M1010_g 0.0101796f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_545 N_A_876_93#_c_624_n N_A_967_193#_M1010_g 0.00154438f $X=9.93 $Y=0.73
+ $X2=0 $Y2=0
cc_546 N_A_876_93#_c_620_n N_A_967_193#_c_795_n 0.0109097f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_547 N_A_876_93#_c_621_n N_A_967_193#_c_795_n 0.00442471f $X=10.735 $Y=1.6
+ $X2=0 $Y2=0
cc_548 N_A_876_93#_c_625_n N_A_967_193#_c_795_n 0.00809844f $X=9.93 $Y=1.6 $X2=0
+ $Y2=0
cc_549 N_A_876_93#_c_620_n N_A_967_193#_c_796_n 0.00147809f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_550 N_A_876_93#_c_625_n N_A_967_193#_c_796_n 0.00440039f $X=9.93 $Y=1.6 $X2=0
+ $Y2=0
cc_551 N_A_876_93#_M1051_g N_A_967_193#_c_797_n 0.0127307f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_552 N_A_876_93#_c_619_n N_A_967_193#_c_797_n 0.00960805f $X=9.93 $Y=0.43
+ $X2=0 $Y2=0
cc_553 N_A_876_93#_c_620_n N_A_967_193#_c_797_n 0.00834488f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_554 N_A_876_93#_c_624_n N_A_967_193#_c_797_n 0.00253712f $X=9.93 $Y=0.73
+ $X2=0 $Y2=0
cc_555 N_A_876_93#_M1044_g N_A_967_193#_c_798_n 0.0272112f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_556 N_A_876_93#_c_629_n N_A_967_193#_c_798_n 0.00604003f $X=9.85 $Y=1.98
+ $X2=0 $Y2=0
cc_557 N_A_876_93#_c_621_n N_A_967_193#_c_798_n 0.0128584f $X=10.735 $Y=1.6
+ $X2=0 $Y2=0
cc_558 N_A_876_93#_M1051_g N_A_967_193#_c_799_n 0.0102957f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_559 N_A_876_93#_M1044_g N_A_967_193#_c_825_n 0.00830878f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_560 N_A_876_93#_M1044_g N_A_967_193#_M1042_g 0.0218299f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_561 N_A_876_93#_M1051_g N_A_967_193#_M1045_g 0.0181172f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_562 N_A_876_93#_c_621_n N_A_967_193#_c_805_n 0.00861195f $X=10.735 $Y=1.6
+ $X2=0 $Y2=0
cc_563 N_A_876_93#_c_626_n N_A_967_193#_c_805_n 0.0194852f $X=10.765 $Y=1.59
+ $X2=0 $Y2=0
cc_564 N_A_876_93#_c_613_n N_A_1147_490#_c_1092_n 0.00164789f $X=6.57 $Y=0.35
+ $X2=0 $Y2=0
cc_565 N_A_876_93#_c_615_n N_A_1147_490#_c_1092_n 0.0644084f $X=7.5 $Y=0.8 $X2=0
+ $Y2=0
cc_566 N_A_876_93#_c_665_p N_A_1147_490#_c_1092_n 0.0115167f $X=6.74 $Y=0.8
+ $X2=0 $Y2=0
cc_567 N_A_876_93#_c_617_n N_A_1147_490#_c_1092_n 0.00542747f $X=8.42 $Y=0.35
+ $X2=0 $Y2=0
cc_568 N_A_876_93#_c_617_n N_A_1147_490#_c_1094_n 0.00439765f $X=8.42 $Y=0.35
+ $X2=0 $Y2=0
cc_569 N_A_876_93#_c_637_p N_A_1147_490#_c_1094_n 0.0569981f $X=9.765 $Y=0.73
+ $X2=0 $Y2=0
cc_570 N_A_876_93#_c_669_p N_A_1147_490#_c_1094_n 0.00842615f $X=8.59 $Y=0.73
+ $X2=0 $Y2=0
cc_571 N_A_876_93#_c_620_n N_A_1147_490#_c_1094_n 0.0101043f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_572 N_A_876_93#_c_620_n N_A_1147_490#_c_1095_n 0.0189871f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_573 N_A_876_93#_c_629_n N_A_1147_490#_c_1095_n 0.0352733f $X=9.85 $Y=1.98
+ $X2=0 $Y2=0
cc_574 N_A_876_93#_c_625_n N_A_1147_490#_c_1095_n 0.0251978f $X=9.93 $Y=1.6
+ $X2=0 $Y2=0
cc_575 N_A_876_93#_M1029_d N_A_1147_490#_c_1109_n 0.00595816f $X=9.71 $Y=1.835
+ $X2=0 $Y2=0
cc_576 N_A_876_93#_c_629_n N_A_1147_490#_c_1109_n 0.0115129f $X=9.85 $Y=1.98
+ $X2=0 $Y2=0
cc_577 N_A_876_93#_M1044_g N_A_1147_490#_c_1110_n 0.00117311f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_578 N_A_876_93#_c_629_n N_A_1147_490#_c_1110_n 0.0418163f $X=9.85 $Y=1.98
+ $X2=0 $Y2=0
cc_579 N_A_876_93#_M1044_g N_A_1147_490#_c_1111_n 0.0117459f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_580 N_A_876_93#_c_621_n N_A_1147_490#_c_1111_n 0.0430269f $X=10.735 $Y=1.6
+ $X2=0 $Y2=0
cc_581 N_A_876_93#_c_626_n N_A_1147_490#_c_1111_n 0.009413f $X=10.765 $Y=1.59
+ $X2=0 $Y2=0
cc_582 N_A_876_93#_c_629_n N_A_1147_490#_c_1112_n 0.0135568f $X=9.85 $Y=1.98
+ $X2=0 $Y2=0
cc_583 N_A_876_93#_c_621_n N_A_1147_490#_c_1112_n 0.0131219f $X=10.735 $Y=1.6
+ $X2=0 $Y2=0
cc_584 N_A_876_93#_M1051_g N_A_1147_490#_c_1096_n 0.00448139f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_585 N_A_876_93#_c_619_n N_A_1147_490#_c_1096_n 0.00262944f $X=9.93 $Y=0.43
+ $X2=0 $Y2=0
cc_586 N_A_876_93#_c_620_n N_A_1147_490#_c_1096_n 0.010196f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_587 N_A_876_93#_c_624_n N_A_1147_490#_c_1096_n 0.00681237f $X=9.93 $Y=0.73
+ $X2=0 $Y2=0
cc_588 N_A_876_93#_M1044_g N_A_1147_490#_c_1097_n 0.00344273f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_589 N_A_876_93#_M1051_g N_A_1147_490#_c_1097_n 0.00985831f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_590 N_A_876_93#_c_621_n N_A_1147_490#_c_1097_n 0.0246103f $X=10.735 $Y=1.6
+ $X2=0 $Y2=0
cc_591 N_A_876_93#_c_626_n N_A_1147_490#_c_1097_n 0.00923468f $X=10.765 $Y=1.59
+ $X2=0 $Y2=0
cc_592 N_A_876_93#_c_613_n N_A_1147_490#_c_1098_n 0.00339737f $X=6.57 $Y=0.35
+ $X2=0 $Y2=0
cc_593 N_A_876_93#_c_615_n N_A_1147_490#_c_1100_n 0.0146155f $X=7.5 $Y=0.8 $X2=0
+ $Y2=0
cc_594 N_A_876_93#_c_616_n N_A_1147_490#_c_1100_n 0.00768154f $X=7.585 $Y=0.715
+ $X2=0 $Y2=0
cc_595 N_A_876_93#_c_617_n N_A_1147_490#_c_1100_n 0.0259929f $X=8.42 $Y=0.35
+ $X2=0 $Y2=0
cc_596 N_A_876_93#_c_636_p N_A_1147_490#_c_1100_n 0.00211237f $X=8.505 $Y=0.645
+ $X2=0 $Y2=0
cc_597 N_A_876_93#_c_669_p N_A_1147_490#_c_1100_n 0.0135888f $X=8.59 $Y=0.73
+ $X2=0 $Y2=0
cc_598 N_A_876_93#_M1051_g N_A_1147_490#_c_1101_n 0.0157314f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_599 N_A_876_93#_c_620_n N_A_1147_490#_c_1101_n 0.00669386f $X=9.93 $Y=1.435
+ $X2=0 $Y2=0
cc_600 N_A_876_93#_c_621_n N_A_1147_490#_c_1101_n 0.0201562f $X=10.735 $Y=1.6
+ $X2=0 $Y2=0
cc_601 N_A_876_93#_c_626_n N_A_1147_490#_c_1101_n 0.0106529f $X=10.765 $Y=1.59
+ $X2=0 $Y2=0
cc_602 N_A_876_93#_M1044_g N_A_1147_490#_c_1114_n 0.00135051f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_603 N_A_876_93#_c_613_n N_A_1147_490#_c_1102_n 0.00196586f $X=6.57 $Y=0.35
+ $X2=0 $Y2=0
cc_604 N_A_876_93#_c_614_n N_A_1147_490#_c_1102_n 0.00345307f $X=6.655 $Y=0.715
+ $X2=0 $Y2=0
cc_605 N_A_876_93#_M1032_g N_RESET_B_M1041_g 5.52563e-19 $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_606 N_A_876_93#_c_622_n N_RESET_B_M1041_g 5.2369e-19 $X=4.545 $Y=0.35 $X2=0
+ $Y2=0
cc_607 N_A_876_93#_c_623_n N_RESET_B_M1041_g 0.00428363f $X=4.545 $Y=0.63 $X2=0
+ $Y2=0
cc_608 N_A_876_93#_c_613_n N_RESET_B_c_1288_n 0.041722f $X=6.57 $Y=0.35 $X2=0
+ $Y2=0
cc_609 N_A_876_93#_c_622_n N_RESET_B_c_1288_n 0.00249662f $X=4.545 $Y=0.35 $X2=0
+ $Y2=0
cc_610 N_A_876_93#_c_623_n N_RESET_B_c_1288_n 0.0193123f $X=4.545 $Y=0.63 $X2=0
+ $Y2=0
cc_611 N_A_876_93#_M1032_g N_RESET_B_c_1302_n 0.0162052f $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_612 N_A_876_93#_c_613_n N_RESET_B_M1005_g 0.00443749f $X=6.57 $Y=0.35 $X2=0
+ $Y2=0
cc_613 N_A_876_93#_c_614_n N_RESET_B_M1005_g 0.003242f $X=6.655 $Y=0.715 $X2=0
+ $Y2=0
cc_614 N_A_876_93#_c_615_n N_RESET_B_M1005_g 0.0135141f $X=7.5 $Y=0.8 $X2=0
+ $Y2=0
cc_615 N_A_876_93#_c_616_n N_RESET_B_M1005_g 0.0040992f $X=7.585 $Y=0.715 $X2=0
+ $Y2=0
cc_616 N_A_876_93#_M1032_g N_RESET_B_c_1292_n 0.0167373f $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_617 N_A_876_93#_M1032_g N_RESET_B_c_1311_n 0.00165392f $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_618 N_A_876_93#_M1029_d N_RESET_B_c_1313_n 0.00403646f $X=9.71 $Y=1.835 $X2=0
+ $Y2=0
cc_619 N_A_876_93#_M1044_g N_RESET_B_c_1313_n 0.00378765f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_620 N_A_876_93#_c_629_n N_RESET_B_c_1313_n 0.0170987f $X=9.85 $Y=1.98 $X2=0
+ $Y2=0
cc_621 N_A_876_93#_c_621_n N_RESET_B_c_1313_n 0.00158216f $X=10.735 $Y=1.6 $X2=0
+ $Y2=0
cc_622 N_A_876_93#_c_625_n N_RESET_B_c_1313_n 0.00577392f $X=9.93 $Y=1.6 $X2=0
+ $Y2=0
cc_623 N_A_876_93#_M1032_g N_RESET_B_c_1297_n 0.0462143f $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_624 N_A_876_93#_M1032_g N_RESET_B_c_1298_n 0.00356364f $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_625 N_A_876_93#_c_616_n N_A_911_219#_M1000_g 0.00464978f $X=7.585 $Y=0.715
+ $X2=0 $Y2=0
cc_626 N_A_876_93#_c_617_n N_A_911_219#_M1000_g 0.0113089f $X=8.42 $Y=0.35 $X2=0
+ $Y2=0
cc_627 N_A_876_93#_c_636_p N_A_911_219#_M1000_g 0.00405082f $X=8.505 $Y=0.645
+ $X2=0 $Y2=0
cc_628 N_A_876_93#_c_669_p N_A_911_219#_M1000_g 0.00116289f $X=8.59 $Y=0.73
+ $X2=0 $Y2=0
cc_629 N_A_876_93#_c_617_n N_A_911_219#_M1021_g 0.00389352f $X=8.42 $Y=0.35
+ $X2=0 $Y2=0
cc_630 N_A_876_93#_c_636_p N_A_911_219#_M1021_g 0.00564384f $X=8.505 $Y=0.645
+ $X2=0 $Y2=0
cc_631 N_A_876_93#_c_637_p N_A_911_219#_M1021_g 0.00842229f $X=9.765 $Y=0.73
+ $X2=0 $Y2=0
cc_632 N_A_876_93#_c_669_p N_A_911_219#_M1021_g 0.00237414f $X=8.59 $Y=0.73
+ $X2=0 $Y2=0
cc_633 N_A_876_93#_M1032_g N_A_911_219#_c_1560_n 0.00233985f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_634 N_A_876_93#_M1032_g N_A_911_219#_c_1562_n 0.00114045f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_635 N_A_876_93#_M1032_g N_A_911_219#_c_1555_n 0.00516707f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_636 N_A_876_93#_M1051_g N_A_2168_439#_c_1855_n 0.00454537f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_637 N_A_876_93#_M1051_g N_A_2168_439#_c_1856_n 0.00140967f $X=11.08 $Y=0.915
+ $X2=0 $Y2=0
cc_638 N_A_876_93#_M1044_g N_A_2168_439#_c_1879_n 0.00261241f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_639 N_A_876_93#_M1032_g N_VPWR_c_2206_n 0.00378843f $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_640 N_A_876_93#_M1029_d N_VPWR_c_2191_n 0.00233022f $X=9.71 $Y=1.835 $X2=0
+ $Y2=0
cc_641 N_A_876_93#_M1032_g N_VPWR_c_2191_n 0.00519032f $X=4.48 $Y=1.305 $X2=0
+ $Y2=0
cc_642 N_A_876_93#_M1032_g N_A_342_261#_c_2422_n 0.0107319f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_643 N_A_876_93#_M1032_g N_A_342_261#_c_2413_n 0.0126909f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_644 N_A_876_93#_M1032_g N_A_342_261#_c_2414_n 0.00245967f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_645 N_A_876_93#_M1032_g N_A_342_261#_c_2415_n 0.00948659f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_646 N_A_876_93#_M1044_g N_A_2081_439#_c_2552_n 0.0084067f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_647 N_A_876_93#_M1044_g N_A_2081_439#_c_2555_n 0.00273774f $X=10.765 $Y=2.405
+ $X2=0 $Y2=0
cc_648 N_A_876_93#_c_615_n N_VGND_M1005_d 0.010182f $X=7.5 $Y=0.8 $X2=0 $Y2=0
cc_649 N_A_876_93#_c_637_p N_VGND_M1021_d 0.0117478f $X=9.765 $Y=0.73 $X2=0
+ $Y2=0
cc_650 N_A_876_93#_c_613_n N_VGND_c_2683_n 0.011083f $X=6.57 $Y=0.35 $X2=0 $Y2=0
cc_651 N_A_876_93#_c_614_n N_VGND_c_2683_n 0.00581049f $X=6.655 $Y=0.715 $X2=0
+ $Y2=0
cc_652 N_A_876_93#_c_615_n N_VGND_c_2683_n 0.0184457f $X=7.5 $Y=0.8 $X2=0 $Y2=0
cc_653 N_A_876_93#_c_616_n N_VGND_c_2683_n 0.0056646f $X=7.585 $Y=0.715 $X2=0
+ $Y2=0
cc_654 N_A_876_93#_c_618_n N_VGND_c_2683_n 0.0108372f $X=7.67 $Y=0.35 $X2=0
+ $Y2=0
cc_655 N_A_876_93#_c_617_n N_VGND_c_2684_n 0.0101302f $X=8.42 $Y=0.35 $X2=0
+ $Y2=0
cc_656 N_A_876_93#_c_636_p N_VGND_c_2684_n 0.00151347f $X=8.505 $Y=0.645 $X2=0
+ $Y2=0
cc_657 N_A_876_93#_c_637_p N_VGND_c_2684_n 0.0237698f $X=9.765 $Y=0.73 $X2=0
+ $Y2=0
cc_658 N_A_876_93#_c_613_n N_VGND_c_2688_n 0.12409f $X=6.57 $Y=0.35 $X2=0 $Y2=0
cc_659 N_A_876_93#_c_615_n N_VGND_c_2688_n 0.00309923f $X=7.5 $Y=0.8 $X2=0 $Y2=0
cc_660 N_A_876_93#_c_622_n N_VGND_c_2688_n 0.0214369f $X=4.545 $Y=0.35 $X2=0
+ $Y2=0
cc_661 N_A_876_93#_c_615_n N_VGND_c_2694_n 0.00389189f $X=7.5 $Y=0.8 $X2=0 $Y2=0
cc_662 N_A_876_93#_c_617_n N_VGND_c_2694_n 0.0567024f $X=8.42 $Y=0.35 $X2=0
+ $Y2=0
cc_663 N_A_876_93#_c_618_n N_VGND_c_2694_n 0.0113826f $X=7.67 $Y=0.35 $X2=0
+ $Y2=0
cc_664 N_A_876_93#_c_637_p N_VGND_c_2694_n 0.00413351f $X=9.765 $Y=0.73 $X2=0
+ $Y2=0
cc_665 N_A_876_93#_c_637_p N_VGND_c_2695_n 0.00813591f $X=9.765 $Y=0.73 $X2=0
+ $Y2=0
cc_666 N_A_876_93#_c_619_n N_VGND_c_2695_n 0.019758f $X=9.93 $Y=0.43 $X2=0 $Y2=0
cc_667 N_A_876_93#_M1010_d N_VGND_c_2698_n 0.00229659f $X=9.79 $Y=0.235 $X2=0
+ $Y2=0
cc_668 N_A_876_93#_M1051_g N_VGND_c_2698_n 9.39239e-19 $X=11.08 $Y=0.915 $X2=0
+ $Y2=0
cc_669 N_A_876_93#_c_613_n N_VGND_c_2698_n 0.0679736f $X=6.57 $Y=0.35 $X2=0
+ $Y2=0
cc_670 N_A_876_93#_c_615_n N_VGND_c_2698_n 0.0139256f $X=7.5 $Y=0.8 $X2=0 $Y2=0
cc_671 N_A_876_93#_c_617_n N_VGND_c_2698_n 0.0345619f $X=8.42 $Y=0.35 $X2=0
+ $Y2=0
cc_672 N_A_876_93#_c_618_n N_VGND_c_2698_n 0.00656134f $X=7.67 $Y=0.35 $X2=0
+ $Y2=0
cc_673 N_A_876_93#_c_637_p N_VGND_c_2698_n 0.0239728f $X=9.765 $Y=0.73 $X2=0
+ $Y2=0
cc_674 N_A_876_93#_c_619_n N_VGND_c_2698_n 0.012508f $X=9.93 $Y=0.43 $X2=0 $Y2=0
cc_675 N_A_876_93#_c_622_n N_VGND_c_2698_n 0.0112452f $X=4.545 $Y=0.35 $X2=0
+ $Y2=0
cc_676 N_A_876_93#_M1032_g N_noxref_39_c_2894_n 9.89873e-19 $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_677 N_A_876_93#_c_622_n N_noxref_39_c_2894_n 0.0370171f $X=4.545 $Y=0.35
+ $X2=0 $Y2=0
cc_678 N_A_876_93#_c_623_n N_noxref_39_c_2894_n 0.00398163f $X=4.545 $Y=0.63
+ $X2=0 $Y2=0
cc_679 N_A_876_93#_M1032_g N_A_824_219#_c_2941_n 0.0150947f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_680 N_A_876_93#_c_613_n N_A_824_219#_c_2941_n 0.0292037f $X=6.57 $Y=0.35
+ $X2=0 $Y2=0
cc_681 N_A_876_93#_c_622_n N_A_824_219#_c_2941_n 0.0248086f $X=4.545 $Y=0.35
+ $X2=0 $Y2=0
cc_682 N_A_876_93#_c_623_n N_A_824_219#_c_2941_n 0.00446668f $X=4.545 $Y=0.63
+ $X2=0 $Y2=0
cc_683 N_A_876_93#_c_613_n N_A_824_219#_c_2942_n 0.0279535f $X=6.57 $Y=0.35
+ $X2=0 $Y2=0
cc_684 N_A_876_93#_M1032_g N_A_824_219#_c_2943_n 0.00102833f $X=4.48 $Y=1.305
+ $X2=0 $Y2=0
cc_685 N_A_876_93#_c_613_n N_A_824_219#_c_2944_n 0.0149241f $X=6.57 $Y=0.35
+ $X2=0 $Y2=0
cc_686 N_A_876_93#_c_665_p A_1303_119# 0.00145611f $X=6.74 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_687 N_A_876_93#_c_636_p A_1661_87# 0.00225487f $X=8.505 $Y=0.645 $X2=-0.19
+ $Y2=-0.245
cc_688 N_A_876_93#_c_669_p A_1661_87# 0.00221959f $X=8.59 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_689 N_A_876_93#_c_637_p A_1880_47# 0.00352317f $X=9.765 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_690 N_A_967_193#_c_828_n N_A_1147_490#_c_1104_n 0.00114316f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_691 N_A_967_193#_c_836_n N_A_1147_490#_c_1104_n 0.0129874f $X=5.99 $Y=2.05
+ $X2=0 $Y2=0
cc_692 N_A_967_193#_M1028_g N_A_1147_490#_c_1105_n 0.0121603f $X=5.025 $Y=2.665
+ $X2=0 $Y2=0
cc_693 N_A_967_193#_c_791_n N_A_1147_490#_c_1105_n 0.0129874f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_694 N_A_967_193#_c_835_n N_A_1147_490#_c_1105_n 3.15928e-19 $X=6.005 $Y=1.97
+ $X2=0 $Y2=0
cc_695 N_A_967_193#_c_828_n N_A_1147_490#_c_1091_n 0.0104313f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_696 N_A_967_193#_c_835_n N_A_1147_490#_c_1091_n 0.00118353f $X=6.005 $Y=1.97
+ $X2=0 $Y2=0
cc_697 N_A_967_193#_c_836_n N_A_1147_490#_c_1091_n 0.023793f $X=5.99 $Y=2.05
+ $X2=0 $Y2=0
cc_698 N_A_967_193#_c_828_n N_A_1147_490#_c_1093_n 0.0139102f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_699 N_A_967_193#_c_829_n N_A_1147_490#_c_1093_n 0.0471828f $X=7.725 $Y=2.895
+ $X2=0 $Y2=0
cc_700 N_A_967_193#_c_830_n N_A_1147_490#_c_1093_n 0.015156f $X=8.42 $Y=2.98
+ $X2=0 $Y2=0
cc_701 N_A_967_193#_c_832_n N_A_1147_490#_c_1093_n 0.0446769f $X=8.505 $Y=2.895
+ $X2=0 $Y2=0
cc_702 N_A_967_193#_c_808_n N_A_1147_490#_c_1093_n 0.0254083f $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_703 N_A_967_193#_M1057_g N_A_1147_490#_c_1094_n 0.0154637f $X=9.325 $Y=0.655
+ $X2=0 $Y2=0
cc_704 N_A_967_193#_M1010_g N_A_1147_490#_c_1094_n 9.87159e-19 $X=9.715 $Y=0.655
+ $X2=0 $Y2=0
cc_705 N_A_967_193#_c_796_n N_A_1147_490#_c_1094_n 0.00743529f $X=9.79 $Y=1.42
+ $X2=0 $Y2=0
cc_706 N_A_967_193#_c_808_n N_A_1147_490#_c_1094_n 0.0134111f $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_707 N_A_967_193#_c_809_n N_A_1147_490#_c_1094_n 0.0469999f $X=9.1 $Y=1.51
+ $X2=0 $Y2=0
cc_708 N_A_967_193#_M1025_g N_A_1147_490#_c_1095_n 0.0103798f $X=9.275 $Y=2.465
+ $X2=0 $Y2=0
cc_709 N_A_967_193#_M1057_g N_A_1147_490#_c_1095_n 0.00439211f $X=9.325 $Y=0.655
+ $X2=0 $Y2=0
cc_710 N_A_967_193#_M1029_g N_A_1147_490#_c_1095_n 0.0206121f $X=9.635 $Y=2.465
+ $X2=0 $Y2=0
cc_711 N_A_967_193#_M1010_g N_A_1147_490#_c_1095_n 0.00118084f $X=9.715 $Y=0.655
+ $X2=0 $Y2=0
cc_712 N_A_967_193#_c_796_n N_A_1147_490#_c_1095_n 0.0153686f $X=9.79 $Y=1.42
+ $X2=0 $Y2=0
cc_713 N_A_967_193#_c_798_n N_A_1147_490#_c_1095_n 5.60842e-19 $X=10.255
+ $Y=2.985 $X2=0 $Y2=0
cc_714 N_A_967_193#_c_809_n N_A_1147_490#_c_1095_n 0.0238596f $X=9.1 $Y=1.51
+ $X2=0 $Y2=0
cc_715 N_A_967_193#_M1029_g N_A_1147_490#_c_1109_n 0.00854145f $X=9.635 $Y=2.465
+ $X2=0 $Y2=0
cc_716 N_A_967_193#_c_798_n N_A_1147_490#_c_1109_n 0.00375393f $X=10.255
+ $Y=2.985 $X2=0 $Y2=0
cc_717 N_A_967_193#_c_826_n N_A_1147_490#_c_1109_n 0.00408698f $X=10.33 $Y=3.06
+ $X2=0 $Y2=0
cc_718 N_A_967_193#_M1025_g N_A_1147_490#_c_1184_n 0.00125403f $X=9.275 $Y=2.465
+ $X2=0 $Y2=0
cc_719 N_A_967_193#_M1029_g N_A_1147_490#_c_1184_n 0.00155755f $X=9.635 $Y=2.465
+ $X2=0 $Y2=0
cc_720 N_A_967_193#_M1029_g N_A_1147_490#_c_1110_n 0.00203204f $X=9.635 $Y=2.465
+ $X2=0 $Y2=0
cc_721 N_A_967_193#_c_798_n N_A_1147_490#_c_1110_n 0.0201468f $X=10.255 $Y=2.985
+ $X2=0 $Y2=0
cc_722 N_A_967_193#_c_798_n N_A_1147_490#_c_1111_n 0.00442675f $X=10.255
+ $Y=2.985 $X2=0 $Y2=0
cc_723 N_A_967_193#_c_798_n N_A_1147_490#_c_1112_n 0.00473587f $X=10.255
+ $Y=2.985 $X2=0 $Y2=0
cc_724 N_A_967_193#_c_797_n N_A_1147_490#_c_1096_n 0.00567348f $X=10.255
+ $Y=1.345 $X2=0 $Y2=0
cc_725 N_A_967_193#_c_799_n N_A_1147_490#_c_1096_n 0.0065164f $X=11.55 $Y=0.18
+ $X2=0 $Y2=0
cc_726 N_A_967_193#_M1042_g N_A_1147_490#_c_1097_n 0.0034796f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_727 N_A_967_193#_c_797_n N_A_1147_490#_c_1101_n 0.00201979f $X=10.255
+ $Y=1.345 $X2=0 $Y2=0
cc_728 N_A_967_193#_M1045_g N_A_1147_490#_c_1101_n 0.00167593f $X=11.625
+ $Y=0.915 $X2=0 $Y2=0
cc_729 N_A_967_193#_M1042_g N_A_1147_490#_c_1114_n 0.0164492f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_730 N_A_967_193#_M1045_g N_A_1147_490#_c_1114_n 0.00160833f $X=11.625
+ $Y=0.915 $X2=0 $Y2=0
cc_731 N_A_967_193#_M1015_g N_RESET_B_c_1288_n 0.00129703f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_732 N_A_967_193#_c_828_n N_RESET_B_M1005_g 0.0121631f $X=7.64 $Y=1.97 $X2=0
+ $Y2=0
cc_733 N_A_967_193#_c_803_n N_RESET_B_M1054_g 0.00495156f $X=14.5 $Y=0.18 $X2=0
+ $Y2=0
cc_734 N_A_967_193#_c_812_n N_RESET_B_M1054_g 0.00111755f $X=12.855 $Y=0.43
+ $X2=0 $Y2=0
cc_735 N_A_967_193#_c_814_n N_RESET_B_M1054_g 0.00168671f $X=14.5 $Y=0.487 $X2=0
+ $Y2=0
cc_736 N_A_967_193#_M1028_g N_RESET_B_c_1311_n 0.00241705f $X=5.025 $Y=2.665
+ $X2=0 $Y2=0
cc_737 N_A_967_193#_c_791_n N_RESET_B_c_1311_n 0.0163362f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_738 N_A_967_193#_c_792_n N_RESET_B_c_1311_n 0.00326086f $X=5.1 $Y=2.142 $X2=0
+ $Y2=0
cc_739 N_A_967_193#_c_828_n N_RESET_B_c_1311_n 0.0149852f $X=7.64 $Y=1.97 $X2=0
+ $Y2=0
cc_740 N_A_967_193#_c_835_n N_RESET_B_c_1311_n 0.00793652f $X=6.005 $Y=1.97
+ $X2=0 $Y2=0
cc_741 N_A_967_193#_M1025_g N_RESET_B_c_1313_n 0.0110001f $X=9.275 $Y=2.465
+ $X2=0 $Y2=0
cc_742 N_A_967_193#_M1029_g N_RESET_B_c_1313_n 0.00686428f $X=9.635 $Y=2.465
+ $X2=0 $Y2=0
cc_743 N_A_967_193#_c_798_n N_RESET_B_c_1313_n 0.00339426f $X=10.255 $Y=2.985
+ $X2=0 $Y2=0
cc_744 N_A_967_193#_c_825_n N_RESET_B_c_1313_n 7.93409e-19 $X=11.235 $Y=3.06
+ $X2=0 $Y2=0
cc_745 N_A_967_193#_M1042_g N_RESET_B_c_1313_n 0.00302943f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_746 N_A_967_193#_c_828_n N_RESET_B_c_1313_n 0.016659f $X=7.64 $Y=1.97 $X2=0
+ $Y2=0
cc_747 N_A_967_193#_c_829_n N_RESET_B_c_1313_n 0.0197545f $X=7.725 $Y=2.895
+ $X2=0 $Y2=0
cc_748 N_A_967_193#_c_830_n N_RESET_B_c_1313_n 0.0135422f $X=8.42 $Y=2.98 $X2=0
+ $Y2=0
cc_749 N_A_967_193#_c_832_n N_RESET_B_c_1313_n 0.0241844f $X=8.505 $Y=2.895
+ $X2=0 $Y2=0
cc_750 N_A_967_193#_c_828_n N_RESET_B_c_1314_n 0.00225868f $X=7.64 $Y=1.97 $X2=0
+ $Y2=0
cc_751 N_A_967_193#_c_829_n N_RESET_B_c_1314_n 0.0016978f $X=7.725 $Y=2.895
+ $X2=0 $Y2=0
cc_752 N_A_967_193#_c_828_n N_RESET_B_c_1318_n 0.0103071f $X=7.64 $Y=1.97 $X2=0
+ $Y2=0
cc_753 N_A_967_193#_c_829_n N_RESET_B_c_1318_n 0.0109272f $X=7.725 $Y=2.895
+ $X2=0 $Y2=0
cc_754 N_A_967_193#_c_828_n N_RESET_B_c_1319_n 0.0221256f $X=7.64 $Y=1.97 $X2=0
+ $Y2=0
cc_755 N_A_967_193#_c_829_n N_RESET_B_c_1319_n 0.00568187f $X=7.725 $Y=2.895
+ $X2=0 $Y2=0
cc_756 N_A_967_193#_c_808_n N_A_911_219#_M1000_g 2.70371e-19 $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_757 N_A_967_193#_c_829_n N_A_911_219#_M1002_g 0.00356685f $X=7.725 $Y=2.895
+ $X2=0 $Y2=0
cc_758 N_A_967_193#_c_830_n N_A_911_219#_M1002_g 0.00669315f $X=8.42 $Y=2.98
+ $X2=0 $Y2=0
cc_759 N_A_967_193#_c_832_n N_A_911_219#_M1002_g 0.00555672f $X=8.505 $Y=2.895
+ $X2=0 $Y2=0
cc_760 N_A_967_193#_c_808_n N_A_911_219#_M1002_g 0.00102254f $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_761 N_A_967_193#_c_808_n N_A_911_219#_c_1546_n 0.00526248f $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_762 N_A_967_193#_M1057_g N_A_911_219#_M1021_g 0.0212194f $X=9.325 $Y=0.655
+ $X2=0 $Y2=0
cc_763 N_A_967_193#_c_796_n N_A_911_219#_M1021_g 0.00218407f $X=9.79 $Y=1.42
+ $X2=0 $Y2=0
cc_764 N_A_967_193#_c_808_n N_A_911_219#_M1021_g 0.00106386f $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_765 N_A_967_193#_c_809_n N_A_911_219#_M1021_g 0.00226808f $X=9.1 $Y=1.51
+ $X2=0 $Y2=0
cc_766 N_A_967_193#_M1025_g N_A_911_219#_M1009_g 0.0141759f $X=9.275 $Y=2.465
+ $X2=0 $Y2=0
cc_767 N_A_967_193#_c_832_n N_A_911_219#_M1009_g 0.0226862f $X=8.505 $Y=2.895
+ $X2=0 $Y2=0
cc_768 N_A_967_193#_c_808_n N_A_911_219#_M1009_g 9.99418e-19 $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_769 N_A_967_193#_c_809_n N_A_911_219#_M1009_g 0.00937645f $X=9.1 $Y=1.51
+ $X2=0 $Y2=0
cc_770 N_A_967_193#_c_796_n N_A_911_219#_c_1550_n 0.0188731f $X=9.79 $Y=1.42
+ $X2=0 $Y2=0
cc_771 N_A_967_193#_c_808_n N_A_911_219#_c_1550_n 6.3561e-19 $X=8.59 $Y=1.51
+ $X2=0 $Y2=0
cc_772 N_A_967_193#_c_809_n N_A_911_219#_c_1550_n 0.00371192f $X=9.1 $Y=1.51
+ $X2=0 $Y2=0
cc_773 N_A_967_193#_M1028_g N_A_911_219#_c_1560_n 5.89459e-19 $X=5.025 $Y=2.665
+ $X2=0 $Y2=0
cc_774 N_A_967_193#_M1015_g N_A_911_219#_c_1551_n 0.0111421f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_775 N_A_967_193#_c_791_n N_A_911_219#_c_1551_n 0.00389581f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_776 N_A_967_193#_c_792_n N_A_911_219#_c_1551_n 9.95394e-19 $X=5.1 $Y=2.142
+ $X2=0 $Y2=0
cc_777 N_A_967_193#_M1028_g N_A_911_219#_c_1561_n 0.0113089f $X=5.025 $Y=2.665
+ $X2=0 $Y2=0
cc_778 N_A_967_193#_c_791_n N_A_911_219#_c_1561_n 0.0104566f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_779 N_A_967_193#_c_792_n N_A_911_219#_c_1561_n 0.00114407f $X=5.1 $Y=2.142
+ $X2=0 $Y2=0
cc_780 N_A_967_193#_c_792_n N_A_911_219#_c_1562_n 0.00180261f $X=5.1 $Y=2.142
+ $X2=0 $Y2=0
cc_781 N_A_967_193#_M1015_g N_A_911_219#_c_1552_n 0.0022453f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_782 N_A_967_193#_M1015_g N_A_911_219#_c_1553_n 4.52138e-19 $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_783 N_A_967_193#_M1028_g N_A_911_219#_c_1553_n 0.00340983f $X=5.025 $Y=2.665
+ $X2=0 $Y2=0
cc_784 N_A_967_193#_c_791_n N_A_911_219#_c_1553_n 0.0174409f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_785 N_A_967_193#_c_835_n N_A_911_219#_c_1553_n 0.0229425f $X=6.005 $Y=1.97
+ $X2=0 $Y2=0
cc_786 N_A_967_193#_c_836_n N_A_911_219#_c_1553_n 0.00369219f $X=5.99 $Y=2.05
+ $X2=0 $Y2=0
cc_787 N_A_967_193#_c_791_n N_A_911_219#_c_1554_n 0.00305321f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_788 N_A_967_193#_c_828_n N_A_911_219#_c_1554_n 0.0969495f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_789 N_A_967_193#_c_835_n N_A_911_219#_c_1554_n 0.0225071f $X=6.005 $Y=1.97
+ $X2=0 $Y2=0
cc_790 N_A_967_193#_c_836_n N_A_911_219#_c_1554_n 0.00295632f $X=5.99 $Y=2.05
+ $X2=0 $Y2=0
cc_791 N_A_967_193#_c_791_n N_A_911_219#_c_1565_n 0.00407408f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_792 N_A_967_193#_c_828_n N_A_911_219#_c_1565_n 0.0119853f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_793 N_A_967_193#_c_835_n N_A_911_219#_c_1565_n 0.0195166f $X=6.005 $Y=1.97
+ $X2=0 $Y2=0
cc_794 N_A_967_193#_c_828_n N_A_911_219#_c_1619_n 0.0033119f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_795 N_A_967_193#_M1015_g N_A_911_219#_c_1555_n 0.00439537f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_796 N_A_967_193#_M1015_g N_A_911_219#_c_1556_n 0.00135954f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_797 N_A_967_193#_c_828_n N_A_911_219#_c_1622_n 0.00253475f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_798 N_A_967_193#_c_829_n N_A_911_219#_c_1622_n 0.0142061f $X=7.725 $Y=2.895
+ $X2=0 $Y2=0
cc_799 N_A_967_193#_c_831_n N_A_911_219#_c_1622_n 0.0139102f $X=7.81 $Y=2.98
+ $X2=0 $Y2=0
cc_800 N_A_967_193#_c_828_n N_A_911_219#_c_1568_n 0.0255743f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_801 N_A_967_193#_c_828_n N_A_911_219#_c_1557_n 0.00245628f $X=7.64 $Y=1.97
+ $X2=0 $Y2=0
cc_802 N_A_967_193#_M1045_g N_A_2388_115#_c_1729_n 0.0351778f $X=11.625 $Y=0.915
+ $X2=0 $Y2=0
cc_803 N_A_967_193#_c_802_n N_A_2388_115#_c_1729_n 0.00654454f $X=12.69 $Y=0.18
+ $X2=0 $Y2=0
cc_804 N_A_967_193#_c_812_n N_A_2388_115#_c_1729_n 2.3257e-19 $X=12.855 $Y=0.43
+ $X2=0 $Y2=0
cc_805 N_A_967_193#_c_811_n N_A_2388_115#_c_1746_n 0.00771307f $X=12.855 $Y=0.35
+ $X2=0 $Y2=0
cc_806 N_A_967_193#_c_812_n N_A_2388_115#_c_1746_n 9.92375e-19 $X=12.855 $Y=0.43
+ $X2=0 $Y2=0
cc_807 N_A_967_193#_c_814_n N_A_2388_115#_c_1746_n 0.0271337f $X=14.5 $Y=0.487
+ $X2=0 $Y2=0
cc_808 N_A_967_193#_c_811_n N_A_2388_115#_c_1733_n 0.00860154f $X=12.855 $Y=0.35
+ $X2=0 $Y2=0
cc_809 N_A_967_193#_c_812_n N_A_2388_115#_c_1733_n 0.00112873f $X=12.855 $Y=0.43
+ $X2=0 $Y2=0
cc_810 N_A_967_193#_c_814_n N_A_2388_115#_c_1734_n 0.0137064f $X=14.5 $Y=0.487
+ $X2=0 $Y2=0
cc_811 N_A_967_193#_c_815_n N_A_2388_115#_c_1734_n 0.00123001f $X=15.085
+ $Y=0.485 $X2=0 $Y2=0
cc_812 N_A_967_193#_c_818_n N_A_2388_115#_c_1734_n 0.00508318f $X=14.85 $Y=1.24
+ $X2=0 $Y2=0
cc_813 N_A_967_193#_c_803_n N_A_2168_439#_c_1839_n 0.00495156f $X=14.5 $Y=0.18
+ $X2=0 $Y2=0
cc_814 N_A_967_193#_c_813_n N_A_2168_439#_c_1839_n 2.24354e-19 $X=14.665 $Y=0.43
+ $X2=0 $Y2=0
cc_815 N_A_967_193#_c_814_n N_A_2168_439#_c_1839_n 0.00168671f $X=14.5 $Y=0.487
+ $X2=0 $Y2=0
cc_816 N_A_967_193#_c_815_n N_A_2168_439#_c_1839_n 0.00229599f $X=15.085
+ $Y=0.485 $X2=0 $Y2=0
cc_817 N_A_967_193#_c_810_n N_A_2168_439#_M1019_g 0.00809023f $X=15.085 $Y=1.93
+ $X2=0 $Y2=0
cc_818 N_A_967_193#_c_799_n N_A_2168_439#_c_1855_n 0.00596695f $X=11.55 $Y=0.18
+ $X2=0 $Y2=0
cc_819 N_A_967_193#_M1045_g N_A_2168_439#_c_1855_n 0.0226557f $X=11.625 $Y=0.915
+ $X2=0 $Y2=0
cc_820 N_A_967_193#_c_802_n N_A_2168_439#_c_1855_n 0.00312209f $X=12.69 $Y=0.18
+ $X2=0 $Y2=0
cc_821 N_A_967_193#_M1042_g N_A_2168_439#_c_1874_n 0.00960962f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_822 N_A_967_193#_M1045_g N_A_2168_439#_c_1856_n 0.00579323f $X=11.625
+ $Y=0.915 $X2=0 $Y2=0
cc_823 N_A_967_193#_M1042_g N_A_2168_439#_c_1876_n 0.00415241f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_824 N_A_967_193#_c_818_n N_A_2168_439#_c_1859_n 0.00591312f $X=14.85 $Y=1.24
+ $X2=0 $Y2=0
cc_825 N_A_967_193#_M1026_s N_A_2168_439#_c_1860_n 0.00508077f $X=14.94 $Y=0.235
+ $X2=0 $Y2=0
cc_826 N_A_967_193#_c_813_n N_A_2168_439#_c_1860_n 9.6494e-19 $X=14.665 $Y=0.43
+ $X2=0 $Y2=0
cc_827 N_A_967_193#_c_814_n N_A_2168_439#_c_1860_n 3.43233e-19 $X=14.5 $Y=0.487
+ $X2=0 $Y2=0
cc_828 N_A_967_193#_c_815_n N_A_2168_439#_c_1860_n 0.0519493f $X=15.085 $Y=0.485
+ $X2=0 $Y2=0
cc_829 N_A_967_193#_c_816_n N_A_2168_439#_c_1860_n 0.00400978f $X=14.85 $Y=1.405
+ $X2=0 $Y2=0
cc_830 N_A_967_193#_c_817_n N_A_2168_439#_c_1860_n 0.0385179f $X=15.085 $Y=1.405
+ $X2=0 $Y2=0
cc_831 N_A_967_193#_c_818_n N_A_2168_439#_c_1860_n 0.0126659f $X=14.85 $Y=1.24
+ $X2=0 $Y2=0
cc_832 N_A_967_193#_c_814_n N_A_2168_439#_c_1861_n 0.00687613f $X=14.5 $Y=0.487
+ $X2=0 $Y2=0
cc_833 N_A_967_193#_c_825_n N_A_2168_439#_c_1879_n 0.00126273f $X=11.235 $Y=3.06
+ $X2=0 $Y2=0
cc_834 N_A_967_193#_M1042_g N_A_2168_439#_c_1879_n 0.00620478f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_835 N_A_967_193#_M1042_g N_A_2168_439#_c_1880_n 0.00205837f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_836 N_A_967_193#_c_816_n N_A_2168_439#_c_1863_n 0.00132226f $X=14.85 $Y=1.405
+ $X2=0 $Y2=0
cc_837 N_A_967_193#_c_817_n N_A_2168_439#_c_1863_n 0.0255696f $X=15.085 $Y=1.405
+ $X2=0 $Y2=0
cc_838 N_A_967_193#_c_817_n N_A_2168_439#_c_1866_n 3.49205e-19 $X=15.085
+ $Y=1.405 $X2=0 $Y2=0
cc_839 N_A_967_193#_c_818_n N_A_2168_439#_c_1866_n 0.0139346f $X=14.85 $Y=1.24
+ $X2=0 $Y2=0
cc_840 N_A_967_193#_c_803_n N_CLK_M1026_g 0.031402f $X=14.5 $Y=0.18 $X2=0 $Y2=0
cc_841 N_A_967_193#_c_815_n N_CLK_M1026_g 0.00847086f $X=15.085 $Y=0.485 $X2=0
+ $Y2=0
cc_842 N_A_967_193#_c_816_n N_CLK_M1026_g 0.0214279f $X=14.85 $Y=1.405 $X2=0
+ $Y2=0
cc_843 N_A_967_193#_c_817_n N_CLK_M1026_g 0.00181527f $X=15.085 $Y=1.405 $X2=0
+ $Y2=0
cc_844 N_A_967_193#_c_810_n N_CLK_M1052_g 0.0299055f $X=15.085 $Y=1.93 $X2=0
+ $Y2=0
cc_845 N_A_967_193#_c_815_n N_CLK_M1027_g 0.00120041f $X=15.085 $Y=0.485 $X2=0
+ $Y2=0
cc_846 N_A_967_193#_c_817_n N_CLK_M1027_g 2.64121e-19 $X=15.085 $Y=1.405 $X2=0
+ $Y2=0
cc_847 N_A_967_193#_c_810_n N_CLK_M1055_g 0.00403175f $X=15.085 $Y=1.93 $X2=0
+ $Y2=0
cc_848 N_A_967_193#_c_810_n N_CLK_c_2085_n 0.0156558f $X=15.085 $Y=1.93 $X2=0
+ $Y2=0
cc_849 N_A_967_193#_c_817_n N_CLK_c_2085_n 0.0205799f $X=15.085 $Y=1.405 $X2=0
+ $Y2=0
cc_850 N_A_967_193#_c_810_n N_CLK_c_2086_n 0.0021084f $X=15.085 $Y=1.93 $X2=0
+ $Y2=0
cc_851 N_A_967_193#_c_817_n N_CLK_c_2086_n 0.00728284f $X=15.085 $Y=1.405 $X2=0
+ $Y2=0
cc_852 N_A_967_193#_M1025_g N_VPWR_c_2195_n 0.0210336f $X=9.275 $Y=2.465 $X2=0
+ $Y2=0
cc_853 N_A_967_193#_M1029_g N_VPWR_c_2195_n 0.00232677f $X=9.635 $Y=2.465 $X2=0
+ $Y2=0
cc_854 N_A_967_193#_c_796_n N_VPWR_c_2195_n 0.00596338f $X=9.79 $Y=1.42 $X2=0
+ $Y2=0
cc_855 N_A_967_193#_c_830_n N_VPWR_c_2195_n 0.0100097f $X=8.42 $Y=2.98 $X2=0
+ $Y2=0
cc_856 N_A_967_193#_c_832_n N_VPWR_c_2195_n 0.0480401f $X=8.505 $Y=2.895 $X2=0
+ $Y2=0
cc_857 N_A_967_193#_c_809_n N_VPWR_c_2195_n 0.023551f $X=9.1 $Y=1.51 $X2=0 $Y2=0
cc_858 N_A_967_193#_c_810_n N_VPWR_c_2198_n 0.0369704f $X=15.085 $Y=1.93 $X2=0
+ $Y2=0
cc_859 N_A_967_193#_c_830_n N_VPWR_c_2200_n 0.0483946f $X=8.42 $Y=2.98 $X2=0
+ $Y2=0
cc_860 N_A_967_193#_c_831_n N_VPWR_c_2200_n 0.0114622f $X=7.81 $Y=2.98 $X2=0
+ $Y2=0
cc_861 N_A_967_193#_c_810_n N_VPWR_c_2202_n 0.0220321f $X=15.085 $Y=1.93 $X2=0
+ $Y2=0
cc_862 N_A_967_193#_M1028_g N_VPWR_c_2206_n 0.00517164f $X=5.025 $Y=2.665 $X2=0
+ $Y2=0
cc_863 N_A_967_193#_M1025_g N_VPWR_c_2207_n 0.00486043f $X=9.275 $Y=2.465 $X2=0
+ $Y2=0
cc_864 N_A_967_193#_M1029_g N_VPWR_c_2207_n 0.0035993f $X=9.635 $Y=2.465 $X2=0
+ $Y2=0
cc_865 N_A_967_193#_c_826_n N_VPWR_c_2207_n 0.0244315f $X=10.33 $Y=3.06 $X2=0
+ $Y2=0
cc_866 N_A_967_193#_M1028_g N_VPWR_c_2191_n 0.00519032f $X=5.025 $Y=2.665 $X2=0
+ $Y2=0
cc_867 N_A_967_193#_M1025_g N_VPWR_c_2191_n 0.00814425f $X=9.275 $Y=2.465 $X2=0
+ $Y2=0
cc_868 N_A_967_193#_M1029_g N_VPWR_c_2191_n 0.00627252f $X=9.635 $Y=2.465 $X2=0
+ $Y2=0
cc_869 N_A_967_193#_c_825_n N_VPWR_c_2191_n 0.0308185f $X=11.235 $Y=3.06 $X2=0
+ $Y2=0
cc_870 N_A_967_193#_c_826_n N_VPWR_c_2191_n 0.0058694f $X=10.33 $Y=3.06 $X2=0
+ $Y2=0
cc_871 N_A_967_193#_c_830_n N_VPWR_c_2191_n 0.0293671f $X=8.42 $Y=2.98 $X2=0
+ $Y2=0
cc_872 N_A_967_193#_c_831_n N_VPWR_c_2191_n 0.00657784f $X=7.81 $Y=2.98 $X2=0
+ $Y2=0
cc_873 N_A_967_193#_c_810_n N_VPWR_c_2191_n 0.0125808f $X=15.085 $Y=1.93 $X2=0
+ $Y2=0
cc_874 N_A_967_193#_M1028_g N_A_342_261#_c_2422_n 5.03128e-19 $X=5.025 $Y=2.665
+ $X2=0 $Y2=0
cc_875 N_A_967_193#_c_792_n N_A_342_261#_c_2413_n 0.0012461f $X=5.1 $Y=2.142
+ $X2=0 $Y2=0
cc_876 N_A_967_193#_M1015_g N_A_342_261#_c_2414_n 0.00491952f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_877 N_A_967_193#_c_791_n N_A_342_261#_c_2414_n 0.011767f $X=5.825 $Y=2.142
+ $X2=0 $Y2=0
cc_878 N_A_967_193#_c_792_n N_A_342_261#_c_2414_n 0.00993017f $X=5.1 $Y=2.142
+ $X2=0 $Y2=0
cc_879 N_A_967_193#_M1015_g N_A_342_261#_c_2416_n 0.0171862f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_880 N_A_967_193#_c_798_n N_A_2081_439#_c_2552_n 0.00606218f $X=10.255
+ $Y=2.985 $X2=0 $Y2=0
cc_881 N_A_967_193#_M1042_g N_A_2081_439#_c_2552_n 0.00417858f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_882 N_A_967_193#_c_825_n N_A_2081_439#_c_2553_n 0.0103459f $X=11.235 $Y=3.06
+ $X2=0 $Y2=0
cc_883 N_A_967_193#_M1042_g N_A_2081_439#_c_2554_n 0.00235434f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_884 N_A_967_193#_c_825_n N_A_2081_439#_c_2555_n 0.0169947f $X=11.235 $Y=3.06
+ $X2=0 $Y2=0
cc_885 N_A_967_193#_M1042_g N_A_2081_439#_c_2555_n 0.00811813f $X=11.31 $Y=2.355
+ $X2=0 $Y2=0
cc_886 N_A_967_193#_c_810_n N_A_2523_397#_c_2584_n 0.0121616f $X=15.085 $Y=1.93
+ $X2=0 $Y2=0
cc_887 N_A_967_193#_c_817_n N_A_2523_397#_c_2584_n 4.03902e-19 $X=15.085
+ $Y=1.405 $X2=0 $Y2=0
cc_888 N_A_967_193#_c_810_n N_A_2523_397#_c_2587_n 0.0714654f $X=15.085 $Y=1.93
+ $X2=0 $Y2=0
cc_889 N_A_967_193#_M1057_g N_VGND_c_2684_n 0.00708683f $X=9.325 $Y=0.655 $X2=0
+ $Y2=0
cc_890 N_A_967_193#_M1045_g N_VGND_c_2685_n 0.00856041f $X=11.625 $Y=0.915 $X2=0
+ $Y2=0
cc_891 N_A_967_193#_c_802_n N_VGND_c_2685_n 0.0259201f $X=12.69 $Y=0.18 $X2=0
+ $Y2=0
cc_892 N_A_967_193#_c_811_n N_VGND_c_2685_n 0.0250186f $X=12.855 $Y=0.35 $X2=0
+ $Y2=0
cc_893 N_A_967_193#_c_812_n N_VGND_c_2685_n 0.00760374f $X=12.855 $Y=0.43 $X2=0
+ $Y2=0
cc_894 N_A_967_193#_c_815_n N_VGND_c_2686_n 0.0157205f $X=15.085 $Y=0.485 $X2=0
+ $Y2=0
cc_895 N_A_967_193#_c_802_n N_VGND_c_2690_n 0.0527574f $X=12.69 $Y=0.18 $X2=0
+ $Y2=0
cc_896 N_A_967_193#_c_811_n N_VGND_c_2690_n 0.0199384f $X=12.855 $Y=0.35 $X2=0
+ $Y2=0
cc_897 N_A_967_193#_c_814_n N_VGND_c_2690_n 0.135113f $X=14.5 $Y=0.487 $X2=0
+ $Y2=0
cc_898 N_A_967_193#_M1057_g N_VGND_c_2695_n 0.00426565f $X=9.325 $Y=0.655 $X2=0
+ $Y2=0
cc_899 N_A_967_193#_M1010_g N_VGND_c_2695_n 0.00416934f $X=9.715 $Y=0.655 $X2=0
+ $Y2=0
cc_900 N_A_967_193#_c_800_n N_VGND_c_2695_n 0.0595572f $X=10.33 $Y=0.18 $X2=0
+ $Y2=0
cc_901 N_A_967_193#_M1026_s N_VGND_c_2698_n 0.002305f $X=14.94 $Y=0.235 $X2=0
+ $Y2=0
cc_902 N_A_967_193#_M1057_g N_VGND_c_2698_n 0.00721123f $X=9.325 $Y=0.655 $X2=0
+ $Y2=0
cc_903 N_A_967_193#_M1010_g N_VGND_c_2698_n 0.00600684f $X=9.715 $Y=0.655 $X2=0
+ $Y2=0
cc_904 N_A_967_193#_c_799_n N_VGND_c_2698_n 0.0431249f $X=11.55 $Y=0.18 $X2=0
+ $Y2=0
cc_905 N_A_967_193#_c_800_n N_VGND_c_2698_n 0.0104031f $X=10.33 $Y=0.18 $X2=0
+ $Y2=0
cc_906 N_A_967_193#_c_802_n N_VGND_c_2698_n 0.0260478f $X=12.69 $Y=0.18 $X2=0
+ $Y2=0
cc_907 N_A_967_193#_c_803_n N_VGND_c_2698_n 0.0439564f $X=14.5 $Y=0.18 $X2=0
+ $Y2=0
cc_908 N_A_967_193#_c_806_n N_VGND_c_2698_n 0.00416972f $X=11.625 $Y=0.18 $X2=0
+ $Y2=0
cc_909 N_A_967_193#_c_807_n N_VGND_c_2698_n 0.00778385f $X=12.855 $Y=0.18 $X2=0
+ $Y2=0
cc_910 N_A_967_193#_c_811_n N_VGND_c_2698_n 0.01095f $X=12.855 $Y=0.35 $X2=0
+ $Y2=0
cc_911 N_A_967_193#_c_814_n N_VGND_c_2698_n 0.0763668f $X=14.5 $Y=0.487 $X2=0
+ $Y2=0
cc_912 N_A_967_193#_M1015_g N_A_824_219#_c_2941_n 0.00824316f $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_913 N_A_967_193#_M1015_g N_A_824_219#_c_2944_n 2.13168e-19 $X=4.91 $Y=1.305
+ $X2=0 $Y2=0
cc_914 N_A_1147_490#_c_1102_n N_RESET_B_c_1288_n 0.00881852f $X=6.35 $Y=1.125
+ $X2=0 $Y2=0
cc_915 N_A_1147_490#_c_1104_n N_RESET_B_M1043_g 0.00758113f $X=6.365 $Y=2.525
+ $X2=0 $Y2=0
cc_916 N_A_1147_490#_c_1092_n N_RESET_B_M1005_g 0.0130892f $X=7.85 $Y=1.15 $X2=0
+ $Y2=0
cc_917 N_A_1147_490#_c_1098_n N_RESET_B_M1005_g 0.00102347f $X=6.35 $Y=1.15
+ $X2=0 $Y2=0
cc_918 N_A_1147_490#_c_1102_n N_RESET_B_M1005_g 0.0516466f $X=6.35 $Y=1.125
+ $X2=0 $Y2=0
cc_919 N_A_1147_490#_c_1091_n N_RESET_B_c_1311_n 0.00259619f $X=6.44 $Y=2.45
+ $X2=0 $Y2=0
cc_920 N_A_1147_490#_M1002_s N_RESET_B_c_1313_n 0.00297368f $X=7.93 $Y=1.875
+ $X2=0 $Y2=0
cc_921 N_A_1147_490#_M1042_d N_RESET_B_c_1313_n 0.0039379f $X=11.385 $Y=1.935
+ $X2=0 $Y2=0
cc_922 N_A_1147_490#_c_1093_n N_RESET_B_c_1313_n 0.0237758f $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_923 N_A_1147_490#_c_1095_n N_RESET_B_c_1313_n 0.0234299f $X=9.5 $Y=2.895
+ $X2=0 $Y2=0
cc_924 N_A_1147_490#_c_1109_n N_RESET_B_c_1313_n 0.0126921f $X=10.115 $Y=2.98
+ $X2=0 $Y2=0
cc_925 N_A_1147_490#_c_1110_n N_RESET_B_c_1313_n 0.0176424f $X=10.2 $Y=2.895
+ $X2=0 $Y2=0
cc_926 N_A_1147_490#_c_1111_n N_RESET_B_c_1313_n 0.0214481f $X=11.08 $Y=2.03
+ $X2=0 $Y2=0
cc_927 N_A_1147_490#_c_1114_n N_RESET_B_c_1313_n 0.0139003f $X=11.165 $Y=2.08
+ $X2=0 $Y2=0
cc_928 N_A_1147_490#_c_1091_n N_RESET_B_c_1318_n 0.00758113f $X=6.44 $Y=2.45
+ $X2=0 $Y2=0
cc_929 N_A_1147_490#_c_1099_n N_RESET_B_c_1318_n 0.0516466f $X=6.35 $Y=1.29
+ $X2=0 $Y2=0
cc_930 N_A_1147_490#_c_1091_n N_RESET_B_c_1319_n 0.00144432f $X=6.44 $Y=2.45
+ $X2=0 $Y2=0
cc_931 N_A_1147_490#_c_1093_n N_A_911_219#_c_1543_n 0.0131866f $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_932 N_A_1147_490#_c_1100_n N_A_911_219#_c_1543_n 0.00572384f $X=8.015
+ $Y=0.855 $X2=0 $Y2=0
cc_933 N_A_1147_490#_c_1092_n N_A_911_219#_M1000_g 5.78457e-19 $X=7.85 $Y=1.15
+ $X2=0 $Y2=0
cc_934 N_A_1147_490#_c_1093_n N_A_911_219#_M1000_g 0.00555232f $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_935 N_A_1147_490#_c_1094_n N_A_911_219#_M1000_g 0.00789001f $X=9.415 $Y=1.08
+ $X2=0 $Y2=0
cc_936 N_A_1147_490#_c_1100_n N_A_911_219#_M1000_g 0.016213f $X=8.015 $Y=0.855
+ $X2=0 $Y2=0
cc_937 N_A_1147_490#_c_1093_n N_A_911_219#_M1002_g 0.0195313f $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_938 N_A_1147_490#_c_1094_n N_A_911_219#_c_1546_n 0.00119926f $X=9.415 $Y=1.08
+ $X2=0 $Y2=0
cc_939 N_A_1147_490#_c_1094_n N_A_911_219#_M1021_g 0.0114672f $X=9.415 $Y=1.08
+ $X2=0 $Y2=0
cc_940 N_A_1147_490#_c_1100_n N_A_911_219#_M1021_g 0.00229777f $X=8.015 $Y=0.855
+ $X2=0 $Y2=0
cc_941 N_A_1147_490#_c_1093_n N_A_911_219#_M1009_g 9.94249e-19 $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_942 N_A_1147_490#_c_1093_n N_A_911_219#_c_1549_n 0.0047893f $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_943 N_A_1147_490#_c_1098_n N_A_911_219#_c_1551_n 0.00518802f $X=6.35 $Y=1.15
+ $X2=0 $Y2=0
cc_944 N_A_1147_490#_c_1099_n N_A_911_219#_c_1551_n 0.00353702f $X=6.35 $Y=1.29
+ $X2=0 $Y2=0
cc_945 N_A_1147_490#_c_1091_n N_A_911_219#_c_1552_n 0.00178512f $X=6.44 $Y=2.45
+ $X2=0 $Y2=0
cc_946 N_A_1147_490#_c_1099_n N_A_911_219#_c_1552_n 0.00130336f $X=6.35 $Y=1.29
+ $X2=0 $Y2=0
cc_947 N_A_1147_490#_c_1091_n N_A_911_219#_c_1553_n 0.00593585f $X=6.44 $Y=2.45
+ $X2=0 $Y2=0
cc_948 N_A_1147_490#_c_1091_n N_A_911_219#_c_1554_n 0.0122168f $X=6.44 $Y=2.45
+ $X2=0 $Y2=0
cc_949 N_A_1147_490#_c_1092_n N_A_911_219#_c_1554_n 0.046762f $X=7.85 $Y=1.15
+ $X2=0 $Y2=0
cc_950 N_A_1147_490#_c_1098_n N_A_911_219#_c_1554_n 0.024097f $X=6.35 $Y=1.15
+ $X2=0 $Y2=0
cc_951 N_A_1147_490#_c_1099_n N_A_911_219#_c_1554_n 0.00443958f $X=6.35 $Y=1.29
+ $X2=0 $Y2=0
cc_952 N_A_1147_490#_c_1104_n N_A_911_219#_c_1565_n 0.0157355f $X=6.365 $Y=2.525
+ $X2=0 $Y2=0
cc_953 N_A_1147_490#_c_1105_n N_A_911_219#_c_1565_n 0.00718943f $X=5.885
+ $Y=2.525 $X2=0 $Y2=0
cc_954 N_A_1147_490#_c_1091_n N_A_911_219#_c_1565_n 0.00450492f $X=6.44 $Y=2.45
+ $X2=0 $Y2=0
cc_955 N_A_1147_490#_c_1103_n N_A_911_219#_c_1566_n 0.00243485f $X=5.81 $Y=2.6
+ $X2=0 $Y2=0
cc_956 N_A_1147_490#_c_1104_n N_A_911_219#_c_1566_n 0.00538873f $X=6.365
+ $Y=2.525 $X2=0 $Y2=0
cc_957 N_A_1147_490#_c_1103_n N_A_911_219#_c_1653_n 9.11999e-19 $X=5.81 $Y=2.6
+ $X2=0 $Y2=0
cc_958 N_A_1147_490#_c_1092_n N_A_911_219#_c_1568_n 0.0235511f $X=7.85 $Y=1.15
+ $X2=0 $Y2=0
cc_959 N_A_1147_490#_c_1093_n N_A_911_219#_c_1568_n 0.0217731f $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_960 N_A_1147_490#_c_1092_n N_A_911_219#_c_1557_n 0.00900288f $X=7.85 $Y=1.15
+ $X2=0 $Y2=0
cc_961 N_A_1147_490#_c_1093_n N_A_911_219#_c_1557_n 0.00142037f $X=8.075 $Y=2.02
+ $X2=0 $Y2=0
cc_962 N_A_1147_490#_c_1097_n N_A_2388_115#_c_1736_n 5.40467e-19 $X=11.165
+ $Y=1.915 $X2=0 $Y2=0
cc_963 N_A_1147_490#_c_1101_n N_A_2168_439#_M1051_d 0.00265622f $X=11.165
+ $Y=1.17 $X2=-0.19 $Y2=-0.245
cc_964 N_A_1147_490#_c_1111_n N_A_2168_439#_M1044_d 0.00373773f $X=11.08 $Y=2.03
+ $X2=0 $Y2=0
cc_965 N_A_1147_490#_c_1114_n N_A_2168_439#_M1044_d 0.00143183f $X=11.165
+ $Y=2.08 $X2=0 $Y2=0
cc_966 N_A_1147_490#_c_1096_n N_A_2168_439#_c_1855_n 0.0139162f $X=10.785
+ $Y=0.74 $X2=0 $Y2=0
cc_967 N_A_1147_490#_c_1101_n N_A_2168_439#_c_1855_n 0.0044527f $X=11.165
+ $Y=1.17 $X2=0 $Y2=0
cc_968 N_A_1147_490#_M1042_d N_A_2168_439#_c_1874_n 0.00588487f $X=11.385
+ $Y=1.935 $X2=0 $Y2=0
cc_969 N_A_1147_490#_c_1114_n N_A_2168_439#_c_1874_n 0.0128543f $X=11.165
+ $Y=2.08 $X2=0 $Y2=0
cc_970 N_A_1147_490#_c_1097_n N_A_2168_439#_c_1856_n 0.0165442f $X=11.165
+ $Y=1.915 $X2=0 $Y2=0
cc_971 N_A_1147_490#_c_1101_n N_A_2168_439#_c_1856_n 0.00593205f $X=11.165
+ $Y=1.17 $X2=0 $Y2=0
cc_972 N_A_1147_490#_c_1114_n N_A_2168_439#_c_1876_n 0.0253514f $X=11.165
+ $Y=2.08 $X2=0 $Y2=0
cc_973 N_A_1147_490#_c_1111_n N_A_2168_439#_c_1879_n 0.00496444f $X=11.08
+ $Y=2.03 $X2=0 $Y2=0
cc_974 N_A_1147_490#_c_1114_n N_A_2168_439#_c_1879_n 0.00790462f $X=11.165
+ $Y=2.08 $X2=0 $Y2=0
cc_975 N_A_1147_490#_c_1097_n N_A_2168_439#_c_1880_n 0.00599428f $X=11.165
+ $Y=1.915 $X2=0 $Y2=0
cc_976 N_A_1147_490#_c_1103_n N_VPWR_c_2194_n 0.0215433f $X=5.81 $Y=2.6 $X2=0
+ $Y2=0
cc_977 N_A_1147_490#_c_1104_n N_VPWR_c_2194_n 0.00616387f $X=6.365 $Y=2.525
+ $X2=0 $Y2=0
cc_978 N_A_1147_490#_c_1095_n N_VPWR_c_2195_n 0.0692829f $X=9.5 $Y=2.895 $X2=0
+ $Y2=0
cc_979 N_A_1147_490#_c_1184_n N_VPWR_c_2195_n 0.0128808f $X=9.585 $Y=2.98 $X2=0
+ $Y2=0
cc_980 N_A_1147_490#_c_1104_n N_VPWR_c_2200_n 0.00335648f $X=6.365 $Y=2.525
+ $X2=0 $Y2=0
cc_981 N_A_1147_490#_c_1103_n N_VPWR_c_2206_n 0.00486043f $X=5.81 $Y=2.6 $X2=0
+ $Y2=0
cc_982 N_A_1147_490#_c_1109_n N_VPWR_c_2207_n 0.0410341f $X=10.115 $Y=2.98 $X2=0
+ $Y2=0
cc_983 N_A_1147_490#_c_1184_n N_VPWR_c_2207_n 0.00925931f $X=9.585 $Y=2.98 $X2=0
+ $Y2=0
cc_984 N_A_1147_490#_c_1103_n N_VPWR_c_2191_n 0.00588254f $X=5.81 $Y=2.6 $X2=0
+ $Y2=0
cc_985 N_A_1147_490#_c_1104_n N_VPWR_c_2191_n 0.00396575f $X=6.365 $Y=2.525
+ $X2=0 $Y2=0
cc_986 N_A_1147_490#_c_1109_n N_VPWR_c_2191_n 0.0253219f $X=10.115 $Y=2.98 $X2=0
+ $Y2=0
cc_987 N_A_1147_490#_c_1184_n N_VPWR_c_2191_n 0.0064524f $X=9.585 $Y=2.98 $X2=0
+ $Y2=0
cc_988 N_A_1147_490#_c_1095_n A_1870_367# 0.00860146f $X=9.5 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_989 N_A_1147_490#_c_1184_n A_1870_367# 0.00237462f $X=9.585 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_990 N_A_1147_490#_c_1110_n N_A_2081_439#_c_2552_n 0.0410255f $X=10.2 $Y=2.895
+ $X2=0 $Y2=0
cc_991 N_A_1147_490#_c_1111_n N_A_2081_439#_c_2552_n 0.0153675f $X=11.08 $Y=2.03
+ $X2=0 $Y2=0
cc_992 N_A_1147_490#_c_1109_n N_A_2081_439#_c_2553_n 0.0141092f $X=10.115
+ $Y=2.98 $X2=0 $Y2=0
cc_993 N_A_1147_490#_c_1094_n N_VGND_M1021_d 0.00566574f $X=9.415 $Y=1.08 $X2=0
+ $Y2=0
cc_994 N_A_1147_490#_c_1096_n N_VGND_c_2695_n 0.00739145f $X=10.785 $Y=0.74
+ $X2=0 $Y2=0
cc_995 N_A_1147_490#_c_1096_n N_VGND_c_2698_n 0.00896868f $X=10.785 $Y=0.74
+ $X2=0 $Y2=0
cc_996 N_A_1147_490#_c_1098_n N_A_824_219#_c_2942_n 0.0130623f $X=6.35 $Y=1.15
+ $X2=0 $Y2=0
cc_997 N_A_1147_490#_c_1099_n N_A_824_219#_c_2942_n 9.50186e-19 $X=6.35 $Y=1.29
+ $X2=0 $Y2=0
cc_998 N_A_1147_490#_c_1102_n N_A_824_219#_c_2942_n 0.00237631f $X=6.35 $Y=1.125
+ $X2=0 $Y2=0
cc_999 N_A_1147_490#_c_1102_n N_A_824_219#_c_2944_n 0.00282534f $X=6.35 $Y=1.125
+ $X2=0 $Y2=0
cc_1000 N_A_1147_490#_c_1094_n A_1661_87# 0.00185339f $X=9.415 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_1001 N_A_1147_490#_c_1094_n A_1880_47# 0.00143193f $X=9.415 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_1002 N_RESET_B_c_1311_n N_A_911_219#_M1006_d 0.00608559f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1003 N_RESET_B_c_1313_n N_A_911_219#_M1002_g 0.00718921f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1004 N_RESET_B_c_1313_n N_A_911_219#_M1009_g 0.0121332f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1005 N_RESET_B_c_1311_n N_A_911_219#_c_1561_n 0.0371566f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1006 N_RESET_B_c_1311_n N_A_911_219#_c_1562_n 0.0125676f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1007 N_RESET_B_c_1311_n N_A_911_219#_c_1553_n 0.00861089f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1008 N_RESET_B_M1005_g N_A_911_219#_c_1554_n 0.0121418f $X=6.83 $Y=0.805
+ $X2=0 $Y2=0
cc_1009 N_RESET_B_c_1311_n N_A_911_219#_c_1565_n 0.0437026f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1010 N_RESET_B_c_1314_n N_A_911_219#_c_1565_n 3.28223e-19 $X=7.105 $Y=2.405
+ $X2=0 $Y2=0
cc_1011 N_RESET_B_c_1318_n N_A_911_219#_c_1565_n 0.0016559f $X=6.92 $Y=2.35
+ $X2=0 $Y2=0
cc_1012 N_RESET_B_c_1319_n N_A_911_219#_c_1565_n 0.00768209f $X=6.92 $Y=2.35
+ $X2=0 $Y2=0
cc_1013 N_RESET_B_M1043_g N_A_911_219#_c_1566_n 0.00421471f $X=6.8 $Y=2.885
+ $X2=0 $Y2=0
cc_1014 N_RESET_B_M1043_g N_A_911_219#_c_1619_n 0.0122284f $X=6.8 $Y=2.885 $X2=0
+ $Y2=0
cc_1015 N_RESET_B_M1049_g N_A_911_219#_c_1619_n 0.0090114f $X=7.16 $Y=2.885
+ $X2=0 $Y2=0
cc_1016 N_RESET_B_c_1311_n N_A_911_219#_c_1619_n 0.00655905f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1017 N_RESET_B_c_1313_n N_A_911_219#_c_1619_n 0.00254728f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1018 N_RESET_B_c_1314_n N_A_911_219#_c_1619_n 0.00258123f $X=7.105 $Y=2.405
+ $X2=0 $Y2=0
cc_1019 N_RESET_B_c_1318_n N_A_911_219#_c_1619_n 2.05922e-19 $X=6.92 $Y=2.35
+ $X2=0 $Y2=0
cc_1020 N_RESET_B_c_1319_n N_A_911_219#_c_1619_n 0.0167307f $X=6.92 $Y=2.35
+ $X2=0 $Y2=0
cc_1021 N_RESET_B_c_1293_n N_A_911_219#_c_1555_n 4.59109e-19 $X=4.03 $Y=1.625
+ $X2=0 $Y2=0
cc_1022 N_RESET_B_c_1311_n N_A_911_219#_c_1567_n 0.00910342f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1023 N_RESET_B_M1043_g N_A_911_219#_c_1622_n 0.00105898f $X=6.8 $Y=2.885
+ $X2=0 $Y2=0
cc_1024 N_RESET_B_M1049_g N_A_911_219#_c_1622_n 0.00489679f $X=7.16 $Y=2.885
+ $X2=0 $Y2=0
cc_1025 N_RESET_B_c_1313_n N_A_911_219#_c_1622_n 0.00751655f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1026 N_RESET_B_M1005_g N_A_911_219#_c_1568_n 7.60322e-19 $X=6.83 $Y=0.805
+ $X2=0 $Y2=0
cc_1027 N_RESET_B_c_1313_n N_A_911_219#_c_1568_n 7.25494e-19 $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1028 N_RESET_B_M1005_g N_A_911_219#_c_1557_n 0.00662185f $X=6.83 $Y=0.805
+ $X2=0 $Y2=0
cc_1029 N_RESET_B_c_1313_n N_A_2388_115#_M1037_d 0.00190347f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1030 N_RESET_B_M1038_g N_A_2388_115#_c_1738_n 0.00597725f $X=13.52 $Y=2.8
+ $X2=0 $Y2=0
cc_1031 N_RESET_B_M1036_g N_A_2388_115#_c_1738_n 5.53294e-19 $X=13.88 $Y=2.8
+ $X2=0 $Y2=0
cc_1032 N_RESET_B_c_1296_n N_A_2388_115#_c_1738_n 4.85115e-19 $X=13.52 $Y=1.7
+ $X2=0 $Y2=0
cc_1033 N_RESET_B_c_1313_n N_A_2388_115#_c_1738_n 0.0497875f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1034 N_RESET_B_c_1316_n N_A_2388_115#_c_1738_n 0.00519122f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1035 N_RESET_B_M1054_g N_A_2388_115#_c_1746_n 0.0134417f $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1036 N_RESET_B_M1038_g N_A_2388_115#_c_1739_n 0.00762341f $X=13.52 $Y=2.8
+ $X2=0 $Y2=0
cc_1037 N_RESET_B_M1036_g N_A_2388_115#_c_1739_n 0.0013214f $X=13.88 $Y=2.8
+ $X2=0 $Y2=0
cc_1038 N_RESET_B_c_1313_n N_A_2388_115#_c_1740_n 0.0194407f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1039 N_RESET_B_c_1313_n N_A_2388_115#_c_1741_n 0.00426141f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1040 N_RESET_B_M1054_g N_A_2388_115#_c_1733_n 0.00479215f $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1041 N_RESET_B_c_1313_n N_A_2168_439#_M1044_d 0.00426168f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1042 N_RESET_B_c_1313_n N_A_2168_439#_M1037_g 0.00286958f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1043 N_RESET_B_c_1316_n N_A_2168_439#_M1037_g 9.29081e-19 $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1044 N_RESET_B_c_1320_n N_A_2168_439#_M1037_g 0.0106184f $X=13.88 $Y=2.265
+ $X2=0 $Y2=0
cc_1045 N_RESET_B_M1054_g N_A_2168_439#_c_1839_n 0.0465889f $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1046 N_RESET_B_c_1320_n N_A_2168_439#_c_1841_n 0.00324605f $X=13.88 $Y=2.265
+ $X2=0 $Y2=0
cc_1047 N_RESET_B_M1036_g N_A_2168_439#_M1019_g 0.0167077f $X=13.88 $Y=2.8 $X2=0
+ $Y2=0
cc_1048 N_RESET_B_c_1296_n N_A_2168_439#_M1019_g 0.00943348f $X=13.52 $Y=1.7
+ $X2=0 $Y2=0
cc_1049 N_RESET_B_c_1315_n N_A_2168_439#_M1019_g 0.00541727f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1050 N_RESET_B_c_1316_n N_A_2168_439#_M1019_g 0.0106178f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1051 N_RESET_B_c_1320_n N_A_2168_439#_M1019_g 0.0181356f $X=13.88 $Y=2.265
+ $X2=0 $Y2=0
cc_1052 N_RESET_B_c_1313_n N_A_2168_439#_c_1874_n 0.0209187f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1053 N_RESET_B_c_1313_n N_A_2168_439#_c_1876_n 0.0146265f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1054 N_RESET_B_c_1313_n N_A_2168_439#_c_1877_n 0.011912f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1055 N_RESET_B_M1054_g N_A_2168_439#_c_1938_n 0.00121316f $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1056 N_RESET_B_M1054_g N_A_2168_439#_c_1857_n 0.0184118f $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1057 N_RESET_B_c_1306_n N_A_2168_439#_c_1857_n 0.0106184f $X=13.52 $Y=2.1
+ $X2=0 $Y2=0
cc_1058 N_RESET_B_c_1313_n N_A_2168_439#_c_1879_n 0.0100144f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1059 N_RESET_B_M1054_g N_A_2168_439#_c_1862_n 0.0136429f $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1060 N_RESET_B_c_1296_n N_A_2168_439#_c_1862_n 0.00532141f $X=13.52 $Y=1.7
+ $X2=0 $Y2=0
cc_1061 N_RESET_B_M1054_g N_A_2168_439#_c_1863_n 5.09934e-19 $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1062 N_RESET_B_M1054_g N_A_2168_439#_c_1866_n 0.00219464f $X=13.335 $Y=0.915
+ $X2=0 $Y2=0
cc_1063 N_RESET_B_c_1313_n N_VPWR_M1009_d 0.0130079f $X=14.015 $Y=2.405 $X2=0
+ $Y2=0
cc_1064 N_RESET_B_c_1299_n N_VPWR_c_2193_n 0.00623553f $X=3.6 $Y=2.345 $X2=0
+ $Y2=0
cc_1065 N_RESET_B_M1043_g N_VPWR_c_2194_n 0.00801732f $X=6.8 $Y=2.885 $X2=0
+ $Y2=0
cc_1066 N_RESET_B_c_1311_n N_VPWR_c_2194_n 0.00231493f $X=6.815 $Y=2.405 $X2=0
+ $Y2=0
cc_1067 N_RESET_B_c_1313_n N_VPWR_c_2195_n 0.0423883f $X=14.015 $Y=2.405 $X2=0
+ $Y2=0
cc_1068 N_RESET_B_M1038_g N_VPWR_c_2196_n 0.00252391f $X=13.52 $Y=2.8 $X2=0
+ $Y2=0
cc_1069 N_RESET_B_c_1313_n N_VPWR_c_2196_n 0.00203166f $X=14.015 $Y=2.405 $X2=0
+ $Y2=0
cc_1070 N_RESET_B_M1038_g N_VPWR_c_2197_n 0.00163177f $X=13.52 $Y=2.8 $X2=0
+ $Y2=0
cc_1071 N_RESET_B_M1036_g N_VPWR_c_2197_n 0.00934419f $X=13.88 $Y=2.8 $X2=0
+ $Y2=0
cc_1072 N_RESET_B_c_1313_n N_VPWR_c_2197_n 6.28884e-19 $X=14.015 $Y=2.405 $X2=0
+ $Y2=0
cc_1073 N_RESET_B_c_1315_n N_VPWR_c_2197_n 0.00464341f $X=14.16 $Y=2.405 $X2=0
+ $Y2=0
cc_1074 N_RESET_B_c_1316_n N_VPWR_c_2197_n 0.0153312f $X=14.16 $Y=2.405 $X2=0
+ $Y2=0
cc_1075 N_RESET_B_M1043_g N_VPWR_c_2200_n 0.00397042f $X=6.8 $Y=2.885 $X2=0
+ $Y2=0
cc_1076 N_RESET_B_M1049_g N_VPWR_c_2200_n 0.00392332f $X=7.16 $Y=2.885 $X2=0
+ $Y2=0
cc_1077 N_RESET_B_c_1299_n N_VPWR_c_2206_n 0.00377843f $X=3.6 $Y=2.345 $X2=0
+ $Y2=0
cc_1078 N_RESET_B_c_1302_n N_VPWR_c_2206_n 0.00377907f $X=3.99 $Y=2.345 $X2=0
+ $Y2=0
cc_1079 N_RESET_B_M1038_g N_VPWR_c_2208_n 0.00473334f $X=13.52 $Y=2.8 $X2=0
+ $Y2=0
cc_1080 N_RESET_B_M1036_g N_VPWR_c_2208_n 0.00418439f $X=13.88 $Y=2.8 $X2=0
+ $Y2=0
cc_1081 N_RESET_B_c_1299_n N_VPWR_c_2191_n 0.006036f $X=3.6 $Y=2.345 $X2=0 $Y2=0
cc_1082 N_RESET_B_c_1302_n N_VPWR_c_2191_n 0.00676694f $X=3.99 $Y=2.345 $X2=0
+ $Y2=0
cc_1083 N_RESET_B_M1043_g N_VPWR_c_2191_n 0.00683083f $X=6.8 $Y=2.885 $X2=0
+ $Y2=0
cc_1084 N_RESET_B_M1049_g N_VPWR_c_2191_n 0.00678531f $X=7.16 $Y=2.885 $X2=0
+ $Y2=0
cc_1085 N_RESET_B_M1038_g N_VPWR_c_2191_n 0.00957559f $X=13.52 $Y=2.8 $X2=0
+ $Y2=0
cc_1086 N_RESET_B_M1036_g N_VPWR_c_2191_n 0.00402597f $X=13.88 $Y=2.8 $X2=0
+ $Y2=0
cc_1087 N_RESET_B_c_1316_n N_VPWR_c_2191_n 0.0121256f $X=14.16 $Y=2.405 $X2=0
+ $Y2=0
cc_1088 N_RESET_B_c_1311_n N_A_342_261#_M1048_d 0.00124344f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1089 N_RESET_B_c_1312_n N_A_342_261#_M1048_d 0.00123465f $X=4.225 $Y=2.405
+ $X2=0 $Y2=0
cc_1090 N_RESET_B_c_1298_n N_A_342_261#_M1048_d 6.87532e-19 $X=4.03 $Y=1.79
+ $X2=0 $Y2=0
cc_1091 N_RESET_B_c_1286_n N_A_342_261#_c_2412_n 0.0054062f $X=3.675 $Y=2.27
+ $X2=0 $Y2=0
cc_1092 N_RESET_B_c_1294_n N_A_342_261#_c_2412_n 0.00106989f $X=4.03 $Y=2.195
+ $X2=0 $Y2=0
cc_1093 N_RESET_B_c_1298_n N_A_342_261#_c_2412_n 0.00885661f $X=4.03 $Y=1.79
+ $X2=0 $Y2=0
cc_1094 N_RESET_B_c_1299_n N_A_342_261#_c_2421_n 0.0101095f $X=3.6 $Y=2.345
+ $X2=0 $Y2=0
cc_1095 N_RESET_B_c_1286_n N_A_342_261#_c_2421_n 0.00100477f $X=3.675 $Y=2.27
+ $X2=0 $Y2=0
cc_1096 N_RESET_B_c_1302_n N_A_342_261#_c_2421_n 0.00112446f $X=3.99 $Y=2.345
+ $X2=0 $Y2=0
cc_1097 N_RESET_B_c_1312_n N_A_342_261#_c_2421_n 0.00110457f $X=4.225 $Y=2.405
+ $X2=0 $Y2=0
cc_1098 N_RESET_B_c_1298_n N_A_342_261#_c_2421_n 0.00710053f $X=4.03 $Y=1.79
+ $X2=0 $Y2=0
cc_1099 N_RESET_B_c_1299_n N_A_342_261#_c_2422_n 0.0110328f $X=3.6 $Y=2.345
+ $X2=0 $Y2=0
cc_1100 N_RESET_B_c_1285_n N_A_342_261#_c_2422_n 0.00178753f $X=3.865 $Y=2.27
+ $X2=0 $Y2=0
cc_1101 N_RESET_B_c_1302_n N_A_342_261#_c_2422_n 0.0106079f $X=3.99 $Y=2.345
+ $X2=0 $Y2=0
cc_1102 N_RESET_B_c_1295_n N_A_342_261#_c_2422_n 5.10219e-19 $X=4.03 $Y=2.27
+ $X2=0 $Y2=0
cc_1103 N_RESET_B_c_1311_n N_A_342_261#_c_2422_n 0.00670633f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1104 N_RESET_B_c_1312_n N_A_342_261#_c_2422_n 0.00350252f $X=4.225 $Y=2.405
+ $X2=0 $Y2=0
cc_1105 N_RESET_B_c_1298_n N_A_342_261#_c_2422_n 0.0146528f $X=4.03 $Y=1.79
+ $X2=0 $Y2=0
cc_1106 N_RESET_B_c_1299_n N_A_342_261#_c_2489_n 0.0052893f $X=3.6 $Y=2.345
+ $X2=0 $Y2=0
cc_1107 N_RESET_B_c_1302_n N_A_342_261#_c_2413_n 2.74071e-19 $X=3.99 $Y=2.345
+ $X2=0 $Y2=0
cc_1108 N_RESET_B_c_1295_n N_A_342_261#_c_2413_n 8.01826e-19 $X=4.03 $Y=2.27
+ $X2=0 $Y2=0
cc_1109 N_RESET_B_c_1311_n N_A_342_261#_c_2413_n 0.0224024f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1110 N_RESET_B_c_1312_n N_A_342_261#_c_2413_n 0.00264827f $X=4.225 $Y=2.405
+ $X2=0 $Y2=0
cc_1111 N_RESET_B_c_1298_n N_A_342_261#_c_2413_n 0.0199554f $X=4.03 $Y=1.79
+ $X2=0 $Y2=0
cc_1112 N_RESET_B_c_1311_n N_A_342_261#_c_2414_n 0.023388f $X=6.815 $Y=2.405
+ $X2=0 $Y2=0
cc_1113 N_RESET_B_c_1294_n N_A_342_261#_c_2415_n 0.0010467f $X=4.03 $Y=2.195
+ $X2=0 $Y2=0
cc_1114 N_RESET_B_c_1298_n N_A_342_261#_c_2415_n 0.0136966f $X=4.03 $Y=1.79
+ $X2=0 $Y2=0
cc_1115 N_RESET_B_c_1313_n A_1673_375# 0.00263244f $X=14.015 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_1116 N_RESET_B_c_1313_n A_1870_367# 0.00502061f $X=14.015 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_1117 N_RESET_B_c_1313_n N_A_2081_439#_M1044_s 0.00188511f $X=14.015 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_1118 N_RESET_B_c_1313_n N_A_2081_439#_c_2552_n 0.0181936f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1119 N_RESET_B_c_1313_n N_A_2081_439#_c_2554_n 0.00727962f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1120 N_RESET_B_c_1313_n N_A_2081_439#_c_2555_n 0.0135295f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1121 N_RESET_B_c_1313_n N_A_2523_397#_M1037_s 0.00210586f $X=14.015 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_1122 N_RESET_B_c_1306_n N_A_2523_397#_c_2582_n 0.00243519f $X=13.52 $Y=2.1
+ $X2=0 $Y2=0
cc_1123 N_RESET_B_c_1313_n N_A_2523_397#_c_2582_n 0.0223542f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1124 N_RESET_B_c_1316_n N_A_2523_397#_c_2582_n 0.0103857f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1125 N_RESET_B_c_1306_n N_A_2523_397#_c_2583_n 0.00444842f $X=13.52 $Y=2.1
+ $X2=0 $Y2=0
cc_1126 N_RESET_B_c_1306_n N_A_2523_397#_c_2584_n 0.009582f $X=13.52 $Y=2.1
+ $X2=0 $Y2=0
cc_1127 N_RESET_B_c_1296_n N_A_2523_397#_c_2584_n 0.00342537f $X=13.52 $Y=1.7
+ $X2=0 $Y2=0
cc_1128 N_RESET_B_c_1313_n N_A_2523_397#_c_2584_n 0.00894877f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1129 N_RESET_B_c_1315_n N_A_2523_397#_c_2584_n 0.00221939f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1130 N_RESET_B_c_1316_n N_A_2523_397#_c_2584_n 0.0430878f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1131 N_RESET_B_c_1320_n N_A_2523_397#_c_2584_n 0.00666923f $X=13.88 $Y=2.265
+ $X2=0 $Y2=0
cc_1132 N_RESET_B_c_1296_n N_A_2523_397#_c_2585_n 0.00558927f $X=13.52 $Y=1.7
+ $X2=0 $Y2=0
cc_1133 N_RESET_B_c_1315_n N_A_2523_397#_c_2587_n 0.0062291f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1134 N_RESET_B_c_1316_n N_A_2523_397#_c_2587_n 0.0211152f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1135 N_RESET_B_c_1289_n N_VGND_c_2682_n 0.0113547f $X=3.915 $Y=0.18 $X2=0
+ $Y2=0
cc_1136 N_RESET_B_c_1288_n N_VGND_c_2683_n 0.011854f $X=6.755 $Y=0.18 $X2=0
+ $Y2=0
cc_1137 N_RESET_B_c_1289_n N_VGND_c_2688_n 0.0691484f $X=3.915 $Y=0.18 $X2=0
+ $Y2=0
cc_1138 N_RESET_B_c_1288_n N_VGND_c_2698_n 0.0785957f $X=6.755 $Y=0.18 $X2=0
+ $Y2=0
cc_1139 N_RESET_B_c_1289_n N_VGND_c_2698_n 0.00640313f $X=3.915 $Y=0.18 $X2=0
+ $Y2=0
cc_1140 N_RESET_B_c_1293_n N_noxref_39_c_2889_n 0.00368504f $X=4.03 $Y=1.625
+ $X2=0 $Y2=0
cc_1141 N_RESET_B_c_1292_n N_noxref_39_c_2891_n 0.00200577f $X=3.94 $Y=0.9 $X2=0
+ $Y2=0
cc_1142 N_RESET_B_c_1293_n N_noxref_39_c_2891_n 0.0018102f $X=4.03 $Y=1.625
+ $X2=0 $Y2=0
cc_1143 N_RESET_B_M1041_g N_noxref_39_c_2892_n 0.00425508f $X=3.84 $Y=0.54 $X2=0
+ $Y2=0
cc_1144 N_RESET_B_c_1292_n N_noxref_39_c_2892_n 0.00425668f $X=3.94 $Y=0.9 $X2=0
+ $Y2=0
cc_1145 N_RESET_B_M1041_g N_noxref_39_c_2894_n 0.0139499f $X=3.84 $Y=0.54 $X2=0
+ $Y2=0
cc_1146 N_RESET_B_c_1288_n N_noxref_39_c_2894_n 0.00483809f $X=6.755 $Y=0.18
+ $X2=0 $Y2=0
cc_1147 N_RESET_B_c_1292_n N_noxref_39_c_2894_n 0.0131707f $X=3.94 $Y=0.9 $X2=0
+ $Y2=0
cc_1148 N_RESET_B_c_1288_n N_A_824_219#_c_2941_n 0.00241014f $X=6.755 $Y=0.18
+ $X2=0 $Y2=0
cc_1149 N_RESET_B_c_1288_n N_A_824_219#_c_2943_n 0.00349538f $X=6.755 $Y=0.18
+ $X2=0 $Y2=0
cc_1150 N_RESET_B_c_1292_n N_A_824_219#_c_2943_n 0.00253041f $X=3.94 $Y=0.9
+ $X2=0 $Y2=0
cc_1151 N_RESET_B_c_1293_n N_A_824_219#_c_2943_n 0.00752376f $X=4.03 $Y=1.625
+ $X2=0 $Y2=0
cc_1152 N_RESET_B_c_1297_n N_A_824_219#_c_2943_n 6.921e-19 $X=4.03 $Y=1.79 $X2=0
+ $Y2=0
cc_1153 N_RESET_B_c_1298_n N_A_824_219#_c_2943_n 0.00757334f $X=4.03 $Y=1.79
+ $X2=0 $Y2=0
cc_1154 N_A_911_219#_c_1566_n N_VPWR_M1003_d 6.46074e-19 $X=6.455 $Y=2.7 $X2=0
+ $Y2=0
cc_1155 N_A_911_219#_c_1619_n N_VPWR_M1003_d 0.00397447f $X=7.21 $Y=2.785 $X2=0
+ $Y2=0
cc_1156 N_A_911_219#_c_1653_n N_VPWR_M1003_d 0.00521329f $X=6.54 $Y=2.785 $X2=0
+ $Y2=0
cc_1157 N_A_911_219#_c_1565_n N_VPWR_c_2194_n 0.0194564f $X=6.37 $Y=2.47 $X2=0
+ $Y2=0
cc_1158 N_A_911_219#_c_1653_n N_VPWR_c_2194_n 0.0110159f $X=6.54 $Y=2.785 $X2=0
+ $Y2=0
cc_1159 N_A_911_219#_M1009_g N_VPWR_c_2195_n 0.0091923f $X=8.65 $Y=2.295 $X2=0
+ $Y2=0
cc_1160 N_A_911_219#_M1009_g N_VPWR_c_2200_n 0.00385726f $X=8.65 $Y=2.295 $X2=0
+ $Y2=0
cc_1161 N_A_911_219#_c_1619_n N_VPWR_c_2200_n 0.0158767f $X=7.21 $Y=2.785 $X2=0
+ $Y2=0
cc_1162 N_A_911_219#_c_1653_n N_VPWR_c_2200_n 0.00492112f $X=6.54 $Y=2.785 $X2=0
+ $Y2=0
cc_1163 N_A_911_219#_c_1622_n N_VPWR_c_2200_n 0.0139044f $X=7.335 $Y=2.785 $X2=0
+ $Y2=0
cc_1164 N_A_911_219#_c_1560_n N_VPWR_c_2206_n 0.00611391f $X=4.81 $Y=2.665 $X2=0
+ $Y2=0
cc_1165 N_A_911_219#_M1049_d N_VPWR_c_2191_n 0.00445132f $X=7.235 $Y=2.675 $X2=0
+ $Y2=0
cc_1166 N_A_911_219#_M1009_g N_VPWR_c_2191_n 0.00426651f $X=8.65 $Y=2.295 $X2=0
+ $Y2=0
cc_1167 N_A_911_219#_c_1560_n N_VPWR_c_2191_n 0.00650468f $X=4.81 $Y=2.665 $X2=0
+ $Y2=0
cc_1168 N_A_911_219#_c_1561_n N_VPWR_c_2191_n 0.0213833f $X=5.505 $Y=2.47 $X2=0
+ $Y2=0
cc_1169 N_A_911_219#_c_1565_n N_VPWR_c_2191_n 0.0129253f $X=6.37 $Y=2.47 $X2=0
+ $Y2=0
cc_1170 N_A_911_219#_c_1619_n N_VPWR_c_2191_n 0.0205282f $X=7.21 $Y=2.785 $X2=0
+ $Y2=0
cc_1171 N_A_911_219#_c_1653_n N_VPWR_c_2191_n 0.00575654f $X=6.54 $Y=2.785 $X2=0
+ $Y2=0
cc_1172 N_A_911_219#_c_1567_n N_VPWR_c_2191_n 0.00707863f $X=5.59 $Y=2.47 $X2=0
+ $Y2=0
cc_1173 N_A_911_219#_c_1622_n N_VPWR_c_2191_n 0.00932251f $X=7.335 $Y=2.785
+ $X2=0 $Y2=0
cc_1174 N_A_911_219#_c_1551_n N_A_342_261#_M1015_d 0.00990086f $X=5.505 $Y=1.32
+ $X2=0 $Y2=0
cc_1175 N_A_911_219#_c_1560_n N_A_342_261#_c_2422_n 0.0154734f $X=4.81 $Y=2.665
+ $X2=0 $Y2=0
cc_1176 N_A_911_219#_c_1560_n N_A_342_261#_c_2413_n 0.0101975f $X=4.81 $Y=2.665
+ $X2=0 $Y2=0
cc_1177 N_A_911_219#_c_1562_n N_A_342_261#_c_2413_n 0.0124128f $X=4.905 $Y=2.47
+ $X2=0 $Y2=0
cc_1178 N_A_911_219#_c_1551_n N_A_342_261#_c_2414_n 0.00470077f $X=5.505 $Y=1.32
+ $X2=0 $Y2=0
cc_1179 N_A_911_219#_c_1561_n N_A_342_261#_c_2414_n 0.0240572f $X=5.505 $Y=2.47
+ $X2=0 $Y2=0
cc_1180 N_A_911_219#_c_1562_n N_A_342_261#_c_2414_n 0.0111236f $X=4.905 $Y=2.47
+ $X2=0 $Y2=0
cc_1181 N_A_911_219#_c_1553_n N_A_342_261#_c_2414_n 0.0125335f $X=5.59 $Y=2.385
+ $X2=0 $Y2=0
cc_1182 N_A_911_219#_c_1555_n N_A_342_261#_c_2414_n 0.0116283f $X=4.86 $Y=1.385
+ $X2=0 $Y2=0
cc_1183 N_A_911_219#_c_1555_n N_A_342_261#_c_2415_n 5.00719e-19 $X=4.86 $Y=1.385
+ $X2=0 $Y2=0
cc_1184 N_A_911_219#_c_1551_n N_A_342_261#_c_2416_n 0.0191954f $X=5.505 $Y=1.32
+ $X2=0 $Y2=0
cc_1185 N_A_911_219#_c_1553_n N_A_342_261#_c_2416_n 0.0227878f $X=5.59 $Y=2.385
+ $X2=0 $Y2=0
cc_1186 N_A_911_219#_c_1556_n N_A_342_261#_c_2416_n 0.0106375f $X=5.59 $Y=1.63
+ $X2=0 $Y2=0
cc_1187 N_A_911_219#_c_1561_n A_1020_491# 0.00781194f $X=5.505 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_1188 N_A_911_219#_c_1567_n A_1020_491# 0.00296637f $X=5.59 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_1189 N_A_911_219#_c_1619_n A_1375_535# 0.00220461f $X=7.21 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1190 N_A_911_219#_M1021_g N_VGND_c_2684_n 0.00158723f $X=8.62 $Y=0.755 $X2=0
+ $Y2=0
cc_1191 N_A_911_219#_M1000_g N_VGND_c_2694_n 8.5177e-19 $X=8.23 $Y=0.755 $X2=0
+ $Y2=0
cc_1192 N_A_911_219#_M1021_g N_VGND_c_2694_n 0.00311088f $X=8.62 $Y=0.755 $X2=0
+ $Y2=0
cc_1193 N_A_911_219#_M1021_g N_VGND_c_2698_n 0.00367659f $X=8.62 $Y=0.755 $X2=0
+ $Y2=0
cc_1194 N_A_911_219#_c_1555_n N_A_824_219#_c_2941_n 0.0603427f $X=4.86 $Y=1.385
+ $X2=0 $Y2=0
cc_1195 N_A_911_219#_c_1554_n N_A_824_219#_c_2942_n 0.011992f $X=7.48 $Y=1.63
+ $X2=0 $Y2=0
cc_1196 N_A_911_219#_c_1551_n N_A_824_219#_c_2944_n 0.0171057f $X=5.505 $Y=1.32
+ $X2=0 $Y2=0
cc_1197 N_A_911_219#_c_1554_n N_A_824_219#_c_2944_n 0.00358109f $X=7.48 $Y=1.63
+ $X2=0 $Y2=0
cc_1198 N_A_2388_115#_c_1738_n N_A_2168_439#_M1037_g 0.00766138f $X=13.14
+ $Y=2.53 $X2=0 $Y2=0
cc_1199 N_A_2388_115#_c_1740_n N_A_2168_439#_M1037_g 9.42915e-19 $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1200 N_A_2388_115#_c_1741_n N_A_2168_439#_M1037_g 0.00661606f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1201 N_A_2388_115#_c_1735_n N_A_2168_439#_M1037_g 0.00452932f $X=12.275
+ $Y=2.185 $X2=0 $Y2=0
cc_1202 N_A_2388_115#_c_1746_n N_A_2168_439#_c_1839_n 0.0120541f $X=13.89
+ $Y=0.975 $X2=0 $Y2=0
cc_1203 N_A_2388_115#_c_1734_n N_A_2168_439#_c_1839_n 0.00923711f $X=14.055
+ $Y=0.87 $X2=0 $Y2=0
cc_1204 N_A_2388_115#_c_1746_n N_A_2168_439#_c_1840_n 0.00162939f $X=13.89
+ $Y=0.975 $X2=0 $Y2=0
cc_1205 N_A_2388_115#_c_1734_n N_A_2168_439#_c_1840_n 0.00546738f $X=14.055
+ $Y=0.87 $X2=0 $Y2=0
cc_1206 N_A_2388_115#_c_1729_n N_A_2168_439#_c_1855_n 0.00856388f $X=12.015
+ $Y=1.235 $X2=0 $Y2=0
cc_1207 N_A_2388_115#_M1018_g N_A_2168_439#_c_1874_n 4.45208e-19 $X=12.365
+ $Y=2.885 $X2=0 $Y2=0
cc_1208 N_A_2388_115#_c_1740_n N_A_2168_439#_c_1874_n 0.0131871f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1209 N_A_2388_115#_c_1741_n N_A_2168_439#_c_1874_n 0.00184515f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1210 N_A_2388_115#_c_1729_n N_A_2168_439#_c_1856_n 0.0098168f $X=12.015
+ $Y=1.235 $X2=0 $Y2=0
cc_1211 N_A_2388_115#_c_1730_n N_A_2168_439#_c_1856_n 0.0242019f $X=12.305
+ $Y=1.4 $X2=0 $Y2=0
cc_1212 N_A_2388_115#_c_1732_n N_A_2168_439#_c_1856_n 0.00960491f $X=12.47
+ $Y=1.135 $X2=0 $Y2=0
cc_1213 N_A_2388_115#_c_1736_n N_A_2168_439#_c_1856_n 0.0157277f $X=12.185
+ $Y=1.4 $X2=0 $Y2=0
cc_1214 N_A_2388_115#_c_1740_n N_A_2168_439#_c_1876_n 0.0163662f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1215 N_A_2388_115#_c_1735_n N_A_2168_439#_c_1876_n 0.0134788f $X=12.275
+ $Y=2.185 $X2=0 $Y2=0
cc_1216 N_A_2388_115#_c_1730_n N_A_2168_439#_c_1877_n 0.0241017f $X=12.305
+ $Y=1.4 $X2=0 $Y2=0
cc_1217 N_A_2388_115#_c_1738_n N_A_2168_439#_c_1877_n 0.00341922f $X=13.14
+ $Y=2.53 $X2=0 $Y2=0
cc_1218 N_A_2388_115#_c_1731_n N_A_2168_439#_c_1877_n 0.00757017f $X=12.69
+ $Y=1.135 $X2=0 $Y2=0
cc_1219 N_A_2388_115#_c_1740_n N_A_2168_439#_c_1877_n 0.0128444f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1220 N_A_2388_115#_c_1741_n N_A_2168_439#_c_1877_n 9.63138e-19 $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1221 N_A_2388_115#_c_1733_n N_A_2168_439#_c_1877_n 0.00103775f $X=12.775
+ $Y=0.975 $X2=0 $Y2=0
cc_1222 N_A_2388_115#_c_1735_n N_A_2168_439#_c_1877_n 0.0145274f $X=12.275
+ $Y=2.185 $X2=0 $Y2=0
cc_1223 N_A_2388_115#_c_1736_n N_A_2168_439#_c_1877_n 0.0058871f $X=12.185
+ $Y=1.4 $X2=0 $Y2=0
cc_1224 N_A_2388_115#_c_1735_n N_A_2168_439#_c_1938_n 9.58794e-19 $X=12.275
+ $Y=2.185 $X2=0 $Y2=0
cc_1225 N_A_2388_115#_c_1746_n N_A_2168_439#_c_1857_n 9.57564e-19 $X=13.89
+ $Y=0.975 $X2=0 $Y2=0
cc_1226 N_A_2388_115#_c_1733_n N_A_2168_439#_c_1857_n 8.05223e-19 $X=12.775
+ $Y=0.975 $X2=0 $Y2=0
cc_1227 N_A_2388_115#_c_1735_n N_A_2168_439#_c_1857_n 0.0068951f $X=12.275
+ $Y=2.185 $X2=0 $Y2=0
cc_1228 N_A_2388_115#_c_1736_n N_A_2168_439#_c_1857_n 0.00357567f $X=12.185
+ $Y=1.4 $X2=0 $Y2=0
cc_1229 N_A_2388_115#_c_1730_n N_A_2168_439#_c_1858_n 0.0101082f $X=12.305
+ $Y=1.4 $X2=0 $Y2=0
cc_1230 N_A_2388_115#_c_1746_n N_A_2168_439#_c_1858_n 0.00940644f $X=13.89
+ $Y=0.975 $X2=0 $Y2=0
cc_1231 N_A_2388_115#_c_1733_n N_A_2168_439#_c_1858_n 0.0116024f $X=12.775
+ $Y=0.975 $X2=0 $Y2=0
cc_1232 N_A_2388_115#_c_1736_n N_A_2168_439#_c_1858_n 0.0024195f $X=12.185
+ $Y=1.4 $X2=0 $Y2=0
cc_1233 N_A_2388_115#_c_1734_n N_A_2168_439#_c_1861_n 0.0139106f $X=14.055
+ $Y=0.87 $X2=0 $Y2=0
cc_1234 N_A_2388_115#_c_1746_n N_A_2168_439#_c_1862_n 0.0315956f $X=13.89
+ $Y=0.975 $X2=0 $Y2=0
cc_1235 N_A_2388_115#_c_1734_n N_A_2168_439#_c_1862_n 0.00782921f $X=14.055
+ $Y=0.87 $X2=0 $Y2=0
cc_1236 N_A_2388_115#_c_1734_n N_A_2168_439#_c_1863_n 0.00633107f $X=14.055
+ $Y=0.87 $X2=0 $Y2=0
cc_1237 N_A_2388_115#_M1018_g N_VPWR_c_2196_n 0.010302f $X=12.365 $Y=2.885 $X2=0
+ $Y2=0
cc_1238 N_A_2388_115#_c_1738_n N_VPWR_c_2196_n 0.0227507f $X=13.14 $Y=2.53 $X2=0
+ $Y2=0
cc_1239 N_A_2388_115#_c_1739_n N_VPWR_c_2196_n 0.0124053f $X=13.305 $Y=2.8 $X2=0
+ $Y2=0
cc_1240 N_A_2388_115#_c_1739_n N_VPWR_c_2197_n 0.010811f $X=13.305 $Y=2.8 $X2=0
+ $Y2=0
cc_1241 N_A_2388_115#_M1018_g N_VPWR_c_2207_n 0.00424635f $X=12.365 $Y=2.885
+ $X2=0 $Y2=0
cc_1242 N_A_2388_115#_c_1738_n N_VPWR_c_2207_n 0.00118595f $X=13.14 $Y=2.53
+ $X2=0 $Y2=0
cc_1243 N_A_2388_115#_c_1740_n N_VPWR_c_2207_n 0.00144139f $X=12.275 $Y=2.35
+ $X2=0 $Y2=0
cc_1244 N_A_2388_115#_c_1738_n N_VPWR_c_2208_n 0.00485687f $X=13.14 $Y=2.53
+ $X2=0 $Y2=0
cc_1245 N_A_2388_115#_c_1739_n N_VPWR_c_2208_n 0.0180077f $X=13.305 $Y=2.8 $X2=0
+ $Y2=0
cc_1246 N_A_2388_115#_M1018_g N_VPWR_c_2191_n 0.0085805f $X=12.365 $Y=2.885
+ $X2=0 $Y2=0
cc_1247 N_A_2388_115#_c_1738_n N_VPWR_c_2191_n 0.01182f $X=13.14 $Y=2.53 $X2=0
+ $Y2=0
cc_1248 N_A_2388_115#_c_1739_n N_VPWR_c_2191_n 0.0122962f $X=13.305 $Y=2.8 $X2=0
+ $Y2=0
cc_1249 N_A_2388_115#_c_1740_n N_VPWR_c_2191_n 0.00263247f $X=12.275 $Y=2.35
+ $X2=0 $Y2=0
cc_1250 N_A_2388_115#_M1018_g N_A_2081_439#_c_2554_n 0.0034909f $X=12.365
+ $Y=2.885 $X2=0 $Y2=0
cc_1251 N_A_2388_115#_c_1740_n N_A_2081_439#_c_2554_n 0.0101956f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1252 N_A_2388_115#_c_1741_n N_A_2081_439#_c_2554_n 0.00190976f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1253 N_A_2388_115#_M1037_d N_A_2523_397#_c_2582_n 0.00496606f $X=13.05
+ $Y=1.985 $X2=0 $Y2=0
cc_1254 N_A_2388_115#_c_1738_n N_A_2523_397#_c_2582_n 0.0455287f $X=13.14
+ $Y=2.53 $X2=0 $Y2=0
cc_1255 N_A_2388_115#_c_1740_n N_A_2523_397#_c_2582_n 0.00630305f $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1256 N_A_2388_115#_c_1741_n N_A_2523_397#_c_2582_n 7.61571e-19 $X=12.275
+ $Y=2.35 $X2=0 $Y2=0
cc_1257 N_A_2388_115#_c_1735_n N_A_2523_397#_c_2582_n 0.00107199f $X=12.275
+ $Y=2.185 $X2=0 $Y2=0
cc_1258 N_A_2388_115#_M1037_d N_A_2523_397#_c_2583_n 0.00147792f $X=13.05
+ $Y=1.985 $X2=0 $Y2=0
cc_1259 N_A_2388_115#_c_1738_n N_A_2523_397#_c_2584_n 0.00125731f $X=13.14
+ $Y=2.53 $X2=0 $Y2=0
cc_1260 N_A_2388_115#_c_1731_n N_VGND_M1011_d 0.00773021f $X=12.69 $Y=1.135
+ $X2=0 $Y2=0
cc_1261 N_A_2388_115#_c_1732_n N_VGND_M1011_d 0.00481048f $X=12.47 $Y=1.135
+ $X2=0 $Y2=0
cc_1262 N_A_2388_115#_c_1746_n N_VGND_M1011_d 0.0118757f $X=13.89 $Y=0.975 $X2=0
+ $Y2=0
cc_1263 N_A_2388_115#_c_1733_n N_VGND_M1011_d 0.00834166f $X=12.775 $Y=0.975
+ $X2=0 $Y2=0
cc_1264 N_A_2388_115#_c_1729_n N_VGND_c_2685_n 0.00633384f $X=12.015 $Y=1.235
+ $X2=0 $Y2=0
cc_1265 N_A_2388_115#_c_1731_n N_VGND_c_2685_n 0.00300524f $X=12.69 $Y=1.135
+ $X2=0 $Y2=0
cc_1266 N_A_2388_115#_c_1732_n N_VGND_c_2685_n 0.0244573f $X=12.47 $Y=1.135
+ $X2=0 $Y2=0
cc_1267 N_A_2388_115#_c_1736_n N_VGND_c_2685_n 0.00148018f $X=12.185 $Y=1.4
+ $X2=0 $Y2=0
cc_1268 N_A_2388_115#_c_1729_n N_VGND_c_2698_n 8.38936e-19 $X=12.015 $Y=1.235
+ $X2=0 $Y2=0
cc_1269 N_A_2388_115#_c_1746_n A_2682_141# 0.00356853f $X=13.89 $Y=0.975
+ $X2=-0.19 $Y2=-0.245
cc_1270 N_A_2168_439#_c_1860_n N_CLK_M1026_g 0.0181798f $X=16.015 $Y=0.975 $X2=0
+ $Y2=0
cc_1271 N_A_2168_439#_M1046_g N_CLK_M1027_g 0.0371463f $X=16.09 $Y=0.655 $X2=0
+ $Y2=0
cc_1272 N_A_2168_439#_c_1860_n N_CLK_M1027_g 0.0142078f $X=16.015 $Y=0.975 $X2=0
+ $Y2=0
cc_1273 N_A_2168_439#_c_1865_n N_CLK_M1027_g 0.00147457f $X=16.18 $Y=1.255 $X2=0
+ $Y2=0
cc_1274 N_A_2168_439#_M1033_g N_CLK_M1055_g 0.0198497f $X=16.09 $Y=2.415 $X2=0
+ $Y2=0
cc_1275 N_A_2168_439#_M1033_g N_CLK_c_2085_n 0.00329784f $X=16.09 $Y=2.415 $X2=0
+ $Y2=0
cc_1276 N_A_2168_439#_c_1860_n N_CLK_c_2085_n 0.0168106f $X=16.015 $Y=0.975
+ $X2=0 $Y2=0
cc_1277 N_A_2168_439#_c_1864_n N_CLK_c_2085_n 0.0157409f $X=16.18 $Y=1.42 $X2=0
+ $Y2=0
cc_1278 N_A_2168_439#_c_1867_n N_CLK_c_2085_n 0.00147094f $X=16.525 $Y=1.42
+ $X2=0 $Y2=0
cc_1279 N_A_2168_439#_c_1864_n N_CLK_c_2086_n 0.00119764f $X=16.18 $Y=1.42 $X2=0
+ $Y2=0
cc_1280 N_A_2168_439#_c_1867_n N_CLK_c_2086_n 0.0172607f $X=16.525 $Y=1.42 $X2=0
+ $Y2=0
cc_1281 N_A_2168_439#_M1001_g N_A_3416_137#_M1012_g 0.0154566f $X=17.8 $Y=0.895
+ $X2=0 $Y2=0
cc_1282 N_A_2168_439#_M1039_g N_A_3416_137#_M1053_g 0.0166304f $X=17.8 $Y=2.155
+ $X2=0 $Y2=0
cc_1283 N_A_2168_439#_M1031_g N_A_3416_137#_c_2133_n 0.00169897f $X=16.45
+ $Y=0.655 $X2=0 $Y2=0
cc_1284 N_A_2168_439#_c_1847_n N_A_3416_137#_c_2133_n 0.00717458f $X=17.365
+ $Y=1.33 $X2=0 $Y2=0
cc_1285 N_A_2168_439#_M1022_g N_A_3416_137#_c_2133_n 0.0148544f $X=17.44
+ $Y=0.895 $X2=0 $Y2=0
cc_1286 N_A_2168_439#_M1001_g N_A_3416_137#_c_2133_n 0.00197812f $X=17.8
+ $Y=0.895 $X2=0 $Y2=0
cc_1287 N_A_2168_439#_c_1853_n N_A_3416_137#_c_2133_n 0.00230932f $X=17.44
+ $Y=1.33 $X2=0 $Y2=0
cc_1288 N_A_2168_439#_M1007_g N_A_3416_137#_c_2134_n 0.0023197f $X=16.45
+ $Y=2.415 $X2=0 $Y2=0
cc_1289 N_A_2168_439#_M1034_g N_A_3416_137#_c_2134_n 0.0201599f $X=17.44
+ $Y=2.155 $X2=0 $Y2=0
cc_1290 N_A_2168_439#_M1039_g N_A_3416_137#_c_2134_n 0.0028674f $X=17.8 $Y=2.155
+ $X2=0 $Y2=0
cc_1291 N_A_2168_439#_M1034_g N_A_3416_137#_c_2135_n 0.0106629f $X=17.44
+ $Y=2.155 $X2=0 $Y2=0
cc_1292 N_A_2168_439#_c_1850_n N_A_3416_137#_c_2135_n 0.0122117f $X=17.725
+ $Y=1.33 $X2=0 $Y2=0
cc_1293 N_A_2168_439#_M1039_g N_A_3416_137#_c_2135_n 0.0157309f $X=17.8 $Y=2.155
+ $X2=0 $Y2=0
cc_1294 N_A_2168_439#_c_1853_n N_A_3416_137#_c_2135_n 0.00707746f $X=17.44
+ $Y=1.33 $X2=0 $Y2=0
cc_1295 N_A_2168_439#_c_1854_n N_A_3416_137#_c_2135_n 0.0100329f $X=17.8 $Y=1.33
+ $X2=0 $Y2=0
cc_1296 N_A_2168_439#_c_1847_n N_A_3416_137#_c_2136_n 0.00974531f $X=17.365
+ $Y=1.33 $X2=0 $Y2=0
cc_1297 N_A_2168_439#_M1034_g N_A_3416_137#_c_2136_n 0.00516568f $X=17.44
+ $Y=2.155 $X2=0 $Y2=0
cc_1298 N_A_2168_439#_c_1853_n N_A_3416_137#_c_2136_n 2.35411e-19 $X=17.44
+ $Y=1.33 $X2=0 $Y2=0
cc_1299 N_A_2168_439#_c_1854_n N_A_3416_137#_c_2137_n 0.0103406f $X=17.8 $Y=1.33
+ $X2=0 $Y2=0
cc_1300 N_A_2168_439#_M1019_g N_VPWR_c_2197_n 0.00272121f $X=14.31 $Y=2.8 $X2=0
+ $Y2=0
cc_1301 N_A_2168_439#_M1033_g N_VPWR_c_2198_n 0.0223586f $X=16.09 $Y=2.415 $X2=0
+ $Y2=0
cc_1302 N_A_2168_439#_M1007_g N_VPWR_c_2198_n 0.00386758f $X=16.45 $Y=2.415
+ $X2=0 $Y2=0
cc_1303 N_A_2168_439#_c_1864_n N_VPWR_c_2198_n 0.00102733f $X=16.18 $Y=1.42
+ $X2=0 $Y2=0
cc_1304 N_A_2168_439#_M1039_g N_VPWR_c_2199_n 0.0124152f $X=17.8 $Y=2.155 $X2=0
+ $Y2=0
cc_1305 N_A_2168_439#_M1019_g N_VPWR_c_2202_n 0.00473334f $X=14.31 $Y=2.8 $X2=0
+ $Y2=0
cc_1306 N_A_2168_439#_M1033_g N_VPWR_c_2209_n 0.00445056f $X=16.09 $Y=2.415
+ $X2=0 $Y2=0
cc_1307 N_A_2168_439#_M1007_g N_VPWR_c_2209_n 0.00502664f $X=16.45 $Y=2.415
+ $X2=0 $Y2=0
cc_1308 N_A_2168_439#_M1034_g N_VPWR_c_2209_n 0.00312414f $X=17.44 $Y=2.155
+ $X2=0 $Y2=0
cc_1309 N_A_2168_439#_M1039_g N_VPWR_c_2209_n 0.00312414f $X=17.8 $Y=2.155 $X2=0
+ $Y2=0
cc_1310 N_A_2168_439#_M1019_g N_VPWR_c_2191_n 0.00835478f $X=14.31 $Y=2.8 $X2=0
+ $Y2=0
cc_1311 N_A_2168_439#_M1033_g N_VPWR_c_2191_n 0.00796275f $X=16.09 $Y=2.415
+ $X2=0 $Y2=0
cc_1312 N_A_2168_439#_M1007_g N_VPWR_c_2191_n 0.010303f $X=16.45 $Y=2.415 $X2=0
+ $Y2=0
cc_1313 N_A_2168_439#_M1034_g N_VPWR_c_2191_n 0.00410284f $X=17.44 $Y=2.155
+ $X2=0 $Y2=0
cc_1314 N_A_2168_439#_M1039_g N_VPWR_c_2191_n 0.00410284f $X=17.8 $Y=2.155 $X2=0
+ $Y2=0
cc_1315 N_A_2168_439#_c_1879_n N_A_2081_439#_c_2552_n 0.0184558f $X=11.26
+ $Y=2.57 $X2=0 $Y2=0
cc_1316 N_A_2168_439#_c_1874_n N_A_2081_439#_c_2555_n 0.0255271f $X=11.79
+ $Y=2.51 $X2=0 $Y2=0
cc_1317 N_A_2168_439#_c_1879_n N_A_2081_439#_c_2555_n 0.0195211f $X=11.26
+ $Y=2.57 $X2=0 $Y2=0
cc_1318 N_A_2168_439#_M1037_g N_A_2523_397#_c_2582_n 0.0087186f $X=12.975
+ $Y=2.195 $X2=0 $Y2=0
cc_1319 N_A_2168_439#_c_1876_n N_A_2523_397#_c_2582_n 0.00296012f $X=11.875
+ $Y=2.425 $X2=0 $Y2=0
cc_1320 N_A_2168_439#_c_1877_n N_A_2523_397#_c_2582_n 0.0296143f $X=12.72
+ $Y=1.83 $X2=0 $Y2=0
cc_1321 N_A_2168_439#_c_1857_n N_A_2523_397#_c_2582_n 8.89472e-19 $X=12.885
+ $Y=1.66 $X2=0 $Y2=0
cc_1322 N_A_2168_439#_c_1862_n N_A_2523_397#_c_2582_n 0.00500548f $X=14.055
+ $Y=1.405 $X2=0 $Y2=0
cc_1323 N_A_2168_439#_M1037_g N_A_2523_397#_c_2583_n 0.00374223f $X=12.975
+ $Y=2.195 $X2=0 $Y2=0
cc_1324 N_A_2168_439#_M1019_g N_A_2523_397#_c_2584_n 0.0158993f $X=14.31 $Y=2.8
+ $X2=0 $Y2=0
cc_1325 N_A_2168_439#_c_1862_n N_A_2523_397#_c_2584_n 0.0777081f $X=14.055
+ $Y=1.405 $X2=0 $Y2=0
cc_1326 N_A_2168_439#_c_1866_n N_A_2523_397#_c_2584_n 0.00402216f $X=14.22
+ $Y=1.31 $X2=0 $Y2=0
cc_1327 N_A_2168_439#_c_1877_n N_A_2523_397#_c_2585_n 0.0140445f $X=12.72
+ $Y=1.83 $X2=0 $Y2=0
cc_1328 N_A_2168_439#_c_1857_n N_A_2523_397#_c_2585_n 7.11062e-19 $X=12.885
+ $Y=1.66 $X2=0 $Y2=0
cc_1329 N_A_2168_439#_c_1862_n N_A_2523_397#_c_2585_n 0.0123289f $X=14.055
+ $Y=1.405 $X2=0 $Y2=0
cc_1330 N_A_2168_439#_M1019_g N_A_2523_397#_c_2586_n 0.00510283f $X=14.31 $Y=2.8
+ $X2=0 $Y2=0
cc_1331 N_A_2168_439#_M1019_g N_A_2523_397#_c_2587_n 0.0210129f $X=14.31 $Y=2.8
+ $X2=0 $Y2=0
cc_1332 N_A_2168_439#_M1033_g N_Q_N_c_2634_n 0.00398253f $X=16.09 $Y=2.415 $X2=0
+ $Y2=0
cc_1333 N_A_2168_439#_M1007_g N_Q_N_c_2634_n 0.00448422f $X=16.45 $Y=2.415 $X2=0
+ $Y2=0
cc_1334 N_A_2168_439#_c_1847_n N_Q_N_c_2634_n 0.00151161f $X=17.365 $Y=1.33
+ $X2=0 $Y2=0
cc_1335 N_A_2168_439#_M1007_g N_Q_N_c_2635_n 0.0225194f $X=16.45 $Y=2.415 $X2=0
+ $Y2=0
cc_1336 N_A_2168_439#_M1034_g N_Q_N_c_2635_n 0.00278664f $X=17.44 $Y=2.155 $X2=0
+ $Y2=0
cc_1337 N_A_2168_439#_M1031_g N_Q_N_c_2631_n 0.0030176f $X=16.45 $Y=0.655 $X2=0
+ $Y2=0
cc_1338 N_A_2168_439#_c_1847_n N_Q_N_c_2631_n 0.0157433f $X=17.365 $Y=1.33 $X2=0
+ $Y2=0
cc_1339 N_A_2168_439#_M1034_g N_Q_N_c_2631_n 0.00281971f $X=17.44 $Y=2.155 $X2=0
+ $Y2=0
cc_1340 N_A_2168_439#_c_1864_n N_Q_N_c_2631_n 0.0150719f $X=16.18 $Y=1.42 $X2=0
+ $Y2=0
cc_1341 N_A_2168_439#_c_1865_n N_Q_N_c_2631_n 0.00476004f $X=16.18 $Y=1.255
+ $X2=0 $Y2=0
cc_1342 N_A_2168_439#_c_1867_n N_Q_N_c_2631_n 0.00951916f $X=16.525 $Y=1.42
+ $X2=0 $Y2=0
cc_1343 N_A_2168_439#_M1046_g N_Q_N_c_2632_n 0.00233112f $X=16.09 $Y=0.655 $X2=0
+ $Y2=0
cc_1344 N_A_2168_439#_M1031_g N_Q_N_c_2632_n 0.014553f $X=16.45 $Y=0.655 $X2=0
+ $Y2=0
cc_1345 N_A_2168_439#_M1022_g N_Q_N_c_2632_n 0.00430775f $X=17.44 $Y=0.895 $X2=0
+ $Y2=0
cc_1346 N_A_2168_439#_M1046_g Q_N 2.05581e-19 $X=16.09 $Y=0.655 $X2=0 $Y2=0
cc_1347 N_A_2168_439#_M1031_g Q_N 0.00709729f $X=16.45 $Y=0.655 $X2=0 $Y2=0
cc_1348 N_A_2168_439#_c_1847_n Q_N 0.00183f $X=17.365 $Y=1.33 $X2=0 $Y2=0
cc_1349 N_A_2168_439#_c_1860_n N_VGND_M1027_d 0.00814128f $X=16.015 $Y=0.975
+ $X2=0 $Y2=0
cc_1350 N_A_2168_439#_c_1855_n N_VGND_c_2685_n 0.0201156f $X=11.79 $Y=0.74 $X2=0
+ $Y2=0
cc_1351 N_A_2168_439#_M1046_g N_VGND_c_2686_n 0.0133134f $X=16.09 $Y=0.655 $X2=0
+ $Y2=0
cc_1352 N_A_2168_439#_M1031_g N_VGND_c_2686_n 0.00245447f $X=16.45 $Y=0.655
+ $X2=0 $Y2=0
cc_1353 N_A_2168_439#_c_1860_n N_VGND_c_2686_n 0.0166287f $X=16.015 $Y=0.975
+ $X2=0 $Y2=0
cc_1354 N_A_2168_439#_M1001_g N_VGND_c_2687_n 0.0093704f $X=17.8 $Y=0.895 $X2=0
+ $Y2=0
cc_1355 N_A_2168_439#_c_1855_n N_VGND_c_2695_n 0.0178642f $X=11.79 $Y=0.74 $X2=0
+ $Y2=0
cc_1356 N_A_2168_439#_M1046_g N_VGND_c_2696_n 0.00486043f $X=16.09 $Y=0.655
+ $X2=0 $Y2=0
cc_1357 N_A_2168_439#_M1031_g N_VGND_c_2696_n 0.00466554f $X=16.45 $Y=0.655
+ $X2=0 $Y2=0
cc_1358 N_A_2168_439#_M1022_g N_VGND_c_2696_n 0.00371502f $X=17.44 $Y=0.895
+ $X2=0 $Y2=0
cc_1359 N_A_2168_439#_M1001_g N_VGND_c_2696_n 0.00385058f $X=17.8 $Y=0.895 $X2=0
+ $Y2=0
cc_1360 N_A_2168_439#_M1046_g N_VGND_c_2698_n 0.00814425f $X=16.09 $Y=0.655
+ $X2=0 $Y2=0
cc_1361 N_A_2168_439#_M1031_g N_VGND_c_2698_n 0.00907206f $X=16.45 $Y=0.655
+ $X2=0 $Y2=0
cc_1362 N_A_2168_439#_M1022_g N_VGND_c_2698_n 0.00453162f $X=17.44 $Y=0.895
+ $X2=0 $Y2=0
cc_1363 N_A_2168_439#_M1001_g N_VGND_c_2698_n 0.00453162f $X=17.8 $Y=0.895 $X2=0
+ $Y2=0
cc_1364 N_A_2168_439#_c_1855_n N_VGND_c_2698_n 0.0221088f $X=11.79 $Y=0.74 $X2=0
+ $Y2=0
cc_1365 N_A_2168_439#_c_1855_n A_2340_141# 0.00132284f $X=11.79 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_1366 N_A_2168_439#_c_1856_n A_2340_141# 0.00251505f $X=11.875 $Y=1.745
+ $X2=-0.19 $Y2=-0.245
cc_1367 N_A_2168_439#_c_1860_n A_3075_47# 0.00476445f $X=16.015 $Y=0.975
+ $X2=-0.19 $Y2=-0.245
cc_1368 N_CLK_M1052_g N_VPWR_c_2198_n 0.00386758f $X=15.3 $Y=2.415 $X2=0 $Y2=0
cc_1369 N_CLK_M1055_g N_VPWR_c_2198_n 0.0221859f $X=15.66 $Y=2.415 $X2=0 $Y2=0
cc_1370 N_CLK_c_2085_n N_VPWR_c_2198_n 0.00287647f $X=15.595 $Y=1.46 $X2=0 $Y2=0
cc_1371 N_CLK_M1052_g N_VPWR_c_2202_n 0.00502664f $X=15.3 $Y=2.415 $X2=0 $Y2=0
cc_1372 N_CLK_M1055_g N_VPWR_c_2202_n 0.00445056f $X=15.66 $Y=2.415 $X2=0 $Y2=0
cc_1373 N_CLK_M1052_g N_VPWR_c_2191_n 0.010303f $X=15.3 $Y=2.415 $X2=0 $Y2=0
cc_1374 N_CLK_M1055_g N_VPWR_c_2191_n 0.00796275f $X=15.66 $Y=2.415 $X2=0 $Y2=0
cc_1375 N_CLK_M1052_g N_A_2523_397#_c_2584_n 4.28954e-19 $X=15.3 $Y=2.415 $X2=0
+ $Y2=0
cc_1376 N_CLK_M1052_g N_A_2523_397#_c_2587_n 0.00214794f $X=15.3 $Y=2.415 $X2=0
+ $Y2=0
cc_1377 N_CLK_M1026_g N_VGND_c_2686_n 0.0024971f $X=15.3 $Y=0.655 $X2=0 $Y2=0
cc_1378 N_CLK_M1027_g N_VGND_c_2686_n 0.0137365f $X=15.66 $Y=0.655 $X2=0 $Y2=0
cc_1379 N_CLK_M1026_g N_VGND_c_2690_n 0.00547815f $X=15.3 $Y=0.655 $X2=0 $Y2=0
cc_1380 N_CLK_M1027_g N_VGND_c_2690_n 0.00486043f $X=15.66 $Y=0.655 $X2=0 $Y2=0
cc_1381 N_CLK_M1026_g N_VGND_c_2698_n 0.0101319f $X=15.3 $Y=0.655 $X2=0 $Y2=0
cc_1382 N_CLK_M1027_g N_VGND_c_2698_n 0.00814425f $X=15.66 $Y=0.655 $X2=0 $Y2=0
cc_1383 N_A_3416_137#_M1053_g N_VPWR_c_2199_n 0.0300646f $X=18.345 $Y=2.465
+ $X2=0 $Y2=0
cc_1384 N_A_3416_137#_M1058_g N_VPWR_c_2199_n 0.00468428f $X=18.705 $Y=2.465
+ $X2=0 $Y2=0
cc_1385 N_A_3416_137#_c_2134_n N_VPWR_c_2199_n 0.0203141f $X=17.225 $Y=1.98
+ $X2=0 $Y2=0
cc_1386 N_A_3416_137#_c_2135_n N_VPWR_c_2199_n 0.0275493f $X=18.41 $Y=1.47 $X2=0
+ $Y2=0
cc_1387 N_A_3416_137#_c_2137_n N_VPWR_c_2199_n 5.79521e-19 $X=18.705 $Y=1.47
+ $X2=0 $Y2=0
cc_1388 N_A_3416_137#_M1053_g N_VPWR_c_2210_n 0.00486043f $X=18.345 $Y=2.465
+ $X2=0 $Y2=0
cc_1389 N_A_3416_137#_M1058_g N_VPWR_c_2210_n 0.00549284f $X=18.705 $Y=2.465
+ $X2=0 $Y2=0
cc_1390 N_A_3416_137#_M1053_g N_VPWR_c_2191_n 0.00814425f $X=18.345 $Y=2.465
+ $X2=0 $Y2=0
cc_1391 N_A_3416_137#_M1058_g N_VPWR_c_2191_n 0.0107611f $X=18.705 $Y=2.465
+ $X2=0 $Y2=0
cc_1392 N_A_3416_137#_c_2134_n N_VPWR_c_2191_n 0.0128958f $X=17.225 $Y=1.98
+ $X2=0 $Y2=0
cc_1393 N_A_3416_137#_c_2134_n N_Q_N_c_2631_n 0.057812f $X=17.225 $Y=1.98 $X2=0
+ $Y2=0
cc_1394 N_A_3416_137#_c_2136_n N_Q_N_c_2631_n 0.0216849f $X=17.225 $Y=1.47 $X2=0
+ $Y2=0
cc_1395 N_A_3416_137#_c_2133_n N_Q_N_c_2632_n 0.0425814f $X=17.225 $Y=0.895
+ $X2=0 $Y2=0
cc_1396 N_A_3416_137#_M1012_g N_Q_c_2665_n 0.00323857f $X=18.345 $Y=0.685 $X2=0
+ $Y2=0
cc_1397 N_A_3416_137#_M1053_g N_Q_c_2665_n 0.00430008f $X=18.345 $Y=2.465 $X2=0
+ $Y2=0
cc_1398 N_A_3416_137#_M1020_g N_Q_c_2665_n 0.0238324f $X=18.705 $Y=0.685 $X2=0
+ $Y2=0
cc_1399 N_A_3416_137#_M1058_g N_Q_c_2665_n 0.0300568f $X=18.705 $Y=2.465 $X2=0
+ $Y2=0
cc_1400 N_A_3416_137#_c_2135_n N_Q_c_2665_n 0.0250026f $X=18.41 $Y=1.47 $X2=0
+ $Y2=0
cc_1401 N_A_3416_137#_c_2137_n N_Q_c_2665_n 0.0121537f $X=18.705 $Y=1.47 $X2=0
+ $Y2=0
cc_1402 N_A_3416_137#_M1012_g N_VGND_c_2687_n 0.0221425f $X=18.345 $Y=0.685
+ $X2=0 $Y2=0
cc_1403 N_A_3416_137#_M1020_g N_VGND_c_2687_n 0.00336955f $X=18.705 $Y=0.685
+ $X2=0 $Y2=0
cc_1404 N_A_3416_137#_c_2133_n N_VGND_c_2687_n 0.0137622f $X=17.225 $Y=0.895
+ $X2=0 $Y2=0
cc_1405 N_A_3416_137#_c_2135_n N_VGND_c_2687_n 0.0275493f $X=18.41 $Y=1.47 $X2=0
+ $Y2=0
cc_1406 N_A_3416_137#_c_2137_n N_VGND_c_2687_n 5.79521e-19 $X=18.705 $Y=1.47
+ $X2=0 $Y2=0
cc_1407 N_A_3416_137#_c_2133_n N_VGND_c_2696_n 0.00619475f $X=17.225 $Y=0.895
+ $X2=0 $Y2=0
cc_1408 N_A_3416_137#_M1012_g N_VGND_c_2697_n 0.00461019f $X=18.345 $Y=0.685
+ $X2=0 $Y2=0
cc_1409 N_A_3416_137#_M1020_g N_VGND_c_2697_n 0.00520813f $X=18.705 $Y=0.685
+ $X2=0 $Y2=0
cc_1410 N_A_3416_137#_M1012_g N_VGND_c_2698_n 0.00803623f $X=18.345 $Y=0.685
+ $X2=0 $Y2=0
cc_1411 N_A_3416_137#_M1020_g N_VGND_c_2698_n 0.0104f $X=18.705 $Y=0.685 $X2=0
+ $Y2=0
cc_1412 N_A_3416_137#_c_2133_n N_VGND_c_2698_n 0.00970591f $X=17.225 $Y=0.895
+ $X2=0 $Y2=0
cc_1413 A_125_491# N_VPWR_c_2191_n 0.00899413f $X=0.625 $Y=2.455 $X2=18.96
+ $Y2=3.33
cc_1414 N_VPWR_c_2191_n A_342_491# 0.010279f $X=18.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1415 N_VPWR_c_2191_n N_A_342_261#_M1014_d 0.0022543f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1416 N_VPWR_c_2191_n N_A_342_261#_M1048_d 0.00225781f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1417 N_VPWR_c_2192_n N_A_342_261#_c_2410_n 0.0105911f $X=1.125 $Y=2.805 $X2=0
+ $Y2=0
cc_1418 N_VPWR_c_2192_n N_A_342_261#_c_2411_n 0.0125256f $X=1.125 $Y=2.805 $X2=0
+ $Y2=0
cc_1419 N_VPWR_c_2193_n N_A_342_261#_c_2440_n 0.018058f $X=3.06 $Y=2.805 $X2=0
+ $Y2=0
cc_1420 N_VPWR_c_2205_n N_A_342_261#_c_2440_n 0.0178561f $X=2.895 $Y=3.33 $X2=0
+ $Y2=0
cc_1421 N_VPWR_c_2191_n N_A_342_261#_c_2440_n 0.0124703f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1422 N_VPWR_c_2193_n N_A_342_261#_c_2412_n 0.0234047f $X=3.06 $Y=2.805 $X2=0
+ $Y2=0
cc_1423 N_VPWR_M1023_d N_A_342_261#_c_2421_n 0.00257422f $X=2.92 $Y=2.455 $X2=0
+ $Y2=0
cc_1424 N_VPWR_c_2193_n N_A_342_261#_c_2421_n 0.0149798f $X=3.06 $Y=2.805 $X2=0
+ $Y2=0
cc_1425 N_VPWR_c_2206_n N_A_342_261#_c_2422_n 0.0354956f $X=5.86 $Y=3.33 $X2=0
+ $Y2=0
cc_1426 N_VPWR_c_2191_n N_A_342_261#_c_2422_n 0.0335044f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1427 N_VPWR_M1023_d N_A_342_261#_c_2489_n 0.00350184f $X=2.92 $Y=2.455 $X2=0
+ $Y2=0
cc_1428 N_VPWR_c_2193_n N_A_342_261#_c_2489_n 0.0224397f $X=3.06 $Y=2.805 $X2=0
+ $Y2=0
cc_1429 N_VPWR_c_2206_n N_A_342_261#_c_2489_n 0.00596366f $X=5.86 $Y=3.33 $X2=0
+ $Y2=0
cc_1430 N_VPWR_c_2191_n N_A_342_261#_c_2489_n 0.0060058f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1431 N_VPWR_c_2191_n A_506_491# 0.010279f $X=18.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1432 N_VPWR_c_2191_n A_735_491# 0.00201892f $X=18.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1433 N_VPWR_c_2191_n A_1020_491# 0.00779746f $X=18.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1434 N_VPWR_c_2191_n A_1375_535# 0.00195399f $X=18.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1435 N_VPWR_c_2191_n A_1870_367# 0.0039513f $X=18.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1436 N_VPWR_c_2191_n N_A_2081_439#_M1018_s 0.00232217f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1437 N_VPWR_c_2207_n N_A_2081_439#_c_2553_n 0.0159903f $X=12.495 $Y=3.33
+ $X2=0 $Y2=0
cc_1438 N_VPWR_c_2191_n N_A_2081_439#_c_2553_n 0.00852175f $X=18.96 $Y=3.33
+ $X2=0 $Y2=0
cc_1439 N_VPWR_c_2207_n N_A_2081_439#_c_2555_n 0.0936459f $X=12.495 $Y=3.33
+ $X2=0 $Y2=0
cc_1440 N_VPWR_c_2191_n N_A_2081_439#_c_2555_n 0.056634f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1441 N_VPWR_c_2197_n N_A_2523_397#_c_2586_n 0.0125556f $X=14.095 $Y=2.865
+ $X2=0 $Y2=0
cc_1442 N_VPWR_c_2202_n N_A_2523_397#_c_2586_n 0.0177637f $X=15.71 $Y=3.33 $X2=0
+ $Y2=0
cc_1443 N_VPWR_c_2191_n N_A_2523_397#_c_2586_n 0.0122287f $X=18.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1444 N_VPWR_c_2198_n N_Q_N_c_2635_n 0.0369704f $X=15.875 $Y=2.125 $X2=0 $Y2=0
cc_1445 N_VPWR_c_2209_n N_Q_N_c_2635_n 0.0220321f $X=17.965 $Y=3.33 $X2=0 $Y2=0
cc_1446 N_VPWR_c_2191_n N_Q_N_c_2635_n 0.0125808f $X=18.96 $Y=3.33 $X2=0 $Y2=0
cc_1447 N_VPWR_c_2191_n A_3684_367# 0.00899413f $X=18.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1448 N_VPWR_c_2191_n N_Q_M1058_d 0.0023218f $X=18.96 $Y=3.33 $X2=0 $Y2=0
cc_1449 N_VPWR_c_2199_n N_Q_c_2665_n 0.0418217f $X=18.13 $Y=1.98 $X2=0 $Y2=0
cc_1450 N_VPWR_c_2210_n N_Q_c_2665_n 0.019758f $X=18.96 $Y=3.33 $X2=0 $Y2=0
cc_1451 N_VPWR_c_2191_n N_Q_c_2665_n 0.012508f $X=18.96 $Y=3.33 $X2=0 $Y2=0
cc_1452 N_A_342_261#_c_2422_n A_735_491# 0.00499711f $X=4.375 $Y=2.837 $X2=-0.19
+ $Y2=-0.245
cc_1453 N_A_342_261#_c_2407_n N_noxref_37_c_2854_n 0.0270263f $X=1.07 $Y=2.145
+ $X2=0 $Y2=0
cc_1454 N_A_342_261#_c_2408_n N_noxref_37_c_2854_n 0.0130585f $X=1.685 $Y=1.15
+ $X2=0 $Y2=0
cc_1455 N_A_342_261#_c_2408_n N_noxref_37_c_2855_n 0.00496156f $X=1.685 $Y=1.15
+ $X2=0 $Y2=0
cc_1456 N_A_342_261#_c_2410_n N_noxref_37_c_2855_n 0.0388355f $X=2.075 $Y=2.23
+ $X2=0 $Y2=0
cc_1457 N_A_342_261#_c_2439_n N_noxref_37_c_2855_n 0.0204355f $X=1.85 $Y=1.45
+ $X2=0 $Y2=0
cc_1458 N_A_342_261#_c_2412_n N_noxref_37_c_2855_n 0.0528431f $X=3.405 $Y=2.23
+ $X2=0 $Y2=0
cc_1459 N_A_342_261#_c_2417_n N_noxref_37_c_2855_n 0.0260797f $X=2.24 $Y=2.23
+ $X2=0 $Y2=0
cc_1460 N_A_342_261#_c_2407_n N_noxref_37_c_2856_n 0.0127005f $X=1.07 $Y=2.145
+ $X2=0 $Y2=0
cc_1461 N_A_342_261#_c_2410_n N_noxref_37_c_2856_n 0.0127932f $X=2.075 $Y=2.23
+ $X2=0 $Y2=0
cc_1462 N_A_342_261#_c_2439_n N_noxref_39_c_2888_n 0.0124162f $X=1.85 $Y=1.45
+ $X2=0 $Y2=0
cc_1463 N_A_342_261#_c_2408_n N_noxref_39_c_2890_n 0.00637892f $X=1.685 $Y=1.15
+ $X2=0 $Y2=0
cc_1464 N_Q_N_c_2632_n N_VGND_c_2686_n 0.0167815f $X=16.665 $Y=0.43 $X2=0 $Y2=0
cc_1465 N_Q_N_c_2632_n N_VGND_c_2696_n 0.0232759f $X=16.665 $Y=0.43 $X2=0 $Y2=0
cc_1466 N_Q_N_M1031_d N_VGND_c_2698_n 0.0023218f $X=16.525 $Y=0.235 $X2=0 $Y2=0
cc_1467 N_Q_N_c_2632_n N_VGND_c_2698_n 0.0143828f $X=16.665 $Y=0.43 $X2=0 $Y2=0
cc_1468 N_Q_c_2665_n N_VGND_c_2687_n 0.0287733f $X=18.92 $Y=0.43 $X2=0 $Y2=0
cc_1469 N_Q_c_2665_n N_VGND_c_2697_n 0.019758f $X=18.92 $Y=0.43 $X2=0 $Y2=0
cc_1470 N_Q_c_2665_n N_VGND_c_2698_n 0.0125705f $X=18.92 $Y=0.43 $X2=0 $Y2=0
cc_1471 A_116_47# N_VGND_c_2698_n 0.00307274f $X=0.58 $Y=0.235 $X2=18.96 $Y2=0
cc_1472 N_VGND_M1041_s N_noxref_39_c_2892_n 0.00176502f $X=3.44 $Y=0.215 $X2=0
+ $Y2=0
cc_1473 N_VGND_c_2682_n N_noxref_39_c_2892_n 0.00497259f $X=3.565 $Y=0.38 $X2=0
+ $Y2=0
cc_1474 N_VGND_c_2688_n N_noxref_39_c_2892_n 0.00213516f $X=6.995 $Y=0 $X2=0
+ $Y2=0
cc_1475 N_VGND_c_2698_n N_noxref_39_c_2892_n 0.00474902f $X=18.96 $Y=0 $X2=0
+ $Y2=0
cc_1476 N_VGND_M1041_s N_noxref_39_c_2893_n 0.00210986f $X=3.44 $Y=0.215 $X2=0
+ $Y2=0
cc_1477 N_VGND_c_2682_n N_noxref_39_c_2893_n 0.00880633f $X=3.565 $Y=0.38 $X2=0
+ $Y2=0
cc_1478 N_VGND_c_2693_n N_noxref_39_c_2893_n 0.00103404f $X=3.48 $Y=0 $X2=0
+ $Y2=0
cc_1479 N_VGND_c_2698_n N_noxref_39_c_2893_n 0.00230244f $X=18.96 $Y=0 $X2=0
+ $Y2=0
cc_1480 N_VGND_c_2682_n N_noxref_39_c_2894_n 0.0208116f $X=3.565 $Y=0.38 $X2=0
+ $Y2=0
cc_1481 N_VGND_c_2688_n N_noxref_39_c_2894_n 0.0248299f $X=6.995 $Y=0 $X2=0
+ $Y2=0
cc_1482 N_VGND_c_2698_n N_noxref_39_c_2894_n 0.0130041f $X=18.96 $Y=0 $X2=0
+ $Y2=0
cc_1483 N_VGND_c_2698_n A_1880_47# 0.00282558f $X=18.96 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1484 N_VGND_c_2698_n A_3075_47# 0.00899413f $X=18.96 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1485 N_VGND_c_2698_n A_3233_47# 0.00899413f $X=18.96 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1486 N_noxref_37_c_2855_n N_noxref_39_c_2888_n 0.0167261f $X=2.905 $Y=1.88
+ $X2=0 $Y2=0
cc_1487 N_noxref_37_c_2855_n N_noxref_39_c_2889_n 0.00496145f $X=2.905 $Y=1.88
+ $X2=0 $Y2=0
cc_1488 N_noxref_37_c_2857_n N_noxref_39_c_2889_n 0.0167678f $X=3.07 $Y=1.58
+ $X2=0 $Y2=0
cc_1489 N_noxref_39_c_2889_n N_A_824_219#_c_2943_n 0.00673996f $X=3.415 $Y=1.15
+ $X2=0 $Y2=0
cc_1490 N_noxref_39_c_2891_n N_A_824_219#_c_2943_n 0.00585985f $X=3.5 $Y=1.065
+ $X2=0 $Y2=0
cc_1491 N_noxref_39_c_2894_n N_A_824_219#_c_2943_n 0.00746964f $X=4.055 $Y=0.505
+ $X2=0 $Y2=0
