* File: sky130_fd_sc_lp__mux2i_2.pex.spice
* Created: Wed Sep  2 10:01:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2I_2%S 3 7 11 15 19 23 25 27 31 32 34 37 38 39 48
+ 53
c104 53 0 1.03504e-19 $X=2.47 $Y=1.495
c105 32 0 1.86637e-20 $X=1.85 $Y=1.537
r106 52 53 57.0789 $w=2.28e-07 $l=2.7e-07 $layer=POLY_cond $X=2.2 $Y=1.495
+ $X2=2.47 $Y2=1.495
r107 38 39 19.0044 $w=2.63e-07 $l=4.37e-07 $layer=LI1_cond $X=1.2 $Y=1.987
+ $X2=1.637 $Y2=1.987
r108 37 56 2.89663 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=0.7 $Y=1.987 $X2=0.79
+ $Y2=1.987
r109 37 38 17.5258 $w=2.63e-07 $l=4.03e-07 $layer=LI1_cond $X=0.797 $Y=1.987
+ $X2=1.2 $Y2=1.987
r110 37 56 0.304419 $w=2.63e-07 $l=7e-09 $layer=LI1_cond $X=0.797 $Y=1.987
+ $X2=0.79 $Y2=1.987
r111 35 52 19.0263 $w=2.28e-07 $l=9e-08 $layer=POLY_cond $X=2.11 $Y=1.495
+ $X2=2.2 $Y2=1.495
r112 35 50 14.7982 $w=2.28e-07 $l=7e-08 $layer=POLY_cond $X=2.11 $Y=1.495
+ $X2=2.04 $Y2=1.495
r113 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.51 $X2=2.11 $Y2=1.51
r114 32 34 11.307 $w=2.63e-07 $l=2.6e-07 $layer=LI1_cond $X=1.85 $Y=1.537
+ $X2=2.11 $Y2=1.537
r115 31 39 4.40896 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.765 $Y=1.855
+ $X2=1.765 $Y2=1.987
r116 30 32 7.24806 $w=2.65e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.765 $Y=1.67
+ $X2=1.85 $Y2=1.537
r117 30 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.765 $Y=1.67
+ $X2=1.765 $Y2=1.855
r118 28 48 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.695 $Y=1.51
+ $X2=0.75 $Y2=1.51
r119 28 45 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.695 $Y=1.51
+ $X2=0.56 $Y2=1.51
r120 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.695
+ $Y=1.51 $X2=0.695 $Y2=1.51
r121 25 37 4.2484 $w=1.8e-07 $l=1.32e-07 $layer=LI1_cond $X=0.7 $Y=1.855 $X2=0.7
+ $Y2=1.987
r122 25 27 21.2576 $w=1.78e-07 $l=3.45e-07 $layer=LI1_cond $X=0.7 $Y=1.855
+ $X2=0.7 $Y2=1.51
r123 21 53 33.8246 $w=2.28e-07 $l=1.6e-07 $layer=POLY_cond $X=2.63 $Y=1.495
+ $X2=2.47 $Y2=1.495
r124 21 23 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.63 $Y=1.495
+ $X2=2.63 $Y2=2.465
r125 17 53 12.5943 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.47 $Y=1.345
+ $X2=2.47 $Y2=1.495
r126 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.47 $Y=1.345
+ $X2=2.47 $Y2=0.655
r127 13 52 12.5943 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.2 $Y=1.675
+ $X2=2.2 $Y2=1.495
r128 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.2 $Y=1.675
+ $X2=2.2 $Y2=2.465
r129 9 50 12.5943 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.04 $Y=1.345
+ $X2=2.04 $Y2=1.495
r130 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.04 $Y=1.345
+ $X2=2.04 $Y2=0.655
r131 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.75 $Y=1.345
+ $X2=0.75 $Y2=1.51
r132 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.75 $Y=1.345
+ $X2=0.75 $Y2=0.655
r133 1 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.675
+ $X2=0.56 $Y2=1.51
r134 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.56 $Y=1.675
+ $X2=0.56 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%A_44_367# 1 2 9 13 17 21 25 29 33 36 37 39
+ 42 46
c76 39 0 1.03504e-19 $X=1.27 $Y=1.5
c77 13 0 7.30391e-20 $X=1.18 $Y=2.465
r78 40 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.27 $Y=1.5 $X2=1.61
+ $Y2=1.5
r79 40 43 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.27 $Y=1.5 $X2=1.18
+ $Y2=1.5
r80 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.5 $X2=1.27 $Y2=1.5
r81 37 39 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.13 $Y=1.5 $X2=1.27
+ $Y2=1.5
r82 36 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.045 $Y=1.415
+ $X2=1.13 $Y2=1.5
r83 35 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.045 $Y=1.155
+ $X2=1.045 $Y2=1.415
r84 34 42 4.08752 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.63 $Y=1.07
+ $X2=0.405 $Y2=1.07
r85 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.96 $Y=1.07
+ $X2=1.045 $Y2=1.155
r86 33 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.96 $Y=1.07
+ $X2=0.63 $Y2=1.07
r87 29 31 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.31 $Y=1.98 $X2=0.31
+ $Y2=2.91
r88 27 42 2.70057 $w=3.55e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.31 $Y=1.155
+ $X2=0.405 $Y2=1.07
r89 27 29 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=0.31 $Y=1.155
+ $X2=0.31 $Y2=1.98
r90 23 42 2.70057 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.405 $Y=0.985
+ $X2=0.405 $Y2=1.07
r91 23 25 15.0174 $w=4.48e-07 $l=5.65e-07 $layer=LI1_cond $X=0.405 $Y=0.985
+ $X2=0.405 $Y2=0.42
r92 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.665
+ $X2=1.61 $Y2=1.5
r93 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.61 $Y=1.665 $X2=1.61
+ $Y2=2.465
r94 15 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.335
+ $X2=1.61 $Y2=1.5
r95 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.61 $Y=1.335
+ $X2=1.61 $Y2=0.655
r96 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.5
r97 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.18 $Y=1.665 $X2=1.18
+ $Y2=2.465
r98 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.335
+ $X2=1.18 $Y2=1.5
r99 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.18 $Y=1.335 $X2=1.18
+ $Y2=0.655
r100 2 31 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.835 $X2=0.345 $Y2=2.91
r101 2 29 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.835 $X2=0.345 $Y2=1.98
r102 1 25 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.41
+ $Y=0.235 $X2=0.535 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%A0 3 7 11 15 17 18 26
c59 26 0 2.929e-20 $X=4.19 $Y=1.51
c60 7 0 4.83235e-20 $X=3.76 $Y=2.465
r61 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.1 $Y=1.51 $X2=4.19
+ $Y2=1.51
r62 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=1.51 $X2=4.1 $Y2=1.51
r63 21 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.76 $Y=1.51 $X2=4.1
+ $Y2=1.51
r64 18 25 16.3115 $w=3.23e-07 $l=4.6e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.1 $Y2=1.587
r65 17 25 0.709196 $w=3.23e-07 $l=2e-08 $layer=LI1_cond $X=4.08 $Y=1.587 $X2=4.1
+ $Y2=1.587
r66 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.675
+ $X2=4.19 $Y2=1.51
r67 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.19 $Y=1.675
+ $X2=4.19 $Y2=2.465
r68 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.345
+ $X2=4.19 $Y2=1.51
r69 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.19 $Y=1.345
+ $X2=4.19 $Y2=0.765
r70 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.76 $Y=1.675
+ $X2=3.76 $Y2=1.51
r71 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.76 $Y=1.675 $X2=3.76
+ $Y2=2.465
r72 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.76 $Y=1.345
+ $X2=3.76 $Y2=1.51
r73 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.76 $Y=1.345 $X2=3.76
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%A1 3 7 9 13 17 19 20 21 24
c49 21 0 2.929e-20 $X=5.52 $Y=1.665
r50 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.12 $Y=1.51
+ $X2=5.12 $Y2=1.675
r51 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.51 $X2=5.12 $Y2=1.51
r52 24 27 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.12 $Y=1.42 $X2=5.12
+ $Y2=1.51
r53 24 25 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.12 $Y=1.42 $X2=5.12
+ $Y2=1.345
r54 21 28 14.1839 $w=3.23e-07 $l=4e-07 $layer=LI1_cond $X=5.52 $Y=1.587 $X2=5.12
+ $Y2=1.587
r55 20 28 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=5.04 $Y=1.587 $X2=5.12
+ $Y2=1.587
r56 17 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.21 $Y=0.765
+ $X2=5.21 $Y2=1.345
r57 13 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.05 $Y=2.465
+ $X2=5.05 $Y2=1.675
r58 10 19 5.30422 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=4.775 $Y=1.42
+ $X2=4.66 $Y2=1.42
r59 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.42
+ $X2=5.12 $Y2=1.42
r60 9 10 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.955 $Y=1.42
+ $X2=4.775 $Y2=1.42
r61 5 19 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=4.7 $Y=1.345
+ $X2=4.66 $Y2=1.42
r62 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.7 $Y=1.345 $X2=4.7
+ $Y2=0.765
r63 1 19 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=4.62 $Y=1.495
+ $X2=4.66 $Y2=1.42
r64 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=4.62 $Y=1.495 $X2=4.62
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%VPWR 1 2 3 14 17 20 23 29 35 36 39 42
r70 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r71 42 45 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.96 $Y=3.045
+ $X2=2.96 $Y2=3.33
r72 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 36 46 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=3.12 $Y2=3.33
r74 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 33 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=2.96 $Y2=3.33
r76 33 35 156.251 $w=1.68e-07 $l=2.395e-06 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=5.52 $Y2=3.33
r77 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 29 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.96 $Y2=3.33
r79 29 31 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.64 $Y2=3.33
r80 28 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 28 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.875 $Y2=3.33
r84 25 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.04 $Y=3.33 $X2=1.68
+ $Y2=3.33
r85 23 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r86 23 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 21 31 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 20 27 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.74 $Y=3.33 $X2=1.68
+ $Y2=3.33
r89 19 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.07 $Y2=3.33
r90 19 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r91 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.905 $Y=3.045
+ $X2=1.905 $Y2=3.33
r92 12 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r93 12 14 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.375
r94 3 42 600 $w=1.7e-07 $l=1.33141e-06 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.96 $Y2=3.045
r95 2 17 600 $w=1.7e-07 $l=1.31541e-06 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.835 $X2=1.905 $Y2=3.045
r96 1 14 300 $w=1.7e-07 $l=6.48999e-07 $layer=licon1_PDIFF $count=2 $X=0.635
+ $Y=1.835 $X2=0.875 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%A_251_367# 1 2 7 9 13 16 20
c49 7 0 5.43754e-20 $X=3.305 $Y=2.685
r50 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.39 $Y=2.685
+ $X2=3.39 $Y2=2.99
r51 16 18 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.395 $Y=2.375
+ $X2=1.395 $Y2=2.685
r52 11 13 24.0733 $w=2.23e-07 $l=4.7e-07 $layer=LI1_cond $X=4.852 $Y=2.905
+ $X2=4.852 $Y2=2.435
r53 10 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=2.99
+ $X2=3.39 $Y2=2.99
r54 9 11 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.74 $Y=2.99
+ $X2=4.852 $Y2=2.905
r55 9 10 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=4.74 $Y=2.99
+ $X2=3.475 $Y2=2.99
r56 8 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=2.685
+ $X2=1.395 $Y2=2.685
r57 7 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=2.685
+ $X2=3.39 $Y2=2.685
r58 7 8 113.845 $w=1.68e-07 $l=1.745e-06 $layer=LI1_cond $X=3.305 $Y=2.685
+ $X2=1.56 $Y2=2.685
r59 2 13 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=4.695
+ $Y=1.835 $X2=4.835 $Y2=2.435
r60 1 16 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=1.255
+ $Y=1.835 $X2=1.395 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%A_455_367# 1 2 9 11 12 15
r30 13 15 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=3.94 $Y=2.43
+ $X2=3.94 $Y2=2.57
r31 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.81 $Y=2.345
+ $X2=3.94 $Y2=2.43
r32 11 12 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.81 $Y=2.345
+ $X2=2.58 $Y2=2.345
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=2.26
+ $X2=2.58 $Y2=2.345
r34 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=2.26
+ $X2=2.415 $Y2=2.005
r35 2 15 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.835 $X2=3.975 $Y2=2.57
r36 1 9 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%Y 1 2 3 4 5 6 19 21 27 29 31 33 35 39 41 45
+ 46 49 50 63
c88 45 0 4.83235e-20 $X=4.405 $Y=2.095
r89 50 63 8.28896 $w=5.08e-07 $l=1.1e-07 $layer=LI1_cond $X=3.6 $Y=1.835
+ $X2=3.71 $Y2=1.835
r90 50 60 1.28989 $w=5.08e-07 $l=5.5e-08 $layer=LI1_cond $X=3.6 $Y=1.835
+ $X2=3.545 $Y2=1.835
r91 50 60 3.28461 $w=3.3e-07 $l=2.55e-07 $layer=LI1_cond $X=3.545 $Y=1.58
+ $X2=3.545 $Y2=1.835
r92 49 60 9.96732 $w=5.08e-07 $l=4.25e-07 $layer=LI1_cond $X=3.12 $Y=1.835
+ $X2=3.545 $Y2=1.835
r93 41 50 9.03645 $w=4.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.545 $Y=1.245
+ $X2=3.545 $Y2=1.58
r94 41 43 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.545 $Y=1.245
+ $X2=3.545 $Y2=1.105
r95 37 39 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=5.46 $Y=1.075
+ $X2=5.46 $Y2=0.495
r96 33 48 2.79092 $w=2.95e-07 $l=9e-08 $layer=LI1_cond $X=5.282 $Y=2.1 $X2=5.282
+ $Y2=2.01
r97 33 35 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=5.282 $Y=2.1
+ $X2=5.282 $Y2=2.46
r98 32 46 7.01393 $w=2.25e-07 $l=1.90526e-07 $layer=LI1_cond $X=4.65 $Y=1.16
+ $X2=4.485 $Y2=1.105
r99 31 37 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.33 $Y=1.16
+ $X2=5.46 $Y2=1.075
r100 31 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.33 $Y=1.16
+ $X2=4.65 $Y2=1.16
r101 30 45 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=4.57 $Y=2.01
+ $X2=4.405 $Y2=2.01
r102 29 48 4.55851 $w=1.8e-07 $l=1.47e-07 $layer=LI1_cond $X=5.135 $Y=2.01
+ $X2=5.282 $Y2=2.01
r103 29 30 34.8131 $w=1.78e-07 $l=5.65e-07 $layer=LI1_cond $X=5.135 $Y=2.01
+ $X2=4.57 $Y2=2.01
r104 25 46 0.00725833 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=4.485 $Y=0.965
+ $X2=4.485 $Y2=1.105
r105 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.485 $Y=0.965
+ $X2=4.485 $Y2=0.69
r106 21 45 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.24 $Y=2.005
+ $X2=4.405 $Y2=2.01
r107 21 63 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.24 $Y=2.005
+ $X2=3.71 $Y2=2.005
r108 20 43 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=1.105
+ $X2=3.545 $Y2=1.105
r109 19 46 7.01393 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=1.105
+ $X2=4.485 $Y2=1.105
r110 19 20 25.1068 $w=2.78e-07 $l=6.1e-07 $layer=LI1_cond $X=4.32 $Y=1.105
+ $X2=3.71 $Y2=1.105
r111 6 48 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=5.125
+ $Y=1.835 $X2=5.265 $Y2=2.005
r112 6 35 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.835 $X2=5.265 $Y2=2.46
r113 5 45 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=4.265
+ $Y=1.835 $X2=4.405 $Y2=2.095
r114 4 60 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.835 $X2=3.545 $Y2=1.995
r115 3 39 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.345 $X2=5.425 $Y2=0.495
r116 2 27 91 $w=1.7e-07 $l=4.41503e-07 $layer=licon1_NDIFF $count=2 $X=4.265
+ $Y=0.345 $X2=4.485 $Y2=0.69
r117 1 43 182 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.345 $X2=3.545 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%VGND 1 2 3 12 17 18 20 23 24 26 27 28 41 42
r59 41 42 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r60 38 41 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=5.52
+ $Y2=0
r61 38 39 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 36 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r63 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 32 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r65 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 28 42 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=5.52
+ $Y2=0
r67 28 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r68 26 35 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.68
+ $Y2=0
r69 26 27 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.81
+ $Y2=0
r70 25 38 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r71 25 27 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.81
+ $Y2=0
r72 23 31 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.72
+ $Y2=0
r73 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.965
+ $Y2=0
r74 22 35 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=1.68
+ $Y2=0
r75 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=0.965
+ $Y2=0
r76 18 20 40.0736 $w=2.18e-07 $l=7.65e-07 $layer=LI1_cond $X=1.92 $Y=0.785
+ $X2=2.685 $Y2=0.785
r77 15 18 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=1.81 $Y=0.675
+ $X2=1.92 $Y2=0.785
r78 15 17 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=1.81 $Y=0.675
+ $X2=1.81 $Y2=0.38
r79 14 27 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0
r80 14 17 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.38
r81 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=0.085
+ $X2=0.965 $Y2=0
r82 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.965 $Y=0.085
+ $X2=0.965 $Y2=0.36
r83 3 20 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.235 $X2=2.685 $Y2=0.78
r84 2 17 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.685
+ $Y=0.235 $X2=1.825 $Y2=0.38
r85 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.825
+ $Y=0.235 $X2=0.965 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%A_251_47# 1 2 9 11 12 14 15 17
r45 15 17 44.6555 $w=1.88e-07 $l=7.65e-07 $layer=LI1_cond $X=3.21 $Y=0.7
+ $X2=3.975 $Y2=0.7
r46 13 15 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=3.115 $Y=0.795
+ $X2=3.21 $Y2=0.7
r47 13 14 15.7608 $w=1.88e-07 $l=2.7e-07 $layer=LI1_cond $X=3.115 $Y=0.795
+ $X2=3.115 $Y2=1.065
r48 11 14 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.02 $Y=1.15
+ $X2=3.115 $Y2=1.065
r49 11 12 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=3.02 $Y=1.15
+ $X2=1.53 $Y2=1.15
r50 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.415 $Y=1.065
+ $X2=1.53 $Y2=1.15
r51 7 9 32.3185 $w=2.28e-07 $l=6.45e-07 $layer=LI1_cond $X=1.415 $Y=1.065
+ $X2=1.415 $Y2=0.42
r52 2 17 182 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.345 $X2=3.975 $Y2=0.71
r53 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.255
+ $Y=0.235 $X2=1.395 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_2%A_423_47# 1 2 7 11 16
r31 14 16 8.52828 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=0.38
+ $X2=2.42 $Y2=0.38
r32 9 11 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=4.995 $Y=0.435
+ $X2=4.995 $Y2=0.47
r33 7 9 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.83 $Y=0.345
+ $X2=4.995 $Y2=0.435
r34 7 16 148.495 $w=1.78e-07 $l=2.41e-06 $layer=LI1_cond $X=4.83 $Y=0.345
+ $X2=2.42 $Y2=0.345
r35 2 11 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=4.775
+ $Y=0.345 $X2=4.995 $Y2=0.47
r36 1 14 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.255 $Y2=0.38
.ends

