* File: sky130_fd_sc_lp__a2111o_0.spice
* Created: Fri Aug 28 09:45:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111o_0.pex.spice"
.subckt sky130_fd_sc_lp__a2111o_0  VNB VPB D1 C1 B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_80_159#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_80_159#_M1001_d N_D1_M1001_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_C1_M1007_g N_A_80_159#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1386 AS=0.0588 PD=1.08 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_80_159#_M1004_d N_B1_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1386 PD=0.7 PS=1.08 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1010 A_582_47# N_A1_M1010_g N_A_80_159#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A2_M1011_g A_582_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_80_159#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 A_312_476# N_D1_M1002_g N_A_80_159#_M1002_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.81 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1009 A_390_476# N_C1_M1009_g A_312_476# VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=19.9955 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1003 N_A_468_476#_M1003_d N_B1_M1003_g A_390_476# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1584 AS=0.0768 PD=1.135 PS=0.88 NRD=33.0763 NRS=19.9955 M=1 R=4.26667
+ SA=75001 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_468_476#_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1584 PD=0.92 PS=1.135 NRD=0 NRS=33.0763 M=1 R=4.26667
+ SA=75001.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_468_476#_M1000_d N_A2_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a2111o_0.pxi.spice"
*
.ends
*
*
