* File: sky130_fd_sc_lp__a41o_1.pxi.spice
* Created: Wed Sep  2 09:28:55 2020
* 
x_PM_SKY130_FD_SC_LP__A41O_1%A_113_237# N_A_113_237#_M1010_d
+ N_A_113_237#_M1011_s N_A_113_237#_M1008_g N_A_113_237#_c_62_n
+ N_A_113_237#_M1001_g N_A_113_237#_c_63_n N_A_113_237#_c_64_n
+ N_A_113_237#_c_76_p N_A_113_237#_c_108_p N_A_113_237#_c_65_n
+ N_A_113_237#_c_66_n N_A_113_237#_c_70_n N_A_113_237#_c_85_p
+ PM_SKY130_FD_SC_LP__A41O_1%A_113_237#
x_PM_SKY130_FD_SC_LP__A41O_1%B1 N_B1_M1010_g N_B1_M1011_g B1 B1 N_B1_c_120_n
+ N_B1_c_121_n PM_SKY130_FD_SC_LP__A41O_1%B1
x_PM_SKY130_FD_SC_LP__A41O_1%A1 N_A1_M1005_g N_A1_c_154_n N_A1_M1002_g A1 A1 A1
+ N_A1_c_156_n PM_SKY130_FD_SC_LP__A41O_1%A1
x_PM_SKY130_FD_SC_LP__A41O_1%A2 N_A2_M1000_g N_A2_M1003_g A2 A2 A2 N_A2_c_190_n
+ N_A2_c_191_n PM_SKY130_FD_SC_LP__A41O_1%A2
x_PM_SKY130_FD_SC_LP__A41O_1%A3 N_A3_M1004_g N_A3_M1009_g A3 A3 A3 N_A3_c_223_n
+ N_A3_c_224_n PM_SKY130_FD_SC_LP__A41O_1%A3
x_PM_SKY130_FD_SC_LP__A41O_1%A4 N_A4_c_256_n N_A4_M1007_g N_A4_M1006_g A4
+ N_A4_c_259_n PM_SKY130_FD_SC_LP__A41O_1%A4
x_PM_SKY130_FD_SC_LP__A41O_1%X N_X_M1001_s N_X_M1008_s X X X X X X X N_X_c_279_n
+ PM_SKY130_FD_SC_LP__A41O_1%X
x_PM_SKY130_FD_SC_LP__A41O_1%VPWR N_VPWR_M1008_d N_VPWR_M1005_d N_VPWR_M1009_d
+ N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n
+ VPWR N_VPWR_c_298_n N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_292_n
+ N_VPWR_c_302_n N_VPWR_c_303_n PM_SKY130_FD_SC_LP__A41O_1%VPWR
x_PM_SKY130_FD_SC_LP__A41O_1%A_346_367# N_A_346_367#_M1011_d
+ N_A_346_367#_M1003_d N_A_346_367#_M1006_d N_A_346_367#_c_375_n
+ N_A_346_367#_c_348_n N_A_346_367#_c_349_n N_A_346_367#_c_379_n
+ N_A_346_367#_c_350_n N_A_346_367#_c_351_n N_A_346_367#_c_352_n
+ PM_SKY130_FD_SC_LP__A41O_1%A_346_367#
x_PM_SKY130_FD_SC_LP__A41O_1%VGND N_VGND_M1001_d N_VGND_M1007_d N_VGND_c_385_n
+ N_VGND_c_386_n VGND N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n
+ N_VGND_c_390_n PM_SKY130_FD_SC_LP__A41O_1%VGND
cc_1 VNB N_A_113_237#_M1008_g 0.0091365f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_2 VNB N_A_113_237#_c_62_n 0.0223684f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.185
cc_3 VNB N_A_113_237#_c_63_n 0.00338266f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.35
cc_4 VNB N_A_113_237#_c_64_n 0.0480979f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.35
cc_5 VNB N_A_113_237#_c_65_n 0.00638943f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.69
cc_6 VNB N_A_113_237#_c_66_n 2.94739e-19 $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.69
cc_7 VNB N_B1_M1011_g 0.00867994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB B1 0.00761973f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_9 VNB N_B1_c_120_n 0.04631f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.655
cc_10 VNB N_B1_c_121_n 0.021652f $X=-0.19 $Y=-0.245 $X2=0.842 $Y2=1.605
cc_11 VNB N_A1_M1005_g 0.00705582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_c_154_n 0.0173085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A1 0.00135578f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_14 VNB N_A1_c_156_n 0.040921f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.955
cc_15 VNB N_A2_M1003_g 0.00881095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A2 0.00581686f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_17 VNB N_A2_c_190_n 0.0328143f $X=-0.19 $Y=-0.245 $X2=0.842 $Y2=1.605
cc_18 VNB N_A2_c_191_n 0.0155803f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.35
cc_19 VNB N_A3_M1009_g 0.00774896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A3 0.00745973f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_21 VNB N_A3_c_223_n 0.0285375f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.69
cc_22 VNB N_A3_c_224_n 0.0172487f $X=-0.19 $Y=-0.245 $X2=1.422 $Y2=1.775
cc_23 VNB N_A4_c_256_n 0.0226103f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.235
cc_24 VNB N_A4_M1006_g 0.0116295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB A4 0.0202977f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_26 VNB N_A4_c_259_n 0.0424276f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.655
cc_27 VNB N_X_c_279_n 0.0713003f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.69
cc_28 VNB N_VPWR_c_292_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_385_n 0.0134879f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.515
cc_30 VNB N_VGND_c_386_n 0.0350086f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.465
cc_31 VNB N_VGND_c_387_n 0.0612483f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.35
cc_32 VNB N_VGND_c_388_n 0.0204132f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=0.87
cc_33 VNB N_VGND_c_389_n 0.0159665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_390_n 0.233322f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.35
cc_35 VPB N_A_113_237#_M1008_g 0.0282539f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.465
cc_36 VPB N_A_113_237#_c_65_n 0.0127632f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.69
cc_37 VPB N_A_113_237#_c_66_n 0.00355348f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.69
cc_38 VPB N_A_113_237#_c_70_n 0.0151384f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.98
cc_39 VPB N_B1_M1011_g 0.0234317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A1_M1005_g 0.0213983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A2_M1003_g 0.0214003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A3_M1009_g 0.0189942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A4_M1006_g 0.0247156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_X_c_279_n 0.0688374f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.69
cc_45 VPB N_VPWR_c_293_n 0.0171727f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.655
cc_46 VPB N_VPWR_c_294_n 0.00183691f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.35
cc_47 VPB N_VPWR_c_295_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.422 $Y2=1.98
cc_48 VPB N_VPWR_c_296_n 0.0213315f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=0.87
cc_49 VPB N_VPWR_c_297_n 0.00516749f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=0.42
cc_50 VPB N_VPWR_c_298_n 0.0295039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_299_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_300_n 0.0186881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_292_n 0.0606097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_302_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_303_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_346_367#_c_348_n 0.0120706f $X=-0.19 $Y=1.655 $X2=0.842 $Y2=1.35
cc_57 VPB N_A_346_367#_c_349_n 0.00537394f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.35
cc_58 VPB N_A_346_367#_c_350_n 0.0123332f $X=-0.19 $Y=1.655 $X2=1.422 $Y2=1.98
cc_59 VPB N_A_346_367#_c_351_n 0.0465671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_346_367#_c_352_n 0.00326453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 N_A_113_237#_c_63_n N_B1_M1011_g 0.0019258f $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_113_237#_c_65_n N_B1_M1011_g 0.00611255f $X=1.275 $Y=1.69 $X2=0 $Y2=0
cc_63 N_A_113_237#_c_70_n N_B1_M1011_g 0.00442794f $X=1.44 $Y=1.98 $X2=0 $Y2=0
cc_64 N_A_113_237#_c_63_n B1 0.0182129f $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_65 N_A_113_237#_c_64_n B1 0.0017866f $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_66 N_A_113_237#_c_76_p B1 0.0545883f $X=1.725 $Y=0.955 $X2=0 $Y2=0
cc_67 N_A_113_237#_c_65_n B1 0.0364943f $X=1.275 $Y=1.69 $X2=0 $Y2=0
cc_68 N_A_113_237#_c_63_n N_B1_c_120_n 8.90177e-19 $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_69 N_A_113_237#_c_64_n N_B1_c_120_n 0.0161526f $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_70 N_A_113_237#_c_76_p N_B1_c_120_n 0.00765392f $X=1.725 $Y=0.955 $X2=0 $Y2=0
cc_71 N_A_113_237#_c_65_n N_B1_c_120_n 0.00786716f $X=1.275 $Y=1.69 $X2=0 $Y2=0
cc_72 N_A_113_237#_c_63_n N_B1_c_121_n 0.00327397f $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_73 N_A_113_237#_c_76_p N_B1_c_121_n 0.0142704f $X=1.725 $Y=0.955 $X2=0 $Y2=0
cc_74 N_A_113_237#_c_76_p N_A1_c_154_n 5.49694e-19 $X=1.725 $Y=0.955 $X2=0 $Y2=0
cc_75 N_A_113_237#_c_85_p N_A1_c_154_n 0.00385454f $X=1.82 $Y=0.42 $X2=0 $Y2=0
cc_76 N_A_113_237#_M1010_d A1 0.00788225f $X=1.68 $Y=0.235 $X2=0 $Y2=0
cc_77 N_A_113_237#_c_76_p A1 0.0142756f $X=1.725 $Y=0.955 $X2=0 $Y2=0
cc_78 N_A_113_237#_c_85_p A1 0.0362276f $X=1.82 $Y=0.42 $X2=0 $Y2=0
cc_79 N_A_113_237#_M1008_g N_X_c_279_n 0.0310712f $X=0.64 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A_113_237#_c_62_n N_X_c_279_n 0.00488643f $X=0.68 $Y=1.185 $X2=0 $Y2=0
cc_81 N_A_113_237#_c_63_n N_X_c_279_n 0.0414257f $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_82 N_A_113_237#_c_64_n N_X_c_279_n 0.0122211f $X=0.835 $Y=1.35 $X2=0 $Y2=0
cc_83 N_A_113_237#_c_66_n N_X_c_279_n 0.0147231f $X=0.945 $Y=1.69 $X2=0 $Y2=0
cc_84 N_A_113_237#_M1008_g N_VPWR_c_293_n 0.0058595f $X=0.64 $Y=2.465 $X2=0
+ $Y2=0
cc_85 N_A_113_237#_c_64_n N_VPWR_c_293_n 9.40382e-19 $X=0.835 $Y=1.35 $X2=0
+ $Y2=0
cc_86 N_A_113_237#_c_65_n N_VPWR_c_293_n 0.00615025f $X=1.275 $Y=1.69 $X2=0
+ $Y2=0
cc_87 N_A_113_237#_c_66_n N_VPWR_c_293_n 0.0168876f $X=0.945 $Y=1.69 $X2=0 $Y2=0
cc_88 N_A_113_237#_c_70_n N_VPWR_c_293_n 0.0692919f $X=1.44 $Y=1.98 $X2=0 $Y2=0
cc_89 N_A_113_237#_M1008_g N_VPWR_c_296_n 0.00579312f $X=0.64 $Y=2.465 $X2=0
+ $Y2=0
cc_90 N_A_113_237#_c_70_n N_VPWR_c_298_n 0.0190529f $X=1.44 $Y=1.98 $X2=0 $Y2=0
cc_91 N_A_113_237#_M1011_s N_VPWR_c_292_n 0.00249946f $X=1.315 $Y=1.835 $X2=0
+ $Y2=0
cc_92 N_A_113_237#_M1008_g N_VPWR_c_292_n 0.0128077f $X=0.64 $Y=2.465 $X2=0
+ $Y2=0
cc_93 N_A_113_237#_c_70_n N_VPWR_c_292_n 0.0113912f $X=1.44 $Y=1.98 $X2=0 $Y2=0
cc_94 N_A_113_237#_c_65_n N_A_346_367#_c_349_n 0.00842668f $X=1.275 $Y=1.69
+ $X2=0 $Y2=0
cc_95 N_A_113_237#_c_70_n N_A_346_367#_c_349_n 0.00513286f $X=1.44 $Y=1.98 $X2=0
+ $Y2=0
cc_96 N_A_113_237#_c_63_n N_VGND_M1001_d 5.75986e-19 $X=0.835 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_113_237#_c_76_p N_VGND_M1001_d 0.0150363f $X=1.725 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_113_237#_c_108_p N_VGND_M1001_d 0.00155015f $X=0.945 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_99 N_A_113_237#_c_85_p N_VGND_c_387_n 0.0121325f $X=1.82 $Y=0.42 $X2=0 $Y2=0
cc_100 N_A_113_237#_c_62_n N_VGND_c_388_n 0.00564095f $X=0.68 $Y=1.185 $X2=0
+ $Y2=0
cc_101 N_A_113_237#_c_62_n N_VGND_c_389_n 0.0142455f $X=0.68 $Y=1.185 $X2=0
+ $Y2=0
cc_102 N_A_113_237#_c_64_n N_VGND_c_389_n 7.76243e-19 $X=0.835 $Y=1.35 $X2=0
+ $Y2=0
cc_103 N_A_113_237#_c_76_p N_VGND_c_389_n 0.0445861f $X=1.725 $Y=0.955 $X2=0
+ $Y2=0
cc_104 N_A_113_237#_c_108_p N_VGND_c_389_n 0.0123177f $X=0.945 $Y=0.955 $X2=0
+ $Y2=0
cc_105 N_A_113_237#_M1010_d N_VGND_c_390_n 0.0122133f $X=1.68 $Y=0.235 $X2=0
+ $Y2=0
cc_106 N_A_113_237#_c_62_n N_VGND_c_390_n 0.0105114f $X=0.68 $Y=1.185 $X2=0
+ $Y2=0
cc_107 N_A_113_237#_c_85_p N_VGND_c_390_n 0.00692023f $X=1.82 $Y=0.42 $X2=0
+ $Y2=0
cc_108 N_B1_c_121_n N_A1_c_154_n 0.011334f $X=1.535 $Y=1.185 $X2=0 $Y2=0
cc_109 B1 A1 0.01855f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_B1_c_120_n A1 8.90331e-19 $X=1.635 $Y=1.35 $X2=0 $Y2=0
cc_111 N_B1_c_121_n A1 0.00270573f $X=1.535 $Y=1.185 $X2=0 $Y2=0
cc_112 N_B1_M1011_g N_A1_c_156_n 0.0260655f $X=1.655 $Y=2.465 $X2=0 $Y2=0
cc_113 B1 N_A1_c_156_n 0.00158518f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B1_c_120_n N_A1_c_156_n 0.0216465f $X=1.635 $Y=1.35 $X2=0 $Y2=0
cc_115 N_B1_M1011_g N_VPWR_c_293_n 0.00400223f $X=1.655 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B1_M1011_g N_VPWR_c_294_n 0.00144284f $X=1.655 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B1_M1011_g N_VPWR_c_298_n 0.00585385f $X=1.655 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B1_M1011_g N_VPWR_c_292_n 0.0120903f $X=1.655 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B1_M1011_g N_A_346_367#_c_349_n 0.00132667f $X=1.655 $Y=2.465 $X2=0
+ $Y2=0
cc_120 B1 N_A_346_367#_c_349_n 0.0106005f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_121 N_B1_c_120_n N_A_346_367#_c_349_n 0.00147518f $X=1.635 $Y=1.35 $X2=0
+ $Y2=0
cc_122 N_B1_c_121_n N_VGND_c_387_n 0.00486043f $X=1.535 $Y=1.185 $X2=0 $Y2=0
cc_123 N_B1_c_121_n N_VGND_c_389_n 0.0153744f $X=1.535 $Y=1.185 $X2=0 $Y2=0
cc_124 N_B1_c_121_n N_VGND_c_390_n 0.00875669f $X=1.535 $Y=1.185 $X2=0 $Y2=0
cc_125 N_A1_M1005_g N_A2_M1003_g 0.00945196f $X=2.085 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A1_c_156_n N_A2_M1003_g 0.00119553f $X=2.315 $Y=1.365 $X2=0 $Y2=0
cc_127 N_A1_c_154_n A2 0.00654243f $X=2.315 $Y=1.185 $X2=0 $Y2=0
cc_128 A1 A2 0.0867814f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_129 N_A1_c_156_n N_A2_c_190_n 0.0431028f $X=2.315 $Y=1.365 $X2=0 $Y2=0
cc_130 N_A1_c_154_n N_A2_c_191_n 0.0431028f $X=2.315 $Y=1.185 $X2=0 $Y2=0
cc_131 A1 N_A2_c_191_n 0.00111324f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_132 N_A1_M1005_g N_VPWR_c_294_n 0.018307f $X=2.085 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A1_M1005_g N_VPWR_c_298_n 0.00486043f $X=2.085 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A1_M1005_g N_VPWR_c_292_n 0.0082726f $X=2.085 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A1_M1005_g N_A_346_367#_c_348_n 0.0168914f $X=2.085 $Y=2.465 $X2=0
+ $Y2=0
cc_136 A1 N_A_346_367#_c_348_n 0.0211027f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_137 N_A1_c_156_n N_A_346_367#_c_348_n 0.0067002f $X=2.315 $Y=1.365 $X2=0
+ $Y2=0
cc_138 N_A1_c_154_n N_VGND_c_387_n 0.00445971f $X=2.315 $Y=1.185 $X2=0 $Y2=0
cc_139 A1 N_VGND_c_387_n 0.00882826f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_140 N_A1_c_154_n N_VGND_c_389_n 8.32463e-19 $X=2.315 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A1_c_154_n N_VGND_c_390_n 0.00763243f $X=2.315 $Y=1.185 $X2=0 $Y2=0
cc_142 A1 N_VGND_c_390_n 0.00914594f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A2_M1003_g N_A3_M1009_g 0.0271157f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_144 A2 A3 0.0953814f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_145 N_A2_c_190_n A3 0.00235973f $X=2.765 $Y=1.35 $X2=0 $Y2=0
cc_146 N_A2_c_191_n A3 0.00268387f $X=2.765 $Y=1.185 $X2=0 $Y2=0
cc_147 A2 N_A3_c_223_n 2.88215e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_148 N_A2_c_190_n N_A3_c_223_n 0.0204266f $X=2.765 $Y=1.35 $X2=0 $Y2=0
cc_149 A2 N_A3_c_224_n 0.00229153f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_150 N_A2_c_191_n N_A3_c_224_n 0.0330969f $X=2.765 $Y=1.185 $X2=0 $Y2=0
cc_151 N_A2_M1003_g N_VPWR_c_294_n 0.0171444f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A2_M1003_g N_VPWR_c_295_n 7.17596e-19 $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A2_M1003_g N_VPWR_c_299_n 0.00486043f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A2_M1003_g N_VPWR_c_292_n 0.0082726f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A2_M1003_g N_A_346_367#_c_348_n 0.0175743f $X=2.855 $Y=2.465 $X2=0
+ $Y2=0
cc_156 A2 N_A_346_367#_c_348_n 0.0267356f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A2_c_190_n N_A_346_367#_c_348_n 0.00125478f $X=2.765 $Y=1.35 $X2=0
+ $Y2=0
cc_158 A2 N_VGND_c_387_n 0.0101834f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A2_c_191_n N_VGND_c_387_n 0.00384307f $X=2.765 $Y=1.185 $X2=0 $Y2=0
cc_160 A2 N_VGND_c_390_n 0.0112623f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_161 N_A2_c_191_n N_VGND_c_390_n 0.00564664f $X=2.765 $Y=1.185 $X2=0 $Y2=0
cc_162 A2 A_478_47# 0.00611827f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_163 A2 A_550_47# 0.00666359f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_164 A3 N_A4_c_256_n 0.025456f $X=3.035 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_165 N_A3_c_224_n N_A4_c_256_n 0.0324042f $X=3.305 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A3_M1009_g N_A4_M1006_g 0.0233828f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_167 A3 A4 0.0264094f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_168 N_A3_c_223_n A4 2.15932e-19 $X=3.305 $Y=1.35 $X2=0 $Y2=0
cc_169 A3 N_A4_c_259_n 0.00787909f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_170 N_A3_c_223_n N_A4_c_259_n 0.021443f $X=3.305 $Y=1.35 $X2=0 $Y2=0
cc_171 N_A3_M1009_g N_VPWR_c_294_n 7.67382e-19 $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A3_M1009_g N_VPWR_c_295_n 0.0134639f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A3_M1009_g N_VPWR_c_299_n 0.00564095f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A3_M1009_g N_VPWR_c_292_n 0.00950825f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A3_M1009_g N_A_346_367#_c_350_n 0.0147433f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_176 A3 N_A_346_367#_c_350_n 0.0402185f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A3_c_223_n N_A_346_367#_c_350_n 9.47144e-19 $X=3.305 $Y=1.35 $X2=0
+ $Y2=0
cc_178 A3 N_A_346_367#_c_352_n 0.015162f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_179 N_A3_c_223_n N_A_346_367#_c_352_n 3.51912e-19 $X=3.305 $Y=1.35 $X2=0
+ $Y2=0
cc_180 A3 N_VGND_c_387_n 0.0214915f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_181 N_A3_c_224_n N_VGND_c_387_n 0.00384307f $X=3.305 $Y=1.185 $X2=0 $Y2=0
cc_182 A3 N_VGND_c_390_n 0.0231323f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A3_c_224_n N_VGND_c_390_n 0.00610266f $X=3.305 $Y=1.185 $X2=0 $Y2=0
cc_184 A3 A_550_47# 0.00699873f $X=3.035 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_185 A3 A_658_47# 0.00454243f $X=3.035 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_186 N_A4_M1006_g N_VPWR_c_295_n 0.0154114f $X=3.755 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A4_M1006_g N_VPWR_c_300_n 0.00564095f $X=3.755 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A4_M1006_g N_VPWR_c_292_n 0.0104902f $X=3.755 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A4_M1006_g N_A_346_367#_c_350_n 0.0204172f $X=3.755 $Y=2.465 $X2=0
+ $Y2=0
cc_190 A4 N_A_346_367#_c_350_n 0.0236959f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A4_c_259_n N_A_346_367#_c_350_n 0.00697869f $X=3.95 $Y=1.35 $X2=0 $Y2=0
cc_192 N_A4_c_256_n N_VGND_c_386_n 0.00636314f $X=3.755 $Y=1.185 $X2=0 $Y2=0
cc_193 A4 N_VGND_c_386_n 0.0217129f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A4_c_259_n N_VGND_c_386_n 0.00593911f $X=3.95 $Y=1.35 $X2=0 $Y2=0
cc_195 N_A4_c_256_n N_VGND_c_387_n 0.00580023f $X=3.755 $Y=1.185 $X2=0 $Y2=0
cc_196 N_A4_c_256_n N_VGND_c_390_n 0.011782f $X=3.755 $Y=1.185 $X2=0 $Y2=0
cc_197 N_X_c_279_n N_VPWR_c_296_n 0.0322284f $X=0.465 $Y=0.42 $X2=0 $Y2=0
cc_198 N_X_M1008_s N_VPWR_c_292_n 0.00215158f $X=0.3 $Y=1.835 $X2=0 $Y2=0
cc_199 N_X_c_279_n N_VPWR_c_292_n 0.0186864f $X=0.465 $Y=0.42 $X2=0 $Y2=0
cc_200 N_X_c_279_n N_VGND_c_388_n 0.0335785f $X=0.465 $Y=0.42 $X2=0 $Y2=0
cc_201 N_X_M1001_s N_VGND_c_390_n 0.00336915f $X=0.34 $Y=0.235 $X2=0 $Y2=0
cc_202 N_X_c_279_n N_VGND_c_390_n 0.0187779f $X=0.465 $Y=0.42 $X2=0 $Y2=0
cc_203 N_VPWR_c_292_n N_A_346_367#_M1011_d 0.0041489f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_204 N_VPWR_c_292_n N_A_346_367#_M1003_d 0.00467071f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_292_n N_A_346_367#_M1006_d 0.00302127f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_298_n N_A_346_367#_c_375_n 0.0136943f $X=2.135 $Y=3.33 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_292_n N_A_346_367#_c_375_n 0.00866972f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_208 N_VPWR_M1005_d N_A_346_367#_c_348_n 0.00565231f $X=2.16 $Y=1.835 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_294_n N_A_346_367#_c_348_n 0.0447396f $X=2.3 $Y=2.11 $X2=0 $Y2=0
cc_210 N_VPWR_c_299_n N_A_346_367#_c_379_n 0.0131621f $X=3.355 $Y=3.33 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_292_n N_A_346_367#_c_379_n 0.00808656f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_212 N_VPWR_M1009_d N_A_346_367#_c_350_n 0.00218982f $X=3.36 $Y=1.835 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_295_n N_A_346_367#_c_350_n 0.017285f $X=3.52 $Y=2.11 $X2=0 $Y2=0
cc_214 N_VPWR_c_300_n N_A_346_367#_c_351_n 0.0185207f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_292_n N_A_346_367#_c_351_n 0.010808f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VGND_c_390_n A_478_47# 0.00612418f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_217 N_VGND_c_390_n A_550_47# 0.00926526f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_218 N_VGND_c_390_n A_658_47# 0.00338869f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
