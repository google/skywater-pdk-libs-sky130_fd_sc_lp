* File: sky130_fd_sc_lp__o31ai_lp.pex.spice
* Created: Wed Sep  2 10:25:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31AI_LP%A1 2 7 9 11 14 16 17 21 22 23
r37 21 23 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.275
+ $X2=0.402 $Y2=1.11
r38 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.275 $X2=0.385 $Y2=1.275
r39 16 17 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r40 16 22 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.275
r41 12 14 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.51 $Y=0.855
+ $X2=0.73 $Y2=0.855
r42 9 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.73 $Y=0.78 $X2=0.73
+ $Y2=0.855
r43 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.73 $Y=0.78 $X2=0.73
+ $Y2=0.495
r44 5 7 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.56 $Y=1.905 $X2=0.56
+ $Y2=2.595
r45 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=0.93 $X2=0.51
+ $Y2=0.855
r46 3 23 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.51 $Y=0.93 $X2=0.51
+ $Y2=1.11
r47 2 5 46.5327 $w=3.18e-07 $l=3.77829e-07 $layer=POLY_cond $X=0.402 $Y=1.598
+ $X2=0.56 $Y2=1.905
r48 1 21 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.292
+ $X2=0.402 $Y2=1.275
r49 1 2 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=0.402 $Y=1.292
+ $X2=0.402 $Y2=1.598
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_LP%A2 3 7 11 12 13 14 15 16 22 23
c49 22 0 1.32025e-19 $X=1.09 $Y=1.43
r50 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09
+ $Y=1.43 $X2=1.09 $Y2=1.43
r51 15 16 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=2.405
+ $X2=1.12 $Y2=2.775
r52 14 15 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=2.035
+ $X2=1.12 $Y2=2.405
r53 13 14 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=2.035
r54 13 23 6.94421 $w=3.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.43
r55 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.09 $Y=1.77
+ $X2=1.09 $Y2=1.43
r56 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.77
+ $X2=1.09 $Y2=1.935
r57 10 22 43.0552 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.265
+ $X2=1.09 $Y2=1.43
r58 7 10 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.16 $Y=0.495 $X2=1.16
+ $Y2=1.265
r59 3 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.05 $Y=2.595
+ $X2=1.05 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_LP%A3 3 7 11 12 13 16 17
r41 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.39 $X2=1.66 $Y2=1.39
r42 13 17 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.66 $Y=1.665
+ $X2=1.66 $Y2=1.39
r43 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.66 $Y=1.73
+ $X2=1.66 $Y2=1.39
r44 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.73
+ $X2=1.66 $Y2=1.895
r45 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.225
+ $X2=1.66 $Y2=1.39
r46 7 10 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.75 $Y=0.495
+ $X2=1.75 $Y2=1.225
r47 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.62 $Y=2.595 $X2=1.62
+ $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_LP%B1 3 7 11 12 13 16 17
r36 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.39 $X2=2.23 $Y2=1.39
r37 13 17 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=2.22 $Y2=1.39
r38 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=1.73
+ $X2=2.23 $Y2=1.39
r39 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.73
+ $X2=2.23 $Y2=1.895
r40 10 16 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.225
+ $X2=2.23 $Y2=1.39
r41 7 10 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.18 $Y=0.495
+ $X2=2.18 $Y2=1.225
r42 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.19 $Y=2.595 $X2=2.19
+ $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_LP%VPWR 1 2 7 9 13 15 17 19 32
r35 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 20 28 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r43 20 22 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 19 31 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.585 $Y2=3.33
r45 19 25 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 17 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 13 31 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.455 $Y=3.245
+ $X2=2.585 $Y2=3.33
r49 13 15 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.455 $Y=3.245
+ $X2=2.455 $Y2=2.905
r50 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.295 $Y=2.24
+ $X2=0.295 $Y2=2.95
r51 7 28 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r52 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.95
r53 2 15 600 $w=1.7e-07 $l=8.77211e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.095 $X2=2.455 $Y2=2.905
r54 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.095 $X2=0.295 $Y2=2.95
r55 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.095 $X2=0.295 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_LP%Y 1 2 9 12 16 18 19 20 25 31
r36 20 25 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=2.405
+ $X2=2.585 $Y2=2.405
r37 20 25 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.57 $Y=2.405
+ $X2=2.585 $Y2=2.405
r38 19 20 20.5435 $w=2.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.16 $Y=2.405
+ $X2=2.57 $Y2=2.405
r39 19 26 5.51168 $w=2.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.16 $Y=2.405
+ $X2=2.05 $Y2=2.405
r40 18 26 5.11717 $w=2.3e-07 $l=2.43e-07 $layer=LI1_cond $X=1.807 $Y=2.405
+ $X2=2.05 $Y2=2.405
r41 18 31 4.06913 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.807 $Y=2.405
+ $X2=1.807 $Y2=2.24
r42 14 16 5.07033 $w=4.58e-07 $l=1.95e-07 $layer=LI1_cond $X=2.475 $Y=0.495
+ $X2=2.67 $Y2=0.495
r43 12 20 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.67 $Y=2.29
+ $X2=2.67 $Y2=2.405
r44 11 16 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.67 $Y=0.725 $X2=2.67
+ $Y2=0.495
r45 11 12 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=2.67 $Y=0.725
+ $X2=2.67 $Y2=2.29
r46 7 18 2.83606 $w=4.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.807 $Y=2.52
+ $X2=1.807 $Y2=2.405
r47 7 9 9.37134 $w=4.83e-07 $l=3.8e-07 $layer=LI1_cond $X=1.807 $Y=2.52
+ $X2=1.807 $Y2=2.9
r48 2 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.095 $X2=1.885 $Y2=2.24
r49 2 9 600 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.095 $X2=1.885 $Y2=2.9
r50 1 14 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=2.255
+ $Y=0.285 $X2=2.475 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_LP%VGND 1 2 7 9 13 16 17 18 28 29
r33 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r34 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 26 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r36 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r37 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r38 23 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r39 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r40 20 32 4.48049 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.3 $Y2=0
r41 20 22 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=1.2 $Y2=0
r42 18 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r43 18 23 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r44 16 22 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.2
+ $Y2=0
r45 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.455
+ $Y2=0
r46 15 25 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.68
+ $Y2=0
r47 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.455
+ $Y2=0
r48 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=0.085
+ $X2=1.455 $Y2=0
r49 11 13 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.455 $Y=0.085
+ $X2=1.455 $Y2=0.48
r50 7 32 3.28569 $w=3.3e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.435 $Y=0.085
+ $X2=0.3 $Y2=0
r51 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.435 $Y=0.085
+ $X2=0.435 $Y2=0.495
r52 2 13 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=1.235
+ $Y=0.285 $X2=1.455 $Y2=0.48
r53 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.29
+ $Y=0.285 $X2=0.435 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_LP%A_161_57# 1 2 9 11 12 15
c35 11 0 1.32025e-19 $X=1.8 $Y=0.96
r36 13 15 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.965 $Y=0.875
+ $X2=1.965 $Y2=0.495
r37 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.8 $Y=0.96
+ $X2=1.965 $Y2=0.875
r38 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.8 $Y=0.96 $X2=1.11
+ $Y2=0.96
r39 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.945 $Y=0.875
+ $X2=1.11 $Y2=0.96
r40 7 9 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.945 $Y=0.875
+ $X2=0.945 $Y2=0.495
r41 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.285 $X2=1.965 $Y2=0.495
r42 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.805
+ $Y=0.285 $X2=0.945 $Y2=0.495
.ends

