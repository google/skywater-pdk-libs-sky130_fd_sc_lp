* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 X a_88_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_88_269# B1 a_250_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR A1 a_264_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND A3 a_250_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_250_69# B2 a_88_269# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND A1 a_250_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_358_367# A3 a_88_269# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 X a_88_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_264_367# A2 a_358_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_250_69# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_88_269# B2 a_604_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_604_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
