* File: sky130_fd_sc_lp__xor2_lp.spice
* Created: Wed Sep  2 10:41:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor2_lp.pex.spice"
.subckt sky130_fd_sc_lp__xor2_lp  VNB VPB A B X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_114_119# N_A_84_93#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1012 N_X_M1012_d N_A_84_93#_M1012_g A_114_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 A_272_119# N_B_M1000_g N_X_M1012_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75001.2 A=0.063
+ P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g A_272_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0979125 AS=0.0441 PD=1.035 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1007 A_446_68# N_B_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0979125 PD=0.66 PS=1.035 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.9 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_84_93#_M1003_d N_B_M1003_g A_446_68# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_610_68# N_A_M1008_g N_A_84_93#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g A_610_68# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_159_419#_M1004_d N_A_84_93#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.3 PD=1.28 PS=2.6 NRD=0 NRS=2.9353 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_159_419#_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1005 N_A_159_419#_M1005_d N_B_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1010 A_590_412# N_B_M1010_g N_A_84_93#_M1010_s VPB PHIGHVT L=0.25 W=1 AD=0.105
+ AS=0.285 PD=1.21 PS=2.57 NRD=9.8303 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g A_590_412# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.105 PD=2.57 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125001 SB=125000 A=0.25
+ P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__xor2_lp.pxi.spice"
*
.ends
*
*
