* File: sky130_fd_sc_lp__o311ai_1.pex.spice
* Created: Wed Sep  2 10:23:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311AI_1%A1 3 7 9 10 14
c25 10 0 7.50033e-20 $X=0.72 $Y=1.665
r26 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.7 $Y=1.51 $X2=0.7
+ $Y2=1.675
r27 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.7 $Y=1.51 $X2=0.7
+ $Y2=1.345
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.51 $X2=0.7 $Y2=1.51
r29 10 15 0.569108 $w=4.03e-07 $l=2e-08 $layer=LI1_cond $X=0.72 $Y=1.547 $X2=0.7
+ $Y2=1.547
r30 9 15 13.0895 $w=4.03e-07 $l=4.6e-07 $layer=LI1_cond $X=0.24 $Y=1.547 $X2=0.7
+ $Y2=1.547
r31 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.79 $Y=2.465
+ $X2=0.79 $Y2=1.675
r32 3 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.79 $Y=0.655
+ $X2=0.79 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%A2 3 7 9 10 11 12 18 19
c35 7 0 7.50033e-20 $X=1.23 $Y=2.465
r36 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.24 $Y=1.51
+ $X2=1.24 $Y2=1.675
r37 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.24 $Y=1.51
+ $X2=1.24 $Y2=1.345
r38 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.24
+ $Y=1.51 $X2=1.24 $Y2=1.51
r39 11 12 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=2.405
+ $X2=1.192 $Y2=2.775
r40 10 11 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=2.035
+ $X2=1.192 $Y2=2.405
r41 9 10 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=1.665
+ $X2=1.192 $Y2=2.035
r42 9 19 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=1.192 $Y=1.665
+ $X2=1.192 $Y2=1.51
r43 7 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.23 $Y=2.465
+ $X2=1.23 $Y2=1.675
r44 3 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.22 $Y=0.655
+ $X2=1.22 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%A3 3 7 9 12 13
r32 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.51
+ $X2=1.78 $Y2=1.675
r33 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.51
+ $X2=1.78 $Y2=1.345
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=1.51 $X2=1.78 $Y2=1.51
r35 9 13 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.51
r36 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=0.655
+ $X2=1.73 $Y2=1.345
r37 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.69 $Y=2.465
+ $X2=1.69 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%B1 3 7 9 15 16
r34 14 16 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.32 $Y=1.51 $X2=2.5
+ $Y2=1.51
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.51 $X2=2.32 $Y2=1.51
r36 11 14 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.23 $Y=1.51 $X2=2.32
+ $Y2=1.51
r37 9 15 4.23887 $w=4.33e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=2.32 $Y2=1.562
r38 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=1.345 $X2=2.5
+ $Y2=1.51
r39 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.5 $Y=1.345 $X2=2.5
+ $Y2=0.655
r40 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.675
+ $X2=2.23 $Y2=1.51
r41 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.23 $Y=1.675 $X2=2.23
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%C1 3 7 9 10 16
r23 13 16 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.86 $Y=1.375
+ $X2=3.09 $Y2=1.375
r24 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=1.295
+ $X2=3.105 $Y2=1.665
r25 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.375 $X2=3.09 $Y2=1.375
r26 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.86 $Y=1.54
+ $X2=2.86 $Y2=1.375
r27 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.86 $Y=1.54 $X2=2.86
+ $Y2=2.465
r28 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.86 $Y=1.21
+ $X2=2.86 $Y2=1.375
r29 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.86 $Y=1.21 $X2=2.86
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%VPWR 1 2 9 15 18 19 20 22 32 33 36
r41 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.74 $Y=3.33
+ $X2=0.575 $Y2=3.33
r46 27 29 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=0.74 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 25 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.41 $Y=3.33
+ $X2=0.575 $Y2=3.33
r50 22 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.41 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 20 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 20 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 18 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r55 17 32 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r57 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r58 13 15 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=2.395
r59 9 12 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.575 $Y=2.005
+ $X2=0.575 $Y2=2.95
r60 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.575 $Y=3.245
+ $X2=0.575 $Y2=3.33
r61 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.575 $Y=3.245
+ $X2=0.575 $Y2=2.95
r62 2 15 300 $w=1.7e-07 $l=6.69328e-07 $layer=licon1_PDIFF $count=2 $X=2.305
+ $Y=1.835 $X2=2.545 $Y2=2.395
r63 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.45
+ $Y=1.835 $X2=0.575 $Y2=2.95
r64 1 9 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.45
+ $Y=1.835 $X2=0.575 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%Y 1 2 3 10 12 17 21 24 25 26 41
r41 40 41 5.90032 $w=1.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.67 $Y=2.03
+ $X2=2.575 $Y2=2.03
r42 26 38 4.26246 $w=3.63e-07 $l=1.35e-07 $layer=LI1_cond $X=3.092 $Y=2.775
+ $X2=3.092 $Y2=2.91
r43 25 26 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.092 $Y=2.405
+ $X2=3.092 $Y2=2.775
r44 24 40 24.9545 $w=1.78e-07 $l=4.05e-07 $layer=LI1_cond $X=3.075 $Y=2.03
+ $X2=2.67 $Y2=2.03
r45 24 25 7.58733 $w=5.33e-07 $l=2.85e-07 $layer=LI1_cond $X=3.092 $Y=2.12
+ $X2=3.092 $Y2=2.405
r46 21 23 18.6775 $w=6.63e-07 $l=6.6e-07 $layer=LI1_cond $X=2.907 $Y=0.38
+ $X2=2.907 $Y2=1.04
r47 17 40 0.384081 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.67 $Y=1.94 $X2=2.67
+ $Y2=2.03
r48 17 23 52.5359 $w=1.88e-07 $l=9e-07 $layer=LI1_cond $X=2.67 $Y=1.94 $X2=2.67
+ $Y2=1.04
r49 15 19 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=2.035
+ $X2=1.96 $Y2=2.035
r50 15 41 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.125 $Y=2.035
+ $X2=2.575 $Y2=2.035
r51 10 19 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=2.12 $X2=1.96
+ $Y2=2.035
r52 10 12 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.96 $Y=2.12
+ $X2=1.96 $Y2=2.51
r53 3 24 400 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.835 $X2=3.075 $Y2=2.035
r54 3 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.835 $X2=3.075 $Y2=2.91
r55 2 19 600 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=1.835 $X2=1.96 $Y2=2.035
r56 2 12 300 $w=1.7e-07 $l=7.66322e-07 $layer=licon1_PDIFF $count=2 $X=1.765
+ $Y=1.835 $X2=1.96 $Y2=2.51
r57 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.935
+ $Y=0.235 $X2=3.075 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r36 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r39 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 21 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r42 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r43 21 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r44 19 28 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=1.2
+ $Y2=0
r45 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=1.475
+ $Y2=0
r46 18 31 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=0 $X2=1.68
+ $Y2=0
r47 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=0 $X2=1.475
+ $Y2=0
r48 16 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.24
+ $Y2=0
r49 16 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.54
+ $Y2=0
r50 15 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=1.2
+ $Y2=0
r51 15 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.54
+ $Y2=0
r52 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=0.085
+ $X2=1.475 $Y2=0
r53 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0.085
+ $X2=1.475 $Y2=0.36
r54 7 17 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.54 $Y=0.085
+ $X2=0.54 $Y2=0
r55 7 9 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.54 $Y=0.085
+ $X2=0.54 $Y2=0.38
r56 2 13 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=1.295
+ $Y=0.235 $X2=1.475 $Y2=0.36
r57 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.45
+ $Y=0.235 $X2=0.575 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_1%A_173_47# 1 2 9 11 12 15
r26 13 15 11.5587 $w=5.93e-07 $l=5.75e-07 $layer=LI1_cond $X=2.107 $Y=1.005
+ $X2=2.107 $Y2=0.43
r27 11 13 10.0057 $w=1.7e-07 $l=3.36829e-07 $layer=LI1_cond $X=1.81 $Y=1.09
+ $X2=2.107 $Y2=1.005
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.81 $Y=1.09
+ $X2=1.14 $Y2=1.09
r29 7 12 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.99 $Y=1.005
+ $X2=1.14 $Y2=1.09
r30 7 9 22.0885 $w=2.98e-07 $l=5.75e-07 $layer=LI1_cond $X=0.99 $Y=1.005
+ $X2=0.99 $Y2=0.43
r31 2 15 45.5 $w=1.7e-07 $l=5.6921e-07 $layer=licon1_NDIFF $count=4 $X=1.805
+ $Y=0.235 $X2=2.285 $Y2=0.43
r32 1 9 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=0.865
+ $Y=0.235 $X2=1.005 $Y2=0.43
.ends

