* NGSPICE file created from sky130_fd_sc_lp__nand4b_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand4b_lp A_N B C D VGND VNB VPB VPWR Y
M1000 a_173_47# a_87_231# Y VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_87_231# A_N VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=8.65e+11p ps=7.73e+06u
M1002 a_509_47# A_N VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.512e+11p ps=1.56e+06u
M1003 VPWR B Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1004 VPWR D Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_329_47# C a_251_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1006 VGND D a_329_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_87_231# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_251_47# B a_173_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_87_231# A_N a_509_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends

