# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.365000 1.805000 1.775000 2.190000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.225000 0.255000 10.465000 3.075000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 1.895000 7.635000 1.915000 ;
        RECT 3.975000 1.915000 6.085000 1.935000 ;
        RECT 3.975000 1.935000 4.305000 2.155000 ;
        RECT 4.135000 0.985000 4.825000 1.235000 ;
        RECT 4.135000 1.235000 4.305000 1.765000 ;
        RECT 4.135000 1.765000 7.635000 1.895000 ;
        RECT 5.905000 1.245000 7.635000 1.765000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.925000 0.855000 1.405000 ;
        RECT 0.545000 0.840000 0.855000 0.925000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 11.040000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 11.230000 3.520000 ;
        RECT  8.145000 1.445000  9.185000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.090000  0.410000  0.405000 0.740000 ;
      RECT  0.090000  0.740000  0.260000 1.575000 ;
      RECT  0.090000  1.575000  0.845000 1.825000 ;
      RECT  0.090000  1.825000  0.365000 2.975000 ;
      RECT  0.575000  0.085000  0.905000 0.670000 ;
      RECT  0.585000  2.315000  0.795000 3.245000 ;
      RECT  1.025000  0.840000  1.355000 1.455000 ;
      RECT  1.025000  1.455000  2.125000 1.635000 ;
      RECT  1.025000  1.635000  1.195000 2.315000 ;
      RECT  1.025000  2.315000  1.235000 2.985000 ;
      RECT  1.075000  0.415000  1.355000 0.840000 ;
      RECT  1.545000  0.085000  1.840000 0.970000 ;
      RECT  1.545000  2.360000  1.875000 3.245000 ;
      RECT  1.945000  1.635000  2.125000 1.845000 ;
      RECT  2.010000  0.640000  2.235000 1.005000 ;
      RECT  2.010000  1.005000  2.465000 1.175000 ;
      RECT  2.045000  2.095000  2.465000 2.265000 ;
      RECT  2.045000  2.265000  2.235000 2.690000 ;
      RECT  2.295000  1.175000  2.465000 2.095000 ;
      RECT  2.405000  0.615000  2.815000 0.835000 ;
      RECT  2.405000  2.435000  2.815000 2.710000 ;
      RECT  2.645000  0.835000  2.815000 1.555000 ;
      RECT  2.645000  1.555000  3.945000 1.725000 ;
      RECT  2.645000  1.725000  2.815000 2.435000 ;
      RECT  3.070000  1.015000  3.955000 1.185000 ;
      RECT  3.070000  1.185000  3.400000 1.385000 ;
      RECT  3.070000  1.895000  3.805000 2.155000 ;
      RECT  3.195000  0.085000  3.525000 0.845000 ;
      RECT  3.195000  2.360000  3.465000 3.245000 ;
      RECT  3.615000  1.355000  3.945000 1.555000 ;
      RECT  3.635000  2.155000  3.805000 2.360000 ;
      RECT  3.635000  2.360000  3.995000 2.690000 ;
      RECT  3.785000  0.280000  4.100000 0.610000 ;
      RECT  3.785000  0.610000  3.955000 1.015000 ;
      RECT  4.165000  2.360000  4.745000 3.245000 ;
      RECT  4.485000  2.105000  4.745000 2.360000 ;
      RECT  4.895000  0.085000  5.225000 0.815000 ;
      RECT  4.915000  2.105000  5.245000 2.855000 ;
      RECT  4.915000  2.855000  6.835000 3.055000 ;
      RECT  5.405000  1.205000  5.735000 1.595000 ;
      RECT  5.435000  2.170000  5.710000 2.515000 ;
      RECT  5.435000  2.515000  7.385000 2.685000 ;
      RECT  5.785000  0.255000  6.115000 0.865000 ;
      RECT  5.785000  0.865000  8.535000 1.035000 ;
      RECT  5.925000  2.105000  8.195000 2.265000 ;
      RECT  5.925000  2.265000  6.350000 2.345000 ;
      RECT  6.255000  2.095000  8.195000 2.105000 ;
      RECT  7.030000  0.085000  7.360000 0.665000 ;
      RECT  7.055000  2.435000  7.385000 2.515000 ;
      RECT  7.555000  2.435000  7.785000 3.245000 ;
      RECT  7.625000  0.445000  9.065000 0.615000 ;
      RECT  7.625000  0.615000  7.955000 0.695000 ;
      RECT  7.955000  2.265000  8.195000 2.690000 ;
      RECT  7.975000  1.035000  8.535000 1.465000 ;
      RECT  7.975000  1.465000  8.195000 2.095000 ;
      RECT  8.285000  0.795000  8.535000 0.865000 ;
      RECT  8.365000  1.670000  8.565000 3.245000 ;
      RECT  8.735000  0.615000  9.065000 3.075000 ;
      RECT  9.235000  0.255000  9.515000 1.185000 ;
      RECT  9.235000  1.185000 10.055000 1.515000 ;
      RECT  9.235000  1.515000  9.505000 2.635000 ;
      RECT  9.685000  0.085000 10.055000 0.545000 ;
      RECT  9.725000  1.975000  9.935000 3.245000 ;
      RECT  9.745000  0.545000 10.055000 1.015000 ;
      RECT 10.635000  0.085000 10.935000 1.095000 ;
      RECT 10.635000  1.815000 10.935000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.210000  1.285000 1.380000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.210000  5.605000 1.380000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
    LAYER met1 ;
      RECT 1.055000 1.180000 1.345000 1.225000 ;
      RECT 1.055000 1.225000 5.665000 1.365000 ;
      RECT 1.055000 1.365000 1.345000 1.410000 ;
      RECT 5.375000 1.180000 5.665000 1.225000 ;
      RECT 5.375000 1.365000 5.665000 1.410000 ;
  END
END sky130_fd_sc_lp__dfstp_2
END LIBRARY
