* NGSPICE file created from sky130_fd_sc_lp__o211a_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o211a_lp A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_606_47# a_232_419# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.045e+11p ps=3.13e+06u
M1001 X a_232_419# a_606_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1002 a_27_144# A2 VGND VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1003 a_232_419# A2 a_134_419# VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=2.4e+11p ps=2.48e+06u
M1004 X a_232_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=9.6e+11p ps=7.92e+06u
M1005 a_232_419# C1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_232_419# C1 a_318_144# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1007 VPWR B1 a_232_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_318_144# B1 a_27_144# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_134_419# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_27_144# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

