* File: sky130_fd_sc_lp__buflp_2.spice
* Created: Fri Aug 28 10:12:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buflp_2.pex.spice"
.subckt sky130_fd_sc_lp__buflp_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_98_21#_M1003_g N_A_128_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2982 AS=0.1176 PD=2.39 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6
+ SA=75000.3 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1005 N_A_128_47#_M1003_s N_A_98_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.7
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1006 N_A_128_47#_M1006_d N_A_98_21#_M1006_g N_X_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A_98_21#_M1007_g N_A_128_47#_M1006_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1708 AS=0.147 PD=1.6 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 A_516_47# N_A_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0854 PD=0.63 PS=0.8 NRD=14.28 NRS=2.856 M=1 R=2.8 SA=75002.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_98_21#_M1010_d N_A_M1010_g A_516_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_128_367#_M1001_d N_A_98_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4473 PD=1.54 PS=3.23 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75000.3 SB=75002 A=0.189 P=2.82 MULT=1
MM1000 N_A_128_367#_M1001_d N_A_98_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1004 N_A_128_367#_M1004_d N_A_98_21#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1009 N_A_128_367#_M1004_d N_A_98_21#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.343317 PD=1.54 PS=2.28789 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75001.6 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1002 A_509_377# N_A_M1002_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.174383 PD=0.88 PS=1.16211 NRD=19.9955 NRS=36.1495 M=1 R=4.26667
+ SA=75002.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_98_21#_M1011_d N_A_M1011_g A_509_377# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75002.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__buflp_2.pxi.spice"
*
.ends
*
*
