* File: sky130_fd_sc_lp__maj3_4.pex.spice
* Created: Wed Sep  2 09:59:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MAJ3_4%C 3 6 10 14 17 18 19 21 25 26 28 31 33 42
c89 26 0 1.9317e-19 $X=2.815 $Y=1.44
c90 14 0 2.76993e-19 $X=2.725 $Y=2.465
r91 31 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.35
+ $X2=0.605 $Y2=1.515
r92 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.35
+ $X2=0.605 $Y2=1.185
r93 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.35 $X2=0.605 $Y2=1.35
r94 28 42 3.44013 $w=3.33e-07 $l=1e-07 $layer=LI1_cond $X=0.72 $Y=1.347 $X2=0.82
+ $Y2=1.347
r95 28 32 3.95615 $w=3.33e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.347
+ $X2=0.605 $Y2=1.347
r96 26 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.44
+ $X2=2.815 $Y2=1.605
r97 26 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.44
+ $X2=2.815 $Y2=1.275
r98 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.815
+ $Y=1.44 $X2=2.815 $Y2=1.44
r99 22 25 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.57 $Y=1.44
+ $X2=2.815 $Y2=1.44
r100 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=1.605
+ $X2=2.57 $Y2=1.44
r101 20 21 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.57 $Y=1.605
+ $X2=2.57 $Y2=2.225
r102 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.485 $Y=2.31
+ $X2=2.57 $Y2=2.225
r103 18 19 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=2.485 $Y=2.31
+ $X2=0.905 $Y2=2.31
r104 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.82 $Y=2.225
+ $X2=0.905 $Y2=2.31
r105 16 42 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.82 $Y=1.515
+ $X2=0.82 $Y2=1.347
r106 16 17 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.82 $Y=1.515
+ $X2=0.82 $Y2=2.225
r107 14 37 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.725 $Y=2.465
+ $X2=2.725 $Y2=1.605
r108 10 36 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.725 $Y=0.655
+ $X2=2.725 $Y2=1.275
r109 6 34 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.695 $Y=2.465
+ $X2=0.695 $Y2=1.515
r110 3 33 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.695 $Y=0.655
+ $X2=0.695 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_4%A 1 3 6 8 10 13 15 16 24
r45 22 24 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.25 $Y=1.35
+ $X2=1.515 $Y2=1.35
r46 19 22 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.35
+ $X2=1.25 $Y2=1.35
r47 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.25 $Y=1.295
+ $X2=1.25 $Y2=1.665
r48 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.35 $X2=1.25 $Y2=1.35
r49 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.515
+ $X2=1.515 $Y2=1.35
r50 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.515 $Y=1.515
+ $X2=1.515 $Y2=2.465
r51 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.185
+ $X2=1.515 $Y2=1.35
r52 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.515 $Y=1.185
+ $X2=1.515 $Y2=0.655
r53 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.515
+ $X2=1.085 $Y2=1.35
r54 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.085 $Y=1.515
+ $X2=1.085 $Y2=2.465
r55 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.185
+ $X2=1.085 $Y2=1.35
r56 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.085 $Y=1.185
+ $X2=1.085 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_4%B 1 3 6 8 10 13 15 22
c44 15 0 1.9317e-19 $X=2.16 $Y=1.295
r45 20 22 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.14 $Y=1.35
+ $X2=2.335 $Y2=1.35
r46 17 20 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.905 $Y=1.35
+ $X2=2.14 $Y2=1.35
r47 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.35 $X2=2.14 $Y2=1.35
r48 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.515
+ $X2=2.335 $Y2=1.35
r49 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.335 $Y=1.515
+ $X2=2.335 $Y2=2.465
r50 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.185
+ $X2=2.335 $Y2=1.35
r51 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.335 $Y=1.185
+ $X2=2.335 $Y2=0.655
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.515
+ $X2=1.905 $Y2=1.35
r53 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.905 $Y=1.515
+ $X2=1.905 $Y2=2.465
r54 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.185
+ $X2=1.905 $Y2=1.35
r55 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.905 $Y=1.185
+ $X2=1.905 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_4%A_65_367# 1 2 3 4 15 19 23 27 31 35 39 43 49
+ 53 55 56 58 59 61 65 67 68 70 71 76 83 84 96
c165 61 0 1.98867e-19 $X=2.12 $Y=1.96
c166 19 0 1.6164e-19 $X=3.38 $Y=0.655
r167 93 94 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.275 $Y=1.44
+ $X2=4.315 $Y2=1.44
r168 92 93 81.3105 $w=3.3e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.44
+ $X2=4.275 $Y2=1.44
r169 91 92 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=3.725 $Y=1.44
+ $X2=3.81 $Y2=1.44
r170 87 89 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=3.295 $Y=1.44
+ $X2=3.38 $Y2=1.44
r171 83 84 9.30866 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.322 $Y=1.96
+ $X2=0.322 $Y2=1.795
r172 77 96 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.505 $Y=1.44
+ $X2=4.745 $Y2=1.44
r173 77 94 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.505 $Y=1.44
+ $X2=4.315 $Y2=1.44
r174 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.505
+ $Y=1.44 $X2=4.505 $Y2=1.44
r175 74 91 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.485 $Y=1.44
+ $X2=3.725 $Y2=1.44
r176 74 89 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=3.485 $Y=1.44
+ $X2=3.38 $Y2=1.44
r177 73 76 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.485 $Y=1.44
+ $X2=4.505 $Y2=1.44
r178 73 74 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.485
+ $Y=1.44 $X2=3.485 $Y2=1.44
r179 71 73 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.33 $Y=1.44
+ $X2=3.485 $Y2=1.44
r180 70 71 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.245 $Y=1.275
+ $X2=3.33 $Y2=1.44
r181 69 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.245 $Y=1
+ $X2=3.245 $Y2=1.275
r182 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.16 $Y=0.915
+ $X2=3.245 $Y2=1
r183 67 68 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.16 $Y=0.915
+ $X2=2.285 $Y2=0.915
r184 63 68 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=0.915
+ $X2=2.285 $Y2=0.915
r185 63 85 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.12 $Y=0.915
+ $X2=1.71 $Y2=0.915
r186 63 65 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.12 $Y=0.83
+ $X2=2.12 $Y2=0.38
r187 59 61 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.795 $Y=1.92
+ $X2=2.12 $Y2=1.92
r188 58 59 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.71 $Y=1.795
+ $X2=1.795 $Y2=1.92
r189 57 85 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1 $X2=1.71
+ $Y2=0.915
r190 57 58 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.71 $Y=1 $X2=1.71
+ $Y2=1.795
r191 55 85 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=0.915
+ $X2=1.71 $Y2=0.915
r192 55 56 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=1.625 $Y=0.915
+ $X2=0.645 $Y2=0.915
r193 51 56 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.48 $Y=0.915
+ $X2=0.645 $Y2=0.915
r194 51 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.48 $Y=0.915
+ $X2=0.175 $Y2=0.915
r195 51 53 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.48 $Y=0.83 $X2=0.48
+ $Y2=0.43
r196 47 83 1.72338 $w=4.63e-07 $l=6.7e-08 $layer=LI1_cond $X=0.322 $Y=2.027
+ $X2=0.322 $Y2=1.96
r197 47 49 22.4554 $w=4.63e-07 $l=8.73e-07 $layer=LI1_cond $X=0.322 $Y=2.027
+ $X2=0.322 $Y2=2.9
r198 45 79 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=1
+ $X2=0.175 $Y2=0.915
r199 45 84 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.175 $Y=1
+ $X2=0.175 $Y2=1.795
r200 41 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.605
+ $X2=4.745 $Y2=1.44
r201 41 43 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.745 $Y=1.605
+ $X2=4.745 $Y2=2.465
r202 37 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.275
+ $X2=4.745 $Y2=1.44
r203 37 39 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.745 $Y=1.275
+ $X2=4.745 $Y2=0.655
r204 33 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.605
+ $X2=4.315 $Y2=1.44
r205 33 35 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.315 $Y=1.605
+ $X2=4.315 $Y2=2.465
r206 29 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.275 $Y=1.275
+ $X2=4.275 $Y2=1.44
r207 29 31 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.275 $Y=1.275
+ $X2=4.275 $Y2=0.655
r208 25 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.275
+ $X2=3.81 $Y2=1.44
r209 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.81 $Y=1.275
+ $X2=3.81 $Y2=0.655
r210 21 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.725 $Y=1.605
+ $X2=3.725 $Y2=1.44
r211 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.725 $Y=1.605
+ $X2=3.725 $Y2=2.465
r212 17 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.275
+ $X2=3.38 $Y2=1.44
r213 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.38 $Y=1.275
+ $X2=3.38 $Y2=0.655
r214 13 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.605
+ $X2=3.295 $Y2=1.44
r215 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.295 $Y=1.605
+ $X2=3.295 $Y2=2.465
r216 4 61 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.835 $X2=2.12 $Y2=1.96
r217 3 83 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.47 $Y2=1.96
r218 3 49 400 $w=1.7e-07 $l=1.13519e-06 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.47 $Y2=2.9
r219 2 65 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.98
+ $Y=0.235 $X2=2.12 $Y2=0.38
r220 1 53 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=0.335
+ $Y=0.235 $X2=0.48 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_4%VPWR 1 2 3 4 15 19 25 27 29 32 33 34 36 48 52
+ 58 61 65
r67 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r68 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r69 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r70 56 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r71 56 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r72 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r73 53 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.02 $Y2=3.33
r74 53 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 52 64 3.96406 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=5.077 $Y2=3.33
r76 52 55 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 48 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.02 $Y2=3.33
r80 48 50 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r81 44 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r82 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r83 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 41 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.3 $Y2=3.33
r85 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.68 $Y2=3.33
r86 39 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r87 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=1.3 $Y2=3.33
r89 36 38 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 34 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r91 34 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 34 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 32 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33 $X2=3
+ $Y2=3.33
r95 31 50 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r96 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33 $X2=3
+ $Y2=3.33
r97 27 64 3.1791 $w=2.5e-07 $l=1.17346e-07 $layer=LI1_cond $X=5 $Y=3.245
+ $X2=5.077 $Y2=3.33
r98 27 29 43.5623 $w=2.48e-07 $l=9.45e-07 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=2.3
r99 23 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=3.33
r100 23 25 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=2.3
r101 19 22 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=3 $Y=1.96 $X2=3
+ $Y2=2.93
r102 17 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=3.33
r103 17 22 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.93
r104 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=3.245 $X2=1.3
+ $Y2=3.33
r105 13 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.3 $Y=3.245
+ $X2=1.3 $Y2=2.835
r106 4 29 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=2.3
r107 3 25 300 $w=1.7e-07 $l=5.6438e-07 $layer=licon1_PDIFF $count=2 $X=3.8
+ $Y=1.835 $X2=4.02 $Y2=2.3
r108 2 22 400 $w=1.7e-07 $l=1.19081e-06 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.835 $X2=3 $Y2=2.93
r109 2 19 400 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.835 $X2=3 $Y2=1.96
r110 1 15 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.835 $X2=1.3 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_4%X 1 2 3 4 15 21 23 24 25 26 29 33 37 39 41 42
+ 45 46
c67 26 0 1.6164e-19 $X=3.68 $Y=1.01
c68 24 0 7.81255e-20 $X=3.675 $Y=1.87
r69 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.665
r70 44 46 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.04 $Y=1.785
+ $X2=5.04 $Y2=1.665
r71 43 45 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=5.04 $Y=1.095 $X2=5.04
+ $Y2=1.295
r72 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.695 $Y=1.87
+ $X2=4.53 $Y2=1.87
r73 39 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.925 $Y=1.87
+ $X2=5.04 $Y2=1.785
r74 39 40 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.925 $Y=1.87
+ $X2=4.695 $Y2=1.87
r75 38 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=1.01
+ $X2=4.49 $Y2=1.01
r76 37 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.925 $Y=1.01
+ $X2=5.04 $Y2=1.095
r77 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.925 $Y=1.01
+ $X2=4.655 $Y2=1.01
r78 33 35 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=4.53 $Y=1.96
+ $X2=4.53 $Y2=2.9
r79 31 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=1.955
+ $X2=4.53 $Y2=1.87
r80 31 33 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=4.53 $Y=1.955
+ $X2=4.53 $Y2=1.96
r81 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.925
+ $X2=4.49 $Y2=1.01
r82 27 29 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.49 $Y=0.925
+ $X2=4.49 $Y2=0.43
r83 25 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=1.01
+ $X2=4.49 $Y2=1.01
r84 25 26 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.325 $Y=1.01
+ $X2=3.68 $Y2=1.01
r85 23 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=1.87
+ $X2=4.53 $Y2=1.87
r86 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.365 $Y=1.87
+ $X2=3.675 $Y2=1.87
r87 19 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.595 $Y=0.925
+ $X2=3.68 $Y2=1.01
r88 19 21 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.595 $Y=0.925
+ $X2=3.595 $Y2=0.43
r89 15 17 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=3.51 $Y=1.96
+ $X2=3.51 $Y2=2.9
r90 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.51 $Y=1.955
+ $X2=3.675 $Y2=1.87
r91 13 15 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.51 $Y=1.955
+ $X2=3.51 $Y2=1.96
r92 4 35 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.835 $X2=4.53 $Y2=2.9
r93 4 33 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.835 $X2=4.53 $Y2=1.96
r94 3 17 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=2.9
r95 3 15 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=1.835 $X2=3.51 $Y2=1.96
r96 2 29 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=4.35
+ $Y=0.235 $X2=4.49 $Y2=0.43
r97 1 21 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.235 $X2=3.595 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_4%VGND 1 2 3 4 15 19 23 25 27 30 31 33 34 35 37
+ 52 57 61
r75 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r76 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r77 55 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r78 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r79 52 60 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5.057
+ $Y2=0
r80 52 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.56
+ $Y2=0
r81 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r82 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r83 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r84 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r85 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r86 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.3
+ $Y2=0
r87 42 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.68
+ $Y2=0
r88 40 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r89 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r90 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.3
+ $Y2=0
r91 37 39 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.24
+ $Y2=0
r92 35 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r93 35 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r94 35 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r95 33 50 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.86 $Y=0 $X2=3.6
+ $Y2=0
r96 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.86 $Y=0 $X2=3.985
+ $Y2=0
r97 32 54 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=4.56
+ $Y2=0
r98 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=3.985
+ $Y2=0
r99 30 47 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.64
+ $Y2=0
r100 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.94
+ $Y2=0
r101 29 50 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.6
+ $Y2=0
r102 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.94
+ $Y2=0
r103 25 60 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5 $Y=0.085
+ $X2=5.057 $Y2=0
r104 25 27 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.48
r105 21 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=0.085
+ $X2=3.985 $Y2=0
r106 21 23 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=3.985 $Y=0.085
+ $X2=3.985 $Y2=0.48
r107 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0
r108 17 19 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.43
r109 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0.085 $X2=1.3
+ $Y2=0
r110 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.3 $Y=0.085
+ $X2=1.3 $Y2=0.43
r111 4 27 182 $w=1.7e-07 $l=3.22684e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.235 $X2=5 $Y2=0.48
r112 3 23 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.025 $Y2=0.48
r113 2 19 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.94 $Y2=0.43
r114 1 15 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.235 $X2=1.3 $Y2=0.43
.ends

