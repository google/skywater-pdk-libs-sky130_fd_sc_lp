* NGSPICE file created from sky130_fd_sc_lp__and2b_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and2b_m A_N B VGND VNB VPB VPWR X
M1000 VPWR A_N a_35_70# VPB phighvt w=420000u l=150000u
+  ad=3.99e+11p pd=3.58e+06u as=1.113e+11p ps=1.37e+06u
M1001 X a_255_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1002 a_338_47# a_35_70# a_255_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1003 VPWR B a_255_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1004 X a_255_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.289e+11p ps=2.77e+06u
M1005 VGND B a_338_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_255_47# a_35_70# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_35_70# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

