* File: sky130_fd_sc_lp__o31a_2.spice
* Created: Fri Aug 28 11:15:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31a_2.pex.spice"
.subckt sky130_fd_sc_lp__o31a_2  VNB VPB A1 A2 A3 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_85_21#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A_85_21#_M1011_g N_X_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1007 N_A_355_47#_M1007_d N_A1_M1007_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.2604 PD=1.2 PS=1.46 NRD=1.428 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_355_47#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.9
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_A_355_47#_M1004_d N_A3_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1003 N_A_85_21#_M1003_d N_B1_M1003_g N_A_355_47#_M1004_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.147 PD=2.21 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_85_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_85_21#_M1008_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.36855 AS=0.1764 PD=1.845 PS=1.54 NRD=14.0658 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1001 A_355_367# N_A1_M1001_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.36855 PD=1.47 PS=1.845 NRD=7.8012 NRS=33.6082 M=1 R=8.4
+ SA=75001.4 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1006 A_427_367# N_A2_M1006_g A_355_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75001.7
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1005 N_A_85_21#_M1005_d N_A3_M1005_g A_427_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=9.3772 NRS=21.8867 M=1 R=8.4
+ SA=75002.3 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g N_A_85_21#_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3654 AS=0.2457 PD=3.1 PS=1.65 NRD=3.9006 NRS=7.8012 M=1 R=8.4 SA=75002.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o31a_2.pxi.spice"
*
.ends
*
*
