* File: sky130_fd_sc_lp__a32oi_lp.pex.spice
* Created: Fri Aug 28 10:02:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32OI_LP%B2 3 5 7 11 12 13 17
c39 12 0 6.50813e-20 $X=0.72 $Y=1.295
c40 7 0 1.0851e-19 $X=0.69 $Y=2.545
c41 3 0 5.59169e-20 $X=0.625 $Y=0.445
r42 12 13 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.69 $Y=1.285
+ $X2=0.69 $Y2=1.665
r43 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.285 $X2=0.69 $Y2=1.285
r44 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.69 $Y=1.625
+ $X2=0.69 $Y2=1.285
r45 10 17 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.69 $Y=1.12
+ $X2=0.69 $Y2=1.285
r46 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.69 $Y=1.79
+ $X2=0.69 $Y2=1.625
r47 5 7 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.69 $Y=1.79 $X2=0.69
+ $Y2=2.545
r48 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.625 $Y=0.445
+ $X2=0.625 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%B1 1 3 8 12 15 16 17 18 19 23
c59 18 0 5.59169e-20 $X=1.2 $Y=1.295
c60 8 0 6.50813e-20 $X=1.22 $Y=2.545
r61 18 19 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.23 $Y=1.275
+ $X2=1.23 $Y2=1.665
r62 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=1.275 $X2=1.23 $Y2=1.275
r63 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.23 $Y=1.615
+ $X2=1.23 $Y2=1.275
r64 16 17 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.615
+ $X2=1.23 $Y2=1.78
r65 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.11
+ $X2=1.23 $Y2=1.275
r66 10 12 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.015 $Y=0.805
+ $X2=1.14 $Y2=0.805
r67 8 17 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.22 $Y=2.545
+ $X2=1.22 $Y2=1.78
r68 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.14 $Y=0.88 $X2=1.14
+ $Y2=0.805
r69 4 15 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.14 $Y=0.88 $X2=1.14
+ $Y2=1.11
r70 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.015 $Y=0.73
+ $X2=1.015 $Y2=0.805
r71 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.015 $Y=0.73 $X2=1.015
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%A1 3 7 9 10 11 12 13 14 15 21
c54 21 0 2.64121e-20 $X=1.77 $Y=0.93
c55 11 0 2.73563e-19 $X=1.77 $Y=1.435
c56 9 0 1.8299e-20 $X=1.77 $Y=0.765
c57 3 0 6.83464e-20 $X=1.75 $Y=2.545
r58 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=0.93 $X2=1.77 $Y2=0.93
r59 14 15 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.755 $Y=1.295
+ $X2=1.755 $Y2=1.665
r60 14 22 11.6845 $w=3.58e-07 $l=3.65e-07 $layer=LI1_cond $X=1.755 $Y=1.295
+ $X2=1.755 $Y2=0.93
r61 13 22 0.160062 $w=3.58e-07 $l=5e-09 $layer=LI1_cond $X=1.755 $Y=0.925
+ $X2=1.755 $Y2=0.93
r62 12 13 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.755 $Y=0.555
+ $X2=1.755 $Y2=0.925
r63 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.77 $Y=1.27
+ $X2=1.77 $Y2=0.93
r64 10 11 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.27
+ $X2=1.77 $Y2=1.435
r65 9 21 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=0.765
+ $X2=1.77 $Y2=0.93
r66 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.71 $Y=0.445 $X2=1.71
+ $Y2=0.765
r67 3 11 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.75 $Y=2.545
+ $X2=1.75 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%A2 3 7 9 12
c34 3 0 4.93603e-20 $X=2.28 $Y=2.545
r35 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.615
+ $X2=2.31 $Y2=1.78
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.615
+ $X2=2.31 $Y2=1.45
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.615 $X2=2.31 $Y2=1.615
r38 9 13 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=2.31 $Y2=1.615
r39 7 14 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=1.45
r40 3 15 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.28 $Y=2.545
+ $X2=2.28 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%A3 3 7 9 10 14
r26 14 17 31.8314 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=0.975
+ $X2=2.75 $Y2=1.14
r27 14 16 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=0.975
+ $X2=2.75 $Y2=0.81
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.73
+ $Y=0.975 $X2=2.73 $Y2=0.975
r29 10 15 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.12 $Y=0.975
+ $X2=2.73 $Y2=0.975
r30 9 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=0.975 $X2=2.73
+ $Y2=0.975
r31 7 17 349.077 $w=2.5e-07 $l=1.405e-06 $layer=POLY_cond $X=2.81 $Y=2.545
+ $X2=2.81 $Y2=1.14
r32 3 16 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.64 $Y=0.445
+ $X2=2.64 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%A_56_409# 1 2 3 12 14 15 17 19 20 21 24
c57 21 0 1.84788e-19 $X=1.65 $Y=2.045
c58 20 0 1.97286e-19 $X=2.38 $Y=2.045
c59 17 0 4.93603e-20 $X=1.485 $Y=2.895
r60 24 26 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.545 $Y=2.19
+ $X2=2.545 $Y2=2.9
r61 22 24 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=2.545 $Y=2.13
+ $X2=2.545 $Y2=2.19
r62 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.38 $Y=2.045
+ $X2=2.545 $Y2=2.13
r63 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.38 $Y=2.045
+ $X2=1.65 $Y2=2.045
r64 17 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=2.895
+ $X2=1.485 $Y2=2.98
r65 17 19 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.485 $Y=2.895
+ $X2=1.485 $Y2=2.19
r66 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.485 $Y=2.13
+ $X2=1.65 $Y2=2.045
r67 16 19 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.485 $Y=2.13
+ $X2=1.485 $Y2=2.19
r68 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=2.98
+ $X2=1.485 $Y2=2.98
r69 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.32 $Y=2.98
+ $X2=0.59 $Y2=2.98
r70 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.425 $Y=2.895
+ $X2=0.59 $Y2=2.98
r71 10 12 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.425 $Y=2.895
+ $X2=0.425 $Y2=2.485
r72 3 26 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=2.045 $X2=2.545 $Y2=2.9
r73 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=2.045 $X2=2.545 $Y2=2.19
r74 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=2.045 $X2=1.485 $Y2=2.9
r75 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=2.045 $X2=1.485 $Y2=2.19
r76 1 12 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=2.045 $X2=0.425 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%Y 1 2 7 9 10 13 17 20 21 22 27
c54 9 0 6.83464e-20 $X=0.79 $Y=2.055
c55 7 0 1.8299e-20 $X=1.065 $Y=0.845
r56 21 22 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r57 20 27 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=0.845
+ $X2=0.235 $Y2=0.93
r58 20 21 17.0247 $w=2.18e-07 $l=3.25e-07 $layer=LI1_cond $X=0.235 $Y=0.97
+ $X2=0.235 $Y2=1.295
r59 20 27 2.09535 $w=2.18e-07 $l=4e-08 $layer=LI1_cond $X=0.235 $Y=0.97
+ $X2=0.235 $Y2=0.93
r60 19 22 15.9771 $w=2.18e-07 $l=3.05e-07 $layer=LI1_cond $X=0.235 $Y=1.97
+ $X2=0.235 $Y2=1.665
r61 15 17 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.23 $Y=0.76
+ $X2=1.23 $Y2=0.47
r62 11 13 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.955 $Y=2.14
+ $X2=0.955 $Y2=2.19
r63 10 19 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.345 $Y=2.055
+ $X2=0.235 $Y2=1.97
r64 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.79 $Y=2.055
+ $X2=0.955 $Y2=2.14
r65 9 10 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.79 $Y=2.055
+ $X2=0.345 $Y2=2.055
r66 8 20 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.345 $Y=0.845
+ $X2=0.235 $Y2=0.845
r67 7 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.065 $Y=0.845
+ $X2=1.23 $Y2=0.76
r68 7 8 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.065 $Y=0.845
+ $X2=0.345 $Y2=0.845
r69 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.815
+ $Y=2.045 $X2=0.955 $Y2=2.19
r70 1 17 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%VPWR 1 2 9 11 13 18 19 20 29 35
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 29 34 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=3.175 $Y2=3.33
r42 29 31 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 23 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 20 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 20 24 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 20 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 18 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=2.015 $Y2=3.33
r50 17 31 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=3.33
+ $X2=2.015 $Y2=3.33
r52 13 16 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=3.115 $Y=2.19
+ $X2=3.115 $Y2=2.9
r53 11 34 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.115 $Y=3.245
+ $X2=3.175 $Y2=3.33
r54 11 16 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=3.115 $Y=3.245
+ $X2=3.115 $Y2=2.9
r55 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=3.245
+ $X2=2.015 $Y2=3.33
r56 7 9 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.015 $Y=3.245
+ $X2=2.015 $Y2=2.475
r57 2 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=2.045 $X2=3.075 $Y2=2.9
r58 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=2.045 $X2=3.075 $Y2=2.19
r59 1 9 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=1.875
+ $Y=2.045 $X2=2.015 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_LP%VGND 1 2 7 9 13 16 17 18 28 29
c41 29 0 2.64121e-20 $X=3.12 $Y=0
r42 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 26 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r45 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r47 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r48 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 20 32 4.50939 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.287
+ $Y2=0
r50 20 22 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.72
+ $Y2=0
r51 18 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r52 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r53 16 25 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.64
+ $Y2=0
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.855
+ $Y2=0
r55 15 28 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.12
+ $Y2=0
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.855
+ $Y2=0
r57 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r58 11 13 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.42
r59 7 32 3.25678 $w=3.3e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.41 $Y=0.085
+ $X2=0.287 $Y2=0
r60 7 9 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.41 $Y=0.085 $X2=0.41
+ $Y2=0.395
r61 2 13 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.855 $Y2=0.42
r62 1 9 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.265
+ $Y=0.235 $X2=0.41 $Y2=0.395
.ends

