* File: sky130_fd_sc_lp__and2b_m.spice
* Created: Fri Aug 28 10:05:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2b_m.pex.spice"
.subckt sky130_fd_sc_lp__and2b_m  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_N_M1007_g N_A_35_70#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_338_47# N_A_35_70#_M1002_g N_A_255_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g A_338_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_255_47#_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_35_70#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 N_A_255_47#_M1006_d N_A_35_70#_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=42.1974 M=1 R=2.8
+ SA=75000.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_255_47#_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0588 PD=0.98 PS=0.7 NRD=121.943 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_255_47#_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.1176 PD=1.37 PS=0.98 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__and2b_m.pxi.spice"
*
.ends
*
*
