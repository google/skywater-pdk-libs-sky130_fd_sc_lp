* File: sky130_fd_sc_lp__a31oi_m.pxi.spice
* Created: Fri Aug 28 10:00:34 2020
* 
x_PM_SKY130_FD_SC_LP__A31OI_M%A3 N_A3_c_63_n N_A3_c_64_n N_A3_c_65_n N_A3_c_71_n
+ N_A3_c_72_n N_A3_c_73_n N_A3_M1007_g N_A3_c_66_n N_A3_M1006_g N_A3_c_67_n A3
+ A3 A3 A3 A3 N_A3_c_69_n PM_SKY130_FD_SC_LP__A31OI_M%A3
x_PM_SKY130_FD_SC_LP__A31OI_M%A2 N_A2_M1003_g N_A2_M1004_g N_A2_c_100_n
+ N_A2_c_105_n A2 A2 A2 A2 A2 N_A2_c_102_n PM_SKY130_FD_SC_LP__A31OI_M%A2
x_PM_SKY130_FD_SC_LP__A31OI_M%A1 N_A1_M1005_g N_A1_M1000_g N_A1_c_144_n
+ N_A1_c_149_n A1 A1 A1 A1 A1 N_A1_c_146_n PM_SKY130_FD_SC_LP__A31OI_M%A1
x_PM_SKY130_FD_SC_LP__A31OI_M%B1 N_B1_c_198_n N_B1_M1001_g N_B1_c_199_n
+ N_B1_M1002_g N_B1_c_200_n N_B1_c_195_n N_B1_c_202_n B1 B1 B1 N_B1_c_197_n
+ PM_SKY130_FD_SC_LP__A31OI_M%B1
x_PM_SKY130_FD_SC_LP__A31OI_M%VPWR N_VPWR_M1007_s N_VPWR_M1003_d N_VPWR_c_244_n
+ N_VPWR_c_245_n N_VPWR_c_246_n N_VPWR_c_247_n N_VPWR_c_248_n N_VPWR_c_249_n
+ VPWR N_VPWR_c_250_n N_VPWR_c_243_n PM_SKY130_FD_SC_LP__A31OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A31OI_M%A_169_500# N_A_169_500#_M1007_d
+ N_A_169_500#_M1000_d N_A_169_500#_c_290_n N_A_169_500#_c_277_n
+ N_A_169_500#_c_278_n N_A_169_500#_c_295_n
+ PM_SKY130_FD_SC_LP__A31OI_M%A_169_500#
x_PM_SKY130_FD_SC_LP__A31OI_M%Y N_Y_M1005_d N_Y_M1001_d N_Y_c_305_n N_Y_c_302_n
+ N_Y_c_299_n N_Y_c_300_n Y PM_SKY130_FD_SC_LP__A31OI_M%Y
x_PM_SKY130_FD_SC_LP__A31OI_M%VGND N_VGND_M1006_s N_VGND_M1002_d N_VGND_c_332_n
+ N_VGND_c_333_n N_VGND_c_334_n VGND N_VGND_c_335_n N_VGND_c_336_n
+ N_VGND_c_337_n N_VGND_c_338_n PM_SKY130_FD_SC_LP__A31OI_M%VGND
cc_1 VNB N_A3_c_63_n 0.00316927f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.24
cc_2 VNB N_A3_c_64_n 0.0456239f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.015
cc_3 VNB N_A3_c_65_n 0.0264706f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.015
cc_4 VNB N_A3_c_66_n 0.0185413f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=0.94
cc_5 VNB N_A3_c_67_n 0.0253241f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_6 VNB A3 0.0103629f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_A3_c_69_n 0.0388328f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_8 VNB N_A2_M1004_g 0.0351582f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.39
cc_9 VNB N_A2_c_100_n 0.0126902f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=0.62
cc_10 VNB A2 0.00792552f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.09
cc_11 VNB N_A2_c_102_n 0.020439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1005_g 0.0381837f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.015
cc_13 VNB N_A1_c_144_n 0.0108513f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=0.62
cc_14 VNB A1 0.00476924f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.09
cc_15 VNB N_A1_c_146_n 0.0185306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_M1002_g 0.0387833f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.71
cc_17 VNB N_B1_c_195_n 0.0211577f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_18 VNB B1 0.00157892f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_B1_c_197_n 0.0184035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_243_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_21 VNB N_Y_c_299_n 0.0184635f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_22 VNB N_Y_c_300_n 0.00591456f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_23 VNB Y 0.0310039f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_24 VNB N_VGND_c_332_n 0.0233004f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.71
cc_25 VNB N_VGND_c_333_n 0.0146092f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=0.62
cc_26 VNB N_VGND_c_334_n 0.0231892f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.09
cc_27 VNB N_VGND_c_335_n 0.0177361f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_VGND_c_336_n 0.0453356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_337_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_338_n 0.215501f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_31 VPB N_A3_c_63_n 0.0401529f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.24
cc_32 VPB N_A3_c_71_n 0.0360863f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.315
cc_33 VPB N_A3_c_72_n 0.0119234f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.315
cc_34 VPB N_A3_c_73_n 0.0189893f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.39
cc_35 VPB A3 0.0343192f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_36 VPB N_A2_M1003_g 0.0381818f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=1.015
cc_37 VPB N_A2_c_100_n 0.0142865f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_38 VPB N_A2_c_105_n 0.0183796f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_39 VPB A2 0.00351152f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.09
cc_40 VPB N_A1_M1000_g 0.0356208f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.39
cc_41 VPB N_A1_c_144_n 0.0122162f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_42 VPB N_A1_c_149_n 0.0165215f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_43 VPB A1 0.00152328f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.09
cc_44 VPB N_B1_c_198_n 0.021217f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.61
cc_45 VPB N_B1_c_199_n 0.0216126f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.315
cc_46 VPB N_B1_c_200_n 0.018841f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_47 VPB N_B1_c_195_n 0.00447422f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_48 VPB N_B1_c_202_n 0.0179202f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_49 VPB B1 0.00587327f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_50 VPB N_VPWR_c_244_n 0.0217005f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.71
cc_51 VPB N_VPWR_c_245_n 0.00527219f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.09
cc_52 VPB N_VPWR_c_246_n 0.0145539f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_53 VPB N_VPWR_c_247_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_54 VPB N_VPWR_c_248_n 0.0158991f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_55 VPB N_VPWR_c_249_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_56 VPB N_VPWR_c_250_n 0.0393882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_243_n 0.0770647f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.665
cc_58 VPB N_A_169_500#_c_277_n 0.0155761f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_59 VPB N_A_169_500#_c_278_n 0.00569047f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_60 VPB N_Y_c_302_n 0.0297138f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.62
cc_61 VPB Y 0.0407623f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_62 N_A3_c_63_n N_A2_M1003_g 0.00199395f $X=0.36 $Y=2.24 $X2=0 $Y2=0
cc_63 N_A3_c_71_n N_A2_M1003_g 0.0215139f $X=0.695 $Y=2.315 $X2=0 $Y2=0
cc_64 N_A3_c_66_n N_A2_M1004_g 0.0489031f $X=0.87 $Y=0.94 $X2=0 $Y2=0
cc_65 N_A3_c_69_n N_A2_M1004_g 0.00164362f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_66 N_A3_c_67_n N_A2_c_100_n 0.00440099f $X=0.27 $Y=1.61 $X2=0 $Y2=0
cc_67 N_A3_c_63_n N_A2_c_105_n 0.00440099f $X=0.36 $Y=2.24 $X2=0 $Y2=0
cc_68 N_A3_c_63_n A2 0.00179918f $X=0.36 $Y=2.24 $X2=0 $Y2=0
cc_69 N_A3_c_66_n A2 0.011193f $X=0.87 $Y=0.94 $X2=0 $Y2=0
cc_70 N_A3_c_69_n A2 0.00558561f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_71 A3 N_A2_c_102_n 0.00342905f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_72 N_A3_c_69_n N_A2_c_102_n 0.00440099f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A3_c_72_n N_VPWR_c_244_n 0.0101374f $X=0.435 $Y=2.315 $X2=0 $Y2=0
cc_74 N_A3_c_73_n N_VPWR_c_244_n 0.0100076f $X=0.77 $Y=2.39 $X2=0 $Y2=0
cc_75 N_A3_c_73_n N_VPWR_c_245_n 7.3042e-19 $X=0.77 $Y=2.39 $X2=0 $Y2=0
cc_76 N_A3_c_73_n N_VPWR_c_248_n 0.00455951f $X=0.77 $Y=2.39 $X2=0 $Y2=0
cc_77 N_A3_c_73_n N_VPWR_c_243_n 0.00447788f $X=0.77 $Y=2.39 $X2=0 $Y2=0
cc_78 A3 N_VPWR_c_243_n 0.00780715f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_79 N_A3_c_71_n N_A_169_500#_c_278_n 0.00257058f $X=0.695 $Y=2.315 $X2=0 $Y2=0
cc_80 A3 N_A_169_500#_c_278_n 0.00545759f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A3_c_64_n N_VGND_c_332_n 0.00986778f $X=0.795 $Y=1.015 $X2=0 $Y2=0
cc_82 N_A3_c_66_n N_VGND_c_332_n 0.00968764f $X=0.87 $Y=0.94 $X2=0 $Y2=0
cc_83 N_A3_c_66_n N_VGND_c_336_n 0.00455951f $X=0.87 $Y=0.94 $X2=0 $Y2=0
cc_84 N_A3_c_66_n N_VGND_c_338_n 0.00447788f $X=0.87 $Y=0.94 $X2=0 $Y2=0
cc_85 A3 N_VGND_c_338_n 0.00780715f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A2_M1004_g N_A1_M1005_g 0.0252403f $X=1.23 $Y=0.62 $X2=0 $Y2=0
cc_87 A2 N_A1_M1005_g 0.00508683f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_88 N_A2_M1003_g N_A1_M1000_g 0.0333954f $X=1.2 $Y=2.71 $X2=0 $Y2=0
cc_89 A2 N_A1_M1000_g 7.29839e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A2_c_100_n N_A1_c_144_n 0.0252403f $X=1.14 $Y=1.835 $X2=0 $Y2=0
cc_91 N_A2_c_105_n N_A1_c_149_n 0.0252403f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_92 N_A2_M1004_g A1 0.00445121f $X=1.23 $Y=0.62 $X2=0 $Y2=0
cc_93 A2 A1 0.0711308f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_94 N_A2_c_102_n N_A1_c_146_n 0.0252403f $X=1.14 $Y=1.495 $X2=0 $Y2=0
cc_95 N_A2_M1003_g N_VPWR_c_244_n 7.36388e-19 $X=1.2 $Y=2.71 $X2=0 $Y2=0
cc_96 N_A2_M1003_g N_VPWR_c_245_n 0.00793595f $X=1.2 $Y=2.71 $X2=0 $Y2=0
cc_97 N_A2_M1003_g N_VPWR_c_248_n 0.00455951f $X=1.2 $Y=2.71 $X2=0 $Y2=0
cc_98 N_A2_M1003_g N_VPWR_c_243_n 0.00447788f $X=1.2 $Y=2.71 $X2=0 $Y2=0
cc_99 N_A2_M1003_g N_A_169_500#_c_277_n 0.0112605f $X=1.2 $Y=2.71 $X2=0 $Y2=0
cc_100 N_A2_c_105_n N_A_169_500#_c_277_n 0.00104857f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_101 A2 N_A_169_500#_c_277_n 0.0137645f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_102 N_A2_c_105_n N_A_169_500#_c_278_n 0.00315551f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_103 A2 N_A_169_500#_c_278_n 0.00106241f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 N_A2_M1004_g N_VGND_c_332_n 0.00112191f $X=1.23 $Y=0.62 $X2=0 $Y2=0
cc_105 A2 N_VGND_c_332_n 0.011188f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_106 N_A2_M1004_g N_VGND_c_336_n 0.00423474f $X=1.23 $Y=0.62 $X2=0 $Y2=0
cc_107 A2 N_VGND_c_336_n 0.00563313f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A2_M1004_g N_VGND_c_338_n 0.00533081f $X=1.23 $Y=0.62 $X2=0 $Y2=0
cc_109 A2 N_VGND_c_338_n 0.007657f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_110 A2 A_189_82# 0.00437911f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_111 N_A1_M1000_g N_B1_c_199_n 0.00817109f $X=1.63 $Y=2.71 $X2=0 $Y2=0
cc_112 N_A1_c_149_n N_B1_c_199_n 0.00633822f $X=1.68 $Y=2 $X2=0 $Y2=0
cc_113 A1 N_B1_c_199_n 5.67385e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_114 N_A1_M1005_g N_B1_M1002_g 0.0127243f $X=1.59 $Y=0.62 $X2=0 $Y2=0
cc_115 A1 N_B1_M1002_g 0.00437276f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_116 N_A1_M1000_g N_B1_c_200_n 0.0222213f $X=1.63 $Y=2.71 $X2=0 $Y2=0
cc_117 N_A1_c_144_n N_B1_c_195_n 0.0113346f $X=1.68 $Y=1.835 $X2=0 $Y2=0
cc_118 N_A1_c_149_n N_B1_c_202_n 0.0113346f $X=1.68 $Y=2 $X2=0 $Y2=0
cc_119 A1 B1 0.0241896f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_120 N_A1_c_146_n B1 0.00155416f $X=1.68 $Y=1.495 $X2=0 $Y2=0
cc_121 N_A1_M1000_g B1 3.91157e-19 $X=1.63 $Y=2.71 $X2=0 $Y2=0
cc_122 N_A1_c_144_n B1 4.10178e-19 $X=1.68 $Y=1.835 $X2=0 $Y2=0
cc_123 N_A1_c_149_n B1 7.76629e-19 $X=1.68 $Y=2 $X2=0 $Y2=0
cc_124 A1 B1 0.0164127f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A1_M1005_g N_B1_c_197_n 0.00331856f $X=1.59 $Y=0.62 $X2=0 $Y2=0
cc_126 A1 N_B1_c_197_n 0.00259466f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_127 N_A1_c_146_n N_B1_c_197_n 0.0113346f $X=1.68 $Y=1.495 $X2=0 $Y2=0
cc_128 N_A1_M1000_g N_VPWR_c_245_n 0.00815163f $X=1.63 $Y=2.71 $X2=0 $Y2=0
cc_129 N_A1_M1000_g N_VPWR_c_250_n 0.00455951f $X=1.63 $Y=2.71 $X2=0 $Y2=0
cc_130 N_A1_M1000_g N_VPWR_c_243_n 0.00447788f $X=1.63 $Y=2.71 $X2=0 $Y2=0
cc_131 N_A1_M1000_g N_A_169_500#_c_277_n 0.012493f $X=1.63 $Y=2.71 $X2=0 $Y2=0
cc_132 N_A1_c_149_n N_A_169_500#_c_277_n 0.00473865f $X=1.68 $Y=2 $X2=0 $Y2=0
cc_133 A1 N_A_169_500#_c_277_n 0.0105919f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_134 A1 N_Y_M1005_d 0.00455774f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_135 N_A1_M1005_g N_Y_c_305_n 0.0010315f $X=1.59 $Y=0.62 $X2=0 $Y2=0
cc_136 A1 N_Y_c_305_n 0.0205537f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_A1_M1005_g N_Y_c_300_n 6.65953e-19 $X=1.59 $Y=0.62 $X2=0 $Y2=0
cc_138 A1 N_Y_c_300_n 0.0125801f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_A1_M1005_g N_VGND_c_334_n 8.61044e-19 $X=1.59 $Y=0.62 $X2=0 $Y2=0
cc_140 A1 N_VGND_c_334_n 0.00137773f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A1_M1005_g N_VGND_c_336_n 0.00481722f $X=1.59 $Y=0.62 $X2=0 $Y2=0
cc_142 A1 N_VGND_c_336_n 0.00398853f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A1_M1005_g N_VGND_c_338_n 0.00533081f $X=1.59 $Y=0.62 $X2=0 $Y2=0
cc_144 A1 N_VGND_c_338_n 0.00566862f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_145 N_B1_c_198_n N_VPWR_c_245_n 0.0011975f $X=2.06 $Y=2.39 $X2=0 $Y2=0
cc_146 N_B1_c_198_n N_VPWR_c_250_n 0.00548708f $X=2.06 $Y=2.39 $X2=0 $Y2=0
cc_147 N_B1_c_198_n N_VPWR_c_243_n 0.00533081f $X=2.06 $Y=2.39 $X2=0 $Y2=0
cc_148 N_B1_c_200_n N_A_169_500#_c_277_n 0.00250539f $X=2.16 $Y=2.315 $X2=0
+ $Y2=0
cc_149 N_B1_M1002_g N_Y_c_305_n 2.41059e-19 $X=2.31 $Y=0.62 $X2=0 $Y2=0
cc_150 N_B1_c_198_n N_Y_c_302_n 4.585e-19 $X=2.06 $Y=2.39 $X2=0 $Y2=0
cc_151 N_B1_c_200_n N_Y_c_302_n 0.0020933f $X=2.16 $Y=2.315 $X2=0 $Y2=0
cc_152 N_B1_c_202_n N_Y_c_302_n 0.00264668f $X=2.22 $Y=1.88 $X2=0 $Y2=0
cc_153 B1 N_Y_c_302_n 0.00555428f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_154 N_B1_M1002_g N_Y_c_299_n 0.0161923f $X=2.31 $Y=0.62 $X2=0 $Y2=0
cc_155 B1 N_Y_c_299_n 0.00845871f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B1_c_197_n N_Y_c_299_n 3.67359e-19 $X=2.22 $Y=1.375 $X2=0 $Y2=0
cc_157 B1 N_Y_c_300_n 0.00799148f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_B1_c_197_n N_Y_c_300_n 0.00170321f $X=2.22 $Y=1.375 $X2=0 $Y2=0
cc_159 N_B1_c_198_n Y 0.00153177f $X=2.06 $Y=2.39 $X2=0 $Y2=0
cc_160 N_B1_c_199_n Y 0.00911377f $X=2.16 $Y=2.24 $X2=0 $Y2=0
cc_161 N_B1_M1002_g Y 0.0224119f $X=2.31 $Y=0.62 $X2=0 $Y2=0
cc_162 B1 Y 0.0303555f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_163 B1 Y 0.0182805f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_164 N_B1_M1002_g N_VGND_c_334_n 0.0102495f $X=2.31 $Y=0.62 $X2=0 $Y2=0
cc_165 N_B1_M1002_g N_VGND_c_336_n 0.00455951f $X=2.31 $Y=0.62 $X2=0 $Y2=0
cc_166 N_B1_M1002_g N_VGND_c_338_n 0.00447788f $X=2.31 $Y=0.62 $X2=0 $Y2=0
cc_167 N_VPWR_c_248_n N_A_169_500#_c_290_n 0.00389976f $X=1.25 $Y=3.33 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_243_n N_A_169_500#_c_290_n 0.00535446f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_169 N_VPWR_M1003_d N_A_169_500#_c_277_n 0.00177921f $X=1.275 $Y=2.5 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_245_n N_A_169_500#_c_277_n 0.0158947f $X=1.415 $Y=2.795 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_243_n N_A_169_500#_c_277_n 0.0128809f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_250_n N_A_169_500#_c_295_n 0.00415318f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_243_n N_A_169_500#_c_295_n 0.00600028f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_250_n N_Y_c_302_n 0.0135693f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_175 N_VPWR_c_243_n N_Y_c_302_n 0.0179049f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_176 N_A_169_500#_c_277_n N_Y_c_302_n 0.00138245f $X=1.76 $Y=2.425 $X2=0 $Y2=0
cc_177 N_A_169_500#_c_277_n Y 0.00480525f $X=1.76 $Y=2.425 $X2=0 $Y2=0
cc_178 N_Y_c_299_n N_VGND_c_334_n 0.0238409f $X=2.555 $Y=0.925 $X2=0 $Y2=0
cc_179 N_Y_c_305_n N_VGND_c_336_n 0.00512596f $X=2.075 $Y=0.685 $X2=0 $Y2=0
cc_180 N_Y_c_305_n N_VGND_c_338_n 0.00676033f $X=2.075 $Y=0.685 $X2=0 $Y2=0
cc_181 N_Y_c_299_n N_VGND_c_338_n 0.0083624f $X=2.555 $Y=0.925 $X2=0 $Y2=0
