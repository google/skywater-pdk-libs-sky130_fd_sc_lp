* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor2_2 A B VGND VNB VPB VPWR Y
X0 Y a_162_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_162_367# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_545_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Y B a_545_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_162_367# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND B a_555_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR A a_545_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_555_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_27_47# B a_162_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_545_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR B a_162_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_162_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR A a_162_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND A a_555_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_555_65# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_555_65# a_162_367# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VPWR a_162_367# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 Y a_162_367# a_555_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
