* File: sky130_fd_sc_lp__fa_lp.pxi.spice
* Created: Fri Aug 28 10:35:07 2020
* 
x_PM_SKY130_FD_SC_LP__FA_LP%A_84_209# N_A_84_209#_M1007_d N_A_84_209#_M1011_d
+ N_A_84_209#_M1014_g N_A_84_209#_M1018_g N_A_84_209#_M1005_g
+ N_A_84_209#_M1010_g N_A_84_209#_c_189_n N_A_84_209#_M1023_g
+ N_A_84_209#_c_190_n N_A_84_209#_c_191_n N_A_84_209#_c_192_n
+ N_A_84_209#_c_208_n N_A_84_209#_c_193_n N_A_84_209#_c_213_p
+ N_A_84_209#_c_291_p N_A_84_209#_c_209_n N_A_84_209#_c_210_n
+ N_A_84_209#_c_221_p N_A_84_209#_c_222_p N_A_84_209#_c_224_p
+ N_A_84_209#_c_194_n N_A_84_209#_c_195_n N_A_84_209#_c_196_n
+ N_A_84_209#_c_197_n N_A_84_209#_c_198_n N_A_84_209#_c_199_n
+ N_A_84_209#_c_200_n N_A_84_209#_c_201_n N_A_84_209#_c_202_n
+ PM_SKY130_FD_SC_LP__FA_LP%A_84_209#
x_PM_SKY130_FD_SC_LP__FA_LP%B N_B_c_382_n N_B_M1007_g N_B_c_383_n N_B_M1011_g
+ N_B_c_384_n N_B_M1015_g N_B_c_385_n N_B_c_401_n N_B_M1016_g N_B_c_402_n
+ N_B_c_386_n N_B_M1024_g N_B_c_403_n N_B_M1000_g N_B_c_387_n N_B_M1012_g
+ N_B_M1025_g N_B_c_405_n N_B_c_388_n N_B_c_389_n N_B_c_390_n N_B_c_391_n
+ N_B_c_436_n N_B_c_438_n N_B_c_392_n N_B_c_393_n N_B_c_394_n N_B_c_440_n
+ N_B_c_441_n B N_B_c_396_n N_B_c_397_n PM_SKY130_FD_SC_LP__FA_LP%B
x_PM_SKY130_FD_SC_LP__FA_LP%CIN N_CIN_c_574_n N_CIN_M1002_g N_CIN_M1027_g
+ N_CIN_M1004_g N_CIN_M1028_g N_CIN_M1022_g N_CIN_M1009_g N_CIN_c_577_n
+ N_CIN_c_578_n N_CIN_c_590_n N_CIN_c_579_n N_CIN_c_592_n N_CIN_c_580_n
+ N_CIN_c_581_n N_CIN_c_582_n CIN N_CIN_c_584_n N_CIN_c_585_n
+ PM_SKY130_FD_SC_LP__FA_LP%CIN
x_PM_SKY130_FD_SC_LP__FA_LP%A N_A_c_727_n N_A_M1029_g N_A_c_729_n N_A_c_730_n
+ N_A_c_731_n N_A_M1021_g N_A_M1019_g N_A_M1020_g N_A_M1008_g N_A_c_752_n
+ N_A_M1003_g N_A_c_736_n N_A_M1013_g N_A_M1017_g N_A_c_739_n N_A_c_740_n
+ N_A_c_741_n N_A_c_742_n N_A_c_743_n N_A_c_744_n A A N_A_c_745_n N_A_c_746_n
+ N_A_c_747_n N_A_c_748_n PM_SKY130_FD_SC_LP__FA_LP%A
x_PM_SKY130_FD_SC_LP__FA_LP%A_1574_141# N_A_1574_141#_M1010_d
+ N_A_1574_141#_M1023_d N_A_1574_141#_c_894_n N_A_1574_141#_M1006_g
+ N_A_1574_141#_c_895_n N_A_1574_141#_c_896_n N_A_1574_141#_M1001_g
+ N_A_1574_141#_c_897_n N_A_1574_141#_M1026_g N_A_1574_141#_c_898_n
+ N_A_1574_141#_c_899_n N_A_1574_141#_c_909_n N_A_1574_141#_c_900_n
+ N_A_1574_141#_c_912_n N_A_1574_141#_c_901_n N_A_1574_141#_c_923_n
+ N_A_1574_141#_c_913_n N_A_1574_141#_c_902_n N_A_1574_141#_c_903_n
+ N_A_1574_141#_c_904_n N_A_1574_141#_c_953_n N_A_1574_141#_c_905_n
+ N_A_1574_141#_c_906_n PM_SKY130_FD_SC_LP__FA_LP%A_1574_141#
x_PM_SKY130_FD_SC_LP__FA_LP%COUT N_COUT_M1018_s N_COUT_M1014_s COUT COUT COUT
+ COUT COUT COUT COUT COUT PM_SKY130_FD_SC_LP__FA_LP%COUT
x_PM_SKY130_FD_SC_LP__FA_LP%VPWR N_VPWR_M1014_d N_VPWR_M1029_d N_VPWR_M1016_d
+ N_VPWR_M1028_d N_VPWR_M1017_d N_VPWR_c_1014_n N_VPWR_c_1015_n N_VPWR_c_1016_n
+ N_VPWR_c_1017_n N_VPWR_c_1018_n N_VPWR_c_1019_n N_VPWR_c_1020_n
+ N_VPWR_c_1021_n N_VPWR_c_1022_n N_VPWR_c_1023_n N_VPWR_c_1024_n VPWR
+ N_VPWR_c_1025_n N_VPWR_c_1026_n N_VPWR_c_1013_n N_VPWR_c_1028_n
+ N_VPWR_c_1029_n PM_SKY130_FD_SC_LP__FA_LP%VPWR
x_PM_SKY130_FD_SC_LP__FA_LP%A_245_409# N_A_245_409#_M1029_s N_A_245_409#_M1011_s
+ N_A_245_409#_c_1125_n N_A_245_409#_c_1126_n N_A_245_409#_c_1127_n
+ N_A_245_409#_c_1128_n N_A_245_409#_c_1129_n N_A_245_409#_c_1130_n
+ PM_SKY130_FD_SC_LP__FA_LP%A_245_409#
x_PM_SKY130_FD_SC_LP__FA_LP%A_458_409# N_A_458_409#_M1021_d N_A_458_409#_M1027_d
+ N_A_458_409#_c_1168_n N_A_458_409#_c_1169_n N_A_458_409#_c_1170_n
+ N_A_458_409#_c_1174_n PM_SKY130_FD_SC_LP__FA_LP%A_458_409#
x_PM_SKY130_FD_SC_LP__FA_LP%A_1049_419# N_A_1049_419#_M1000_d
+ N_A_1049_419#_M1003_d N_A_1049_419#_c_1209_n N_A_1049_419#_c_1205_n
+ N_A_1049_419#_c_1211_n N_A_1049_419#_c_1206_n
+ PM_SKY130_FD_SC_LP__FA_LP%A_1049_419#
x_PM_SKY130_FD_SC_LP__FA_LP%SUM N_SUM_M1026_d N_SUM_M1001_d N_SUM_c_1242_n
+ N_SUM_c_1239_n SUM SUM SUM PM_SKY130_FD_SC_LP__FA_LP%SUM
x_PM_SKY130_FD_SC_LP__FA_LP%VGND N_VGND_M1005_d N_VGND_M1019_d N_VGND_M1015_d
+ N_VGND_M1004_d N_VGND_M1013_d N_VGND_c_1263_n N_VGND_c_1264_n N_VGND_c_1265_n
+ N_VGND_c_1266_n N_VGND_c_1267_n N_VGND_c_1268_n N_VGND_c_1269_n
+ N_VGND_c_1270_n N_VGND_c_1271_n N_VGND_c_1272_n N_VGND_c_1273_n VGND
+ N_VGND_c_1274_n N_VGND_c_1275_n N_VGND_c_1276_n N_VGND_c_1277_n
+ N_VGND_c_1278_n N_VGND_c_1279_n N_VGND_c_1280_n N_VGND_c_1281_n
+ PM_SKY130_FD_SC_LP__FA_LP%VGND
x_PM_SKY130_FD_SC_LP__FA_LP%A_355_141# N_A_355_141#_M1019_s N_A_355_141#_M1002_d
+ N_A_355_141#_c_1391_n N_A_355_141#_c_1392_n N_A_355_141#_c_1393_n
+ N_A_355_141#_c_1394_n PM_SKY130_FD_SC_LP__FA_LP%A_355_141#
x_PM_SKY130_FD_SC_LP__FA_LP%A_1005_141# N_A_1005_141#_M1024_d
+ N_A_1005_141#_M1008_d N_A_1005_141#_c_1430_n N_A_1005_141#_c_1431_n
+ N_A_1005_141#_c_1432_n N_A_1005_141#_c_1439_n N_A_1005_141#_c_1433_n
+ N_A_1005_141#_c_1434_n N_A_1005_141#_c_1435_n
+ PM_SKY130_FD_SC_LP__FA_LP%A_1005_141#
cc_1 VNB N_A_84_209#_M1018_g 0.0240902f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.635
cc_2 VNB N_A_84_209#_M1005_g 0.021505f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.635
cc_3 VNB N_A_84_209#_M1010_g 0.0211871f $X=-0.19 $Y=-0.245 $X2=7.795 $Y2=0.915
cc_4 VNB N_A_84_209#_c_189_n 0.0342932f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=1.76
cc_5 VNB N_A_84_209#_c_190_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.21
cc_6 VNB N_A_84_209#_c_191_n 0.0759782f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.21
cc_7 VNB N_A_84_209#_c_192_n 0.0261627f $X=-0.19 $Y=-0.245 $X2=2.775 $Y2=1.63
cc_8 VNB N_A_84_209#_c_193_n 0.00669818f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=1.545
cc_9 VNB N_A_84_209#_c_194_n 0.00227164f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=0.915
cc_10 VNB N_A_84_209#_c_195_n 0.00319857f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=1.465
cc_11 VNB N_A_84_209#_c_196_n 0.021465f $X=-0.19 $Y=-0.245 $X2=6.45 $Y2=1.55
cc_12 VNB N_A_84_209#_c_197_n 0.00272316f $X=-0.19 $Y=-0.245 $X2=5.06 $Y2=1.55
cc_13 VNB N_A_84_209#_c_198_n 0.00809192f $X=-0.19 $Y=-0.245 $X2=7.845 $Y2=1.47
cc_14 VNB N_A_84_209#_c_199_n 0.00204046f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=1.63
cc_15 VNB N_A_84_209#_c_200_n 0.0130769f $X=-0.19 $Y=-0.245 $X2=6.535 $Y2=1.285
cc_16 VNB N_A_84_209#_c_201_n 0.0146399f $X=-0.19 $Y=-0.245 $X2=7.26 $Y2=1.417
cc_17 VNB N_A_84_209#_c_202_n 0.00383335f $X=-0.19 $Y=-0.245 $X2=7.43 $Y2=1.417
cc_18 VNB N_B_c_382_n 0.0167737f $X=-0.19 $Y=-0.245 $X2=3.275 $Y2=0.705
cc_19 VNB N_B_c_383_n 0.0436974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_c_384_n 0.0161477f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.415
cc_21 VNB N_B_c_385_n 0.00325329f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.635
cc_22 VNB N_B_c_386_n 0.0156539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_387_n 0.015402f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=2.595
cc_24 VNB N_B_c_388_n 0.0230978f $X=-0.19 $Y=-0.245 $X2=3.25 $Y2=0.942
cc_25 VNB N_B_c_389_n 0.00729538f $X=-0.19 $Y=-0.245 $X2=3.255 $Y2=1.83
cc_26 VNB N_B_c_390_n 0.00182671f $X=-0.19 $Y=-0.245 $X2=3.695 $Y2=2.54
cc_27 VNB N_B_c_391_n 0.00915997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_392_n 0.00156735f $X=-0.19 $Y=-0.245 $X2=6.62 $Y2=1.285
cc_29 VNB N_B_c_393_n 0.00799019f $X=-0.19 $Y=-0.245 $X2=7.43 $Y2=1.47
cc_30 VNB N_B_c_394_n 0.00233498f $X=-0.19 $Y=-0.245 $X2=7.845 $Y2=1.47
cc_31 VNB B 0.00387651f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=1.63
cc_32 VNB N_B_c_396_n 0.0584113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_c_397_n 0.014428f $X=-0.19 $Y=-0.245 $X2=7.43 $Y2=1.417
cc_34 VNB N_CIN_c_574_n 0.0162902f $X=-0.19 $Y=-0.245 $X2=3.275 $Y2=0.705
cc_35 VNB N_CIN_M1004_g 0.0386246f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.635
cc_36 VNB N_CIN_M1022_g 0.0353977f $X=-0.19 $Y=-0.245 $X2=7.795 $Y2=0.915
cc_37 VNB N_CIN_c_577_n 0.0168476f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.21
cc_38 VNB N_CIN_c_578_n 0.0184657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_CIN_c_579_n 0.00297178f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.63
cc_40 VNB N_CIN_c_580_n 0.0115579f $X=-0.19 $Y=-0.245 $X2=3.255 $Y2=1.83
cc_41 VNB N_CIN_c_581_n 0.00180961f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=1.915
cc_42 VNB N_CIN_c_582_n 0.00857711f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=2.45
cc_43 VNB CIN 0.00327042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_CIN_c_584_n 0.0465576f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=1
cc_45 VNB N_CIN_c_585_n 0.0143797f $X=-0.19 $Y=-0.245 $X2=7.26 $Y2=1.285
cc_46 VNB N_A_c_727_n 0.054994f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=2.095
cc_47 VNB N_A_M1029_g 0.016278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_c_729_n 0.072192f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.715
cc_49 VNB N_A_c_730_n 0.0113868f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.415
cc_50 VNB N_A_c_731_n 0.0145636f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.415
cc_51 VNB N_A_M1021_g 0.0177393f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.635
cc_52 VNB N_A_M1019_g 0.0188895f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.635
cc_53 VNB N_A_M1020_g 0.0456974f $X=-0.19 $Y=-0.245 $X2=7.795 $Y2=0.915
cc_54 VNB N_A_M1008_g 0.0385295f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.21
cc_55 VNB N_A_c_736_n 0.145451f $X=-0.19 $Y=-0.245 $X2=2.775 $Y2=1.63
cc_56 VNB N_A_M1013_g 0.00994473f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=0.942
cc_57 VNB N_A_M1017_g 0.0166566f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=2.582
cc_58 VNB N_A_c_739_n 0.00739381f $X=-0.19 $Y=-0.245 $X2=3.695 $Y2=2.54
cc_59 VNB N_A_c_740_n 0.00871625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_c_741_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=4.89 $Y2=0.915
cc_61 VNB N_A_c_742_n 0.0146952f $X=-0.19 $Y=-0.245 $X2=6.45 $Y2=1.55
cc_62 VNB N_A_c_743_n 0.0164602f $X=-0.19 $Y=-0.245 $X2=7.26 $Y2=1.285
cc_63 VNB N_A_c_744_n 0.0199084f $X=-0.19 $Y=-0.245 $X2=6.62 $Y2=1.285
cc_64 VNB N_A_c_745_n 0.00406307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_c_746_n 0.293138f $X=-0.19 $Y=-0.245 $X2=3.415 $Y2=0.87
cc_66 VNB N_A_c_747_n 0.0887847f $X=-0.19 $Y=-0.245 $X2=6.535 $Y2=1.285
cc_67 VNB N_A_c_748_n 0.0151373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1574_141#_c_894_n 0.0151368f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.715
cc_69 VNB N_A_1574_141#_c_895_n 0.00814236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1574_141#_c_896_n 0.00923997f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=1.045
cc_71 VNB N_A_1574_141#_c_897_n 0.0183145f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=0.635
cc_72 VNB N_A_1574_141#_c_898_n 0.017889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1574_141#_c_899_n 0.0202677f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=1.76
cc_74 VNB N_A_1574_141#_c_900_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=7.945
+ $Y2=2.595
cc_75 VNB N_A_1574_141#_c_901_n 0.0295239f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.21
cc_76 VNB N_A_1574_141#_c_902_n 0.0026182f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=1.545
cc_77 VNB N_A_1574_141#_c_903_n 0.00978788f $X=-0.19 $Y=-0.245 $X2=3.25
+ $Y2=0.942
cc_78 VNB N_A_1574_141#_c_904_n 0.0128158f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=2.45
cc_79 VNB N_A_1574_141#_c_905_n 0.00203096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1574_141#_c_906_n 0.01366f $X=-0.19 $Y=-0.245 $X2=4.89 $Y2=0.915
cc_81 VNB COUT 0.0245031f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.715
cc_82 VNB COUT 0.0347976f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=2.595
cc_83 VNB N_VPWR_c_1013_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_SUM_c_1239_n 0.0289562f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.635
cc_85 VNB SUM 0.0248036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB SUM 0.0138548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1263_n 0.00610239f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.635
cc_88 VNB N_VGND_c_1264_n 0.00336798f $X=-0.19 $Y=-0.245 $X2=7.795 $Y2=1.305
cc_89 VNB N_VGND_c_1265_n 0.0131868f $X=-0.19 $Y=-0.245 $X2=7.795 $Y2=0.915
cc_90 VNB N_VGND_c_1266_n 0.00255393f $X=-0.19 $Y=-0.245 $X2=7.795 $Y2=0.915
cc_91 VNB N_VGND_c_1267_n 0.00306649f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=2.595
cc_92 VNB N_VGND_c_1268_n 0.0125496f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.21
cc_93 VNB N_VGND_c_1269_n 0.0180008f $X=-0.19 $Y=-0.245 $X2=2.775 $Y2=1.63
cc_94 VNB N_VGND_c_1270_n 0.00740028f $X=-0.19 $Y=-0.245 $X2=3.25 $Y2=0.942
cc_95 VNB N_VGND_c_1271_n 0.0155086f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=1.83
cc_96 VNB N_VGND_c_1272_n 0.0196283f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=2.582
cc_97 VNB N_VGND_c_1273_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.695 $Y2=2.582
cc_98 VNB N_VGND_c_1274_n 0.031123f $X=-0.19 $Y=-0.245 $X2=4.89 $Y2=0.915
cc_99 VNB N_VGND_c_1275_n 0.0701323f $X=-0.19 $Y=-0.245 $X2=5.06 $Y2=1.55
cc_100 VNB N_VGND_c_1276_n 0.0950063f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=1.83
cc_101 VNB N_VGND_c_1277_n 0.0297101f $X=-0.19 $Y=-0.245 $X2=7.43 $Y2=1.417
cc_102 VNB N_VGND_c_1278_n 0.516205f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.21
cc_103 VNB N_VGND_c_1279_n 0.00951394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1280_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1281_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_355_141#_c_1391_n 0.00861273f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=2.415
cc_107 VNB N_A_355_141#_c_1392_n 0.0383468f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=1.045
cc_108 VNB N_A_355_141#_c_1393_n 0.00485915f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=0.635
cc_109 VNB N_A_355_141#_c_1394_n 0.0103469f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=0.635
cc_110 VNB N_A_1005_141#_c_1430_n 3.49958e-19 $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=2.415
cc_111 VNB N_A_1005_141#_c_1431_n 0.00590991f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=2.415
cc_112 VNB N_A_1005_141#_c_1432_n 0.00290651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1005_141#_c_1433_n 0.00918254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1005_141#_c_1434_n 0.00583699f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=0.635
cc_115 VNB N_A_1005_141#_c_1435_n 0.0030827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VPB N_A_84_209#_M1014_g 0.0401774f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.415
cc_117 VPB N_A_84_209#_c_189_n 0.006941f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=1.76
cc_118 VPB N_A_84_209#_M1023_g 0.0352236f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=2.595
cc_119 VPB N_A_84_209#_c_191_n 0.0169859f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.21
cc_120 VPB N_A_84_209#_c_192_n 0.0182462f $X=-0.19 $Y=1.655 $X2=2.775 $Y2=1.63
cc_121 VPB N_A_84_209#_c_208_n 0.0048444f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.63
cc_122 VPB N_A_84_209#_c_209_n 0.016182f $X=-0.19 $Y=1.655 $X2=3.255 $Y2=1.83
cc_123 VPB N_A_84_209#_c_210_n 0.00611493f $X=-0.19 $Y=1.655 $X2=3.34 $Y2=2.45
cc_124 VPB N_A_84_209#_c_199_n 0.00717489f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=1.63
cc_125 VPB N_B_c_383_n 0.00432091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_B_M1011_g 0.0461098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_B_c_385_n 0.0123292f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.635
cc_128 VPB N_B_c_401_n 0.0207312f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.635
cc_129 VPB N_B_c_402_n 0.0235267f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=0.635
cc_130 VPB N_B_c_403_n 0.0199918f $X=-0.19 $Y=1.655 $X2=7.795 $Y2=0.915
cc_131 VPB N_B_M1025_g 0.0233355f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.21
cc_132 VPB N_B_c_405_n 0.00792076f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.63
cc_133 VPB N_B_c_390_n 0.00793135f $X=-0.19 $Y=1.655 $X2=3.695 $Y2=2.54
cc_134 VPB N_B_c_392_n 0.00250562f $X=-0.19 $Y=1.655 $X2=6.62 $Y2=1.285
cc_135 VPB N_B_c_393_n 0.0214132f $X=-0.19 $Y=1.655 $X2=7.43 $Y2=1.47
cc_136 VPB N_CIN_M1027_g 0.0279596f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.415
cc_137 VPB N_CIN_M1028_g 0.0321975f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=0.635
cc_138 VPB N_CIN_M1009_g 0.024845f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=2.595
cc_139 VPB N_CIN_c_578_n 0.018136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_CIN_c_590_n 0.0202274f $X=-0.19 $Y=1.655 $X2=2.775 $Y2=1.63
cc_141 VPB N_CIN_c_579_n 0.0076944f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.63
cc_142 VPB N_CIN_c_592_n 0.0180089f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=1.055
cc_143 VPB N_CIN_c_580_n 0.0231702f $X=-0.19 $Y=1.655 $X2=3.255 $Y2=1.83
cc_144 VPB N_CIN_c_581_n 0.00117056f $X=-0.19 $Y=1.655 $X2=3.34 $Y2=1.915
cc_145 VPB N_CIN_c_582_n 0.0205858f $X=-0.19 $Y=1.655 $X2=3.34 $Y2=2.45
cc_146 VPB CIN 0.00295066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_CIN_c_584_n 0.0777061f $X=-0.19 $Y=1.655 $X2=4.975 $Y2=1
cc_148 VPB N_A_M1029_g 0.0483045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_M1021_g 0.0455802f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.635
cc_150 VPB N_A_M1008_g 0.0113401f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.21
cc_151 VPB N_A_c_752_n 0.0381571f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.21
cc_152 VPB N_A_M1017_g 0.0399118f $X=-0.19 $Y=1.655 $X2=3.425 $Y2=2.582
cc_153 VPB N_A_1574_141#_M1001_g 0.0332877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_1574_141#_c_899_n 0.00521587f $X=-0.19 $Y=1.655 $X2=7.945
+ $Y2=1.76
cc_155 VPB N_A_1574_141#_c_909_n 0.0147042f $X=-0.19 $Y=1.655 $X2=7.945
+ $Y2=2.595
cc_156 VPB N_A_1574_141#_c_902_n 0.00270571f $X=-0.19 $Y=1.655 $X2=2.86
+ $Y2=1.545
cc_157 VPB N_A_1574_141#_c_905_n 6.65629e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB COUT 0.0525041f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=2.595
cc_159 VPB N_VPWR_c_1014_n 0.019905f $X=-0.19 $Y=1.655 $X2=7.795 $Y2=0.915
cc_160 VPB N_VPWR_c_1015_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1016_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.21
cc_162 VPB N_VPWR_c_1017_n 0.00284591f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=1.055
cc_163 VPB N_VPWR_c_1018_n 0.00928226f $X=-0.19 $Y=1.655 $X2=3.255 $Y2=1.83
cc_164 VPB N_VPWR_c_1019_n 0.0203774f $X=-0.19 $Y=1.655 $X2=3.695 $Y2=2.582
cc_165 VPB N_VPWR_c_1020_n 0.00497896f $X=-0.19 $Y=1.655 $X2=3.695 $Y2=2.54
cc_166 VPB N_VPWR_c_1021_n 0.0621101f $X=-0.19 $Y=1.655 $X2=4.89 $Y2=0.915
cc_167 VPB N_VPWR_c_1022_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.605 $Y2=0.915
cc_168 VPB N_VPWR_c_1023_n 0.0968504f $X=-0.19 $Y=1.655 $X2=4.975 $Y2=1.465
cc_169 VPB N_VPWR_c_1024_n 0.00356964f $X=-0.19 $Y=1.655 $X2=6.45 $Y2=1.55
cc_170 VPB N_VPWR_c_1025_n 0.0171673f $X=-0.19 $Y=1.655 $X2=3.415 $Y2=0.87
cc_171 VPB N_VPWR_c_1026_n 0.018365f $X=-0.19 $Y=1.655 $X2=7.875 $Y2=1.47
cc_172 VPB N_VPWR_c_1013_n 0.0702151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1028_n 0.0266443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1029_n 0.00510127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_245_409#_c_1125_n 0.0112128f $X=-0.19 $Y=1.655 $X2=0.545
+ $Y2=2.415
cc_176 VPB N_A_245_409#_c_1126_n 0.00241151f $X=-0.19 $Y=1.655 $X2=0.595
+ $Y2=0.635
cc_177 VPB N_A_245_409#_c_1127_n 0.00502875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_245_409#_c_1128_n 0.0109099f $X=-0.19 $Y=1.655 $X2=0.955
+ $Y2=1.045
cc_179 VPB N_A_245_409#_c_1129_n 0.00514915f $X=-0.19 $Y=1.655 $X2=7.795
+ $Y2=1.305
cc_180 VPB N_A_245_409#_c_1130_n 0.00587628f $X=-0.19 $Y=1.655 $X2=7.795
+ $Y2=0.915
cc_181 VPB N_A_458_409#_c_1168_n 0.00996687f $X=-0.19 $Y=1.655 $X2=0.545
+ $Y2=2.415
cc_182 VPB N_A_458_409#_c_1169_n 0.00723305f $X=-0.19 $Y=1.655 $X2=0.595
+ $Y2=1.045
cc_183 VPB N_A_458_409#_c_1170_n 0.00245219f $X=-0.19 $Y=1.655 $X2=0.595
+ $Y2=0.635
cc_184 VPB N_SUM_c_1242_n 0.0454269f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.635
cc_185 VPB N_SUM_c_1239_n 0.0198953f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.635
cc_186 N_A_84_209#_c_193_n N_B_c_382_n 0.00360117f $X=2.86 $Y=1.545 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_84_209#_c_213_p N_B_c_382_n 0.00847215f $X=3.25 $Y=0.942 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_84_209#_c_194_n N_B_c_382_n 0.00408938f $X=3.605 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A_84_209#_c_193_n N_B_c_383_n 0.00220719f $X=2.86 $Y=1.545 $X2=0 $Y2=0
cc_190 N_A_84_209#_c_209_n N_B_c_383_n 0.00463745f $X=3.255 $Y=1.83 $X2=0 $Y2=0
cc_191 N_A_84_209#_c_194_n N_B_c_383_n 0.0045237f $X=3.605 $Y=0.915 $X2=0 $Y2=0
cc_192 N_A_84_209#_c_199_n N_B_c_383_n 0.00364086f $X=2.86 $Y=1.63 $X2=0 $Y2=0
cc_193 N_A_84_209#_c_209_n N_B_M1011_g 0.00862459f $X=3.255 $Y=1.83 $X2=0 $Y2=0
cc_194 N_A_84_209#_c_210_n N_B_M1011_g 0.0196314f $X=3.34 $Y=2.45 $X2=0 $Y2=0
cc_195 N_A_84_209#_c_221_p N_B_M1011_g 0.00874322f $X=3.425 $Y=2.582 $X2=0 $Y2=0
cc_196 N_A_84_209#_c_222_p N_B_M1011_g 0.0109435f $X=3.695 $Y=2.54 $X2=0 $Y2=0
cc_197 N_A_84_209#_c_199_n N_B_M1011_g 5.20642e-19 $X=2.86 $Y=1.63 $X2=0 $Y2=0
cc_198 N_A_84_209#_c_224_p N_B_c_384_n 0.0117318f $X=4.89 $Y=0.915 $X2=0 $Y2=0
cc_199 N_A_84_209#_c_195_n N_B_c_384_n 9.88971e-19 $X=4.975 $Y=1.465 $X2=0 $Y2=0
cc_200 N_A_84_209#_c_222_p N_B_c_401_n 3.06813e-19 $X=3.695 $Y=2.54 $X2=0 $Y2=0
cc_201 N_A_84_209#_c_196_n N_B_c_402_n 0.00109936f $X=6.45 $Y=1.55 $X2=0 $Y2=0
cc_202 N_A_84_209#_c_197_n N_B_c_402_n 7.25218e-19 $X=5.06 $Y=1.55 $X2=0 $Y2=0
cc_203 N_A_84_209#_c_224_p N_B_c_386_n 0.00868286f $X=4.89 $Y=0.915 $X2=0 $Y2=0
cc_204 N_A_84_209#_c_195_n N_B_c_386_n 0.0067129f $X=4.975 $Y=1.465 $X2=0 $Y2=0
cc_205 N_A_84_209#_c_193_n N_B_c_389_n 0.0250169f $X=2.86 $Y=1.545 $X2=0 $Y2=0
cc_206 N_A_84_209#_c_213_p N_B_c_389_n 0.00867105f $X=3.25 $Y=0.942 $X2=0 $Y2=0
cc_207 N_A_84_209#_c_209_n N_B_c_389_n 0.0225087f $X=3.255 $Y=1.83 $X2=0 $Y2=0
cc_208 N_A_84_209#_c_194_n N_B_c_389_n 0.024899f $X=3.605 $Y=0.915 $X2=0 $Y2=0
cc_209 N_A_84_209#_c_209_n N_B_c_390_n 0.0126566f $X=3.255 $Y=1.83 $X2=0 $Y2=0
cc_210 N_A_84_209#_c_210_n N_B_c_390_n 0.0124245f $X=3.34 $Y=2.45 $X2=0 $Y2=0
cc_211 N_A_84_209#_c_199_n N_B_c_390_n 0.00520243f $X=2.86 $Y=1.63 $X2=0 $Y2=0
cc_212 N_A_84_209#_c_224_p N_B_c_391_n 0.033482f $X=4.89 $Y=0.915 $X2=0 $Y2=0
cc_213 N_A_84_209#_M1011_d N_B_c_436_n 0.00224566f $X=3.555 $Y=2.095 $X2=0 $Y2=0
cc_214 N_A_84_209#_c_222_p N_B_c_436_n 0.013055f $X=3.695 $Y=2.54 $X2=0 $Y2=0
cc_215 N_A_84_209#_M1023_g N_B_c_438_n 0.0209795f $X=7.945 $Y=2.595 $X2=0 $Y2=0
cc_216 N_A_84_209#_c_224_p N_B_c_394_n 0.00896178f $X=4.89 $Y=0.915 $X2=0 $Y2=0
cc_217 N_A_84_209#_c_222_p N_B_c_440_n 0.00175265f $X=3.695 $Y=2.54 $X2=0 $Y2=0
cc_218 N_A_84_209#_c_210_n N_B_c_441_n 0.0016727f $X=3.34 $Y=2.45 $X2=0 $Y2=0
cc_219 N_A_84_209#_c_224_p B 0.0188116f $X=4.89 $Y=0.915 $X2=0 $Y2=0
cc_220 N_A_84_209#_c_195_n B 0.0191752f $X=4.975 $Y=1.465 $X2=0 $Y2=0
cc_221 N_A_84_209#_c_197_n B 0.00752359f $X=5.06 $Y=1.55 $X2=0 $Y2=0
cc_222 N_A_84_209#_c_224_p N_B_c_396_n 0.00400199f $X=4.89 $Y=0.915 $X2=0 $Y2=0
cc_223 N_A_84_209#_c_195_n N_B_c_396_n 0.00896345f $X=4.975 $Y=1.465 $X2=0 $Y2=0
cc_224 N_A_84_209#_c_197_n N_B_c_396_n 0.00520891f $X=5.06 $Y=1.55 $X2=0 $Y2=0
cc_225 N_A_84_209#_c_224_p N_CIN_c_574_n 0.0124103f $X=4.89 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_84_209#_c_194_n N_CIN_c_574_n 0.00564206f $X=3.605 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_84_209#_c_210_n N_CIN_M1027_g 7.36645e-19 $X=3.34 $Y=2.45 $X2=0 $Y2=0
cc_228 N_A_84_209#_c_222_p N_CIN_M1027_g 0.00564645f $X=3.695 $Y=2.54 $X2=0
+ $Y2=0
cc_229 N_A_84_209#_c_195_n N_CIN_M1004_g 0.00335462f $X=4.975 $Y=1.465 $X2=0
+ $Y2=0
cc_230 N_A_84_209#_c_196_n N_CIN_M1004_g 0.00282299f $X=6.45 $Y=1.55 $X2=0 $Y2=0
cc_231 N_A_84_209#_M1010_g N_CIN_M1022_g 0.0134329f $X=7.795 $Y=0.915 $X2=0
+ $Y2=0
cc_232 N_A_84_209#_c_189_n N_CIN_M1022_g 0.0147851f $X=7.945 $Y=1.76 $X2=0 $Y2=0
cc_233 N_A_84_209#_c_198_n N_CIN_M1022_g 0.0015461f $X=7.845 $Y=1.47 $X2=0 $Y2=0
cc_234 N_A_84_209#_M1023_g N_CIN_M1009_g 0.0452099f $X=7.945 $Y=2.595 $X2=0
+ $Y2=0
cc_235 N_A_84_209#_c_224_p N_CIN_c_577_n 0.00350648f $X=4.89 $Y=0.915 $X2=0
+ $Y2=0
cc_236 N_A_84_209#_c_196_n N_CIN_c_578_n 0.0158834f $X=6.45 $Y=1.55 $X2=0 $Y2=0
cc_237 N_A_84_209#_c_196_n N_CIN_c_590_n 0.0934164f $X=6.45 $Y=1.55 $X2=0 $Y2=0
cc_238 N_A_84_209#_c_197_n N_CIN_c_590_n 0.0137842f $X=5.06 $Y=1.55 $X2=0 $Y2=0
cc_239 N_A_84_209#_c_200_n N_CIN_c_590_n 0.0117766f $X=6.535 $Y=1.285 $X2=0
+ $Y2=0
cc_240 N_A_84_209#_c_201_n N_CIN_c_590_n 0.00626929f $X=7.26 $Y=1.417 $X2=0
+ $Y2=0
cc_241 N_A_84_209#_c_197_n N_CIN_c_579_n 0.00133162f $X=5.06 $Y=1.55 $X2=0 $Y2=0
cc_242 N_A_84_209#_c_189_n N_CIN_c_592_n 0.00350848f $X=7.945 $Y=1.76 $X2=0
+ $Y2=0
cc_243 N_A_84_209#_M1023_g N_CIN_c_592_n 0.0161481f $X=7.945 $Y=2.595 $X2=0
+ $Y2=0
cc_244 N_A_84_209#_c_201_n N_CIN_c_592_n 0.00695228f $X=7.26 $Y=1.417 $X2=0
+ $Y2=0
cc_245 N_A_84_209#_c_202_n N_CIN_c_592_n 0.0540634f $X=7.43 $Y=1.417 $X2=0 $Y2=0
cc_246 N_A_84_209#_c_197_n N_CIN_c_580_n 2.03566e-19 $X=5.06 $Y=1.55 $X2=0 $Y2=0
cc_247 N_A_84_209#_c_189_n N_CIN_c_581_n 0.0012945f $X=7.945 $Y=1.76 $X2=0 $Y2=0
cc_248 N_A_84_209#_c_198_n N_CIN_c_581_n 0.00159672f $X=7.845 $Y=1.47 $X2=0
+ $Y2=0
cc_249 N_A_84_209#_c_189_n N_CIN_c_582_n 0.0196943f $X=7.945 $Y=1.76 $X2=0 $Y2=0
cc_250 N_A_84_209#_c_200_n CIN 0.00603641f $X=6.535 $Y=1.285 $X2=0 $Y2=0
cc_251 N_A_84_209#_c_201_n CIN 0.0217347f $X=7.26 $Y=1.417 $X2=0 $Y2=0
cc_252 N_A_84_209#_c_202_n CIN 0.00687283f $X=7.43 $Y=1.417 $X2=0 $Y2=0
cc_253 N_A_84_209#_c_196_n N_CIN_c_584_n 0.0238504f $X=6.45 $Y=1.55 $X2=0 $Y2=0
cc_254 N_A_84_209#_c_200_n N_CIN_c_584_n 0.00750594f $X=6.535 $Y=1.285 $X2=0
+ $Y2=0
cc_255 N_A_84_209#_c_201_n N_CIN_c_584_n 0.00606568f $X=7.26 $Y=1.417 $X2=0
+ $Y2=0
cc_256 N_A_84_209#_c_202_n N_CIN_c_584_n 2.97621e-19 $X=7.43 $Y=1.417 $X2=0
+ $Y2=0
cc_257 N_A_84_209#_M1005_g N_A_c_727_n 0.0136159f $X=0.955 $Y=0.635 $X2=0 $Y2=0
cc_258 N_A_84_209#_c_190_n N_A_c_727_n 3.45975e-19 $X=0.865 $Y=1.21 $X2=0 $Y2=0
cc_259 N_A_84_209#_c_192_n N_A_M1029_g 0.0158571f $X=2.775 $Y=1.63 $X2=0 $Y2=0
cc_260 N_A_84_209#_c_192_n N_A_c_731_n 0.00199111f $X=2.775 $Y=1.63 $X2=0 $Y2=0
cc_261 N_A_84_209#_c_192_n N_A_M1021_g 0.016754f $X=2.775 $Y=1.63 $X2=0 $Y2=0
cc_262 N_A_84_209#_c_199_n N_A_M1021_g 0.00763904f $X=2.86 $Y=1.63 $X2=0 $Y2=0
cc_263 N_A_84_209#_c_192_n N_A_M1020_g 0.0014603f $X=2.775 $Y=1.63 $X2=0 $Y2=0
cc_264 N_A_84_209#_c_193_n N_A_M1020_g 0.0065806f $X=2.86 $Y=1.545 $X2=0 $Y2=0
cc_265 N_A_84_209#_c_291_p N_A_M1020_g 0.00827832f $X=2.945 $Y=0.942 $X2=0 $Y2=0
cc_266 N_A_84_209#_c_194_n N_A_M1020_g 4.42998e-19 $X=3.605 $Y=0.915 $X2=0 $Y2=0
cc_267 N_A_84_209#_c_189_n N_A_M1008_g 0.0270775f $X=7.945 $Y=1.76 $X2=0 $Y2=0
cc_268 N_A_84_209#_c_198_n N_A_M1008_g 0.00391475f $X=7.845 $Y=1.47 $X2=0 $Y2=0
cc_269 N_A_84_209#_c_200_n N_A_M1008_g 0.0011999f $X=6.535 $Y=1.285 $X2=0 $Y2=0
cc_270 N_A_84_209#_c_202_n N_A_M1008_g 0.0186487f $X=7.43 $Y=1.417 $X2=0 $Y2=0
cc_271 N_A_84_209#_M1023_g N_A_c_752_n 0.0479252f $X=7.945 $Y=2.595 $X2=0 $Y2=0
cc_272 N_A_84_209#_c_198_n N_A_c_752_n 6.21385e-19 $X=7.845 $Y=1.47 $X2=0 $Y2=0
cc_273 N_A_84_209#_M1010_g N_A_c_736_n 0.00660574f $X=7.795 $Y=0.915 $X2=0 $Y2=0
cc_274 N_A_84_209#_c_190_n N_A_c_739_n 0.00107752f $X=0.865 $Y=1.21 $X2=0 $Y2=0
cc_275 N_A_84_209#_c_191_n N_A_c_739_n 0.0136159f $X=0.865 $Y=1.21 $X2=0 $Y2=0
cc_276 N_A_84_209#_c_193_n N_A_c_740_n 0.00281668f $X=2.86 $Y=1.545 $X2=0 $Y2=0
cc_277 N_A_84_209#_c_224_p N_A_c_746_n 0.00317285f $X=4.89 $Y=0.915 $X2=0 $Y2=0
cc_278 N_A_84_209#_M1010_g N_A_c_747_n 0.018361f $X=7.795 $Y=0.915 $X2=0 $Y2=0
cc_279 N_A_84_209#_M1023_g N_A_1574_141#_c_912_n 0.00751144f $X=7.945 $Y=2.595
+ $X2=0 $Y2=0
cc_280 N_A_84_209#_M1023_g N_A_1574_141#_c_913_n 0.00423236f $X=7.945 $Y=2.595
+ $X2=0 $Y2=0
cc_281 N_A_84_209#_M1010_g N_A_1574_141#_c_904_n 0.00981734f $X=7.795 $Y=0.915
+ $X2=0 $Y2=0
cc_282 N_A_84_209#_c_189_n N_A_1574_141#_c_904_n 0.00319978f $X=7.945 $Y=1.76
+ $X2=0 $Y2=0
cc_283 N_A_84_209#_c_198_n N_A_1574_141#_c_904_n 0.00984148f $X=7.845 $Y=1.47
+ $X2=0 $Y2=0
cc_284 N_A_84_209#_M1018_g COUT 0.0102968f $X=0.595 $Y=0.635 $X2=0 $Y2=0
cc_285 N_A_84_209#_M1005_g COUT 0.00124947f $X=0.955 $Y=0.635 $X2=0 $Y2=0
cc_286 N_A_84_209#_c_191_n COUT 0.00341555f $X=0.865 $Y=1.21 $X2=0 $Y2=0
cc_287 N_A_84_209#_M1014_g COUT 0.0308438f $X=0.545 $Y=2.415 $X2=0 $Y2=0
cc_288 N_A_84_209#_M1018_g COUT 0.00736383f $X=0.595 $Y=0.635 $X2=0 $Y2=0
cc_289 N_A_84_209#_c_190_n COUT 0.0271129f $X=0.865 $Y=1.21 $X2=0 $Y2=0
cc_290 N_A_84_209#_c_191_n COUT 0.0273279f $X=0.865 $Y=1.21 $X2=0 $Y2=0
cc_291 N_A_84_209#_c_208_n COUT 0.00979969f $X=1.03 $Y=1.63 $X2=0 $Y2=0
cc_292 N_A_84_209#_M1014_g N_VPWR_c_1014_n 0.0278602f $X=0.545 $Y=2.415 $X2=0
+ $Y2=0
cc_293 N_A_84_209#_c_191_n N_VPWR_c_1014_n 0.00356371f $X=0.865 $Y=1.21 $X2=0
+ $Y2=0
cc_294 N_A_84_209#_c_208_n N_VPWR_c_1014_n 0.0233646f $X=1.03 $Y=1.63 $X2=0
+ $Y2=0
cc_295 N_A_84_209#_M1023_g N_VPWR_c_1023_n 0.0090344f $X=7.945 $Y=2.595 $X2=0
+ $Y2=0
cc_296 N_A_84_209#_M1011_d N_VPWR_c_1013_n 0.00225465f $X=3.555 $Y=2.095 $X2=0
+ $Y2=0
cc_297 N_A_84_209#_M1014_g N_VPWR_c_1013_n 0.00800793f $X=0.545 $Y=2.415 $X2=0
+ $Y2=0
cc_298 N_A_84_209#_M1023_g N_VPWR_c_1013_n 0.0154451f $X=7.945 $Y=2.595 $X2=0
+ $Y2=0
cc_299 N_A_84_209#_M1014_g N_VPWR_c_1028_n 0.00791861f $X=0.545 $Y=2.415 $X2=0
+ $Y2=0
cc_300 N_A_84_209#_M1014_g N_A_245_409#_c_1125_n 0.00198025f $X=0.545 $Y=2.415
+ $X2=0 $Y2=0
cc_301 N_A_84_209#_c_192_n N_A_245_409#_c_1126_n 0.0480591f $X=2.775 $Y=1.63
+ $X2=0 $Y2=0
cc_302 N_A_84_209#_M1014_g N_A_245_409#_c_1127_n 3.95513e-19 $X=0.545 $Y=2.415
+ $X2=0 $Y2=0
cc_303 N_A_84_209#_c_192_n N_A_245_409#_c_1127_n 0.0265557f $X=2.775 $Y=1.63
+ $X2=0 $Y2=0
cc_304 N_A_84_209#_c_192_n N_A_245_409#_c_1128_n 0.0153104f $X=2.775 $Y=1.63
+ $X2=0 $Y2=0
cc_305 N_A_84_209#_c_209_n N_A_245_409#_c_1128_n 0.0102347f $X=3.255 $Y=1.83
+ $X2=0 $Y2=0
cc_306 N_A_84_209#_c_199_n N_A_245_409#_c_1128_n 0.0143947f $X=2.86 $Y=1.63
+ $X2=0 $Y2=0
cc_307 N_A_84_209#_c_192_n N_A_245_409#_c_1130_n 0.0126154f $X=2.775 $Y=1.63
+ $X2=0 $Y2=0
cc_308 N_A_84_209#_c_199_n N_A_245_409#_c_1130_n 8.9643e-19 $X=2.86 $Y=1.63
+ $X2=0 $Y2=0
cc_309 N_A_84_209#_M1011_d N_A_458_409#_c_1169_n 0.00332313f $X=3.555 $Y=2.095
+ $X2=0 $Y2=0
cc_310 N_A_84_209#_c_221_p N_A_458_409#_c_1169_n 0.00813115f $X=3.425 $Y=2.582
+ $X2=0 $Y2=0
cc_311 N_A_84_209#_c_222_p N_A_458_409#_c_1169_n 0.0208086f $X=3.695 $Y=2.54
+ $X2=0 $Y2=0
cc_312 N_A_84_209#_c_222_p N_A_458_409#_c_1174_n 0.0138075f $X=3.695 $Y=2.54
+ $X2=0 $Y2=0
cc_313 N_A_84_209#_M1023_g N_A_1049_419#_c_1205_n 0.00423236f $X=7.945 $Y=2.595
+ $X2=0 $Y2=0
cc_314 N_A_84_209#_M1023_g N_A_1049_419#_c_1206_n 0.00751144f $X=7.945 $Y=2.595
+ $X2=0 $Y2=0
cc_315 N_A_84_209#_c_224_p N_VGND_M1015_d 0.00802243f $X=4.89 $Y=0.915 $X2=0
+ $Y2=0
cc_316 N_A_84_209#_M1018_g N_VGND_c_1263_n 0.00179293f $X=0.595 $Y=0.635 $X2=0
+ $Y2=0
cc_317 N_A_84_209#_M1005_g N_VGND_c_1263_n 0.00779381f $X=0.955 $Y=0.635 $X2=0
+ $Y2=0
cc_318 N_A_84_209#_M1005_g N_VGND_c_1264_n 0.00436629f $X=0.955 $Y=0.635 $X2=0
+ $Y2=0
cc_319 N_A_84_209#_c_190_n N_VGND_c_1264_n 0.00622446f $X=0.865 $Y=1.21 $X2=0
+ $Y2=0
cc_320 N_A_84_209#_c_192_n N_VGND_c_1265_n 0.072159f $X=2.775 $Y=1.63 $X2=0
+ $Y2=0
cc_321 N_A_84_209#_c_193_n N_VGND_c_1265_n 0.0135588f $X=2.86 $Y=1.545 $X2=0
+ $Y2=0
cc_322 N_A_84_209#_c_190_n N_VGND_c_1266_n 0.00796091f $X=0.865 $Y=1.21 $X2=0
+ $Y2=0
cc_323 N_A_84_209#_c_191_n N_VGND_c_1266_n 0.00158326f $X=0.865 $Y=1.21 $X2=0
+ $Y2=0
cc_324 N_A_84_209#_c_192_n N_VGND_c_1266_n 0.0132443f $X=2.775 $Y=1.63 $X2=0
+ $Y2=0
cc_325 N_A_84_209#_c_193_n N_VGND_c_1267_n 0.00994785f $X=2.86 $Y=1.545 $X2=0
+ $Y2=0
cc_326 N_A_84_209#_c_291_p N_VGND_c_1267_n 0.0177344f $X=2.945 $Y=0.942 $X2=0
+ $Y2=0
cc_327 N_A_84_209#_c_194_n N_VGND_c_1267_n 0.00389014f $X=3.605 $Y=0.915 $X2=0
+ $Y2=0
cc_328 N_A_84_209#_c_224_p N_VGND_c_1268_n 0.0248851f $X=4.89 $Y=0.915 $X2=0
+ $Y2=0
cc_329 N_A_84_209#_M1005_g N_VGND_c_1271_n 0.00548338f $X=0.955 $Y=0.635 $X2=0
+ $Y2=0
cc_330 N_A_84_209#_c_190_n N_VGND_c_1271_n 0.00185662f $X=0.865 $Y=1.21 $X2=0
+ $Y2=0
cc_331 N_A_84_209#_M1018_g N_VGND_c_1274_n 0.00514022f $X=0.595 $Y=0.635 $X2=0
+ $Y2=0
cc_332 N_A_84_209#_M1005_g N_VGND_c_1274_n 0.00447026f $X=0.955 $Y=0.635 $X2=0
+ $Y2=0
cc_333 N_A_84_209#_M1018_g N_VGND_c_1278_n 0.00528353f $X=0.595 $Y=0.635 $X2=0
+ $Y2=0
cc_334 N_A_84_209#_M1005_g N_VGND_c_1278_n 0.00443817f $X=0.955 $Y=0.635 $X2=0
+ $Y2=0
cc_335 N_A_84_209#_M1010_g N_VGND_c_1278_n 9.68004e-19 $X=7.795 $Y=0.915 $X2=0
+ $Y2=0
cc_336 N_A_84_209#_c_224_p N_VGND_c_1278_n 0.0176895f $X=4.89 $Y=0.915 $X2=0
+ $Y2=0
cc_337 N_A_84_209#_c_224_p N_A_355_141#_M1002_d 0.00738232f $X=4.89 $Y=0.915
+ $X2=0 $Y2=0
cc_338 N_A_84_209#_c_213_p N_A_355_141#_c_1392_n 0.0111998f $X=3.25 $Y=0.942
+ $X2=0 $Y2=0
cc_339 N_A_84_209#_c_291_p N_A_355_141#_c_1392_n 0.00566421f $X=2.945 $Y=0.942
+ $X2=0 $Y2=0
cc_340 N_A_84_209#_c_224_p N_A_355_141#_c_1392_n 0.00966425f $X=4.89 $Y=0.915
+ $X2=0 $Y2=0
cc_341 N_A_84_209#_c_194_n N_A_355_141#_c_1392_n 0.0234966f $X=3.605 $Y=0.915
+ $X2=0 $Y2=0
cc_342 N_A_84_209#_c_224_p N_A_355_141#_c_1394_n 0.0234417f $X=4.89 $Y=0.915
+ $X2=0 $Y2=0
cc_343 N_A_84_209#_c_193_n A_577_141# 8.05715e-19 $X=2.86 $Y=1.545 $X2=-0.19
+ $Y2=-0.245
cc_344 N_A_84_209#_c_213_p A_577_141# 0.00643501f $X=3.25 $Y=0.942 $X2=-0.19
+ $Y2=-0.245
cc_345 N_A_84_209#_c_196_n N_A_1005_141#_c_1431_n 0.0487289f $X=6.45 $Y=1.55
+ $X2=0 $Y2=0
cc_346 N_A_84_209#_c_195_n N_A_1005_141#_c_1432_n 0.0133676f $X=4.975 $Y=1.465
+ $X2=0 $Y2=0
cc_347 N_A_84_209#_c_196_n N_A_1005_141#_c_1432_n 0.0137879f $X=6.45 $Y=1.55
+ $X2=0 $Y2=0
cc_348 N_A_84_209#_c_196_n N_A_1005_141#_c_1439_n 0.00669981f $X=6.45 $Y=1.55
+ $X2=0 $Y2=0
cc_349 N_A_84_209#_c_200_n N_A_1005_141#_c_1439_n 0.012909f $X=6.535 $Y=1.285
+ $X2=0 $Y2=0
cc_350 N_A_84_209#_c_201_n N_A_1005_141#_c_1439_n 0.0544155f $X=7.26 $Y=1.417
+ $X2=0 $Y2=0
cc_351 N_A_84_209#_c_196_n N_A_1005_141#_c_1434_n 0.0131356f $X=6.45 $Y=1.55
+ $X2=0 $Y2=0
cc_352 N_A_84_209#_c_200_n N_A_1005_141#_c_1434_n 0.00614786f $X=6.535 $Y=1.285
+ $X2=0 $Y2=0
cc_353 N_A_84_209#_M1010_g N_A_1005_141#_c_1435_n 0.00494775f $X=7.795 $Y=0.915
+ $X2=0 $Y2=0
cc_354 N_A_84_209#_c_198_n N_A_1005_141#_c_1435_n 0.0141931f $X=7.845 $Y=1.47
+ $X2=0 $Y2=0
cc_355 N_A_84_209#_c_202_n N_A_1005_141#_c_1435_n 0.00103143f $X=7.43 $Y=1.417
+ $X2=0 $Y2=0
cc_356 N_B_c_382_n N_CIN_c_574_n 0.0140925f $X=3.2 $Y=1.235 $X2=-0.19 $Y2=-0.245
cc_357 N_B_c_384_n N_CIN_c_574_n 0.0178471f $X=4.36 $Y=1.2 $X2=-0.19 $Y2=-0.245
cc_358 N_B_M1011_g N_CIN_M1027_g 0.0270539f $X=3.43 $Y=2.595 $X2=0 $Y2=0
cc_359 N_B_c_405_n N_CIN_M1027_g 0.0352107f $X=4.59 $Y=1.945 $X2=0 $Y2=0
cc_360 N_B_c_440_n N_CIN_M1027_g 0.0165985f $X=4.04 $Y=2.217 $X2=0 $Y2=0
cc_361 N_B_c_441_n N_CIN_M1027_g 0.00677919f $X=4.21 $Y=2.217 $X2=0 $Y2=0
cc_362 N_B_c_386_n N_CIN_M1004_g 0.0105472f $X=4.95 $Y=1.2 $X2=0 $Y2=0
cc_363 N_B_c_403_n N_CIN_M1028_g 0.0240782f $X=5.12 $Y=2.02 $X2=0 $Y2=0
cc_364 N_B_c_438_n N_CIN_M1028_g 0.0170819f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_365 N_B_c_387_n N_CIN_M1022_g 0.0426498f $X=8.745 $Y=1.215 $X2=0 $Y2=0
cc_366 N_B_c_397_n N_CIN_M1022_g 0.00816644f $X=8.985 $Y=1.605 $X2=0 $Y2=0
cc_367 N_B_M1025_g N_CIN_M1009_g 0.0741666f $X=8.965 $Y=2.595 $X2=0 $Y2=0
cc_368 N_B_c_438_n N_CIN_M1009_g 0.0146919f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_369 N_B_c_392_n N_CIN_M1009_g 0.00277055f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_370 N_B_c_383_n N_CIN_c_577_n 0.00632664f $X=3.43 $Y=1.715 $X2=0 $Y2=0
cc_371 N_B_c_391_n N_CIN_c_577_n 0.00674779f $X=4.435 $Y=1.32 $X2=0 $Y2=0
cc_372 N_B_c_394_n N_CIN_c_577_n 0.00543898f $X=3.69 $Y=1.4 $X2=0 $Y2=0
cc_373 B N_CIN_c_577_n 2.60362e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_374 N_B_c_396_n N_CIN_c_577_n 0.00659214f $X=4.6 $Y=1.4 $X2=0 $Y2=0
cc_375 N_B_c_402_n N_CIN_c_578_n 0.0240782f $X=4.995 $Y=1.945 $X2=0 $Y2=0
cc_376 N_B_c_396_n N_CIN_c_578_n 0.0105472f $X=4.6 $Y=1.4 $X2=0 $Y2=0
cc_377 N_B_c_385_n N_CIN_c_590_n 0.00117564f $X=4.54 $Y=1.87 $X2=0 $Y2=0
cc_378 N_B_c_402_n N_CIN_c_590_n 0.0186344f $X=4.995 $Y=1.945 $X2=0 $Y2=0
cc_379 N_B_c_405_n N_CIN_c_590_n 0.00435122f $X=4.59 $Y=1.945 $X2=0 $Y2=0
cc_380 N_B_c_438_n N_CIN_c_590_n 0.143814f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_381 B N_CIN_c_590_n 0.00828328f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_382 N_B_c_396_n N_CIN_c_590_n 0.00432183f $X=4.6 $Y=1.4 $X2=0 $Y2=0
cc_383 N_B_c_385_n N_CIN_c_579_n 0.00776182f $X=4.54 $Y=1.87 $X2=0 $Y2=0
cc_384 N_B_c_405_n N_CIN_c_579_n 0.00339124f $X=4.59 $Y=1.945 $X2=0 $Y2=0
cc_385 N_B_c_390_n N_CIN_c_579_n 0.0265669f $X=3.69 $Y=2.1 $X2=0 $Y2=0
cc_386 N_B_c_391_n N_CIN_c_579_n 0.0287842f $X=4.435 $Y=1.32 $X2=0 $Y2=0
cc_387 N_B_c_438_n N_CIN_c_579_n 0.0200725f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_388 N_B_c_440_n N_CIN_c_579_n 0.0159528f $X=4.04 $Y=2.217 $X2=0 $Y2=0
cc_389 B N_CIN_c_579_n 0.00877784f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_390 N_B_c_396_n N_CIN_c_579_n 0.00102515f $X=4.6 $Y=1.4 $X2=0 $Y2=0
cc_391 N_B_c_438_n N_CIN_c_592_n 0.0741149f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_392 N_B_c_383_n N_CIN_c_580_n 0.0270539f $X=3.43 $Y=1.715 $X2=0 $Y2=0
cc_393 N_B_c_385_n N_CIN_c_580_n 0.0178371f $X=4.54 $Y=1.87 $X2=0 $Y2=0
cc_394 N_B_c_391_n N_CIN_c_580_n 0.00165219f $X=4.435 $Y=1.32 $X2=0 $Y2=0
cc_395 N_B_c_441_n N_CIN_c_580_n 7.53603e-19 $X=4.21 $Y=2.217 $X2=0 $Y2=0
cc_396 N_B_c_438_n N_CIN_c_581_n 0.0209544f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_397 N_B_c_392_n N_CIN_c_581_n 0.0244151f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_398 N_B_c_393_n N_CIN_c_581_n 0.00114936f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_399 N_B_c_438_n N_CIN_c_582_n 2.98577e-19 $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_400 N_B_c_392_n N_CIN_c_582_n 0.00114961f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_401 N_B_c_393_n N_CIN_c_582_n 0.0201104f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_402 N_B_c_438_n CIN 0.021361f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_403 N_B_c_438_n N_CIN_c_584_n 0.00754888f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_404 N_B_c_383_n N_CIN_c_585_n 0.00638099f $X=3.43 $Y=1.715 $X2=0 $Y2=0
cc_405 N_B_c_385_n N_CIN_c_585_n 7.14372e-19 $X=4.54 $Y=1.87 $X2=0 $Y2=0
cc_406 N_B_c_390_n N_CIN_c_585_n 0.00685829f $X=3.69 $Y=2.1 $X2=0 $Y2=0
cc_407 N_B_c_391_n N_CIN_c_585_n 0.0081418f $X=4.435 $Y=1.32 $X2=0 $Y2=0
cc_408 N_B_c_394_n N_CIN_c_585_n 0.00275315f $X=3.69 $Y=1.4 $X2=0 $Y2=0
cc_409 B N_CIN_c_585_n 6.28208e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_410 N_B_c_396_n N_CIN_c_585_n 0.00535795f $X=4.6 $Y=1.4 $X2=0 $Y2=0
cc_411 N_B_c_382_n N_A_M1020_g 0.035969f $X=3.2 $Y=1.235 $X2=0 $Y2=0
cc_412 N_B_c_438_n N_A_c_752_n 0.0170819f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_413 N_B_c_387_n N_A_c_736_n 0.00673512f $X=8.745 $Y=1.215 $X2=0 $Y2=0
cc_414 N_B_c_387_n N_A_M1013_g 0.0169715f $X=8.745 $Y=1.215 $X2=0 $Y2=0
cc_415 N_B_M1025_g N_A_M1017_g 0.0636383f $X=8.965 $Y=2.595 $X2=0 $Y2=0
cc_416 N_B_c_392_n N_A_M1017_g 9.24329e-19 $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_417 N_B_c_393_n N_A_M1017_g 0.0205836f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_418 N_B_c_397_n N_A_M1017_g 0.00718057f $X=8.985 $Y=1.605 $X2=0 $Y2=0
cc_419 N_B_c_387_n N_A_c_743_n 0.0083899f $X=8.745 $Y=1.215 $X2=0 $Y2=0
cc_420 N_B_c_388_n N_A_c_744_n 0.00832349f $X=8.925 $Y=1.29 $X2=0 $Y2=0
cc_421 N_B_c_382_n N_A_c_746_n 0.00491612f $X=3.2 $Y=1.235 $X2=0 $Y2=0
cc_422 N_B_c_384_n N_A_c_746_n 0.00611177f $X=4.36 $Y=1.2 $X2=0 $Y2=0
cc_423 N_B_c_386_n N_A_c_746_n 0.00611071f $X=4.95 $Y=1.2 $X2=0 $Y2=0
cc_424 N_B_c_438_n N_A_1574_141#_M1023_d 0.00358198f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_425 N_B_M1025_g N_A_1574_141#_c_912_n 0.00164029f $X=8.965 $Y=2.595 $X2=0
+ $Y2=0
cc_426 N_B_c_388_n N_A_1574_141#_c_901_n 0.0226471f $X=8.925 $Y=1.29 $X2=0 $Y2=0
cc_427 N_B_c_392_n N_A_1574_141#_c_901_n 0.0203656f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_428 N_B_c_393_n N_A_1574_141#_c_901_n 0.00149607f $X=8.985 $Y=1.77 $X2=0
+ $Y2=0
cc_429 N_B_c_397_n N_A_1574_141#_c_901_n 0.00333259f $X=8.985 $Y=1.605 $X2=0
+ $Y2=0
cc_430 N_B_M1025_g N_A_1574_141#_c_923_n 0.0168956f $X=8.965 $Y=2.595 $X2=0
+ $Y2=0
cc_431 N_B_c_438_n N_A_1574_141#_c_923_n 0.0414917f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_432 N_B_c_393_n N_A_1574_141#_c_923_n 2.45226e-19 $X=8.985 $Y=1.77 $X2=0
+ $Y2=0
cc_433 N_B_c_438_n N_A_1574_141#_c_913_n 0.0162949f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_434 N_B_M1025_g N_A_1574_141#_c_902_n 6.33721e-19 $X=8.965 $Y=2.595 $X2=0
+ $Y2=0
cc_435 N_B_c_392_n N_A_1574_141#_c_902_n 0.0357316f $X=8.985 $Y=1.77 $X2=0 $Y2=0
cc_436 N_B_c_393_n N_A_1574_141#_c_902_n 0.00179708f $X=8.985 $Y=1.77 $X2=0
+ $Y2=0
cc_437 N_B_c_397_n N_A_1574_141#_c_902_n 0.00385914f $X=8.985 $Y=1.605 $X2=0
+ $Y2=0
cc_438 N_B_c_387_n N_A_1574_141#_c_904_n 0.00297076f $X=8.745 $Y=1.215 $X2=0
+ $Y2=0
cc_439 N_B_c_438_n N_VPWR_M1016_d 0.00331357f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_440 N_B_c_438_n N_VPWR_M1028_d 0.0386431f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_441 N_B_c_401_n N_VPWR_c_1016_n 0.0169043f $X=4.59 $Y=2.02 $X2=0 $Y2=0
cc_442 N_B_c_403_n N_VPWR_c_1016_n 0.0174655f $X=5.12 $Y=2.02 $X2=0 $Y2=0
cc_443 N_B_c_438_n N_VPWR_c_1016_n 0.0164319f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_444 N_B_c_403_n N_VPWR_c_1017_n 0.00106763f $X=5.12 $Y=2.02 $X2=0 $Y2=0
cc_445 N_B_M1011_g N_VPWR_c_1021_n 0.00599941f $X=3.43 $Y=2.595 $X2=0 $Y2=0
cc_446 N_B_c_401_n N_VPWR_c_1021_n 0.008763f $X=4.59 $Y=2.02 $X2=0 $Y2=0
cc_447 N_B_M1025_g N_VPWR_c_1023_n 0.00710941f $X=8.965 $Y=2.595 $X2=0 $Y2=0
cc_448 N_B_c_403_n N_VPWR_c_1025_n 0.00840199f $X=5.12 $Y=2.02 $X2=0 $Y2=0
cc_449 N_B_M1011_g N_VPWR_c_1013_n 0.00935477f $X=3.43 $Y=2.595 $X2=0 $Y2=0
cc_450 N_B_c_401_n N_VPWR_c_1013_n 0.0148063f $X=4.59 $Y=2.02 $X2=0 $Y2=0
cc_451 N_B_c_403_n N_VPWR_c_1013_n 0.0136763f $X=5.12 $Y=2.02 $X2=0 $Y2=0
cc_452 N_B_M1025_g N_VPWR_c_1013_n 0.00886776f $X=8.965 $Y=2.595 $X2=0 $Y2=0
cc_453 N_B_M1011_g N_A_245_409#_c_1128_n 0.00117132f $X=3.43 $Y=2.595 $X2=0
+ $Y2=0
cc_454 N_B_M1011_g N_A_245_409#_c_1129_n 0.00285467f $X=3.43 $Y=2.595 $X2=0
+ $Y2=0
cc_455 N_B_c_438_n N_A_458_409#_M1027_d 0.00524856f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_456 N_B_c_441_n N_A_458_409#_M1027_d 0.00225826f $X=4.21 $Y=2.217 $X2=0 $Y2=0
cc_457 N_B_M1011_g N_A_458_409#_c_1169_n 0.0158203f $X=3.43 $Y=2.595 $X2=0 $Y2=0
cc_458 N_B_c_401_n N_A_458_409#_c_1169_n 0.00205525f $X=4.59 $Y=2.02 $X2=0 $Y2=0
cc_459 N_B_c_440_n N_A_458_409#_c_1169_n 0.00412823f $X=4.04 $Y=2.217 $X2=0
+ $Y2=0
cc_460 N_B_c_441_n N_A_458_409#_c_1169_n 5.08945e-19 $X=4.21 $Y=2.217 $X2=0
+ $Y2=0
cc_461 N_B_M1011_g N_A_458_409#_c_1174_n 7.3358e-19 $X=3.43 $Y=2.595 $X2=0 $Y2=0
cc_462 N_B_c_401_n N_A_458_409#_c_1174_n 0.00420124f $X=4.59 $Y=2.02 $X2=0 $Y2=0
cc_463 N_B_c_441_n N_A_458_409#_c_1174_n 0.0207636f $X=4.21 $Y=2.217 $X2=0 $Y2=0
cc_464 N_B_c_438_n N_A_1049_419#_M1000_d 0.00358644f $X=8.82 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_465 N_B_c_438_n N_A_1049_419#_M1003_d 0.00352464f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_466 N_B_c_403_n N_A_1049_419#_c_1209_n 0.00751144f $X=5.12 $Y=2.02 $X2=0
+ $Y2=0
cc_467 N_B_c_438_n N_A_1049_419#_c_1205_n 0.142891f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_468 N_B_c_403_n N_A_1049_419#_c_1211_n 0.00423889f $X=5.12 $Y=2.02 $X2=0
+ $Y2=0
cc_469 N_B_c_438_n N_A_1049_419#_c_1211_n 0.0162949f $X=8.82 $Y=2.25 $X2=0 $Y2=0
cc_470 N_B_c_438_n A_1720_419# 0.00618276f $X=8.82 $Y=2.25 $X2=-0.19 $Y2=-0.245
cc_471 N_B_c_384_n N_VGND_c_1268_n 8.19597e-19 $X=4.36 $Y=1.2 $X2=0 $Y2=0
cc_472 N_B_c_386_n N_VGND_c_1268_n 8.19597e-19 $X=4.95 $Y=1.2 $X2=0 $Y2=0
cc_473 N_B_c_387_n N_VGND_c_1270_n 9.32276e-19 $X=8.745 $Y=1.215 $X2=0 $Y2=0
cc_474 N_B_c_384_n N_VGND_c_1278_n 9.68004e-19 $X=4.36 $Y=1.2 $X2=0 $Y2=0
cc_475 N_B_c_386_n N_VGND_c_1278_n 9.68003e-19 $X=4.95 $Y=1.2 $X2=0 $Y2=0
cc_476 N_B_c_387_n N_VGND_c_1278_n 9.68004e-19 $X=8.745 $Y=1.215 $X2=0 $Y2=0
cc_477 N_B_c_382_n N_A_355_141#_c_1392_n 0.00163241f $X=3.2 $Y=1.235 $X2=0 $Y2=0
cc_478 N_B_c_384_n N_A_355_141#_c_1394_n 8.19597e-19 $X=4.36 $Y=1.2 $X2=0 $Y2=0
cc_479 N_B_c_386_n N_A_1005_141#_c_1430_n 0.00472369f $X=4.95 $Y=1.2 $X2=0 $Y2=0
cc_480 N_B_c_386_n N_A_1005_141#_c_1432_n 7.02148e-19 $X=4.95 $Y=1.2 $X2=0 $Y2=0
cc_481 N_B_c_386_n N_A_1005_141#_c_1433_n 8.19597e-19 $X=4.95 $Y=1.2 $X2=0 $Y2=0
cc_482 N_CIN_c_592_n N_A_M1008_g 0.00431006f $X=8.28 $Y=1.9 $X2=0 $Y2=0
cc_483 CIN N_A_M1008_g 0.00160564f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_484 N_CIN_c_584_n N_A_M1008_g 0.0221634f $X=6.915 $Y=1.755 $X2=0 $Y2=0
cc_485 N_CIN_c_592_n N_A_c_752_n 0.0104926f $X=8.28 $Y=1.9 $X2=0 $Y2=0
cc_486 CIN N_A_c_752_n 2.77228e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_487 N_CIN_M1022_g N_A_c_736_n 0.00630385f $X=8.355 $Y=0.915 $X2=0 $Y2=0
cc_488 N_CIN_c_574_n N_A_c_746_n 0.00491612f $X=3.77 $Y=1.2 $X2=0 $Y2=0
cc_489 N_CIN_M1004_g N_A_c_746_n 0.0065768f $X=5.54 $Y=0.915 $X2=0 $Y2=0
cc_490 N_CIN_M1009_g N_A_1574_141#_c_912_n 0.00861375f $X=8.475 $Y=2.595 $X2=0
+ $Y2=0
cc_491 N_CIN_M1022_g N_A_1574_141#_c_901_n 0.0069519f $X=8.355 $Y=0.915 $X2=0
+ $Y2=0
cc_492 N_CIN_c_581_n N_A_1574_141#_c_901_n 0.0156264f $X=8.445 $Y=1.77 $X2=0
+ $Y2=0
cc_493 N_CIN_c_582_n N_A_1574_141#_c_901_n 0.00118654f $X=8.445 $Y=1.77 $X2=0
+ $Y2=0
cc_494 N_CIN_M1009_g N_A_1574_141#_c_923_n 0.0136108f $X=8.475 $Y=2.595 $X2=0
+ $Y2=0
cc_495 N_CIN_M1009_g N_A_1574_141#_c_913_n 0.0016877f $X=8.475 $Y=2.595 $X2=0
+ $Y2=0
cc_496 N_CIN_M1022_g N_A_1574_141#_c_904_n 0.0182374f $X=8.355 $Y=0.915 $X2=0
+ $Y2=0
cc_497 N_CIN_c_592_n N_A_1574_141#_c_904_n 0.00403843f $X=8.28 $Y=1.9 $X2=0
+ $Y2=0
cc_498 N_CIN_c_581_n N_A_1574_141#_c_904_n 0.00531193f $X=8.445 $Y=1.77 $X2=0
+ $Y2=0
cc_499 N_CIN_M1027_g N_VPWR_c_1016_n 0.00109572f $X=3.96 $Y=2.595 $X2=0 $Y2=0
cc_500 N_CIN_M1028_g N_VPWR_c_1016_n 0.00118445f $X=5.65 $Y=2.595 $X2=0 $Y2=0
cc_501 N_CIN_M1028_g N_VPWR_c_1017_n 0.0103571f $X=5.65 $Y=2.595 $X2=0 $Y2=0
cc_502 N_CIN_M1027_g N_VPWR_c_1021_n 0.00599906f $X=3.96 $Y=2.595 $X2=0 $Y2=0
cc_503 N_CIN_M1009_g N_VPWR_c_1023_n 0.00701311f $X=8.475 $Y=2.595 $X2=0 $Y2=0
cc_504 N_CIN_M1028_g N_VPWR_c_1025_n 0.00629498f $X=5.65 $Y=2.595 $X2=0 $Y2=0
cc_505 N_CIN_M1027_g N_VPWR_c_1013_n 0.00820224f $X=3.96 $Y=2.595 $X2=0 $Y2=0
cc_506 N_CIN_M1028_g N_VPWR_c_1013_n 0.00702131f $X=5.65 $Y=2.595 $X2=0 $Y2=0
cc_507 N_CIN_M1009_g N_VPWR_c_1013_n 0.00878098f $X=8.475 $Y=2.595 $X2=0 $Y2=0
cc_508 N_CIN_M1027_g N_A_458_409#_c_1169_n 0.0150373f $X=3.96 $Y=2.595 $X2=0
+ $Y2=0
cc_509 N_CIN_M1027_g N_A_458_409#_c_1174_n 0.00834402f $X=3.96 $Y=2.595 $X2=0
+ $Y2=0
cc_510 N_CIN_M1028_g N_A_1049_419#_c_1209_n 0.0126416f $X=5.65 $Y=2.595 $X2=0
+ $Y2=0
cc_511 N_CIN_M1028_g N_A_1049_419#_c_1205_n 0.0157453f $X=5.65 $Y=2.595 $X2=0
+ $Y2=0
cc_512 N_CIN_M1028_g N_A_1049_419#_c_1211_n 0.0016877f $X=5.65 $Y=2.595 $X2=0
+ $Y2=0
cc_513 N_CIN_M1004_g N_VGND_c_1269_n 0.00708812f $X=5.54 $Y=0.915 $X2=0 $Y2=0
cc_514 N_CIN_M1004_g N_VGND_c_1278_n 8.13123e-19 $X=5.54 $Y=0.915 $X2=0 $Y2=0
cc_515 N_CIN_M1022_g N_VGND_c_1278_n 9.68004e-19 $X=8.355 $Y=0.915 $X2=0 $Y2=0
cc_516 N_CIN_c_574_n N_A_355_141#_c_1392_n 0.00167972f $X=3.77 $Y=1.2 $X2=0
+ $Y2=0
cc_517 N_CIN_c_574_n N_A_355_141#_c_1394_n 0.00218115f $X=3.77 $Y=1.2 $X2=0
+ $Y2=0
cc_518 N_CIN_M1004_g N_A_1005_141#_c_1431_n 0.0159448f $X=5.54 $Y=0.915 $X2=0
+ $Y2=0
cc_519 N_CIN_c_578_n N_A_1005_141#_c_1431_n 0.00256946f $X=5.465 $Y=1.48 $X2=0
+ $Y2=0
cc_520 N_CIN_c_584_n N_A_1005_141#_c_1439_n 0.00157801f $X=6.915 $Y=1.755 $X2=0
+ $Y2=0
cc_521 N_CIN_M1004_g N_A_1005_141#_c_1433_n 0.0037504f $X=5.54 $Y=0.915 $X2=0
+ $Y2=0
cc_522 N_CIN_M1004_g N_A_1005_141#_c_1434_n 0.00351859f $X=5.54 $Y=0.915 $X2=0
+ $Y2=0
cc_523 N_CIN_c_584_n N_A_1005_141#_c_1434_n 9.35709e-19 $X=6.915 $Y=1.755 $X2=0
+ $Y2=0
cc_524 N_A_c_736_n N_A_1574_141#_c_894_n 0.00827182f $X=9.145 $Y=0.18 $X2=0
+ $Y2=0
cc_525 N_A_c_742_n N_A_1574_141#_c_896_n 0.00998944f $X=9.315 $Y=0.9 $X2=0 $Y2=0
cc_526 N_A_M1017_g N_A_1574_141#_M1001_g 0.015773f $X=9.485 $Y=2.595 $X2=0 $Y2=0
cc_527 N_A_c_743_n N_A_1574_141#_c_898_n 0.006013f $X=9.425 $Y=1.215 $X2=0 $Y2=0
cc_528 N_A_M1017_g N_A_1574_141#_c_899_n 0.0207482f $X=9.485 $Y=2.595 $X2=0
+ $Y2=0
cc_529 N_A_c_742_n N_A_1574_141#_c_901_n 0.00356777f $X=9.315 $Y=0.9 $X2=0 $Y2=0
cc_530 N_A_c_744_n N_A_1574_141#_c_901_n 0.00587133f $X=9.425 $Y=1.365 $X2=0
+ $Y2=0
cc_531 N_A_M1017_g N_A_1574_141#_c_923_n 0.00820963f $X=9.485 $Y=2.595 $X2=0
+ $Y2=0
cc_532 N_A_M1017_g N_A_1574_141#_c_902_n 0.0297081f $X=9.485 $Y=2.595 $X2=0
+ $Y2=0
cc_533 N_A_M1017_g N_A_1574_141#_c_903_n 0.00596068f $X=9.485 $Y=2.595 $X2=0
+ $Y2=0
cc_534 N_A_c_744_n N_A_1574_141#_c_903_n 0.00475625f $X=9.425 $Y=1.365 $X2=0
+ $Y2=0
cc_535 N_A_c_736_n N_A_1574_141#_c_904_n 0.00579918f $X=9.145 $Y=0.18 $X2=0
+ $Y2=0
cc_536 N_A_M1017_g N_A_1574_141#_c_953_n 6.26406e-19 $X=9.485 $Y=2.595 $X2=0
+ $Y2=0
cc_537 N_A_c_744_n N_A_1574_141#_c_953_n 0.00611229f $X=9.425 $Y=1.365 $X2=0
+ $Y2=0
cc_538 N_A_M1017_g N_A_1574_141#_c_905_n 0.00181818f $X=9.485 $Y=2.595 $X2=0
+ $Y2=0
cc_539 N_A_c_744_n N_A_1574_141#_c_906_n 0.0207482f $X=9.425 $Y=1.365 $X2=0
+ $Y2=0
cc_540 N_A_M1029_g N_VPWR_c_1014_n 0.00431088f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_541 N_A_M1029_g N_VPWR_c_1015_n 0.0208668f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_542 N_A_M1021_g N_VPWR_c_1015_n 0.0256986f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_543 N_A_M1017_g N_VPWR_c_1018_n 0.00301415f $X=9.485 $Y=2.595 $X2=0 $Y2=0
cc_544 N_A_M1029_g N_VPWR_c_1019_n 0.00769046f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_545 N_A_M1021_g N_VPWR_c_1021_n 0.00767656f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_546 N_A_c_752_n N_VPWR_c_1023_n 0.00701311f $X=7.415 $Y=2 $X2=0 $Y2=0
cc_547 N_A_M1017_g N_VPWR_c_1023_n 0.00843169f $X=9.485 $Y=2.595 $X2=0 $Y2=0
cc_548 N_A_M1029_g N_VPWR_c_1013_n 0.0143431f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_549 N_A_M1021_g N_VPWR_c_1013_n 0.014306f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_550 N_A_c_752_n N_VPWR_c_1013_n 0.0102835f $X=7.415 $Y=2 $X2=0 $Y2=0
cc_551 N_A_M1017_g N_VPWR_c_1013_n 0.012855f $X=9.485 $Y=2.595 $X2=0 $Y2=0
cc_552 N_A_M1029_g N_A_245_409#_c_1125_n 0.0179336f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_553 N_A_M1021_g N_A_245_409#_c_1125_n 9.61614e-19 $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_554 N_A_M1029_g N_A_245_409#_c_1126_n 0.0178912f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_555 N_A_M1021_g N_A_245_409#_c_1126_n 0.017012f $X=2.165 $Y=2.545 $X2=0 $Y2=0
cc_556 N_A_M1029_g N_A_245_409#_c_1127_n 0.00378193f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_557 N_A_M1021_g N_A_245_409#_c_1128_n 9.8644e-19 $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_558 N_A_M1021_g N_A_245_409#_c_1129_n 0.00533849f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_559 N_A_M1029_g N_A_245_409#_c_1130_n 8.11481e-19 $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_560 N_A_M1021_g N_A_245_409#_c_1130_n 0.0134167f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_561 N_A_M1021_g N_A_458_409#_c_1168_n 0.0102071f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_562 N_A_M1021_g N_A_458_409#_c_1170_n 0.0059434f $X=2.165 $Y=2.545 $X2=0
+ $Y2=0
cc_563 N_A_c_752_n N_A_1049_419#_c_1205_n 0.0176783f $X=7.415 $Y=2 $X2=0 $Y2=0
cc_564 N_A_c_752_n N_A_1049_419#_c_1206_n 0.0180525f $X=7.415 $Y=2 $X2=0 $Y2=0
cc_565 N_A_c_727_n N_VGND_c_1263_n 0.0131084f $X=1.585 $Y=1.255 $X2=0 $Y2=0
cc_566 N_A_c_730_n N_VGND_c_1263_n 0.00930002f $X=1.66 $Y=0.18 $X2=0 $Y2=0
cc_567 N_A_M1019_g N_VGND_c_1263_n 0.00119534f $X=2.215 $Y=0.915 $X2=0 $Y2=0
cc_568 N_A_c_727_n N_VGND_c_1264_n 0.00948351f $X=1.585 $Y=1.255 $X2=0 $Y2=0
cc_569 N_A_c_727_n N_VGND_c_1265_n 0.00417405f $X=1.585 $Y=1.255 $X2=0 $Y2=0
cc_570 N_A_c_731_n N_VGND_c_1265_n 0.0102367f $X=2.04 $Y=1.33 $X2=0 $Y2=0
cc_571 N_A_M1019_g N_VGND_c_1265_n 0.00830626f $X=2.215 $Y=0.915 $X2=0 $Y2=0
cc_572 N_A_M1020_g N_VGND_c_1265_n 5.22374e-19 $X=2.81 $Y=0.915 $X2=0 $Y2=0
cc_573 N_A_c_739_n N_VGND_c_1265_n 0.00457393f $X=1.635 $Y=1.33 $X2=0 $Y2=0
cc_574 N_A_c_740_n N_VGND_c_1265_n 0.00843499f $X=2.165 $Y=1.33 $X2=0 $Y2=0
cc_575 N_A_c_727_n N_VGND_c_1266_n 9.56008e-19 $X=1.585 $Y=1.255 $X2=0 $Y2=0
cc_576 N_A_c_739_n N_VGND_c_1266_n 0.00275299f $X=1.635 $Y=1.33 $X2=0 $Y2=0
cc_577 N_A_c_727_n N_VGND_c_1267_n 7.22847e-19 $X=1.585 $Y=1.255 $X2=0 $Y2=0
cc_578 N_A_M1019_g N_VGND_c_1267_n 0.00979267f $X=2.215 $Y=0.915 $X2=0 $Y2=0
cc_579 N_A_M1020_g N_VGND_c_1267_n 0.00498019f $X=2.81 $Y=0.915 $X2=0 $Y2=0
cc_580 N_A_c_746_n N_VGND_c_1268_n 0.0252872f $X=6.905 $Y=0.35 $X2=0 $Y2=0
cc_581 N_A_c_746_n N_VGND_c_1269_n 0.0257761f $X=6.905 $Y=0.35 $X2=0 $Y2=0
cc_582 N_A_c_748_n N_VGND_c_1269_n 0.0101612f $X=6.905 $Y=0.555 $X2=0 $Y2=0
cc_583 N_A_c_736_n N_VGND_c_1270_n 0.00716616f $X=9.145 $Y=0.18 $X2=0 $Y2=0
cc_584 N_A_M1013_g N_VGND_c_1270_n 0.0195749f $X=9.22 $Y=0.54 $X2=0 $Y2=0
cc_585 N_A_c_742_n N_VGND_c_1270_n 0.00335009f $X=9.315 $Y=0.9 $X2=0 $Y2=0
cc_586 N_A_c_744_n N_VGND_c_1270_n 0.00470622f $X=9.425 $Y=1.365 $X2=0 $Y2=0
cc_587 N_A_c_727_n N_VGND_c_1271_n 0.00871212f $X=1.585 $Y=1.255 $X2=0 $Y2=0
cc_588 N_A_c_746_n N_VGND_c_1272_n 0.0224546f $X=6.905 $Y=0.35 $X2=0 $Y2=0
cc_589 N_A_c_730_n N_VGND_c_1275_n 0.0693424f $X=1.66 $Y=0.18 $X2=0 $Y2=0
cc_590 N_A_c_745_n N_VGND_c_1276_n 0.0202218f $X=7.07 $Y=0.43 $X2=0 $Y2=0
cc_591 N_A_c_746_n N_VGND_c_1276_n 0.102117f $X=6.905 $Y=0.35 $X2=0 $Y2=0
cc_592 N_A_c_748_n N_VGND_c_1276_n 0.016303f $X=6.905 $Y=0.555 $X2=0 $Y2=0
cc_593 N_A_c_729_n N_VGND_c_1278_n 0.0288382f $X=2.735 $Y=0.18 $X2=0 $Y2=0
cc_594 N_A_c_730_n N_VGND_c_1278_n 0.00506533f $X=1.66 $Y=0.18 $X2=0 $Y2=0
cc_595 N_A_c_736_n N_VGND_c_1278_n 0.0751547f $X=9.145 $Y=0.18 $X2=0 $Y2=0
cc_596 N_A_c_741_n N_VGND_c_1278_n 0.00373782f $X=2.81 $Y=0.18 $X2=0 $Y2=0
cc_597 N_A_c_745_n N_VGND_c_1278_n 0.0110116f $X=7.07 $Y=0.43 $X2=0 $Y2=0
cc_598 N_A_c_746_n N_VGND_c_1278_n 0.0923818f $X=6.905 $Y=0.35 $X2=0 $Y2=0
cc_599 N_A_c_747_n N_VGND_c_1278_n 0.0142265f $X=7.44 $Y=0.35 $X2=0 $Y2=0
cc_600 N_A_c_748_n N_VGND_c_1278_n 0.0158949f $X=6.905 $Y=0.555 $X2=0 $Y2=0
cc_601 N_A_c_727_n N_A_355_141#_c_1391_n 0.00590077f $X=1.585 $Y=1.255 $X2=0
+ $Y2=0
cc_602 N_A_M1019_g N_A_355_141#_c_1391_n 0.00550334f $X=2.215 $Y=0.915 $X2=0
+ $Y2=0
cc_603 N_A_M1020_g N_A_355_141#_c_1391_n 0.00214849f $X=2.81 $Y=0.915 $X2=0
+ $Y2=0
cc_604 N_A_c_739_n N_A_355_141#_c_1391_n 0.00196411f $X=1.635 $Y=1.33 $X2=0
+ $Y2=0
cc_605 N_A_c_729_n N_A_355_141#_c_1392_n 0.010501f $X=2.735 $Y=0.18 $X2=0 $Y2=0
cc_606 N_A_M1019_g N_A_355_141#_c_1392_n 0.00342153f $X=2.215 $Y=0.915 $X2=0
+ $Y2=0
cc_607 N_A_M1020_g N_A_355_141#_c_1392_n 0.016153f $X=2.81 $Y=0.915 $X2=0 $Y2=0
cc_608 N_A_c_746_n N_A_355_141#_c_1392_n 0.0166039f $X=6.905 $Y=0.35 $X2=0 $Y2=0
cc_609 N_A_c_727_n N_A_355_141#_c_1393_n 0.00320362f $X=1.585 $Y=1.255 $X2=0
+ $Y2=0
cc_610 N_A_c_729_n N_A_355_141#_c_1393_n 0.00791974f $X=2.735 $Y=0.18 $X2=0
+ $Y2=0
cc_611 N_A_c_746_n N_A_355_141#_c_1394_n 0.00761373f $X=6.905 $Y=0.35 $X2=0
+ $Y2=0
cc_612 N_A_M1008_g N_A_1005_141#_c_1439_n 0.0113171f $X=7.365 $Y=0.915 $X2=0
+ $Y2=0
cc_613 N_A_c_745_n N_A_1005_141#_c_1439_n 0.0243847f $X=7.07 $Y=0.43 $X2=0 $Y2=0
cc_614 N_A_c_746_n N_A_1005_141#_c_1439_n 0.00257451f $X=6.905 $Y=0.35 $X2=0
+ $Y2=0
cc_615 N_A_c_747_n N_A_1005_141#_c_1439_n 0.00186776f $X=7.44 $Y=0.35 $X2=0
+ $Y2=0
cc_616 N_A_c_748_n N_A_1005_141#_c_1439_n 0.0381778f $X=6.905 $Y=0.555 $X2=0
+ $Y2=0
cc_617 N_A_c_746_n N_A_1005_141#_c_1433_n 0.00775351f $X=6.905 $Y=0.35 $X2=0
+ $Y2=0
cc_618 N_A_c_746_n N_A_1005_141#_c_1434_n 0.00415742f $X=6.905 $Y=0.35 $X2=0
+ $Y2=0
cc_619 N_A_M1008_g N_A_1005_141#_c_1435_n 0.00926578f $X=7.365 $Y=0.915 $X2=0
+ $Y2=0
cc_620 N_A_c_736_n N_A_1005_141#_c_1435_n 0.00343986f $X=9.145 $Y=0.18 $X2=0
+ $Y2=0
cc_621 N_A_1574_141#_M1001_g N_VPWR_c_1018_n 0.0233718f $X=10.015 $Y=2.595 $X2=0
+ $Y2=0
cc_622 N_A_1574_141#_c_909_n N_VPWR_c_1018_n 5.34541e-19 $X=9.985 $Y=1.89 $X2=0
+ $Y2=0
cc_623 N_A_1574_141#_c_902_n N_VPWR_c_1018_n 0.0149392f $X=9.4 $Y=2.515 $X2=0
+ $Y2=0
cc_624 N_A_1574_141#_c_905_n N_VPWR_c_1018_n 0.00765767f $X=9.985 $Y=1.385 $X2=0
+ $Y2=0
cc_625 N_A_1574_141#_c_912_n N_VPWR_c_1023_n 0.0176422f $X=8.21 $Y=2.79 $X2=0
+ $Y2=0
cc_626 N_A_1574_141#_c_923_n N_VPWR_c_1023_n 0.0167557f $X=9.315 $Y=2.6 $X2=0
+ $Y2=0
cc_627 N_A_1574_141#_M1001_g N_VPWR_c_1026_n 0.00840199f $X=10.015 $Y=2.595
+ $X2=0 $Y2=0
cc_628 N_A_1574_141#_M1023_d N_VPWR_c_1013_n 0.0022543f $X=8.07 $Y=2.095 $X2=0
+ $Y2=0
cc_629 N_A_1574_141#_M1001_g N_VPWR_c_1013_n 0.0145244f $X=10.015 $Y=2.595 $X2=0
+ $Y2=0
cc_630 N_A_1574_141#_c_912_n N_VPWR_c_1013_n 0.0123981f $X=8.21 $Y=2.79 $X2=0
+ $Y2=0
cc_631 N_A_1574_141#_c_923_n N_VPWR_c_1013_n 0.0287336f $X=9.315 $Y=2.6 $X2=0
+ $Y2=0
cc_632 N_A_1574_141#_c_913_n N_A_1049_419#_c_1205_n 0.0126166f $X=8.375 $Y=2.6
+ $X2=0 $Y2=0
cc_633 N_A_1574_141#_c_912_n N_A_1049_419#_c_1206_n 0.0249726f $X=8.21 $Y=2.79
+ $X2=0 $Y2=0
cc_634 N_A_1574_141#_c_923_n A_1720_419# 0.0035945f $X=9.315 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_635 N_A_1574_141#_c_923_n A_1818_419# 0.00858555f $X=9.315 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_636 N_A_1574_141#_M1001_g N_SUM_c_1242_n 0.0240298f $X=10.015 $Y=2.595 $X2=0
+ $Y2=0
cc_637 N_A_1574_141#_c_909_n N_SUM_c_1242_n 4.72208e-19 $X=9.985 $Y=1.89 $X2=0
+ $Y2=0
cc_638 N_A_1574_141#_M1001_g N_SUM_c_1239_n 0.004938f $X=10.015 $Y=2.595 $X2=0
+ $Y2=0
cc_639 N_A_1574_141#_c_898_n N_SUM_c_1239_n 0.00448208f $X=9.985 $Y=1.22 $X2=0
+ $Y2=0
cc_640 N_A_1574_141#_c_905_n N_SUM_c_1239_n 0.0486291f $X=9.985 $Y=1.385 $X2=0
+ $Y2=0
cc_641 N_A_1574_141#_c_906_n N_SUM_c_1239_n 0.0154176f $X=9.985 $Y=1.385 $X2=0
+ $Y2=0
cc_642 N_A_1574_141#_c_894_n SUM 0.00156037f $X=9.705 $Y=0.825 $X2=0 $Y2=0
cc_643 N_A_1574_141#_c_897_n SUM 0.0114628f $X=10.065 $Y=0.825 $X2=0 $Y2=0
cc_644 N_A_1574_141#_c_900_n SUM 0.00251815f $X=10.065 $Y=0.9 $X2=0 $Y2=0
cc_645 N_A_1574_141#_c_898_n SUM 0.0053642f $X=9.985 $Y=1.22 $X2=0 $Y2=0
cc_646 N_A_1574_141#_c_900_n SUM 0.00762252f $X=10.065 $Y=0.9 $X2=0 $Y2=0
cc_647 N_A_1574_141#_c_906_n SUM 4.74761e-19 $X=9.985 $Y=1.385 $X2=0 $Y2=0
cc_648 N_A_1574_141#_c_894_n N_VGND_c_1270_n 0.00362216f $X=9.705 $Y=0.825 $X2=0
+ $Y2=0
cc_649 N_A_1574_141#_c_901_n N_VGND_c_1270_n 0.00159286f $X=9.315 $Y=1.305 $X2=0
+ $Y2=0
cc_650 N_A_1574_141#_c_903_n N_VGND_c_1270_n 0.00444822f $X=9.82 $Y=1.305 $X2=0
+ $Y2=0
cc_651 N_A_1574_141#_c_953_n N_VGND_c_1270_n 0.00727853f $X=9.4 $Y=1.305 $X2=0
+ $Y2=0
cc_652 N_A_1574_141#_c_904_n N_VGND_c_1276_n 0.00673673f $X=8.14 $Y=0.905 $X2=0
+ $Y2=0
cc_653 N_A_1574_141#_c_894_n N_VGND_c_1277_n 0.00495161f $X=9.705 $Y=0.825 $X2=0
+ $Y2=0
cc_654 N_A_1574_141#_c_897_n N_VGND_c_1277_n 0.0046526f $X=10.065 $Y=0.825 $X2=0
+ $Y2=0
cc_655 N_A_1574_141#_c_894_n N_VGND_c_1278_n 0.00966152f $X=9.705 $Y=0.825 $X2=0
+ $Y2=0
cc_656 N_A_1574_141#_c_895_n N_VGND_c_1278_n 6.16811e-19 $X=9.99 $Y=0.9 $X2=0
+ $Y2=0
cc_657 N_A_1574_141#_c_897_n N_VGND_c_1278_n 0.00919106f $X=10.065 $Y=0.825
+ $X2=0 $Y2=0
cc_658 N_A_1574_141#_c_904_n N_VGND_c_1278_n 0.0095376f $X=8.14 $Y=0.905 $X2=0
+ $Y2=0
cc_659 N_A_1574_141#_c_904_n N_A_1005_141#_c_1435_n 0.0209787f $X=8.14 $Y=0.905
+ $X2=0 $Y2=0
cc_660 COUT N_VPWR_c_1014_n 0.0685263f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_661 COUT N_VPWR_c_1013_n 0.0117582f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_662 COUT N_VPWR_c_1028_n 0.0123222f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_663 COUT N_VGND_c_1263_n 0.0163608f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_664 COUT N_VGND_c_1274_n 0.0154682f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_665 COUT N_VGND_c_1278_n 0.0152006f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_666 N_VPWR_c_1013_n N_A_245_409#_M1011_s 0.00379821f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_1014_n N_A_245_409#_c_1125_n 0.0673848f $X=0.81 $Y=2.06 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_1015_n N_A_245_409#_c_1125_n 0.0540304f $X=1.9 $Y=2.41 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_1019_n N_A_245_409#_c_1125_n 0.0220321f $X=1.735 $Y=3.33 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_1013_n N_A_245_409#_c_1125_n 0.0125808f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_671 N_VPWR_M1029_d N_A_245_409#_c_1126_n 0.00180746f $X=1.76 $Y=2.045 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_1015_n N_A_245_409#_c_1126_n 0.0163515f $X=1.9 $Y=2.41 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_1014_n N_A_245_409#_c_1127_n 0.0121616f $X=0.81 $Y=2.06 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_1015_n N_A_245_409#_c_1130_n 0.00136426f $X=1.9 $Y=2.41 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_1013_n N_A_458_409#_M1027_d 0.00566776f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_1015_n N_A_458_409#_c_1168_n 0.0296179f $X=1.9 $Y=2.41 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_1016_n N_A_458_409#_c_1169_n 0.00907331f $X=4.855 $Y=2.815 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_1021_n N_A_458_409#_c_1169_n 0.101755f $X=4.69 $Y=3.33 $X2=0
+ $Y2=0
cc_679 N_VPWR_c_1013_n N_A_458_409#_c_1169_n 0.0651465f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_680 N_VPWR_c_1015_n N_A_458_409#_c_1170_n 0.0119061f $X=1.9 $Y=2.41 $X2=0
+ $Y2=0
cc_681 N_VPWR_c_1021_n N_A_458_409#_c_1170_n 0.0220111f $X=4.69 $Y=3.33 $X2=0
+ $Y2=0
cc_682 N_VPWR_c_1013_n N_A_458_409#_c_1170_n 0.0126218f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_683 N_VPWR_c_1016_n N_A_458_409#_c_1174_n 0.0190578f $X=4.855 $Y=2.815 $X2=0
+ $Y2=0
cc_684 N_VPWR_c_1013_n N_A_1049_419#_M1000_d 0.0022543f $X=10.32 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_685 N_VPWR_c_1013_n N_A_1049_419#_M1003_d 0.0022543f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_686 N_VPWR_c_1016_n N_A_1049_419#_c_1209_n 0.0250055f $X=4.855 $Y=2.815 $X2=0
+ $Y2=0
cc_687 N_VPWR_c_1017_n N_A_1049_419#_c_1209_n 0.0131781f $X=5.915 $Y=2.95 $X2=0
+ $Y2=0
cc_688 N_VPWR_c_1025_n N_A_1049_419#_c_1209_n 0.0176422f $X=5.75 $Y=3.33 $X2=0
+ $Y2=0
cc_689 N_VPWR_c_1013_n N_A_1049_419#_c_1209_n 0.0123981f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_690 N_VPWR_M1028_d N_A_1049_419#_c_1205_n 0.0477083f $X=5.775 $Y=2.095 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_1017_n N_A_1049_419#_c_1205_n 0.019543f $X=5.915 $Y=2.95 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_1023_n N_A_1049_419#_c_1205_n 0.0238172f $X=9.665 $Y=3.33 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_1025_n N_A_1049_419#_c_1205_n 0.00317549f $X=5.75 $Y=3.33 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_1013_n N_A_1049_419#_c_1205_n 0.0457621f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_1016_n N_A_1049_419#_c_1211_n 0.0119061f $X=4.855 $Y=2.815 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_1023_n N_A_1049_419#_c_1206_n 0.0176422f $X=9.665 $Y=3.33 $X2=0
+ $Y2=0
cc_697 N_VPWR_c_1013_n N_A_1049_419#_c_1206_n 0.0123981f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_698 N_VPWR_c_1013_n A_1720_419# 0.00282558f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_699 N_VPWR_c_1013_n A_1818_419# 0.00317813f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_700 N_VPWR_c_1013_n N_SUM_M1001_d 0.0023218f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_701 N_VPWR_c_1018_n N_SUM_c_1242_n 0.0642065f $X=9.75 $Y=2.24 $X2=0 $Y2=0
cc_702 N_VPWR_c_1026_n N_SUM_c_1242_n 0.0214436f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_703 N_VPWR_c_1013_n N_SUM_c_1242_n 0.0134754f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_704 N_A_245_409#_c_1128_n N_A_458_409#_M1021_d 0.00561832f $X=2.825 $Y=2.18
+ $X2=-0.19 $Y2=1.655
cc_705 N_A_245_409#_c_1130_n N_A_458_409#_M1021_d 0.00318829f $X=2.33 $Y=1.98
+ $X2=-0.19 $Y2=1.655
cc_706 N_A_245_409#_c_1128_n N_A_458_409#_c_1168_n 0.0139082f $X=2.825 $Y=2.18
+ $X2=0 $Y2=0
cc_707 N_A_245_409#_c_1129_n N_A_458_409#_c_1168_n 0.0178286f $X=2.99 $Y=2.405
+ $X2=0 $Y2=0
cc_708 N_A_245_409#_c_1130_n N_A_458_409#_c_1168_n 0.00733762f $X=2.33 $Y=1.98
+ $X2=0 $Y2=0
cc_709 N_A_245_409#_M1011_s N_A_458_409#_c_1169_n 0.0156046f $X=2.845 $Y=2.095
+ $X2=0 $Y2=0
cc_710 N_A_245_409#_c_1128_n N_A_458_409#_c_1169_n 0.00689394f $X=2.825 $Y=2.18
+ $X2=0 $Y2=0
cc_711 N_A_245_409#_c_1129_n N_A_458_409#_c_1169_n 0.0179393f $X=2.99 $Y=2.405
+ $X2=0 $Y2=0
cc_712 SUM N_VGND_c_1270_n 0.00777878f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_713 SUM N_VGND_c_1277_n 0.018672f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_714 SUM N_VGND_c_1278_n 0.0132289f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_715 N_VGND_c_1263_n N_A_355_141#_c_1391_n 0.0403367f $X=1.29 $Y=0.58 $X2=0
+ $Y2=0
cc_716 N_VGND_c_1265_n N_A_355_141#_c_1391_n 0.0260497f $X=2.265 $Y=1.28 $X2=0
+ $Y2=0
cc_717 N_VGND_c_1267_n N_A_355_141#_c_1391_n 0.0125869f $X=2.43 $Y=0.915 $X2=0
+ $Y2=0
cc_718 N_VGND_c_1267_n N_A_355_141#_c_1392_n 0.0234001f $X=2.43 $Y=0.915 $X2=0
+ $Y2=0
cc_719 N_VGND_c_1275_n N_A_355_141#_c_1392_n 0.0826331f $X=4.49 $Y=0 $X2=0 $Y2=0
cc_720 N_VGND_c_1278_n N_A_355_141#_c_1392_n 0.0580629f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_721 N_VGND_c_1263_n N_A_355_141#_c_1393_n 0.014265f $X=1.29 $Y=0.58 $X2=0
+ $Y2=0
cc_722 N_VGND_c_1275_n N_A_355_141#_c_1393_n 0.0167482f $X=4.49 $Y=0 $X2=0 $Y2=0
cc_723 N_VGND_c_1278_n N_A_355_141#_c_1393_n 0.0110904f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_724 N_VGND_c_1268_n N_A_355_141#_c_1394_n 0.0204369f $X=4.655 $Y=0.485 $X2=0
+ $Y2=0
cc_725 N_VGND_c_1275_n N_A_355_141#_c_1394_n 0.0157794f $X=4.49 $Y=0 $X2=0 $Y2=0
cc_726 N_VGND_c_1278_n N_A_355_141#_c_1394_n 0.0107479f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_727 N_VGND_M1004_d N_A_1005_141#_c_1431_n 0.00977412f $X=5.615 $Y=0.705 $X2=0
+ $Y2=0
cc_728 N_VGND_c_1269_n N_A_1005_141#_c_1431_n 0.0209601f $X=5.755 $Y=0.85 $X2=0
+ $Y2=0
cc_729 N_VGND_M1004_d N_A_1005_141#_c_1439_n 0.0278972f $X=5.615 $Y=0.705 $X2=0
+ $Y2=0
cc_730 N_VGND_c_1278_n N_A_1005_141#_c_1439_n 0.00929174f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_731 N_VGND_c_1268_n N_A_1005_141#_c_1433_n 0.0204369f $X=4.655 $Y=0.485 $X2=0
+ $Y2=0
cc_732 N_VGND_c_1269_n N_A_1005_141#_c_1433_n 0.0382104f $X=5.755 $Y=0.85 $X2=0
+ $Y2=0
cc_733 N_VGND_c_1272_n N_A_1005_141#_c_1433_n 0.0162125f $X=5.59 $Y=0 $X2=0
+ $Y2=0
cc_734 N_VGND_c_1278_n N_A_1005_141#_c_1433_n 0.0108853f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_735 N_VGND_M1004_d N_A_1005_141#_c_1434_n 0.0123612f $X=5.615 $Y=0.705 $X2=0
+ $Y2=0
cc_736 N_VGND_c_1269_n N_A_1005_141#_c_1434_n 0.00622561f $X=5.755 $Y=0.85 $X2=0
+ $Y2=0
cc_737 N_VGND_c_1278_n N_A_1005_141#_c_1434_n 0.00564953f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_738 N_VGND_c_1276_n N_A_1005_141#_c_1435_n 0.00558302f $X=9.27 $Y=0 $X2=0
+ $Y2=0
cc_739 N_VGND_c_1278_n N_A_1005_141#_c_1435_n 0.00792972f $X=10.32 $Y=0 $X2=0
+ $Y2=0
