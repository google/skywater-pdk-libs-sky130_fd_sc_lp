* File: sky130_fd_sc_lp__a311oi_m.pxi.spice
* Created: Wed Sep  2 09:26:05 2020
* 
x_PM_SKY130_FD_SC_LP__A311OI_M%A3 N_A3_c_77_n N_A3_c_84_n N_A3_c_85_n
+ N_A3_M1006_g N_A3_c_78_n N_A3_M1001_g N_A3_c_79_n N_A3_c_80_n A3 A3 A3 A3 A3
+ A3 A3 N_A3_c_82_n PM_SKY130_FD_SC_LP__A311OI_M%A3
x_PM_SKY130_FD_SC_LP__A311OI_M%A2 N_A2_c_124_n N_A2_M1008_g N_A2_M1004_g
+ N_A2_c_128_n N_A2_c_129_n N_A2_c_130_n A2 A2 A2 A2 A2 N_A2_c_127_n
+ PM_SKY130_FD_SC_LP__A311OI_M%A2
x_PM_SKY130_FD_SC_LP__A311OI_M%A1 N_A1_M1009_g N_A1_M1000_g N_A1_c_183_n
+ N_A1_c_184_n A1 A1 A1 N_A1_c_181_n PM_SKY130_FD_SC_LP__A311OI_M%A1
x_PM_SKY130_FD_SC_LP__A311OI_M%B1 N_B1_M1002_g N_B1_M1007_g N_B1_c_226_n
+ N_B1_c_227_n N_B1_c_228_n N_B1_c_229_n N_B1_c_234_n B1 B1 B1 N_B1_c_231_n
+ PM_SKY130_FD_SC_LP__A311OI_M%B1
x_PM_SKY130_FD_SC_LP__A311OI_M%C1 N_C1_c_277_n N_C1_M1005_g N_C1_M1003_g
+ N_C1_c_278_n N_C1_c_279_n N_C1_c_284_n N_C1_c_285_n N_C1_c_280_n C1 C1 C1 C1
+ N_C1_c_282_n PM_SKY130_FD_SC_LP__A311OI_M%C1
x_PM_SKY130_FD_SC_LP__A311OI_M%VPWR N_VPWR_M1006_s N_VPWR_M1004_d N_VPWR_c_322_n
+ N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n VPWR
+ N_VPWR_c_327_n N_VPWR_c_321_n PM_SKY130_FD_SC_LP__A311OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A311OI_M%A_191_535# N_A_191_535#_M1006_d
+ N_A_191_535#_M1000_d N_A_191_535#_c_363_n N_A_191_535#_c_364_n
+ N_A_191_535#_c_365_n N_A_191_535#_c_366_n
+ PM_SKY130_FD_SC_LP__A311OI_M%A_191_535#
x_PM_SKY130_FD_SC_LP__A311OI_M%Y N_Y_M1009_d N_Y_M1005_d N_Y_M1003_d N_Y_c_407_n
+ N_Y_c_400_n Y Y Y Y Y Y N_Y_c_405_n Y N_Y_c_403_n
+ PM_SKY130_FD_SC_LP__A311OI_M%Y
x_PM_SKY130_FD_SC_LP__A311OI_M%VGND N_VGND_M1001_s N_VGND_M1002_d N_VGND_c_442_n
+ N_VGND_c_443_n N_VGND_c_444_n VGND N_VGND_c_445_n N_VGND_c_446_n
+ N_VGND_c_447_n N_VGND_c_448_n PM_SKY130_FD_SC_LP__A311OI_M%VGND
cc_1 VNB N_A3_c_77_n 0.0159782f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.085
cc_2 VNB N_A3_c_78_n 0.0187829f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.785
cc_3 VNB N_A3_c_79_n 0.0428155f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.86
cc_4 VNB N_A3_c_80_n 0.0199744f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.455
cc_5 VNB A3 0.0100176f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_6 VNB N_A3_c_82_n 0.0359062f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.95
cc_7 VNB N_A2_c_124_n 0.020588f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.16
cc_8 VNB N_A2_M1008_g 0.0317239f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.235
cc_9 VNB A2 0.00351306f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.86
cc_10 VNB N_A2_c_127_n 0.0261966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_M1009_g 0.0545982f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.16
cc_12 VNB A1 0.0042485f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.935
cc_13 VNB N_A1_c_181_n 0.0150669f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_14 VNB N_B1_c_226_n 0.015312f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.465
cc_15 VNB N_B1_c_227_n 0.0139026f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.465
cc_16 VNB N_B1_c_228_n 0.0180326f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.935
cc_17 VNB N_B1_c_229_n 0.0213433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB B1 0.00125055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_231_n 0.0184324f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_20 VNB N_C1_c_277_n 0.019508f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.455
cc_21 VNB N_C1_c_278_n 0.0256725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C1_c_279_n 0.0122344f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.785
cc_23 VNB N_C1_c_280_n 0.0393578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB C1 0.00530689f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.29
cc_25 VNB N_C1_c_282_n 0.00796429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_321_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_400_n 0.00675004f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.86
cc_28 VNB Y 0.0313905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB Y 0.0383179f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.95
cc_30 VNB N_Y_c_403_n 0.00850378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_442_n 0.0107731f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.885
cc_32 VNB N_VGND_c_443_n 0.00572882f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.785
cc_33 VNB N_VGND_c_444_n 0.00100404f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.935
cc_34 VNB N_VGND_c_445_n 0.0502858f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.29
cc_35 VNB N_VGND_c_446_n 0.0251131f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_36 VNB N_VGND_c_447_n 0.222538f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_37 VNB N_VGND_c_448_n 0.00460801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A3_c_77_n 0.0354989f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.085
cc_39 VPB N_A3_c_84_n 0.0273841f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.16
cc_40 VPB N_A3_c_85_n 0.0168378f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.16
cc_41 VPB N_A3_M1006_g 0.0370433f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=2.885
cc_42 VPB A3 0.0256009f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_43 VPB N_A2_c_128_n 0.0181263f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.86
cc_44 VPB N_A2_c_129_n 0.0297628f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_45 VPB N_A2_c_130_n 0.0293087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB A2 0.00341539f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.86
cc_47 VPB N_A2_c_127_n 0.00179459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A1_M1000_g 0.0344578f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=2.885
cc_49 VPB N_A1_c_183_n 0.0232625f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.465
cc_50 VPB N_A1_c_184_n 0.0164978f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.86
cc_51 VPB A1 7.47878e-19 $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_52 VPB N_A1_c_181_n 0.00307112f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_53 VPB N_B1_M1007_g 0.0478781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B1_c_229_n 0.00402608f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B1_c_234_n 0.0185986f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.86
cc_56 VPB B1 0.00656907f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_C1_M1003_g 0.0370895f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=2.885
cc_58 VPB N_C1_c_284_n 0.0256668f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_59 VPB N_C1_c_285_n 0.0304034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB C1 0.00817188f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.29
cc_61 VPB N_C1_c_282_n 0.00754249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_322_n 0.0107725f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=2.885
cc_63 VPB N_VPWR_c_323_n 0.00485511f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.785
cc_64 VPB N_VPWR_c_324_n 0.00482866f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_65 VPB N_VPWR_c_325_n 0.0299798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_326_n 0.00362661f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.29
cc_67 VPB N_VPWR_c_327_n 0.0502744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_321_n 0.0509835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_191_535#_c_363_n 6.7104e-19 $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.785
cc_70 VPB N_A_191_535#_c_364_n 0.00936666f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.465
cc_71 VPB N_A_191_535#_c_365_n 0.00320773f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.86
cc_72 VPB N_A_191_535#_c_366_n 0.00899229f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_73 VPB Y 0.00944387f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_74 VPB N_Y_c_405_n 0.0165143f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.95
cc_75 VPB Y 0.0484965f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.95
cc_76 N_A3_c_79_n N_A2_c_124_n 7.36453e-19 $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_77 A3 N_A2_c_124_n 0.00536736f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_78 N_A3_c_82_n N_A2_c_124_n 0.00963178f $X=0.61 $Y=0.95 $X2=0 $Y2=0
cc_79 N_A3_c_78_n N_A2_M1008_g 0.0510476f $X=0.92 $Y=0.785 $X2=0 $Y2=0
cc_80 A3 N_A2_M1008_g 7.53733e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_81 N_A3_c_82_n N_A2_M1008_g 0.00519142f $X=0.61 $Y=0.95 $X2=0 $Y2=0
cc_82 N_A3_c_77_n N_A2_c_129_n 0.00359324f $X=0.52 $Y=2.085 $X2=0 $Y2=0
cc_83 N_A3_c_84_n N_A2_c_129_n 0.0149105f $X=0.805 $Y=2.16 $X2=0 $Y2=0
cc_84 A3 N_A2_c_129_n 0.00141709f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A3_M1006_g N_A2_c_130_n 0.0302262f $X=0.88 $Y=2.885 $X2=0 $Y2=0
cc_86 N_A3_c_77_n A2 9.86688e-19 $X=0.52 $Y=2.085 $X2=0 $Y2=0
cc_87 N_A3_c_84_n A2 2.69421e-19 $X=0.805 $Y=2.16 $X2=0 $Y2=0
cc_88 N_A3_c_78_n A2 0.0035736f $X=0.92 $Y=0.785 $X2=0 $Y2=0
cc_89 A3 A2 0.0878193f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A3_c_82_n A2 0.00116697f $X=0.61 $Y=0.95 $X2=0 $Y2=0
cc_91 N_A3_c_77_n N_A2_c_127_n 0.0104801f $X=0.52 $Y=2.085 $X2=0 $Y2=0
cc_92 N_A3_c_80_n N_A2_c_127_n 0.00876553f $X=0.61 $Y=1.455 $X2=0 $Y2=0
cc_93 A3 N_VPWR_M1006_s 0.0107975f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_94 N_A3_M1006_g N_VPWR_c_323_n 0.00722131f $X=0.88 $Y=2.885 $X2=0 $Y2=0
cc_95 A3 N_VPWR_c_323_n 0.00546724f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_96 N_A3_M1006_g N_VPWR_c_325_n 0.00585385f $X=0.88 $Y=2.885 $X2=0 $Y2=0
cc_97 A3 N_VPWR_c_325_n 0.0072891f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_98 N_A3_M1006_g N_VPWR_c_321_n 0.0124078f $X=0.88 $Y=2.885 $X2=0 $Y2=0
cc_99 A3 N_VPWR_c_321_n 0.00949689f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A3_M1006_g N_A_191_535#_c_363_n 3.77206e-19 $X=0.88 $Y=2.885 $X2=0
+ $Y2=0
cc_101 A3 N_A_191_535#_c_363_n 0.00363011f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_102 N_A3_M1006_g N_A_191_535#_c_365_n 0.00137775f $X=0.88 $Y=2.885 $X2=0
+ $Y2=0
cc_103 A3 N_A_191_535#_c_365_n 0.0139875f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_104 A3 N_VGND_M1001_s 0.0112865f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_105 N_A3_c_78_n N_VGND_c_443_n 0.00747537f $X=0.92 $Y=0.785 $X2=0 $Y2=0
cc_106 A3 N_VGND_c_443_n 0.00692518f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_107 N_A3_c_78_n N_VGND_c_445_n 0.00565115f $X=0.92 $Y=0.785 $X2=0 $Y2=0
cc_108 A3 N_VGND_c_445_n 0.00782722f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_109 N_A3_c_78_n N_VGND_c_447_n 0.0118165f $X=0.92 $Y=0.785 $X2=0 $Y2=0
cc_110 N_A3_c_79_n N_VGND_c_447_n 0.00300234f $X=0.92 $Y=0.86 $X2=0 $Y2=0
cc_111 A3 N_VGND_c_447_n 0.00949689f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A2_M1008_g N_A1_M1009_g 0.0712765f $X=1.28 $Y=0.465 $X2=0 $Y2=0
cc_113 A2 N_A1_M1009_g 0.00419539f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_114 N_A2_c_127_n N_A1_M1009_g 0.0112546f $X=1.15 $Y=1.34 $X2=0 $Y2=0
cc_115 N_A2_c_129_n N_A1_M1000_g 0.00867821f $X=1.275 $Y=2.415 $X2=0 $Y2=0
cc_116 N_A2_c_130_n N_A1_M1000_g 0.0224311f $X=1.275 $Y=2.565 $X2=0 $Y2=0
cc_117 N_A2_c_128_n N_A1_c_183_n 0.0135757f $X=1.15 $Y=1.845 $X2=0 $Y2=0
cc_118 N_A2_c_129_n N_A1_c_184_n 0.0135757f $X=1.275 $Y=2.415 $X2=0 $Y2=0
cc_119 N_A2_c_124_n A1 3.04263e-19 $X=1.28 $Y=1.145 $X2=0 $Y2=0
cc_120 A2 A1 0.0389504f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A2_c_127_n A1 0.0031133f $X=1.15 $Y=1.34 $X2=0 $Y2=0
cc_122 A2 N_A1_c_181_n 0.00204304f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A2_c_127_n N_A1_c_181_n 0.0135757f $X=1.15 $Y=1.34 $X2=0 $Y2=0
cc_124 N_A2_c_130_n N_VPWR_c_324_n 0.00285763f $X=1.275 $Y=2.565 $X2=0 $Y2=0
cc_125 N_A2_c_130_n N_VPWR_c_325_n 0.00456613f $X=1.275 $Y=2.565 $X2=0 $Y2=0
cc_126 N_A2_c_130_n N_VPWR_c_321_n 0.00599853f $X=1.275 $Y=2.565 $X2=0 $Y2=0
cc_127 N_A2_c_130_n N_A_191_535#_c_363_n 6.39777e-19 $X=1.275 $Y=2.565 $X2=0
+ $Y2=0
cc_128 N_A2_c_130_n N_A_191_535#_c_364_n 0.015054f $X=1.275 $Y=2.565 $X2=0 $Y2=0
cc_129 A2 N_A_191_535#_c_364_n 0.00368754f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_130 N_A2_c_128_n N_A_191_535#_c_365_n 0.00264496f $X=1.15 $Y=1.845 $X2=0
+ $Y2=0
cc_131 N_A2_c_130_n N_A_191_535#_c_365_n 0.00248499f $X=1.275 $Y=2.565 $X2=0
+ $Y2=0
cc_132 A2 N_A_191_535#_c_365_n 0.00733121f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_133 N_A2_c_130_n N_A_191_535#_c_366_n 5.18854e-19 $X=1.275 $Y=2.565 $X2=0
+ $Y2=0
cc_134 A2 N_Y_c_407_n 0.00349937f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_135 A2 N_Y_c_400_n 0.00656335f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_136 N_A2_M1008_g N_VGND_c_445_n 0.00469388f $X=1.28 $Y=0.465 $X2=0 $Y2=0
cc_137 A2 N_VGND_c_445_n 0.00541982f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_138 N_A2_M1008_g N_VGND_c_447_n 0.00766989f $X=1.28 $Y=0.465 $X2=0 $Y2=0
cc_139 A2 N_VGND_c_447_n 0.00705042f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_140 A2 A_199_51# 0.00318989f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_141 N_A1_M1000_g N_B1_M1007_g 0.0328691f $X=1.74 $Y=2.885 $X2=0 $Y2=0
cc_142 N_A1_c_183_n N_B1_M1007_g 0.0174728f $X=1.69 $Y=2.04 $X2=0 $Y2=0
cc_143 A1 N_B1_M1007_g 7.32753e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A1_M1009_g N_B1_c_226_n 0.0214587f $X=1.64 $Y=0.465 $X2=0 $Y2=0
cc_145 N_A1_M1009_g N_B1_c_228_n 0.0219056f $X=1.64 $Y=0.465 $X2=0 $Y2=0
cc_146 A1 N_B1_c_229_n 0.00107341f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A1_c_181_n N_B1_c_229_n 0.0106544f $X=1.69 $Y=1.7 $X2=0 $Y2=0
cc_148 N_A1_c_183_n N_B1_c_234_n 0.0106544f $X=1.69 $Y=2.04 $X2=0 $Y2=0
cc_149 N_A1_M1009_g B1 3.79887e-19 $X=1.64 $Y=0.465 $X2=0 $Y2=0
cc_150 N_A1_c_183_n B1 0.00161969f $X=1.69 $Y=2.04 $X2=0 $Y2=0
cc_151 A1 B1 0.0425437f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A1_c_181_n B1 0.00125338f $X=1.69 $Y=1.7 $X2=0 $Y2=0
cc_153 A1 N_B1_c_231_n 0.00222059f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A1_M1000_g N_VPWR_c_324_n 0.00274937f $X=1.74 $Y=2.885 $X2=0 $Y2=0
cc_155 N_A1_M1000_g N_VPWR_c_327_n 0.00428423f $X=1.74 $Y=2.885 $X2=0 $Y2=0
cc_156 N_A1_M1000_g N_VPWR_c_321_n 0.00593521f $X=1.74 $Y=2.885 $X2=0 $Y2=0
cc_157 N_A1_M1000_g N_A_191_535#_c_364_n 0.010073f $X=1.74 $Y=2.885 $X2=0 $Y2=0
cc_158 N_A1_c_184_n N_A_191_535#_c_364_n 0.00313343f $X=1.69 $Y=2.205 $X2=0
+ $Y2=0
cc_159 A1 N_A_191_535#_c_364_n 0.0102146f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A1_M1000_g N_A_191_535#_c_366_n 0.00954051f $X=1.74 $Y=2.885 $X2=0
+ $Y2=0
cc_161 N_A1_c_184_n N_A_191_535#_c_366_n 0.00167937f $X=1.69 $Y=2.205 $X2=0
+ $Y2=0
cc_162 N_A1_M1009_g N_Y_c_400_n 0.00239046f $X=1.64 $Y=0.465 $X2=0 $Y2=0
cc_163 A1 N_Y_c_400_n 0.00131454f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A1_c_181_n N_Y_c_400_n 0.00230534f $X=1.69 $Y=1.7 $X2=0 $Y2=0
cc_165 N_A1_M1009_g N_VGND_c_444_n 0.00148754f $X=1.64 $Y=0.465 $X2=0 $Y2=0
cc_166 N_A1_M1009_g N_VGND_c_445_n 0.00565115f $X=1.64 $Y=0.465 $X2=0 $Y2=0
cc_167 N_A1_M1009_g N_VGND_c_447_n 0.0106402f $X=1.64 $Y=0.465 $X2=0 $Y2=0
cc_168 N_B1_c_226_n N_C1_c_277_n 0.0140864f $X=2.105 $Y=0.785 $X2=-0.19
+ $Y2=-0.245
cc_169 N_B1_c_227_n N_C1_c_279_n 0.0105225f $X=2.105 $Y=0.935 $X2=0 $Y2=0
cc_170 N_B1_M1007_g N_C1_c_284_n 0.00773724f $X=2.17 $Y=2.885 $X2=0 $Y2=0
cc_171 N_B1_c_234_n N_C1_c_284_n 0.0087078f $X=2.23 $Y=1.88 $X2=0 $Y2=0
cc_172 B1 N_C1_c_284_n 8.0658e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_B1_M1007_g N_C1_c_285_n 0.0687299f $X=2.17 $Y=2.885 $X2=0 $Y2=0
cc_174 N_B1_c_228_n N_C1_c_280_n 0.00724161f $X=2.23 $Y=1.21 $X2=0 $Y2=0
cc_175 B1 N_C1_c_280_n 3.30393e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_176 N_B1_c_231_n N_C1_c_280_n 0.010432f $X=2.23 $Y=1.375 $X2=0 $Y2=0
cc_177 N_B1_M1007_g C1 0.00267649f $X=2.17 $Y=2.885 $X2=0 $Y2=0
cc_178 B1 C1 0.0549401f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_179 N_B1_c_231_n C1 0.0053354f $X=2.23 $Y=1.375 $X2=0 $Y2=0
cc_180 N_B1_c_229_n N_C1_c_282_n 0.0087078f $X=2.23 $Y=1.715 $X2=0 $Y2=0
cc_181 B1 N_C1_c_282_n 2.86229e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_B1_M1007_g N_VPWR_c_327_n 0.00553654f $X=2.17 $Y=2.885 $X2=0 $Y2=0
cc_183 N_B1_M1007_g N_VPWR_c_321_n 0.00997093f $X=2.17 $Y=2.885 $X2=0 $Y2=0
cc_184 N_B1_M1007_g N_A_191_535#_c_366_n 0.011389f $X=2.17 $Y=2.885 $X2=0 $Y2=0
cc_185 N_B1_c_234_n N_A_191_535#_c_366_n 4.17533e-19 $X=2.23 $Y=1.88 $X2=0 $Y2=0
cc_186 B1 N_A_191_535#_c_366_n 0.00222091f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B1_c_226_n N_Y_c_407_n 2.03427e-19 $X=2.105 $Y=0.785 $X2=0 $Y2=0
cc_188 N_B1_c_226_n N_Y_c_403_n 0.00680482f $X=2.105 $Y=0.785 $X2=0 $Y2=0
cc_189 N_B1_c_227_n N_Y_c_403_n 0.00979311f $X=2.105 $Y=0.935 $X2=0 $Y2=0
cc_190 B1 N_Y_c_403_n 0.0103973f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_191 N_B1_c_231_n N_Y_c_403_n 0.00332531f $X=2.23 $Y=1.375 $X2=0 $Y2=0
cc_192 N_B1_c_226_n N_VGND_c_444_n 0.00851777f $X=2.105 $Y=0.785 $X2=0 $Y2=0
cc_193 N_B1_c_227_n N_VGND_c_444_n 2.77104e-19 $X=2.105 $Y=0.935 $X2=0 $Y2=0
cc_194 N_B1_c_226_n N_VGND_c_445_n 0.00345529f $X=2.105 $Y=0.785 $X2=0 $Y2=0
cc_195 N_B1_c_226_n N_VGND_c_447_n 0.00421603f $X=2.105 $Y=0.785 $X2=0 $Y2=0
cc_196 N_C1_M1003_g N_VPWR_c_327_n 0.00585385f $X=2.53 $Y=2.885 $X2=0 $Y2=0
cc_197 N_C1_M1003_g N_VPWR_c_321_n 0.010759f $X=2.53 $Y=2.885 $X2=0 $Y2=0
cc_198 C1 N_VPWR_c_321_n 0.00353887f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_199 N_C1_M1003_g N_A_191_535#_c_366_n 0.00171778f $X=2.53 $Y=2.885 $X2=0
+ $Y2=0
cc_200 C1 N_A_191_535#_c_366_n 0.00121927f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_201 N_C1_c_277_n Y 4.26254e-19 $X=2.5 $Y=0.785 $X2=0 $Y2=0
cc_202 N_C1_c_278_n Y 0.01731f $X=2.785 $Y=0.86 $X2=0 $Y2=0
cc_203 N_C1_c_285_n Y 0.00374273f $X=2.695 $Y=2.27 $X2=0 $Y2=0
cc_204 C1 Y 0.0172109f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_205 N_C1_M1003_g Y 0.00556098f $X=2.53 $Y=2.885 $X2=0 $Y2=0
cc_206 N_C1_c_278_n Y 0.0383549f $X=2.785 $Y=0.86 $X2=0 $Y2=0
cc_207 C1 Y 0.09227f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_208 N_C1_c_277_n N_Y_c_403_n 0.00817602f $X=2.5 $Y=0.785 $X2=0 $Y2=0
cc_209 N_C1_c_278_n N_Y_c_403_n 0.00184154f $X=2.785 $Y=0.86 $X2=0 $Y2=0
cc_210 N_C1_c_279_n N_Y_c_403_n 0.00674951f $X=2.575 $Y=0.86 $X2=0 $Y2=0
cc_211 C1 N_Y_c_403_n 0.0142921f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_212 N_C1_c_277_n N_VGND_c_444_n 0.0116358f $X=2.5 $Y=0.785 $X2=0 $Y2=0
cc_213 N_C1_c_277_n N_VGND_c_446_n 0.00345529f $X=2.5 $Y=0.785 $X2=0 $Y2=0
cc_214 N_C1_c_277_n N_VGND_c_447_n 0.00539236f $X=2.5 $Y=0.785 $X2=0 $Y2=0
cc_215 N_VPWR_c_321_n N_A_191_535#_M1006_d 0.00374715f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_216 N_VPWR_c_321_n N_A_191_535#_M1000_d 0.0024615f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_325_n N_A_191_535#_c_363_n 0.00756903f $X=1.42 $Y=3.33 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_321_n N_A_191_535#_c_363_n 0.00753735f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_324_n N_A_191_535#_c_364_n 0.0132188f $X=1.525 $Y=2.97 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_325_n N_A_191_535#_c_364_n 0.00318349f $X=1.42 $Y=3.33 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_327_n N_A_191_535#_c_364_n 0.00260523f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_321_n N_A_191_535#_c_364_n 0.0101207f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_327_n N_A_191_535#_c_366_n 0.00944217f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_321_n N_A_191_535#_c_366_n 0.0112873f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_321_n A_449_535# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_226 N_VPWR_c_321_n N_Y_M1003_d 0.00251773f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_227 N_VPWR_c_327_n Y 0.0172678f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_228 N_VPWR_c_321_n Y 0.0142354f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_c_327_n N_Y_c_405_n 0.00819846f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_230 N_VPWR_c_321_n N_Y_c_405_n 0.00634055f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_231 N_A_191_535#_c_366_n Y 0.00385365f $X=1.955 $Y=2.54 $X2=0 $Y2=0
cc_232 N_Y_c_403_n N_VGND_c_444_n 0.0193682f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_233 N_Y_c_407_n N_VGND_c_445_n 0.00711705f $X=1.855 $Y=0.53 $X2=0 $Y2=0
cc_234 N_Y_c_403_n N_VGND_c_445_n 0.00271048f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_235 Y N_VGND_c_446_n 0.0232709f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_236 N_Y_c_403_n N_VGND_c_446_n 0.00271048f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_237 N_Y_c_407_n N_VGND_c_447_n 0.00679726f $X=1.855 $Y=0.53 $X2=0 $Y2=0
cc_238 Y N_VGND_c_447_n 0.02078f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_239 N_Y_c_403_n N_VGND_c_447_n 0.0100561f $X=2.63 $Y=0.61 $X2=0 $Y2=0
