* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_367_491# a_27_75# a_453_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VGND a_1812_379# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_1953_496# a_2002_42# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_1024_367# a_840_119# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR RESET_B a_367_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VGND CLK a_840_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1812_379# a_1024_367# a_1953_496# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_453_491# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1374_362# a_840_119# a_1812_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_300_75# D a_367_491# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1246_463# a_1024_367# a_1430_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_840_119# a_1024_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND a_840_119# a_1024_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_1812_379# a_2352_327# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1332_463# a_1374_362# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND a_1246_463# a_1374_362# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 a_1374_362# a_1024_367# a_1812_379# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 a_217_75# a_27_75# a_300_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_840_119# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR RESET_B a_2002_42# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_1502_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 Q a_2352_327# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 VPWR RESET_B a_1246_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_27_75# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_840_119# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_27_75# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_367_491# SCE a_488_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_367_491# a_1024_367# a_1246_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_1430_119# a_1374_362# a_1502_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_217_75# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_2002_42# a_1812_379# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 VPWR a_1812_379# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_2138_68# a_1812_379# a_2002_42# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VPWR SCE a_295_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X34 a_295_491# D a_367_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 Q a_2352_327# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 a_1246_463# a_840_119# a_1332_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 VPWR a_1812_379# a_2352_327# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X38 a_1812_379# a_840_119# a_1960_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND RESET_B a_2138_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_488_81# SCD a_217_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 VPWR a_1246_463# a_1374_362# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X42 a_367_491# a_840_119# a_1246_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_1960_68# a_2002_42# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
