* NGSPICE file created from sky130_fd_sc_lp__a211o_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a211o_0 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_80_172# C1 VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=5.208e+11p ps=4.16e+06u
M1001 a_265_60# A2 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1002 a_80_172# A1 a_265_60# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B1 a_80_172# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_487_482# B1 a_224_482# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=3.488e+11p ps=3.65e+06u
M1005 a_80_172# C1 a_487_482# VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1006 a_224_482# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.744e+11p ps=3.73e+06u
M1007 VGND a_80_172# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 VPWR A2 a_224_482# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_80_172# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
.ends

