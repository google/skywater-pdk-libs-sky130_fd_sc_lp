* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_267_47# B1 a_591_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_356_367# A3 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR A1 a_267_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_267_367# A2 a_356_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_591_47# C1 a_80_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_267_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND A1 a_267_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND A3 a_267_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
