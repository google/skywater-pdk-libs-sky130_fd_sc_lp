* NGSPICE file created from sky130_fd_sc_lp__and4bb_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4bb_m A_N B_N C D VGND VNB VPB VPWR X
M1000 VGND A_N a_54_55# VNB nshort w=420000u l=150000u
+  ad=3.003e+11p pd=3.11e+06u as=1.113e+11p ps=1.37e+06u
M1001 a_223_55# B_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1002 VGND D a_595_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1003 VPWR a_223_55# a_332_125# VPB phighvt w=420000u l=150000u
+  ad=4.809e+11p pd=5.65e+06u as=2.352e+11p ps=2.8e+06u
M1004 a_415_125# a_54_55# a_332_125# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1005 X a_332_125# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 a_595_125# C a_487_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1007 VPWR D a_332_125# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_332_125# a_54_55# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_332_125# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1010 VPWR A_N a_54_55# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 a_332_125# C VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_223_55# B_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 a_487_125# a_223_55# a_415_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

