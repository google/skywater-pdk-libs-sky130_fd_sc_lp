* File: sky130_fd_sc_lp__nand3b_4.pex.spice
* Created: Fri Aug 28 10:49:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3B_4%A_N 1 3 4 6 7 8 13
r35 13 15 13.0438 $w=3.88e-07 $l=1.05e-07 $layer=POLY_cond $X=0.685 $Y=1.52
+ $X2=0.79 $Y2=1.52
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.685
+ $Y=1.485 $X2=0.685 $Y2=1.485
r37 11 13 21.1186 $w=3.88e-07 $l=1.7e-07 $layer=POLY_cond $X=0.515 $Y=1.52
+ $X2=0.685 $Y2=1.52
r38 8 14 9.73836 $w=2.03e-07 $l=1.8e-07 $layer=LI1_cond $X=0.702 $Y=1.665
+ $X2=0.702 $Y2=1.485
r39 7 14 10.2794 $w=2.03e-07 $l=1.9e-07 $layer=LI1_cond $X=0.702 $Y=1.295
+ $X2=0.702 $Y2=1.485
r40 4 15 25.1189 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=0.79 $Y=1.72 $X2=0.79
+ $Y2=1.52
r41 4 6 239.393 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.79 $Y=1.72 $X2=0.79
+ $Y2=2.465
r42 1 11 25.1189 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=0.515 $Y=1.32 $X2=0.515
+ $Y2=1.52
r43 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.515 $Y=1.32
+ $X2=0.515 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%A_35_74# 1 2 9 11 13 16 18 20 23 25 27 30
+ 32 34 37 42 45 47 50 56 57 59 61
c124 57 0 6.17957e-20 $X=2.585 $Y=1.4
c125 56 0 1.90858e-19 $X=2.585 $Y=1.4
c126 25 0 5.86634e-20 $X=2.325 $Y=1.185
r127 73 74 32.6558 $w=3.69e-07 $l=2.5e-07 $layer=POLY_cond $X=2.325 $Y=1.375
+ $X2=2.575 $Y2=1.375
r128 72 73 23.5122 $w=3.69e-07 $l=1.8e-07 $layer=POLY_cond $X=2.145 $Y=1.375
+ $X2=2.325 $Y2=1.375
r129 71 72 32.6558 $w=3.69e-07 $l=2.5e-07 $layer=POLY_cond $X=1.895 $Y=1.375
+ $X2=2.145 $Y2=1.375
r130 70 71 23.5122 $w=3.69e-07 $l=1.8e-07 $layer=POLY_cond $X=1.715 $Y=1.375
+ $X2=1.895 $Y2=1.375
r131 67 68 23.5122 $w=3.69e-07 $l=1.8e-07 $layer=POLY_cond $X=1.285 $Y=1.375
+ $X2=1.465 $Y2=1.375
r132 65 67 7.8374 $w=3.69e-07 $l=6e-08 $layer=POLY_cond $X=1.225 $Y=1.375
+ $X2=1.285 $Y2=1.375
r133 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.4 $X2=1.225 $Y2=1.4
r134 61 62 5.39863 $w=6.03e-07 $l=8.5e-08 $layer=LI1_cond $X=0.437 $Y=2.005
+ $X2=0.437 $Y2=1.92
r135 57 74 1.30623 $w=3.69e-07 $l=1e-08 $layer=POLY_cond $X=2.585 $Y=1.375
+ $X2=2.575 $Y2=1.375
r136 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.585
+ $Y=1.4 $X2=2.585 $Y2=1.4
r137 54 70 19.5935 $w=3.69e-07 $l=1.5e-07 $layer=POLY_cond $X=1.565 $Y=1.375
+ $X2=1.715 $Y2=1.375
r138 54 68 13.0623 $w=3.69e-07 $l=1e-07 $layer=POLY_cond $X=1.565 $Y=1.375
+ $X2=1.465 $Y2=1.375
r139 53 56 55.184 $w=2.03e-07 $l=1.02e-06 $layer=LI1_cond $X=1.565 $Y=1.417
+ $X2=2.585 $Y2=1.417
r140 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.565
+ $Y=1.4 $X2=1.565 $Y2=1.4
r141 51 64 4.65982 $w=2.05e-07 $l=1.73e-07 $layer=LI1_cond $X=1.32 $Y=1.417
+ $X2=1.147 $Y2=1.417
r142 51 53 13.255 $w=2.03e-07 $l=2.45e-07 $layer=LI1_cond $X=1.32 $Y=1.417
+ $X2=1.565 $Y2=1.417
r143 50 64 2.74741 $w=3.45e-07 $l=1.02e-07 $layer=LI1_cond $X=1.147 $Y=1.315
+ $X2=1.147 $Y2=1.417
r144 49 50 9.18614 $w=3.43e-07 $l=2.75e-07 $layer=LI1_cond $X=1.147 $Y=1.04
+ $X2=1.147 $Y2=1.315
r145 48 59 2.98021 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.405 $Y=0.955
+ $X2=0.27 $Y2=0.955
r146 47 49 7.89393 $w=1.7e-07 $l=2.10247e-07 $layer=LI1_cond $X=0.975 $Y=0.955
+ $X2=1.147 $Y2=1.04
r147 47 48 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.975 $Y=0.955
+ $X2=0.405 $Y2=0.955
r148 43 61 4.29007 $w=6.03e-07 $l=2.17e-07 $layer=LI1_cond $X=0.437 $Y=2.222
+ $X2=0.437 $Y2=2.005
r149 43 45 13.6017 $w=6.03e-07 $l=6.88e-07 $layer=LI1_cond $X=0.437 $Y=2.222
+ $X2=0.437 $Y2=2.91
r150 42 62 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.27 $Y=1.065
+ $X2=0.27 $Y2=1.92
r151 39 59 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.04
+ $X2=0.27 $Y2=0.955
r152 39 42 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.27 $Y=1.04
+ $X2=0.27 $Y2=1.065
r153 35 59 3.52026 $w=2.65e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.265 $Y=0.87
+ $X2=0.27 $Y2=0.955
r154 35 37 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.265 $Y=0.87
+ $X2=0.265 $Y2=0.525
r155 32 57 22.206 $w=3.69e-07 $l=2.61534e-07 $layer=POLY_cond $X=2.755 $Y=1.185
+ $X2=2.585 $Y2=1.375
r156 32 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.755 $Y=1.185
+ $X2=2.755 $Y2=0.655
r157 28 74 23.9013 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.575 $Y=1.565
+ $X2=2.575 $Y2=1.375
r158 28 30 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.575 $Y=1.565
+ $X2=2.575 $Y2=2.465
r159 25 73 23.9013 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.325 $Y=1.185
+ $X2=2.325 $Y2=1.375
r160 25 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.325 $Y=1.185
+ $X2=2.325 $Y2=0.655
r161 21 72 23.9013 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.145 $Y=1.565
+ $X2=2.145 $Y2=1.375
r162 21 23 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.145 $Y=1.565
+ $X2=2.145 $Y2=2.465
r163 18 71 23.9013 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.895 $Y=1.185
+ $X2=1.895 $Y2=1.375
r164 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.895 $Y=1.185
+ $X2=1.895 $Y2=0.655
r165 14 70 23.9013 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.715 $Y=1.565
+ $X2=1.715 $Y2=1.375
r166 14 16 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.715 $Y=1.565
+ $X2=1.715 $Y2=2.465
r167 11 68 23.9013 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.465 $Y=1.185
+ $X2=1.465 $Y2=1.375
r168 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.465 $Y=1.185
+ $X2=1.465 $Y2=0.655
r169 7 67 23.9013 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.285 $Y=1.565
+ $X2=1.285 $Y2=1.375
r170 7 9 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.285 $Y=1.565
+ $X2=1.285 $Y2=2.465
r171 2 61 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.45
+ $Y=1.835 $X2=0.575 $Y2=2.005
r172 2 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.45
+ $Y=1.835 $X2=0.575 $Y2=2.91
r173 1 42 182 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.37 $X2=0.3 $Y2=1.065
r174 1 37 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.37 $X2=0.3 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 45 48
c87 22 0 2.98258e-20 $X=4.405 $Y=1.725
c88 6 0 1.90858e-19 $X=3.185 $Y=0.655
r89 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.57
+ $Y=1.51 $X2=4.57 $Y2=1.51
r90 45 47 12.7194 $w=3.6e-07 $l=9.5e-08 $layer=POLY_cond $X=4.475 $Y=1.535
+ $X2=4.57 $Y2=1.535
r91 44 45 9.37222 $w=3.6e-07 $l=7e-08 $layer=POLY_cond $X=4.405 $Y=1.535
+ $X2=4.475 $Y2=1.535
r92 43 44 48.2 $w=3.6e-07 $l=3.6e-07 $layer=POLY_cond $X=4.045 $Y=1.535
+ $X2=4.405 $Y2=1.535
r93 42 43 9.37222 $w=3.6e-07 $l=7e-08 $layer=POLY_cond $X=3.975 $Y=1.535
+ $X2=4.045 $Y2=1.535
r94 40 42 11.3806 $w=3.6e-07 $l=8.5e-08 $layer=POLY_cond $X=3.89 $Y=1.535
+ $X2=3.975 $Y2=1.535
r95 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.89
+ $Y=1.51 $X2=3.89 $Y2=1.51
r96 38 40 36.8194 $w=3.6e-07 $l=2.75e-07 $layer=POLY_cond $X=3.615 $Y=1.535
+ $X2=3.89 $Y2=1.535
r97 37 38 20.0833 $w=3.6e-07 $l=1.5e-07 $layer=POLY_cond $X=3.465 $Y=1.535
+ $X2=3.615 $Y2=1.535
r98 36 37 37.4889 $w=3.6e-07 $l=2.8e-07 $layer=POLY_cond $X=3.185 $Y=1.535
+ $X2=3.465 $Y2=1.535
r99 31 48 0.324632 $w=3.53e-07 $l=1e-08 $layer=LI1_cond $X=4.56 $Y=1.582
+ $X2=4.57 $Y2=1.582
r100 30 31 15.5823 $w=3.53e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.582
+ $X2=4.56 $Y2=1.582
r101 30 41 6.168 $w=3.53e-07 $l=1.9e-07 $layer=LI1_cond $X=4.08 $Y=1.582
+ $X2=3.89 $Y2=1.582
r102 29 41 9.41432 $w=3.53e-07 $l=2.9e-07 $layer=LI1_cond $X=3.6 $Y=1.582
+ $X2=3.89 $Y2=1.582
r103 25 45 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.475 $Y=1.345
+ $X2=4.475 $Y2=1.535
r104 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.475 $Y=1.345
+ $X2=4.475 $Y2=0.655
r105 22 44 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.405 $Y=1.725
+ $X2=4.405 $Y2=1.535
r106 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.405 $Y=1.725
+ $X2=4.405 $Y2=2.465
r107 18 43 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.045 $Y=1.345
+ $X2=4.045 $Y2=1.535
r108 18 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.045 $Y=1.345
+ $X2=4.045 $Y2=0.655
r109 15 42 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.975 $Y=1.725
+ $X2=3.975 $Y2=1.535
r110 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.975 $Y=1.725
+ $X2=3.975 $Y2=2.465
r111 11 38 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.615 $Y=1.345
+ $X2=3.615 $Y2=1.535
r112 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.615 $Y=1.345
+ $X2=3.615 $Y2=0.655
r113 8 37 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.465 $Y=1.725
+ $X2=3.465 $Y2=1.535
r114 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.465 $Y=1.725
+ $X2=3.465 $Y2=2.465
r115 4 36 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.185 $Y=1.345
+ $X2=3.185 $Y2=1.535
r116 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.185 $Y=1.345
+ $X2=3.185 $Y2=0.655
r117 1 36 20.0833 $w=3.6e-07 $l=2.54165e-07 $layer=POLY_cond $X=3.035 $Y=1.725
+ $X2=3.185 $Y2=1.535
r118 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.035 $Y=1.725
+ $X2=3.035 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%C 3 7 11 15 19 23 27 31 33 34 35 36 37 62
c76 37 0 2.98258e-20 $X=6.96 $Y=1.665
r77 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.815
+ $Y=1.51 $X2=6.815 $Y2=1.51
r78 60 62 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.715 $Y=1.51
+ $X2=6.815 $Y2=1.51
r79 59 60 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=6.31 $Y=1.51
+ $X2=6.715 $Y2=1.51
r80 58 59 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=6.285 $Y=1.51
+ $X2=6.31 $Y2=1.51
r81 56 58 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.135 $Y=1.51
+ $X2=6.285 $Y2=1.51
r82 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.135
+ $Y=1.51 $X2=6.135 $Y2=1.51
r83 54 56 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=5.88 $Y=1.51
+ $X2=6.135 $Y2=1.51
r84 53 54 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.855 $Y=1.51
+ $X2=5.88 $Y2=1.51
r85 51 53 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.795 $Y=1.51
+ $X2=5.855 $Y2=1.51
r86 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.795
+ $Y=1.51 $X2=5.795 $Y2=1.51
r87 48 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.455 $Y=1.51
+ $X2=5.795 $Y2=1.51
r88 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.455
+ $Y=1.51 $X2=5.455 $Y2=1.51
r89 46 48 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=5.45 $Y=1.51
+ $X2=5.455 $Y2=1.51
r90 45 46 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.425 $Y=1.51
+ $X2=5.45 $Y2=1.51
r91 43 45 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=5.02 $Y=1.51
+ $X2=5.425 $Y2=1.51
r92 37 63 4.70716 $w=3.53e-07 $l=1.45e-07 $layer=LI1_cond $X=6.96 $Y=1.582
+ $X2=6.815 $Y2=1.582
r93 36 63 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=6.48 $Y=1.582
+ $X2=6.815 $Y2=1.582
r94 36 57 11.1998 $w=3.53e-07 $l=3.45e-07 $layer=LI1_cond $X=6.48 $Y=1.582
+ $X2=6.135 $Y2=1.582
r95 35 57 4.38253 $w=3.53e-07 $l=1.35e-07 $layer=LI1_cond $X=6 $Y=1.582
+ $X2=6.135 $Y2=1.582
r96 35 52 6.65495 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=6 $Y=1.582
+ $X2=5.795 $Y2=1.582
r97 34 52 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=5.52 $Y=1.582
+ $X2=5.795 $Y2=1.582
r98 34 49 2.11011 $w=3.53e-07 $l=6.5e-08 $layer=LI1_cond $X=5.52 $Y=1.582
+ $X2=5.455 $Y2=1.582
r99 33 49 13.4722 $w=3.53e-07 $l=4.15e-07 $layer=LI1_cond $X=5.04 $Y=1.582
+ $X2=5.455 $Y2=1.582
r100 29 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.345
+ $X2=6.715 $Y2=1.51
r101 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.715 $Y=1.345
+ $X2=6.715 $Y2=0.655
r102 25 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.31 $Y=1.675
+ $X2=6.31 $Y2=1.51
r103 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.31 $Y=1.675
+ $X2=6.31 $Y2=2.465
r104 21 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.285 $Y=1.345
+ $X2=6.285 $Y2=1.51
r105 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.285 $Y=1.345
+ $X2=6.285 $Y2=0.655
r106 17 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.88 $Y=1.675
+ $X2=5.88 $Y2=1.51
r107 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.88 $Y=1.675
+ $X2=5.88 $Y2=2.465
r108 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.855 $Y=1.345
+ $X2=5.855 $Y2=1.51
r109 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.855 $Y=1.345
+ $X2=5.855 $Y2=0.655
r110 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.45 $Y=1.675
+ $X2=5.45 $Y2=1.51
r111 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.45 $Y=1.675
+ $X2=5.45 $Y2=2.465
r112 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.425 $Y=1.345
+ $X2=5.425 $Y2=1.51
r113 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.425 $Y=1.345
+ $X2=5.425 $Y2=0.655
r114 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.02 $Y=1.675
+ $X2=5.02 $Y2=1.51
r115 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.02 $Y=1.675
+ $X2=5.02 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%VPWR 1 2 3 4 5 6 7 24 30 34 38 40 44 46 50
+ 52 56 60 65 66 67 68 69 78 85 86 89 92 95 98 101
r106 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r107 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 86 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r113 83 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.525 $Y2=3.33
r114 83 85 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 82 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r116 82 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r117 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r118 79 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.665 $Y2=3.33
r119 79 81 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.83 $Y=3.33 $X2=6
+ $Y2=3.33
r120 78 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.36 $Y=3.33
+ $X2=6.525 $Y2=3.33
r121 78 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.36 $Y=3.33 $X2=6
+ $Y2=3.33
r122 77 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r123 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 73 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 69 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 69 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 69 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 67 76 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.68 $Y2=3.33
r130 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.93 $Y2=3.33
r131 65 72 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 65 66 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=1.047 $Y2=3.33
r133 64 76 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=1.68 $Y2=3.33
r134 64 66 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=1.047 $Y2=3.33
r135 60 63 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=6.525 $Y=2.015
+ $X2=6.525 $Y2=2.95
r136 58 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=3.245
+ $X2=6.525 $Y2=3.33
r137 58 63 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.525 $Y=3.245
+ $X2=6.525 $Y2=2.95
r138 54 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=3.245
+ $X2=5.665 $Y2=3.33
r139 54 56 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.665 $Y=3.245
+ $X2=5.665 $Y2=2.385
r140 53 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=4.7 $Y2=3.33
r141 52 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=5.665 $Y2=3.33
r142 52 53 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=4.865 $Y2=3.33
r143 48 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=3.245 $X2=4.7
+ $Y2=3.33
r144 48 50 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=4.7 $Y=3.245
+ $X2=4.7 $Y2=2.375
r145 47 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=3.715 $Y2=3.33
r146 46 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=3.33
+ $X2=4.7 $Y2=3.33
r147 46 47 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.535 $Y=3.33
+ $X2=3.88 $Y2=3.33
r148 42 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=3.245
+ $X2=3.715 $Y2=3.33
r149 42 44 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=3.715 $Y=3.245
+ $X2=3.715 $Y2=2.38
r150 41 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=3.33
+ $X2=2.79 $Y2=3.33
r151 40 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=3.715 $Y2=3.33
r152 40 41 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=2.955 $Y2=3.33
r153 36 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=3.33
r154 36 38 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=2.78
r155 35 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.93 $Y2=3.33
r156 34 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.79 $Y2=3.33
r157 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.095 $Y2=3.33
r158 30 33 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.93 $Y=2.2
+ $X2=1.93 $Y2=2.97
r159 28 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r160 28 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.97
r161 24 27 38.5545 $w=2.73e-07 $l=9.2e-07 $layer=LI1_cond $X=1.047 $Y=2.05
+ $X2=1.047 $Y2=2.97
r162 22 66 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.047 $Y=3.245
+ $X2=1.047 $Y2=3.33
r163 22 27 11.5244 $w=2.73e-07 $l=2.75e-07 $layer=LI1_cond $X=1.047 $Y=3.245
+ $X2=1.047 $Y2=2.97
r164 7 63 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.385
+ $Y=1.835 $X2=6.525 $Y2=2.95
r165 7 60 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=6.385
+ $Y=1.835 $X2=6.525 $Y2=2.015
r166 6 56 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=5.525
+ $Y=1.835 $X2=5.665 $Y2=2.385
r167 5 50 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=4.48
+ $Y=1.835 $X2=4.7 $Y2=2.375
r168 4 44 300 $w=1.7e-07 $l=6.26418e-07 $layer=licon1_PDIFF $count=2 $X=3.54
+ $Y=1.835 $X2=3.715 $Y2=2.38
r169 3 38 600 $w=1.7e-07 $l=1.01258e-06 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.835 $X2=2.79 $Y2=2.78
r170 2 33 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=2.97
r171 2 30 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=2.2
r172 1 27 400 $w=1.7e-07 $l=1.22864e-06 $layer=licon1_PDIFF $count=1 $X=0.865
+ $Y=1.835 $X2=1.06 $Y2=2.97
r173 1 24 400 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_PDIFF $count=1 $X=0.865
+ $Y=1.835 $X2=1.06 $Y2=2.05
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%Y 1 2 3 4 5 6 7 8 27 33 35 36 37 38 43 45
+ 47 48 51 53 57 59 61 63 65 67 69 72 73 83 88 91 97 99
c123 83 0 6.17957e-20 $X=3.062 $Y=1.352
r124 106 107 0.192126 $w=7.62e-07 $l=1.2e-08 $layer=LI1_cond $X=3.25 $Y=2.09
+ $X2=3.262 $Y2=2.09
r125 99 101 11.2394 $w=7.62e-07 $l=7.02e-07 $layer=LI1_cond $X=2.36 $Y=2.09
+ $X2=3.062 $Y2=2.09
r126 84 101 6.57024 $w=2.85e-07 $l=4e-07 $layer=LI1_cond $X=3.062 $Y=1.69
+ $X2=3.062 $Y2=2.09
r127 84 88 1.01091 $w=2.83e-07 $l=2.5e-08 $layer=LI1_cond $X=3.062 $Y=1.69
+ $X2=3.062 $Y2=1.665
r128 83 97 3.24541 $w=2.85e-07 $l=5.7e-08 $layer=LI1_cond $X=3.062 $Y=1.352
+ $X2=3.062 $Y2=1.295
r129 73 107 7.78155 $w=2.35e-07 $l=4e-07 $layer=LI1_cond $X=3.262 $Y=2.49
+ $X2=3.262 $Y2=2.09
r130 73 106 2.08136 $w=7.62e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=2.09
+ $X2=3.25 $Y2=2.09
r131 73 101 0.928609 $w=7.62e-07 $l=5.8e-08 $layer=LI1_cond $X=3.12 $Y=2.09
+ $X2=3.062 $Y2=2.09
r132 73 91 2.07227 $w=2.93e-07 $l=4e-08 $layer=LI1_cond $X=3.262 $Y=2.49
+ $X2=3.262 $Y2=2.53
r133 73 88 1.2131 $w=2.83e-07 $l=3e-08 $layer=LI1_cond $X=3.062 $Y=1.635
+ $X2=3.062 $Y2=1.665
r134 72 97 0.801878 $w=2.13e-07 $l=1.4e-08 $layer=LI1_cond $X=3.062 $Y=1.281
+ $X2=3.062 $Y2=1.295
r135 72 94 12.6582 $w=2.13e-07 $l=2.21e-07 $layer=LI1_cond $X=3.062 $Y=1.281
+ $X2=3.062 $Y2=1.06
r136 72 73 10.8774 $w=2.83e-07 $l=2.69e-07 $layer=LI1_cond $X=3.062 $Y=1.366
+ $X2=3.062 $Y2=1.635
r137 72 83 0.566112 $w=2.83e-07 $l=1.4e-08 $layer=LI1_cond $X=3.062 $Y=1.366
+ $X2=3.062 $Y2=1.352
r138 61 71 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.095 $Y=2.1
+ $X2=6.095 $Y2=2.015
r139 61 63 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=6.095 $Y=2.1
+ $X2=6.095 $Y2=2.91
r140 60 69 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=5.33 $Y=2.015
+ $X2=5.182 $Y2=2.015
r141 59 71 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6 $Y=2.015 $X2=6.095
+ $Y2=2.015
r142 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6 $Y=2.015 $X2=5.33
+ $Y2=2.015
r143 55 69 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.182 $Y=2.1
+ $X2=5.182 $Y2=2.015
r144 55 57 31.6434 $w=2.93e-07 $l=8.1e-07 $layer=LI1_cond $X=5.182 $Y=2.1
+ $X2=5.182 $Y2=2.91
r145 54 67 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=4.365 $Y=2.015
+ $X2=4.207 $Y2=2.015
r146 53 69 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=5.035 $Y=2.015
+ $X2=5.182 $Y2=2.015
r147 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.035 $Y=2.015
+ $X2=4.365 $Y2=2.015
r148 49 67 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.207 $Y=2.1
+ $X2=4.207 $Y2=2.015
r149 49 51 29.6342 $w=3.13e-07 $l=8.1e-07 $layer=LI1_cond $X=4.207 $Y=2.1
+ $X2=4.207 $Y2=2.91
r150 48 107 10.6698 $w=7.62e-07 $l=1.50911e-07 $layer=LI1_cond $X=3.38 $Y=2.015
+ $X2=3.262 $Y2=2.09
r151 47 67 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=4.05 $Y=2.015
+ $X2=4.207 $Y2=2.015
r152 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.05 $Y=2.015
+ $X2=3.38 $Y2=2.015
r153 46 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.635 $Y=1.06
+ $X2=2.54 $Y2=1.06
r154 45 94 2.0603 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=2.92 $Y=1.06
+ $X2=3.062 $Y2=1.06
r155 45 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.92 $Y=1.06
+ $X2=2.635 $Y2=1.06
r156 41 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.975
+ $X2=2.54 $Y2=1.06
r157 41 43 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.54 $Y=0.975
+ $X2=2.54 $Y2=0.76
r158 37 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.445 $Y=1.06
+ $X2=2.54 $Y2=1.06
r159 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.445 $Y=1.06
+ $X2=1.775 $Y2=1.06
r160 35 99 7.31617 $w=7.62e-07 $l=3.16961e-07 $layer=LI1_cond $X=2.265 $Y=1.817
+ $X2=2.36 $Y2=2.09
r161 35 36 30.2799 $w=2.53e-07 $l=6.7e-07 $layer=LI1_cond $X=2.265 $Y=1.817
+ $X2=1.595 $Y2=1.817
r162 31 38 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.645 $Y=0.975
+ $X2=1.775 $Y2=1.06
r163 31 33 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=1.645 $Y=0.975
+ $X2=1.645 $Y2=0.76
r164 27 29 45.6175 $w=2.38e-07 $l=9.5e-07 $layer=LI1_cond $X=1.475 $Y=1.96
+ $X2=1.475 $Y2=2.91
r165 25 36 6.82464 $w=2.55e-07 $l=1.78168e-07 $layer=LI1_cond $X=1.475 $Y=1.945
+ $X2=1.595 $Y2=1.817
r166 25 27 0.720277 $w=2.38e-07 $l=1.5e-08 $layer=LI1_cond $X=1.475 $Y=1.945
+ $X2=1.475 $Y2=1.96
r167 8 71 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=5.955
+ $Y=1.835 $X2=6.095 $Y2=2.095
r168 8 63 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.955
+ $Y=1.835 $X2=6.095 $Y2=2.91
r169 7 69 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.835 $X2=5.235 $Y2=2.095
r170 7 57 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.835 $X2=5.235 $Y2=2.91
r171 6 67 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=4.05
+ $Y=1.835 $X2=4.19 $Y2=2.095
r172 6 51 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.05
+ $Y=1.835 $X2=4.19 $Y2=2.91
r173 5 106 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=1.835 $X2=3.25 $Y2=2.095
r174 5 91 300 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=2 $X=3.11
+ $Y=1.835 $X2=3.25 $Y2=2.53
r175 4 99 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=2.22
+ $Y=1.835 $X2=2.36 $Y2=2.475
r176 4 99 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.835 $X2=2.36 $Y2=1.96
r177 3 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.91
r178 3 27 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=1.96
r179 2 43 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.235 $X2=2.54 $Y2=0.76
r180 1 33 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.235 $X2=1.68 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%VGND 1 2 3 4 15 19 23 25 27 30 31 32 34 46
+ 50 56 59 63
r98 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r99 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r100 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 54 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r102 54 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r103 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r104 51 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=0 $X2=6.07
+ $Y2=0
r105 51 53 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.235 $Y=0 $X2=6.48
+ $Y2=0
r106 50 62 4.42457 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.8 $Y=0 $X2=7 $Y2=0
r107 50 53 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.8 $Y=0 $X2=6.48
+ $Y2=0
r108 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r109 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r110 46 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.905 $Y=0 $X2=6.07
+ $Y2=0
r111 46 48 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=5.52 $Y2=0
r112 45 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r113 44 45 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r114 42 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r115 41 44 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r116 41 42 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r117 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r118 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r119 37 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r120 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r121 34 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r122 34 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0
+ $X2=0.24 $Y2=0
r123 32 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r124 32 42 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=1.2
+ $Y2=0
r125 30 44 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.04
+ $Y2=0
r126 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.21
+ $Y2=0
r127 29 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.52 $Y2=0
r128 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=0 $X2=5.21
+ $Y2=0
r129 25 62 3.05295 $w=2.95e-07 $l=1.08305e-07 $layer=LI1_cond $X=6.947 $Y=0.085
+ $X2=7 $Y2=0
r130 25 27 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=6.947 $Y=0.085
+ $X2=6.947 $Y2=0.38
r131 21 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0
r132 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0.36
r133 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=0.085
+ $X2=5.21 $Y2=0
r134 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.21 $Y=0.085
+ $X2=5.21 $Y2=0.38
r135 13 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r136 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.585
r137 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.79
+ $Y=0.235 $X2=6.93 $Y2=0.38
r138 3 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.93
+ $Y=0.235 $X2=6.07 $Y2=0.36
r139 2 19 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.085
+ $Y=0.235 $X2=5.21 $Y2=0.38
r140 1 15 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%A_225_47# 1 2 3 4 5 18 20 21 24 28 32 37 39
+ 41 43
c82 39 0 5.86634e-20 $X=2.97 $Y=0.36
r83 33 41 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.995 $Y=0.35
+ $X2=3.83 $Y2=0.35
r84 32 43 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=0.35
+ $X2=4.69 $Y2=0.35
r85 32 33 30.9378 $w=1.88e-07 $l=5.3e-07 $layer=LI1_cond $X=4.525 $Y=0.35
+ $X2=3.995 $Y2=0.35
r86 29 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0.35
+ $X2=2.97 $Y2=0.35
r87 28 41 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=0.35
+ $X2=3.83 $Y2=0.35
r88 28 29 30.9378 $w=1.88e-07 $l=5.3e-07 $layer=LI1_cond $X=3.665 $Y=0.35
+ $X2=3.135 $Y2=0.35
r89 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0.34
+ $X2=2.11 $Y2=0.34
r90 24 39 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.805 $Y=0.34
+ $X2=2.97 $Y2=0.35
r91 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.805 $Y=0.34
+ $X2=2.275 $Y2=0.34
r92 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0.34
+ $X2=2.11 $Y2=0.34
r93 20 21 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.945 $Y=0.34
+ $X2=1.345 $Y2=0.34
r94 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.215 $Y=0.425
+ $X2=1.345 $Y2=0.34
r95 16 18 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=1.215 $Y=0.425
+ $X2=1.215 $Y2=0.535
r96 5 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.55
+ $Y=0.235 $X2=4.69 $Y2=0.38
r97 4 41 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.69
+ $Y=0.235 $X2=3.83 $Y2=0.36
r98 3 39 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.83
+ $Y=0.235 $X2=2.97 $Y2=0.36
r99 2 37 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.97
+ $Y=0.235 $X2=2.11 $Y2=0.36
r100 1 18 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_4%A_652_47# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
r53 31 33 33.0367 $w=2.23e-07 $l=6.45e-07 $layer=LI1_cond $X=6.517 $Y=1.065
+ $X2=6.517 $Y2=0.42
r54 30 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.735 $Y=1.15
+ $X2=5.64 $Y2=1.15
r55 29 31 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=6.405 $Y=1.15
+ $X2=6.517 $Y2=1.065
r56 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.405 $Y=1.15
+ $X2=5.735 $Y2=1.15
r57 25 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=1.065
+ $X2=5.64 $Y2=1.15
r58 25 27 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=5.64 $Y=1.065
+ $X2=5.64 $Y2=0.42
r59 24 35 4.47804 $w=2.25e-07 $l=1.19373e-07 $layer=LI1_cond $X=4.355 $Y=1.15
+ $X2=4.26 $Y2=1.095
r60 23 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.545 $Y=1.15
+ $X2=5.64 $Y2=1.15
r61 23 24 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=5.545 $Y=1.15
+ $X2=4.355 $Y2=1.15
r62 19 35 1.9579 $w=1.9e-07 $l=1.4e-07 $layer=LI1_cond $X=4.26 $Y=0.955 $X2=4.26
+ $Y2=1.095
r63 19 21 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=4.26 $Y=0.955
+ $X2=4.26 $Y2=0.78
r64 17 35 4.47804 $w=2.25e-07 $l=9.5e-08 $layer=LI1_cond $X=4.165 $Y=1.095
+ $X2=4.26 $Y2=1.095
r65 17 18 27.5763 $w=2.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.165 $Y=1.095
+ $X2=3.495 $Y2=1.095
r66 13 18 6.11365 $w=2.74e-07 $l=1.81384e-07 $layer=LI1_cond $X=3.4 $Y=0.955
+ $X2=3.495 $Y2=1.095
r67 13 15 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=3.4 $Y=0.955
+ $X2=3.4 $Y2=0.78
r68 4 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.36
+ $Y=0.235 $X2=6.5 $Y2=0.42
r69 3 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.5
+ $Y=0.235 $X2=5.64 $Y2=0.42
r70 2 21 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=4.12
+ $Y=0.235 $X2=4.26 $Y2=0.78
r71 1 15 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=3.26
+ $Y=0.235 $X2=3.4 $Y2=0.78
.ends

