* File: sky130_fd_sc_lp__a32o_lp.pxi.spice
* Created: Wed Sep  2 09:27:55 2020
* 
x_PM_SKY130_FD_SC_LP__A32O_LP%B2 N_B2_M1006_g N_B2_M1001_g N_B2_c_76_n
+ N_B2_c_77_n N_B2_c_82_n B2 N_B2_c_78_n N_B2_c_79_n
+ PM_SKY130_FD_SC_LP__A32O_LP%B2
x_PM_SKY130_FD_SC_LP__A32O_LP%B1 N_B1_M1010_g N_B1_c_112_n N_B1_M1000_g
+ N_B1_c_108_n N_B1_c_109_n B1 N_B1_c_111_n PM_SKY130_FD_SC_LP__A32O_LP%B1
x_PM_SKY130_FD_SC_LP__A32O_LP%A1 N_A1_M1008_g N_A1_M1007_g N_A1_c_153_n
+ N_A1_c_154_n N_A1_c_159_n A1 N_A1_c_155_n N_A1_c_156_n
+ PM_SKY130_FD_SC_LP__A32O_LP%A1
x_PM_SKY130_FD_SC_LP__A32O_LP%A2 N_A2_M1011_g N_A2_c_201_n N_A2_M1012_g
+ N_A2_c_197_n N_A2_c_198_n A2 A2 A2 N_A2_c_200_n PM_SKY130_FD_SC_LP__A32O_LP%A2
x_PM_SKY130_FD_SC_LP__A32O_LP%A3 N_A3_M1009_g N_A3_M1003_g A3 N_A3_c_244_n
+ PM_SKY130_FD_SC_LP__A32O_LP%A3
x_PM_SKY130_FD_SC_LP__A32O_LP%A_137_419# N_A_137_419#_M1010_d
+ N_A_137_419#_M1006_d N_A_137_419#_c_281_n N_A_137_419#_M1005_g
+ N_A_137_419#_M1002_g N_A_137_419#_c_283_n N_A_137_419#_M1004_g
+ N_A_137_419#_c_298_n N_A_137_419#_c_295_n N_A_137_419#_c_296_n
+ N_A_137_419#_c_285_n N_A_137_419#_c_286_n N_A_137_419#_c_287_n
+ N_A_137_419#_c_288_n N_A_137_419#_c_289_n N_A_137_419#_c_290_n
+ N_A_137_419#_c_291_n N_A_137_419#_c_292_n N_A_137_419#_c_293_n
+ PM_SKY130_FD_SC_LP__A32O_LP%A_137_419#
x_PM_SKY130_FD_SC_LP__A32O_LP%A_30_419# N_A_30_419#_M1006_s N_A_30_419#_M1000_d
+ N_A_30_419#_M1012_d N_A_30_419#_c_390_n N_A_30_419#_c_395_n
+ N_A_30_419#_c_391_n N_A_30_419#_c_397_n N_A_30_419#_c_404_n
+ N_A_30_419#_c_401_n N_A_30_419#_c_406_n PM_SKY130_FD_SC_LP__A32O_LP%A_30_419#
x_PM_SKY130_FD_SC_LP__A32O_LP%VPWR N_VPWR_M1007_d N_VPWR_M1003_d N_VPWR_c_440_n
+ N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n VPWR N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_439_n N_VPWR_c_447_n PM_SKY130_FD_SC_LP__A32O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A32O_LP%X N_X_M1002_d N_X_M1004_d X X X X X X X
+ PM_SKY130_FD_SC_LP__A32O_LP%X
x_PM_SKY130_FD_SC_LP__A32O_LP%VGND N_VGND_M1001_s N_VGND_M1009_d N_VGND_c_506_n
+ N_VGND_c_507_n N_VGND_c_508_n VGND N_VGND_c_509_n N_VGND_c_510_n
+ N_VGND_c_511_n N_VGND_c_512_n PM_SKY130_FD_SC_LP__A32O_LP%VGND
cc_1 VNB N_B2_c_76_n 0.0216299f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.235
cc_2 VNB N_B2_c_77_n 0.0191034f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.74
cc_3 VNB N_B2_c_78_n 0.0170897f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_4 VNB N_B2_c_79_n 0.0258946f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_5 VNB N_B1_c_108_n 0.0185972f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.235
cc_6 VNB N_B1_c_109_n 0.0147879f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.74
cc_7 VNB B1 0.00611839f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.905
cc_8 VNB N_B1_c_111_n 0.0176707f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_9 VNB N_A1_c_153_n 0.018412f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.235
cc_10 VNB N_A1_c_154_n 0.0179472f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.74
cc_11 VNB N_A1_c_155_n 0.0167497f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_12 VNB N_A1_c_156_n 0.00294366f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_13 VNB N_A2_c_197_n 0.0175392f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.235
cc_14 VNB N_A2_c_198_n 0.0163639f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.74
cc_15 VNB A2 0.00493854f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.905
cc_16 VNB N_A2_c_200_n 0.0157387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_M1009_g 0.0391379f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_18 VNB A3 0.00310189f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.235
cc_19 VNB N_A3_c_244_n 0.0236715f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_20 VNB N_A_137_419#_c_281_n 0.0164444f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.915
cc_21 VNB N_A_137_419#_M1002_g 0.0178043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_137_419#_c_283_n 0.0172917f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_23 VNB N_A_137_419#_M1004_g 0.0159985f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.4
cc_24 VNB N_A_137_419#_c_285_n 0.00104921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_137_419#_c_286_n 0.0314623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_137_419#_c_287_n 0.00662092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_137_419#_c_288_n 0.0013348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_137_419#_c_289_n 0.00174367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_137_419#_c_290_n 0.029654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_137_419#_c_291_n 0.00243016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_137_419#_c_292_n 0.00108937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_137_419#_c_293_n 0.0568263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_439_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.0582901f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.915
cc_35 VNB N_VGND_c_506_n 0.0158851f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.915
cc_36 VNB N_VGND_c_507_n 0.0497917f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.235
cc_37 VNB N_VGND_c_508_n 0.0227238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_509_n 0.0654219f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.57
cc_39 VNB N_VGND_c_510_n 0.0333408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_511_n 0.290733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_512_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_B2_M1006_g 0.0359013f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.595
cc_43 VPB N_B2_c_77_n 0.00631765f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.74
cc_44 VPB N_B2_c_82_n 0.0144588f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.905
cc_45 VPB N_B2_c_79_n 0.0145083f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.4
cc_46 VPB N_B1_c_112_n 0.0116807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B1_M1000_g 0.0277452f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.915
cc_48 VPB N_B1_c_109_n 0.00489048f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.74
cc_49 VPB B1 0.00386728f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.905
cc_50 VPB N_A1_M1007_g 0.0284456f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.915
cc_51 VPB N_A1_c_154_n 0.00593531f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.74
cc_52 VPB N_A1_c_159_n 0.0138958f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.905
cc_53 VPB N_A1_c_156_n 7.56276e-19 $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.4
cc_54 VPB N_A2_c_201_n 0.0128849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A2_M1012_g 0.0286324f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.915
cc_56 VPB N_A2_c_198_n 0.0054117f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.74
cc_57 VPB A2 0.00262925f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.905
cc_58 VPB N_A3_M1003_g 0.0366767f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.915
cc_59 VPB A3 0.00318476f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.235
cc_60 VPB N_A3_c_244_n 0.0343239f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.4
cc_61 VPB N_A_137_419#_M1004_g 0.060478f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.4
cc_62 VPB N_A_137_419#_c_295_n 0.0219473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_137_419#_c_296_n 0.00993484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_137_419#_c_289_n 0.00331746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_30_419#_c_390_n 0.0334046f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_66 VPB N_A_30_419#_c_391_n 0.0071976f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.4
cc_67 VPB N_VPWR_c_440_n 0.002833f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.235
cc_68 VPB N_VPWR_c_441_n 0.00832351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_442_n 0.0422809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_443_n 0.00506702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_444_n 0.0237058f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_445_n 0.0329154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_439_n 0.0469352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_447_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB X 0.0555816f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.915
cc_76 N_B2_c_82_n N_B1_c_112_n 0.0177796f $X=0.52 $Y=1.905 $X2=0 $Y2=0
cc_77 N_B2_M1006_g N_B1_M1000_g 0.044871f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_78 N_B2_c_76_n N_B1_c_108_n 0.0177796f $X=0.52 $Y=1.235 $X2=0 $Y2=0
cc_79 N_B2_c_77_n N_B1_c_109_n 0.0177796f $X=0.52 $Y=1.74 $X2=0 $Y2=0
cc_80 N_B2_c_78_n B1 8.513e-19 $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_81 N_B2_c_79_n B1 0.0403261f $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_82 N_B2_c_78_n N_B1_c_111_n 0.0177796f $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_83 N_B2_c_79_n N_B1_c_111_n 8.4747e-19 $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_84 N_B2_M1006_g N_A_137_419#_c_298_n 0.00980901f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_85 N_B2_M1006_g N_A_137_419#_c_296_n 0.00484805f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_86 N_B2_c_79_n N_A_137_419#_c_296_n 0.00199742f $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_87 N_B2_M1006_g N_A_30_419#_c_390_n 0.0199864f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_88 N_B2_c_82_n N_A_30_419#_c_390_n 0.00213543f $X=0.52 $Y=1.905 $X2=0 $Y2=0
cc_89 N_B2_c_79_n N_A_30_419#_c_390_n 0.0287632f $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_90 N_B2_M1006_g N_A_30_419#_c_395_n 0.0167335f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_91 N_B2_M1006_g N_A_30_419#_c_391_n 6.00691e-19 $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_92 N_B2_M1006_g N_A_30_419#_c_397_n 8.38214e-19 $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_93 N_B2_M1006_g N_VPWR_c_442_n 0.00599906f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_94 N_B2_M1006_g N_VPWR_c_439_n 0.00882257f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_95 N_B2_c_76_n N_VGND_c_507_n 0.0125217f $X=0.52 $Y=1.235 $X2=0 $Y2=0
cc_96 N_B2_c_78_n N_VGND_c_507_n 0.00466416f $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_97 N_B2_c_79_n N_VGND_c_507_n 0.0253051f $X=0.52 $Y=1.4 $X2=0 $Y2=0
cc_98 N_B2_c_76_n N_VGND_c_509_n 0.0031218f $X=0.52 $Y=1.235 $X2=0 $Y2=0
cc_99 N_B2_c_76_n N_VGND_c_511_n 0.00376215f $X=0.52 $Y=1.235 $X2=0 $Y2=0
cc_100 N_B1_M1000_g N_A1_M1007_g 0.0456085f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_101 N_B1_c_108_n N_A1_c_153_n 0.0124338f $X=1.09 $Y=1.235 $X2=0 $Y2=0
cc_102 N_B1_c_109_n N_A1_c_154_n 0.0117589f $X=1.09 $Y=1.74 $X2=0 $Y2=0
cc_103 N_B1_c_112_n N_A1_c_159_n 0.0117589f $X=1.09 $Y=1.905 $X2=0 $Y2=0
cc_104 B1 N_A1_c_155_n 0.00410596f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_105 N_B1_c_111_n N_A1_c_155_n 0.0117589f $X=1.09 $Y=1.4 $X2=0 $Y2=0
cc_106 B1 N_A1_c_156_n 0.0514906f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B1_c_111_n N_A1_c_156_n 7.5249e-19 $X=1.09 $Y=1.4 $X2=0 $Y2=0
cc_108 N_B1_M1000_g N_A_137_419#_c_298_n 0.0100859f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_109 N_B1_c_112_n N_A_137_419#_c_295_n 0.00103139f $X=1.09 $Y=1.905 $X2=0
+ $Y2=0
cc_110 N_B1_M1000_g N_A_137_419#_c_295_n 0.0146437f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_111 B1 N_A_137_419#_c_295_n 0.024121f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_112 N_B1_c_112_n N_A_137_419#_c_296_n 0.00107953f $X=1.09 $Y=1.905 $X2=0
+ $Y2=0
cc_113 N_B1_M1000_g N_A_137_419#_c_296_n 0.00216399f $X=1.09 $Y=2.595 $X2=0
+ $Y2=0
cc_114 B1 N_A_137_419#_c_296_n 0.0053728f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_115 N_B1_c_108_n N_A_137_419#_c_285_n 0.00596098f $X=1.09 $Y=1.235 $X2=0
+ $Y2=0
cc_116 B1 N_A_137_419#_c_285_n 0.010476f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B1_c_111_n N_A_137_419#_c_285_n 0.00170912f $X=1.09 $Y=1.4 $X2=0 $Y2=0
cc_118 N_B1_c_108_n N_A_137_419#_c_287_n 8.68172e-19 $X=1.09 $Y=1.235 $X2=0
+ $Y2=0
cc_119 N_B1_M1000_g N_A_30_419#_c_390_n 0.00101601f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_120 N_B1_M1000_g N_A_30_419#_c_395_n 0.015535f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_121 N_B1_M1000_g N_A_30_419#_c_397_n 0.00545394f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_122 N_B1_M1000_g N_A_30_419#_c_401_n 0.00473007f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_123 N_B1_M1000_g N_VPWR_c_440_n 0.00110172f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_124 N_B1_M1000_g N_VPWR_c_442_n 0.00599906f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_125 N_B1_M1000_g N_VPWR_c_439_n 0.00796144f $X=1.09 $Y=2.595 $X2=0 $Y2=0
cc_126 N_B1_c_108_n N_VGND_c_507_n 0.00144874f $X=1.09 $Y=1.235 $X2=0 $Y2=0
cc_127 N_B1_c_108_n N_VGND_c_509_n 0.00375548f $X=1.09 $Y=1.235 $X2=0 $Y2=0
cc_128 N_B1_c_108_n N_VGND_c_511_n 0.00447875f $X=1.09 $Y=1.235 $X2=0 $Y2=0
cc_129 N_A1_c_159_n N_A2_c_201_n 0.01184f $X=1.66 $Y=1.905 $X2=0 $Y2=0
cc_130 N_A1_M1007_g N_A2_M1012_g 0.0411107f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_131 N_A1_c_153_n N_A2_c_197_n 0.017139f $X=1.66 $Y=1.235 $X2=0 $Y2=0
cc_132 N_A1_c_154_n N_A2_c_198_n 0.01184f $X=1.66 $Y=1.74 $X2=0 $Y2=0
cc_133 N_A1_c_153_n A2 0.00307688f $X=1.66 $Y=1.235 $X2=0 $Y2=0
cc_134 N_A1_c_155_n A2 0.00410205f $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_135 N_A1_c_156_n A2 0.0438819f $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_136 N_A1_c_155_n N_A2_c_200_n 0.01184f $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_137 N_A1_c_156_n N_A2_c_200_n 8.23261e-19 $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_138 N_A1_M1007_g N_A_137_419#_c_298_n 8.85073e-19 $X=1.62 $Y=2.595 $X2=0
+ $Y2=0
cc_139 N_A1_M1007_g N_A_137_419#_c_295_n 0.0153614f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_140 N_A1_c_159_n N_A_137_419#_c_295_n 5.43485e-19 $X=1.66 $Y=1.905 $X2=0
+ $Y2=0
cc_141 N_A1_c_156_n N_A_137_419#_c_295_n 0.0241279f $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_142 N_A1_c_153_n N_A_137_419#_c_285_n 0.00937242f $X=1.66 $Y=1.235 $X2=0
+ $Y2=0
cc_143 N_A1_c_156_n N_A_137_419#_c_285_n 0.00183793f $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_144 N_A1_c_153_n N_A_137_419#_c_286_n 0.00693417f $X=1.66 $Y=1.235 $X2=0
+ $Y2=0
cc_145 N_A1_c_155_n N_A_137_419#_c_286_n 8.97816e-19 $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_146 N_A1_c_156_n N_A_137_419#_c_286_n 0.00871406f $X=1.66 $Y=1.4 $X2=0 $Y2=0
cc_147 N_A1_c_153_n N_A_137_419#_c_287_n 0.00127765f $X=1.66 $Y=1.235 $X2=0
+ $Y2=0
cc_148 N_A1_M1007_g N_A_30_419#_c_395_n 0.00461641f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_149 N_A1_M1007_g N_A_30_419#_c_397_n 0.00569758f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_150 N_A1_M1007_g N_A_30_419#_c_404_n 0.0144834f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_151 N_A1_M1007_g N_A_30_419#_c_401_n 0.00216399f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_152 N_A1_M1007_g N_A_30_419#_c_406_n 6.91099e-19 $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_153 N_A1_M1007_g N_VPWR_c_440_n 0.0106626f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_154 N_A1_M1007_g N_VPWR_c_442_n 0.00642969f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_155 N_A1_M1007_g N_VPWR_c_439_n 0.00729472f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_156 N_A1_c_153_n N_VGND_c_509_n 5.91536e-19 $X=1.66 $Y=1.235 $X2=0 $Y2=0
cc_157 N_A2_c_197_n N_A3_M1009_g 0.016633f $X=2.23 $Y=1.235 $X2=0 $Y2=0
cc_158 A2 N_A3_M1009_g 0.00222727f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_159 N_A2_c_200_n N_A3_M1009_g 0.0117462f $X=2.23 $Y=1.4 $X2=0 $Y2=0
cc_160 N_A2_c_201_n N_A3_M1003_g 0.0117462f $X=2.23 $Y=1.905 $X2=0 $Y2=0
cc_161 N_A2_M1012_g N_A3_M1003_g 0.0434559f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_162 N_A2_c_198_n N_A3_c_244_n 0.0117462f $X=2.23 $Y=1.74 $X2=0 $Y2=0
cc_163 N_A2_c_201_n N_A_137_419#_c_295_n 5.43152e-19 $X=2.23 $Y=1.905 $X2=0
+ $Y2=0
cc_164 N_A2_M1012_g N_A_137_419#_c_295_n 0.0153755f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_165 A2 N_A_137_419#_c_295_n 0.0257713f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_166 N_A2_c_197_n N_A_137_419#_c_285_n 0.00106776f $X=2.23 $Y=1.235 $X2=0
+ $Y2=0
cc_167 N_A2_c_197_n N_A_137_419#_c_286_n 0.00706291f $X=2.23 $Y=1.235 $X2=0
+ $Y2=0
cc_168 A2 N_A_137_419#_c_286_n 0.0226185f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_169 N_A2_c_200_n N_A_137_419#_c_286_n 5.2374e-19 $X=2.23 $Y=1.4 $X2=0 $Y2=0
cc_170 N_A2_c_197_n N_A_137_419#_c_288_n 0.00405509f $X=2.23 $Y=1.235 $X2=0
+ $Y2=0
cc_171 A2 N_A_137_419#_c_288_n 0.0288788f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_172 N_A2_M1012_g N_A_137_419#_c_289_n 0.0035511f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_173 A2 N_A_137_419#_c_289_n 0.0385788f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_174 N_A2_c_200_n N_A_137_419#_c_289_n 0.00302898f $X=2.23 $Y=1.4 $X2=0 $Y2=0
cc_175 A2 N_A_137_419#_c_292_n 0.0139345f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_176 N_A2_c_200_n N_A_137_419#_c_292_n 8.86678e-19 $X=2.23 $Y=1.4 $X2=0 $Y2=0
cc_177 N_A2_M1012_g N_A_30_419#_c_397_n 7.81611e-19 $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_178 N_A2_M1012_g N_A_30_419#_c_404_n 0.0169455f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_179 N_A2_M1012_g N_A_30_419#_c_406_n 0.00973664f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_180 N_A2_M1012_g N_VPWR_c_440_n 0.00487432f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_181 N_A2_M1012_g N_VPWR_c_444_n 0.00718242f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_182 N_A2_M1012_g N_VPWR_c_439_n 0.00926181f $X=2.23 $Y=2.595 $X2=0 $Y2=0
cc_183 N_A2_c_197_n N_VGND_c_509_n 5.76631e-19 $X=2.23 $Y=1.235 $X2=0 $Y2=0
cc_184 A2 A_443_141# 0.0041903f $X=2.075 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_185 A3 N_A_137_419#_M1004_g 0.00140786f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A3_c_244_n N_A_137_419#_M1004_g 0.0102273f $X=3.09 $Y=1.715 $X2=0 $Y2=0
cc_187 N_A3_M1003_g N_A_137_419#_c_295_n 0.0100354f $X=2.76 $Y=2.595 $X2=0 $Y2=0
cc_188 N_A3_M1009_g N_A_137_419#_c_286_n 0.00359332f $X=2.71 $Y=0.915 $X2=0
+ $Y2=0
cc_189 N_A3_M1009_g N_A_137_419#_c_288_n 0.0152693f $X=2.71 $Y=0.915 $X2=0 $Y2=0
cc_190 N_A3_M1009_g N_A_137_419#_c_289_n 0.00910508f $X=2.71 $Y=0.915 $X2=0
+ $Y2=0
cc_191 N_A3_M1003_g N_A_137_419#_c_289_n 0.0105575f $X=2.76 $Y=2.595 $X2=0 $Y2=0
cc_192 A3 N_A_137_419#_c_289_n 0.0225103f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A3_c_244_n N_A_137_419#_c_289_n 0.00932426f $X=3.09 $Y=1.715 $X2=0
+ $Y2=0
cc_194 N_A3_M1009_g N_A_137_419#_c_290_n 0.00767149f $X=2.71 $Y=0.915 $X2=0
+ $Y2=0
cc_195 A3 N_A_137_419#_c_290_n 0.0237223f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A3_c_244_n N_A_137_419#_c_290_n 0.00791336f $X=3.09 $Y=1.715 $X2=0
+ $Y2=0
cc_197 N_A3_M1009_g N_A_137_419#_c_291_n 6.66262e-19 $X=2.71 $Y=0.915 $X2=0
+ $Y2=0
cc_198 N_A3_M1009_g N_A_137_419#_c_292_n 0.00256205f $X=2.71 $Y=0.915 $X2=0
+ $Y2=0
cc_199 N_A3_M1009_g N_A_137_419#_c_293_n 0.0120328f $X=2.71 $Y=0.915 $X2=0 $Y2=0
cc_200 N_A3_M1003_g N_A_30_419#_c_404_n 0.00440321f $X=2.76 $Y=2.595 $X2=0 $Y2=0
cc_201 N_A3_M1003_g N_A_30_419#_c_406_n 0.00870289f $X=2.76 $Y=2.595 $X2=0 $Y2=0
cc_202 N_A3_M1003_g N_VPWR_c_441_n 0.0271942f $X=2.76 $Y=2.595 $X2=0 $Y2=0
cc_203 A3 N_VPWR_c_441_n 0.0250595f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A3_c_244_n N_VPWR_c_441_n 0.00255109f $X=3.09 $Y=1.715 $X2=0 $Y2=0
cc_205 N_A3_M1003_g N_VPWR_c_444_n 0.00939541f $X=2.76 $Y=2.595 $X2=0 $Y2=0
cc_206 N_A3_M1003_g N_VPWR_c_439_n 0.0175663f $X=2.76 $Y=2.595 $X2=0 $Y2=0
cc_207 A3 X 0.00860964f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_208 N_A3_c_244_n X 0.0011325f $X=3.09 $Y=1.715 $X2=0 $Y2=0
cc_209 N_A3_M1009_g N_VGND_c_508_n 0.00367502f $X=2.71 $Y=0.915 $X2=0 $Y2=0
cc_210 N_A3_M1009_g N_VGND_c_509_n 0.00142392f $X=2.71 $Y=0.915 $X2=0 $Y2=0
cc_211 N_A3_M1009_g N_VGND_c_511_n 0.00119433f $X=2.71 $Y=0.915 $X2=0 $Y2=0
cc_212 N_A_137_419#_c_295_n N_A_30_419#_M1000_d 0.00180746f $X=2.575 $Y=2.17
+ $X2=0 $Y2=0
cc_213 N_A_137_419#_c_295_n N_A_30_419#_M1012_d 0.00176391f $X=2.575 $Y=2.17
+ $X2=0 $Y2=0
cc_214 N_A_137_419#_c_298_n N_A_30_419#_c_390_n 0.0302768f $X=0.825 $Y=2.4 $X2=0
+ $Y2=0
cc_215 N_A_137_419#_c_296_n N_A_30_419#_c_390_n 0.0119061f $X=0.99 $Y=2.17 $X2=0
+ $Y2=0
cc_216 N_A_137_419#_M1006_d N_A_30_419#_c_395_n 0.00340092f $X=0.685 $Y=2.095
+ $X2=0 $Y2=0
cc_217 N_A_137_419#_c_298_n N_A_30_419#_c_395_n 0.0152185f $X=0.825 $Y=2.4 $X2=0
+ $Y2=0
cc_218 N_A_137_419#_c_295_n N_A_30_419#_c_395_n 0.00447619f $X=2.575 $Y=2.17
+ $X2=0 $Y2=0
cc_219 N_A_137_419#_c_298_n N_A_30_419#_c_397_n 0.00721503f $X=0.825 $Y=2.4
+ $X2=0 $Y2=0
cc_220 N_A_137_419#_c_295_n N_A_30_419#_c_404_n 0.0628611f $X=2.575 $Y=2.17
+ $X2=0 $Y2=0
cc_221 N_A_137_419#_c_298_n N_A_30_419#_c_401_n 0.0119061f $X=0.825 $Y=2.4 $X2=0
+ $Y2=0
cc_222 N_A_137_419#_c_295_n N_A_30_419#_c_401_n 0.0164738f $X=2.575 $Y=2.17
+ $X2=0 $Y2=0
cc_223 N_A_137_419#_c_295_n N_VPWR_M1007_d 0.00268484f $X=2.575 $Y=2.17
+ $X2=-0.19 $Y2=-0.245
cc_224 N_A_137_419#_M1004_g N_VPWR_c_441_n 0.0233092f $X=3.775 $Y=2.595 $X2=0
+ $Y2=0
cc_225 N_A_137_419#_c_295_n N_VPWR_c_441_n 0.00719944f $X=2.575 $Y=2.17 $X2=0
+ $Y2=0
cc_226 N_A_137_419#_c_289_n N_VPWR_c_441_n 6.9093e-19 $X=2.66 $Y=2.085 $X2=0
+ $Y2=0
cc_227 N_A_137_419#_M1004_g N_VPWR_c_445_n 0.00924499f $X=3.775 $Y=2.595 $X2=0
+ $Y2=0
cc_228 N_A_137_419#_M1006_d N_VPWR_c_439_n 0.00225465f $X=0.685 $Y=2.095 $X2=0
+ $Y2=0
cc_229 N_A_137_419#_M1004_g N_VPWR_c_439_n 0.0182052f $X=3.775 $Y=2.595 $X2=0
+ $Y2=0
cc_230 N_A_137_419#_c_283_n X 0.00852269f $X=3.775 $Y=1.475 $X2=0 $Y2=0
cc_231 N_A_137_419#_M1004_g X 0.061748f $X=3.775 $Y=2.595 $X2=0 $Y2=0
cc_232 N_A_137_419#_c_290_n X 0.0135663f $X=3.355 $Y=1.285 $X2=0 $Y2=0
cc_233 N_A_137_419#_c_291_n X 0.0570295f $X=3.52 $Y=0.43 $X2=0 $Y2=0
cc_234 N_A_137_419#_c_293_n X 0.021256f $X=3.725 $Y=0.43 $X2=0 $Y2=0
cc_235 N_A_137_419#_c_285_n N_VGND_c_507_n 0.0117876f $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_236 N_A_137_419#_c_287_n N_VGND_c_507_n 0.00577797f $X=1.52 $Y=0.545 $X2=0
+ $Y2=0
cc_237 N_A_137_419#_c_286_n N_VGND_c_508_n 0.0139073f $X=2.575 $Y=0.545 $X2=0
+ $Y2=0
cc_238 N_A_137_419#_c_288_n N_VGND_c_508_n 0.0270818f $X=2.66 $Y=1.2 $X2=0 $Y2=0
cc_239 N_A_137_419#_c_290_n N_VGND_c_508_n 0.0196687f $X=3.355 $Y=1.285 $X2=0
+ $Y2=0
cc_240 N_A_137_419#_c_291_n N_VGND_c_508_n 0.0554984f $X=3.52 $Y=0.43 $X2=0
+ $Y2=0
cc_241 N_A_137_419#_c_293_n N_VGND_c_508_n 0.0127598f $X=3.725 $Y=0.43 $X2=0
+ $Y2=0
cc_242 N_A_137_419#_c_286_n N_VGND_c_509_n 0.0346907f $X=2.575 $Y=0.545 $X2=0
+ $Y2=0
cc_243 N_A_137_419#_c_287_n N_VGND_c_509_n 0.01008f $X=1.52 $Y=0.545 $X2=0 $Y2=0
cc_244 N_A_137_419#_c_291_n N_VGND_c_510_n 0.0209793f $X=3.52 $Y=0.43 $X2=0
+ $Y2=0
cc_245 N_A_137_419#_c_293_n N_VGND_c_510_n 0.0100081f $X=3.725 $Y=0.43 $X2=0
+ $Y2=0
cc_246 N_A_137_419#_c_286_n N_VGND_c_511_n 0.0402996f $X=2.575 $Y=0.545 $X2=0
+ $Y2=0
cc_247 N_A_137_419#_c_287_n N_VGND_c_511_n 0.0112907f $X=1.52 $Y=0.545 $X2=0
+ $Y2=0
cc_248 N_A_137_419#_c_291_n N_VGND_c_511_n 0.0124888f $X=3.52 $Y=0.43 $X2=0
+ $Y2=0
cc_249 N_A_137_419#_c_293_n N_VGND_c_511_n 0.00760165f $X=3.725 $Y=0.43 $X2=0
+ $Y2=0
cc_250 N_A_137_419#_c_288_n A_443_141# 0.00432633f $X=2.66 $Y=1.2 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_30_419#_c_404_n N_VPWR_M1007_d 0.00524772f $X=2.33 $Y=2.52 $X2=-0.19
+ $Y2=1.655
cc_252 N_A_30_419#_c_395_n N_VPWR_c_440_n 0.0119061f $X=1.19 $Y=2.98 $X2=0 $Y2=0
cc_253 N_A_30_419#_c_397_n N_VPWR_c_440_n 0.00721503f $X=1.355 $Y=2.75 $X2=0
+ $Y2=0
cc_254 N_A_30_419#_c_404_n N_VPWR_c_440_n 0.0199416f $X=2.33 $Y=2.52 $X2=0 $Y2=0
cc_255 N_A_30_419#_c_395_n N_VPWR_c_442_n 0.0575464f $X=1.19 $Y=2.98 $X2=0 $Y2=0
cc_256 N_A_30_419#_c_391_n N_VPWR_c_442_n 0.0198894f $X=0.46 $Y=2.98 $X2=0 $Y2=0
cc_257 N_A_30_419#_c_404_n N_VPWR_c_442_n 0.00265901f $X=2.33 $Y=2.52 $X2=0
+ $Y2=0
cc_258 N_A_30_419#_c_404_n N_VPWR_c_444_n 0.00341959f $X=2.33 $Y=2.52 $X2=0
+ $Y2=0
cc_259 N_A_30_419#_c_406_n N_VPWR_c_444_n 0.0177783f $X=2.495 $Y=2.75 $X2=0
+ $Y2=0
cc_260 N_A_30_419#_M1006_s N_VPWR_c_439_n 0.0023218f $X=0.15 $Y=2.095 $X2=0
+ $Y2=0
cc_261 N_A_30_419#_M1000_d N_VPWR_c_439_n 0.0022543f $X=1.215 $Y=2.095 $X2=0
+ $Y2=0
cc_262 N_A_30_419#_M1012_d N_VPWR_c_439_n 0.0022543f $X=2.355 $Y=2.095 $X2=0
+ $Y2=0
cc_263 N_A_30_419#_c_395_n N_VPWR_c_439_n 0.037727f $X=1.19 $Y=2.98 $X2=0 $Y2=0
cc_264 N_A_30_419#_c_391_n N_VPWR_c_439_n 0.0125808f $X=0.46 $Y=2.98 $X2=0 $Y2=0
cc_265 N_A_30_419#_c_404_n N_VPWR_c_439_n 0.0119638f $X=2.33 $Y=2.52 $X2=0 $Y2=0
cc_266 N_A_30_419#_c_406_n N_VPWR_c_439_n 0.0124439f $X=2.495 $Y=2.75 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_439_n N_X_M1004_d 0.0023218f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_c_441_n X 0.0282188f $X=3.09 $Y=2.24 $X2=0 $Y2=0
cc_269 N_VPWR_c_445_n X 0.0203976f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_270 N_VPWR_c_439_n X 0.0128489f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_271 X N_VGND_c_510_n 0.0110524f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_272 X N_VGND_c_511_n 0.0117849f $X=3.995 $Y=0.47 $X2=0 $Y2=0
