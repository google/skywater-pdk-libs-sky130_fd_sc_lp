* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 X a_112_65# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VPWR a_112_65# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_726_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_29_65# C1 a_112_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_292_367# B2 a_112_65# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR B1 a_292_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_284_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_112_65# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND A2 a_284_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 X a_112_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR C1 a_112_65# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_284_65# B2 a_29_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_112_65# B2 a_292_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_29_65# B2 a_284_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_284_65# B1 a_29_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VGND A1 a_284_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VPWR a_112_65# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 X a_112_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_284_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VGND a_112_65# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR A1 a_726_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_292_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_112_65# C1 a_29_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_29_65# B1 a_284_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_112_65# A2 a_726_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 X a_112_65# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_726_367# A2 a_112_65# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VGND a_112_65# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
