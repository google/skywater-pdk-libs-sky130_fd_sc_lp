* File: sky130_fd_sc_lp__and2b_lp.spice
* Created: Fri Aug 28 10:05:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2b_lp.pex.spice"
.subckt sky130_fd_sc_lp__and2b_lp  VNB VPB B A_N X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A_N	A_N
* B	B
* VPB	VPB
* VNB	VNB
MM1006 A_138_153# N_A_108_127#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_108_127#_M1003_g A_138_153# VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0504 PD=0.755 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 A_313_153# N_B_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.08225
+ AS=0.07035 PD=0.905 PS=0.755 NRD=40.236 NRS=15.708 M=1 R=2.8 SA=75001.1
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_108_127#_M1004_d N_A_378_159#_M1004_g A_313_153# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.08225 PD=1.41 PS=0.905 NRD=0 NRS=40.236 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_510_47# N_A_N_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_378_159#_M1007_d N_A_N_M1007_g A_510_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_108_127#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.25 W=1
+ AD=0.2425 AS=0.285 PD=1.485 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_108_127#_M1000_d N_B_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.2425 PD=1.28 PS=1.485 NRD=0 NRS=40.3653 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A_378_159#_M1009_g N_A_108_127#_M1000_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.2025 AS=0.14 PD=1.405 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1002 N_A_378_159#_M1002_d N_A_N_M1002_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.2025 PD=2.57 PS=1.405 NRD=0 NRS=24.6053 M=1 R=4 SA=125002
+ SB=125000 A=0.25 P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.937 P=11.27
*
.include "sky130_fd_sc_lp__and2b_lp.pxi.spice"
*
.ends
*
*
