* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__isolatch_lp D SLEEP_B KAPWR VGND VNB VPB VPWR Q
X0 a_419_73# a_458_293# a_521_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_21_179# SLEEP_B a_837_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_281_535# a_21_179# a_419_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_117_535# a_21_179# a_281_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_837_93# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_232_125# a_36_73# a_281_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 KAPWR a_281_535# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_36_73# a_21_179# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR D a_117_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 KAPWR a_21_179# a_36_73# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND D a_232_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_458_293# a_281_535# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_21_179# SLEEP_B KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_410_419# a_458_293# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 a_1284_177# a_281_535# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_281_535# a_36_73# a_410_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_1009_93# a_281_535# a_458_293# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_281_535# a_1284_177# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_521_73# a_458_293# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_281_535# a_1009_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
