* File: sky130_fd_sc_lp__nor3_m.spice
* Created: Wed Sep  2 10:09:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor3_m.pex.spice"
.subckt sky130_fd_sc_lp__nor3_m  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1 A=0.063
+ P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1000 A_123_483# N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.126 PD=0.66 PS=1.44 NRD=30.4759 NRS=16.4101 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1003 A_201_483# N_B_M1003_g A_123_483# VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=30.4759 NRS=30.4759 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_C_M1005_g A_201_483# VPB PHIGHVT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
c_181 A_123_483# 0 6.97414e-20 $X=0.615 $Y=2.415
*
.include "sky130_fd_sc_lp__nor3_m.pxi.spice"
*
.ends
*
*
