* File: sky130_fd_sc_lp__clkbuf_lp.pxi.spice
* Created: Fri Aug 28 10:15:16 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUF_LP%A_94_31# N_A_94_31#_M1003_d N_A_94_31#_M1001_d
+ N_A_94_31#_M1000_g N_A_94_31#_c_35_n N_A_94_31#_M1004_g N_A_94_31#_M1005_g
+ N_A_94_31#_c_37_n N_A_94_31#_c_41_n N_A_94_31#_c_42_n N_A_94_31#_c_43_n
+ N_A_94_31#_c_44_n N_A_94_31#_c_38_n PM_SKY130_FD_SC_LP__CLKBUF_LP%A_94_31#
x_PM_SKY130_FD_SC_LP__CLKBUF_LP%A N_A_c_89_n N_A_M1001_g N_A_c_90_n N_A_M1002_g
+ N_A_c_91_n N_A_M1003_g A A A PM_SKY130_FD_SC_LP__CLKBUF_LP%A
x_PM_SKY130_FD_SC_LP__CLKBUF_LP%X N_X_M1000_s N_X_M1004_s X X X X X X X
+ N_X_c_123_n X PM_SKY130_FD_SC_LP__CLKBUF_LP%X
x_PM_SKY130_FD_SC_LP__CLKBUF_LP%VPWR N_VPWR_M1004_d N_VPWR_c_143_n
+ N_VPWR_c_144_n N_VPWR_c_145_n VPWR N_VPWR_c_146_n N_VPWR_c_142_n
+ PM_SKY130_FD_SC_LP__CLKBUF_LP%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUF_LP%VGND N_VGND_M1005_d N_VGND_c_164_n VGND
+ N_VGND_c_165_n N_VGND_c_166_n N_VGND_c_167_n N_VGND_c_168_n
+ PM_SKY130_FD_SC_LP__CLKBUF_LP%VGND
cc_1 VNB N_A_94_31#_M1000_g 0.0402424f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.495
cc_2 VNB N_A_94_31#_c_35_n 0.0580216f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.835
cc_3 VNB N_A_94_31#_M1005_g 0.0357774f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.495
cc_4 VNB N_A_94_31#_c_37_n 0.0012441f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.33
cc_5 VNB N_A_94_31#_c_38_n 0.068013f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.495
cc_6 VNB N_A_c_89_n 0.0963502f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.285
cc_7 VNB N_A_c_90_n 0.0167868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_91_n 0.0182203f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.495
cc_9 VNB A 0.00224068f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.835
cc_10 VNB N_X_c_123_n 0.0653287f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=1.75
cc_11 VNB N_VPWR_c_142_n 0.103974f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=1.75
cc_12 VNB N_VGND_c_164_n 0.0141206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_165_n 0.0284206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_166_n 0.0331896f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.495
cc_15 VNB N_VGND_c_167_n 0.174162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_168_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.33
cc_17 VPB N_A_94_31#_c_35_n 0.0248541f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.835
cc_18 VPB N_A_94_31#_M1004_g 0.0354785f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.535
cc_19 VPB N_A_94_31#_c_41_n 0.0159709f $X=-0.19 $Y=1.655 $X2=1.535 $Y2=1.75
cc_20 VPB N_A_94_31#_c_42_n 0.00271353f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.75
cc_21 VPB N_A_94_31#_c_43_n 0.0501169f $X=-0.19 $Y=1.655 $X2=1.7 $Y2=2.18
cc_22 VPB N_A_94_31#_c_44_n 0.0283749f $X=-0.19 $Y=1.655 $X2=2.1 $Y2=1.665
cc_23 VPB N_A_94_31#_c_38_n 0.00128442f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.495
cc_24 VPB N_A_c_89_n 0.00168305f $X=-0.19 $Y=1.655 $X2=1.92 $Y2=0.285
cc_25 VPB N_A_M1001_g 0.0464991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB X 0.0374576f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.835
cc_27 VPB X 0.0190631f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.535
cc_28 VPB N_X_c_123_n 0.00946326f $X=-0.19 $Y=1.655 $X2=1.535 $Y2=1.75
cc_29 VPB N_VPWR_c_143_n 0.00675703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_144_n 0.0219971f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.835
cc_31 VPB N_VPWR_c_145_n 0.00556335f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.535
cc_32 VPB N_VPWR_c_146_n 0.0408627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_142_n 0.077677f $X=-0.19 $Y=1.655 $X2=1.535 $Y2=1.75
cc_34 N_A_94_31#_c_35_n N_A_c_89_n 0.0306391f $X=0.66 $Y=1.835 $X2=-0.19
+ $Y2=-0.245
cc_35 N_A_94_31#_c_37_n N_A_c_89_n 0.00261829f $X=0.905 $Y=1.33 $X2=-0.19
+ $Y2=-0.245
cc_36 N_A_94_31#_c_41_n N_A_c_89_n 0.00766318f $X=1.535 $Y=1.75 $X2=-0.19
+ $Y2=-0.245
cc_37 N_A_94_31#_c_44_n N_A_c_89_n 0.00749697f $X=2.1 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_38 N_A_94_31#_c_38_n N_A_c_89_n 0.0051575f $X=2.06 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_39 N_A_94_31#_M1004_g N_A_M1001_g 0.0160946f $X=0.66 $Y=2.535 $X2=0 $Y2=0
cc_40 N_A_94_31#_c_41_n N_A_M1001_g 0.0147045f $X=1.535 $Y=1.75 $X2=0 $Y2=0
cc_41 N_A_94_31#_c_43_n N_A_M1001_g 0.0332734f $X=1.7 $Y=2.18 $X2=0 $Y2=0
cc_42 N_A_94_31#_c_44_n N_A_M1001_g 0.00405169f $X=2.1 $Y=1.665 $X2=0 $Y2=0
cc_43 N_A_94_31#_M1005_g N_A_c_90_n 0.022004f $X=0.905 $Y=0.495 $X2=0 $Y2=0
cc_44 N_A_94_31#_c_38_n N_A_c_91_n 0.022913f $X=2.06 $Y=0.495 $X2=0 $Y2=0
cc_45 N_A_94_31#_c_35_n A 0.00133496f $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_46 N_A_94_31#_M1005_g A 0.00232976f $X=0.905 $Y=0.495 $X2=0 $Y2=0
cc_47 N_A_94_31#_c_37_n A 0.0121778f $X=0.905 $Y=1.33 $X2=0 $Y2=0
cc_48 N_A_94_31#_c_41_n A 0.0247098f $X=1.535 $Y=1.75 $X2=0 $Y2=0
cc_49 N_A_94_31#_c_38_n A 0.0672651f $X=2.06 $Y=0.495 $X2=0 $Y2=0
cc_50 N_A_94_31#_c_35_n X 0.00258773f $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_51 N_A_94_31#_M1004_g X 0.0241219f $X=0.66 $Y=2.535 $X2=0 $Y2=0
cc_52 N_A_94_31#_M1004_g X 0.00732788f $X=0.66 $Y=2.535 $X2=0 $Y2=0
cc_53 N_A_94_31#_M1000_g N_X_c_123_n 0.0258113f $X=0.545 $Y=0.495 $X2=0 $Y2=0
cc_54 N_A_94_31#_c_35_n N_X_c_123_n 0.0226459f $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_55 N_A_94_31#_M1005_g N_X_c_123_n 0.00344883f $X=0.905 $Y=0.495 $X2=0 $Y2=0
cc_56 N_A_94_31#_c_37_n N_X_c_123_n 0.0297326f $X=0.905 $Y=1.33 $X2=0 $Y2=0
cc_57 N_A_94_31#_c_42_n N_X_c_123_n 0.0108953f $X=1.07 $Y=1.75 $X2=0 $Y2=0
cc_58 N_A_94_31#_c_35_n N_VPWR_c_143_n 0.00221364f $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_59 N_A_94_31#_M1004_g N_VPWR_c_143_n 0.0244058f $X=0.66 $Y=2.535 $X2=0 $Y2=0
cc_60 N_A_94_31#_c_41_n N_VPWR_c_143_n 0.00150469f $X=1.535 $Y=1.75 $X2=0 $Y2=0
cc_61 N_A_94_31#_c_42_n N_VPWR_c_143_n 0.0262399f $X=1.07 $Y=1.75 $X2=0 $Y2=0
cc_62 N_A_94_31#_c_43_n N_VPWR_c_143_n 0.0384439f $X=1.7 $Y=2.18 $X2=0 $Y2=0
cc_63 N_A_94_31#_M1004_g N_VPWR_c_144_n 0.00754485f $X=0.66 $Y=2.535 $X2=0 $Y2=0
cc_64 N_A_94_31#_c_43_n N_VPWR_c_146_n 0.020789f $X=1.7 $Y=2.18 $X2=0 $Y2=0
cc_65 N_A_94_31#_M1004_g N_VPWR_c_142_n 0.0139836f $X=0.66 $Y=2.535 $X2=0 $Y2=0
cc_66 N_A_94_31#_c_43_n N_VPWR_c_142_n 0.0125177f $X=1.7 $Y=2.18 $X2=0 $Y2=0
cc_67 N_A_94_31#_M1000_g N_VGND_c_164_n 0.002112f $X=0.545 $Y=0.495 $X2=0 $Y2=0
cc_68 N_A_94_31#_c_35_n N_VGND_c_164_n 6.10645e-19 $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_69 N_A_94_31#_M1005_g N_VGND_c_164_n 0.0130921f $X=0.905 $Y=0.495 $X2=0 $Y2=0
cc_70 N_A_94_31#_c_37_n N_VGND_c_164_n 0.00481421f $X=0.905 $Y=1.33 $X2=0 $Y2=0
cc_71 N_A_94_31#_M1000_g N_VGND_c_165_n 0.00502664f $X=0.545 $Y=0.495 $X2=0
+ $Y2=0
cc_72 N_A_94_31#_M1005_g N_VGND_c_165_n 0.00445056f $X=0.905 $Y=0.495 $X2=0
+ $Y2=0
cc_73 N_A_94_31#_c_38_n N_VGND_c_166_n 0.0167213f $X=2.06 $Y=0.495 $X2=0 $Y2=0
cc_74 N_A_94_31#_M1000_g N_VGND_c_167_n 0.0100902f $X=0.545 $Y=0.495 $X2=0 $Y2=0
cc_75 N_A_94_31#_M1005_g N_VGND_c_167_n 0.00796275f $X=0.905 $Y=0.495 $X2=0
+ $Y2=0
cc_76 N_A_94_31#_c_38_n N_VGND_c_167_n 0.0095959f $X=2.06 $Y=0.495 $X2=0 $Y2=0
cc_77 N_A_M1001_g N_VPWR_c_143_n 0.0139346f $X=1.435 $Y=2.535 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_VPWR_c_146_n 0.00845216f $X=1.435 $Y=2.535 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_VPWR_c_142_n 0.0167829f $X=1.435 $Y=2.535 $X2=0 $Y2=0
cc_80 N_A_c_90_n N_VGND_c_164_n 0.00934749f $X=1.485 $Y=0.815 $X2=0 $Y2=0
cc_81 A N_VGND_c_164_n 0.0211991f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_82 N_A_c_90_n N_VGND_c_166_n 0.00423858f $X=1.485 $Y=0.815 $X2=0 $Y2=0
cc_83 N_A_c_91_n N_VGND_c_166_n 0.00507383f $X=1.845 $Y=0.815 $X2=0 $Y2=0
cc_84 A N_VGND_c_166_n 0.00851294f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A_c_90_n N_VGND_c_167_n 0.00716149f $X=1.485 $Y=0.815 $X2=0 $Y2=0
cc_86 N_A_c_91_n N_VGND_c_167_n 0.0101244f $X=1.845 $Y=0.815 $X2=0 $Y2=0
cc_87 A N_VGND_c_167_n 0.0108483f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_88 A A_312_57# 0.00133334f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_89 X N_VPWR_c_143_n 0.0442231f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_90 X N_VPWR_c_143_n 0.0255914f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_91 X N_VPWR_c_144_n 0.0243021f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_92 X N_VPWR_c_142_n 0.016239f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_93 N_X_c_123_n N_VGND_c_164_n 0.0155263f $X=0.33 $Y=0.495 $X2=0 $Y2=0
cc_94 N_X_c_123_n N_VGND_c_165_n 0.0247291f $X=0.33 $Y=0.495 $X2=0 $Y2=0
cc_95 N_X_c_123_n N_VGND_c_167_n 0.0141285f $X=0.33 $Y=0.495 $X2=0 $Y2=0
