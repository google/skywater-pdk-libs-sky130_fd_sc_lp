* File: sky130_fd_sc_lp__invkapwr_2.pex.spice
* Created: Fri Aug 28 10:39:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVKAPWR_2%A 3 7 11 15 19 21 22 33 34
r48 34 35 11.5066 $w=3.77e-07 $l=9e-08 $layer=POLY_cond $X=1.355 $Y=1.485
+ $X2=1.445 $Y2=1.485
r49 32 34 12.1459 $w=3.77e-07 $l=9.5e-08 $layer=POLY_cond $X=1.26 $Y=1.485
+ $X2=1.355 $Y2=1.485
r50 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=1.46 $X2=1.26 $Y2=1.46
r51 30 32 31.3236 $w=3.77e-07 $l=2.45e-07 $layer=POLY_cond $X=1.015 $Y=1.485
+ $X2=1.26 $Y2=1.485
r52 29 30 11.5066 $w=3.77e-07 $l=9e-08 $layer=POLY_cond $X=0.925 $Y=1.485
+ $X2=1.015 $Y2=1.485
r53 27 29 0.639257 $w=3.77e-07 $l=5e-09 $layer=POLY_cond $X=0.92 $Y=1.485
+ $X2=0.925 $Y2=1.485
r54 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.46 $X2=0.92 $Y2=1.46
r55 25 27 54.3369 $w=3.77e-07 $l=4.25e-07 $layer=POLY_cond $X=0.495 $Y=1.485
+ $X2=0.92 $Y2=1.485
r56 22 33 2.06408 $w=3.33e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=1.377 $X2=1.26
+ $Y2=1.377
r57 22 28 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=1.2 $Y=1.377
+ $X2=0.92 $Y2=1.377
r58 21 28 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=0.72 $Y=1.377 $X2=0.92
+ $Y2=1.377
r59 17 35 24.4204 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.445 $Y=1.295
+ $X2=1.445 $Y2=1.485
r60 17 19 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.445 $Y=1.295
+ $X2=1.445 $Y2=0.56
r61 13 34 24.4204 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.355 $Y=1.675
+ $X2=1.355 $Y2=1.485
r62 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.355 $Y=1.675
+ $X2=1.355 $Y2=2.465
r63 9 30 24.4204 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.015 $Y=1.295
+ $X2=1.015 $Y2=1.485
r64 9 11 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.015 $Y=1.295
+ $X2=1.015 $Y2=0.56
r65 5 29 24.4204 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.925 $Y=1.675
+ $X2=0.925 $Y2=1.485
r66 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.925 $Y=1.675
+ $X2=0.925 $Y2=2.465
r67 1 25 24.4204 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.675
+ $X2=0.495 $Y2=1.485
r68 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.495 $Y=1.675
+ $X2=0.495 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_2%Y 1 2 3 12 16 17 20 26 28 30 31 33 34 38
r55 34 38 15.2875 $w=1.83e-07 $l=2.55e-07 $layer=LI1_cond $X=1.687 $Y=1.295
+ $X2=1.687 $Y2=1.04
r56 33 38 3.55727 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=1.687 $Y=0.94
+ $X2=1.687 $Y2=1.04
r57 32 34 25.1794 $w=1.83e-07 $l=4.2e-07 $layer=LI1_cond $X=1.687 $Y=1.715
+ $X2=1.687 $Y2=1.295
r58 31 33 9.73502 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.325 $Y=0.94
+ $X2=1.595 $Y2=0.94
r59 29 30 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.27 $Y=1.8 $X2=1.14
+ $Y2=1.8
r60 28 32 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=1.595 $Y=1.8
+ $X2=1.687 $Y2=1.715
r61 28 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.595 $Y=1.8
+ $X2=1.27 $Y2=1.8
r62 24 31 6.84722 $w=2e-07 $l=1.55142e-07 $layer=LI1_cond $X=1.212 $Y=0.84
+ $X2=1.325 $Y2=0.94
r63 24 26 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=1.212 $Y=0.84
+ $X2=1.212 $Y2=0.56
r64 20 22 39.0058 $w=2.58e-07 $l=8.8e-07 $layer=LI1_cond $X=1.14 $Y=2 $X2=1.14
+ $Y2=2.88
r65 18 30 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.885
+ $X2=1.14 $Y2=1.8
r66 18 20 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.14 $Y=1.885
+ $X2=1.14 $Y2=2
r67 16 30 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.01 $Y=1.8 $X2=1.14
+ $Y2=1.8
r68 16 17 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.01 $Y=1.8 $X2=0.41
+ $Y2=1.8
r69 12 14 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=0.282 $Y=2 $X2=0.282
+ $Y2=2.88
r70 10 17 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.282 $Y=1.885
+ $X2=0.41 $Y2=1.8
r71 10 12 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=0.282 $Y=1.885
+ $X2=0.282 $Y2=2
r72 3 22 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=1 $Y=1.835
+ $X2=1.14 $Y2=2.88
r73 3 20 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2
r74 2 14 400 $w=1.7e-07 $l=1.10574e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=2.88
r75 2 12 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=2
r76 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.35 $X2=1.23 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_2%KAPWR 1 2 7 10 18 22 28
r23 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.565 $Y=2.81
+ $X2=1.565 $Y2=2.81
r24 18 21 26.6644 $w=2.53e-07 $l=5.9e-07 $layer=LI1_cond $X=1.567 $Y=2.22
+ $X2=1.567 $Y2=2.81
r25 14 28 0.141782 $w=2.55e-07 $l=2.45e-07 $layer=MET1_cond $X=0.705 $Y=2.817
+ $X2=0.95 $Y2=2.817
r26 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.705 $Y=2.81
+ $X2=0.705 $Y2=2.81
r27 10 13 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=0.71 $Y=2.22
+ $X2=0.71 $Y2=2.81
r28 7 22 0.350115 $w=2.55e-07 $l=6.05e-07 $layer=MET1_cond $X=0.96 $Y=2.817
+ $X2=1.565 $Y2=2.817
r29 7 28 0.00578702 $w=2.55e-07 $l=1e-08 $layer=MET1_cond $X=0.96 $Y=2.817
+ $X2=0.95 $Y2=2.817
r30 2 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.91
r31 2 18 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.22
r32 1 13 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.91
r33 1 10 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_2%VGND 1 2 9 11 13 15 17 22 28 32
r22 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r23 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r24 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r25 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r26 23 28 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.782
+ $Y2=0
r27 23 25 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.2
+ $Y2=0
r28 22 31 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.707
+ $Y2=0
r29 22 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.2
+ $Y2=0
r30 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r31 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r32 17 28 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.782
+ $Y2=0
r33 17 19 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.24
+ $Y2=0
r34 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r35 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r36 11 31 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.707 $Y2=0
r37 11 13 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0.56
r38 7 28 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=0.085
+ $X2=0.782 $Y2=0
r39 7 9 18.5563 $w=2.93e-07 $l=4.75e-07 $layer=LI1_cond $X=0.782 $Y=0.085
+ $X2=0.782 $Y2=0.56
r40 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.35 $X2=1.66 $Y2=0.56
r41 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.675
+ $Y=0.35 $X2=0.8 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_2%VPWR 1 8 14
r23 5 14 0.0081048 $w=1.92e-06 $l=1.22e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.96 $Y2=3.208
r24 5 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33 $X2=1.68
+ $Y2=3.33
r25 4 8 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.68
+ $Y2=3.33
r26 4 5 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r27 1 14 6.64328e-05 $w=1.92e-06 $l=1e-09 $layer=MET1_cond $X=0.96 $Y=3.207
+ $X2=0.96 $Y2=3.208
.ends

