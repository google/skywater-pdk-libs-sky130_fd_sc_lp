# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.210000 1.850000 1.515000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.020000 1.210000 5.330000 1.245000 ;
        RECT 2.020000 1.245000 3.250000 1.515000 ;
        RECT 3.035000 1.075000 5.330000 1.210000 ;
        RECT 5.070000 1.245000 5.330000 1.515000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.420000 1.415000 4.770000 1.645000 ;
        RECT 3.420000 1.645000 4.235000 1.765000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  2.116800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 0.255000 0.795000 0.870000 ;
        RECT 0.575000 0.870000 5.670000 0.895000 ;
        RECT 0.575000 0.895000 2.865000 1.040000 ;
        RECT 1.465000 0.255000 1.655000 0.870000 ;
        RECT 2.325000 0.255000 2.545000 0.725000 ;
        RECT 2.325000 0.725000 5.670000 0.870000 ;
        RECT 3.115000 0.255000 3.445000 0.725000 ;
        RECT 3.545000 1.935000 5.670000 1.985000 ;
        RECT 3.545000 1.985000 4.735000 2.155000 ;
        RECT 3.975000 0.255000 4.305000 0.725000 ;
        RECT 4.405000 1.815000 5.670000 1.935000 ;
        RECT 4.835000 0.255000 5.165000 0.725000 ;
        RECT 5.500000 0.895000 5.670000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.105000  0.085000 0.405000 1.040000 ;
      RECT 0.105000  1.705000 3.015000 1.875000 ;
      RECT 0.105000  1.875000 0.365000 3.075000 ;
      RECT 0.535000  2.105000 0.865000 3.245000 ;
      RECT 0.965000  0.085000 1.295000 0.700000 ;
      RECT 1.035000  1.875000 1.225000 3.075000 ;
      RECT 1.395000  2.105000 1.725000 3.245000 ;
      RECT 1.825000  0.085000 2.155000 0.700000 ;
      RECT 1.895000  1.875000 2.085000 3.075000 ;
      RECT 2.255000  2.055000 2.585000 2.675000 ;
      RECT 2.255000  2.675000 5.105000 3.075000 ;
      RECT 2.715000  0.085000 2.945000 0.555000 ;
      RECT 2.755000  1.875000 3.015000 2.325000 ;
      RECT 2.755000  2.325000 5.615000 2.495000 ;
      RECT 3.615000  0.085000 3.805000 0.555000 ;
      RECT 4.475000  0.085000 4.665000 0.555000 ;
      RECT 5.285000  2.155000 5.615000 2.325000 ;
      RECT 5.285000  2.495000 5.615000 3.075000 ;
      RECT 5.335000  0.085000 5.595000 0.555000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__nor3_4
END LIBRARY
