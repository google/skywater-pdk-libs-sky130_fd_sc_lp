* File: sky130_fd_sc_lp__fa_m.pxi.spice
* Created: Wed Sep  2 09:53:36 2020
* 
x_PM_SKY130_FD_SC_LP__FA_M%A_80_241# N_A_80_241#_M1007_d N_A_80_241#_M1005_d
+ N_A_80_241#_M1024_g N_A_80_241#_M1021_g N_A_80_241#_M1027_g
+ N_A_80_241#_M1016_g N_A_80_241#_c_143_n N_A_80_241#_c_154_p
+ N_A_80_241#_c_144_n N_A_80_241#_c_145_n N_A_80_241#_c_146_n
+ N_A_80_241#_c_147_n N_A_80_241#_c_148_n N_A_80_241#_c_149_n
+ PM_SKY130_FD_SC_LP__FA_M%A_80_241#
x_PM_SKY130_FD_SC_LP__FA_M%B N_B_M1007_g N_B_M1005_g N_B_M1009_g N_B_c_244_n
+ N_B_M1004_g N_B_c_236_n N_B_c_237_n N_B_M1023_g N_B_M1006_g N_B_M1022_g
+ N_B_M1015_g N_B_c_240_n N_B_c_241_n N_B_c_242_n N_B_c_252_n N_B_c_253_n
+ N_B_c_254_n N_B_c_255_n N_B_c_256_n N_B_c_257_n B B B N_B_c_258_n N_B_c_259_n
+ N_B_c_260_n N_B_c_261_n N_B_c_262_n PM_SKY130_FD_SC_LP__FA_M%B
x_PM_SKY130_FD_SC_LP__FA_M%CIN N_CIN_M1008_g N_CIN_M1025_g N_CIN_c_380_n
+ N_CIN_c_381_n N_CIN_M1017_g N_CIN_M1014_g N_CIN_c_383_n N_CIN_M1000_g
+ N_CIN_M1011_g N_CIN_c_385_n N_CIN_c_386_n CIN N_CIN_c_387_n N_CIN_c_388_n
+ PM_SKY130_FD_SC_LP__FA_M%CIN
x_PM_SKY130_FD_SC_LP__FA_M%A N_A_M1013_g N_A_M1002_g N_A_c_452_n N_A_c_453_n
+ N_A_M1010_g N_A_M1026_g N_A_c_456_n N_A_M1018_g N_A_M1003_g N_A_c_458_n
+ N_A_M1012_g N_A_M1020_g N_A_c_460_n N_A_c_461_n A A A N_A_c_463_n N_A_c_464_n
+ PM_SKY130_FD_SC_LP__FA_M%A
x_PM_SKY130_FD_SC_LP__FA_M%A_1101_119# N_A_1101_119#_M1027_d
+ N_A_1101_119#_M1016_d N_A_1101_119#_c_569_n N_A_1101_119#_M1019_g
+ N_A_1101_119#_M1001_g N_A_1101_119#_c_570_n N_A_1101_119#_c_571_n
+ N_A_1101_119#_c_572_n N_A_1101_119#_c_573_n N_A_1101_119#_c_580_n
+ N_A_1101_119#_c_574_n N_A_1101_119#_c_575_n N_A_1101_119#_c_576_n
+ PM_SKY130_FD_SC_LP__FA_M%A_1101_119#
x_PM_SKY130_FD_SC_LP__FA_M%COUT N_COUT_M1021_s N_COUT_M1024_s N_COUT_c_627_n
+ COUT COUT COUT COUT COUT PM_SKY130_FD_SC_LP__FA_M%COUT
x_PM_SKY130_FD_SC_LP__FA_M%VPWR N_VPWR_M1024_d N_VPWR_M1010_d N_VPWR_M1006_s
+ N_VPWR_M1014_d N_VPWR_M1020_d N_VPWR_c_640_n N_VPWR_c_641_n N_VPWR_c_642_n
+ N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n N_VPWR_c_646_n N_VPWR_c_647_n
+ N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n N_VPWR_c_651_n VPWR
+ N_VPWR_c_652_n N_VPWR_c_653_n N_VPWR_c_639_n N_VPWR_c_655_n
+ PM_SKY130_FD_SC_LP__FA_M%VPWR
x_PM_SKY130_FD_SC_LP__FA_M%A_385_367# N_A_385_367#_M1025_d N_A_385_367#_M1004_d
+ N_A_385_367#_c_740_n N_A_385_367#_c_741_n N_A_385_367#_c_742_n
+ PM_SKY130_FD_SC_LP__FA_M%A_385_367#
x_PM_SKY130_FD_SC_LP__FA_M%A_843_391# N_A_843_391#_M1006_d N_A_843_391#_M1003_d
+ N_A_843_391#_c_761_n N_A_843_391#_c_762_n N_A_843_391#_c_763_n
+ N_A_843_391#_c_764_n PM_SKY130_FD_SC_LP__FA_M%A_843_391#
x_PM_SKY130_FD_SC_LP__FA_M%SUM N_SUM_M1019_d N_SUM_M1001_d N_SUM_c_784_n SUM SUM
+ SUM SUM SUM PM_SKY130_FD_SC_LP__FA_M%SUM
x_PM_SKY130_FD_SC_LP__FA_M%VGND N_VGND_M1021_d N_VGND_M1026_d N_VGND_M1023_s
+ N_VGND_M1017_d N_VGND_M1012_d N_VGND_c_798_n N_VGND_c_799_n N_VGND_c_800_n
+ N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n N_VGND_c_804_n N_VGND_c_844_n
+ N_VGND_c_805_n N_VGND_c_806_n N_VGND_c_807_n N_VGND_c_808_n N_VGND_c_809_n
+ N_VGND_c_810_n N_VGND_c_811_n N_VGND_c_812_n VGND N_VGND_c_813_n
+ N_VGND_c_814_n PM_SKY130_FD_SC_LP__FA_M%VGND
x_PM_SKY130_FD_SC_LP__FA_M%A_385_125# N_A_385_125#_M1008_d N_A_385_125#_M1009_d
+ N_A_385_125#_c_883_n N_A_385_125#_c_898_n N_A_385_125#_c_884_n
+ PM_SKY130_FD_SC_LP__FA_M%A_385_125#
x_PM_SKY130_FD_SC_LP__FA_M%A_843_119# N_A_843_119#_M1023_d N_A_843_119#_M1018_d
+ N_A_843_119#_c_917_n N_A_843_119#_c_909_n N_A_843_119#_c_910_n
+ N_A_843_119#_c_919_n PM_SKY130_FD_SC_LP__FA_M%A_843_119#
cc_1 VNB N_A_80_241#_M1024_g 0.00734606f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.045
cc_2 VNB N_A_80_241#_M1021_g 0.0245049f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.835
cc_3 VNB N_A_80_241#_M1027_g 0.0246727f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=0.805
cc_4 VNB N_A_80_241#_M1016_g 0.00216594f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=2.165
cc_5 VNB N_A_80_241#_c_143_n 0.0240334f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.45
cc_6 VNB N_A_80_241#_c_144_n 0.00220909f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.98
cc_7 VNB N_A_80_241#_c_145_n 0.0607362f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_8 VNB N_A_80_241#_c_146_n 0.0350534f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_9 VNB N_A_80_241#_c_147_n 0.00313074f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.37
cc_10 VNB N_A_80_241#_c_148_n 0.0388327f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.37
cc_11 VNB N_A_80_241#_c_149_n 0.002861f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.45
cc_12 VNB N_B_M1007_g 0.0342438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_M1009_g 0.0484172f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.045
cc_14 VNB N_B_c_236_n 0.00999198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_237_n 0.0214962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1023_g 0.0472233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_M1022_g 0.0378152f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.98
cc_18 VNB N_B_c_240_n 0.00338523f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_19 VNB N_B_c_241_n 0.00584094f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_20 VNB N_B_c_242_n 0.0049077f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_21 VNB N_CIN_M1008_g 0.0369557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_CIN_M1017_g 0.0395333f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.205
cc_23 VNB N_CIN_M1000_g 0.0370182f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=1.615
cc_24 VNB N_A_M1013_g 0.0506834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_c_452_n 0.0679716f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.535
cc_26 VNB N_A_c_453_n 0.012503f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.045
cc_27 VNB N_A_M1010_g 0.0177401f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.205
cc_28 VNB N_A_M1026_g 0.0121865f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=0.805
cc_29 VNB N_A_c_456_n 0.189096f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=0.805
cc_30 VNB N_A_M1018_g 0.0553337f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=2.165
cc_31 VNB N_A_c_458_n 0.124501f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.365
cc_32 VNB N_A_M1012_g 0.053511f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.535
cc_33 VNB N_A_c_460_n 0.0137598f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_34 VNB N_A_c_461_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB A 0.00354893f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.37
cc_36 VNB N_A_c_463_n 0.0451035f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.37
cc_37 VNB N_A_c_464_n 0.00569926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1101_119#_c_569_n 0.0235065f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=2.045
cc_39 VNB N_A_1101_119#_c_570_n 0.00375784f $X=-0.19 $Y=-0.245 $X2=5.43
+ $Y2=0.805
cc_40 VNB N_A_1101_119#_c_571_n 0.00997374f $X=-0.19 $Y=-0.245 $X2=5.43
+ $Y2=0.805
cc_41 VNB N_A_1101_119#_c_572_n 0.00291173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1101_119#_c_573_n 0.0390569f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=1.615
cc_43 VNB N_A_1101_119#_c_574_n 2.7762e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1101_119#_c_575_n 0.0214163f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.45
cc_45 VNB N_A_1101_119#_c_576_n 0.0215052f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_46 VNB N_COUT_c_627_n 0.0162969f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.205
cc_47 VNB COUT 0.0313128f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.835
cc_48 VNB N_VPWR_c_639_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_SUM_c_784_n 0.0113784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB SUM 0.034122f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.835
cc_51 VNB N_VGND_c_798_n 0.0200314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_799_n 0.0137671f $X=-0.19 $Y=-0.245 $X2=5.43 $Y2=2.165
cc_53 VNB N_VGND_c_800_n 0.0176069f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.45
cc_54 VNB N_VGND_c_801_n 0.00335285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_802_n 0.0196633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_803_n 0.0242526f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_57 VNB N_VGND_c_804_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_58 VNB N_VGND_c_805_n 0.041006f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.45
cc_59 VNB N_VGND_c_806_n 0.00226387f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.37
cc_60 VNB N_VGND_c_807_n 0.0281107f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.535
cc_61 VNB N_VGND_c_808_n 0.00279655f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.45
cc_62 VNB N_VGND_c_809_n 0.0158898f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.615
cc_63 VNB N_VGND_c_810_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_811_n 0.053314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_812_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_813_n 0.0247812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_814_n 0.395816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_385_125#_c_883_n 0.0123698f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.535
cc_69 VNB N_A_385_125#_c_884_n 0.00316673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_843_119#_c_909_n 0.00711356f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.205
cc_71 VNB N_A_843_119#_c_910_n 0.00391136f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.835
cc_72 VPB N_A_80_241#_M1024_g 0.0259917f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.045
cc_73 VPB N_A_80_241#_M1016_g 0.0261038f $X=-0.19 $Y=1.655 $X2=5.43 $Y2=2.165
cc_74 VPB N_A_80_241#_c_144_n 0.00388096f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.98
cc_75 VPB N_B_M1007_g 0.0298134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_B_c_244_n 0.0178768f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.205
cc_77 VPB N_B_c_236_n 0.00596434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_B_c_237_n 0.0112931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_B_M1006_g 0.0281561f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=0.92
cc_80 VPB N_B_M1022_g 0.0337962f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.98
cc_81 VPB N_B_c_240_n 0.00309079f $X=-0.19 $Y=1.655 $X2=5.45 $Y2=1.45
cc_82 VPB N_B_c_241_n 8.27806e-19 $X=-0.19 $Y=1.655 $X2=5.45 $Y2=1.45
cc_83 VPB N_B_c_242_n 3.59711e-19 $X=-0.19 $Y=1.655 $X2=5.45 $Y2=1.45
cc_84 VPB N_B_c_252_n 0.00118164f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.37
cc_85 VPB N_B_c_253_n 0.0130629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_B_c_254_n 0.00961713f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.45
cc_87 VPB N_B_c_255_n 0.0440461f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.535
cc_88 VPB N_B_c_256_n 0.0376816f $X=-0.19 $Y=1.655 $X2=5.45 $Y2=1.45
cc_89 VPB N_B_c_257_n 0.0160719f $X=-0.19 $Y=1.655 $X2=5.45 $Y2=1.615
cc_90 VPB N_B_c_258_n 0.0462783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_B_c_259_n 0.0400087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_B_c_260_n 0.0565122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_B_c_261_n 0.0325454f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_B_c_262_n 0.00949182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_CIN_M1008_g 0.0363596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_CIN_c_380_n 0.171336f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.535
cc_97 VPB N_CIN_c_381_n 0.0217847f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.045
cc_98 VPB N_CIN_M1017_g 0.0734958f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.205
cc_99 VPB N_CIN_c_383_n 0.0944918f $X=-0.19 $Y=1.655 $X2=5.43 $Y2=1.285
cc_100 VPB N_CIN_M1000_g 0.0588957f $X=-0.19 $Y=1.655 $X2=5.43 $Y2=1.615
cc_101 VPB N_CIN_c_385_n 0.0164403f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.365
cc_102 VPB N_CIN_c_386_n 0.00749069f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=0.92
cc_103 VPB N_CIN_c_387_n 0.0162535f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.98
cc_104 VPB N_CIN_c_388_n 0.00924407f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.98
cc_105 VPB N_A_M1013_g 0.0233289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_M1010_g 0.0227755f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.205
cc_107 VPB N_A_M1018_g 0.0236011f $X=-0.19 $Y=1.655 $X2=5.43 $Y2=2.165
cc_108 VPB N_A_M1012_g 0.0262193f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.535
cc_109 VPB N_A_1101_119#_M1001_g 0.0240902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_1101_119#_c_570_n 0.0176536f $X=-0.19 $Y=1.655 $X2=5.43 $Y2=0.805
cc_111 VPB N_A_1101_119#_c_572_n 0.00256849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_1101_119#_c_580_n 0.00748839f $X=-0.19 $Y=1.655 $X2=1.635
+ $Y2=1.535
cc_113 VPB N_A_1101_119#_c_574_n 0.00548423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB COUT 0.0416298f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.835
cc_115 VPB N_VPWR_c_640_n 0.0371476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_641_n 0.019653f $X=-0.19 $Y=1.655 $X2=5.43 $Y2=2.165
cc_117 VPB N_VPWR_c_642_n 0.00883768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_643_n 8.47464e-19 $X=-0.19 $Y=1.655 $X2=1.635 $Y2=0.92
cc_119 VPB N_VPWR_c_644_n 0.0357885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_645_n 0.0241889f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.98
cc_121 VPB N_VPWR_c_646_n 0.0063612f $X=-0.19 $Y=1.655 $X2=1.8 $Y2=1.45
cc_122 VPB N_VPWR_c_647_n 0.00443729f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.37
cc_123 VPB N_VPWR_c_648_n 0.00164942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_649_n 0.00533485f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.45
cc_125 VPB N_VPWR_c_650_n 0.148335f $X=-0.19 $Y=1.655 $X2=5.45 $Y2=1.285
cc_126 VPB N_VPWR_c_651_n 0.00324402f $X=-0.19 $Y=1.655 $X2=5.45 $Y2=1.615
cc_127 VPB N_VPWR_c_652_n 0.0176897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_653_n 0.0226221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_639_n 0.0953278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_655_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_385_367#_c_740_n 0.00598165f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=1.535
cc_132 VPB N_A_385_367#_c_741_n 0.00322664f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=2.045
cc_133 VPB N_A_385_367#_c_742_n 0.00224547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_843_391#_c_761_n 0.00136805f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=2.045
cc_135 VPB N_A_843_391#_c_762_n 0.011008f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.205
cc_136 VPB N_A_843_391#_c_763_n 0.00421427f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.835
cc_137 VPB N_A_843_391#_c_764_n 0.00123105f $X=-0.19 $Y=1.655 $X2=5.43 $Y2=1.285
cc_138 VPB SUM 0.04226f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.835
cc_139 N_A_80_241#_c_143_n N_B_M1007_g 0.0144354f $X=1.47 $Y=1.45 $X2=0 $Y2=0
cc_140 N_A_80_241#_c_154_p N_B_M1007_g 0.0132254f $X=1.635 $Y=0.92 $X2=0 $Y2=0
cc_141 N_A_80_241#_c_144_n N_B_M1007_g 0.0076035f $X=1.635 $Y=1.98 $X2=0 $Y2=0
cc_142 N_A_80_241#_c_149_n N_B_M1007_g 0.00363367f $X=1.635 $Y=1.45 $X2=0 $Y2=0
cc_143 N_A_80_241#_c_145_n N_B_M1009_g 0.0104138f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_144 N_A_80_241#_c_145_n N_B_c_236_n 0.0116888f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_145 N_A_80_241#_c_145_n N_B_c_237_n 0.0267887f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_146 N_A_80_241#_c_145_n N_B_M1023_g 0.0140169f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_147 N_A_80_241#_c_145_n N_B_c_240_n 0.00273107f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_148 N_A_80_241#_c_145_n N_B_c_241_n 0.009504f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_149 N_A_80_241#_c_145_n N_B_c_242_n 0.00713f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_150 N_A_80_241#_c_144_n N_B_c_253_n 0.0138628f $X=1.635 $Y=1.98 $X2=0 $Y2=0
cc_151 N_A_80_241#_M1016_g N_B_c_255_n 4.80386e-19 $X=5.43 $Y=2.165 $X2=0 $Y2=0
cc_152 N_A_80_241#_c_154_p N_CIN_M1008_g 0.0110062f $X=1.635 $Y=0.92 $X2=0 $Y2=0
cc_153 N_A_80_241#_c_144_n N_CIN_M1008_g 0.00555026f $X=1.635 $Y=1.98 $X2=0
+ $Y2=0
cc_154 N_A_80_241#_c_145_n N_CIN_M1008_g 0.0148906f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_155 N_A_80_241#_c_149_n N_CIN_M1008_g 0.00363367f $X=1.635 $Y=1.45 $X2=0
+ $Y2=0
cc_156 N_A_80_241#_c_145_n N_CIN_M1017_g 0.0105827f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_157 N_A_80_241#_M1016_g N_CIN_c_383_n 0.00201695f $X=5.43 $Y=2.165 $X2=0
+ $Y2=0
cc_158 N_A_80_241#_M1027_g N_CIN_M1000_g 0.0188072f $X=5.43 $Y=0.805 $X2=0 $Y2=0
cc_159 N_A_80_241#_M1016_g N_CIN_M1000_g 0.0215643f $X=5.43 $Y=2.165 $X2=0 $Y2=0
cc_160 N_A_80_241#_c_146_n N_CIN_M1000_g 0.0209578f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_161 N_A_80_241#_M1024_g N_A_M1013_g 0.0174292f $X=0.475 $Y=2.045 $X2=0 $Y2=0
cc_162 N_A_80_241#_M1021_g N_A_M1013_g 0.0158568f $X=0.63 $Y=0.835 $X2=0 $Y2=0
cc_163 N_A_80_241#_c_143_n N_A_M1013_g 0.0186515f $X=1.47 $Y=1.45 $X2=0 $Y2=0
cc_164 N_A_80_241#_c_154_p N_A_M1013_g 0.00243786f $X=1.635 $Y=0.92 $X2=0 $Y2=0
cc_165 N_A_80_241#_c_147_n N_A_M1013_g 9.79826e-19 $X=0.61 $Y=1.37 $X2=0 $Y2=0
cc_166 N_A_80_241#_c_148_n N_A_M1013_g 0.0211904f $X=0.61 $Y=1.37 $X2=0 $Y2=0
cc_167 N_A_80_241#_c_145_n N_A_M1010_g 0.0115445f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_168 N_A_80_241#_M1027_g N_A_M1018_g 0.0215351f $X=5.43 $Y=0.805 $X2=0 $Y2=0
cc_169 N_A_80_241#_M1016_g N_A_M1018_g 0.0248243f $X=5.43 $Y=2.165 $X2=0 $Y2=0
cc_170 N_A_80_241#_c_145_n N_A_M1018_g 0.0101275f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_171 N_A_80_241#_c_146_n N_A_M1018_g 0.022218f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_172 N_A_80_241#_M1027_g N_A_c_458_n 0.0104164f $X=5.43 $Y=0.805 $X2=0 $Y2=0
cc_173 N_A_80_241#_c_154_p N_A_c_460_n 9.21836e-19 $X=1.635 $Y=0.92 $X2=0 $Y2=0
cc_174 N_A_80_241#_c_145_n N_A_c_460_n 0.0024114f $X=5.45 $Y=1.45 $X2=0 $Y2=0
cc_175 N_A_80_241#_M1007_d N_A_c_464_n 0.00191751f $X=1.495 $Y=0.625 $X2=0 $Y2=0
cc_176 N_A_80_241#_c_154_p N_A_c_464_n 0.0156527f $X=1.635 $Y=0.92 $X2=0 $Y2=0
cc_177 N_A_80_241#_M1027_g N_A_1101_119#_c_571_n 0.00542921f $X=5.43 $Y=0.805
+ $X2=0 $Y2=0
cc_178 N_A_80_241#_c_145_n N_A_1101_119#_c_571_n 0.00162117f $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_179 N_A_80_241#_c_146_n N_A_1101_119#_c_571_n 0.00105959f $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_180 N_A_80_241#_M1016_g N_A_1101_119#_c_572_n 0.00329008f $X=5.43 $Y=2.165
+ $X2=0 $Y2=0
cc_181 N_A_80_241#_c_145_n N_A_1101_119#_c_572_n 0.0128545f $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_182 N_A_80_241#_c_146_n N_A_1101_119#_c_572_n 0.00354731f $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_183 N_A_80_241#_M1016_g N_A_1101_119#_c_580_n 0.00172382f $X=5.43 $Y=2.165
+ $X2=0 $Y2=0
cc_184 N_A_80_241#_c_145_n N_A_1101_119#_c_580_n 0.00145571f $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_185 N_A_80_241#_c_146_n N_A_1101_119#_c_580_n 7.60101e-19 $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_186 N_A_80_241#_c_148_n N_COUT_c_627_n 0.00482706f $X=0.61 $Y=1.37 $X2=0
+ $Y2=0
cc_187 N_A_80_241#_M1021_g COUT 0.00564061f $X=0.63 $Y=0.835 $X2=0 $Y2=0
cc_188 N_A_80_241#_c_147_n COUT 0.0228107f $X=0.61 $Y=1.37 $X2=0 $Y2=0
cc_189 N_A_80_241#_c_148_n COUT 0.0249493f $X=0.61 $Y=1.37 $X2=0 $Y2=0
cc_190 N_A_80_241#_M1024_g N_VPWR_c_640_n 0.00709812f $X=0.475 $Y=2.045 $X2=0
+ $Y2=0
cc_191 N_A_80_241#_c_143_n N_VPWR_c_640_n 0.00602035f $X=1.47 $Y=1.45 $X2=0
+ $Y2=0
cc_192 N_A_80_241#_c_147_n N_VPWR_c_640_n 0.00503554f $X=0.61 $Y=1.37 $X2=0
+ $Y2=0
cc_193 N_A_80_241#_c_148_n N_VPWR_c_640_n 0.00231964f $X=0.61 $Y=1.37 $X2=0
+ $Y2=0
cc_194 N_A_80_241#_M1016_g N_VPWR_c_644_n 0.0113387f $X=5.43 $Y=2.165 $X2=0
+ $Y2=0
cc_195 N_A_80_241#_c_145_n N_VPWR_c_647_n 0.00637856f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_196 N_A_80_241#_c_145_n N_A_385_367#_c_740_n 0.0615696f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_197 N_A_80_241#_c_144_n N_A_385_367#_c_741_n 0.00771601f $X=1.635 $Y=1.98
+ $X2=0 $Y2=0
cc_198 N_A_80_241#_c_145_n N_A_385_367#_c_741_n 0.0162494f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_199 N_A_80_241#_c_145_n N_A_385_367#_c_742_n 0.0152619f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_200 N_A_80_241#_M1016_g N_A_843_391#_c_762_n 0.00241866f $X=5.43 $Y=2.165
+ $X2=0 $Y2=0
cc_201 N_A_80_241#_c_145_n N_A_843_391#_c_762_n 0.0612212f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_202 N_A_80_241#_c_146_n N_A_843_391#_c_762_n 8.85824e-19 $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_203 N_A_80_241#_c_145_n N_A_843_391#_c_763_n 0.0166894f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_204 N_A_80_241#_M1016_g N_A_843_391#_c_764_n 7.11755e-19 $X=5.43 $Y=2.165
+ $X2=0 $Y2=0
cc_205 N_A_80_241#_M1021_g N_VGND_c_798_n 0.00322999f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_206 N_A_80_241#_c_143_n N_VGND_c_798_n 0.00735359f $X=1.47 $Y=1.45 $X2=0
+ $Y2=0
cc_207 N_A_80_241#_c_148_n N_VGND_c_798_n 6.93622e-19 $X=0.61 $Y=1.37 $X2=0
+ $Y2=0
cc_208 N_A_80_241#_c_145_n N_VGND_c_800_n 0.00795516f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_209 N_A_80_241#_M1027_g N_VGND_c_801_n 0.0011413f $X=5.43 $Y=0.805 $X2=0
+ $Y2=0
cc_210 N_A_80_241#_M1021_g N_VGND_c_803_n 0.00415323f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_211 N_A_80_241#_M1021_g N_VGND_c_814_n 0.00469432f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_212 N_A_80_241#_M1027_g N_VGND_c_814_n 9.39239e-19 $X=5.43 $Y=0.805 $X2=0
+ $Y2=0
cc_213 N_A_80_241#_c_145_n N_A_385_125#_c_883_n 0.0685339f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_214 N_A_80_241#_c_154_p N_A_385_125#_c_884_n 0.0180988f $X=1.635 $Y=0.92
+ $X2=0 $Y2=0
cc_215 N_A_80_241#_c_145_n N_A_385_125#_c_884_n 0.024377f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_216 N_A_80_241#_M1027_g N_A_843_119#_c_909_n 0.00218937f $X=5.43 $Y=0.805
+ $X2=0 $Y2=0
cc_217 N_A_80_241#_c_145_n N_A_843_119#_c_909_n 0.0599491f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_218 N_A_80_241#_c_146_n N_A_843_119#_c_909_n 8.77827e-19 $X=5.45 $Y=1.45
+ $X2=0 $Y2=0
cc_219 N_A_80_241#_c_145_n N_A_843_119#_c_910_n 0.014395f $X=5.45 $Y=1.45 $X2=0
+ $Y2=0
cc_220 N_B_M1007_g N_CIN_M1008_g 0.0691081f $X=1.42 $Y=0.835 $X2=0 $Y2=0
cc_221 N_B_c_252_n N_CIN_M1008_g 9.92836e-19 $X=1.25 $Y=2.79 $X2=0 $Y2=0
cc_222 N_B_c_253_n N_CIN_M1008_g 0.0157639f $X=2.135 $Y=2.425 $X2=0 $Y2=0
cc_223 N_B_c_257_n N_CIN_M1008_g 0.00683111f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_224 N_B_M1006_g N_CIN_c_380_n 0.00201695f $X=4.14 $Y=2.165 $X2=0 $Y2=0
cc_225 N_B_c_253_n N_CIN_c_380_n 2.26873e-19 $X=2.135 $Y=2.425 $X2=0 $Y2=0
cc_226 N_B_c_257_n N_CIN_c_380_n 0.00297086f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_227 N_B_c_259_n N_CIN_c_380_n 0.0193612f $X=3.525 $Y=2.7 $X2=0 $Y2=0
cc_228 N_B_c_261_n N_CIN_c_380_n 0.0406679f $X=3.5 $Y=2.805 $X2=0 $Y2=0
cc_229 N_B_M1023_g N_CIN_M1017_g 0.0613729f $X=4.14 $Y=0.805 $X2=0 $Y2=0
cc_230 N_B_c_255_n N_CIN_M1017_g 0.0146954f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_231 N_B_c_255_n N_CIN_c_383_n 0.0189515f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_232 N_B_M1022_g N_CIN_M1000_g 0.163472f $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_233 N_B_c_255_n N_CIN_M1000_g 0.0121531f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_234 N_B_c_253_n N_CIN_c_387_n 0.00359083f $X=2.135 $Y=2.425 $X2=0 $Y2=0
cc_235 N_B_c_257_n N_CIN_c_387_n 0.00634211f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_236 N_B_c_258_n N_CIN_c_387_n 0.0138137f $X=1.42 $Y=2.79 $X2=0 $Y2=0
cc_237 N_B_c_252_n N_CIN_c_388_n 0.0141105f $X=1.25 $Y=2.79 $X2=0 $Y2=0
cc_238 N_B_c_253_n N_CIN_c_388_n 0.0257092f $X=2.135 $Y=2.425 $X2=0 $Y2=0
cc_239 N_B_c_257_n N_CIN_c_388_n 0.0222788f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_240 N_B_c_258_n N_CIN_c_388_n 0.00339887f $X=1.42 $Y=2.79 $X2=0 $Y2=0
cc_241 N_B_M1007_g N_A_M1013_g 0.116596f $X=1.42 $Y=0.835 $X2=0 $Y2=0
cc_242 N_B_c_254_n N_A_M1013_g 0.00401163f $X=1.415 $Y=2.425 $X2=0 $Y2=0
cc_243 N_B_c_258_n N_A_M1013_g 0.00276667f $X=1.42 $Y=2.79 $X2=0 $Y2=0
cc_244 N_B_M1007_g N_A_c_452_n 0.00740131f $X=1.42 $Y=0.835 $X2=0 $Y2=0
cc_245 N_B_M1009_g N_A_M1010_g 0.0226866f $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_246 N_B_c_257_n N_A_M1010_g 0.00540179f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_247 N_B_c_261_n N_A_M1010_g 0.00143235f $X=3.5 $Y=2.805 $X2=0 $Y2=0
cc_248 N_B_M1009_g N_A_M1026_g 0.0154075f $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_249 N_B_M1009_g N_A_c_456_n 0.00907339f $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_250 N_B_M1023_g N_A_c_456_n 0.0104164f $X=4.14 $Y=0.805 $X2=0 $Y2=0
cc_251 N_B_c_255_n N_A_M1018_g 4.80386e-19 $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_252 N_B_M1022_g N_A_c_458_n 0.0104164f $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_253 N_B_M1022_g N_A_M1012_g 0.12656f $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_254 N_B_M1009_g N_A_c_463_n 4.92694e-19 $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_255 N_B_M1007_g N_A_c_464_n 0.0126992f $X=1.42 $Y=0.835 $X2=0 $Y2=0
cc_256 N_B_M1022_g N_A_1101_119#_c_571_n 0.00273707f $X=6.26 $Y=0.805 $X2=0
+ $Y2=0
cc_257 N_B_M1022_g N_A_1101_119#_c_572_n 0.00406858f $X=6.26 $Y=0.805 $X2=0
+ $Y2=0
cc_258 N_B_M1022_g N_A_1101_119#_c_573_n 0.0184418f $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_259 N_B_M1022_g N_A_1101_119#_c_580_n 0.00213148f $X=6.26 $Y=0.805 $X2=0
+ $Y2=0
cc_260 N_B_M1007_g N_VPWR_c_640_n 0.00103634f $X=1.42 $Y=0.835 $X2=0 $Y2=0
cc_261 N_B_c_252_n N_VPWR_c_640_n 0.0235091f $X=1.25 $Y=2.79 $X2=0 $Y2=0
cc_262 N_B_c_254_n N_VPWR_c_640_n 0.0119492f $X=1.415 $Y=2.425 $X2=0 $Y2=0
cc_263 N_B_c_258_n N_VPWR_c_640_n 0.00884002f $X=1.42 $Y=2.79 $X2=0 $Y2=0
cc_264 N_B_c_244_n N_VPWR_c_641_n 0.00785419f $X=2.945 $Y=1.665 $X2=0 $Y2=0
cc_265 N_B_c_236_n N_VPWR_c_641_n 2.94442e-19 $X=3.36 $Y=1.59 $X2=0 $Y2=0
cc_266 N_B_c_237_n N_VPWR_c_641_n 0.0048091f $X=4.065 $Y=1.59 $X2=0 $Y2=0
cc_267 N_B_c_255_n N_VPWR_c_641_n 0.00547321f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_268 N_B_c_259_n N_VPWR_c_641_n 0.00440824f $X=3.525 $Y=2.7 $X2=0 $Y2=0
cc_269 N_B_c_260_n N_VPWR_c_641_n 0.0173918f $X=3.525 $Y=2.535 $X2=0 $Y2=0
cc_270 N_B_c_261_n N_VPWR_c_641_n 0.065383f $X=3.5 $Y=2.805 $X2=0 $Y2=0
cc_271 N_B_M1006_g N_VPWR_c_642_n 0.0114177f $X=4.14 $Y=2.165 $X2=0 $Y2=0
cc_272 N_B_c_255_n N_VPWR_c_642_n 0.0350758f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_273 N_B_M1022_g N_VPWR_c_644_n 0.0154471f $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_274 N_B_c_255_n N_VPWR_c_644_n 0.0890462f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_275 N_B_c_256_n N_VPWR_c_644_n 0.00426207f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_276 N_B_M1022_g N_VPWR_c_645_n 0.0036275f $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_277 N_B_c_255_n N_VPWR_c_645_n 0.00844246f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_278 N_B_c_256_n N_VPWR_c_645_n 0.00625232f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_279 N_B_c_244_n N_VPWR_c_646_n 0.00320791f $X=2.945 $Y=1.665 $X2=0 $Y2=0
cc_280 N_B_c_257_n N_VPWR_c_646_n 0.00706295f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_281 N_B_c_260_n N_VPWR_c_646_n 2.57983e-19 $X=3.525 $Y=2.535 $X2=0 $Y2=0
cc_282 N_B_c_261_n N_VPWR_c_646_n 0.0268617f $X=3.5 $Y=2.805 $X2=0 $Y2=0
cc_283 N_B_c_237_n N_VPWR_c_647_n 0.00282749f $X=4.065 $Y=1.59 $X2=0 $Y2=0
cc_284 N_B_M1006_g N_VPWR_c_647_n 0.00101299f $X=4.14 $Y=2.165 $X2=0 $Y2=0
cc_285 N_B_c_255_n N_VPWR_c_647_n 0.012749f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_286 N_B_c_259_n N_VPWR_c_647_n 0.00263784f $X=3.525 $Y=2.7 $X2=0 $Y2=0
cc_287 N_B_c_260_n N_VPWR_c_647_n 0.00656853f $X=3.525 $Y=2.535 $X2=0 $Y2=0
cc_288 N_B_c_255_n N_VPWR_c_648_n 0.0129606f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_289 N_B_M1022_g N_VPWR_c_649_n 0.00182906f $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_290 N_B_c_252_n N_VPWR_c_650_n 0.00925924f $X=1.25 $Y=2.79 $X2=0 $Y2=0
cc_291 N_B_c_256_n N_VPWR_c_650_n 0.00807533f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_292 N_B_c_257_n N_VPWR_c_650_n 0.0079474f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_293 N_B_c_258_n N_VPWR_c_650_n 0.00955224f $X=1.42 $Y=2.79 $X2=0 $Y2=0
cc_294 N_B_c_261_n N_VPWR_c_650_n 0.182217f $X=3.5 $Y=2.805 $X2=0 $Y2=0
cc_295 N_B_c_252_n N_VPWR_c_639_n 0.0108904f $X=1.25 $Y=2.79 $X2=0 $Y2=0
cc_296 N_B_c_253_n N_VPWR_c_639_n 0.0121795f $X=2.135 $Y=2.425 $X2=0 $Y2=0
cc_297 N_B_c_256_n N_VPWR_c_639_n 0.011167f $X=6.35 $Y=2.91 $X2=0 $Y2=0
cc_298 N_B_c_257_n N_VPWR_c_639_n 0.00557914f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_299 N_B_c_258_n N_VPWR_c_639_n 0.0127824f $X=1.42 $Y=2.79 $X2=0 $Y2=0
cc_300 N_B_c_261_n N_VPWR_c_639_n 0.136291f $X=3.5 $Y=2.805 $X2=0 $Y2=0
cc_301 N_B_c_244_n N_A_385_367#_c_740_n 0.0109591f $X=2.945 $Y=1.665 $X2=0 $Y2=0
cc_302 N_B_c_257_n N_A_385_367#_c_740_n 0.00417946f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_303 N_B_c_253_n N_A_385_367#_c_741_n 0.0117621f $X=2.135 $Y=2.425 $X2=0 $Y2=0
cc_304 N_B_c_257_n N_A_385_367#_c_741_n 0.00185041f $X=2.22 $Y=2.425 $X2=0 $Y2=0
cc_305 N_B_c_236_n N_A_385_367#_c_742_n 0.00351337f $X=3.36 $Y=1.59 $X2=0 $Y2=0
cc_306 N_B_c_260_n N_A_385_367#_c_742_n 0.00876196f $X=3.525 $Y=2.535 $X2=0
+ $Y2=0
cc_307 N_B_M1006_g N_A_843_391#_c_761_n 0.0017418f $X=4.14 $Y=2.165 $X2=0 $Y2=0
cc_308 N_B_M1006_g N_A_843_391#_c_763_n 0.00551383f $X=4.14 $Y=2.165 $X2=0 $Y2=0
cc_309 N_B_M1009_g N_VGND_c_799_n 0.00345216f $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_310 N_B_c_237_n N_VGND_c_800_n 8.27465e-19 $X=4.065 $Y=1.59 $X2=0 $Y2=0
cc_311 N_B_M1023_g N_VGND_c_800_n 0.00367548f $X=4.14 $Y=0.805 $X2=0 $Y2=0
cc_312 N_B_M1023_g N_VGND_c_801_n 6.94973e-19 $X=4.14 $Y=0.805 $X2=0 $Y2=0
cc_313 N_B_M1009_g N_VGND_c_814_n 9.49986e-19 $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_314 N_B_M1023_g N_VGND_c_814_n 9.39239e-19 $X=4.14 $Y=0.805 $X2=0 $Y2=0
cc_315 N_B_M1022_g N_VGND_c_814_n 9.39239e-19 $X=6.26 $Y=0.805 $X2=0 $Y2=0
cc_316 N_B_M1009_g N_A_385_125#_c_883_n 0.016098f $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_317 N_B_c_236_n N_A_385_125#_c_883_n 8.31844e-19 $X=3.36 $Y=1.59 $X2=0 $Y2=0
cc_318 N_B_M1009_g N_A_385_125#_c_884_n 6.2538e-19 $X=2.945 $Y=0.835 $X2=0 $Y2=0
cc_319 N_B_M1023_g N_A_843_119#_c_910_n 0.00516145f $X=4.14 $Y=0.805 $X2=0 $Y2=0
cc_320 N_CIN_M1008_g N_A_c_452_n 0.00740131f $X=1.85 $Y=0.835 $X2=0 $Y2=0
cc_321 N_CIN_c_380_n N_A_M1010_g 0.00143578f $X=4.495 $Y=3.15 $X2=0 $Y2=0
cc_322 N_CIN_M1008_g N_A_M1026_g 0.0139657f $X=1.85 $Y=0.835 $X2=0 $Y2=0
cc_323 N_CIN_M1017_g N_A_c_456_n 0.0103107f $X=4.57 $Y=0.805 $X2=0 $Y2=0
cc_324 N_CIN_M1017_g N_A_M1018_g 0.0629986f $X=4.57 $Y=0.805 $X2=0 $Y2=0
cc_325 N_CIN_c_383_n N_A_M1018_g 0.00201695f $X=5.825 $Y=3.15 $X2=0 $Y2=0
cc_326 N_CIN_M1000_g N_A_c_458_n 0.00991962f $X=5.9 $Y=0.805 $X2=0 $Y2=0
cc_327 N_CIN_M1008_g N_A_c_460_n 0.0401025f $X=1.85 $Y=0.835 $X2=0 $Y2=0
cc_328 N_CIN_M1008_g N_A_c_463_n 0.00109563f $X=1.85 $Y=0.835 $X2=0 $Y2=0
cc_329 N_CIN_M1008_g N_A_c_464_n 0.013157f $X=1.85 $Y=0.835 $X2=0 $Y2=0
cc_330 N_CIN_M1000_g N_A_1101_119#_c_571_n 0.017234f $X=5.9 $Y=0.805 $X2=0 $Y2=0
cc_331 N_CIN_M1000_g N_A_1101_119#_c_572_n 0.0181891f $X=5.9 $Y=0.805 $X2=0
+ $Y2=0
cc_332 N_CIN_M1000_g N_A_1101_119#_c_573_n 0.00243077f $X=5.9 $Y=0.805 $X2=0
+ $Y2=0
cc_333 N_CIN_M1000_g N_A_1101_119#_c_580_n 0.0115494f $X=5.9 $Y=0.805 $X2=0
+ $Y2=0
cc_334 N_CIN_M1017_g N_VPWR_c_642_n 0.0147067f $X=4.57 $Y=0.805 $X2=0 $Y2=0
cc_335 N_CIN_M1017_g N_VPWR_c_643_n 6.65496e-19 $X=4.57 $Y=0.805 $X2=0 $Y2=0
cc_336 N_CIN_M1000_g N_VPWR_c_644_n 0.0118409f $X=5.9 $Y=0.805 $X2=0 $Y2=0
cc_337 N_CIN_c_381_n N_VPWR_c_650_n 0.0963201f $X=2.035 $Y=3.15 $X2=0 $Y2=0
cc_338 N_CIN_c_388_n N_VPWR_c_650_n 0.0222841f $X=1.87 $Y=2.9 $X2=0 $Y2=0
cc_339 N_CIN_c_380_n N_VPWR_c_639_n 0.0587652f $X=4.495 $Y=3.15 $X2=0 $Y2=0
cc_340 N_CIN_c_381_n N_VPWR_c_639_n 0.0107987f $X=2.035 $Y=3.15 $X2=0 $Y2=0
cc_341 N_CIN_c_383_n N_VPWR_c_639_n 0.0340769f $X=5.825 $Y=3.15 $X2=0 $Y2=0
cc_342 N_CIN_c_386_n N_VPWR_c_639_n 0.00375056f $X=4.57 $Y=3.15 $X2=0 $Y2=0
cc_343 N_CIN_c_388_n N_VPWR_c_639_n 0.0125559f $X=1.87 $Y=2.9 $X2=0 $Y2=0
cc_344 N_CIN_M1008_g N_A_385_367#_c_741_n 9.83941e-19 $X=1.85 $Y=0.835 $X2=0
+ $Y2=0
cc_345 N_CIN_M1017_g N_A_843_391#_c_761_n 9.4709e-19 $X=4.57 $Y=0.805 $X2=0
+ $Y2=0
cc_346 N_CIN_M1017_g N_A_843_391#_c_762_n 0.0119084f $X=4.57 $Y=0.805 $X2=0
+ $Y2=0
cc_347 N_CIN_M1017_g N_VGND_c_801_n 0.00773664f $X=4.57 $Y=0.805 $X2=0 $Y2=0
cc_348 N_CIN_M1017_g N_VGND_c_814_n 7.88961e-19 $X=4.57 $Y=0.805 $X2=0 $Y2=0
cc_349 N_CIN_M1000_g N_VGND_c_814_n 9.39239e-19 $X=5.9 $Y=0.805 $X2=0 $Y2=0
cc_350 N_CIN_M1008_g N_A_385_125#_c_884_n 0.00227433f $X=1.85 $Y=0.835 $X2=0
+ $Y2=0
cc_351 N_CIN_M1017_g N_A_843_119#_c_909_n 0.0135964f $X=4.57 $Y=0.805 $X2=0
+ $Y2=0
cc_352 N_A_M1012_g N_A_1101_119#_M1001_g 0.0136913f $X=6.62 $Y=0.805 $X2=0 $Y2=0
cc_353 N_A_c_458_n N_A_1101_119#_c_571_n 0.00431159f $X=6.545 $Y=0.18 $X2=0
+ $Y2=0
cc_354 N_A_M1012_g N_A_1101_119#_c_573_n 0.0186515f $X=6.62 $Y=0.805 $X2=0 $Y2=0
cc_355 N_A_M1012_g N_A_1101_119#_c_574_n 0.00277702f $X=6.62 $Y=0.805 $X2=0
+ $Y2=0
cc_356 N_A_M1012_g N_A_1101_119#_c_575_n 0.043786f $X=6.62 $Y=0.805 $X2=0 $Y2=0
cc_357 N_A_M1012_g N_A_1101_119#_c_576_n 0.0135433f $X=6.62 $Y=0.805 $X2=0 $Y2=0
cc_358 N_A_M1013_g N_VPWR_c_640_n 0.00754175f $X=1.06 $Y=0.835 $X2=0 $Y2=0
cc_359 N_A_M1018_g N_VPWR_c_643_n 0.00123209f $X=5 $Y=0.805 $X2=0 $Y2=0
cc_360 N_A_M1018_g N_VPWR_c_644_n 0.00847061f $X=5 $Y=0.805 $X2=0 $Y2=0
cc_361 N_A_M1012_g N_VPWR_c_644_n 0.0094046f $X=6.62 $Y=0.805 $X2=0 $Y2=0
cc_362 N_A_M1010_g N_VPWR_c_646_n 0.00726707f $X=2.28 $Y=2.045 $X2=0 $Y2=0
cc_363 N_A_M1012_g N_VPWR_c_649_n 0.00890308f $X=6.62 $Y=0.805 $X2=0 $Y2=0
cc_364 N_A_M1010_g N_A_385_367#_c_740_n 0.0123816f $X=2.28 $Y=2.045 $X2=0 $Y2=0
cc_365 N_A_M1010_g N_A_385_367#_c_741_n 2.96346e-19 $X=2.28 $Y=2.045 $X2=0 $Y2=0
cc_366 N_A_M1018_g N_A_843_391#_c_762_n 0.0119084f $X=5 $Y=0.805 $X2=0 $Y2=0
cc_367 N_A_M1018_g N_A_843_391#_c_764_n 9.4709e-19 $X=5 $Y=0.805 $X2=0 $Y2=0
cc_368 N_A_c_453_n N_VGND_c_798_n 0.0120891f $X=1.135 $Y=0.18 $X2=0 $Y2=0
cc_369 N_A_c_464_n N_VGND_c_798_n 0.0276317f $X=2.058 $Y=0.452 $X2=0 $Y2=0
cc_370 N_A_M1026_g N_VGND_c_799_n 0.00118099f $X=2.36 $Y=0.835 $X2=0 $Y2=0
cc_371 N_A_c_456_n N_VGND_c_799_n 0.0166369f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_372 A N_VGND_c_799_n 0.0223886f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_373 N_A_c_463_n N_VGND_c_799_n 0.0027103f $X=2.33 $Y=0.18 $X2=0 $Y2=0
cc_374 N_A_c_456_n N_VGND_c_800_n 0.0183754f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_375 N_A_c_456_n N_VGND_c_801_n 0.0173284f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_376 N_A_M1018_g N_VGND_c_801_n 0.0207826f $X=5 $Y=0.805 $X2=0 $Y2=0
cc_377 N_A_c_461_n N_VGND_c_801_n 0.00460513f $X=5 $Y=0.18 $X2=0 $Y2=0
cc_378 N_A_c_458_n N_VGND_c_802_n 0.0174933f $X=6.545 $Y=0.18 $X2=0 $Y2=0
cc_379 N_A_M1026_g N_VGND_c_844_n 0.00529664f $X=2.36 $Y=0.835 $X2=0 $Y2=0
cc_380 N_A_c_456_n N_VGND_c_844_n 0.00209921f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_381 N_A_c_453_n N_VGND_c_805_n 0.0396845f $X=1.135 $Y=0.18 $X2=0 $Y2=0
cc_382 A N_VGND_c_805_n 0.0265057f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_383 N_A_c_464_n N_VGND_c_805_n 0.0603444f $X=2.058 $Y=0.452 $X2=0 $Y2=0
cc_384 N_A_c_456_n N_VGND_c_807_n 0.0323518f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_385 N_A_c_456_n N_VGND_c_809_n 0.0189055f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_386 N_A_c_461_n N_VGND_c_811_n 0.0574859f $X=5 $Y=0.18 $X2=0 $Y2=0
cc_387 N_A_c_452_n N_VGND_c_814_n 0.0242175f $X=2.165 $Y=0.18 $X2=0 $Y2=0
cc_388 N_A_c_453_n N_VGND_c_814_n 0.0107428f $X=1.135 $Y=0.18 $X2=0 $Y2=0
cc_389 N_A_c_456_n N_VGND_c_814_n 0.0699675f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_390 N_A_c_458_n N_VGND_c_814_n 0.0704551f $X=6.545 $Y=0.18 $X2=0 $Y2=0
cc_391 N_A_c_461_n N_VGND_c_814_n 0.00749832f $X=5 $Y=0.18 $X2=0 $Y2=0
cc_392 A N_VGND_c_814_n 0.01454f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_393 N_A_c_463_n N_VGND_c_814_n 0.00795132f $X=2.33 $Y=0.18 $X2=0 $Y2=0
cc_394 N_A_c_464_n N_VGND_c_814_n 0.0320939f $X=2.058 $Y=0.452 $X2=0 $Y2=0
cc_395 N_A_c_464_n A_227_125# 0.00403009f $X=2.058 $Y=0.452 $X2=-0.19 $Y2=-0.245
cc_396 A N_A_385_125#_M1008_d 0.00193032f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_397 N_A_c_464_n N_A_385_125#_M1008_d 8.66345e-19 $X=2.058 $Y=0.452 $X2=-0.19
+ $Y2=-0.245
cc_398 N_A_M1026_g N_A_385_125#_c_883_n 0.00752544f $X=2.36 $Y=0.835 $X2=0 $Y2=0
cc_399 N_A_c_460_n N_A_385_125#_c_883_n 0.00222426f $X=2.36 $Y=1.23 $X2=0 $Y2=0
cc_400 A N_A_385_125#_c_883_n 0.00412315f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_401 N_A_c_463_n N_A_385_125#_c_883_n 9.1249e-19 $X=2.33 $Y=0.18 $X2=0 $Y2=0
cc_402 N_A_c_456_n N_A_385_125#_c_898_n 0.00349426f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_403 N_A_M1026_g N_A_385_125#_c_884_n 0.00627022f $X=2.36 $Y=0.835 $X2=0 $Y2=0
cc_404 N_A_c_460_n N_A_385_125#_c_884_n 0.00349129f $X=2.36 $Y=1.23 $X2=0 $Y2=0
cc_405 A N_A_385_125#_c_884_n 0.0136914f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_406 N_A_c_463_n N_A_385_125#_c_884_n 3.13248e-19 $X=2.33 $Y=0.18 $X2=0 $Y2=0
cc_407 N_A_c_464_n N_A_385_125#_c_884_n 0.00536565f $X=2.058 $Y=0.452 $X2=0
+ $Y2=0
cc_408 N_A_c_456_n N_A_843_119#_c_917_n 0.00323202f $X=4.925 $Y=0.18 $X2=0 $Y2=0
cc_409 N_A_M1018_g N_A_843_119#_c_909_n 0.0138674f $X=5 $Y=0.805 $X2=0 $Y2=0
cc_410 N_A_c_458_n N_A_843_119#_c_919_n 0.00263199f $X=6.545 $Y=0.18 $X2=0 $Y2=0
cc_411 N_A_1101_119#_c_580_n N_VPWR_c_644_n 0.0256003f $X=5.88 $Y=2.08 $X2=0
+ $Y2=0
cc_412 N_A_1101_119#_M1001_g N_VPWR_c_649_n 0.00394083f $X=7.205 $Y=2.165 $X2=0
+ $Y2=0
cc_413 N_A_1101_119#_c_570_n N_VPWR_c_649_n 0.00337541f $X=7.092 $Y=1.795 $X2=0
+ $Y2=0
cc_414 N_A_1101_119#_c_574_n N_VPWR_c_649_n 6.79568e-19 $X=7.07 $Y=1.29 $X2=0
+ $Y2=0
cc_415 N_A_1101_119#_M1001_g N_VPWR_c_639_n 0.00387136f $X=7.205 $Y=2.165 $X2=0
+ $Y2=0
cc_416 N_A_1101_119#_c_572_n N_A_843_391#_c_762_n 0.00699064f $X=5.88 $Y=1.915
+ $X2=0 $Y2=0
cc_417 N_A_1101_119#_c_572_n N_A_843_391#_c_764_n 0.00110213f $X=5.88 $Y=1.915
+ $X2=0 $Y2=0
cc_418 N_A_1101_119#_c_580_n N_A_843_391#_c_764_n 0.0110398f $X=5.88 $Y=2.08
+ $X2=0 $Y2=0
cc_419 N_A_1101_119#_c_574_n N_SUM_c_784_n 0.00301371f $X=7.07 $Y=1.29 $X2=0
+ $Y2=0
cc_420 N_A_1101_119#_c_575_n N_SUM_c_784_n 0.00475335f $X=7.07 $Y=1.29 $X2=0
+ $Y2=0
cc_421 N_A_1101_119#_c_576_n N_SUM_c_784_n 0.00335402f $X=7.092 $Y=1.125 $X2=0
+ $Y2=0
cc_422 N_A_1101_119#_c_574_n SUM 0.0475752f $X=7.07 $Y=1.29 $X2=0 $Y2=0
cc_423 N_A_1101_119#_c_575_n SUM 0.0287265f $X=7.07 $Y=1.29 $X2=0 $Y2=0
cc_424 N_A_1101_119#_c_576_n SUM 0.00483137f $X=7.092 $Y=1.125 $X2=0 $Y2=0
cc_425 N_A_1101_119#_c_573_n N_VGND_c_802_n 0.012026f $X=6.985 $Y=1.21 $X2=0
+ $Y2=0
cc_426 N_A_1101_119#_c_575_n N_VGND_c_802_n 3.61281e-19 $X=7.07 $Y=1.29 $X2=0
+ $Y2=0
cc_427 N_A_1101_119#_c_576_n N_VGND_c_802_n 0.00314874f $X=7.092 $Y=1.125 $X2=0
+ $Y2=0
cc_428 N_A_1101_119#_c_571_n N_VGND_c_811_n 0.00557805f $X=5.88 $Y=1.295 $X2=0
+ $Y2=0
cc_429 N_A_1101_119#_c_576_n N_VGND_c_813_n 0.00416091f $X=7.092 $Y=1.125 $X2=0
+ $Y2=0
cc_430 N_A_1101_119#_c_571_n N_VGND_c_814_n 0.00920022f $X=5.88 $Y=1.295 $X2=0
+ $Y2=0
cc_431 N_A_1101_119#_c_576_n N_VGND_c_814_n 0.00477801f $X=7.092 $Y=1.125 $X2=0
+ $Y2=0
cc_432 N_A_1101_119#_c_571_n N_A_843_119#_c_909_n 0.0075828f $X=5.88 $Y=1.295
+ $X2=0 $Y2=0
cc_433 COUT N_VPWR_c_640_n 0.0548272f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_434 COUT N_VPWR_c_652_n 0.00563668f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_435 COUT N_VPWR_c_639_n 0.00642236f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_436 N_COUT_c_627_n N_VGND_c_803_n 0.00581815f $X=0.415 $Y=0.86 $X2=0 $Y2=0
cc_437 N_COUT_c_627_n N_VGND_c_814_n 0.0102363f $X=0.415 $Y=0.86 $X2=0 $Y2=0
cc_438 N_VPWR_M1010_d N_A_385_367#_c_740_n 0.00731913f $X=2.355 $Y=1.835 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_641_n N_A_385_367#_c_740_n 0.00725056f $X=3.82 $Y=2.35 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_646_n N_A_385_367#_c_740_n 0.0242771f $X=2.65 $Y=2.15 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_641_n N_A_385_367#_c_742_n 0.0148992f $X=3.82 $Y=2.35 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_647_n N_A_385_367#_c_742_n 6.22467e-19 $X=3.93 $Y=2.35 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_642_n N_A_843_391#_c_761_n 0.0144312f $X=4.68 $Y=2.51 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_642_n N_A_843_391#_c_762_n 0.00627406f $X=4.68 $Y=2.51 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_643_n N_A_843_391#_c_762_n 0.0144312f $X=4.785 $Y=2.23 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_644_n N_A_843_391#_c_762_n 0.00627406f $X=6.67 $Y=2.51 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_644_n N_A_843_391#_c_764_n 0.0144312f $X=6.67 $Y=2.51 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_649_n SUM 0.0296f $X=6.835 $Y=2.23 $X2=0 $Y2=0
cc_449 N_VPWR_c_653_n SUM 0.00563668f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_450 N_VPWR_c_639_n SUM 0.00642236f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_451 N_SUM_c_784_n N_VGND_c_813_n 0.00579262f $X=7.43 $Y=0.84 $X2=0 $Y2=0
cc_452 N_SUM_c_784_n N_VGND_c_814_n 0.0112973f $X=7.43 $Y=0.84 $X2=0 $Y2=0
cc_453 N_VGND_M1026_d N_A_385_125#_c_883_n 0.00413587f $X=2.435 $Y=0.625 $X2=0
+ $Y2=0
cc_454 N_VGND_c_844_n N_A_385_125#_c_883_n 0.0209187f $X=2.76 $Y=0.74 $X2=0
+ $Y2=0
cc_455 N_VGND_c_800_n N_A_385_125#_c_898_n 0.00528386f $X=3.925 $Y=0.74 $X2=0
+ $Y2=0
cc_456 N_VGND_c_807_n N_A_385_125#_c_898_n 0.00300513f $X=3.82 $Y=0 $X2=0 $Y2=0
cc_457 N_VGND_c_814_n N_A_385_125#_c_898_n 0.00494077f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_809_n N_A_843_119#_c_917_n 0.00287f $X=4.62 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_814_n N_A_843_119#_c_917_n 0.00458436f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_460 N_VGND_M1017_d N_A_843_119#_c_909_n 0.00180746f $X=4.645 $Y=0.595 $X2=0
+ $Y2=0
cc_461 N_VGND_c_801_n N_A_843_119#_c_909_n 0.0163515f $X=4.785 $Y=0.72 $X2=0
+ $Y2=0
cc_462 N_VGND_c_811_n N_A_843_119#_c_919_n 0.00287035f $X=6.73 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_c_814_n N_A_843_119#_c_919_n 0.00458436f $X=7.44 $Y=0 $X2=0 $Y2=0
