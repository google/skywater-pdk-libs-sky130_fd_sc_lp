* File: sky130_fd_sc_lp__o32a_0.pxi.spice
* Created: Wed Sep  2 10:25:51 2020
* 
x_PM_SKY130_FD_SC_LP__O32A_0%A_97_309# N_A_97_309#_M1007_d N_A_97_309#_M1002_d
+ N_A_97_309#_M1000_g N_A_97_309#_M1011_g N_A_97_309#_c_91_n N_A_97_309#_c_92_n
+ N_A_97_309#_c_86_n N_A_97_309#_c_87_n N_A_97_309#_c_94_n N_A_97_309#_c_95_n
+ N_A_97_309#_c_96_n N_A_97_309#_c_97_n N_A_97_309#_c_88_n N_A_97_309#_c_99_n
+ N_A_97_309#_c_89_n PM_SKY130_FD_SC_LP__O32A_0%A_97_309#
x_PM_SKY130_FD_SC_LP__O32A_0%A1 N_A1_M1005_g N_A1_c_171_n N_A1_M1003_g
+ N_A1_c_167_n N_A1_c_168_n N_A1_c_174_n A1 A1 A1 N_A1_c_170_n
+ PM_SKY130_FD_SC_LP__O32A_0%A1
x_PM_SKY130_FD_SC_LP__O32A_0%A2 N_A2_M1010_g N_A2_M1009_g N_A2_c_220_n
+ N_A2_c_225_n A2 A2 N_A2_c_222_n PM_SKY130_FD_SC_LP__O32A_0%A2
x_PM_SKY130_FD_SC_LP__O32A_0%A3 N_A3_M1002_g N_A3_M1001_g N_A3_c_263_n
+ N_A3_c_268_n A3 A3 N_A3_c_265_n PM_SKY130_FD_SC_LP__O32A_0%A3
x_PM_SKY130_FD_SC_LP__O32A_0%B2 N_B2_M1004_g N_B2_M1007_g N_B2_c_304_n
+ N_B2_c_309_n B2 B2 N_B2_c_306_n PM_SKY130_FD_SC_LP__O32A_0%B2
x_PM_SKY130_FD_SC_LP__O32A_0%B1 N_B1_M1008_g N_B1_M1006_g N_B1_c_344_n
+ N_B1_c_350_n B1 B1 B1 N_B1_c_345_n N_B1_c_346_n N_B1_c_347_n
+ PM_SKY130_FD_SC_LP__O32A_0%B1
x_PM_SKY130_FD_SC_LP__O32A_0%X N_X_M1000_s N_X_M1011_s X X X X X X X N_X_c_377_n
+ X PM_SKY130_FD_SC_LP__O32A_0%X
x_PM_SKY130_FD_SC_LP__O32A_0%VPWR N_VPWR_M1011_d N_VPWR_M1008_d N_VPWR_c_396_n
+ N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n VPWR N_VPWR_c_400_n
+ N_VPWR_c_401_n N_VPWR_c_395_n N_VPWR_c_403_n PM_SKY130_FD_SC_LP__O32A_0%VPWR
x_PM_SKY130_FD_SC_LP__O32A_0%VGND N_VGND_M1000_d N_VGND_M1010_d N_VGND_c_432_n
+ N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n VGND N_VGND_c_436_n
+ N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n PM_SKY130_FD_SC_LP__O32A_0%VGND
x_PM_SKY130_FD_SC_LP__O32A_0%A_271_85# N_A_271_85#_M1005_d N_A_271_85#_M1001_d
+ N_A_271_85#_M1006_d N_A_271_85#_c_482_n N_A_271_85#_c_473_n
+ N_A_271_85#_c_474_n N_A_271_85#_c_494_n N_A_271_85#_c_475_n
+ N_A_271_85#_c_476_n N_A_271_85#_c_477_n N_A_271_85#_c_478_n
+ PM_SKY130_FD_SC_LP__O32A_0%A_271_85#
cc_1 VNB N_A_97_309#_M1000_g 0.0563853f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.635
cc_2 VNB N_A_97_309#_c_86_n 0.00439064f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.71
cc_3 VNB N_A_97_309#_c_87_n 0.0152248f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.71
cc_4 VNB N_A_97_309#_c_88_n 0.00572706f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=2.025
cc_5 VNB N_A_97_309#_c_89_n 0.00411479f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.69
cc_6 VNB N_A1_M1005_g 0.0237478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A1_c_167_n 0.0212971f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.725
cc_8 VNB N_A1_c_168_n 0.00432246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A1 0.00758422f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.025
cc_10 VNB N_A1_c_170_n 0.0158823f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.215
cc_11 VNB N_A2_M1010_g 0.0304136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_220_n 0.0187711f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.215
cc_13 VNB A2 0.00492682f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.725
cc_14 VNB N_A2_c_222_n 0.0152049f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.215
cc_15 VNB N_A3_M1001_g 0.0299489f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.545
cc_16 VNB N_A3_c_263_n 0.0187669f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.215
cc_17 VNB A3 0.00532635f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.725
cc_18 VNB N_A3_c_265_n 0.0153231f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.215
cc_19 VNB N_B2_M1007_g 0.0292071f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.545
cc_20 VNB N_B2_c_304_n 0.0191347f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.215
cc_21 VNB B2 0.00682372f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.725
cc_22 VNB N_B2_c_306_n 0.0159732f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.215
cc_23 VNB N_B1_c_344_n 0.00141645f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.635
cc_24 VNB N_B1_c_345_n 0.0801152f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.71
cc_25 VNB N_B1_c_346_n 0.032003f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.71
cc_26 VNB N_B1_c_347_n 0.0206825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0492713f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.635
cc_28 VNB N_X_c_377_n 0.0201243f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.71
cc_29 VNB N_VPWR_c_395_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=2.12
cc_30 VNB N_VGND_c_432_n 0.0142437f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.635
cc_31 VNB N_VGND_c_433_n 0.0128028f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.725
cc_32 VNB N_VGND_c_434_n 0.0253838f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.545
cc_33 VNB N_VGND_c_435_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.05
cc_34 VNB N_VGND_c_436_n 0.0201223f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=2.12
cc_35 VNB N_VGND_c_437_n 0.0424912f $X=-0.19 $Y=-0.245 $X2=3.065 $Y2=2.12
cc_36 VNB N_VGND_c_438_n 0.243016f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=2.12
cc_37 VNB N_VGND_c_439_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.12
cc_38 VNB N_A_271_85#_c_473_n 0.0202947f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.725
cc_39 VNB N_A_271_85#_c_474_n 0.00280227f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.725
cc_40 VNB N_A_271_85#_c_475_n 0.0209186f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.215
cc_41 VNB N_A_271_85#_c_476_n 0.00237046f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.025
cc_42 VNB N_A_271_85#_c_477_n 0.0132293f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.71
cc_43 VNB N_A_271_85#_c_478_n 0.00251075f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.55
cc_44 VPB N_A_97_309#_M1011_g 0.0273482f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_45 VPB N_A_97_309#_c_91_n 0.0272404f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.05
cc_46 VPB N_A_97_309#_c_92_n 0.0174494f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.215
cc_47 VPB N_A_97_309#_c_87_n 0.00412337f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.71
cc_48 VPB N_A_97_309#_c_94_n 0.0430453f $X=-0.19 $Y=1.655 $X2=2.31 $Y2=2.12
cc_49 VPB N_A_97_309#_c_95_n 0.00104146f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=2.12
cc_50 VPB N_A_97_309#_c_96_n 0.00708705f $X=-0.19 $Y=1.655 $X2=2.465 $Y2=2.55
cc_51 VPB N_A_97_309#_c_97_n 0.0128412f $X=-0.19 $Y=1.655 $X2=3.065 $Y2=2.12
cc_52 VPB N_A_97_309#_c_88_n 0.00294797f $X=-0.19 $Y=1.655 $X2=3.16 $Y2=2.025
cc_53 VPB N_A_97_309#_c_99_n 0.00596531f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=2.12
cc_54 VPB N_A1_c_171_n 0.0191322f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A1_M1003_g 0.0216981f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.635
cc_56 VPB N_A1_c_168_n 0.011004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A1_c_174_n 0.0207693f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.05
cc_58 VPB A1 0.00326993f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.025
cc_59 VPB N_A2_M1009_g 0.0378807f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.545
cc_60 VPB N_A2_c_220_n 0.0020994f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.215
cc_61 VPB N_A2_c_225_n 0.0153256f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_62 VPB A2 0.00365248f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_63 VPB N_A3_M1002_g 0.0395319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A3_c_263_n 0.00209893f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.215
cc_65 VPB N_A3_c_268_n 0.0151302f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_66 VPB A3 0.00295604f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_67 VPB N_B2_M1004_g 0.040982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_B2_c_304_n 0.00214006f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.215
cc_69 VPB N_B2_c_309_n 0.0153155f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_70 VPB B2 0.00322702f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_71 VPB N_B1_M1008_g 0.0250866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B1_c_344_n 0.0229892f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.635
cc_73 VPB N_B1_c_350_n 0.0237823f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_74 VPB N_B1_c_346_n 0.0352682f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.71
cc_75 VPB X 0.0404321f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.635
cc_76 VPB X 0.044603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_396_n 0.010379f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.635
cc_78 VPB N_VPWR_c_397_n 0.0353933f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.725
cc_79 VPB N_VPWR_c_398_n 0.0569131f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.545
cc_80 VPB N_VPWR_c_399_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.05
cc_81 VPB N_VPWR_c_400_n 0.0258564f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.71
cc_82 VPB N_VPWR_c_401_n 0.013281f $X=-0.19 $Y=1.655 $X2=3.065 $Y2=2.12
cc_83 VPB N_VPWR_c_395_n 0.0994729f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=2.12
cc_84 VPB N_VPWR_c_403_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=2.12
cc_85 N_A_97_309#_M1000_g N_A1_M1005_g 0.0172682f $X=0.71 $Y=0.635 $X2=0 $Y2=0
cc_86 N_A_97_309#_c_91_n N_A1_c_171_n 0.00760762f $X=0.65 $Y=2.05 $X2=0 $Y2=0
cc_87 N_A_97_309#_c_86_n N_A1_c_171_n 0.00108052f $X=0.65 $Y=1.71 $X2=0 $Y2=0
cc_88 N_A_97_309#_c_94_n N_A1_c_171_n 0.00727025f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_89 N_A_97_309#_M1011_g N_A1_M1003_g 0.0148973f $X=0.74 $Y=2.725 $X2=0 $Y2=0
cc_90 N_A_97_309#_c_86_n N_A1_c_167_n 2.35974e-19 $X=0.65 $Y=1.71 $X2=0 $Y2=0
cc_91 N_A_97_309#_c_87_n N_A1_c_167_n 0.00637638f $X=0.65 $Y=1.71 $X2=0 $Y2=0
cc_92 N_A_97_309#_c_91_n N_A1_c_168_n 0.00637638f $X=0.65 $Y=2.05 $X2=0 $Y2=0
cc_93 N_A_97_309#_c_94_n N_A1_c_168_n 9.65567e-19 $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_94 N_A_97_309#_c_92_n N_A1_c_174_n 0.00760762f $X=0.65 $Y=2.215 $X2=0 $Y2=0
cc_95 N_A_97_309#_c_94_n N_A1_c_174_n 0.0196523f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_96 N_A_97_309#_M1000_g A1 0.00732287f $X=0.71 $Y=0.635 $X2=0 $Y2=0
cc_97 N_A_97_309#_c_86_n A1 0.0238951f $X=0.65 $Y=1.71 $X2=0 $Y2=0
cc_98 N_A_97_309#_c_87_n A1 0.00196428f $X=0.65 $Y=1.71 $X2=0 $Y2=0
cc_99 N_A_97_309#_c_94_n A1 0.024701f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_100 N_A_97_309#_M1000_g N_A1_c_170_n 0.0232505f $X=0.71 $Y=0.635 $X2=0 $Y2=0
cc_101 N_A_97_309#_c_94_n N_A2_M1009_g 0.0171813f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_102 N_A_97_309#_c_94_n N_A2_c_225_n 0.00126277f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_103 N_A_97_309#_c_94_n A2 0.0292138f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_104 N_A_97_309#_c_94_n N_A3_M1002_g 0.0160188f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_105 N_A_97_309#_c_96_n N_A3_M1002_g 0.00635995f $X=2.465 $Y=2.55 $X2=0 $Y2=0
cc_106 N_A_97_309#_c_94_n N_A3_c_268_n 3.83682e-19 $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_107 N_A_97_309#_c_99_n N_A3_c_268_n 0.00426331f $X=2.475 $Y=2.12 $X2=0 $Y2=0
cc_108 N_A_97_309#_c_94_n A3 0.0234525f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_109 N_A_97_309#_c_99_n A3 0.00391861f $X=2.475 $Y=2.12 $X2=0 $Y2=0
cc_110 N_A_97_309#_c_96_n N_B2_M1004_g 0.00596323f $X=2.465 $Y=2.55 $X2=0 $Y2=0
cc_111 N_A_97_309#_c_97_n N_B2_M1004_g 0.0164069f $X=3.065 $Y=2.12 $X2=0 $Y2=0
cc_112 N_A_97_309#_c_88_n N_B2_M1004_g 0.00336779f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_113 N_A_97_309#_c_88_n N_B2_M1007_g 0.0048906f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_114 N_A_97_309#_c_89_n N_B2_M1007_g 0.0013975f $X=3.075 $Y=0.69 $X2=0 $Y2=0
cc_115 N_A_97_309#_c_97_n N_B2_c_309_n 0.00406107f $X=3.065 $Y=2.12 $X2=0 $Y2=0
cc_116 N_A_97_309#_c_97_n B2 0.0198529f $X=3.065 $Y=2.12 $X2=0 $Y2=0
cc_117 N_A_97_309#_c_88_n B2 0.0511475f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_118 N_A_97_309#_c_99_n B2 0.0106696f $X=2.475 $Y=2.12 $X2=0 $Y2=0
cc_119 N_A_97_309#_c_88_n N_B2_c_306_n 0.00450394f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_120 N_A_97_309#_c_89_n N_B2_c_306_n 0.00235548f $X=3.075 $Y=0.69 $X2=0 $Y2=0
cc_121 N_A_97_309#_c_97_n N_B1_c_344_n 0.00190538f $X=3.065 $Y=2.12 $X2=0 $Y2=0
cc_122 N_A_97_309#_c_88_n N_B1_c_344_n 0.00788472f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_123 N_A_97_309#_c_97_n N_B1_c_350_n 0.0193818f $X=3.065 $Y=2.12 $X2=0 $Y2=0
cc_124 N_A_97_309#_c_88_n N_B1_c_345_n 0.0165531f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_125 N_A_97_309#_c_97_n N_B1_c_346_n 0.0079288f $X=3.065 $Y=2.12 $X2=0 $Y2=0
cc_126 N_A_97_309#_c_88_n N_B1_c_346_n 0.078602f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_127 N_A_97_309#_c_88_n N_B1_c_347_n 0.00499845f $X=3.16 $Y=2.025 $X2=0 $Y2=0
cc_128 N_A_97_309#_c_89_n N_B1_c_347_n 0.00594149f $X=3.075 $Y=0.69 $X2=0 $Y2=0
cc_129 N_A_97_309#_M1000_g X 0.0163415f $X=0.71 $Y=0.635 $X2=0 $Y2=0
cc_130 N_A_97_309#_M1011_g X 0.00572509f $X=0.74 $Y=2.725 $X2=0 $Y2=0
cc_131 N_A_97_309#_c_86_n X 0.0369789f $X=0.65 $Y=1.71 $X2=0 $Y2=0
cc_132 N_A_97_309#_c_87_n X 0.0165074f $X=0.65 $Y=1.71 $X2=0 $Y2=0
cc_133 N_A_97_309#_c_95_n X 0.0157867f $X=0.815 $Y=2.12 $X2=0 $Y2=0
cc_134 N_A_97_309#_M1011_g X 0.00917925f $X=0.74 $Y=2.725 $X2=0 $Y2=0
cc_135 N_A_97_309#_c_92_n X 0.0041452f $X=0.65 $Y=2.215 $X2=0 $Y2=0
cc_136 N_A_97_309#_c_95_n X 0.0113042f $X=0.815 $Y=2.12 $X2=0 $Y2=0
cc_137 N_A_97_309#_M1011_g N_VPWR_c_396_n 0.00970149f $X=0.74 $Y=2.725 $X2=0
+ $Y2=0
cc_138 N_A_97_309#_c_94_n N_VPWR_c_396_n 0.0277457f $X=2.31 $Y=2.12 $X2=0 $Y2=0
cc_139 N_A_97_309#_c_96_n N_VPWR_c_397_n 0.0109443f $X=2.465 $Y=2.55 $X2=0 $Y2=0
cc_140 N_A_97_309#_c_97_n N_VPWR_c_397_n 0.00791465f $X=3.065 $Y=2.12 $X2=0
+ $Y2=0
cc_141 N_A_97_309#_c_96_n N_VPWR_c_398_n 0.0235133f $X=2.465 $Y=2.55 $X2=0 $Y2=0
cc_142 N_A_97_309#_M1011_g N_VPWR_c_400_n 0.00502664f $X=0.74 $Y=2.725 $X2=0
+ $Y2=0
cc_143 N_A_97_309#_M1011_g N_VPWR_c_395_n 0.0106697f $X=0.74 $Y=2.725 $X2=0
+ $Y2=0
cc_144 N_A_97_309#_c_96_n N_VPWR_c_395_n 0.0127519f $X=2.465 $Y=2.55 $X2=0 $Y2=0
cc_145 N_A_97_309#_M1000_g N_VGND_c_432_n 0.00526406f $X=0.71 $Y=0.635 $X2=0
+ $Y2=0
cc_146 N_A_97_309#_M1000_g N_VGND_c_434_n 0.00537957f $X=0.71 $Y=0.635 $X2=0
+ $Y2=0
cc_147 N_A_97_309#_M1000_g N_VGND_c_438_n 0.00528353f $X=0.71 $Y=0.635 $X2=0
+ $Y2=0
cc_148 N_A_97_309#_c_88_n N_A_271_85#_c_473_n 0.00766724f $X=3.16 $Y=2.025 $X2=0
+ $Y2=0
cc_149 N_A_97_309#_c_89_n N_A_271_85#_c_473_n 6.47229e-19 $X=3.075 $Y=0.69 $X2=0
+ $Y2=0
cc_150 N_A_97_309#_c_89_n N_A_271_85#_c_475_n 0.0225397f $X=3.075 $Y=0.69 $X2=0
+ $Y2=0
cc_151 N_A1_M1005_g N_A2_M1010_g 0.0243943f $X=1.28 $Y=0.635 $X2=0 $Y2=0
cc_152 A1 N_A2_M1010_g 0.00107237f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_153 N_A1_c_171_n N_A2_M1009_g 0.00838486f $X=1.28 $Y=2.095 $X2=0 $Y2=0
cc_154 N_A1_c_174_n N_A2_M1009_g 0.0602161f $X=1.43 $Y=2.17 $X2=0 $Y2=0
cc_155 N_A1_c_167_n N_A2_c_220_n 0.013709f $X=1.19 $Y=1.585 $X2=0 $Y2=0
cc_156 N_A1_c_168_n N_A2_c_225_n 0.013709f $X=1.19 $Y=1.75 $X2=0 $Y2=0
cc_157 A1 A2 0.0478f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_158 N_A1_c_170_n A2 0.00436559f $X=1.19 $Y=1.245 $X2=0 $Y2=0
cc_159 A1 N_A2_c_222_n 6.3994e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_160 N_A1_c_170_n N_A2_c_222_n 0.013709f $X=1.19 $Y=1.245 $X2=0 $Y2=0
cc_161 A1 X 0.023822f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_162 N_A1_M1003_g N_VPWR_c_396_n 0.0217917f $X=1.43 $Y=2.725 $X2=0 $Y2=0
cc_163 N_A1_c_174_n N_VPWR_c_396_n 0.00124205f $X=1.43 $Y=2.17 $X2=0 $Y2=0
cc_164 N_A1_M1003_g N_VPWR_c_398_n 0.0053602f $X=1.43 $Y=2.725 $X2=0 $Y2=0
cc_165 N_A1_M1003_g N_VPWR_c_395_n 0.0107416f $X=1.43 $Y=2.725 $X2=0 $Y2=0
cc_166 A1 N_VGND_M1000_d 0.00184152f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_167 N_A1_M1005_g N_VGND_c_432_n 0.00450927f $X=1.28 $Y=0.635 $X2=0 $Y2=0
cc_168 A1 N_VGND_c_432_n 0.0142542f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_169 N_A1_c_170_n N_VGND_c_432_n 5.91804e-19 $X=1.19 $Y=1.245 $X2=0 $Y2=0
cc_170 N_A1_M1005_g N_VGND_c_436_n 0.00512663f $X=1.28 $Y=0.635 $X2=0 $Y2=0
cc_171 N_A1_M1005_g N_VGND_c_438_n 0.00528353f $X=1.28 $Y=0.635 $X2=0 $Y2=0
cc_172 A1 N_VGND_c_438_n 0.0052491f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_173 N_A1_M1005_g N_A_271_85#_c_482_n 0.00363428f $X=1.28 $Y=0.635 $X2=0 $Y2=0
cc_174 A1 N_A_271_85#_c_482_n 3.18716e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_175 N_A1_M1005_g N_A_271_85#_c_474_n 0.00125742f $X=1.28 $Y=0.635 $X2=0 $Y2=0
cc_176 A1 N_A_271_85#_c_474_n 0.0136424f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_177 N_A1_M1005_g N_A_271_85#_c_478_n 0.00476129f $X=1.28 $Y=0.635 $X2=0 $Y2=0
cc_178 N_A2_M1009_g N_A3_M1002_g 0.0725776f $X=1.82 $Y=2.725 $X2=0 $Y2=0
cc_179 N_A2_M1010_g N_A3_M1001_g 0.0173143f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_180 N_A2_c_220_n N_A3_c_263_n 0.0138263f $X=1.73 $Y=1.69 $X2=0 $Y2=0
cc_181 N_A2_c_225_n N_A3_c_268_n 0.0138263f $X=1.73 $Y=1.855 $X2=0 $Y2=0
cc_182 A2 A3 0.0534605f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A2_c_222_n A3 0.00418101f $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_184 A2 N_A3_c_265_n 6.43261e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A2_c_222_n N_A3_c_265_n 0.0138263f $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_186 N_A2_M1009_g N_VPWR_c_398_n 0.0053602f $X=1.82 $Y=2.725 $X2=0 $Y2=0
cc_187 N_A2_M1009_g N_VPWR_c_395_n 0.0103235f $X=1.82 $Y=2.725 $X2=0 $Y2=0
cc_188 N_A2_M1010_g N_VGND_c_433_n 0.00555102f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_189 N_A2_M1010_g N_VGND_c_436_n 0.00512663f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_190 N_A2_M1010_g N_VGND_c_438_n 0.00528353f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_191 N_A2_M1010_g N_A_271_85#_c_482_n 0.00440123f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_192 N_A2_M1010_g N_A_271_85#_c_473_n 0.00945922f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_193 A2 N_A_271_85#_c_473_n 0.0141854f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A2_c_222_n N_A_271_85#_c_473_n 0.00252718f $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_195 N_A2_M1010_g N_A_271_85#_c_474_n 0.00207186f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_196 A2 N_A_271_85#_c_474_n 0.0154106f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A2_c_222_n N_A_271_85#_c_474_n 5.15248e-19 $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_198 N_A2_M1010_g N_A_271_85#_c_494_n 7.9267e-19 $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_199 N_A2_M1010_g N_A_271_85#_c_478_n 0.00400827f $X=1.71 $Y=0.635 $X2=0 $Y2=0
cc_200 N_A3_M1002_g N_B2_M1004_g 0.0220837f $X=2.21 $Y=2.725 $X2=0 $Y2=0
cc_201 N_A3_M1001_g N_B2_M1007_g 0.0218736f $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_202 N_A3_c_263_n N_B2_c_304_n 0.0137828f $X=2.27 $Y=1.69 $X2=0 $Y2=0
cc_203 N_A3_c_268_n N_B2_c_309_n 0.0137828f $X=2.27 $Y=1.855 $X2=0 $Y2=0
cc_204 A3 B2 0.053544f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_205 N_A3_c_265_n B2 0.00448642f $X=2.27 $Y=1.35 $X2=0 $Y2=0
cc_206 A3 N_B2_c_306_n 5.83318e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_207 N_A3_c_265_n N_B2_c_306_n 0.0137828f $X=2.27 $Y=1.35 $X2=0 $Y2=0
cc_208 N_A3_M1002_g N_VPWR_c_398_n 0.0053602f $X=2.21 $Y=2.725 $X2=0 $Y2=0
cc_209 N_A3_M1002_g N_VPWR_c_395_n 0.0105184f $X=2.21 $Y=2.725 $X2=0 $Y2=0
cc_210 N_A3_M1001_g N_VGND_c_433_n 0.00385401f $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_211 N_A3_M1001_g N_VGND_c_437_n 0.00462669f $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_212 N_A3_M1001_g N_VGND_c_438_n 0.00440294f $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_213 N_A3_M1001_g N_A_271_85#_c_482_n 7.4574e-19 $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_214 N_A3_M1001_g N_A_271_85#_c_473_n 0.0144375f $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_215 A3 N_A_271_85#_c_473_n 0.0271251f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_216 N_A3_c_265_n N_A_271_85#_c_473_n 0.00125222f $X=2.27 $Y=1.35 $X2=0 $Y2=0
cc_217 N_A3_M1001_g N_A_271_85#_c_494_n 0.00666911f $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_218 N_A3_M1001_g N_A_271_85#_c_476_n 0.00337159f $X=2.36 $Y=0.635 $X2=0 $Y2=0
cc_219 N_B2_M1004_g N_B1_c_344_n 0.00574715f $X=2.72 $Y=2.725 $X2=0 $Y2=0
cc_220 N_B2_c_304_n N_B1_c_344_n 0.0174123f $X=2.81 $Y=1.69 $X2=0 $Y2=0
cc_221 N_B2_M1004_g N_B1_c_350_n 0.0553792f $X=2.72 $Y=2.725 $X2=0 $Y2=0
cc_222 B2 N_B1_c_345_n 5.6994e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_223 N_B2_c_306_n N_B1_c_345_n 0.0174123f $X=2.81 $Y=1.35 $X2=0 $Y2=0
cc_224 N_B2_M1007_g N_B1_c_347_n 0.0215952f $X=2.79 $Y=0.635 $X2=0 $Y2=0
cc_225 N_B2_M1004_g N_VPWR_c_397_n 0.00273386f $X=2.72 $Y=2.725 $X2=0 $Y2=0
cc_226 N_B2_M1004_g N_VPWR_c_398_n 0.0053602f $X=2.72 $Y=2.725 $X2=0 $Y2=0
cc_227 N_B2_M1004_g N_VPWR_c_395_n 0.0105184f $X=2.72 $Y=2.725 $X2=0 $Y2=0
cc_228 N_B2_M1007_g N_VGND_c_437_n 8.63546e-19 $X=2.79 $Y=0.635 $X2=0 $Y2=0
cc_229 N_B2_M1007_g N_A_271_85#_c_473_n 0.00212009f $X=2.79 $Y=0.635 $X2=0 $Y2=0
cc_230 B2 N_A_271_85#_c_473_n 0.0142547f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_231 N_B2_c_306_n N_A_271_85#_c_473_n 2.73709e-19 $X=2.81 $Y=1.35 $X2=0 $Y2=0
cc_232 N_B2_M1007_g N_A_271_85#_c_475_n 0.0139698f $X=2.79 $Y=0.635 $X2=0 $Y2=0
cc_233 N_B1_M1008_g N_VPWR_c_397_n 0.017337f $X=3.11 $Y=2.725 $X2=0 $Y2=0
cc_234 N_B1_c_350_n N_VPWR_c_397_n 0.00717923f $X=3.29 $Y=2.17 $X2=0 $Y2=0
cc_235 N_B1_c_346_n N_VPWR_c_397_n 0.00421198f $X=3.51 $Y=1.12 $X2=0 $Y2=0
cc_236 N_B1_M1008_g N_VPWR_c_398_n 0.00445056f $X=3.11 $Y=2.725 $X2=0 $Y2=0
cc_237 N_B1_M1008_g N_VPWR_c_395_n 0.00804604f $X=3.11 $Y=2.725 $X2=0 $Y2=0
cc_238 N_B1_c_347_n N_VGND_c_437_n 8.63546e-19 $X=3.445 $Y=0.955 $X2=0 $Y2=0
cc_239 N_B1_c_345_n N_A_271_85#_c_475_n 0.001399f $X=3.51 $Y=1.12 $X2=0 $Y2=0
cc_240 N_B1_c_347_n N_A_271_85#_c_475_n 0.0139359f $X=3.445 $Y=0.955 $X2=0 $Y2=0
cc_241 N_B1_c_345_n N_A_271_85#_c_477_n 0.00218094f $X=3.51 $Y=1.12 $X2=0 $Y2=0
cc_242 N_B1_c_346_n N_A_271_85#_c_477_n 0.0208651f $X=3.51 $Y=1.12 $X2=0 $Y2=0
cc_243 X N_VPWR_c_396_n 3.52044e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_244 X N_VPWR_c_396_n 0.0432003f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_245 X N_VPWR_c_400_n 0.0405511f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_246 X N_VPWR_c_395_n 0.0232167f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_247 N_X_c_377_n N_VGND_c_434_n 0.0141468f $X=0.495 $Y=0.635 $X2=0 $Y2=0
cc_248 N_X_c_377_n N_VGND_c_438_n 0.0170907f $X=0.495 $Y=0.635 $X2=0 $Y2=0
cc_249 N_VGND_c_433_n N_A_271_85#_c_482_n 3.17622e-19 $X=2.035 $Y=0.565 $X2=0
+ $Y2=0
cc_250 N_VGND_c_433_n N_A_271_85#_c_473_n 0.0265277f $X=2.035 $Y=0.565 $X2=0
+ $Y2=0
cc_251 N_VGND_c_438_n N_A_271_85#_c_473_n 0.0146958f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_433_n N_A_271_85#_c_494_n 0.0162247f $X=2.035 $Y=0.565 $X2=0
+ $Y2=0
cc_253 N_VGND_c_437_n N_A_271_85#_c_475_n 0.0652324f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_438_n N_A_271_85#_c_475_n 0.0374769f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_433_n N_A_271_85#_c_476_n 0.0123474f $X=2.035 $Y=0.565 $X2=0
+ $Y2=0
cc_256 N_VGND_c_437_n N_A_271_85#_c_476_n 0.0193554f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_438_n N_A_271_85#_c_476_n 0.010497f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_432_n N_A_271_85#_c_478_n 0.0122667f $X=0.995 $Y=0.55 $X2=0
+ $Y2=0
cc_259 N_VGND_c_433_n N_A_271_85#_c_478_n 0.0188107f $X=2.035 $Y=0.565 $X2=0
+ $Y2=0
cc_260 N_VGND_c_436_n N_A_271_85#_c_478_n 0.0119695f $X=1.87 $Y=0 $X2=0 $Y2=0
cc_261 N_VGND_c_438_n N_A_271_85#_c_478_n 0.0115266f $X=3.6 $Y=0 $X2=0 $Y2=0
