# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__and4bb_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__and4bb_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.785000 1.315000 1.455000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.560000 1.125000 1.890000 1.455000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 1.120000 3.715000 1.790000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.940000 1.120000 4.270000 1.790000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.800000 1.920000 5.190000 3.065000 ;
        RECT 4.815000 0.265000 5.190000 0.675000 ;
        RECT 5.020000 0.675000 5.190000 1.920000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
        RECT 0.905000  0.085000 1.235000 0.605000 ;
        RECT 3.885000  0.085000 4.215000 0.590000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.280000 3.415000 ;
        RECT 0.645000 1.985000 0.975000 3.245000 ;
        RECT 1.965000 2.335000 2.295000 3.245000 ;
        RECT 3.025000 2.685000 3.355000 3.245000 ;
        RECT 4.165000 2.320000 4.495000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.265000 0.445000 1.635000 ;
      RECT 0.115000 1.635000 2.560000 1.805000 ;
      RECT 0.115000 1.805000 0.445000 3.025000 ;
      RECT 1.435000 1.985000 2.970000 2.155000 ;
      RECT 1.435000 2.155000 1.765000 3.065000 ;
      RECT 1.725000 0.265000 2.055000 0.775000 ;
      RECT 1.725000 0.775000 2.970000 0.945000 ;
      RECT 2.230000 1.135000 2.560000 1.635000 ;
      RECT 2.285000 0.265000 3.480000 0.595000 ;
      RECT 2.495000 2.335000 3.965000 2.505000 ;
      RECT 2.495000 2.505000 2.825000 3.065000 ;
      RECT 2.800000 0.945000 2.970000 1.215000 ;
      RECT 2.800000 1.215000 3.130000 1.885000 ;
      RECT 2.800000 1.885000 2.970000 1.985000 ;
      RECT 3.310000 0.595000 3.480000 0.770000 ;
      RECT 3.310000 0.770000 4.620000 0.940000 ;
      RECT 3.635000 1.970000 4.620000 2.140000 ;
      RECT 3.635000 2.140000 3.965000 2.335000 ;
      RECT 3.635000 2.505000 3.965000 3.065000 ;
      RECT 4.450000 0.940000 4.840000 1.610000 ;
      RECT 4.450000 1.610000 4.620000 1.970000 ;
  END
END sky130_fd_sc_lp__and4bb_lp
