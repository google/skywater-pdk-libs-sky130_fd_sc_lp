* File: sky130_fd_sc_lp__a211o_2.pxi.spice
* Created: Wed Sep  2 09:17:33 2020
* 
x_PM_SKY130_FD_SC_LP__A211O_2%A_80_21# N_A_80_21#_M1007_d N_A_80_21#_M1001_d
+ N_A_80_21#_M1006_d N_A_80_21#_M1002_g N_A_80_21#_M1003_g N_A_80_21#_M1004_g
+ N_A_80_21#_M1011_g N_A_80_21#_c_60_n N_A_80_21#_c_72_p N_A_80_21#_c_140_p
+ N_A_80_21#_c_67_n N_A_80_21#_c_94_p N_A_80_21#_c_61_n N_A_80_21#_c_68_n
+ N_A_80_21#_c_62_n N_A_80_21#_c_63_n N_A_80_21#_c_64_n N_A_80_21#_c_89_p
+ PM_SKY130_FD_SC_LP__A211O_2%A_80_21#
x_PM_SKY130_FD_SC_LP__A211O_2%A2 N_A2_c_165_n N_A2_M1005_g N_A2_M1009_g A2
+ N_A2_c_168_n PM_SKY130_FD_SC_LP__A211O_2%A2
x_PM_SKY130_FD_SC_LP__A211O_2%A1 N_A1_M1007_g N_A1_M1000_g A1 N_A1_c_203_n
+ N_A1_c_204_n N_A1_c_205_n PM_SKY130_FD_SC_LP__A211O_2%A1
x_PM_SKY130_FD_SC_LP__A211O_2%B1 N_B1_M1010_g N_B1_M1008_g B1 N_B1_c_241_n
+ N_B1_c_242_n PM_SKY130_FD_SC_LP__A211O_2%B1
x_PM_SKY130_FD_SC_LP__A211O_2%C1 N_C1_c_271_n N_C1_M1001_g N_C1_M1006_g C1
+ N_C1_c_274_n PM_SKY130_FD_SC_LP__A211O_2%C1
x_PM_SKY130_FD_SC_LP__A211O_2%VPWR N_VPWR_M1003_d N_VPWR_M1011_d N_VPWR_M1009_d
+ N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n VPWR
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_294_n N_VPWR_c_303_n
+ N_VPWR_c_304_n PM_SKY130_FD_SC_LP__A211O_2%VPWR
x_PM_SKY130_FD_SC_LP__A211O_2%X N_X_M1002_d N_X_M1003_s X X X X X X X
+ N_X_c_344_n PM_SKY130_FD_SC_LP__A211O_2%X
x_PM_SKY130_FD_SC_LP__A211O_2%A_303_367# N_A_303_367#_M1009_s
+ N_A_303_367#_M1000_d N_A_303_367#_c_361_n N_A_303_367#_c_362_n
+ N_A_303_367#_c_366_n N_A_303_367#_c_367_n N_A_303_367#_c_371_n
+ PM_SKY130_FD_SC_LP__A211O_2%A_303_367#
x_PM_SKY130_FD_SC_LP__A211O_2%VGND N_VGND_M1002_s N_VGND_M1004_s N_VGND_M1010_d
+ N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n VGND N_VGND_c_391_n
+ N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n
+ PM_SKY130_FD_SC_LP__A211O_2%VGND
cc_1 VNB N_A_80_21#_M1002_g 0.0343508f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_80_21#_M1004_g 0.0290292f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_3 VNB N_A_80_21#_c_60_n 0.0050953f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.345
cc_4 VNB N_A_80_21#_c_61_n 0.00740447f $X=-0.19 $Y=-0.245 $X2=3.415 $Y2=0.94
cc_5 VNB N_A_80_21#_c_62_n 0.0228289f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=0.42
cc_6 VNB N_A_80_21#_c_63_n 0.00685481f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.51
cc_7 VNB N_A_80_21#_c_64_n 0.062015f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.51
cc_8 VNB N_A2_c_165_n 0.0190198f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=0.235
cc_9 VNB N_A2_M1009_g 0.00842767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A2 0.00359873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_168_n 0.0419046f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.675
cc_12 VNB N_A1_M1000_g 0.00834293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_203_n 0.0276981f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_14 VNB N_A1_c_204_n 0.00633449f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_15 VNB N_A1_c_205_n 0.0177129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_M1008_g 0.00774559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB B1 0.0080088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_241_n 0.0271379f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_19 VNB N_B1_c_242_n 0.0181648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C1_c_271_n 0.022077f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=0.235
cc_21 VNB N_C1_M1006_g 0.0113687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB C1 0.019205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_c_274_n 0.0516691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_294_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=0.855
cc_25 VNB N_X_c_344_n 0.00553032f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.675
cc_26 VNB N_VGND_c_388_n 0.0108094f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.345
cc_27 VNB N_VGND_c_389_n 0.0493808f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_28 VNB N_VGND_c_390_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_29 VNB N_VGND_c_391_n 0.0300736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_392_n 0.0176034f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=0.855
cc_31 VNB N_VGND_c_393_n 0.210926f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=0.42
cc_32 VNB N_VGND_c_394_n 0.0168265f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.95
cc_33 VNB N_VGND_c_395_n 0.0192665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_396_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.51
cc_35 VPB N_A_80_21#_M1003_g 0.0255346f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_36 VPB N_A_80_21#_M1011_g 0.0223364f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_37 VPB N_A_80_21#_c_67_n 0.0265637f $X=-0.19 $Y=1.655 $X2=3.345 $Y2=1.785
cc_38 VPB N_A_80_21#_c_68_n 0.0466985f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=1.98
cc_39 VPB N_A_80_21#_c_63_n 0.0108234f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.51
cc_40 VPB N_A_80_21#_c_64_n 0.0149297f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.51
cc_41 VPB N_A2_M1009_g 0.0250477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A1_M1000_g 0.0206821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_B1_M1008_g 0.0193402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_C1_M1006_g 0.0245806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_295_n 0.0107835f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.345
cc_46 VPB N_VPWR_c_296_n 0.0653952f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_47 VPB N_VPWR_c_297_n 0.0139719f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.345
cc_48 VPB N_VPWR_c_298_n 0.00500416f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_49 VPB N_VPWR_c_299_n 0.0169856f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=0.94
cc_50 VPB N_VPWR_c_300_n 0.0183524f $X=-0.19 $Y=1.655 $X2=2.53 $Y2=0.42
cc_51 VPB N_VPWR_c_301_n 0.0452282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_294_n 0.0553268f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=0.855
cc_53 VPB N_VPWR_c_303_n 0.00545601f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.51
cc_54 VPB N_VPWR_c_304_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.51
cc_55 VPB N_X_c_344_n 0.00271355f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.675
cc_56 VPB N_A_303_367#_c_361_n 0.00200389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_303_367#_c_362_n 0.00786051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 N_A_80_21#_c_60_n N_A2_c_165_n 0.00470358f $X=1.33 $Y=1.345 $X2=-0.19
+ $Y2=-0.245
cc_59 N_A_80_21#_c_72_p N_A2_c_165_n 0.0144148f $X=2.365 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_60 N_A_80_21#_c_67_n N_A2_M1009_g 0.0146303f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_63_n N_A2_M1009_g 0.0037459f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_64_n N_A2_M1009_g 0.00265087f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_60_n A2 0.011033f $X=1.33 $Y=1.345 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_72_p A2 0.0169121f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_67_n A2 0.0193299f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_63_n A2 0.0143345f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_67 N_A_80_21#_M1004_g N_A2_c_168_n 0.00220312f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_60_n N_A2_c_168_n 0.00163046f $X=1.33 $Y=1.345 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_72_p N_A2_c_168_n 0.00318472f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_67_n N_A2_c_168_n 0.00332142f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_63_n N_A2_c_168_n 0.00133262f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_64_n N_A2_c_168_n 0.00933058f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_67_n N_A1_M1000_g 0.0117401f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_72_p N_A1_c_203_n 0.00175077f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_67_n N_A1_c_203_n 0.00459984f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_89_p N_A1_c_203_n 0.00289427f $X=2.53 $Y=0.94 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_72_p N_A1_c_204_n 0.0217535f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_67_n N_A1_c_204_n 0.0327696f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_89_p N_A1_c_204_n 0.00865234f $X=2.53 $Y=0.94 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_72_p N_A1_c_205_n 0.0125365f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_94_p N_A1_c_205_n 0.0114639f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_67_n N_B1_M1008_g 0.0156967f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_68_n N_B1_M1008_g 0.00390041f $X=3.51 $Y=1.98 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_67_n B1 0.0388724f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_61_n B1 0.0327152f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_89_p B1 0.00123605f $X=2.53 $Y=0.94 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_67_n N_B1_c_241_n 0.00405418f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_61_n N_B1_c_241_n 0.00352542f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_89_p N_B1_c_241_n 3.53661e-19 $X=2.53 $Y=0.94 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_94_p N_B1_c_242_n 0.00912539f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_61_n N_B1_c_242_n 0.0127338f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_61_n N_C1_c_271_n 0.0119242f $X=3.415 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_80_21#_c_67_n N_C1_M1006_g 0.0170761f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_68_n N_C1_M1006_g 0.0254485f $X=3.51 $Y=1.98 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_67_n C1 0.0234044f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_61_n C1 0.0210616f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_67_n N_C1_c_274_n 0.00274682f $X=3.345 $Y=1.785 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_61_n N_C1_c_274_n 0.00608861f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_63_n N_VPWR_M1011_d 5.31253e-19 $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_67_n N_VPWR_M1009_d 0.00301104f $X=3.345 $Y=1.785 $X2=0
+ $Y2=0
cc_101 N_A_80_21#_M1003_g N_VPWR_c_296_n 0.00769005f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_102 N_A_80_21#_M1011_g N_VPWR_c_297_n 0.00338373f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_A_80_21#_c_63_n N_VPWR_c_297_n 0.0138487f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_64_n N_VPWR_c_297_n 0.00171668f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A_80_21#_M1003_g N_VPWR_c_299_n 0.00585385f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_106 N_A_80_21#_M1011_g N_VPWR_c_299_n 0.00585385f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_107 N_A_80_21#_c_68_n N_VPWR_c_301_n 0.0210467f $X=3.51 $Y=1.98 $X2=0 $Y2=0
cc_108 N_A_80_21#_M1006_d N_VPWR_c_294_n 0.00215158f $X=3.37 $Y=1.835 $X2=0
+ $Y2=0
cc_109 N_A_80_21#_M1003_g N_VPWR_c_294_n 0.0114687f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_80_21#_M1011_g N_VPWR_c_294_n 0.0118494f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_c_68_n N_VPWR_c_294_n 0.0125689f $X=3.51 $Y=1.98 $X2=0 $Y2=0
cc_112 N_A_80_21#_M1002_g N_X_c_344_n 0.00768412f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_113 N_A_80_21#_M1003_g N_X_c_344_n 0.0047449f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_80_21#_M1004_g N_X_c_344_n 0.00387303f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_115 N_A_80_21#_M1011_g N_X_c_344_n 0.00264273f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_60_n N_X_c_344_n 0.012097f $X=1.33 $Y=1.345 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_63_n N_X_c_344_n 0.0326026f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_64_n N_X_c_344_n 0.0312522f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_67_n N_A_303_367#_M1009_s 0.00239847f $X=3.345 $Y=1.785
+ $X2=-0.19 $Y2=-0.245
cc_120 N_A_80_21#_c_67_n N_A_303_367#_M1000_d 0.00230018f $X=3.345 $Y=1.785
+ $X2=0 $Y2=0
cc_121 N_A_80_21#_c_67_n N_A_303_367#_c_361_n 0.0211022f $X=3.345 $Y=1.785 $X2=0
+ $Y2=0
cc_122 N_A_80_21#_c_67_n N_A_303_367#_c_366_n 0.0392973f $X=3.345 $Y=1.785 $X2=0
+ $Y2=0
cc_123 N_A_80_21#_c_67_n N_A_303_367#_c_367_n 0.0183639f $X=3.345 $Y=1.785 $X2=0
+ $Y2=0
cc_124 N_A_80_21#_c_67_n A_590_367# 0.00599363f $X=3.345 $Y=1.785 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_80_21#_c_60_n N_VGND_M1004_s 0.00172439f $X=1.33 $Y=1.345 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_72_p N_VGND_M1004_s 0.00897332f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_140_p N_VGND_M1004_s 0.00571468f $X=1.415 $Y=0.94 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_c_61_n N_VGND_M1010_d 0.0034814f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_129 N_A_80_21#_M1002_g N_VGND_c_389_n 0.00708134f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_130 N_A_80_21#_c_94_p N_VGND_c_390_n 0.0273795f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_131 N_A_80_21#_c_61_n N_VGND_c_390_n 0.0167229f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_94_p N_VGND_c_391_n 0.0230625f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_62_n N_VGND_c_392_n 0.0178111f $X=3.51 $Y=0.42 $X2=0 $Y2=0
cc_134 N_A_80_21#_M1007_d N_VGND_c_393_n 0.00521751f $X=2.29 $Y=0.235 $X2=0
+ $Y2=0
cc_135 N_A_80_21#_M1001_d N_VGND_c_393_n 0.00244525f $X=3.37 $Y=0.235 $X2=0
+ $Y2=0
cc_136 N_A_80_21#_M1002_g N_VGND_c_393_n 0.0114687f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_137 N_A_80_21#_M1004_g N_VGND_c_393_n 0.0120404f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_138 N_A_80_21#_c_72_p N_VGND_c_393_n 0.0183388f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_140_p N_VGND_c_393_n 6.06937e-19 $X=1.415 $Y=0.94 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_c_94_p N_VGND_c_393_n 0.0127519f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_61_n N_VGND_c_393_n 0.0124936f $X=3.415 $Y=0.94 $X2=0 $Y2=0
cc_142 N_A_80_21#_c_62_n N_VGND_c_393_n 0.0100304f $X=3.51 $Y=0.42 $X2=0 $Y2=0
cc_143 N_A_80_21#_M1002_g N_VGND_c_394_n 0.00585385f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_M1004_g N_VGND_c_394_n 0.00585385f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_145 N_A_80_21#_M1004_g N_VGND_c_395_n 0.00533336f $X=0.905 $Y=0.655 $X2=0
+ $Y2=0
cc_146 N_A_80_21#_c_72_p N_VGND_c_395_n 0.0262022f $X=2.365 $Y=0.94 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_140_p N_VGND_c_395_n 0.0149065f $X=1.415 $Y=0.94 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_94_p N_VGND_c_395_n 0.0137979f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_63_n N_VGND_c_395_n 0.00632316f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_64_n N_VGND_c_395_n 0.00140412f $X=1.105 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_72_p A_386_47# 0.00324028f $X=2.365 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A2_c_168_n N_A1_M1000_g 0.0314934f $X=1.855 $Y=1.36 $X2=0 $Y2=0
cc_153 A2 N_A1_c_203_n 2.73465e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A2_c_168_n N_A1_c_203_n 0.0439743f $X=1.855 $Y=1.36 $X2=0 $Y2=0
cc_155 A2 N_A1_c_204_n 0.0255156f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_c_168_n N_A1_c_204_n 0.00226574f $X=1.855 $Y=1.36 $X2=0 $Y2=0
cc_157 N_A2_c_165_n N_A1_c_205_n 0.0439743f $X=1.855 $Y=1.195 $X2=0 $Y2=0
cc_158 N_A2_M1009_g N_VPWR_c_297_n 0.00297399f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A2_M1009_g N_VPWR_c_298_n 0.00216724f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_M1009_g N_VPWR_c_300_n 0.00571722f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A2_M1009_g N_VPWR_c_294_n 0.0118478f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A2_M1009_g N_A_303_367#_c_361_n 2.8301e-19 $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A2_M1009_g N_A_303_367#_c_362_n 0.00969654f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A2_M1009_g N_A_303_367#_c_366_n 0.013103f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A2_M1009_g N_A_303_367#_c_371_n 4.56565e-19 $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A2_c_165_n N_VGND_c_391_n 0.00486043f $X=1.855 $Y=1.195 $X2=0 $Y2=0
cc_167 N_A2_c_165_n N_VGND_c_393_n 0.00446329f $X=1.855 $Y=1.195 $X2=0 $Y2=0
cc_168 N_A2_c_165_n N_VGND_c_395_n 0.0180864f $X=1.855 $Y=1.195 $X2=0 $Y2=0
cc_169 N_A1_M1000_g N_B1_M1008_g 0.0226318f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A1_c_203_n B1 3.99867e-19 $X=2.305 $Y=1.35 $X2=0 $Y2=0
cc_171 N_A1_c_204_n B1 0.0216105f $X=2.305 $Y=1.35 $X2=0 $Y2=0
cc_172 N_A1_c_203_n N_B1_c_241_n 0.0215255f $X=2.305 $Y=1.35 $X2=0 $Y2=0
cc_173 N_A1_c_204_n N_B1_c_241_n 4.00674e-19 $X=2.305 $Y=1.35 $X2=0 $Y2=0
cc_174 N_A1_c_205_n N_B1_c_242_n 0.0205014f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A1_M1000_g N_VPWR_c_298_n 0.00354331f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A1_M1000_g N_VPWR_c_301_n 0.00571847f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A1_M1000_g N_VPWR_c_294_n 0.0106896f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A1_M1000_g N_A_303_367#_c_362_n 4.58929e-19 $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A1_M1000_g N_A_303_367#_c_366_n 0.013103f $X=2.395 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1000_g N_A_303_367#_c_367_n 2.8301e-19 $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A1_M1000_g N_A_303_367#_c_371_n 0.00956591f $X=2.395 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A1_c_205_n N_VGND_c_390_n 9.30626e-19 $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A1_c_205_n N_VGND_c_391_n 0.00585385f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_184 N_A1_c_205_n N_VGND_c_393_n 0.00690449f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_185 N_A1_c_205_n N_VGND_c_395_n 0.00253404f $X=2.305 $Y=1.185 $X2=0 $Y2=0
cc_186 N_B1_c_242_n N_C1_c_271_n 0.0316642f $X=2.845 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_187 N_B1_M1008_g N_C1_M1006_g 0.0776565f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_188 B1 C1 0.0265002f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 N_B1_c_241_n C1 2.14743e-19 $X=2.845 $Y=1.35 $X2=0 $Y2=0
cc_190 B1 N_C1_c_274_n 0.00279141f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_191 N_B1_c_241_n N_C1_c_274_n 0.0211059f $X=2.845 $Y=1.35 $X2=0 $Y2=0
cc_192 N_B1_M1008_g N_VPWR_c_301_n 0.00585385f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_193 N_B1_M1008_g N_VPWR_c_294_n 0.0110154f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_194 N_B1_c_242_n N_VGND_c_390_n 0.0120449f $X=2.845 $Y=1.185 $X2=0 $Y2=0
cc_195 N_B1_c_242_n N_VGND_c_391_n 0.00486043f $X=2.845 $Y=1.185 $X2=0 $Y2=0
cc_196 N_B1_c_242_n N_VGND_c_393_n 0.00515226f $X=2.845 $Y=1.185 $X2=0 $Y2=0
cc_197 N_C1_M1006_g N_VPWR_c_301_n 0.0054895f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_198 N_C1_M1006_g N_VPWR_c_294_n 0.011014f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_199 N_C1_c_271_n N_VGND_c_390_n 0.0118451f $X=3.295 $Y=1.185 $X2=0 $Y2=0
cc_200 N_C1_c_271_n N_VGND_c_392_n 0.00486043f $X=3.295 $Y=1.185 $X2=0 $Y2=0
cc_201 N_C1_c_271_n N_VGND_c_393_n 0.00556469f $X=3.295 $Y=1.185 $X2=0 $Y2=0
cc_202 N_VPWR_c_294_n N_X_M1003_s 0.00258346f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_296_n N_X_c_344_n 0.001542f $X=0.26 $Y=1.98 $X2=0 $Y2=0
cc_204 N_VPWR_c_299_n N_X_c_344_n 0.015291f $X=1 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_c_294_n N_X_c_344_n 0.0104192f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_294_n N_A_303_367#_M1009_s 0.00215158f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_207 N_VPWR_c_294_n N_A_303_367#_M1000_d 0.00298853f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_297_n N_A_303_367#_c_361_n 0.014565f $X=1.12 $Y=2.21 $X2=0 $Y2=0
cc_209 N_VPWR_c_297_n N_A_303_367#_c_362_n 0.0644662f $X=1.12 $Y=2.21 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_300_n N_A_303_367#_c_362_n 0.0200241f $X=1.96 $Y=3.33 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_294_n N_A_303_367#_c_362_n 0.0120544f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_M1009_d N_A_303_367#_c_366_n 0.00604565f $X=1.93 $Y=1.835 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_298_n N_A_303_367#_c_366_n 0.0225417f $X=2.125 $Y=2.505 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_301_n N_A_303_367#_c_371_n 0.0182658f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_215 N_VPWR_c_294_n N_A_303_367#_c_371_n 0.0125771f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_294_n A_590_367# 0.0115639f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_217 N_X_c_344_n N_VGND_c_389_n 0.001542f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_218 N_X_M1002_d N_VGND_c_393_n 0.00258346f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_219 N_X_c_344_n N_VGND_c_393_n 0.0104192f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_220 N_X_c_344_n N_VGND_c_394_n 0.015291f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_221 N_VGND_c_393_n A_386_47# 0.00312872f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
