* File: sky130_fd_sc_lp__iso1p_lp2.pex.spice
* Created: Wed Sep  2 09:58:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISO1P_LP2%A 3 7 9 12 14 15 17 24 25
c39 3 0 6.71001e-20 $X=0.66 $Y=0.495
r40 24 26 76.4623 $w=5.4e-07 $l=5.05e-07 $layer=POLY_cond $X=0.855 $Y=1.17
+ $X2=0.855 $Y2=1.675
r41 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.75
+ $Y=1.17 $X2=0.75 $Y2=1.17
r42 17 25 0.462998 $w=7.73e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.392
+ $X2=0.75 $Y2=1.392
r43 15 17 7.40797 $w=7.73e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.392
+ $X2=0.72 $Y2=1.392
r44 14 26 95.9558 $w=1.75e-07 $l=2.4e-07 $layer=POLY_cond $X=1.037 $Y=1.915
+ $X2=1.037 $Y2=1.675
r45 10 24 31.5348 $w=2.7e-07 $l=2.64953e-07 $layer=POLY_cond $X=1.05 $Y=1.005
+ $X2=0.855 $Y2=1.17
r46 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.05 $Y=1.005
+ $X2=1.05 $Y2=0.495
r47 7 14 36.7171 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.075 $Y=2.04
+ $X2=1.075 $Y2=1.915
r48 7 9 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.075 $Y=2.04
+ $X2=1.075 $Y2=2.545
r49 1 24 31.5348 $w=2.7e-07 $l=2.64953e-07 $layer=POLY_cond $X=0.66 $Y=1.005
+ $X2=0.855 $Y2=1.17
r50 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.66 $Y=1.005 $X2=0.66
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1P_LP2%SLEEP 3 6 9 11 13 15 16 17
c50 6 0 1.93391e-19 $X=1.575 $Y=1.665
r51 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.575
+ $Y=1.325 $X2=1.575 $Y2=1.325
r52 17 24 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=1.325
r53 16 24 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.63 $Y=1.295 $X2=1.63
+ $Y2=1.325
r54 11 23 85.7248 $w=2.05e-07 $l=2.65e-07 $layer=POLY_cond $X=1.84 $Y=1.262
+ $X2=1.575 $Y2=1.262
r55 11 13 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=1.84 $Y2=0.495
r56 9 15 177.644 $w=2.5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.535 $Y=2.545
+ $X2=1.535 $Y2=1.83
r57 6 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.665
+ $X2=1.575 $Y2=1.83
r58 6 23 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=1.575 $Y=1.665
+ $X2=1.575 $Y2=1.365
r59 1 23 30.7315 $w=2.05e-07 $l=9.5e-08 $layer=POLY_cond $X=1.48 $Y=1.262
+ $X2=1.575 $Y2=1.262
r60 1 3 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.48 $Y=1.16 $X2=1.48
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1P_LP2%A_137_409# 1 2 9 13 17 23 26 29 33 36 37
+ 41 42 47 49
c84 41 0 1.93391e-19 $X=2.36 $Y=1.03
c85 36 0 6.71001e-20 $X=1.185 $Y=2.025
r86 45 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.81 $Y=2.11
+ $X2=1.185 $Y2=2.11
r87 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.36
+ $Y=1.03 $X2=2.36 $Y2=1.03
r88 39 41 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.36 $Y=0.99 $X2=2.36
+ $Y2=1.03
r89 38 49 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.43 $Y=0.905
+ $X2=1.265 $Y2=0.905
r90 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.195 $Y=0.905
+ $X2=2.36 $Y2=0.99
r91 37 38 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.195 $Y=0.905
+ $X2=1.43 $Y2=0.905
r92 36 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.025
+ $X2=1.185 $Y2=2.11
r93 35 49 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.185 $Y=0.99
+ $X2=1.265 $Y2=0.905
r94 35 36 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=1.185 $Y=0.99
+ $X2=1.185 $Y2=2.025
r95 31 49 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=0.82
+ $X2=1.265 $Y2=0.905
r96 31 33 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.265 $Y=0.82
+ $X2=1.265 $Y2=0.495
r97 29 45 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.81 $Y=2.9
+ $X2=0.81 $Y2=2.195
r98 25 42 58.221 $w=3.35e-07 $l=3.38e-07 $layer=POLY_cond $X=2.362 $Y=1.368
+ $X2=2.362 $Y2=1.03
r99 25 26 32.6064 $w=3.35e-07 $l=1.67e-07 $layer=POLY_cond $X=2.362 $Y=1.368
+ $X2=2.362 $Y2=1.535
r100 22 42 2.58377 $w=3.35e-07 $l=1.5e-08 $layer=POLY_cond $X=2.362 $Y=1.015
+ $X2=2.362 $Y2=1.03
r101 22 23 152.804 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=2.362 $Y=0.94
+ $X2=2.66 $Y2=0.94
r102 19 22 47.1745 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=2.27 $Y=0.94
+ $X2=2.362 $Y2=0.94
r103 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.66 $Y=0.865
+ $X2=2.66 $Y2=0.94
r104 15 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.66 $Y=0.865
+ $X2=2.66 $Y2=0.495
r105 13 26 250.938 $w=2.5e-07 $l=1.01e-06 $layer=POLY_cond $X=2.405 $Y=2.545
+ $X2=2.405 $Y2=1.535
r106 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=0.865
+ $X2=2.27 $Y2=0.94
r107 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.27 $Y=0.865
+ $X2=2.27 $Y2=0.495
r108 2 45 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.81 $Y2=2.19
r109 2 29 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.81 $Y2=2.9
r110 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.285 $X2=1.265 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1P_LP2%KAPWR 1 4 6 12 16
r31 15 18 2.13585 $w=6.98e-07 $l=1.25e-07 $layer=LI1_cond $X=1.985 $Y=2.775
+ $X2=1.985 $Y2=2.9
r32 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.2 $Y=2.775
+ $X2=2.2 $Y2=2.775
r33 12 15 9.9958 $w=6.98e-07 $l=5.85e-07 $layer=LI1_cond $X=1.985 $Y=2.19
+ $X2=1.985 $Y2=2.775
r34 8 9 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.48 $Y=2.775
+ $X2=1.48 $Y2=2.775
r35 6 15 7.37187 $w=2.3e-07 $l=3.5e-07 $layer=LI1_cond $X=1.635 $Y=2.775
+ $X2=1.985 $Y2=2.775
r36 6 8 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.635 $Y=2.775
+ $X2=1.48 $Y2=2.775
r37 4 16 0.333634 $w=2.3e-07 $l=5.2e-07 $layer=MET1_cond $X=1.68 $Y=2.775
+ $X2=2.2 $Y2=2.775
r38 4 9 0.128321 $w=2.3e-07 $l=2e-07 $layer=MET1_cond $X=1.68 $Y=2.775 $X2=1.48
+ $Y2=2.775
r39 1 18 200 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=3 $X=1.66
+ $Y=2.045 $X2=1.8 $Y2=2.9
r40 1 12 200 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=3 $X=1.66
+ $Y=2.045 $X2=1.8 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1P_LP2%X 1 2 9 11 12 13 14 15 16 29
r21 16 40 5.80952 $w=5.23e-07 $l=2.55e-07 $layer=LI1_cond $X=2.972 $Y=1.665
+ $X2=2.972 $Y2=1.92
r22 15 16 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.972 $Y=1.295
+ $X2=2.972 $Y2=1.665
r23 14 15 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.972 $Y=0.925
+ $X2=2.972 $Y2=1.295
r24 13 14 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.972 $Y=0.555
+ $X2=2.972 $Y2=0.925
r25 13 29 1.36695 $w=5.23e-07 $l=6e-08 $layer=LI1_cond $X=2.972 $Y=0.555
+ $X2=2.972 $Y2=0.495
r26 12 48 5.51829 $w=7.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.87 $Y=2.405
+ $X2=2.87 $Y2=2.52
r27 12 44 3.5227 $w=7.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.87 $Y=2.405
+ $X2=2.87 $Y2=2.19
r28 11 44 2.53962 $w=7.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.87 $Y=2.035
+ $X2=2.87 $Y2=2.19
r29 11 40 2.84659 $w=7.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.87 $Y=2.035
+ $X2=2.87 $Y2=1.92
r30 9 48 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.67 $Y=2.9 $X2=2.67
+ $Y2=2.52
r31 2 44 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=2.045 $X2=2.67 $Y2=2.19
r32 2 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=2.045 $X2=2.67 $Y2=2.9
r33 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.285 $X2=2.875 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1P_LP2%VGND 1 2 9 13 16 17 18 23 32 33 36
r36 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r37 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r38 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 30 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.055
+ $Y2=0
r40 30 32 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=3.12
+ $Y2=0
r41 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r42 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.055
+ $Y2=0
r44 23 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r45 22 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 18 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r48 18 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r49 18 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 16 21 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=0.28 $Y=0 $X2=0.24
+ $Y2=0
r51 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0 $X2=0.445
+ $Y2=0
r52 15 25 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.72
+ $Y2=0
r53 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.445
+ $Y2=0
r54 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r55 11 13 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.475
r56 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=0.085
+ $X2=0.445 $Y2=0
r57 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.445 $Y=0.085
+ $X2=0.445 $Y2=0.495
r58 2 13 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.285 $X2=2.055 $Y2=0.475
r59 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.3
+ $Y=0.285 $X2=0.445 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__ISO1P_LP2%VPWR 1 8 14
r19 5 14 0.00453869 $w=3.36e-06 $l=1.22e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.208
r20 5 8 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r21 4 8 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=3.12
+ $Y2=3.33
r22 4 5 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 1 14 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=3.207
+ $X2=1.68 $Y2=3.208
.ends

