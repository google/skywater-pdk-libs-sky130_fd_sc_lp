* File: sky130_fd_sc_lp__xor3_lp.spice
* Created: Wed Sep  2 10:41:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor3_lp.pex.spice"
.subckt sky130_fd_sc_lp__xor3_lp  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_144_113# N_A_M1002_g N_A_57_113#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_M1025_g A_144_113# VNB NSHORT L=0.15 W=0.42 AD=0.1932
+ AS=0.0441 PD=1.34 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75003.1
+ A=0.063 P=1.14 MULT=1
MM1000 A_430_113# N_A_57_113#_M1000_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1932 PD=0.66 PS=1.34 NRD=18.564 NRS=182.856 M=1 R=2.8
+ SA=75001.6 SB=75002 A=0.063 P=1.14 MULT=1
MM1013 N_A_388_419#_M1013_d N_A_57_113#_M1013_g A_430_113# VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_494_419#_M1009_d N_A_580_21#_M1009_g N_A_388_419#_M1013_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.12735 AS=0.0756 PD=1.045 PS=0.78 NRD=22.848 NRS=22.848 M=1
+ R=2.8 SA=75002.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_57_113#_M1006_d N_B_M1006_g N_A_494_419#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.101412 AS=0.12735 PD=1.075 PS=1.045 NRD=53.268 NRS=58.56 M=1 R=2.8
+ SA=75002.8 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1018 N_A_855_66#_M1018_d N_A_580_21#_M1018_g N_A_57_113#_M1006_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.130825 AS=0.101412 PD=1.125 PS=1.075 NRD=22.848 NRS=0 M=1
+ R=2.8 SA=75001.3 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1016 N_A_388_419#_M1016_d N_B_M1016_g N_A_855_66#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.130825 PD=1.41 PS=1.125 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_1245_89# N_B_M1015_g N_A_580_21#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_B_M1010_g A_1245_89# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_1459_406#_M1005_d N_C_M1005_g N_A_494_419#_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0651 AS=0.1407 PD=0.73 PS=1.51 NRD=8.568 NRS=14.28 M=1 R=2.8
+ SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_A_855_66#_M1022_d N_A_1393_300#_M1022_g N_A_1459_406#_M1005_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.1533 AS=0.0651 PD=1.57 PS=0.73 NRD=22.848 NRS=0 M=1
+ R=2.8 SA=75000.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1008 A_1860_141# N_C_M1008_g N_A_1393_300#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1659 PD=0.63 PS=1.63 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75000.3
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g A_1860_141# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0441 PD=0.84 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1011 A_2046_141# N_A_1459_406#_M1011_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_1459_406#_M1004_g A_2046_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_M1023_g N_A_57_113#_M1023_s VPB PHIGHVT L=0.25 W=1
+ AD=0.405 AS=0.285 PD=1.81 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_388_419#_M1003_d N_A_57_113#_M1003_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.405 PD=1.28 PS=1.81 NRD=0 NRS=104.39 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1017 N_A_494_419#_M1017_d N_B_M1017_g N_A_388_419#_M1003_d VPB PHIGHVT L=0.25
+ W=1 AD=0.4075 AS=0.14 PD=1.815 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1019 N_A_57_113#_M1019_d N_A_580_21#_M1019_g N_A_494_419#_M1017_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.31 AS=0.4075 PD=1.62 PS=1.815 NRD=0 NRS=105.375 M=1 R=4
+ SA=125003 SB=125002 A=0.25 P=2.5 MULT=1
MM1020 N_A_855_66#_M1020_d N_B_M1020_g N_A_57_113#_M1019_d VPB PHIGHVT L=0.25
+ W=1 AD=0.145 AS=0.31 PD=1.29 PS=1.62 NRD=1.9503 NRS=66.98 M=1 R=4 SA=125004
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1007 N_A_388_419#_M1007_d N_A_580_21#_M1007_g N_A_855_66#_M1020_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.145 PD=2.57 PS=1.29 NRD=0 NRS=0 M=1 R=4 SA=125004
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1014 N_VPWR_M1014_d N_B_M1014_g N_A_580_21#_M1014_s VPB PHIGHVT L=0.25 W=1
+ AD=0.365 AS=0.375 PD=2.73 PS=2.75 NRD=15.7403 NRS=17.73 M=1 R=4 SA=125000
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1024 N_A_1459_406#_M1024_d N_A_1393_300#_M1024_g N_A_494_419#_M1024_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4
+ SA=125000 SB=125001 A=0.25 P=2.5 MULT=1
MM1012 N_A_855_66#_M1012_d N_C_M1012_g N_A_1459_406#_M1024_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1026 N_VPWR_M1026_d N_C_M1026_g N_A_1393_300#_M1026_s VPB PHIGHVT L=0.25 W=1
+ AD=0.305 AS=0.285 PD=1.61 PS=2.57 NRD=65.01 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1021 N_X_M1021_d N_A_1459_406#_M1021_g N_VPWR_M1026_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.305 PD=2.57 PS=1.61 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX27_noxref VNB VPB NWDIODE A=21.2983 P=26.57
c_116 VNB 0 1.81544e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__xor3_lp.pxi.spice"
*
.ends
*
*
