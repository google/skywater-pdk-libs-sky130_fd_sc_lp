* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ha_lp A B VGND VNB VPB VPWR COUT SUM
X0 a_296_286# B a_743_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_296_286# a_83_153# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VPWR B a_296_286# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_743_125# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_901_125# a_296_286# COUT VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_83_153# B a_493_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 SUM a_83_153# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 VGND a_296_286# a_901_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_296_286# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_113_179# a_83_153# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_83_153# a_296_286# a_369_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_493_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_369_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 SUM a_83_153# a_113_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND A a_369_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_296_286# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
