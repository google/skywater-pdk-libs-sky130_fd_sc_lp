* NGSPICE file created from sky130_fd_sc_lp__a2111oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_253_367# C1 a_157_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.78e+11p pd=3.12e+06u as=4.158e+11p ps=3.18e+06u
M1001 VPWR A1 a_343_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=5.292e+11p pd=3.36e+06u as=8.631e+11p ps=6.41e+06u
M1002 Y D1 VGND VNB nshort w=840000u l=150000u
+  ad=6.846e+11p pd=4.99e+06u as=1.0122e+12p ps=7.45e+06u
M1003 VGND A2 a_499_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1004 a_343_367# B1 a_253_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_157_367# D1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=6.048e+11p ps=3.48e+06u
M1006 a_499_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_343_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

