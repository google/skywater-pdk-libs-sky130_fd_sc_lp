* File: sky130_fd_sc_lp__ha_lp.spice
* Created: Wed Sep  2 09:54:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ha_lp.pex.spice"
.subckt sky130_fd_sc_lp__ha_lp  VNB VPB B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1008 A_113_179# N_A_83_153#_M1008_g N_SUM_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_83_153#_M1006_g A_113_179# VNB NSHORT L=0.15 W=0.42
+ AD=0.11865 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_369_47#_M1005_d N_A_296_286#_M1005_g N_A_83_153#_M1005_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.11865 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_A_369_47#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1015 N_A_369_47#_M1015_d N_A_M1015_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0588 PD=1.4 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 A_743_125# N_B_M1003_g N_A_296_286#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g A_743_125# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1002 A_901_125# N_A_296_286#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_COUT_M1014_d N_A_296_286#_M1014_g A_901_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_83_153#_M1004_g N_SUM_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1013 N_A_83_153#_M1013_d N_A_296_286#_M1013_g N_VPWR_M1004_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.2425 AS=0.14 PD=1.485 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1010 A_493_419# N_B_M1010_g N_A_83_153#_M1013_d VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.2425 PD=1.32 PS=1.485 NRD=20.6653 NRS=40.3653 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_493_419# VPB PHIGHVT L=0.25 W=1 AD=0.165
+ AS=0.16 PD=1.33 PS=1.32 NRD=0 NRS=20.6653 M=1 R=4 SA=125002 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1000 N_A_296_286#_M1000_d N_B_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.165 PD=1.28 PS=1.33 NRD=0 NRS=9.8303 M=1 R=4 SA=125003 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_A_296_286#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1875 AS=0.14 PD=1.375 PS=1.28 NRD=18.715 NRS=0 M=1 R=4 SA=125003
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1012 N_COUT_M1012_d N_A_296_286#_M1012_g N_VPWR_M1011_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1875 PD=2.57 PS=1.375 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125000
+ A=0.25 P=2.5 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5559 P=15.05
c_109 VPB 0 1.51007e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__ha_lp.pxi.spice"
*
.ends
*
*
