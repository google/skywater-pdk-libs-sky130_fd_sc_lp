* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_0 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 SUM a_1059_119# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=8.56e+11p ps=8.58e+06u
M1001 VGND A a_1239_119# VNB nshort w=420000u l=150000u
+  ad=7.1035e+11p pd=7.7e+06u as=1.989e+11p ps=2.16e+06u
M1002 a_781_119# CIN VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1003 a_224_119# A VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_781_457# CIN VPWR VPB phighvt w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1005 a_404_532# CIN a_80_225# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.638e+11p ps=1.62e+06u
M1006 SUM a_1059_119# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 VPWR a_80_225# COUT VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1008 a_781_457# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1239_457# B a_1161_457# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.008e+11p ps=1.32e+06u
M1010 a_218_532# A VPWR VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1011 a_1059_119# a_80_225# a_781_119# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1012 a_1145_119# CIN a_1059_119# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1013 a_781_119# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1239_119# B a_1145_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_1239_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_404_532# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B a_781_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B a_781_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1161_457# CIN a_1059_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.512e+11p ps=1.56e+06u
M1020 a_80_225# B a_224_119# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1021 VPWR B a_404_532# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_382_119# CIN a_80_225# VNB nshort w=420000u l=150000u
+  ad=2.457e+11p pd=2.85e+06u as=0p ps=0u
M1023 a_382_119# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1059_119# a_80_225# a_781_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_80_225# B a_218_532# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_80_225# COUT VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1027 VGND B a_382_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
