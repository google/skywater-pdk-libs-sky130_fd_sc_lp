* File: sky130_fd_sc_lp__dlxbp_lp.pex.spice
* Created: Fri Aug 28 10:28:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%D 1 3 7 11 15 22 23 24 25 30
c41 1 0 1.08557e-19 $X=0.485 $Y=1.85
r42 24 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.735 $Y=1.665
+ $X2=0.735 $Y2=2.035
r43 23 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.735 $Y=1.295
+ $X2=0.735 $Y2=1.665
r44 23 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.735
+ $Y=1.345 $X2=0.735 $Y2=1.345
r45 22 30 6.42035 $w=5e-07 $l=6e-08 $layer=POLY_cond $X=0.67 $Y=1.285 $X2=0.67
+ $Y2=1.345
r46 18 30 37.9871 $w=5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.67 $Y=1.7 $X2=0.67
+ $Y2=1.345
r47 5 22 24.5449 $w=5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=1.135
+ $X2=0.675 $Y2=1.285
r48 5 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.855 $Y=1.135
+ $X2=0.855 $Y2=0.765
r49 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.495 $Y=1.135
+ $X2=0.495 $Y2=0.765
r50 1 18 24.5449 $w=5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.665 $Y=1.85 $X2=0.665
+ $Y2=1.7
r51 1 11 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.845 $Y=1.85
+ $X2=0.845 $Y2=2.725
r52 1 3 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.485 $Y=1.85
+ $X2=0.485 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%GATE 3 7 11 15 17 18 22
c56 22 0 1.56912e-19 $X=1.295 $Y=1.69
c57 3 0 9.31616e-20 $X=1.285 $Y=0.765
r58 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.295
+ $Y=1.69 $X2=1.295 $Y2=1.69
r59 18 23 13.0358 $w=3.03e-07 $l=3.45e-07 $layer=LI1_cond $X=1.237 $Y=2.035
+ $X2=1.237 $Y2=1.69
r60 17 23 0.944625 $w=3.03e-07 $l=2.5e-08 $layer=LI1_cond $X=1.237 $Y=1.665
+ $X2=1.237 $Y2=1.69
r61 13 22 81.4778 $w=3.1e-07 $l=6.1131e-07 $layer=POLY_cond $X=1.675 $Y=2.195
+ $X2=1.44 $Y2=1.69
r62 13 15 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.675 $Y=2.195
+ $X2=1.675 $Y2=2.725
r63 9 22 28.6132 $w=3.1e-07 $l=3.06594e-07 $layer=POLY_cond $X=1.675 $Y=1.525
+ $X2=1.44 $Y2=1.69
r64 9 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.675 $Y=1.525
+ $X2=1.675 $Y2=0.765
r65 5 22 81.4778 $w=3.1e-07 $l=5.64048e-07 $layer=POLY_cond $X=1.315 $Y=2.195
+ $X2=1.44 $Y2=1.69
r66 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.315 $Y=2.195
+ $X2=1.315 $Y2=2.725
r67 1 22 28.6132 $w=3.1e-07 $l=1.55e-07 $layer=POLY_cond $X=1.285 $Y=1.69
+ $X2=1.44 $Y2=1.69
r68 1 3 389.702 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.285 $Y=1.69
+ $X2=1.285 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%A_350_111# 1 2 9 15 19 23 27 31 33 34 36 37
+ 39 43 44 47 49 55 56 65 68 69
c153 69 0 8.94403e-20 $X=4.515 $Y=0.99
c154 44 0 1.16136e-19 $X=4.11 $Y=2
c155 43 0 3.07343e-20 $X=4.11 $Y=2
c156 23 0 1.41808e-19 $X=3.12 $Y=2.695
r157 69 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.515 $Y=0.99
+ $X2=4.515 $Y2=0.825
r158 68 71 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.515 $Y=0.99
+ $X2=4.515 $Y2=1.155
r159 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.515
+ $Y=0.99 $X2=4.515 $Y2=0.99
r160 60 62 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.795 $Y=1.68
+ $X2=2.795 $Y2=1.685
r161 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.68 $X2=2.795 $Y2=1.68
r162 58 60 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.795 $Y=1.42
+ $X2=2.795 $Y2=1.68
r163 56 61 32.1965 $w=5.65e-07 $l=3.4e-07 $layer=POLY_cond $X=2.912 $Y=1.34
+ $X2=2.912 $Y2=1.68
r164 55 58 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.795 $Y=1.34
+ $X2=2.795 $Y2=1.42
r165 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.34 $X2=2.795 $Y2=1.34
r166 49 51 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=1.907 $Y=0.765
+ $X2=1.907 $Y2=0.995
r167 47 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=1.335
+ $X2=4.435 $Y2=1.42
r168 47 71 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.435 $Y=1.335
+ $X2=4.435 $Y2=1.155
r169 44 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.11 $Y=2 $X2=4.11
+ $Y2=2.165
r170 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.11 $Y=2
+ $X2=4.11 $Y2=2
r171 41 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.11 $Y=1.42
+ $X2=4.435 $Y2=1.42
r172 41 43 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.11 $Y=1.505
+ $X2=4.11 $Y2=2
r173 40 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=1.42
+ $X2=2.795 $Y2=1.42
r174 39 41 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=1.42
+ $X2=4.11 $Y2=1.42
r175 39 40 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=3.945 $Y=1.42
+ $X2=2.96 $Y2=1.42
r176 38 53 2.98112 $w=3.2e-07 $l=1.27475e-07 $layer=LI1_cond $X=2.17 $Y=1.685
+ $X2=2.045 $Y2=1.69
r177 37 62 0.903439 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=1.685
+ $X2=2.795 $Y2=1.685
r178 37 38 16.5664 $w=3.18e-07 $l=4.6e-07 $layer=LI1_cond $X=2.63 $Y=1.685
+ $X2=2.17 $Y2=1.685
r179 36 53 4.70099 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=2.005 $Y=1.525
+ $X2=2.045 $Y2=1.69
r180 36 51 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.005 $Y=1.525
+ $X2=2.005 $Y2=0.995
r181 33 34 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=2.732 $Y=2.085
+ $X2=2.732 $Y2=2.235
r182 31 78 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.425 $Y=0.445
+ $X2=4.425 $Y2=0.825
r183 27 76 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.02 $Y=2.695
+ $X2=4.02 $Y2=2.165
r184 21 61 30.5737 $w=2.82e-07 $l=2.78539e-07 $layer=POLY_cond $X=3.12 $Y=1.845
+ $X2=2.912 $Y2=1.68
r185 21 23 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=3.12 $Y=1.845
+ $X2=3.12 $Y2=2.695
r186 17 56 30.5737 $w=2.82e-07 $l=2.52357e-07 $layer=POLY_cond $X=3.095 $Y=1.175
+ $X2=2.912 $Y2=1.34
r187 17 19 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.095 $Y=1.175
+ $X2=3.095 $Y2=0.445
r188 15 34 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.76 $Y=2.695
+ $X2=2.76 $Y2=2.235
r189 11 61 30.5737 $w=2.82e-07 $l=2.77496e-07 $layer=POLY_cond $X=2.705 $Y=1.845
+ $X2=2.912 $Y2=1.68
r190 11 33 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.705 $Y=1.845
+ $X2=2.705 $Y2=2.085
r191 7 56 30.5737 $w=2.82e-07 $l=2.77496e-07 $layer=POLY_cond $X=2.705 $Y=1.175
+ $X2=2.912 $Y2=1.34
r192 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.705 $Y=1.175
+ $X2=2.705 $Y2=0.445
r193 2 53 600 $w=1.7e-07 $l=8.32797e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.405 $X2=2.005 $Y2=1.69
r194 1 49 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.555 $X2=1.89 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%A_27_111# 1 2 11 15 18 20 23 27 28 30 31 32
+ 34 38 40 41 46
c106 23 0 1.08557e-19 $X=1.405 $Y=2.47
c107 18 0 1.47075e-19 $X=3.51 $Y=1.595
r108 41 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=2.03
+ $X2=3.57 $Y2=2.195
r109 41 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=2.03
+ $X2=3.57 $Y2=1.865
r110 40 43 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.57 $Y=2.03 $X2=3.57
+ $Y2=2.11
r111 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=2.03 $X2=3.57 $Y2=2.03
r112 34 36 10.6751 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=0.275 $Y=0.765
+ $X2=0.275 $Y2=0.995
r113 31 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=2.11
+ $X2=3.57 $Y2=2.11
r114 31 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.405 $Y=2.11
+ $X2=3.07 $Y2=2.11
r115 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.985 $Y=2.195
+ $X2=3.07 $Y2=2.11
r116 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.985 $Y=2.195
+ $X2=2.985 $Y2=2.895
r117 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.9 $Y=2.98
+ $X2=2.985 $Y2=2.895
r118 27 28 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=2.9 $Y=2.98
+ $X2=1.575 $Y2=2.98
r119 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.49 $Y=2.895
+ $X2=1.575 $Y2=2.98
r120 25 26 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.49 $Y=2.555
+ $X2=1.49 $Y2=2.895
r121 24 38 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.47
+ $X2=0.27 $Y2=2.47
r122 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=2.47
+ $X2=1.49 $Y2=2.555
r123 23 24 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.405 $Y=2.47
+ $X2=0.435 $Y2=2.47
r124 20 38 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.19 $Y=2.385
+ $X2=0.27 $Y2=2.47
r125 20 36 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=0.19 $Y=2.385
+ $X2=0.19 $Y2=0.995
r126 18 46 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.495 $Y=1.595
+ $X2=3.495 $Y2=1.865
r127 17 18 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.51 $Y=1.445
+ $X2=3.51 $Y2=1.595
r128 15 47 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.63 $Y=2.695
+ $X2=3.63 $Y2=2.195
r129 11 17 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.525 $Y=0.445
+ $X2=3.525 $Y2=1.445
r130 2 38 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.27 $Y2=2.55
r131 1 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.555 $X2=0.28 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%A_469_47# 1 2 9 11 12 15 19 21 22 23 25 26
+ 27 31 34 36 37 40 42 46
c133 46 0 2.58091e-20 $X=3.975 $Y=0.99
c134 36 0 1.47075e-19 $X=3.81 $Y=0.91
c135 26 0 1.41808e-19 $X=2.38 $Y=2.12
c136 23 0 9.31616e-20 $X=1.545 $Y=0.35
c137 15 0 1.24e-19 $X=4.56 $Y=2.805
r138 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=0.99 $X2=3.975 $Y2=0.99
r139 42 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.975 $Y=0.91
+ $X2=3.975 $Y2=0.99
r140 38 40 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.46 $Y=1.26
+ $X2=1.655 $Y2=1.26
r141 36 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=0.91
+ $X2=3.975 $Y2=0.91
r142 36 37 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=3.81 $Y=0.91
+ $X2=2.655 $Y2=0.91
r143 32 34 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.545 $Y=2.205
+ $X2=2.545 $Y2=2.535
r144 29 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.49 $Y=0.825
+ $X2=2.655 $Y2=0.91
r145 29 31 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.49 $Y=0.825
+ $X2=2.49 $Y2=0.47
r146 28 31 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.49 $Y=0.435
+ $X2=2.49 $Y2=0.47
r147 26 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.38 $Y=2.12
+ $X2=2.545 $Y2=2.205
r148 26 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.38 $Y=2.12
+ $X2=1.74 $Y2=2.12
r149 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.655 $Y=2.035
+ $X2=1.74 $Y2=2.12
r150 24 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=1.345
+ $X2=1.655 $Y2=1.26
r151 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.655 $Y=1.345
+ $X2=1.655 $Y2=2.035
r152 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.325 $Y=0.35
+ $X2=2.49 $Y2=0.435
r153 22 23 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.325 $Y=0.35
+ $X2=1.545 $Y2=0.35
r154 21 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=1.175
+ $X2=1.46 $Y2=1.26
r155 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.46 $Y=0.435
+ $X2=1.545 $Y2=0.35
r156 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.46 $Y=0.435
+ $X2=1.46 $Y2=1.175
r157 19 46 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=3.975 $Y=1.395
+ $X2=3.975 $Y2=0.99
r158 18 46 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=0.825
+ $X2=3.975 $Y2=0.99
r159 13 15 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=4.56 $Y=1.545
+ $X2=4.56 $Y2=2.805
r160 12 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.14 $Y=1.47
+ $X2=3.975 $Y2=1.395
r161 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.485 $Y=1.47
+ $X2=4.56 $Y2=1.545
r162 11 12 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.485 $Y=1.47
+ $X2=4.14 $Y2=1.47
r163 9 18 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=3.915 $Y=0.445
+ $X2=3.915 $Y2=0.825
r164 2 34 600 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=2.375 $X2=2.545 $Y2=2.535
r165 1 31 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.235 $X2=2.49 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%A_969_407# 1 2 9 13 17 21 25 29 33 37 39 40
+ 43 47 49 50 53 57 61 64 72 75 77 78 80
c155 40 0 3.39681e-19 $X=7.985 $Y=1.38
c156 13 0 3.07343e-20 $X=4.965 $Y=0.445
r157 90 91 9.55183 $w=3.28e-07 $l=6.5e-08 $layer=POLY_cond $X=7.845 $Y=1.44
+ $X2=7.91 $Y2=1.44
r158 87 88 11.0213 $w=3.28e-07 $l=7.5e-08 $layer=POLY_cond $X=7.3 $Y=1.44
+ $X2=7.375 $Y2=1.44
r159 86 87 41.8811 $w=3.28e-07 $l=2.85e-07 $layer=POLY_cond $X=7.015 $Y=1.44
+ $X2=7.3 $Y2=1.44
r160 85 86 11.0213 $w=3.28e-07 $l=7.5e-08 $layer=POLY_cond $X=6.94 $Y=1.44
+ $X2=7.015 $Y2=1.44
r161 77 79 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.26 $Y=1.95
+ $X2=6.26 $Y2=2.2
r162 77 78 6.24272 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.26 $Y=1.95
+ $X2=6.26 $Y2=1.785
r163 73 90 56.5762 $w=3.28e-07 $l=3.85e-07 $layer=POLY_cond $X=7.46 $Y=1.44
+ $X2=7.845 $Y2=1.44
r164 73 88 12.4909 $w=3.28e-07 $l=8.5e-08 $layer=POLY_cond $X=7.46 $Y=1.44
+ $X2=7.375 $Y2=1.44
r165 72 73 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.46
+ $Y=1.44 $X2=7.46 $Y2=1.44
r166 70 85 23.5122 $w=3.28e-07 $l=1.6e-07 $layer=POLY_cond $X=6.78 $Y=1.44
+ $X2=6.94 $Y2=1.44
r167 69 72 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.78 $Y=1.44
+ $X2=7.46 $Y2=1.44
r168 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.78
+ $Y=1.44 $X2=6.78 $Y2=1.44
r169 67 80 0.105856 $w=3.3e-07 $l=1.33e-07 $layer=LI1_cond $X=6.425 $Y=1.44
+ $X2=6.292 $Y2=1.44
r170 67 69 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.425 $Y=1.44
+ $X2=6.78 $Y2=1.44
r171 65 80 7.19657 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=6.292 $Y=1.605
+ $X2=6.292 $Y2=1.44
r172 65 78 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=6.292 $Y=1.605
+ $X2=6.292 $Y2=1.785
r173 64 80 7.19657 $w=2.17e-07 $l=1.87029e-07 $layer=LI1_cond $X=6.245 $Y=1.275
+ $X2=6.292 $Y2=1.44
r174 64 75 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.245 $Y=1.275
+ $X2=6.245 $Y2=1.095
r175 59 79 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.26 $Y=2.365
+ $X2=6.26 $Y2=2.2
r176 59 61 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=6.26 $Y=2.365
+ $X2=6.26 $Y2=2.9
r177 55 75 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=0.93
+ $X2=6.165 $Y2=1.095
r178 55 57 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.165 $Y=0.93
+ $X2=6.165 $Y2=0.43
r179 53 83 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.01 $Y=2.2
+ $X2=5.01 $Y2=2.365
r180 53 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.01 $Y=2.2
+ $X2=5.01 $Y2=2.035
r181 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=2.2 $X2=5.01 $Y2=2.2
r182 50 79 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=2.2
+ $X2=6.26 $Y2=2.2
r183 50 52 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=6.095 $Y=2.2
+ $X2=5.01 $Y2=2.2
r184 45 49 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=8.27 $Y=1.455
+ $X2=8.252 $Y2=1.38
r185 45 47 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.27 $Y=1.455
+ $X2=8.27 $Y2=2.125
r186 41 49 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=8.235 $Y=1.305
+ $X2=8.252 $Y2=1.38
r187 41 43 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.235 $Y=1.305
+ $X2=8.235 $Y2=0.865
r188 40 91 25.362 $w=3.28e-07 $l=1.00623e-07 $layer=POLY_cond $X=7.985 $Y=1.38
+ $X2=7.91 $Y2=1.44
r189 39 49 5.30422 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=8.16 $Y=1.38
+ $X2=8.252 $Y2=1.38
r190 39 40 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=8.16 $Y=1.38
+ $X2=7.985 $Y2=1.38
r191 35 91 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.91 $Y=1.605
+ $X2=7.91 $Y2=1.44
r192 35 37 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.91 $Y=1.605
+ $X2=7.91 $Y2=2.125
r193 31 90 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.845 $Y=1.275
+ $X2=7.845 $Y2=1.44
r194 31 33 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.845 $Y=1.275
+ $X2=7.845 $Y2=0.865
r195 27 88 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.375 $Y=1.605
+ $X2=7.375 $Y2=1.44
r196 27 29 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.375 $Y=1.605
+ $X2=7.375 $Y2=2.435
r197 23 87 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.3 $Y=1.275
+ $X2=7.3 $Y2=1.44
r198 23 25 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.3 $Y=1.275
+ $X2=7.3 $Y2=0.655
r199 19 86 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.015 $Y=1.605
+ $X2=7.015 $Y2=1.44
r200 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.015 $Y=1.605
+ $X2=7.015 $Y2=2.435
r201 15 85 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.275
+ $X2=6.94 $Y2=1.44
r202 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.94 $Y=1.275
+ $X2=6.94 $Y2=0.655
r203 13 82 815.298 $w=1.5e-07 $l=1.59e-06 $layer=POLY_cond $X=4.965 $Y=0.445
+ $X2=4.965 $Y2=2.035
r204 9 83 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.95 $Y=2.805
+ $X2=4.95 $Y2=2.365
r205 2 77 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.12
+ $Y=1.805 $X2=6.26 $Y2=1.95
r206 2 61 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=6.12
+ $Y=1.805 $X2=6.26 $Y2=2.9
r207 1 57 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=6.025
+ $Y=0.235 $X2=6.165 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%A_798_47# 1 2 9 13 17 21 23 28 29 30 32 33
+ 35 39 47
c106 35 0 1.61717e-19 $X=5.805 $Y=1.44
c107 33 0 1.24e-19 $X=5.03 $Y=1.44
c108 30 0 2.05576e-19 $X=4.625 $Y=1.77
r109 47 48 17.8867 $w=2.56e-07 $l=9.5e-08 $layer=POLY_cond $X=5.95 $Y=1.44
+ $X2=6.045 $Y2=1.44
r110 36 47 27.3008 $w=2.56e-07 $l=1.45e-07 $layer=POLY_cond $X=5.805 $Y=1.44
+ $X2=5.95 $Y2=1.44
r111 36 45 22.5938 $w=2.56e-07 $l=1.2e-07 $layer=POLY_cond $X=5.805 $Y=1.44
+ $X2=5.685 $Y2=1.44
r112 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.805
+ $Y=1.44 $X2=5.805 $Y2=1.44
r113 33 42 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.945 $Y=1.44
+ $X2=4.945 $Y2=1.77
r114 33 35 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=5.03 $Y=1.44
+ $X2=5.805 $Y2=1.44
r115 32 33 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.945 $Y=1.275
+ $X2=4.945 $Y2=1.44
r116 31 32 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=4.945 $Y=0.645
+ $X2=4.945 $Y2=1.275
r117 29 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.86 $Y=1.77
+ $X2=4.945 $Y2=1.77
r118 29 30 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.86 $Y=1.77
+ $X2=4.625 $Y2=1.77
r119 28 39 10.8801 $w=3.42e-07 $l=4.03949e-07 $layer=LI1_cond $X=4.54 $Y=2.575
+ $X2=4.235 $Y2=2.805
r120 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.54 $Y=1.855
+ $X2=4.625 $Y2=1.77
r121 27 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.54 $Y=1.855
+ $X2=4.54 $Y2=2.575
r122 23 31 7.93686 $w=3.5e-07 $l=2.13307e-07 $layer=LI1_cond $X=4.86 $Y=0.47
+ $X2=4.945 $Y2=0.645
r123 23 25 21.4025 $w=3.48e-07 $l=6.5e-07 $layer=LI1_cond $X=4.86 $Y=0.47
+ $X2=4.21 $Y2=0.47
r124 19 48 15.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.605
+ $X2=6.045 $Y2=1.44
r125 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=6.045 $Y=1.605
+ $X2=6.045 $Y2=2.435
r126 15 47 15.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.275
+ $X2=5.95 $Y2=1.44
r127 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.95 $Y=1.275
+ $X2=5.95 $Y2=0.655
r128 11 45 15.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.685 $Y=1.605
+ $X2=5.685 $Y2=1.44
r129 11 13 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=5.685 $Y=1.605
+ $X2=5.685 $Y2=2.435
r130 7 45 17.8867 $w=2.56e-07 $l=2.07123e-07 $layer=POLY_cond $X=5.59 $Y=1.275
+ $X2=5.685 $Y2=1.44
r131 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.59 $Y=1.275
+ $X2=5.59 $Y2=0.655
r132 2 39 600 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=2.375 $X2=4.235 $Y2=2.805
r133 1 25 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.21 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%A_1662_131# 1 2 9 13 17 21 25 29 33 36 42
c52 36 0 2.24197e-19 $X=8.467 $Y=1.47
r53 41 42 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.585 $Y=1.47
+ $X2=9.6 $Y2=1.47
r54 37 39 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.225 $Y=1.47
+ $X2=9.24 $Y2=1.47
r55 34 41 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=9.29 $Y=1.47
+ $X2=9.585 $Y2=1.47
r56 34 39 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=9.29 $Y=1.47 $X2=9.24
+ $Y2=1.47
r57 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.29
+ $Y=1.47 $X2=9.29 $Y2=1.47
r58 31 36 1.52928 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=8.65 $Y=1.47
+ $X2=8.467 $Y2=1.47
r59 31 33 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=8.65 $Y=1.47
+ $X2=9.29 $Y2=1.47
r60 27 36 4.94753 $w=3.47e-07 $l=1.65e-07 $layer=LI1_cond $X=8.467 $Y=1.635
+ $X2=8.467 $Y2=1.47
r61 27 29 9.94574 $w=3.63e-07 $l=3.15e-07 $layer=LI1_cond $X=8.467 $Y=1.635
+ $X2=8.467 $Y2=1.95
r62 23 36 4.94753 $w=3.47e-07 $l=1.73292e-07 $layer=LI1_cond $X=8.45 $Y=1.305
+ $X2=8.467 $Y2=1.47
r63 23 25 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=8.45 $Y=1.305
+ $X2=8.45 $Y2=0.865
r64 19 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.6 $Y=1.635
+ $X2=9.6 $Y2=1.47
r65 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.6 $Y=1.635 $X2=9.6
+ $Y2=2.465
r66 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.585 $Y=1.305
+ $X2=9.585 $Y2=1.47
r67 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=9.585 $Y=1.305
+ $X2=9.585 $Y2=0.685
r68 11 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.24 $Y=1.635
+ $X2=9.24 $Y2=1.47
r69 11 13 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.24 $Y=1.635
+ $X2=9.24 $Y2=2.465
r70 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.225 $Y=1.305
+ $X2=9.225 $Y2=1.47
r71 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=9.225 $Y=1.305
+ $X2=9.225 $Y2=0.685
r72 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.345
+ $Y=1.805 $X2=8.485 $Y2=1.95
r73 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.31
+ $Y=0.655 $X2=8.45 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%VPWR 1 2 3 4 5 18 22 26 30 36 41 42 43 45
+ 54 61 66 73 74 77 80 83 86
r107 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r108 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r109 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 74 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r112 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r113 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.19 $Y=3.33
+ $X2=9.025 $Y2=3.33
r114 71 73 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.19 $Y=3.33
+ $X2=9.84 $Y2=3.33
r115 70 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r117 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 67 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.59 $Y2=3.33
r119 67 69 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 66 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=9.025 $Y2=3.33
r121 66 69 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 65 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r124 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r125 62 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.635 $Y=3.33
+ $X2=5.47 $Y2=3.33
r126 62 64 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.635 $Y=3.33
+ $X2=6 $Y2=3.33
r127 61 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.425 $Y=3.33
+ $X2=7.59 $Y2=3.33
r128 61 64 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=7.425 $Y=3.33
+ $X2=6 $Y2=3.33
r129 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r130 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r131 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.305 $Y=3.33
+ $X2=5.47 $Y2=3.33
r132 54 59 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.305 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 53 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 53 78 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 50 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.06 $Y2=3.33
r137 50 52 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=3.12 $Y2=3.33
r138 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.06 $Y2=3.33
r141 45 47 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.72 $Y2=3.33
r142 43 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r143 43 57 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r144 43 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r145 41 52 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.25 $Y=3.33
+ $X2=3.12 $Y2=3.33
r146 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=3.33
+ $X2=3.415 $Y2=3.33
r147 40 56 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.58 $Y=3.33 $X2=3.6
+ $Y2=3.33
r148 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=3.33
+ $X2=3.415 $Y2=3.33
r149 36 39 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=9.025 $Y=1.98
+ $X2=9.025 $Y2=2.95
r150 34 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.025 $Y=3.245
+ $X2=9.025 $Y2=3.33
r151 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.025 $Y=3.245
+ $X2=9.025 $Y2=2.95
r152 30 33 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=7.59 $Y=2.3 $X2=7.59
+ $Y2=2.92
r153 28 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=3.245
+ $X2=7.59 $Y2=3.33
r154 28 33 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.59 $Y=3.245
+ $X2=7.59 $Y2=2.92
r155 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=3.245
+ $X2=5.47 $Y2=3.33
r156 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.47 $Y=3.245
+ $X2=5.47 $Y2=2.815
r157 20 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=3.245
+ $X2=3.415 $Y2=3.33
r158 20 22 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.415 $Y=3.245
+ $X2=3.415 $Y2=2.705
r159 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=3.33
r160 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=2.9
r161 5 39 400 $w=1.7e-07 $l=1.18057e-06 $layer=licon1_PDIFF $count=1 $X=8.89
+ $Y=1.835 $X2=9.025 $Y2=2.95
r162 5 36 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.89
+ $Y=1.835 $X2=9.025 $Y2=1.98
r163 4 33 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.45
+ $Y=1.805 $X2=7.59 $Y2=2.92
r164 4 30 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=7.45
+ $Y=1.805 $X2=7.59 $Y2=2.3
r165 3 26 600 $w=1.7e-07 $l=5.4399e-07 $layer=licon1_PDIFF $count=1 $X=5.025
+ $Y=2.595 $X2=5.47 $Y2=2.815
r166 2 22 600 $w=1.7e-07 $l=4.26028e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=2.375 $X2=3.415 $Y2=2.705
r167 1 18 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.92
+ $Y=2.405 $X2=1.06 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%Q 1 2 9 11 13 15 16 17 23 24
r66 23 24 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=1.295
+ $X2=7.92 $Y2=1.665
r67 22 24 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.92 $Y=1.785
+ $X2=7.92 $Y2=1.665
r68 21 23 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=7.92 $Y=1.095 $X2=7.92
+ $Y2=1.295
r69 18 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.965 $Y=1.87
+ $X2=6.8 $Y2=1.87
r70 17 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.87
+ $X2=7.92 $Y2=1.785
r71 17 18 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=7.805 $Y=1.87
+ $X2=6.965 $Y2=1.87
r72 15 21 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.01
+ $X2=7.92 $Y2=1.095
r73 15 16 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=7.805 $Y=1.01
+ $X2=6.89 $Y2=1.01
r74 11 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=1.955 $X2=6.8
+ $Y2=1.87
r75 11 13 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=6.8 $Y=1.955
+ $X2=6.8 $Y2=2.9
r76 7 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.725 $Y=0.925
+ $X2=6.89 $Y2=1.01
r77 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.725 $Y=0.925
+ $X2=6.725 $Y2=0.43
r78 2 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.665
+ $Y=1.805 $X2=6.8 $Y2=1.95
r79 2 13 400 $w=1.7e-07 $l=1.16054e-06 $layer=licon1_PDIFF $count=1 $X=6.665
+ $Y=1.805 $X2=6.8 $Y2=2.9
r80 1 9 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=6.58
+ $Y=0.235 $X2=6.725 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%Q_N 1 2 7 8 9 10 11 12 13 22
r15 13 40 4.17552 $w=3.43e-07 $l=1.25e-07 $layer=LI1_cond $X=9.807 $Y=2.775
+ $X2=9.807 $Y2=2.9
r16 12 13 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=9.807 $Y=2.405
+ $X2=9.807 $Y2=2.775
r17 11 12 14.1968 $w=3.43e-07 $l=4.25e-07 $layer=LI1_cond $X=9.807 $Y=1.98
+ $X2=9.807 $Y2=2.405
r18 10 11 10.5223 $w=3.43e-07 $l=3.15e-07 $layer=LI1_cond $X=9.807 $Y=1.665
+ $X2=9.807 $Y2=1.98
r19 9 10 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=9.807 $Y=1.295
+ $X2=9.807 $Y2=1.665
r20 8 9 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=9.807 $Y=0.925
+ $X2=9.807 $Y2=1.295
r21 7 8 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=9.807 $Y=0.555
+ $X2=9.807 $Y2=0.925
r22 7 22 4.17552 $w=3.43e-07 $l=1.25e-07 $layer=LI1_cond $X=9.807 $Y=0.555
+ $X2=9.807 $Y2=0.43
r23 2 40 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=1.835 $X2=9.815 $Y2=2.9
r24 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=1.835 $X2=9.815 $Y2=1.98
r25 1 22 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.265 $X2=9.8 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP%VGND 1 2 3 4 5 18 22 26 32 36 39 40 42 43
+ 44 56 63 68 75 76 79 82 85
c114 76 0 2.58091e-20 $X=9.84 $Y=0
c115 18 0 1.56912e-19 $X=1.07 $Y=0.765
r116 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r117 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r119 76 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=8.88
+ $Y2=0
r120 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r121 73 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.01
+ $Y2=0
r122 73 75 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.84
+ $Y2=0
r123 72 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r124 72 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r125 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r126 69 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.68 $Y=0 $X2=7.515
+ $Y2=0
r127 69 71 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.68 $Y=0 $X2=7.92
+ $Y2=0
r128 68 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=0 $X2=9.01
+ $Y2=0
r129 68 71 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=8.845 $Y=0
+ $X2=7.92 $Y2=0
r130 67 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r131 67 80 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.52 $Y2=0
r132 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r133 64 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=0 $X2=5.375
+ $Y2=0
r134 64 66 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=5.54 $Y=0 $X2=6.96
+ $Y2=0
r135 63 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.35 $Y=0 $X2=7.515
+ $Y2=0
r136 63 66 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.35 $Y=0 $X2=6.96
+ $Y2=0
r137 58 61 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r138 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r139 56 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.375
+ $Y2=0
r140 56 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.04
+ $Y2=0
r141 55 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r142 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r143 52 55 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r144 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r145 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r146 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r147 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r148 44 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r149 44 59 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r150 44 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r151 42 54 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.12
+ $Y2=0
r152 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.31
+ $Y2=0
r153 41 58 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.6
+ $Y2=0
r154 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.31
+ $Y2=0
r155 39 47 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r156 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.03
+ $Y2=0
r157 38 51 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.2
+ $Y2=0
r158 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.03
+ $Y2=0
r159 34 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0
r160 34 36 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0.41
r161 30 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=0.085
+ $X2=7.515 $Y2=0
r162 30 32 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=7.515 $Y=0.085
+ $X2=7.515 $Y2=0.48
r163 26 28 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=5.375 $Y=0.38
+ $X2=5.375 $Y2=0.93
r164 24 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0
r165 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0.38
r166 20 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=0.085
+ $X2=3.31 $Y2=0
r167 20 22 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.31 $Y=0.085
+ $X2=3.31 $Y2=0.43
r168 16 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=0.085
+ $X2=1.03 $Y2=0
r169 16 18 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.03 $Y=0.085
+ $X2=1.03 $Y2=0.765
r170 5 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=8.865
+ $Y=0.265 $X2=9.01 $Y2=0.41
r171 4 32 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.235 $X2=7.515 $Y2=0.48
r172 3 28 182 $w=1.7e-07 $l=8.46079e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.375 $Y2=0.93
r173 3 26 182 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.375 $Y2=0.38
r174 2 22 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.31 $Y2=0.43
r175 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.555 $X2=1.07 $Y2=0.765
.ends

