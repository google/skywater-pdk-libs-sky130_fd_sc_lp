* File: sky130_fd_sc_lp__or2_2.pex.spice
* Created: Fri Aug 28 11:21:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2_2%B 2 5 7 9 12 14 17 19 20 24
c41 14 0 1.9354e-19 $X=0.27 $Y=1.46
r42 19 20 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.245 $Y=0.925
+ $X2=0.245 $Y2=1.295
r43 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=0.955 $X2=0.27 $Y2=0.955
r44 15 17 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.36 $Y=1.765
+ $X2=0.58 $Y2=1.765
r45 13 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=0.955
r46 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.46
r47 12 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.94
+ $X2=0.27 $Y2=0.955
r48 11 12 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.345 $Y=0.79
+ $X2=0.345 $Y2=0.94
r49 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.58 $Y=1.84 $X2=0.58
+ $Y2=1.765
r50 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.58 $Y=1.84 $X2=0.58
+ $Y2=2.16
r51 5 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.51 $Y=0.445
+ $X2=0.51 $Y2=0.79
r52 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.69 $X2=0.36
+ $Y2=1.765
r53 2 14 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=0.36 $Y=1.69 $X2=0.36
+ $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_2%A 3 7 9 12 13
c38 13 0 3.11076e-19 $X=0.81 $Y=1.315
c39 7 0 1.76691e-19 $X=0.94 $Y=2.16
r40 12 15 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.83 $Y=1.315
+ $X2=0.83 $Y2=1.48
r41 12 14 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.83 $Y=1.315
+ $X2=0.83 $Y2=1.15
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.315 $X2=0.81 $Y2=1.315
r43 9 13 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.305 $X2=0.81
+ $Y2=1.305
r44 7 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.94 $Y=2.16 $X2=0.94
+ $Y2=1.48
r45 3 14 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.94 $Y=0.445 $X2=0.94
+ $Y2=1.15
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_2%A_48_390# 1 2 9 13 17 21 25 27 28 31 33 34 36
+ 38 44
c86 44 0 1.98849e-19 $X=1.895 $Y=1.44
c87 28 0 1.9354e-19 $X=0.47 $Y=1.715
c88 25 0 1.76691e-19 $X=0.365 $Y=2.095
c89 9 0 1.12227e-19 $X=1.465 $Y=0.655
r90 43 44 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.465 $Y=1.44
+ $X2=1.895 $Y2=1.44
r91 39 43 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.39 $Y=1.44
+ $X2=1.465 $Y2=1.44
r92 38 40 13.3135 $w=2.52e-07 $l=2.75e-07 $layer=LI1_cond $X=1.33 $Y=1.44
+ $X2=1.33 $Y2=1.715
r93 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.39
+ $Y=1.44 $X2=1.39 $Y2=1.44
r94 36 38 8.1044 $w=2.52e-07 $l=1.79374e-07 $layer=LI1_cond $X=1.3 $Y=1.275
+ $X2=1.33 $Y2=1.44
r95 35 36 19.0404 $w=2.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=0.895 $X2=1.3
+ $Y2=1.275
r96 33 35 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.185 $Y=0.81
+ $X2=1.3 $Y2=0.895
r97 33 34 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.185 $Y=0.81
+ $X2=0.87 $Y2=0.81
r98 29 34 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.87 $Y2=0.81
r99 29 31 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.73 $Y2=0.42
r100 27 40 3.04159 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.185 $Y=1.715
+ $X2=1.33 $Y2=1.715
r101 27 28 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.185 $Y=1.715
+ $X2=0.47 $Y2=1.715
r102 23 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.365 $Y=1.8
+ $X2=0.47 $Y2=1.715
r103 23 25 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.365 $Y=1.8
+ $X2=0.365 $Y2=2.095
r104 19 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.605
+ $X2=1.895 $Y2=1.44
r105 19 21 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.895 $Y=1.605
+ $X2=1.895 $Y2=2.465
r106 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.275
+ $X2=1.895 $Y2=1.44
r107 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.895 $Y=1.275
+ $X2=1.895 $Y2=0.655
r108 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.605
+ $X2=1.465 $Y2=1.44
r109 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.465 $Y=1.605
+ $X2=1.465 $Y2=2.465
r110 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.275
+ $X2=1.465 $Y2=1.44
r111 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.465 $Y=1.275
+ $X2=1.465 $Y2=0.655
r112 2 25 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=1.95 $X2=0.365 $Y2=2.095
r113 1 31 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.235 $X2=0.725 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_2%VPWR 1 2 9 13 14 16 19 21 26 32 36
r28 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 30 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r31 27 32 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.167 $Y2=3.33
r32 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.68 $Y2=3.33
r33 26 35 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.172 $Y2=3.33
r34 26 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 21 32 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=1.167 $Y2=3.33
r37 21 23 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 19 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 19 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 19 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 14 35 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.172 $Y2=3.33
r42 14 16 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=2.48
r43 13 18 10.4482 $w=3.3e-07 $l=2.8e-07 $layer=LI1_cond $X=2.11 $Y=2.26 $X2=2.11
+ $Y2=1.98
r44 13 16 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.11 $Y=2.26
+ $X2=2.11 $Y2=2.48
r45 9 12 10.8302 $w=4.13e-07 $l=3.9e-07 $layer=LI1_cond $X=1.167 $Y=2.135
+ $X2=1.167 $Y2=2.525
r46 7 32 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.167 $Y=3.245
+ $X2=1.167 $Y2=3.33
r47 7 12 19.9942 $w=4.13e-07 $l=7.2e-07 $layer=LI1_cond $X=1.167 $Y=3.245
+ $X2=1.167 $Y2=2.525
r48 2 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.835 $X2=2.11 $Y2=1.98
r49 2 16 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=1.97
+ $Y=1.835 $X2=2.11 $Y2=2.48
r50 1 12 300 $w=1.7e-07 $l=6.82459e-07 $layer=licon1_PDIFF $count=2 $X=1.015
+ $Y=1.95 $X2=1.25 $Y2=2.525
r51 1 9 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.95 $X2=1.155 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_2%X 1 2 9 14 15 17 18 19 20
r25 20 32 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.66 $Y=2.775
+ $X2=1.66 $Y2=2.91
r26 19 20 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=2.405
+ $X2=1.66 $Y2=2.775
r27 18 19 21.2951 $w=2.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.66 $Y=1.98
+ $X2=1.66 $Y2=2.405
r28 16 17 8.02857 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.7 $Y=1.005
+ $X2=1.7 $Y2=1.14
r29 15 18 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.66 $Y=1.925
+ $X2=1.66 $Y2=1.98
r30 14 15 8.82471 $w=2.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.68 $Y=1.765
+ $X2=1.68 $Y2=1.925
r31 14 17 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.73 $Y=1.765
+ $X2=1.73 $Y2=1.14
r32 9 16 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=1.68 $Y=0.42
+ $X2=1.68 $Y2=1.005
r33 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.835 $X2=1.68 $Y2=2.91
r34 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.835 $X2=1.68 $Y2=1.98
r35 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.54
+ $Y=0.235 $X2=1.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_2%VGND 1 2 3 10 12 16 18 19 21 24 26 31 40 44
r41 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.205
+ $Y2=0
r46 32 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.68
+ $Y2=0
r47 31 43 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.172
+ $Y2=0
r48 31 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.68
+ $Y2=0
r49 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r50 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 27 37 4.33874 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.21
+ $Y2=0
r52 27 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.72
+ $Y2=0
r53 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=1.205
+ $Y2=0
r54 26 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.72
+ $Y2=0
r55 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r56 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r57 24 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r58 19 23 9.70217 $w=3.3e-07 $l=2.6e-07 $layer=LI1_cond $X=2.11 $Y=0.67 $X2=2.11
+ $Y2=0.93
r59 19 21 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.11 $Y=0.67
+ $X2=2.11 $Y2=0.38
r60 18 43 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.172 $Y2=0
r61 18 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.38
r62 14 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0
r63 14 16 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0.43
r64 10 37 3.0991 $w=2.9e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.21 $Y2=0
r65 10 12 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.445
r66 3 23 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.11 $Y2=0.93
r67 3 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.11 $Y2=0.38
r68 2 16 182 $w=1.7e-07 $l=2.73998e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.205 $Y2=0.43
r69 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.235 $X2=0.295 $Y2=0.445
.ends

