# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o2bb2ai_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o2bb2ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.450000 1.750000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.210000 1.035000 1.540000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.185000 3.275000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 1.185000 2.735000 1.585000 ;
        RECT 2.505000 1.585000 2.735000 2.995000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.676200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.255000 1.785000 0.650000 ;
        RECT 1.545000 0.650000 1.785000 1.065000 ;
        RECT 1.545000 1.065000 2.100000 1.235000 ;
        RECT 1.930000 1.235000 2.100000 1.755000 ;
        RECT 1.930000 1.755000 2.335000 1.925000 ;
        RECT 1.990000 1.925000 2.335000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.120000  0.085000 0.450000 1.040000 ;
      RECT 0.120000  1.920000 0.450000 3.245000 ;
      RECT 0.620000  1.755000 1.415000 1.925000 ;
      RECT 0.620000  1.925000 0.810000 3.075000 ;
      RECT 0.980000  2.095000 1.820000 3.245000 ;
      RECT 0.985000  0.255000 1.315000 0.820000 ;
      RECT 0.985000  0.820000 1.375000 1.040000 ;
      RECT 1.205000  1.040000 1.375000 1.405000 ;
      RECT 1.205000  1.405000 1.760000 1.675000 ;
      RECT 1.205000  1.675000 1.415000 1.755000 ;
      RECT 1.955000  0.285000 2.285000 0.725000 ;
      RECT 1.955000  0.725000 3.245000 0.895000 ;
      RECT 2.270000  0.895000 3.245000 1.015000 ;
      RECT 2.455000  0.085000 2.785000 0.555000 ;
      RECT 2.915000  1.920000 3.245000 3.245000 ;
      RECT 2.975000  0.265000 3.245000 0.725000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__o2bb2ai_1
END LIBRARY
