* File: sky130_fd_sc_lp__or2b_m.pxi.spice
* Created: Wed Sep  2 10:30:12 2020
* 
x_PM_SKY130_FD_SC_LP__OR2B_M%B_N N_B_N_M1005_g N_B_N_c_68_n N_B_N_c_69_n
+ N_B_N_c_70_n N_B_N_M1002_g N_B_N_c_71_n N_B_N_c_72_n N_B_N_c_77_n B_N B_N B_N
+ N_B_N_c_74_n PM_SKY130_FD_SC_LP__OR2B_M%B_N
x_PM_SKY130_FD_SC_LP__OR2B_M%A_27_496# N_A_27_496#_M1002_s N_A_27_496#_M1005_s
+ N_A_27_496#_M1000_g N_A_27_496#_M1001_g N_A_27_496#_c_107_n
+ N_A_27_496#_c_108_n N_A_27_496#_c_109_n N_A_27_496#_c_118_n
+ N_A_27_496#_c_119_n N_A_27_496#_c_120_n N_A_27_496#_c_110_n
+ N_A_27_496#_c_111_n N_A_27_496#_c_112_n N_A_27_496#_c_113_n
+ N_A_27_496#_c_114_n N_A_27_496#_c_115_n N_A_27_496#_c_116_n
+ PM_SKY130_FD_SC_LP__OR2B_M%A_27_496#
x_PM_SKY130_FD_SC_LP__OR2B_M%A N_A_M1007_g N_A_M1003_g N_A_c_178_n N_A_c_179_n A
+ A N_A_c_182_n PM_SKY130_FD_SC_LP__OR2B_M%A
x_PM_SKY130_FD_SC_LP__OR2B_M%A_224_378# N_A_224_378#_M1000_d
+ N_A_224_378#_M1001_s N_A_224_378#_c_218_n N_A_224_378#_M1004_g
+ N_A_224_378#_M1006_g N_A_224_378#_c_220_n N_A_224_378#_c_229_n
+ N_A_224_378#_c_221_n N_A_224_378#_c_222_n N_A_224_378#_c_223_n
+ N_A_224_378#_c_239_n N_A_224_378#_c_224_n N_A_224_378#_c_225_n
+ N_A_224_378#_c_226_n N_A_224_378#_c_227_n
+ PM_SKY130_FD_SC_LP__OR2B_M%A_224_378#
x_PM_SKY130_FD_SC_LP__OR2B_M%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_281_n
+ N_VPWR_c_282_n VPWR N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n
+ N_VPWR_c_280_n N_VPWR_c_287_n N_VPWR_c_288_n PM_SKY130_FD_SC_LP__OR2B_M%VPWR
x_PM_SKY130_FD_SC_LP__OR2B_M%X N_X_M1006_d N_X_M1004_d X X X X X X X N_X_c_315_n
+ X PM_SKY130_FD_SC_LP__OR2B_M%X
x_PM_SKY130_FD_SC_LP__OR2B_M%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_c_328_n
+ N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n VGND N_VGND_c_332_n
+ N_VGND_c_333_n N_VGND_c_334_n N_VGND_c_335_n PM_SKY130_FD_SC_LP__OR2B_M%VGND
cc_1 VNB N_B_N_c_68_n 0.0279373f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.935
cc_2 VNB N_B_N_c_69_n 0.0160209f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.935
cc_3 VNB N_B_N_c_70_n 0.0221794f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.86
cc_4 VNB N_B_N_c_71_n 0.0354394f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.45
cc_5 VNB N_B_N_c_72_n 0.00339588f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_6 VNB B_N 0.0265698f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_B_N_c_74_n 0.0199218f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_8 VNB N_A_27_496#_M1001_g 0.00761351f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_9 VNB N_A_27_496#_c_107_n 0.0178684f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.12
cc_10 VNB N_A_27_496#_c_108_n 0.0289773f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_A_27_496#_c_109_n 0.0214676f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_12 VNB N_A_27_496#_c_110_n 0.00374454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_496#_c_111_n 0.0127336f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.615
cc_14 VNB N_A_27_496#_c_112_n 0.0139271f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.665
cc_15 VNB N_A_27_496#_c_113_n 0.00883985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_496#_c_114_n 2.19657e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_496#_c_115_n 0.00245841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_496#_c_116_n 0.015631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_M1003_g 0.028558f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.935
cc_20 VNB N_A_c_178_n 0.018414f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.935
cc_21 VNB N_A_c_179_n 0.00891971f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.86
cc_22 VNB N_A_224_378#_c_218_n 0.0234872f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.935
cc_23 VNB N_A_224_378#_M1004_g 0.00739305f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.54
cc_24 VNB N_A_224_378#_c_220_n 0.0231147f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB N_A_224_378#_c_221_n 0.00104616f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_26 VNB N_A_224_378#_c_222_n 0.00409767f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_27 VNB N_A_224_378#_c_223_n 0.00977272f $X=-0.19 $Y=-0.245 $X2=0.312
+ $Y2=1.295
cc_28 VNB N_A_224_378#_c_224_n 0.0010265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_224_378#_c_225_n 0.00295859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_224_378#_c_226_n 0.020177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_224_378#_c_227_n 0.0225611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_280_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB X 0.043944f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.935
cc_34 VNB N_VGND_c_328_n 0.00752162f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.86
cc_35 VNB N_VGND_c_329_n 0.00872824f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.45
cc_36 VNB N_VGND_c_330_n 0.0323609f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VNB N_VGND_c_331_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_VGND_c_332_n 0.0207527f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_39 VNB N_VGND_c_333_n 0.0201649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_334_n 0.19705f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=2.035
cc_41 VNB N_VGND_c_335_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_B_N_M1005_g 0.0441561f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.69
cc_43 VPB N_B_N_c_72_n 0.0260351f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_44 VPB N_B_N_c_77_n 0.019505f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_45 VPB B_N 0.0195644f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_46 VPB N_A_27_496#_M1001_g 0.0242061f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_47 VPB N_A_27_496#_c_118_n 4.08405e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_27_496#_c_119_n 0.00990102f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_49 VPB N_A_27_496#_c_120_n 0.00870687f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_50 VPB N_A_27_496#_c_111_n 0.0156398f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.615
cc_51 VPB N_A_M1003_g 0.0332321f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=0.935
cc_52 VPB A 0.0168154f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_53 VPB N_A_c_182_n 0.0528549f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_54 VPB N_A_224_378#_M1004_g 0.0285771f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=0.54
cc_55 VPB N_A_224_378#_c_229_n 0.00476038f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_56 VPB N_A_224_378#_c_222_n 0.00213706f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_57 VPB N_VPWR_c_281_n 0.0159415f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=0.86
cc_58 VPB N_VPWR_c_282_n 0.0327524f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.45
cc_59 VPB N_VPWR_c_283_n 0.0178394f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_60 VPB N_VPWR_c_284_n 0.0300281f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_61 VPB N_VPWR_c_285_n 0.0197418f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.665
cc_62 VPB N_VPWR_c_280_n 0.0841121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_287_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_288_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB X 0.0160091f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=0.935
cc_66 VPB N_X_c_315_n 0.0387744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB X 0.00510377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 N_B_N_c_70_n N_A_27_496#_c_107_n 0.0112182f $X=0.88 $Y=0.86 $X2=0 $Y2=0
cc_69 N_B_N_c_74_n N_A_27_496#_c_108_n 0.00312139f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_70 N_B_N_M1005_g N_A_27_496#_c_118_n 3.52891e-19 $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_71 N_B_N_M1005_g N_A_27_496#_c_119_n 0.0167585f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_72 N_B_N_c_77_n N_A_27_496#_c_119_n 3.7612e-19 $X=0.385 $Y=2.12 $X2=0 $Y2=0
cc_73 B_N N_A_27_496#_c_119_n 0.00919128f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B_N_c_77_n N_A_27_496#_c_120_n 9.38953e-19 $X=0.385 $Y=2.12 $X2=0 $Y2=0
cc_75 B_N N_A_27_496#_c_120_n 0.0160209f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B_N_c_70_n N_A_27_496#_c_110_n 0.00463703f $X=0.88 $Y=0.86 $X2=0 $Y2=0
cc_77 N_B_N_c_71_n N_A_27_496#_c_111_n 0.0287736f $X=0.385 $Y=1.45 $X2=0 $Y2=0
cc_78 B_N N_A_27_496#_c_111_n 0.0625704f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B_N_c_68_n N_A_27_496#_c_112_n 0.00780307f $X=0.805 $Y=0.935 $X2=0 $Y2=0
cc_80 N_B_N_c_68_n N_A_27_496#_c_113_n 7.64102e-19 $X=0.805 $Y=0.935 $X2=0 $Y2=0
cc_81 N_B_N_c_69_n N_A_27_496#_c_113_n 0.00609344f $X=0.55 $Y=0.935 $X2=0 $Y2=0
cc_82 N_B_N_c_70_n N_A_27_496#_c_113_n 0.00322151f $X=0.88 $Y=0.86 $X2=0 $Y2=0
cc_83 N_B_N_c_68_n N_A_27_496#_c_114_n 0.0159441f $X=0.805 $Y=0.935 $X2=0 $Y2=0
cc_84 N_B_N_c_71_n N_A_27_496#_c_114_n 6.54369e-19 $X=0.385 $Y=1.45 $X2=0 $Y2=0
cc_85 N_B_N_c_68_n N_A_27_496#_c_116_n 0.00977133f $X=0.805 $Y=0.935 $X2=0 $Y2=0
cc_86 N_B_N_c_71_n N_A_27_496#_c_116_n 0.00312139f $X=0.385 $Y=1.45 $X2=0 $Y2=0
cc_87 N_B_N_M1005_g A 0.0051584f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_88 N_B_N_M1005_g N_VPWR_c_281_n 0.0154006f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_89 N_B_N_M1005_g N_VPWR_c_283_n 0.00444095f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_90 N_B_N_M1005_g N_VPWR_c_280_n 0.00442501f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_91 N_B_N_c_70_n N_VGND_c_328_n 0.00309057f $X=0.88 $Y=0.86 $X2=0 $Y2=0
cc_92 N_B_N_c_70_n N_VGND_c_330_n 0.00468586f $X=0.88 $Y=0.86 $X2=0 $Y2=0
cc_93 N_B_N_c_69_n N_VGND_c_334_n 0.00252916f $X=0.55 $Y=0.935 $X2=0 $Y2=0
cc_94 N_B_N_c_70_n N_VGND_c_334_n 0.00566547f $X=0.88 $Y=0.86 $X2=0 $Y2=0
cc_95 N_A_27_496#_c_109_n N_A_M1003_g 0.0649559f $X=1.35 $Y=1.53 $X2=0 $Y2=0
cc_96 N_A_27_496#_c_115_n N_A_M1003_g 4.30219e-19 $X=1.33 $Y=1.025 $X2=0 $Y2=0
cc_97 N_A_27_496#_c_116_n N_A_M1003_g 0.0181459f $X=1.33 $Y=1.025 $X2=0 $Y2=0
cc_98 N_A_27_496#_c_107_n N_A_c_178_n 0.0123877f $X=1.33 $Y=0.86 $X2=0 $Y2=0
cc_99 N_A_27_496#_c_116_n N_A_c_179_n 0.0092653f $X=1.33 $Y=1.025 $X2=0 $Y2=0
cc_100 N_A_27_496#_M1001_g A 0.00948431f $X=1.46 $Y=2.1 $X2=0 $Y2=0
cc_101 N_A_27_496#_c_119_n A 0.00968019f $X=0.66 $Y=2.385 $X2=0 $Y2=0
cc_102 N_A_27_496#_M1001_g N_A_c_182_n 0.00552254f $X=1.46 $Y=2.1 $X2=0 $Y2=0
cc_103 N_A_27_496#_M1001_g N_A_224_378#_c_229_n 0.0128565f $X=1.46 $Y=2.1 $X2=0
+ $Y2=0
cc_104 N_A_27_496#_c_109_n N_A_224_378#_c_229_n 0.00330496f $X=1.35 $Y=1.53
+ $X2=0 $Y2=0
cc_105 N_A_27_496#_c_111_n N_A_224_378#_c_229_n 0.0134175f $X=0.745 $Y=2.3 $X2=0
+ $Y2=0
cc_106 N_A_27_496#_c_115_n N_A_224_378#_c_229_n 0.0056674f $X=1.33 $Y=1.025
+ $X2=0 $Y2=0
cc_107 N_A_27_496#_c_107_n N_A_224_378#_c_221_n 0.00346782f $X=1.33 $Y=0.86
+ $X2=0 $Y2=0
cc_108 N_A_27_496#_c_108_n N_A_224_378#_c_222_n 0.00237934f $X=1.35 $Y=1.38
+ $X2=0 $Y2=0
cc_109 N_A_27_496#_c_109_n N_A_224_378#_c_222_n 0.0101118f $X=1.35 $Y=1.53 $X2=0
+ $Y2=0
cc_110 N_A_27_496#_c_115_n N_A_224_378#_c_222_n 0.0341539f $X=1.33 $Y=1.025
+ $X2=0 $Y2=0
cc_111 N_A_27_496#_c_107_n N_A_224_378#_c_239_n 0.00348663f $X=1.33 $Y=0.86
+ $X2=0 $Y2=0
cc_112 N_A_27_496#_c_113_n N_A_224_378#_c_239_n 0.00109319f $X=0.745 $Y=0.605
+ $X2=0 $Y2=0
cc_113 N_A_27_496#_c_115_n N_A_224_378#_c_239_n 0.00107353f $X=1.33 $Y=1.025
+ $X2=0 $Y2=0
cc_114 N_A_27_496#_c_116_n N_A_224_378#_c_239_n 0.00190762f $X=1.33 $Y=1.025
+ $X2=0 $Y2=0
cc_115 N_A_27_496#_c_115_n N_A_224_378#_c_224_n 0.0144695f $X=1.33 $Y=1.025
+ $X2=0 $Y2=0
cc_116 N_A_27_496#_c_116_n N_A_224_378#_c_224_n 0.00123828f $X=1.33 $Y=1.025
+ $X2=0 $Y2=0
cc_117 N_A_27_496#_c_119_n N_VPWR_c_281_n 0.022211f $X=0.66 $Y=2.385 $X2=0 $Y2=0
cc_118 N_A_27_496#_c_118_n N_VPWR_c_283_n 0.00440258f $X=0.26 $Y=2.625 $X2=0
+ $Y2=0
cc_119 N_A_27_496#_c_118_n N_VPWR_c_280_n 0.00602145f $X=0.26 $Y=2.625 $X2=0
+ $Y2=0
cc_120 N_A_27_496#_c_119_n N_VPWR_c_280_n 0.00674065f $X=0.66 $Y=2.385 $X2=0
+ $Y2=0
cc_121 N_A_27_496#_c_107_n N_VGND_c_328_n 0.00309057f $X=1.33 $Y=0.86 $X2=0
+ $Y2=0
cc_122 N_A_27_496#_c_112_n N_VGND_c_328_n 0.0134055f $X=1.245 $Y=0.945 $X2=0
+ $Y2=0
cc_123 N_A_27_496#_c_116_n N_VGND_c_328_n 0.00140352f $X=1.33 $Y=1.025 $X2=0
+ $Y2=0
cc_124 N_A_27_496#_c_113_n N_VGND_c_330_n 0.00750164f $X=0.745 $Y=0.605 $X2=0
+ $Y2=0
cc_125 N_A_27_496#_c_107_n N_VGND_c_332_n 0.00467915f $X=1.33 $Y=0.86 $X2=0
+ $Y2=0
cc_126 N_A_27_496#_c_107_n N_VGND_c_334_n 0.0052235f $X=1.33 $Y=0.86 $X2=0 $Y2=0
cc_127 N_A_27_496#_c_112_n N_VGND_c_334_n 0.00673221f $X=1.245 $Y=0.945 $X2=0
+ $Y2=0
cc_128 N_A_27_496#_c_113_n N_VGND_c_334_n 0.0104033f $X=0.745 $Y=0.605 $X2=0
+ $Y2=0
cc_129 N_A_27_496#_c_115_n N_VGND_c_334_n 0.00494472f $X=1.33 $Y=1.025 $X2=0
+ $Y2=0
cc_130 N_A_27_496#_c_116_n N_VGND_c_334_n 6.49926e-19 $X=1.33 $Y=1.025 $X2=0
+ $Y2=0
cc_131 N_A_M1003_g N_A_224_378#_c_218_n 0.0205634f $X=1.82 $Y=2.1 $X2=0 $Y2=0
cc_132 N_A_M1003_g N_A_224_378#_M1004_g 0.0218277f $X=1.82 $Y=2.1 $X2=0 $Y2=0
cc_133 N_A_M1003_g N_A_224_378#_c_229_n 0.00428419f $X=1.82 $Y=2.1 $X2=0 $Y2=0
cc_134 A N_A_224_378#_c_229_n 0.0451077f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_135 N_A_c_182_n N_A_224_378#_c_229_n 5.18935e-19 $X=1.82 $Y=2.845 $X2=0 $Y2=0
cc_136 N_A_c_178_n N_A_224_378#_c_221_n 0.00505904f $X=1.8 $Y=0.86 $X2=0 $Y2=0
cc_137 N_A_M1003_g N_A_224_378#_c_222_n 0.0199911f $X=1.82 $Y=2.1 $X2=0 $Y2=0
cc_138 N_A_M1003_g N_A_224_378#_c_223_n 0.00608549f $X=1.82 $Y=2.1 $X2=0 $Y2=0
cc_139 N_A_c_179_n N_A_224_378#_c_223_n 0.00606333f $X=1.8 $Y=1.01 $X2=0 $Y2=0
cc_140 N_A_c_178_n N_A_224_378#_c_239_n 0.00492846f $X=1.8 $Y=0.86 $X2=0 $Y2=0
cc_141 N_A_c_179_n N_A_224_378#_c_224_n 0.00254651f $X=1.8 $Y=1.01 $X2=0 $Y2=0
cc_142 N_A_M1003_g N_A_224_378#_c_225_n 0.00147242f $X=1.82 $Y=2.1 $X2=0 $Y2=0
cc_143 N_A_c_179_n N_A_224_378#_c_226_n 0.0205634f $X=1.8 $Y=1.01 $X2=0 $Y2=0
cc_144 N_A_c_178_n N_A_224_378#_c_227_n 0.0125866f $X=1.8 $Y=0.86 $X2=0 $Y2=0
cc_145 A N_VPWR_c_281_n 0.0182699f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_146 N_A_c_182_n N_VPWR_c_281_n 0.00316108f $X=1.82 $Y=2.845 $X2=0 $Y2=0
cc_147 N_A_M1003_g N_VPWR_c_282_n 0.0196543f $X=1.82 $Y=2.1 $X2=0 $Y2=0
cc_148 A N_VPWR_c_282_n 0.0486407f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_149 A N_VPWR_c_284_n 0.0229626f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_150 N_A_c_182_n N_VPWR_c_284_n 0.0116487f $X=1.82 $Y=2.845 $X2=0 $Y2=0
cc_151 A N_VPWR_c_280_n 0.0228587f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_152 N_A_c_182_n N_VPWR_c_280_n 0.0147442f $X=1.82 $Y=2.845 $X2=0 $Y2=0
cc_153 N_A_c_178_n N_VGND_c_329_n 0.00838092f $X=1.8 $Y=0.86 $X2=0 $Y2=0
cc_154 N_A_c_178_n N_VGND_c_332_n 0.00429772f $X=1.8 $Y=0.86 $X2=0 $Y2=0
cc_155 N_A_c_178_n N_VGND_c_334_n 0.00517579f $X=1.8 $Y=0.86 $X2=0 $Y2=0
cc_156 N_A_c_179_n N_VGND_c_334_n 0.00101167f $X=1.8 $Y=1.01 $X2=0 $Y2=0
cc_157 N_A_224_378#_M1004_g N_VPWR_c_282_n 0.00941023f $X=2.325 $Y=2.1 $X2=0
+ $Y2=0
cc_158 N_A_224_378#_c_220_n N_VPWR_c_282_n 0.00324989f $X=2.292 $Y=1.53 $X2=0
+ $Y2=0
cc_159 N_A_224_378#_c_225_n N_VPWR_c_282_n 0.00250835f $X=2.27 $Y=1.025 $X2=0
+ $Y2=0
cc_160 N_A_224_378#_c_229_n A_307_378# 9.39059e-19 $X=1.595 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_224_378#_c_222_n A_307_378# 4.28993e-19 $X=1.68 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_224_378#_M1004_g X 0.0153407f $X=2.325 $Y=2.1 $X2=0 $Y2=0
cc_163 N_A_224_378#_c_225_n X 0.0475752f $X=2.27 $Y=1.025 $X2=0 $Y2=0
cc_164 N_A_224_378#_c_227_n X 0.0220662f $X=2.292 $Y=0.86 $X2=0 $Y2=0
cc_165 N_A_224_378#_M1004_g N_X_c_315_n 0.00291026f $X=2.325 $Y=2.1 $X2=0 $Y2=0
cc_166 N_A_224_378#_c_220_n X 8.29358e-19 $X=2.292 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A_224_378#_c_223_n N_VGND_c_329_n 0.0125193f $X=2.185 $Y=0.945 $X2=0
+ $Y2=0
cc_168 N_A_224_378#_c_239_n N_VGND_c_329_n 0.00819513f $X=1.68 $Y=0.575 $X2=0
+ $Y2=0
cc_169 N_A_224_378#_c_225_n N_VGND_c_329_n 0.00486161f $X=2.27 $Y=1.025 $X2=0
+ $Y2=0
cc_170 N_A_224_378#_c_226_n N_VGND_c_329_n 0.00264539f $X=2.27 $Y=1.025 $X2=0
+ $Y2=0
cc_171 N_A_224_378#_c_227_n N_VGND_c_329_n 0.00519892f $X=2.292 $Y=0.86 $X2=0
+ $Y2=0
cc_172 N_A_224_378#_c_239_n N_VGND_c_332_n 0.00832525f $X=1.68 $Y=0.575 $X2=0
+ $Y2=0
cc_173 N_A_224_378#_c_227_n N_VGND_c_333_n 0.00495161f $X=2.292 $Y=0.86 $X2=0
+ $Y2=0
cc_174 N_A_224_378#_c_223_n N_VGND_c_334_n 0.00625668f $X=2.185 $Y=0.945 $X2=0
+ $Y2=0
cc_175 N_A_224_378#_c_239_n N_VGND_c_334_n 0.0114781f $X=1.68 $Y=0.575 $X2=0
+ $Y2=0
cc_176 N_A_224_378#_c_225_n N_VGND_c_334_n 0.00308366f $X=2.27 $Y=1.025 $X2=0
+ $Y2=0
cc_177 N_A_224_378#_c_227_n N_VGND_c_334_n 0.0094632f $X=2.292 $Y=0.86 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_282_n X 0.00373336f $X=2.11 $Y=2.035 $X2=0 $Y2=0
cc_179 N_VPWR_c_282_n N_X_c_315_n 0.0538605f $X=2.11 $Y=2.035 $X2=0 $Y2=0
cc_180 N_VPWR_c_285_n N_X_c_315_n 0.00803527f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_280_n N_X_c_315_n 0.00915527f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_182 X N_VGND_c_333_n 0.00592993f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_183 X N_VGND_c_334_n 0.00654783f $X=2.555 $Y=0.47 $X2=0 $Y2=0
