* File: sky130_fd_sc_lp__srsdfxtp_1.pex.spice
* Created: Wed Sep  2 10:39:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%SCE 2 3 5 8 10 11 12 14 17 22 25 26 30 35
+ 38
c102 38 0 1.10134e-19 $X=1.965 $Y=1.345
c103 35 0 1.32023e-19 $X=0.545 $Y=1.15
c104 22 0 1.70902e-19 $X=1.795 $Y=0.925
r105 39 42 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=1.345
+ $X2=1.88 $Y2=1.345
r106 38 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.345
+ $X2=1.965 $Y2=1.18
r107 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.965
+ $Y=1.345 $X2=1.965 $Y2=1.345
r108 30 39 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=1.345
+ $X2=1.965 $Y2=1.345
r109 29 35 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.525 $Y=1.15
+ $X2=0.545 $Y2=1.15
r110 29 32 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.525 $Y=1.15
+ $X2=0.27 $Y2=1.15
r111 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.15 $X2=0.525 $Y2=1.15
r112 26 28 9.76868 $w=2.81e-07 $l=2.25e-07 $layer=LI1_cond $X=0.59 $Y=0.925
+ $X2=0.59 $Y2=1.15
r113 25 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=1.18
+ $X2=1.88 $Y2=1.345
r114 24 25 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.88 $Y=1.01
+ $X2=1.88 $Y2=1.18
r115 23 26 3.67734 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=0.925
+ $X2=0.59 $Y2=0.925
r116 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=0.925
+ $X2=1.88 $Y2=1.01
r117 22 23 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.795 $Y=0.925
+ $X2=0.755 $Y2=0.925
r118 19 21 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.27 $Y=2.2
+ $X2=0.515 $Y2=2.2
r119 17 40 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.905 $Y=0.445
+ $X2=1.905 $Y2=1.18
r120 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.945 $Y=2.275
+ $X2=0.945 $Y2=2.705
r121 11 21 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.59 $Y=2.2
+ $X2=0.515 $Y2=2.2
r122 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.87 $Y=2.2
+ $X2=0.945 $Y2=2.275
r123 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.87 $Y=2.2
+ $X2=0.59 $Y2=2.2
r124 6 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=0.985
+ $X2=0.545 $Y2=1.15
r125 6 8 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.545 $Y=0.985
+ $X2=0.545 $Y2=0.445
r126 3 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.515 $Y=2.275
+ $X2=0.515 $Y2=2.2
r127 3 5 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.515 $Y=2.275
+ $X2=0.515 $Y2=2.705
r128 2 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=2.125
+ $X2=0.27 $Y2=2.2
r129 1 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.315
+ $X2=0.27 $Y2=1.15
r130 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.27 $Y=1.315 $X2=0.27
+ $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_31_477# 1 2 9 13 16 19 21 25 26 31 33
+ 35 43
c91 35 0 1.32023e-19 $X=0.75 $Y=1.72
r92 38 39 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.75 $Y=1.915 $X2=0.75
+ $Y2=1.995
r93 36 43 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.75 $Y=1.72
+ $X2=0.975 $Y2=1.72
r94 35 38 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.75 $Y=1.72
+ $X2=0.75 $Y2=1.915
r95 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.72 $X2=0.75 $Y2=1.72
r96 28 31 4.39026 $w=4.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.17 $Y=0.465
+ $X2=0.33 $Y2=0.465
r97 26 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.915
+ $X2=1.785 $Y2=2.08
r98 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.785
+ $Y=1.915 $X2=1.785 $Y2=1.915
r99 23 38 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=1.915
+ $X2=0.75 $Y2=1.915
r100 23 25 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.915 $Y=1.915
+ $X2=1.785 $Y2=1.915
r101 22 33 2.53056 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.385 $Y=1.995
+ $X2=0.235 $Y2=1.995
r102 21 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=1.995
+ $X2=0.75 $Y2=1.995
r103 21 22 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.585 $Y=1.995
+ $X2=0.385 $Y2=1.995
r104 17 33 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=2.08
+ $X2=0.235 $Y2=1.995
r105 17 19 17.2866 $w=2.98e-07 $l=4.5e-07 $layer=LI1_cond $X=0.235 $Y=2.08
+ $X2=0.235 $Y2=2.53
r106 16 33 3.91525 $w=2.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.17 $Y=1.91
+ $X2=0.235 $Y2=1.995
r107 15 28 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.17 $Y=0.675
+ $X2=0.17 $Y2=0.465
r108 15 16 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=0.17 $Y=0.675
+ $X2=0.17 $Y2=1.91
r109 13 47 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.765 $Y=2.705
+ $X2=1.765 $Y2=2.08
r110 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.555
+ $X2=0.975 $Y2=1.72
r111 7 9 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.975 $Y=1.555
+ $X2=0.975 $Y2=0.445
r112 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=2.385 $X2=0.3 $Y2=2.53
r113 1 31 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.33 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%D 3 7 9 12 13
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.51
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.18
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.425
+ $Y=1.345 $X2=1.425 $Y2=1.345
r39 9 13 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.2 $Y=1.345
+ $X2=1.425 $Y2=1.345
r40 7 14 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.365 $Y=0.445
+ $X2=1.365 $Y2=1.18
r41 3 15 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=1.335 $Y=2.705
+ $X2=1.335 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%SCD 3 7 13 15 18 19 20
c55 20 0 3.51957e-20 $X=2.325 $Y=1.75
c56 19 0 1.4124e-19 $X=2.325 $Y=1.915
c57 13 0 1.35707e-19 $X=2.415 $Y=0.895
c58 7 0 1.25447e-19 $X=2.295 $Y=0.445
r59 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.915
+ $X2=2.325 $Y2=2.08
r60 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.915
+ $X2=2.325 $Y2=1.75
r61 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=1.915 $X2=2.325 $Y2=1.915
r62 15 19 4.75383 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=1.95
+ $X2=2.325 $Y2=1.95
r63 11 13 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.295 $Y=0.895
+ $X2=2.415 $Y2=0.895
r64 9 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.415 $Y=0.97
+ $X2=2.415 $Y2=0.895
r65 9 20 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.415 $Y=0.97
+ $X2=2.415 $Y2=1.75
r66 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.295 $Y=0.82
+ $X2=2.295 $Y2=0.895
r67 5 7 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.295 $Y=0.82
+ $X2=2.295 $Y2=0.445
r68 3 21 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.235 $Y=2.705
+ $X2=2.235 $Y2=2.08
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_570_47# 1 2 7 9 13 15 17 18 20 21 23 24
+ 26 28 30 33 34 37 40 43 44 45 47 48 49 51 52 55 56 57 60 61 67 75 77 78 82 85
+ 89 96
c247 96 0 1.25046e-19 $X=6.52 $Y=1.26
c248 82 0 1.14482e-19 $X=6.455 $Y=1.26
c249 77 0 1.25405e-19 $X=3.57 $Y=0.42
c250 67 0 1.25447e-19 $X=3.17 $Y=0.465
c251 61 0 8.6426e-20 $X=9.255 $Y=1.56
c252 37 0 5.39634e-20 $X=3.76 $Y=2.57
c253 30 0 1.06176e-19 $X=3.085 $Y=1.98
c254 15 0 1.8374e-20 $X=4.545 $Y=2.54
c255 13 0 5.25296e-20 $X=4.285 $Y=0.905
c256 9 0 1.32899e-19 $X=4.47 $Y=2.465
r257 83 96 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=6.455 $Y=1.26
+ $X2=6.52 $Y2=1.26
r258 83 93 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=6.455 $Y=1.26
+ $X2=6.16 $Y2=1.26
r259 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.455
+ $Y=1.26 $X2=6.455 $Y2=1.26
r260 79 82 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.035 $Y=1.26
+ $X2=6.455 $Y2=1.26
r261 76 85 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=3.405 $Y=0.42
+ $X2=3.405 $Y2=0.25
r262 75 77 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0.42
+ $X2=3.57 $Y2=0.42
r263 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.405
+ $Y=0.42 $X2=3.405 $Y2=0.42
r264 67 75 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.17 $Y=0.42
+ $X2=3.405 $Y2=0.42
r265 66 67 2.89329 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.465
+ $X2=3.17 $Y2=0.465
r266 64 66 2.60672 $w=4.18e-07 $l=9.5e-08 $layer=LI1_cond $X=2.99 $Y=0.465
+ $X2=3.085 $Y2=0.465
r267 61 100 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.255 $Y=1.56
+ $X2=9.255 $Y2=1.725
r268 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.255
+ $Y=1.56 $X2=9.255 $Y2=1.56
r269 58 60 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=9.255 $Y=1.255
+ $X2=9.255 $Y2=1.56
r270 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.09 $Y=1.17
+ $X2=9.255 $Y2=1.255
r271 56 57 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=9.09 $Y=1.17
+ $X2=7.78 $Y2=1.17
r272 55 57 8.37092 $w=1.7e-07 $l=2.38747e-07 $layer=LI1_cond $X=7.58 $Y=1.085
+ $X2=7.78 $Y2=1.17
r273 54 55 19.0153 $w=3.98e-07 $l=6.6e-07 $layer=LI1_cond $X=7.58 $Y=0.425
+ $X2=7.58 $Y2=1.085
r274 53 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=0.34
+ $X2=6.035 $Y2=0.34
r275 52 54 8.37092 $w=1.7e-07 $l=2.38747e-07 $layer=LI1_cond $X=7.38 $Y=0.34
+ $X2=7.58 $Y2=0.425
r276 52 53 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=7.38 $Y=0.34
+ $X2=6.12 $Y2=0.34
r277 51 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.035 $Y=1.095
+ $X2=6.035 $Y2=1.26
r278 50 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.035 $Y=0.425
+ $X2=6.035 $Y2=0.34
r279 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.035 $Y=0.425
+ $X2=6.035 $Y2=1.095
r280 48 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=0.34
+ $X2=6.035 $Y2=0.34
r281 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.95 $Y=0.34
+ $X2=5.44 $Y2=0.34
r282 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.355 $Y=0.425
+ $X2=5.44 $Y2=0.34
r283 46 47 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.355 $Y=0.425
+ $X2=5.355 $Y2=0.615
r284 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.27 $Y=0.7
+ $X2=5.355 $Y2=0.615
r285 44 45 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.27 $Y=0.7
+ $X2=4.575 $Y2=0.7
r286 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=0.615
+ $X2=4.575 $Y2=0.7
r287 42 43 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.49 $Y=0.425
+ $X2=4.49 $Y2=0.615
r288 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.405 $Y=0.34
+ $X2=4.49 $Y2=0.425
r289 40 77 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.405 $Y=0.34
+ $X2=3.57 $Y2=0.34
r290 38 89 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=3.76 $Y=2.57
+ $X2=3.76 $Y2=2.465
r291 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=2.57 $X2=3.76 $Y2=2.57
r292 35 73 3.01144 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.455 $Y=2.57
+ $X2=3.33 $Y2=2.57
r293 35 37 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.455 $Y=2.57
+ $X2=3.76 $Y2=2.57
r294 34 73 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=2.405
+ $X2=3.33 $Y2=2.57
r295 33 68 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.33 $Y=2.065
+ $X2=3.085 $Y2=2.065
r296 33 34 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.33 $Y=2.15
+ $X2=3.33 $Y2=2.405
r297 30 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=1.98
+ $X2=3.085 $Y2=2.065
r298 29 66 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.085 $Y=0.675
+ $X2=3.085 $Y2=0.465
r299 29 30 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=3.085 $Y=0.675
+ $X2=3.085 $Y2=1.98
r300 28 100 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.165 $Y=1.965
+ $X2=9.165 $Y2=1.725
r301 24 28 35.9872 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=9.165 $Y=2.09
+ $X2=9.165 $Y2=1.965
r302 24 26 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.165 $Y=2.09
+ $X2=9.165 $Y2=2.595
r303 21 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.52 $Y=1.095
+ $X2=6.52 $Y2=1.26
r304 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.52 $Y=1.095
+ $X2=6.52 $Y2=0.665
r305 18 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.095
+ $X2=6.16 $Y2=1.26
r306 18 20 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.16 $Y=1.095
+ $X2=6.16 $Y2=0.665
r307 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.545 $Y=2.54
+ $X2=4.545 $Y2=2.86
r308 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.285 $Y=0.325
+ $X2=4.285 $Y2=0.905
r309 10 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=2.465
+ $X2=3.76 $Y2=2.465
r310 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.47 $Y=2.465
+ $X2=4.545 $Y2=2.54
r311 9 10 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.47 $Y=2.465
+ $X2=3.925 $Y2=2.465
r312 8 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=0.25
+ $X2=3.405 $Y2=0.25
r313 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.21 $Y=0.25
+ $X2=4.285 $Y2=0.325
r314 7 8 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.21 $Y=0.25 $X2=3.57
+ $Y2=0.25
r315 2 73 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=2.385 $X2=3.29 $Y2=2.57
r316 1 64 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.235 $X2=2.99 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_914_245# 1 2 9 12 16 17 19 20 23 26 27
+ 28 31 34 35 41
c102 34 0 1.25046e-19 $X=5.695 $Y=1.04
c103 31 0 1.5358e-19 $X=5.455 $Y=2.325
c104 20 0 7.12721e-20 $X=4.9 $Y=1.04
c105 17 0 7.06589e-20 $X=4.735 $Y=1.39
r106 35 38 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.5 $Y=2.28 $X2=6.5
+ $Y2=2.42
r107 31 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=2.325
+ $X2=5.455 $Y2=2.49
r108 30 33 7.90247 $w=3.48e-07 $l=2.4e-07 $layer=LI1_cond $X=5.455 $Y=2.28
+ $X2=5.695 $Y2=2.28
r109 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=2.325 $X2=5.455 $Y2=2.325
r110 28 33 2.79879 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=5.78 $Y=2.28
+ $X2=5.695 $Y2=2.28
r111 27 35 0.354467 $w=3.5e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=2.28
+ $X2=6.5 $Y2=2.28
r112 27 28 18.2745 $w=3.48e-07 $l=5.55e-07 $layer=LI1_cond $X=6.335 $Y=2.28
+ $X2=5.78 $Y2=2.28
r113 26 33 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.695 $Y=2.105
+ $X2=5.695 $Y2=2.28
r114 25 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=1.125
+ $X2=5.695 $Y2=1.04
r115 25 26 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.695 $Y=1.125
+ $X2=5.695 $Y2=2.105
r116 21 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=0.955
+ $X2=5.695 $Y2=1.04
r117 21 23 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.695 $Y=0.955
+ $X2=5.695 $Y2=0.8
r118 19 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.61 $Y=1.04
+ $X2=5.695 $Y2=1.04
r119 19 20 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.61 $Y=1.04
+ $X2=4.9 $Y2=1.04
r120 17 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.39
+ $X2=4.735 $Y2=1.225
r121 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.735
+ $Y=1.39 $X2=4.735 $Y2=1.39
r122 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.735 $Y=1.125
+ $X2=4.9 $Y2=1.04
r123 14 16 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.735 $Y=1.125
+ $X2=4.735 $Y2=1.39
r124 12 45 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.365 $Y=2.86
+ $X2=5.365 $Y2=2.49
r125 9 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.675 $Y=0.905
+ $X2=4.675 $Y2=1.225
r126 2 38 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=2.125 $X2=6.5 $Y2=2.42
r127 1 23 182 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_NDIFF $count=1 $X=5.555
+ $Y=0.345 $X2=5.695 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_786_139# 1 2 9 11 13 14 15 18 20 21 23
+ 24 26 30 33 35 36 40 45 46 52
c143 26 0 1.8374e-20 $X=5.995 $Y=2.71
c144 24 0 1.5358e-19 $X=5.11 $Y=1.81
c145 21 0 1.32899e-19 $X=4.235 $Y=1.81
c146 20 0 7.06589e-20 $X=4.595 $Y=1.81
c147 9 0 1.14482e-19 $X=5.48 $Y=0.665
r148 46 56 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=8.175 $Y=2.91
+ $X2=8.175 $Y2=3.15
r149 45 48 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.175 $Y=2.91
+ $X2=8.175 $Y2=2.99
r150 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.175
+ $Y=2.91 $X2=8.175 $Y2=2.91
r151 40 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.08 $Y=2.71
+ $X2=6.08 $Y2=2.99
r152 36 38 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.76 $Y=2.71
+ $X2=4.76 $Y2=2.85
r153 34 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.165 $Y=2.99
+ $X2=6.08 $Y2=2.99
r154 33 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.01 $Y=2.99
+ $X2=8.175 $Y2=2.99
r155 33 34 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=8.01 $Y=2.99
+ $X2=6.165 $Y2=2.99
r156 31 52 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.275 $Y=1.425
+ $X2=5.48 $Y2=1.425
r157 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.275
+ $Y=1.425 $X2=5.275 $Y2=1.425
r158 28 30 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=5.275 $Y=1.725
+ $X2=5.275 $Y2=1.425
r159 27 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=2.71
+ $X2=4.76 $Y2=2.71
r160 26 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=2.71
+ $X2=6.08 $Y2=2.71
r161 26 27 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=5.995 $Y=2.71
+ $X2=4.925 $Y2=2.71
r162 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=1.81
+ $X2=4.76 $Y2=1.81
r163 24 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.11 $Y=1.81
+ $X2=5.275 $Y2=1.725
r164 24 25 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.11 $Y=1.81
+ $X2=4.925 $Y2=1.81
r165 23 36 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=2.625
+ $X2=4.76 $Y2=2.71
r166 22 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=1.895
+ $X2=4.76 $Y2=1.81
r167 22 23 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=4.76 $Y=1.895
+ $X2=4.76 $Y2=2.625
r168 20 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=1.81
+ $X2=4.76 $Y2=1.81
r169 20 21 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.595 $Y=1.81
+ $X2=4.235 $Y2=1.81
r170 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.11 $Y=1.725
+ $X2=4.235 $Y2=1.81
r171 16 18 37.8001 $w=2.48e-07 $l=8.2e-07 $layer=LI1_cond $X=4.11 $Y=1.725
+ $X2=4.11 $Y2=0.905
r172 14 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.01 $Y=3.15
+ $X2=8.175 $Y2=3.15
r173 14 15 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=8.01 $Y=3.15
+ $X2=6.35 $Y2=3.15
r174 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.275 $Y=3.075
+ $X2=6.35 $Y2=3.15
r175 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.275 $Y=3.075
+ $X2=6.275 $Y2=2.545
r176 7 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.48 $Y=1.26
+ $X2=5.48 $Y2=1.425
r177 7 9 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.48 $Y=1.26
+ $X2=5.48 $Y2=0.665
r178 2 38 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=4.62
+ $Y=2.65 $X2=4.76 $Y2=2.85
r179 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.695 $X2=4.07 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_540_21# 1 2 9 12 15 17 21 23 27 29 31
+ 33 35 36 38 40 43 45 49 51 52 53 54 58 59 62 66 68 70 73 75 80 81 82 84 88
c244 82 0 1.20102e-19 $X=10.6 $Y=2.085
c245 62 0 8.6426e-20 $X=10.515 $Y=2.085
c246 52 0 1.60139e-19 $X=3.855 $Y=1.857
c247 21 0 1.25405e-19 $X=3.855 $Y=0.905
r248 84 86 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=10.81 $Y=1.13
+ $X2=10.81 $Y2=1.245
r249 80 81 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=9.235 $Y=2.047
+ $X2=9.405 $Y2=2.047
r250 76 88 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=8.175 $Y=1.93
+ $X2=8.175 $Y2=1.71
r251 75 78 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.175 $Y=1.93
+ $X2=8.175 $Y2=2.01
r252 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.175
+ $Y=1.93 $X2=8.175 $Y2=1.93
r253 72 73 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.265 $Y=1.33
+ $X2=11.265 $Y2=2
r254 71 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.975 $Y=1.245
+ $X2=10.81 $Y2=1.245
r255 70 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.18 $Y=1.245
+ $X2=11.265 $Y2=1.33
r256 70 71 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.18 $Y=1.245
+ $X2=10.975 $Y2=1.245
r257 69 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.685 $Y=2.085
+ $X2=10.6 $Y2=2.085
r258 68 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.18 $Y=2.085
+ $X2=11.265 $Y2=2
r259 68 69 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=11.18 $Y=2.085
+ $X2=10.685 $Y2=2.085
r260 64 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.6 $Y=2.17
+ $X2=10.6 $Y2=2.085
r261 64 66 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=10.6 $Y=2.17
+ $X2=10.6 $Y2=2.405
r262 62 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.515 $Y=2.085
+ $X2=10.6 $Y2=2.085
r263 62 81 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=10.515 $Y=2.085
+ $X2=9.405 $Y2=2.085
r264 61 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.34 $Y=2.01
+ $X2=8.175 $Y2=2.01
r265 61 80 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=8.34 $Y=2.01
+ $X2=9.235 $Y2=2.01
r266 54 56 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.87 $Y=1.71
+ $X2=5.87 $Y2=1.875
r267 47 49 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.775 $Y=0.9
+ $X2=2.975 $Y2=0.9
r268 46 59 12.05 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=7.255 $Y=1.71
+ $X2=7.162 $Y2=1.71
r269 45 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.01 $Y=1.71
+ $X2=8.175 $Y2=1.71
r270 45 46 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=8.01 $Y=1.71
+ $X2=7.255 $Y2=1.71
r271 41 59 12.05 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=7.18 $Y=1.635
+ $X2=7.162 $Y2=1.71
r272 41 43 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.18 $Y=1.635
+ $X2=7.18 $Y2=0.775
r273 38 59 12.05 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=7.145 $Y=1.785
+ $X2=7.162 $Y2=1.71
r274 38 40 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.145 $Y=1.785
+ $X2=7.145 $Y2=2.315
r275 37 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.86 $Y=1.71
+ $X2=6.785 $Y2=1.71
r276 36 59 12.05 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=7.07 $Y=1.71
+ $X2=7.162 $Y2=1.71
r277 36 37 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.07 $Y=1.71
+ $X2=6.86 $Y2=1.71
r278 33 58 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.785 $Y=1.785
+ $X2=6.785 $Y2=1.71
r279 33 35 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.785 $Y=1.785
+ $X2=6.785 $Y2=2.315
r280 32 54 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.945 $Y=1.71
+ $X2=5.87 $Y2=1.71
r281 31 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.71 $Y=1.71
+ $X2=6.785 $Y2=1.71
r282 31 32 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.71 $Y=1.71
+ $X2=5.945 $Y2=1.71
r283 30 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.05 $Y=1.875
+ $X2=4.975 $Y2=1.875
r284 29 56 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.795 $Y=1.875
+ $X2=5.87 $Y2=1.875
r285 29 30 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=5.795 $Y=1.875
+ $X2=5.05 $Y2=1.875
r286 25 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.975 $Y=1.95
+ $X2=4.975 $Y2=1.875
r287 25 27 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.975 $Y=1.95
+ $X2=4.975 $Y2=2.86
r288 24 52 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=3.93 $Y=1.875
+ $X2=3.855 $Y2=1.857
r289 23 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.9 $Y=1.875
+ $X2=4.975 $Y2=1.875
r290 23 24 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=4.9 $Y=1.875
+ $X2=3.93 $Y2=1.875
r291 19 52 5.30422 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=3.855 $Y=1.765
+ $X2=3.855 $Y2=1.857
r292 19 21 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.855 $Y=1.765
+ $X2=3.855 $Y2=0.905
r293 18 51 5.30422 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.15 $Y=1.84
+ $X2=3.025 $Y2=1.84
r294 17 52 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=3.78 $Y=1.84
+ $X2=3.855 $Y2=1.857
r295 17 18 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.78 $Y=1.84
+ $X2=3.15 $Y2=1.84
r296 13 51 20.4101 $w=1.5e-07 $l=9.68246e-08 $layer=POLY_cond $X=3.075 $Y=1.915
+ $X2=3.025 $Y2=1.84
r297 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.075 $Y=1.915
+ $X2=3.075 $Y2=2.705
r298 12 51 20.4101 $w=1.5e-07 $l=9.68246e-08 $layer=POLY_cond $X=2.975 $Y=1.765
+ $X2=3.025 $Y2=1.84
r299 11 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.975 $Y=0.975
+ $X2=2.975 $Y2=0.9
r300 11 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.975 $Y=0.975
+ $X2=2.975 $Y2=1.765
r301 7 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.775 $Y=0.825
+ $X2=2.775 $Y2=0.9
r302 7 9 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.775 $Y=0.825
+ $X2=2.775 $Y2=0.445
r303 2 66 600 $w=1.7e-07 $l=4.25852e-07 $layer=licon1_PDIFF $count=1 $X=10.325
+ $Y=2.095 $X2=10.6 $Y2=2.405
r304 1 84 182 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=1 $X=10.665
+ $Y=0.89 $X2=10.81 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_1319_69# 1 2 3 12 16 18 20 21 22 25 28
+ 31 33 35 40 42 46 47 49 53 54 56 57 60 63 64 65 67 68 69 71 72 74 75 80 82 83
+ 87 90 94
c216 82 0 1.97937e-19 $X=7.282 $Y=1.51
c217 49 0 1.91338e-19 $X=7.125 $Y=1.425
r218 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.715
+ $Y=1.59 $X2=8.715 $Y2=1.59
r219 83 86 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.715 $Y=1.51
+ $X2=8.715 $Y2=1.59
r220 78 80 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=6.965 $Y=0.76
+ $X2=7.125 $Y2=0.76
r221 75 94 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.43 $Y=2.91
+ $X2=12.43 $Y2=2.745
r222 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.43
+ $Y=2.91 $X2=12.43 $Y2=2.91
r223 72 74 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=11.705 $Y=2.91
+ $X2=12.43 $Y2=2.91
r224 71 72 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.62 $Y=2.745
+ $X2=11.705 $Y2=2.91
r225 70 71 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.62 $Y=2.51
+ $X2=11.62 $Y2=2.745
r226 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.535 $Y=2.425
+ $X2=11.62 $Y2=2.51
r227 68 69 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.535 $Y=2.425
+ $X2=11.025 $Y2=2.425
r228 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.94 $Y=2.51
+ $X2=11.025 $Y2=2.425
r229 66 67 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.94 $Y=2.51
+ $X2=10.94 $Y2=2.905
r230 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.855 $Y=2.99
+ $X2=10.94 $Y2=2.905
r231 64 65 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.855 $Y=2.99
+ $X2=10.345 $Y2=2.99
r232 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.26 $Y=2.905
+ $X2=10.345 $Y2=2.99
r233 62 63 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.26 $Y=2.51
+ $X2=10.26 $Y2=2.905
r234 61 90 8.61065 $w=1.7e-07 $l=1.83016e-07 $layer=LI1_cond $X=9.065 $Y=2.425
+ $X2=8.9 $Y2=2.387
r235 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.175 $Y=2.425
+ $X2=10.26 $Y2=2.51
r236 60 61 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=10.175 $Y=2.425
+ $X2=9.065 $Y2=2.425
r237 56 90 8.61065 $w=1.7e-07 $l=1.82565e-07 $layer=LI1_cond $X=8.735 $Y=2.35
+ $X2=8.9 $Y2=2.387
r238 56 57 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=8.735 $Y=2.35
+ $X2=7.525 $Y2=2.35
r239 55 82 2.76166 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=7.525 $Y=1.51
+ $X2=7.282 $Y2=1.51
r240 54 83 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.55 $Y=1.51
+ $X2=8.715 $Y2=1.51
r241 54 55 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=8.55 $Y=1.51
+ $X2=7.525 $Y2=1.51
r242 51 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.36 $Y=2.265
+ $X2=7.525 $Y2=2.35
r243 51 53 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.36 $Y=2.265
+ $X2=7.36 $Y2=2.04
r244 50 82 3.70735 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=7.36 $Y=1.595
+ $X2=7.282 $Y2=1.51
r245 50 53 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.36 $Y=1.595
+ $X2=7.36 $Y2=2.04
r246 49 82 3.70735 $w=2.5e-07 $l=1.94921e-07 $layer=LI1_cond $X=7.125 $Y=1.425
+ $X2=7.282 $Y2=1.51
r247 48 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=0.925
+ $X2=7.125 $Y2=0.76
r248 48 49 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=7.125 $Y=0.925
+ $X2=7.125 $Y2=1.425
r249 45 46 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=12.865 $Y=0.925
+ $X2=12.865 $Y2=1.075
r250 42 44 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=12.34 $Y=1.65
+ $X2=12.34 $Y2=1.91
r251 39 87 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=8.715 $Y=1.395
+ $X2=8.715 $Y2=1.59
r252 39 40 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.715 $Y=1.32
+ $X2=8.805 $Y2=1.32
r253 36 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.445 $Y=1.32
+ $X2=8.715 $Y2=1.32
r254 33 47 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=12.88 $Y=1.725
+ $X2=12.865 $Y2=1.65
r255 33 35 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.88 $Y=1.725
+ $X2=12.88 $Y2=2.155
r256 31 45 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.88 $Y=0.495
+ $X2=12.88 $Y2=0.925
r257 28 47 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=12.85 $Y=1.575
+ $X2=12.865 $Y2=1.65
r258 28 46 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=12.85 $Y=1.575
+ $X2=12.85 $Y2=1.075
r259 26 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.415 $Y=1.65
+ $X2=12.34 $Y2=1.65
r260 25 47 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.775 $Y=1.65
+ $X2=12.865 $Y2=1.65
r261 25 26 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=12.775 $Y=1.65
+ $X2=12.415 $Y2=1.65
r262 23 44 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.34 $Y=1.985
+ $X2=12.34 $Y2=1.91
r263 23 94 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=12.34 $Y=1.985
+ $X2=12.34 $Y2=2.745
r264 21 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.265 $Y=1.91
+ $X2=12.34 $Y2=1.91
r265 21 22 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=12.265 $Y=1.91
+ $X2=11.67 $Y2=1.91
r266 18 22 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=11.545 $Y=1.985
+ $X2=11.67 $Y2=1.91
r267 18 20 117.608 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=11.545 $Y=1.985
+ $X2=11.545 $Y2=2.595
r268 14 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.805 $Y=1.245
+ $X2=8.805 $Y2=1.32
r269 14 16 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.805 $Y=1.245
+ $X2=8.805 $Y2=0.835
r270 10 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.445 $Y=1.245
+ $X2=8.445 $Y2=1.32
r271 10 12 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.445 $Y=1.245
+ $X2=8.445 $Y2=0.835
r272 3 90 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=8.755
+ $Y=2.095 $X2=8.9 $Y2=2.43
r273 2 53 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.22
+ $Y=1.895 $X2=7.36 $Y2=2.04
r274 1 78 182 $w=1.7e-07 $l=5.70767e-07 $layer=licon1_NDIFF $count=1 $X=6.595
+ $Y=0.345 $X2=6.965 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_1493_21# 1 2 9 11 12 15 17 20 21 23 26
+ 27 30 32 34 37 38 39 42 45 52 53 54 58 63
c154 63 0 1.30215e-19 $X=9.705 $Y=0.955
c155 58 0 1.67049e-19 $X=11.23 $Y=0.68
c156 39 0 1.1974e-19 $X=11.69 $Y=2.085
c157 9 0 3.89275e-19 $X=7.54 $Y=0.775
r158 58 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.23 $Y=0.68
+ $X2=11.23 $Y2=0.905
r159 54 56 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=10.39 $Y=0.68
+ $X2=10.39 $Y2=0.83
r160 51 63 9.45098 $w=2.55e-07 $l=5e-08 $layer=POLY_cond $X=9.755 $Y=0.955
+ $X2=9.705 $Y2=0.955
r161 50 53 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=0.932
+ $X2=9.92 $Y2=0.932
r162 50 52 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=0.932
+ $X2=9.59 $Y2=0.932
r163 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.755
+ $Y=0.955 $X2=9.755 $Y2=0.955
r164 45 47 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.135 $Y=0.75
+ $X2=9.135 $Y2=0.83
r165 40 42 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=12 $Y=2.17 $X2=12
+ $Y2=2.325
r166 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.875 $Y=2.085
+ $X2=12 $Y2=2.17
r167 38 39 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=11.875 $Y=2.085
+ $X2=11.69 $Y2=2.085
r168 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.605 $Y=2
+ $X2=11.69 $Y2=2.085
r169 36 37 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=11.605 $Y=0.99
+ $X2=11.605 $Y2=2
r170 35 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.315 $Y=0.905
+ $X2=11.23 $Y2=0.905
r171 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.52 $Y=0.905
+ $X2=11.605 $Y2=0.99
r172 34 35 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.52 $Y=0.905
+ $X2=11.315 $Y2=0.905
r173 33 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.475 $Y=0.68
+ $X2=10.39 $Y2=0.68
r174 32 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.145 $Y=0.68
+ $X2=11.23 $Y2=0.68
r175 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.145 $Y=0.68
+ $X2=10.475 $Y2=0.68
r176 30 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=0.83
+ $X2=10.39 $Y2=0.83
r177 30 53 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.305 $Y=0.83
+ $X2=9.92 $Y2=0.83
r178 29 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.3 $Y=0.83
+ $X2=9.135 $Y2=0.83
r179 29 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.3 $Y=0.83
+ $X2=9.59 $Y2=0.83
r180 24 63 15.178 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.705 $Y=1.12
+ $X2=9.705 $Y2=0.955
r181 24 27 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=9.705 $Y=1.12
+ $X2=9.705 $Y2=1.965
r182 21 27 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=9.655 $Y=2.09
+ $X2=9.655 $Y2=1.965
r183 21 23 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.655 $Y=2.09
+ $X2=9.655 $Y2=2.595
r184 20 63 51.9804 $w=2.55e-07 $l=3.47851e-07 $layer=POLY_cond $X=9.43 $Y=0.79
+ $X2=9.705 $Y2=0.955
r185 19 20 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=9.43 $Y=0.255
+ $X2=9.43 $Y2=0.79
r186 18 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.975 $Y=0.18
+ $X2=7.9 $Y2=0.18
r187 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.355 $Y=0.18
+ $X2=9.43 $Y2=0.255
r188 17 18 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=9.355 $Y=0.18
+ $X2=7.975 $Y2=0.18
r189 13 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.9 $Y=0.255
+ $X2=7.9 $Y2=0.18
r190 13 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.9 $Y=0.255
+ $X2=7.9 $Y2=0.775
r191 11 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.825 $Y=0.18
+ $X2=7.9 $Y2=0.18
r192 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.825 $Y=0.18
+ $X2=7.615 $Y2=0.18
r193 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.54 $Y=0.255
+ $X2=7.615 $Y2=0.18
r194 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.54 $Y=0.255
+ $X2=7.54 $Y2=0.775
r195 2 42 600 $w=1.7e-07 $l=3.8833e-07 $layer=licon1_PDIFF $count=1 $X=11.67
+ $Y=2.095 $X2=11.96 $Y2=2.325
r196 1 45 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=8.88
+ $Y=0.625 $X2=9.135 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%SLEEP_B 3 7 9 11 12 13 19 20 29 31
c66 19 0 1.30215e-19 $X=10.135 $Y=0.415
c67 7 0 1.67049e-19 $X=11.53 $Y=1.1
r68 27 29 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=11.685 $Y=0.485
+ $X2=11.89 $Y2=0.485
r69 24 27 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=11.53 $Y=0.485
+ $X2=11.685 $Y2=0.485
r70 20 31 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=11.685 $Y=0.485
+ $X2=11.685 $Y2=0.34
r71 20 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.685
+ $Y=0.485 $X2=11.685 $Y2=0.485
r72 16 19 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=9.97 $Y=0.415
+ $X2=10.135 $Y2=0.415
r73 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.97
+ $Y=0.415 $X2=9.97 $Y2=0.415
r74 13 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.52 $Y=0.34
+ $X2=11.685 $Y2=0.34
r75 13 19 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=11.52 $Y=0.34
+ $X2=10.135 $Y2=0.34
r76 12 17 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=10.175 $Y=0.415
+ $X2=9.97 $Y2=0.415
r77 9 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.89 $Y=0.65
+ $X2=11.89 $Y2=0.485
r78 9 11 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=11.89 $Y=0.65 $X2=11.89
+ $Y2=1.1
r79 5 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.53 $Y=0.65
+ $X2=11.53 $Y2=0.485
r80 5 7 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=11.53 $Y=0.65
+ $X2=11.53 $Y2=1.1
r81 1 12 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=10.25 $Y=0.58
+ $X2=10.175 $Y2=0.415
r82 1 3 940.926 $w=1.5e-07 $l=1.835e-06 $layer=POLY_cond $X=10.25 $Y=0.58
+ $X2=10.25 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%CLK 3 7 9 10 11 18
c49 18 0 1.20102e-19 $X=10.95 $Y=1.637
c50 3 0 1.1974e-19 $X=10.95 $Y=2.415
r51 16 18 16.814 $w=3.01e-07 $l=1.05e-07 $layer=POLY_cond $X=10.845 $Y=1.637
+ $X2=10.95 $Y2=1.637
r52 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.845
+ $Y=1.665 $X2=10.845 $Y2=1.665
r53 10 11 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=10.32 $Y=1.665
+ $X2=10.8 $Y2=1.665
r54 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.84 $Y=1.665
+ $X2=10.32 $Y2=1.665
r55 5 18 30.4252 $w=3.01e-07 $l=2.70821e-07 $layer=POLY_cond $X=11.14 $Y=1.445
+ $X2=10.95 $Y2=1.637
r56 5 7 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=11.14 $Y=1.445
+ $X2=11.14 $Y2=1.1
r57 1 18 19.0468 $w=1.5e-07 $l=1.93e-07 $layer=POLY_cond $X=10.95 $Y=1.83
+ $X2=10.95 $Y2=1.637
r58 1 3 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=10.95 $Y=1.83
+ $X2=10.95 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_2504_57# 1 2 9 13 17 21 25 26 28
r57 26 31 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=13.332 $Y=1.48
+ $X2=13.332 $Y2=1.645
r58 26 30 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=13.332 $Y=1.48
+ $X2=13.332 $Y2=1.315
r59 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.33
+ $Y=1.48 $X2=13.33 $Y2=1.48
r60 23 28 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.83 $Y=1.48
+ $X2=12.665 $Y2=1.48
r61 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=12.83 $Y=1.48
+ $X2=13.33 $Y2=1.48
r62 19 28 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.665 $Y=1.645
+ $X2=12.665 $Y2=1.48
r63 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.665 $Y=1.645
+ $X2=12.665 $Y2=1.98
r64 15 28 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.665 $Y=1.315
+ $X2=12.665 $Y2=1.48
r65 15 17 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=12.665 $Y=1.315
+ $X2=12.665 $Y2=0.495
r66 13 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=13.425 $Y=2.465
+ $X2=13.425 $Y2=1.645
r67 9 30 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=13.425 $Y=0.705
+ $X2=13.425 $Y2=1.315
r68 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=12.52
+ $Y=1.835 $X2=12.665 $Y2=1.98
r69 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.52
+ $Y=0.285 $X2=12.665 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%VPWR 1 2 3 4 15 19 21 25 29 31 36 44 54
+ 55 58 61 64 71 82
r140 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r141 67 68 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 64 67 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=5.66 $Y=3.05
+ $X2=5.66 $Y2=3.33
r143 62 68 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=5.52 $Y2=3.33
r144 61 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r145 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r146 55 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r147 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r148 52 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.295 $Y=3.33
+ $X2=13.17 $Y2=3.33
r149 52 54 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.295 $Y=3.33
+ $X2=13.68 $Y2=3.33
r150 51 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r151 50 51 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r152 48 82 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.72
+ $Y2=3.33
r153 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r154 47 50 438.417 $w=1.68e-07 $l=6.72e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=12.72 $Y2=3.33
r155 47 48 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r156 45 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=3.33
+ $X2=5.66 $Y2=3.33
r157 45 47 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.825 $Y=3.33
+ $X2=6 $Y2=3.33
r158 44 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=13.17 $Y2=3.33
r159 44 50 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=12.72 $Y2=3.33
r160 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r161 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r162 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r163 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r164 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r165 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r166 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r167 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 36 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.525 $Y2=3.33
r169 36 42 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r170 34 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r171 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r172 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r173 31 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r174 29 51 1.60551 $w=4.9e-07 $l=5.76e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=12.72 $Y2=3.33
r175 29 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.72 $Y2=3.33
r176 25 28 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=13.17 $Y=1.98
+ $X2=13.17 $Y2=2.465
r177 23 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=3.33
r178 23 28 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=2.465
r179 22 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.65 $Y=3.33
+ $X2=2.525 $Y2=3.33
r180 21 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=3.33
+ $X2=5.66 $Y2=3.33
r181 21 22 185.61 $w=1.68e-07 $l=2.845e-06 $layer=LI1_cond $X=5.495 $Y=3.33
+ $X2=2.65 $Y2=3.33
r182 17 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=3.33
r183 17 19 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=2.85
r184 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r185 13 15 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.53
r186 4 28 300 $w=1.7e-07 $l=7.46693e-07 $layer=licon1_PDIFF $count=2 $X=12.955
+ $Y=1.835 $X2=13.21 $Y2=2.465
r187 4 25 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=12.955
+ $Y=1.835 $X2=13.21 $Y2=1.98
r188 3 64 600 $w=1.7e-07 $l=4.97996e-07 $layer=licon1_PDIFF $count=1 $X=5.44
+ $Y=2.65 $X2=5.66 $Y2=3.05
r189 2 19 600 $w=1.7e-07 $l=5.78619e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=2.385 $X2=2.565 $Y2=2.85
r190 1 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=2.385 $X2=0.73 $Y2=2.53
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%A_282_477# 1 2 3 4 15 17 18 19 22 23 24
+ 26 28 29 30 32 33 34 38 40 46 49
c159 40 0 1.10134e-19 $X=1.69 $Y=0.46
c160 23 0 1.4124e-19 $X=2.485 $Y=0.925
r161 49 51 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.64 $Y=0.945
+ $X2=3.64 $Y2=1.135
r162 45 46 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.745 $Y=2.405
+ $X2=2.905 $Y2=2.405
r163 40 42 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.69 $Y=0.46
+ $X2=1.69 $Y2=0.585
r164 36 38 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=4.26 $Y=2.905
+ $X2=4.26 $Y2=2.85
r165 35 38 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=4.26 $Y=2.235
+ $X2=4.26 $Y2=2.85
r166 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.095 $Y=2.15
+ $X2=4.26 $Y2=2.235
r167 33 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.095 $Y=2.15
+ $X2=3.805 $Y2=2.15
r168 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.72 $Y=2.065
+ $X2=3.805 $Y2=2.15
r169 32 51 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.72 $Y=2.065
+ $X2=3.72 $Y2=1.135
r170 29 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.095 $Y=2.99
+ $X2=4.26 $Y2=2.905
r171 29 30 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=4.095 $Y=2.99
+ $X2=2.99 $Y2=2.99
r172 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=2.905
+ $X2=2.99 $Y2=2.99
r173 27 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=2.49
+ $X2=2.905 $Y2=2.405
r174 27 28 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.905 $Y=2.49
+ $X2=2.905 $Y2=2.905
r175 26 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=2.32
+ $X2=2.745 $Y2=2.405
r176 25 44 3.06467 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.745 $Y=1.18
+ $X2=2.745 $Y2=1.01
r177 25 26 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.745 $Y=1.18
+ $X2=2.745 $Y2=2.32
r178 23 44 13.8554 $w=2.53e-07 $l=2.995e-07 $layer=LI1_cond $X=2.485 $Y=0.925
+ $X2=2.745 $Y2=1.01
r179 23 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.485 $Y=0.925
+ $X2=2.305 $Y2=0.925
r180 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=0.84
+ $X2=2.305 $Y2=0.925
r181 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.22 $Y=0.67
+ $X2=2.22 $Y2=0.84
r182 20 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0.585
+ $X2=1.69 $Y2=0.585
r183 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=0.585
+ $X2=2.22 $Y2=0.67
r184 19 20 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.135 $Y=0.585
+ $X2=1.855 $Y2=0.585
r185 17 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.405
+ $X2=2.745 $Y2=2.405
r186 17 18 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.66 $Y=2.405
+ $X2=1.715 $Y2=2.405
r187 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.55 $Y=2.49
+ $X2=1.715 $Y2=2.405
r188 13 15 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=1.55 $Y=2.49 $X2=1.55
+ $Y2=2.53
r189 4 38 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=2.65 $X2=4.26 $Y2=2.85
r190 3 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.385 $X2=1.55 $Y2=2.53
r191 2 49 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=3.495
+ $Y=0.695 $X2=3.64 $Y2=0.945
r192 1 40 182 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.69 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%KAPWR 1 2 7 10 16 17 22
r119 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.82
+ $X2=11.28 $Y2=2.82
r120 11 17 0.787035 $w=2.7e-07 $l=1.44e-06 $layer=MET1_cond $X=9.84 $Y=2.81
+ $X2=11.28 $Y2=2.81
r121 10 11 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=2.82
+ $X2=9.84 $Y2=2.82
r122 7 11 1.57407 $w=2.7e-07 $l=2.88e-06 $layer=MET1_cond $X=6.96 $Y=2.81
+ $X2=9.84 $Y2=2.81
r123 7 22 0.131172 $w=2.7e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=2.81
+ $X2=6.72 $Y2=2.81
r124 2 16 600 $w=1.7e-07 $l=8.98499e-07 $layer=licon1_PDIFF $count=1 $X=11.025
+ $Y=2.095 $X2=11.28 $Y2=2.875
r125 1 10 600 $w=1.7e-07 $l=8.47113e-07 $layer=licon1_PDIFF $count=1 $X=9.78
+ $Y=2.095 $X2=9.92 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%Q 1 2 9 14 15 16 17 23 29
r22 21 29 1.28049 $w=3.58e-07 $l=4e-08 $layer=LI1_cond $X=13.655 $Y=0.965
+ $X2=13.655 $Y2=0.925
r23 17 31 8.28694 $w=3.58e-07 $l=1.58e-07 $layer=LI1_cond $X=13.655 $Y=0.987
+ $X2=13.655 $Y2=1.145
r24 17 21 0.704271 $w=3.58e-07 $l=2.2e-08 $layer=LI1_cond $X=13.655 $Y=0.987
+ $X2=13.655 $Y2=0.965
r25 17 29 0.736283 $w=3.58e-07 $l=2.3e-08 $layer=LI1_cond $X=13.655 $Y=0.902
+ $X2=13.655 $Y2=0.925
r26 16 17 11.1083 $w=3.58e-07 $l=3.47e-07 $layer=LI1_cond $X=13.655 $Y=0.555
+ $X2=13.655 $Y2=0.902
r27 16 23 4.00154 $w=3.58e-07 $l=1.25e-07 $layer=LI1_cond $X=13.655 $Y=0.555
+ $X2=13.655 $Y2=0.43
r28 15 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.75 $Y=1.815
+ $X2=13.75 $Y2=1.145
r29 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=13.655 $Y=1.98
+ $X2=13.655 $Y2=1.815
r30 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=13.655 $Y=1.995
+ $X2=13.655 $Y2=1.98
r31 7 9 29.2913 $w=3.58e-07 $l=9.15e-07 $layer=LI1_cond $X=13.655 $Y=1.995
+ $X2=13.655 $Y2=2.91
r32 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.835 $X2=13.64 $Y2=1.98
r33 2 9 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.835 $X2=13.64 $Y2=2.91
r34 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.5
+ $Y=0.285 $X2=13.64 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFXTP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 46 47
+ 49 50 51 53 58 66 81 87 88 91 94 97 100 111
c154 29 0 5.25296e-20 $X=4.97 $Y=0.28
r155 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r156 98 111 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.72 $Y2=0
r157 97 98 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r158 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r159 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r160 88 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r161 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r162 85 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.295 $Y=0
+ $X2=13.17 $Y2=0
r163 85 87 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.295 $Y=0
+ $X2=13.68 $Y2=0
r164 84 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r165 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r166 81 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.045 $Y=0
+ $X2=13.17 $Y2=0
r167 81 83 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.045 $Y=0
+ $X2=12.72 $Y2=0
r168 80 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r169 79 80 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r170 77 80 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=11.76 $Y2=0
r171 76 79 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=11.76
+ $Y2=0
r172 76 77 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r173 74 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r174 73 74 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r175 71 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.055 $Y=0 $X2=4.93
+ $Y2=0
r176 71 73 186.914 $w=1.68e-07 $l=2.865e-06 $layer=LI1_cond $X=5.055 $Y=0
+ $X2=7.92 $Y2=0
r177 70 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r178 70 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=2.64 $Y2=0
r179 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r180 67 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.56
+ $Y2=0
r181 67 69 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=2.645 $Y=0
+ $X2=4.56 $Y2=0
r182 66 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.93
+ $Y2=0
r183 66 69 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.56
+ $Y2=0
r184 65 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r185 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r186 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r187 62 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r188 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r189 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r190 59 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.76
+ $Y2=0
r191 59 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.2
+ $Y2=0
r192 58 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.56
+ $Y2=0
r193 58 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.16 $Y2=0
r194 56 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r195 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r196 53 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.76
+ $Y2=0
r197 53 55 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.24 $Y2=0
r198 51 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r199 51 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.72 $Y2=0
r200 49 79 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=11.76 $Y2=0
r201 49 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=12.145 $Y2=0
r202 48 83 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=12.27 $Y=0
+ $X2=12.72 $Y2=0
r203 48 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.27 $Y=0
+ $X2=12.145 $Y2=0
r204 46 73 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=7.95 $Y=0 $X2=7.92
+ $Y2=0
r205 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.95 $Y=0 $X2=8.115
+ $Y2=0
r206 45 76 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.28 $Y=0 $X2=8.4
+ $Y2=0
r207 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=0 $X2=8.115
+ $Y2=0
r208 41 43 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=13.17 $Y=0.43
+ $X2=13.17 $Y2=0.98
r209 39 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.17 $Y2=0
r210 39 41 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.17 $Y2=0.43
r211 35 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.145 $Y=0.085
+ $X2=12.145 $Y2=0
r212 35 37 46.7892 $w=2.48e-07 $l=1.015e-06 $layer=LI1_cond $X=12.145 $Y=0.085
+ $X2=12.145 $Y2=1.1
r213 31 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0
r214 31 33 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0.73
r215 27 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0
r216 27 29 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0.28
r217 23 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r218 23 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.44
r219 19 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0
r220 19 21 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.44
r221 6 43 182 $w=1.7e-07 $l=8.12558e-07 $layer=licon1_NDIFF $count=1 $X=12.955
+ $Y=0.285 $X2=13.21 $Y2=0.98
r222 6 41 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=12.955
+ $Y=0.285 $X2=13.21 $Y2=0.43
r223 5 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.965
+ $Y=0.89 $X2=12.105 $Y2=1.1
r224 4 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.565 $X2=8.115 $Y2=0.73
r225 3 29 182 $w=1.7e-07 $l=5.13347e-07 $layer=licon1_NDIFF $count=1 $X=4.75
+ $Y=0.695 $X2=4.97 $Y2=0.28
r226 2 25 182 $w=1.7e-07 $l=2.84561e-07 $layer=licon1_NDIFF $count=1 $X=2.37
+ $Y=0.235 $X2=2.56 $Y2=0.44
r227 1 21 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.235 $X2=0.76 $Y2=0.44
.ends

