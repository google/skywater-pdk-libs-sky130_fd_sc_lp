# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o2bb2a_0
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o2bb2a_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 1.550000 1.295000 2.130000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.860000 1.350000 1.015000 ;
        RECT 1.000000 1.015000 1.610000 1.380000 ;
        RECT 1.105000 0.395000 1.350000 0.860000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.200000 1.155000 3.755000 2.215000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 1.155000 2.990000 1.825000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.380000 0.505000 0.710000 ;
        RECT 0.095000 0.710000 0.325000 2.395000 ;
        RECT 0.095000 2.395000 0.355000 3.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.495000  0.880000 0.715000 1.550000 ;
      RECT 0.525000  2.640000 0.835000 3.245000 ;
      RECT 0.545000  1.550000 0.715000 2.300000 ;
      RECT 0.545000  2.300000 1.175000 2.470000 ;
      RECT 0.675000  0.085000 0.935000 0.690000 ;
      RECT 1.005000  2.470000 1.175000 2.905000 ;
      RECT 1.005000  2.905000 1.975000 3.075000 ;
      RECT 1.345000  2.405000 1.635000 2.735000 ;
      RECT 1.465000  1.745000 2.035000 1.915000 ;
      RECT 1.465000  1.915000 1.635000 2.405000 ;
      RECT 1.520000  0.395000 1.960000 0.725000 ;
      RECT 1.790000  0.725000 1.960000 1.585000 ;
      RECT 1.790000  1.585000 2.035000 1.745000 ;
      RECT 1.805000  2.175000 2.865000 2.345000 ;
      RECT 1.805000  2.345000 1.975000 2.905000 ;
      RECT 2.130000  0.280000 2.375000 0.675000 ;
      RECT 2.145000  2.515000 2.405000 3.245000 ;
      RECT 2.205000  0.675000 2.375000 2.175000 ;
      RECT 2.545000  0.280000 2.830000 0.780000 ;
      RECT 2.545000  0.780000 3.725000 0.950000 ;
      RECT 2.575000  2.345000 2.865000 2.790000 ;
      RECT 3.000000  0.085000 3.260000 0.610000 ;
      RECT 3.325000  2.460000 3.655000 3.245000 ;
      RECT 3.430000  0.280000 3.725000 0.780000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__o2bb2a_0
