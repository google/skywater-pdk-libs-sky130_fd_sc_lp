* NGSPICE file created from sky130_fd_sc_lp__buflp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__buflp_2 A VGND VNB VPB VPWR X
M1000 a_128_367# a_98_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=3.528e+11p ps=3.08e+06u
M1001 a_128_367# a_98_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=9.65e+11p ps=6.68e+06u
M1002 a_509_377# A VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1003 VGND a_98_21# a_128_47# VNB nshort w=840000u l=150000u
+  ad=5.544e+11p pd=4.79e+06u as=5.292e+11p ps=4.62e+06u
M1004 X a_98_21# a_128_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_128_47# a_98_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.94e+11p ps=2.38e+06u
M1006 X a_98_21# a_128_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_128_47# a_98_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_516_47# A VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 VPWR a_98_21# a_128_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_98_21# A a_516_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1011 a_98_21# A a_509_377# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
.ends

