* File: sky130_fd_sc_lp__o32a_2.pxi.spice
* Created: Wed Sep  2 10:26:05 2020
* 
x_PM_SKY130_FD_SC_LP__O32A_2%A_85_21# N_A_85_21#_M1009_d N_A_85_21#_M1005_d
+ N_A_85_21#_M1011_g N_A_85_21#_M1006_g N_A_85_21#_M1013_g N_A_85_21#_M1012_g
+ N_A_85_21#_c_70_n N_A_85_21#_c_122_p N_A_85_21#_c_71_n N_A_85_21#_c_65_n
+ N_A_85_21#_c_66_n N_A_85_21#_c_67_n N_A_85_21#_c_75_n N_A_85_21#_c_101_p
+ PM_SKY130_FD_SC_LP__O32A_2%A_85_21#
x_PM_SKY130_FD_SC_LP__O32A_2%A1 N_A1_M1001_g N_A1_M1000_g A1 N_A1_c_155_n
+ N_A1_c_156_n PM_SKY130_FD_SC_LP__O32A_2%A1
x_PM_SKY130_FD_SC_LP__O32A_2%A2 N_A2_M1004_g N_A2_M1008_g A2 N_A2_c_188_n
+ N_A2_c_189_n PM_SKY130_FD_SC_LP__O32A_2%A2
x_PM_SKY130_FD_SC_LP__O32A_2%A3 N_A3_M1005_g N_A3_M1003_g A3 N_A3_c_221_n
+ N_A3_c_222_n PM_SKY130_FD_SC_LP__O32A_2%A3
x_PM_SKY130_FD_SC_LP__O32A_2%B2 N_B2_M1010_g N_B2_M1009_g B2 N_B2_c_254_n
+ N_B2_c_255_n PM_SKY130_FD_SC_LP__O32A_2%B2
x_PM_SKY130_FD_SC_LP__O32A_2%B1 N_B1_M1007_g N_B1_M1002_g B1 B1 N_B1_c_288_n
+ PM_SKY130_FD_SC_LP__O32A_2%B1
x_PM_SKY130_FD_SC_LP__O32A_2%VPWR N_VPWR_M1006_s N_VPWR_M1012_s N_VPWR_M1002_d
+ N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n
+ VPWR N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_313_n
+ PM_SKY130_FD_SC_LP__O32A_2%VPWR
x_PM_SKY130_FD_SC_LP__O32A_2%X N_X_M1011_s N_X_M1006_d X X X X X X X N_X_c_360_n
+ PM_SKY130_FD_SC_LP__O32A_2%X
x_PM_SKY130_FD_SC_LP__O32A_2%VGND N_VGND_M1011_d N_VGND_M1013_d N_VGND_M1004_d
+ N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n
+ N_VGND_c_387_n VGND N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n
+ N_VGND_c_391_n PM_SKY130_FD_SC_LP__O32A_2%VGND
x_PM_SKY130_FD_SC_LP__O32A_2%A_341_47# N_A_341_47#_M1001_d N_A_341_47#_M1003_d
+ N_A_341_47#_M1007_d N_A_341_47#_c_445_n N_A_341_47#_c_438_n
+ N_A_341_47#_c_440_n N_A_341_47#_c_460_n N_A_341_47#_c_455_n
+ N_A_341_47#_c_441_n N_A_341_47#_c_437_n PM_SKY130_FD_SC_LP__O32A_2%A_341_47#
cc_1 VNB N_A_85_21#_M1011_g 0.0340797f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_2 VNB N_A_85_21#_M1013_g 0.0273582f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.655
cc_3 VNB N_A_85_21#_c_65_n 0.00442802f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.71
cc_4 VNB N_A_85_21#_c_66_n 0.00934122f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.505
cc_5 VNB N_A_85_21#_c_67_n 0.0581007f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.505
cc_6 VNB N_A1_M1000_g 0.00764859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB A1 0.00282816f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_8 VNB N_A1_c_155_n 0.0336336f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.67
cc_9 VNB N_A1_c_156_n 0.0187198f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_10 VNB N_A2_M1008_g 0.00769607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A2 0.00165801f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_12 VNB N_A2_c_188_n 0.0318779f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.67
cc_13 VNB N_A2_c_189_n 0.0188377f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_14 VNB N_A3_M1005_g 0.00862586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A3 0.00422874f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_16 VNB N_A3_c_221_n 0.0303065f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.67
cc_17 VNB N_A3_c_222_n 0.0188359f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_18 VNB N_B2_M1010_g 0.00703781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B2_M1009_g 0.0183962f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.34
cc_20 VNB N_B2_c_254_n 0.0302149f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_21 VNB N_B2_c_255_n 0.00286815f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_22 VNB N_B1_M1007_g 0.0239843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_M1002_g 0.00623472f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.34
cc_24 VNB B1 0.0255496f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_25 VNB N_B1_c_288_n 0.052134f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.655
cc_26 VNB N_VPWR_c_313_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_360_n 0.00558985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_382_n 0.0117031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_383_n 0.0500107f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_30 VNB N_VGND_c_384_n 0.00564356f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.655
cc_31 VNB N_VGND_c_385_n 0.00564356f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.465
cc_32 VNB N_VGND_c_386_n 0.0223974f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=1.77
cc_33 VNB N_VGND_c_387_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.77
cc_34 VNB N_VGND_c_388_n 0.0199547f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=1.98
cc_35 VNB N_VGND_c_389_n 0.0452315f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=0.765
cc_36 VNB N_VGND_c_390_n 0.234247f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=0.76
cc_37 VNB N_VGND_c_391_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.505
cc_38 VNB N_A_341_47#_c_437_n 0.0309037f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=1.925
cc_39 VPB N_A_85_21#_M1006_g 0.0259352f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_40 VPB N_A_85_21#_M1012_g 0.0217193f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.465
cc_41 VPB N_A_85_21#_c_70_n 0.0110285f $X=-0.19 $Y=1.655 $X2=2.7 $Y2=1.77
cc_42 VPB N_A_85_21#_c_71_n 0.00498297f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=1.817
cc_43 VPB N_A_85_21#_c_65_n 5.20539e-19 $X=-0.19 $Y=1.655 $X2=3.57 $Y2=1.71
cc_44 VPB N_A_85_21#_c_66_n 0.00376516f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.505
cc_45 VPB N_A_85_21#_c_67_n 0.0118111f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.505
cc_46 VPB N_A_85_21#_c_75_n 0.00429353f $X=-0.19 $Y=1.655 $X2=2.7 $Y2=1.685
cc_47 VPB N_A1_M1000_g 0.0203074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_M1008_g 0.0190166f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A3_M1005_g 0.0211934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B2_M1010_g 0.0213343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B1_M1002_g 0.0238087f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.34
cc_52 VPB B1 0.01834f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_53 VPB N_VPWR_c_314_n 0.0116772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_315_n 0.0656653f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_55 VPB N_VPWR_c_316_n 0.00183948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_317_n 0.0152774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_318_n 0.0462519f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.77
cc_58 VPB N_VPWR_c_319_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_320_n 0.0645394f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.505
cc_60 VPB N_VPWR_c_321_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.505
cc_61 VPB N_VPWR_c_313_n 0.0516072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_X_c_360_n 0.00270097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 N_A_85_21#_M1012_g N_A1_M1000_g 0.00600671f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_85_21#_c_70_n N_A1_M1000_g 0.0148545f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_65 N_A_85_21#_c_66_n N_A1_M1000_g 0.00371886f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_66 N_A_85_21#_c_67_n N_A1_M1000_g 0.00408309f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_67 N_A_85_21#_M1013_g A1 7.48754e-19 $X=0.93 $Y=0.655 $X2=0 $Y2=0
cc_68 N_A_85_21#_c_70_n A1 0.021399f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_69 N_A_85_21#_c_66_n A1 0.013283f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_70 N_A_85_21#_M1013_g N_A1_c_155_n 0.00393308f $X=0.93 $Y=0.655 $X2=0 $Y2=0
cc_71 N_A_85_21#_c_70_n N_A1_c_155_n 0.00552315f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_72 N_A_85_21#_c_66_n N_A1_c_155_n 0.00117835f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_73 N_A_85_21#_c_67_n N_A1_c_155_n 0.0108874f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_74 N_A_85_21#_M1013_g N_A1_c_156_n 0.017018f $X=0.93 $Y=0.655 $X2=0 $Y2=0
cc_75 N_A_85_21#_c_70_n N_A2_M1008_g 0.0150723f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_76 N_A_85_21#_c_70_n A2 0.0240681f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_77 N_A_85_21#_c_70_n N_A2_c_188_n 0.00126186f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_78 N_A_85_21#_c_70_n N_A3_M1005_g 0.01568f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_79 N_A_85_21#_c_70_n A3 0.015627f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_80 N_A_85_21#_c_75_n A3 0.0129811f $X=2.7 $Y=1.685 $X2=0 $Y2=0
cc_81 N_A_85_21#_c_75_n N_A3_c_221_n 0.00120479f $X=2.7 $Y=1.685 $X2=0 $Y2=0
cc_82 N_A_85_21#_c_71_n N_B2_M1010_g 0.0181523f $X=3.485 $Y=1.817 $X2=0 $Y2=0
cc_83 N_A_85_21#_c_65_n N_B2_M1010_g 0.00300977f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_84 N_A_85_21#_c_75_n N_B2_M1010_g 3.43482e-19 $X=2.7 $Y=1.685 $X2=0 $Y2=0
cc_85 N_A_85_21#_c_65_n N_B2_M1009_g 0.00417507f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_86 N_A_85_21#_c_71_n N_B2_c_254_n 0.00561253f $X=3.485 $Y=1.817 $X2=0 $Y2=0
cc_87 N_A_85_21#_c_65_n N_B2_c_254_n 0.00206348f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_88 N_A_85_21#_c_101_p N_B2_c_254_n 0.00268045f $X=3.57 $Y=0.765 $X2=0 $Y2=0
cc_89 N_A_85_21#_c_71_n N_B2_c_255_n 0.0213351f $X=3.485 $Y=1.817 $X2=0 $Y2=0
cc_90 N_A_85_21#_c_65_n N_B2_c_255_n 0.0245294f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_91 N_A_85_21#_c_75_n N_B2_c_255_n 4.42308e-19 $X=2.7 $Y=1.685 $X2=0 $Y2=0
cc_92 N_A_85_21#_c_65_n N_B1_M1007_g 0.0105325f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_93 N_A_85_21#_c_101_p N_B1_M1007_g 0.00501979f $X=3.57 $Y=0.765 $X2=0 $Y2=0
cc_94 N_A_85_21#_c_71_n N_B1_M1002_g 0.012009f $X=3.485 $Y=1.817 $X2=0 $Y2=0
cc_95 N_A_85_21#_c_65_n N_B1_M1002_g 0.00367676f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_96 N_A_85_21#_c_71_n B1 0.00937373f $X=3.485 $Y=1.817 $X2=0 $Y2=0
cc_97 N_A_85_21#_c_65_n B1 0.0337659f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_98 N_A_85_21#_c_65_n N_B1_c_288_n 0.00790423f $X=3.57 $Y=1.71 $X2=0 $Y2=0
cc_99 N_A_85_21#_c_70_n N_VPWR_M1012_s 0.00240673f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_100 N_A_85_21#_c_66_n N_VPWR_M1012_s 0.00214979f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_101 N_A_85_21#_M1006_g N_VPWR_c_315_n 0.00768196f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_85_21#_M1006_g N_VPWR_c_316_n 7.73831e-19 $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_85_21#_M1012_g N_VPWR_c_316_n 0.0172577f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_85_21#_c_70_n N_VPWR_c_316_n 0.0198926f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_105 N_A_85_21#_c_66_n N_VPWR_c_316_n 0.0223825f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_106 N_A_85_21#_c_67_n N_VPWR_c_316_n 0.00129349f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_107 N_A_85_21#_M1006_g N_VPWR_c_319_n 0.00585385f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_85_21#_M1012_g N_VPWR_c_319_n 0.00486043f $X=0.93 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_A_85_21#_c_122_p N_VPWR_c_320_n 0.0212513f $X=2.865 $Y=1.98 $X2=0 $Y2=0
cc_110 N_A_85_21#_M1005_d N_VPWR_c_313_n 0.00526034f $X=2.675 $Y=1.835 $X2=0
+ $Y2=0
cc_111 N_A_85_21#_M1006_g N_VPWR_c_313_n 0.0114778f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_85_21#_M1012_g N_VPWR_c_313_n 0.00824727f $X=0.93 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_85_21#_c_122_p N_VPWR_c_313_n 0.0127519f $X=2.865 $Y=1.98 $X2=0 $Y2=0
cc_114 N_A_85_21#_M1011_g N_X_c_360_n 0.00733087f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_115 N_A_85_21#_M1006_g N_X_c_360_n 0.00454772f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_85_21#_M1013_g N_X_c_360_n 0.00724702f $X=0.93 $Y=0.655 $X2=0 $Y2=0
cc_117 N_A_85_21#_M1012_g N_X_c_360_n 0.00217088f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_85_21#_c_66_n N_X_c_360_n 0.0325242f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_119 N_A_85_21#_c_67_n N_X_c_360_n 0.029544f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_120 N_A_85_21#_c_70_n A_355_367# 0.00366293f $X=2.7 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_85_21#_c_70_n A_427_367# 0.0105625f $X=2.7 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_85_21#_c_71_n A_643_367# 0.0113119f $X=3.485 $Y=1.817 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_85_21#_M1011_g N_VGND_c_383_n 0.00839485f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_124 N_A_85_21#_M1013_g N_VGND_c_384_n 0.0124106f $X=0.93 $Y=0.655 $X2=0 $Y2=0
cc_125 N_A_85_21#_c_70_n N_VGND_c_384_n 0.00291049f $X=2.7 $Y=1.77 $X2=0 $Y2=0
cc_126 N_A_85_21#_c_66_n N_VGND_c_384_n 0.0131526f $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_127 N_A_85_21#_c_67_n N_VGND_c_384_n 9.13184e-19 $X=1.07 $Y=1.505 $X2=0 $Y2=0
cc_128 N_A_85_21#_M1011_g N_VGND_c_388_n 0.00585385f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_129 N_A_85_21#_M1013_g N_VGND_c_388_n 0.00585385f $X=0.93 $Y=0.655 $X2=0
+ $Y2=0
cc_130 N_A_85_21#_M1009_d N_VGND_c_390_n 0.00257355f $X=3.285 $Y=0.235 $X2=0
+ $Y2=0
cc_131 N_A_85_21#_M1011_g N_VGND_c_390_n 0.0114778f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_132 N_A_85_21#_M1013_g N_VGND_c_390_n 0.0114584f $X=0.93 $Y=0.655 $X2=0 $Y2=0
cc_133 N_A_85_21#_c_70_n N_A_341_47#_c_438_n 0.00484983f $X=2.7 $Y=1.77 $X2=0
+ $Y2=0
cc_134 N_A_85_21#_c_75_n N_A_341_47#_c_438_n 0.00488917f $X=2.7 $Y=1.685 $X2=0
+ $Y2=0
cc_135 N_A_85_21#_c_70_n N_A_341_47#_c_440_n 0.00430921f $X=2.7 $Y=1.77 $X2=0
+ $Y2=0
cc_136 N_A_85_21#_M1009_d N_A_341_47#_c_441_n 0.00412961f $X=3.285 $Y=0.235
+ $X2=0 $Y2=0
cc_137 N_A_85_21#_c_101_p N_A_341_47#_c_441_n 0.0181244f $X=3.57 $Y=0.765 $X2=0
+ $Y2=0
cc_138 N_A_85_21#_c_65_n N_A_341_47#_c_437_n 0.0076449f $X=3.57 $Y=1.71 $X2=0
+ $Y2=0
cc_139 N_A_85_21#_c_101_p N_A_341_47#_c_437_n 0.0261095f $X=3.57 $Y=0.765 $X2=0
+ $Y2=0
cc_140 N_A1_M1000_g N_A2_M1008_g 0.0641255f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_141 A1 A2 0.0239324f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A1_c_155_n A2 3.49821e-19 $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_143 A1 N_A2_c_188_n 0.00223666f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A1_c_155_n N_A2_c_188_n 0.0641255f $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_145 N_A1_c_156_n N_A2_c_189_n 0.0152593f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_146 N_A1_M1000_g N_VPWR_c_316_n 0.027214f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A1_M1000_g N_VPWR_c_320_n 0.00486043f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A1_M1000_g N_VPWR_c_313_n 0.00818711f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A1_c_156_n N_VGND_c_384_n 0.0115657f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_150 N_A1_c_156_n N_VGND_c_386_n 0.0054895f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_151 N_A1_c_156_n N_VGND_c_390_n 0.0106313f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A1_c_156_n N_A_341_47#_c_445_n 0.00843533f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_153 A1 N_A_341_47#_c_440_n 0.00864361f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A1_c_155_n N_A_341_47#_c_440_n 0.0017331f $X=1.61 $Y=1.35 $X2=0 $Y2=0
cc_155 N_A1_c_156_n N_A_341_47#_c_440_n 0.00211924f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_156 N_A2_M1008_g N_A3_M1005_g 0.0565612f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_157 A2 A3 0.024359f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A2_c_188_n A3 0.00173939f $X=2.15 $Y=1.35 $X2=0 $Y2=0
cc_159 A2 N_A3_c_221_n 3.51842e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_c_188_n N_A3_c_221_n 0.0209243f $X=2.15 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A2_c_189_n N_A3_c_222_n 0.0176445f $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A2_M1008_g N_VPWR_c_316_n 0.00650653f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A2_M1008_g N_VPWR_c_320_n 0.00585385f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A2_M1008_g N_VPWR_c_313_n 0.011101f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A2_c_189_n N_VGND_c_385_n 0.00810057f $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A2_c_189_n N_VGND_c_386_n 0.0054895f $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_167 N_A2_c_189_n N_VGND_c_390_n 0.0106628f $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_168 N_A2_c_189_n N_A_341_47#_c_445_n 0.0102095f $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_169 A2 N_A_341_47#_c_438_n 0.0200071f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A2_c_188_n N_A_341_47#_c_438_n 0.00402783f $X=2.15 $Y=1.35 $X2=0 $Y2=0
cc_171 N_A2_c_189_n N_A_341_47#_c_438_n 0.0123033f $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_172 A2 N_A_341_47#_c_440_n 0.00191494f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A2_c_189_n N_A_341_47#_c_440_n 7.3104e-19 $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_174 N_A2_c_189_n N_A_341_47#_c_455_n 7.6739e-19 $X=2.15 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A3_c_222_n N_B2_M1009_g 0.0158135f $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_176 N_A3_M1005_g N_B2_c_254_n 0.0303079f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_177 A3 N_B2_c_254_n 3.49366e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A3_c_221_n N_B2_c_254_n 0.0190731f $X=2.69 $Y=1.35 $X2=0 $Y2=0
cc_179 N_A3_M1005_g N_B2_c_255_n 4.63436e-19 $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_180 A3 N_B2_c_255_n 0.0241348f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A3_c_221_n N_B2_c_255_n 0.00169076f $X=2.69 $Y=1.35 $X2=0 $Y2=0
cc_182 N_A3_M1005_g N_VPWR_c_320_n 0.00585385f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A3_M1005_g N_VPWR_c_313_n 0.0114286f $X=2.6 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A3_c_222_n N_VGND_c_385_n 0.00800696f $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_185 N_A3_c_222_n N_VGND_c_389_n 0.00547432f $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_186 N_A3_c_222_n N_VGND_c_390_n 0.0106257f $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_187 N_A3_c_222_n N_A_341_47#_c_445_n 7.98124e-19 $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_188 A3 N_A_341_47#_c_438_n 0.0250312f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A3_c_221_n N_A_341_47#_c_438_n 0.00463009f $X=2.69 $Y=1.35 $X2=0 $Y2=0
cc_190 N_A3_c_222_n N_A_341_47#_c_438_n 0.0130343f $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_191 N_A3_c_222_n N_A_341_47#_c_460_n 0.00232783f $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A3_c_222_n N_A_341_47#_c_455_n 0.00784611f $X=2.69 $Y=1.185 $X2=0 $Y2=0
cc_193 N_B2_M1009_g N_B1_M1007_g 0.0266175f $X=3.21 $Y=0.655 $X2=0 $Y2=0
cc_194 N_B2_M1010_g N_B1_M1002_g 0.0487307f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_195 N_B2_c_254_n N_B1_c_288_n 0.0204702f $X=3.23 $Y=1.375 $X2=0 $Y2=0
cc_196 N_B2_c_255_n N_B1_c_288_n 2.85575e-19 $X=3.23 $Y=1.375 $X2=0 $Y2=0
cc_197 N_B2_M1010_g N_VPWR_c_320_n 0.00585385f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_198 N_B2_M1010_g N_VPWR_c_313_n 0.011557f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_199 N_B2_M1009_g N_VGND_c_389_n 0.00357877f $X=3.21 $Y=0.655 $X2=0 $Y2=0
cc_200 N_B2_M1009_g N_VGND_c_390_n 0.00550473f $X=3.21 $Y=0.655 $X2=0 $Y2=0
cc_201 N_B2_c_254_n N_A_341_47#_c_438_n 0.00161214f $X=3.23 $Y=1.375 $X2=0 $Y2=0
cc_202 N_B2_c_255_n N_A_341_47#_c_438_n 0.00650161f $X=3.23 $Y=1.375 $X2=0 $Y2=0
cc_203 N_B2_M1009_g N_A_341_47#_c_441_n 0.0124156f $X=3.21 $Y=0.655 $X2=0 $Y2=0
cc_204 N_B1_M1002_g N_VPWR_c_318_n 0.00497867f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_205 B1 N_VPWR_c_318_n 0.0195123f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_206 N_B1_c_288_n N_VPWR_c_318_n 0.00202661f $X=3.93 $Y=1.375 $X2=0 $Y2=0
cc_207 N_B1_M1002_g N_VPWR_c_320_n 0.00585385f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B1_M1002_g N_VPWR_c_313_n 0.0120969f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B1_M1007_g N_VGND_c_389_n 0.00357877f $X=3.68 $Y=0.655 $X2=0 $Y2=0
cc_210 N_B1_M1007_g N_VGND_c_390_n 0.00653509f $X=3.68 $Y=0.655 $X2=0 $Y2=0
cc_211 N_B1_M1007_g N_A_341_47#_c_441_n 0.0108748f $X=3.68 $Y=0.655 $X2=0 $Y2=0
cc_212 N_B1_M1007_g N_A_341_47#_c_437_n 0.0062239f $X=3.68 $Y=0.655 $X2=0 $Y2=0
cc_213 B1 N_A_341_47#_c_437_n 0.021598f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_214 N_B1_c_288_n N_A_341_47#_c_437_n 0.00285168f $X=3.93 $Y=1.375 $X2=0 $Y2=0
cc_215 N_VPWR_c_313_n N_X_M1006_d 0.0041489f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_315_n N_X_c_360_n 0.0015231f $X=0.285 $Y=1.98 $X2=0 $Y2=0
cc_217 N_VPWR_c_319_n N_X_c_360_n 0.0136943f $X=0.98 $Y=3.33 $X2=0 $Y2=0
cc_218 N_VPWR_c_313_n N_X_c_360_n 0.00866972f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_c_313_n A_355_367# 0.00899413f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_220 N_VPWR_c_313_n A_427_367# 0.0167135f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_221 N_VPWR_c_313_n A_643_367# 0.0167135f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_222 N_X_c_360_n N_VGND_c_383_n 0.00112229f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_223 N_X_c_360_n N_VGND_c_388_n 0.0136943f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_224 N_X_M1011_s N_VGND_c_390_n 0.0041489f $X=0.575 $Y=0.235 $X2=0 $Y2=0
cc_225 N_X_c_360_n N_VGND_c_390_n 0.00866972f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_226 N_VGND_c_390_n N_A_341_47#_M1001_d 0.00223559f $X=4.08 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_227 N_VGND_c_390_n N_A_341_47#_M1003_d 0.00220342f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_390_n N_A_341_47#_M1007_d 0.00244485f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_384_n N_A_341_47#_c_445_n 0.036611f $X=1.275 $Y=0.38 $X2=0 $Y2=0
cc_230 N_VGND_c_385_n N_A_341_47#_c_445_n 0.0265115f $X=2.415 $Y=0.575 $X2=0
+ $Y2=0
cc_231 N_VGND_c_386_n N_A_341_47#_c_445_n 0.0189236f $X=2.25 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_390_n N_A_341_47#_c_445_n 0.0123859f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_M1004_d N_A_341_47#_c_438_n 0.0162002f $X=2.135 $Y=0.235 $X2=0
+ $Y2=0
cc_234 N_VGND_c_385_n N_A_341_47#_c_438_n 0.0266856f $X=2.415 $Y=0.575 $X2=0
+ $Y2=0
cc_235 N_VGND_c_384_n N_A_341_47#_c_440_n 0.00995147f $X=1.275 $Y=0.38 $X2=0
+ $Y2=0
cc_236 N_VGND_c_385_n N_A_341_47#_c_460_n 0.0103989f $X=2.415 $Y=0.575 $X2=0
+ $Y2=0
cc_237 N_VGND_c_389_n N_A_341_47#_c_460_n 0.0172109f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_390_n N_A_341_47#_c_460_n 0.0114757f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_385_n N_A_341_47#_c_455_n 0.0157434f $X=2.415 $Y=0.575 $X2=0
+ $Y2=0
cc_240 N_VGND_c_389_n N_A_341_47#_c_441_n 0.0384609f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_390_n N_A_341_47#_c_441_n 0.024616f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_242 N_VGND_c_389_n N_A_341_47#_c_437_n 0.0190394f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_390_n N_A_341_47#_c_437_n 0.010497f $X=4.08 $Y=0 $X2=0 $Y2=0
