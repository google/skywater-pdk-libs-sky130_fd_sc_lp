* File: sky130_fd_sc_lp__nor4_2.spice
* Created: Fri Aug 28 10:57:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4_2.pex.spice"
.subckt sky130_fd_sc_lp__nor4_2  VNB VPB B A C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_B_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75003.4 A=0.126
+ P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75003 A=0.126
+ P=1.98 MULT=1
MM1014 N_VGND_M1010_d N_A_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75002.5 A=0.126
+ P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.84 AD=0.1974
+ AS=0.1176 PD=1.31 PS=1.12 NRD=14.28 NRS=0 M=1 R=5.6 SA=75001.5 SB=75002.1
+ A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1004_d N_C_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84 AD=0.1974
+ AS=0.1176 PD=1.31 PS=1.12 NRD=12.852 NRS=0 M=1 R=5.6 SA=75002.1 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1011_s N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1013 N_Y_M1013_d N_D_M1013_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_C_M1012_g N_Y_M1013_d VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.4 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1007 N_A_157_367#_M1007_d N_B_M1007_g N_A_74_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_157_367#_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6 SB=75003
+ A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1000_d N_A_M1005_g N_A_157_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_157_367#_M1005_s N_B_M1015_g N_A_74_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3402 PD=1.54 PS=1.8 NRD=0 NRS=23.443 M=1 R=8.4
+ SA=75001.5 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1001 N_A_74_367#_M1015_s N_C_M1001_g N_A_553_367#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3402 AS=0.1764 PD=1.8 PS=1.54 NRD=17.1981 NRS=0 M=1 R=8.4
+ SA=75002.2 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_D_M1006_g N_A_553_367#_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1006_d N_D_M1008_g N_A_553_367#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1009 N_A_74_367#_M1009_d N_C_M1009_g N_A_553_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__nor4_2.pxi.spice"
*
.ends
*
*
