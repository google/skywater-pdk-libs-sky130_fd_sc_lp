* File: sky130_fd_sc_lp__o2111ai_m.spice
* Created: Fri Aug 28 11:01:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o2111ai_m  VNB VPB D1 C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 A_213_50# N_D1_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.168 PD=0.63 PS=1.64 NRD=14.28 NRS=38.568 M=1 R=2.8 SA=75000.3 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1004 A_285_50# N_C1_M1004_g A_213_50# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_357_50#_M1005_d N_B1_M1005_g A_285_50# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_357_50#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_357_50#_M1000_d N_A1_M1000_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_D1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.2226 PD=0.7 PS=1.9 NRD=0 NRS=124.287 M=1 R=2.8 SA=75000.5
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_C1_M1009_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.3 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1001 A_443_535# N_A2_M1001_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_443_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o2111ai_m.pxi.spice"
*
.ends
*
*
