* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1162_463# a_934_367# a_1349_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_759_119# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND a_759_119# a_934_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_1770_412# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND a_1770_412# a_2516_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Q_N a_1770_412# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_359_489# SCE a_486_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Q_N a_1770_412# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR RESET_B a_1923_174# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_759_119# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1879_68# a_1923_174# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_359_489# a_27_81# a_445_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_486_81# SCD a_240_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_359_489# a_759_119# a_1162_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1885_496# a_1923_174# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_240_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1770_412# a_759_119# a_1879_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_81# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_759_119# a_934_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND a_2516_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_1770_412# a_934_367# a_1885_496# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_1248_463# a_1290_365# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_1923_174# a_1770_412# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VPWR a_1162_463# a_1290_365# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X24 a_1290_365# a_759_119# a_1770_412# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 a_323_81# D a_359_489# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR a_1770_412# a_2516_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_2067_68# a_1770_412# a_1923_174# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR RESET_B a_1162_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_1162_463# a_759_119# a_1248_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_1290_365# a_934_367# a_1770_412# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X31 Q a_2516_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_359_489# a_934_367# a_1162_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 Q a_2516_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 a_1421_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VPWR a_2516_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 VPWR RESET_B a_359_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 VPWR a_1770_412# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 a_445_489# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 VGND CLK a_759_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_240_81# a_27_81# a_323_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_934_367# a_759_119# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_1349_119# a_1290_365# a_1421_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 VGND a_1162_463# a_1290_365# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X44 VPWR SCE a_287_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X45 a_287_489# D a_359_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X46 VGND RESET_B a_2067_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 a_27_81# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
