* NGSPICE file created from sky130_fd_sc_lp__and2_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and2_2 A B VGND VNB VPB VPWR X
M1000 VPWR B a_46_47# VPB phighvt w=420000u l=150000u
+  ad=8.253e+11p pd=7.69e+06u as=1.176e+11p ps=1.4e+06u
M1001 VPWR a_46_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1002 X a_46_47# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=4.914e+11p ps=4.64e+06u
M1003 a_129_47# A a_46_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1004 X a_46_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_46_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_46_47# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B a_129_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

