* File: sky130_fd_sc_lp__o2111ai_4.pex.spice
* Created: Wed Sep  2 10:13:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111AI_4%D1 3 7 11 15 19 23 27 31 38 42 43 47 56
r76 46 56 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.71 $Y=1.42
+ $X2=1.765 $Y2=1.42
r77 46 54 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.71 $Y=1.42
+ $X2=1.335 $Y2=1.42
r78 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.42 $X2=1.71 $Y2=1.42
r79 43 47 12.5824 $w=3.03e-07 $l=3.33e-07 $layer=LI1_cond $X=1.533 $Y=1.352
+ $X2=1.2 $Y2=1.352
r80 43 45 7.86506 $w=3.05e-07 $l=1.77e-07 $layer=LI1_cond $X=1.533 $Y=1.352
+ $X2=1.71 $Y2=1.352
r81 41 54 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.03 $Y=1.42
+ $X2=1.335 $Y2=1.42
r82 41 52 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.03 $Y=1.42
+ $X2=0.905 $Y2=1.42
r83 40 42 5.45178 $w=3.03e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=1.352
+ $X2=0.945 $Y2=1.352
r84 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.42 $X2=1.03 $Y2=1.42
r85 38 47 3.89186 $w=3.03e-07 $l=1.03e-07 $layer=LI1_cond $X=1.097 $Y=1.352
+ $X2=1.2 $Y2=1.352
r86 38 40 2.5316 $w=3.03e-07 $l=6.7e-08 $layer=LI1_cond $X=1.097 $Y=1.352
+ $X2=1.03 $Y2=1.352
r87 36 52 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.69 $Y=1.42
+ $X2=0.905 $Y2=1.42
r88 36 49 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.69 $Y=1.42
+ $X2=0.475 $Y2=1.42
r89 35 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.69 $Y=1.42
+ $X2=0.945 $Y2=1.42
r90 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.42 $X2=0.69 $Y2=1.42
r91 29 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.585
+ $X2=1.765 $Y2=1.42
r92 29 31 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.765 $Y=1.585
+ $X2=1.765 $Y2=2.465
r93 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.255
+ $X2=1.765 $Y2=1.42
r94 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.765 $Y=1.255
+ $X2=1.765 $Y2=0.655
r95 21 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.585
+ $X2=1.335 $Y2=1.42
r96 21 23 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.335 $Y=1.585
+ $X2=1.335 $Y2=2.465
r97 17 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.255
+ $X2=1.335 $Y2=1.42
r98 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.335 $Y=1.255
+ $X2=1.335 $Y2=0.655
r99 13 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.585
+ $X2=0.905 $Y2=1.42
r100 13 15 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.905 $Y=1.585
+ $X2=0.905 $Y2=2.465
r101 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.255
+ $X2=0.905 $Y2=1.42
r102 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.905 $Y=1.255
+ $X2=0.905 $Y2=0.655
r103 5 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.585
+ $X2=0.475 $Y2=1.42
r104 5 7 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.475 $Y=1.585
+ $X2=0.475 $Y2=2.465
r105 1 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.255
+ $X2=0.475 $Y2=1.42
r106 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.475 $Y=1.255 $X2=0.475
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%C1 3 7 11 15 19 23 27 31 41 45 46 57 58
c86 58 0 1.19089e-19 $X=3.61 $Y=1.42
r87 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.61
+ $Y=1.42 $X2=3.61 $Y2=1.42
r88 55 57 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.485 $Y=1.42
+ $X2=3.61 $Y2=1.42
r89 46 58 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=3.6 $Y=1.33 $X2=3.61
+ $Y2=1.33
r90 44 55 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.27 $Y=1.42
+ $X2=3.485 $Y2=1.42
r91 44 53 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.27 $Y=1.42
+ $X2=3.055 $Y2=1.42
r92 43 45 7.81367 $w=3.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.27 $Y=1.33
+ $X2=3.115 $Y2=1.33
r93 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.42 $X2=3.27 $Y2=1.42
r94 41 46 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=3.29 $Y=1.33 $X2=3.6
+ $Y2=1.33
r95 41 43 0.658539 $w=3.48e-07 $l=2e-08 $layer=LI1_cond $X=3.29 $Y=1.33 $X2=3.27
+ $Y2=1.33
r96 40 53 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.93 $Y=1.42
+ $X2=3.055 $Y2=1.42
r97 40 51 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.93 $Y=1.42
+ $X2=2.625 $Y2=1.42
r98 39 45 11.399 $w=1.78e-07 $l=1.85e-07 $layer=LI1_cond $X=2.93 $Y=1.415
+ $X2=3.115 $Y2=1.415
r99 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.93
+ $Y=1.42 $X2=2.93 $Y2=1.42
r100 36 51 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.25 $Y=1.42
+ $X2=2.625 $Y2=1.42
r101 36 48 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.25 $Y=1.42
+ $X2=2.195 $Y2=1.42
r102 35 39 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.25 $Y=1.415
+ $X2=2.93 $Y2=1.415
r103 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.42 $X2=2.25 $Y2=1.42
r104 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.585
+ $X2=3.485 $Y2=1.42
r105 29 31 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.485 $Y=1.585
+ $X2=3.485 $Y2=2.465
r106 25 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.255
+ $X2=3.485 $Y2=1.42
r107 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.485 $Y=1.255
+ $X2=3.485 $Y2=0.655
r108 21 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.585
+ $X2=3.055 $Y2=1.42
r109 21 23 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.055 $Y=1.585
+ $X2=3.055 $Y2=2.465
r110 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.255
+ $X2=3.055 $Y2=1.42
r111 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.055 $Y=1.255
+ $X2=3.055 $Y2=0.655
r112 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.585
+ $X2=2.625 $Y2=1.42
r113 13 15 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.625 $Y=1.585
+ $X2=2.625 $Y2=2.465
r114 9 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.255
+ $X2=2.625 $Y2=1.42
r115 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.625 $Y=1.255
+ $X2=2.625 $Y2=0.655
r116 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.585
+ $X2=2.195 $Y2=1.42
r117 5 7 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.195 $Y=1.585
+ $X2=2.195 $Y2=2.465
r118 1 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.255
+ $X2=2.195 $Y2=1.42
r119 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.195 $Y=1.255 $X2=2.195
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 45
c85 16 0 1.7599e-19 $X=5.295 $Y=1.185
c86 4 0 1.19089e-19 $X=4.435 $Y=1.185
r87 43 45 2.34436 $w=5.14e-07 $l=2.5e-08 $layer=POLY_cond $X=5.52 $Y=1.457
+ $X2=5.545 $Y2=1.457
r88 41 43 21.0992 $w=5.14e-07 $l=2.25e-07 $layer=POLY_cond $X=5.295 $Y=1.457
+ $X2=5.52 $Y2=1.457
r89 40 41 16.8794 $w=5.14e-07 $l=1.8e-07 $layer=POLY_cond $X=5.115 $Y=1.457
+ $X2=5.295 $Y2=1.457
r90 39 40 23.4436 $w=5.14e-07 $l=2.5e-07 $layer=POLY_cond $X=4.865 $Y=1.457
+ $X2=5.115 $Y2=1.457
r91 38 39 16.8794 $w=5.14e-07 $l=1.8e-07 $layer=POLY_cond $X=4.685 $Y=1.457
+ $X2=4.865 $Y2=1.457
r92 37 38 23.4436 $w=5.14e-07 $l=2.5e-07 $layer=POLY_cond $X=4.435 $Y=1.457
+ $X2=4.685 $Y2=1.457
r93 36 37 16.8794 $w=5.14e-07 $l=1.8e-07 $layer=POLY_cond $X=4.255 $Y=1.457
+ $X2=4.435 $Y2=1.457
r94 34 36 8.90856 $w=5.14e-07 $l=9.5e-08 $layer=POLY_cond $X=4.16 $Y=1.457
+ $X2=4.255 $Y2=1.457
r95 34 35 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.16
+ $Y=1.51 $X2=4.16 $Y2=1.51
r96 28 43 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.52
+ $Y=1.51 $X2=5.52 $Y2=1.51
r97 27 28 14.0044 $w=3.93e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.552
+ $X2=5.52 $Y2=1.552
r98 26 27 14.0044 $w=3.93e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.552
+ $X2=5.04 $Y2=1.552
r99 26 35 11.6703 $w=3.93e-07 $l=4e-07 $layer=LI1_cond $X=4.56 $Y=1.552 $X2=4.16
+ $Y2=1.552
r100 25 35 2.33406 $w=3.93e-07 $l=8e-08 $layer=LI1_cond $X=4.08 $Y=1.552
+ $X2=4.16 $Y2=1.552
r101 22 45 16.8794 $w=5.14e-07 $l=3.50634e-07 $layer=POLY_cond $X=5.725 $Y=1.185
+ $X2=5.545 $Y2=1.457
r102 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.725 $Y=1.185
+ $X2=5.725 $Y2=0.655
r103 19 45 32.1071 $w=1.5e-07 $l=2.68e-07 $layer=POLY_cond $X=5.545 $Y=1.725
+ $X2=5.545 $Y2=1.457
r104 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.545 $Y=1.725
+ $X2=5.545 $Y2=2.465
r105 16 41 32.1071 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.295 $Y=1.185
+ $X2=5.295 $Y2=1.457
r106 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.295 $Y=1.185
+ $X2=5.295 $Y2=0.655
r107 13 40 32.1071 $w=1.5e-07 $l=2.68e-07 $layer=POLY_cond $X=5.115 $Y=1.725
+ $X2=5.115 $Y2=1.457
r108 13 15 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.115 $Y=1.725
+ $X2=5.115 $Y2=2.465
r109 10 39 32.1071 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.865 $Y=1.185
+ $X2=4.865 $Y2=1.457
r110 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.865 $Y=1.185
+ $X2=4.865 $Y2=0.655
r111 7 38 32.1071 $w=1.5e-07 $l=2.68e-07 $layer=POLY_cond $X=4.685 $Y=1.725
+ $X2=4.685 $Y2=1.457
r112 7 9 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.685 $Y=1.725
+ $X2=4.685 $Y2=2.465
r113 4 37 32.1071 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.435 $Y=1.185
+ $X2=4.435 $Y2=1.457
r114 4 6 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.435 $Y=1.185
+ $X2=4.435 $Y2=0.655
r115 1 36 32.1071 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.255 $Y=1.73
+ $X2=4.255 $Y2=1.457
r116 1 3 236.18 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=4.255 $Y=1.73
+ $X2=4.255 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 34 38
+ 39 49
c99 20 0 8.51568e-20 $X=7.015 $Y=0.655
r100 49 50 20.8558 $w=4.16e-07 $l=1.8e-07 $layer=POLY_cond $X=7.265 $Y=1.5
+ $X2=7.445 $Y2=1.5
r101 46 47 20.8558 $w=4.16e-07 $l=1.8e-07 $layer=POLY_cond $X=6.835 $Y=1.5
+ $X2=7.015 $Y2=1.5
r102 45 46 28.9663 $w=4.16e-07 $l=2.5e-07 $layer=POLY_cond $X=6.585 $Y=1.5
+ $X2=6.835 $Y2=1.5
r103 44 45 20.8558 $w=4.16e-07 $l=1.8e-07 $layer=POLY_cond $X=6.405 $Y=1.5
+ $X2=6.585 $Y2=1.5
r104 37 49 8.11058 $w=4.16e-07 $l=7e-08 $layer=POLY_cond $X=7.195 $Y=1.5
+ $X2=7.265 $Y2=1.5
r105 37 47 20.8558 $w=4.16e-07 $l=1.8e-07 $layer=POLY_cond $X=7.195 $Y=1.5
+ $X2=7.015 $Y2=1.5
r106 36 38 4.6788 $w=3.18e-07 $l=6e-08 $layer=LI1_cond $X=7.195 $Y=1.365
+ $X2=7.135 $Y2=1.365
r107 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.195
+ $Y=1.44 $X2=7.195 $Y2=1.44
r108 34 39 5.22201 $w=3.18e-07 $l=1.45e-07 $layer=LI1_cond $X=7.295 $Y=1.365
+ $X2=7.44 $Y2=1.365
r109 34 36 3.60138 $w=3.18e-07 $l=1e-07 $layer=LI1_cond $X=7.295 $Y=1.365
+ $X2=7.195 $Y2=1.365
r110 32 44 26.649 $w=4.16e-07 $l=2.3e-07 $layer=POLY_cond $X=6.175 $Y=1.5
+ $X2=6.405 $Y2=1.5
r111 32 42 2.31731 $w=4.16e-07 $l=2e-08 $layer=POLY_cond $X=6.175 $Y=1.5
+ $X2=6.155 $Y2=1.5
r112 31 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.175 $Y=1.44
+ $X2=7.135 $Y2=1.44
r113 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.175
+ $Y=1.44 $X2=6.175 $Y2=1.44
r114 25 50 26.8236 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.445 $Y=1.275
+ $X2=7.445 $Y2=1.5
r115 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.445 $Y=1.275
+ $X2=7.445 $Y2=0.655
r116 22 49 26.8236 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.265 $Y=1.725
+ $X2=7.265 $Y2=1.5
r117 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.265 $Y=1.725
+ $X2=7.265 $Y2=2.465
r118 18 47 26.8236 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.015 $Y=1.275
+ $X2=7.015 $Y2=1.5
r119 18 20 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.015 $Y=1.275
+ $X2=7.015 $Y2=0.655
r120 15 46 26.8236 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.835 $Y=1.725
+ $X2=6.835 $Y2=1.5
r121 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.835 $Y=1.725
+ $X2=6.835 $Y2=2.465
r122 11 45 26.8236 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.585 $Y=1.275
+ $X2=6.585 $Y2=1.5
r123 11 13 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.585 $Y=1.275
+ $X2=6.585 $Y2=0.655
r124 8 44 26.8236 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.405 $Y=1.725
+ $X2=6.405 $Y2=1.5
r125 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.405 $Y=1.725
+ $X2=6.405 $Y2=2.465
r126 4 42 26.8236 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.155 $Y=1.275
+ $X2=6.155 $Y2=1.5
r127 4 6 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.155 $Y=1.275
+ $X2=6.155 $Y2=0.655
r128 1 42 20.8558 $w=4.16e-07 $l=3.01869e-07 $layer=POLY_cond $X=5.975 $Y=1.725
+ $X2=6.155 $Y2=1.5
r129 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.975 $Y=1.725
+ $X2=5.975 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 41 43
r82 65 66 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=9.505 $Y=1.46
+ $X2=9.525 $Y2=1.46
r83 63 65 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=9.45 $Y=1.46
+ $X2=9.505 $Y2=1.46
r84 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.45
+ $Y=1.46 $X2=9.45 $Y2=1.46
r85 61 63 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=9.095 $Y=1.46
+ $X2=9.45 $Y2=1.46
r86 60 61 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=9.075 $Y=1.46
+ $X2=9.095 $Y2=1.46
r87 58 60 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=8.77 $Y=1.46
+ $X2=9.075 $Y2=1.46
r88 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.77
+ $Y=1.46 $X2=8.77 $Y2=1.46
r89 56 58 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=8.665 $Y=1.46
+ $X2=8.77 $Y2=1.46
r90 55 56 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.645 $Y=1.46
+ $X2=8.665 $Y2=1.46
r91 54 59 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=8.43 $Y=1.567
+ $X2=8.77 $Y2=1.567
r92 53 55 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.43 $Y=1.46
+ $X2=8.645 $Y2=1.46
r93 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.43
+ $Y=1.46 $X2=8.43 $Y2=1.46
r94 51 53 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=8.235 $Y=1.46
+ $X2=8.43 $Y2=1.46
r95 50 51 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.215 $Y=1.46
+ $X2=8.235 $Y2=1.46
r96 47 50 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=8.09 $Y=1.46
+ $X2=8.215 $Y2=1.46
r97 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=1.46 $X2=8.09 $Y2=1.46
r98 44 64 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=9.79 $Y=1.567
+ $X2=9.45 $Y2=1.567
r99 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.79
+ $Y=1.46 $X2=9.79 $Y2=1.46
r100 41 66 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.6 $Y=1.46
+ $X2=9.525 $Y2=1.46
r101 41 43 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=9.6 $Y=1.46
+ $X2=9.79 $Y2=1.46
r102 36 44 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=9.84 $Y=1.567
+ $X2=9.79 $Y2=1.567
r103 35 64 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=9.36 $Y=1.567
+ $X2=9.45 $Y2=1.567
r104 34 35 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.567
+ $X2=9.36 $Y2=1.567
r105 34 59 3.29269 $w=3.83e-07 $l=1.1e-07 $layer=LI1_cond $X=8.88 $Y=1.567
+ $X2=8.77 $Y2=1.567
r106 33 54 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=8.4 $Y=1.567
+ $X2=8.43 $Y2=1.567
r107 33 48 9.27941 $w=3.83e-07 $l=3.1e-07 $layer=LI1_cond $X=8.4 $Y=1.567
+ $X2=8.09 $Y2=1.567
r108 29 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.525 $Y=1.295
+ $X2=9.525 $Y2=1.46
r109 29 31 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=9.525 $Y=1.295
+ $X2=9.525 $Y2=0.655
r110 25 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.505 $Y=1.625
+ $X2=9.505 $Y2=1.46
r111 25 27 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.505 $Y=1.625
+ $X2=9.505 $Y2=2.465
r112 21 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.095 $Y=1.295
+ $X2=9.095 $Y2=1.46
r113 21 23 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=9.095 $Y=1.295
+ $X2=9.095 $Y2=0.655
r114 17 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.075 $Y=1.625
+ $X2=9.075 $Y2=1.46
r115 17 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.075 $Y=1.625
+ $X2=9.075 $Y2=2.465
r116 13 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.665 $Y=1.295
+ $X2=8.665 $Y2=1.46
r117 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.665 $Y=1.295
+ $X2=8.665 $Y2=0.655
r118 9 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.625
+ $X2=8.645 $Y2=1.46
r119 9 11 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.645 $Y=1.625
+ $X2=8.645 $Y2=2.465
r120 5 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=1.295
+ $X2=8.235 $Y2=1.46
r121 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.235 $Y=1.295
+ $X2=8.235 $Y2=0.655
r122 1 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.215 $Y=1.625
+ $X2=8.215 $Y2=1.46
r123 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.215 $Y=1.625
+ $X2=8.215 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%Y 1 2 3 4 5 6 7 8 9 10 11 35 36 40 44 48
+ 52 56 60 64 66 68 70 74 76 80 82 86 88 93 94 95 96 97 103 105 106 112 117 118
+ 119 120 121 133
r146 128 133 0.426831 $w=2.68e-07 $l=1e-08 $layer=LI1_cond $X=0.22 $Y=1.675
+ $X2=0.22 $Y2=1.665
r147 121 143 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=2.775
+ $X2=0.22 $Y2=2.91
r148 120 121 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=2.405
+ $X2=0.22 $Y2=2.775
r149 119 120 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.22 $Y=1.98
+ $X2=0.22 $Y2=2.405
r150 119 134 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=1.98
+ $X2=0.22 $Y2=1.845
r151 118 128 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=1.76
+ $X2=0.22 $Y2=1.675
r152 118 134 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=1.76
+ $X2=0.22 $Y2=1.845
r153 118 133 1.62196 $w=2.68e-07 $l=3.8e-08 $layer=LI1_cond $X=0.22 $Y=1.627
+ $X2=0.22 $Y2=1.665
r154 117 118 14.1708 $w=2.68e-07 $l=3.32e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.627
r155 112 115 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=7.48 $Y=1.79
+ $X2=7.48 $Y2=2.03
r156 106 109 10.2794 $w=2.03e-07 $l=1.9e-07 $layer=LI1_cond $X=6.612 $Y=1.79
+ $X2=6.612 $Y2=1.98
r157 99 101 2.85938 $w=3.2e-07 $l=7.5e-08 $layer=LI1_cond $X=3.952 $Y=2.01
+ $X2=3.952 $Y2=2.085
r158 92 94 3.15794 $w=4.53e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.927
+ $X2=0.775 $Y2=0.927
r159 92 93 7.41179 $w=4.53e-07 $l=9.5e-08 $layer=LI1_cond $X=0.69 $Y=0.927
+ $X2=0.595 $Y2=0.927
r160 90 117 5.97563 $w=2.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.22 $Y=1.155
+ $X2=0.22 $Y2=1.295
r161 89 106 1.83547 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=6.715 $Y=1.79
+ $X2=6.612 $Y2=1.79
r162 88 112 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.315 $Y=1.79
+ $X2=7.48 $Y2=1.79
r163 88 89 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.315 $Y=1.79
+ $X2=6.715 $Y2=1.79
r164 86 111 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.62 $Y=2.56
+ $X2=6.62 $Y2=2.1
r165 83 105 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.855 $Y=2.01
+ $X2=5.76 $Y2=2.01
r166 82 111 4.94607 $w=2.03e-07 $l=9e-08 $layer=LI1_cond $X=6.612 $Y=2.01
+ $X2=6.612 $Y2=2.1
r167 82 109 1.62306 $w=2.03e-07 $l=3e-08 $layer=LI1_cond $X=6.612 $Y=2.01
+ $X2=6.612 $Y2=1.98
r168 82 83 40.3586 $w=1.78e-07 $l=6.55e-07 $layer=LI1_cond $X=6.51 $Y=2.01
+ $X2=5.855 $Y2=2.01
r169 78 105 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=5.76 $Y=2.1 $X2=5.76
+ $Y2=2.01
r170 78 80 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=5.76 $Y=2.1
+ $X2=5.76 $Y2=2.505
r171 77 103 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.995 $Y=2.01
+ $X2=4.9 $Y2=2.01
r172 76 105 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.665 $Y=2.01
+ $X2=5.76 $Y2=2.01
r173 76 77 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=5.665 $Y=2.01
+ $X2=4.995 $Y2=2.01
r174 72 103 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=4.9 $Y=2.1 $X2=4.9
+ $Y2=2.01
r175 72 74 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=4.9 $Y=2.1 $X2=4.9
+ $Y2=2.505
r176 71 99 4.1044 $w=1.8e-07 $l=1.78e-07 $layer=LI1_cond $X=4.13 $Y=2.01
+ $X2=3.952 $Y2=2.01
r177 70 103 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.805 $Y=2.01
+ $X2=4.9 $Y2=2.01
r178 70 71 41.5909 $w=1.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.805 $Y=2.01
+ $X2=4.13 $Y2=2.01
r179 66 101 2.19555 $w=5.25e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.867 $Y=2.1
+ $X2=3.952 $Y2=2.085
r180 66 68 18.4538 $w=5.23e-07 $l=8.1e-07 $layer=LI1_cond $X=3.867 $Y=2.1
+ $X2=3.867 $Y2=2.91
r181 65 97 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.935 $Y=1.76
+ $X2=2.84 $Y2=1.76
r182 64 99 9.53125 $w=3.2e-07 $l=4.55147e-07 $layer=LI1_cond $X=3.605 $Y=1.76
+ $X2=3.952 $Y2=2.01
r183 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.605 $Y=1.76
+ $X2=2.935 $Y2=1.76
r184 60 62 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.84 $Y=1.98
+ $X2=2.84 $Y2=2.91
r185 58 97 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=1.845
+ $X2=2.84 $Y2=1.76
r186 58 60 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=2.84 $Y=1.845
+ $X2=2.84 $Y2=1.98
r187 57 96 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.075 $Y=1.76
+ $X2=1.98 $Y2=1.76
r188 56 97 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.745 $Y=1.76
+ $X2=2.84 $Y2=1.76
r189 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.745 $Y=1.76
+ $X2=2.075 $Y2=1.76
r190 52 54 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.98 $Y=1.98
+ $X2=1.98 $Y2=2.91
r191 50 96 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.845
+ $X2=1.98 $Y2=1.76
r192 50 52 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.98 $Y=1.845
+ $X2=1.98 $Y2=1.98
r193 49 95 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.215 $Y=1.76
+ $X2=1.12 $Y2=1.76
r194 48 96 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.885 $Y=1.76
+ $X2=1.98 $Y2=1.76
r195 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.885 $Y=1.76
+ $X2=1.215 $Y2=1.76
r196 44 46 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.12 $Y=1.98
+ $X2=1.12 $Y2=2.91
r197 42 95 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.845
+ $X2=1.12 $Y2=1.76
r198 42 44 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.12 $Y=1.845
+ $X2=1.12 $Y2=1.98
r199 40 94 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=1.55 $Y=0.865
+ $X2=0.775 $Y2=0.865
r200 37 118 3.05049 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.355 $Y=1.76
+ $X2=0.22 $Y2=1.76
r201 36 95 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.025 $Y=1.76
+ $X2=1.12 $Y2=1.76
r202 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=1.76
+ $X2=0.355 $Y2=1.76
r203 35 90 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.355 $Y=1.07
+ $X2=0.22 $Y2=1.155
r204 35 93 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.355 $Y=1.07
+ $X2=0.595 $Y2=1.07
r205 11 115 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=7.34
+ $Y=1.835 $X2=7.48 $Y2=2.03
r206 10 109 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.835 $X2=6.62 $Y2=1.98
r207 10 86 600 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.835 $X2=6.62 $Y2=2.56
r208 9 105 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=1.835 $X2=5.76 $Y2=2.005
r209 9 80 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=5.62
+ $Y=1.835 $X2=5.76 $Y2=2.505
r210 8 103 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.76
+ $Y=1.835 $X2=4.9 $Y2=2.005
r211 8 74 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=4.76
+ $Y=1.835 $X2=4.9 $Y2=2.505
r212 7 101 200 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=3 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.085
r213 7 68 200 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=3 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.91
r214 6 62 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.91
r215 6 60 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=1.98
r216 5 54 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.91
r217 5 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=1.98
r218 4 46 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.91
r219 4 44 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=1.98
r220 3 143 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r221 3 119 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r222 2 40 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.865
r223 1 92 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%VPWR 1 2 3 4 5 6 7 8 9 30 36 42 46 50 56
+ 60 64 68 70 72 77 78 79 80 82 83 85 86 87 89 108 115 120 126 129 132 135 139
r156 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r157 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r159 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r160 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r161 124 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r162 124 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r163 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r164 121 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=8.86 $Y2=3.33
r165 121 123 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=9.36 $Y2=3.33
r166 120 138 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=9.555 $Y=3.33
+ $X2=9.817 $Y2=3.33
r167 120 123 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=9.555 $Y=3.33
+ $X2=9.36 $Y2=3.33
r168 119 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 119 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r170 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r171 116 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.165 $Y=3.33
+ $X2=8 $Y2=3.33
r172 116 118 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.165 $Y=3.33
+ $X2=8.4 $Y2=3.33
r173 115 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.86 $Y2=3.33
r174 115 118 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.4 $Y2=3.33
r175 114 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r176 113 114 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r177 111 114 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.44 $Y2=3.33
r178 110 113 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.44 $Y2=3.33
r179 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r180 108 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=8 $Y2=3.33
r181 108 113 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.44 $Y2=3.33
r182 104 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r183 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r184 101 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=3.33
+ $X2=3.27 $Y2=3.33
r185 101 103 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r186 100 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r187 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r188 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r189 97 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r190 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r191 94 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r192 94 96 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 92 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r194 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r195 89 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r196 89 91 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r197 87 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r198 87 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r199 87 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r200 85 106 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.165 $Y=3.33
+ $X2=5.04 $Y2=3.33
r201 85 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=3.33
+ $X2=5.33 $Y2=3.33
r202 84 110 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.495 $Y=3.33
+ $X2=5.52 $Y2=3.33
r203 84 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=3.33
+ $X2=5.33 $Y2=3.33
r204 82 103 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.3 $Y=3.33
+ $X2=4.08 $Y2=3.33
r205 82 83 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.3 $Y=3.33
+ $X2=4.467 $Y2=3.33
r206 81 106 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=5.04 $Y2=3.33
r207 81 83 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=4.467 $Y2=3.33
r208 79 99 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.16 $Y2=3.33
r209 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.41 $Y2=3.33
r210 77 96 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.55 $Y2=3.33
r212 76 99 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=2.16 $Y2=3.33
r213 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.55 $Y2=3.33
r214 72 75 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=9.72 $Y=2.015
+ $X2=9.72 $Y2=2.95
r215 70 138 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=9.72 $Y=3.245
+ $X2=9.817 $Y2=3.33
r216 70 75 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.72 $Y=3.245
+ $X2=9.72 $Y2=2.95
r217 66 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=3.245
+ $X2=8.86 $Y2=3.33
r218 66 68 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=8.86 $Y=3.245
+ $X2=8.86 $Y2=2.385
r219 62 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8 $Y=3.245 $X2=8
+ $Y2=3.33
r220 62 64 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8 $Y=3.245 $X2=8
+ $Y2=2.8
r221 58 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=3.245
+ $X2=5.33 $Y2=3.33
r222 58 60 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=5.33 $Y=3.245
+ $X2=5.33 $Y2=2.39
r223 54 83 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.467 $Y=3.245
+ $X2=4.467 $Y2=3.33
r224 54 56 29.4131 $w=3.33e-07 $l=8.55e-07 $layer=LI1_cond $X=4.467 $Y=3.245
+ $X2=4.467 $Y2=2.39
r225 50 53 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=3.27 $Y=2.1
+ $X2=3.27 $Y2=2.95
r226 48 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=3.245
+ $X2=3.27 $Y2=3.33
r227 48 53 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.27 $Y=3.245
+ $X2=3.27 $Y2=2.95
r228 47 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=2.41 $Y2=3.33
r229 46 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=3.27 $Y2=3.33
r230 46 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=2.575 $Y2=3.33
r231 42 45 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=2.41 $Y=2.1
+ $X2=2.41 $Y2=2.95
r232 40 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=3.245
+ $X2=2.41 $Y2=3.33
r233 40 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.41 $Y=3.245
+ $X2=2.41 $Y2=2.95
r234 36 39 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=1.55 $Y=2.1
+ $X2=1.55 $Y2=2.95
r235 34 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=3.33
r236 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=2.95
r237 30 33 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.69 $Y=2.1
+ $X2=0.69 $Y2=2.95
r238 28 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r239 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.95
r240 9 75 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.58
+ $Y=1.835 $X2=9.72 $Y2=2.95
r241 9 72 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=9.58
+ $Y=1.835 $X2=9.72 $Y2=2.015
r242 8 68 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=8.72
+ $Y=1.835 $X2=8.86 $Y2=2.385
r243 7 64 600 $w=1.7e-07 $l=1.0256e-06 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.835 $X2=8 $Y2=2.8
r244 6 60 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=1.835 $X2=5.33 $Y2=2.39
r245 5 56 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=4.33
+ $Y=1.835 $X2=4.47 $Y2=2.39
r246 4 53 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.95
r247 4 50 400 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.1
r248 3 45 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.95
r249 3 42 400 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.1
r250 2 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.95
r251 2 36 400 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.1
r252 1 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
r253 1 30 400 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.1
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%A_1210_367# 1 2 3 4 15 17 18 21 26 27 29
+ 30 33 35 37 39 41 45
r62 37 47 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.29 $Y=2.1 $X2=9.29
+ $Y2=2.015
r63 37 39 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=9.29 $Y=2.1 $X2=9.29
+ $Y2=2.91
r64 36 43 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.525 $Y=2.015
+ $X2=8.395 $Y2=2.015
r65 35 47 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.195 $Y=2.015
+ $X2=9.29 $Y2=2.015
r66 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.195 $Y=2.015
+ $X2=8.525 $Y2=2.015
r67 31 45 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=8.43 $Y=2.495
+ $X2=8.395 $Y2=2.41
r68 31 33 24.2249 $w=1.88e-07 $l=4.15e-07 $layer=LI1_cond $X=8.43 $Y=2.495
+ $X2=8.43 $Y2=2.91
r69 30 45 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=2.325
+ $X2=8.395 $Y2=2.41
r70 29 43 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=2.1
+ $X2=8.395 $Y2=2.015
r71 29 30 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=8.395 $Y=2.1
+ $X2=8.395 $Y2=2.325
r72 28 41 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.215 $Y=2.41
+ $X2=7.05 $Y2=2.41
r73 27 45 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.265 $Y=2.41
+ $X2=8.395 $Y2=2.41
r74 27 28 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=8.265 $Y=2.41
+ $X2=7.215 $Y2=2.41
r75 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.05 $Y=2.895
+ $X2=7.05 $Y2=2.56
r76 23 41 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.05 $Y=2.495
+ $X2=7.05 $Y2=2.41
r77 23 26 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=7.05 $Y=2.495
+ $X2=7.05 $Y2=2.56
r78 19 41 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=7.015 $Y=2.325
+ $X2=7.05 $Y2=2.41
r79 19 21 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=7.015 $Y=2.325
+ $X2=7.015 $Y2=2.21
r80 17 24 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=6.885 $Y=2.985
+ $X2=7.05 $Y2=2.895
r81 17 18 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=6.885 $Y=2.985
+ $X2=6.355 $Y2=2.985
r82 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=6.19 $Y=2.895
+ $X2=6.355 $Y2=2.985
r83 13 15 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.19 $Y=2.895
+ $X2=6.19 $Y2=2.39
r84 4 47 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=9.15
+ $Y=1.835 $X2=9.29 $Y2=2.095
r85 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.15
+ $Y=1.835 $X2=9.29 $Y2=2.91
r86 3 45 600 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=1 $X=8.29
+ $Y=1.835 $X2=8.43 $Y2=2.435
r87 3 43 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=8.29 $Y=1.835
+ $X2=8.43 $Y2=2.015
r88 3 33 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.29
+ $Y=1.835 $X2=8.43 $Y2=2.91
r89 2 26 300 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=2 $X=6.91
+ $Y=1.835 $X2=7.05 $Y2=2.56
r90 2 21 600 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=6.91
+ $Y=1.835 $X2=7.05 $Y2=2.21
r91 1 15 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=6.05
+ $Y=1.835 $X2=6.19 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%A_27_47# 1 2 3 4 5 16 20 24 25 28 31 38
r57 38 40 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=2.845 $Y=0.82
+ $X2=2.845 $Y2=1.07
r58 31 33 0.41907 $w=3.28e-07 $l=1.2e-08 $layer=LI1_cond $X=0.26 $Y=0.38
+ $X2=0.26 $Y2=0.392
r59 28 38 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=3.7 $Y=0.82
+ $X2=2.945 $Y2=0.82
r60 24 40 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.745 $Y=1.07 $X2=2.845
+ $Y2=1.07
r61 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.745 $Y=1.07
+ $X2=2.075 $Y2=1.07
r62 21 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.965 $Y=0.985
+ $X2=2.075 $Y2=1.07
r63 21 23 3.92878 $w=2.18e-07 $l=7.5e-08 $layer=LI1_cond $X=1.965 $Y=0.985
+ $X2=1.965 $Y2=0.91
r64 20 36 3.85427 $w=2.2e-07 $l=1.38e-07 $layer=LI1_cond $X=1.965 $Y=0.53
+ $X2=1.965 $Y2=0.392
r65 20 23 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=1.965 $Y=0.53
+ $X2=1.965 $Y2=0.91
r66 17 33 1.82517 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=0.392
+ $X2=0.26 $Y2=0.392
r67 17 19 29.1254 $w=2.73e-07 $l=6.95e-07 $layer=LI1_cond $X=0.425 $Y=0.392
+ $X2=1.12 $Y2=0.392
r68 16 36 3.07225 $w=2.75e-07 $l=1.1e-07 $layer=LI1_cond $X=1.855 $Y=0.392
+ $X2=1.965 $Y2=0.392
r69 16 19 30.8017 $w=2.73e-07 $l=7.35e-07 $layer=LI1_cond $X=1.855 $Y=0.392
+ $X2=1.12 $Y2=0.392
r70 5 28 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.82
r71 4 38 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.82
r72 3 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.42
r73 3 23 182 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.91
r74 2 19 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.4
r75 1 31 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%A_454_47# 1 2 3 4 13 19 23 29 31
c49 29 0 1.7599e-19 $X=4.65 $Y=0.38
r50 23 26 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=2.41 $Y=0.37 $X2=2.41
+ $Y2=0.38
r51 20 29 7.66117 $w=2e-07 $l=1.79374e-07 $layer=LI1_cond $X=4.815 $Y=0.34
+ $X2=4.65 $Y2=0.37
r52 19 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.345 $Y=0.34
+ $X2=5.51 $Y2=0.34
r53 19 20 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.345 $Y=0.34
+ $X2=4.815 $Y2=0.34
r54 14 23 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0.37
+ $X2=2.41 $Y2=0.37
r55 14 16 34.8238 $w=2.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.575 $Y=0.37
+ $X2=3.27 $Y2=0.37
r56 13 29 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=0.37 $X2=4.65
+ $Y2=0.37
r57 13 16 60.8791 $w=2.28e-07 $l=1.215e-06 $layer=LI1_cond $X=4.485 $Y=0.37
+ $X2=3.27 $Y2=0.37
r58 4 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.37
+ $Y=0.235 $X2=5.51 $Y2=0.38
r59 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.51
+ $Y=0.235 $X2=4.65 $Y2=0.38
r60 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.38
r61 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%A_819_47# 1 2 3 4 5 6 7 24 26 27 30 32 36
+ 38 42 44 48 50 54 56 60 62 63 64 69 71
c95 38 0 8.51568e-20 $X=6.705 $Y=1.1
r96 69 70 3.99065 $w=4.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.84 $Y=0.95
+ $X2=7.84 $Y2=1.09
r97 64 66 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=6.835 $Y=0.95
+ $X2=6.835 $Y2=1.1
r98 64 65 4.62437 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=6.835 $Y=0.95
+ $X2=6.835 $Y2=0.865
r99 58 60 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=9.775 $Y=1.005
+ $X2=9.775 $Y2=0.42
r100 57 71 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.975 $Y=1.09
+ $X2=8.88 $Y2=1.09
r101 56 58 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.645 $Y=1.09
+ $X2=9.775 $Y2=1.005
r102 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.645 $Y=1.09
+ $X2=8.975 $Y2=1.09
r103 52 71 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.88 $Y=1.005
+ $X2=8.88 $Y2=1.09
r104 52 54 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=8.88 $Y=1.005
+ $X2=8.88 $Y2=0.42
r105 51 70 6.19161 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=8.115 $Y=1.09
+ $X2=7.84 $Y2=1.09
r106 50 71 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.785 $Y=1.09
+ $X2=8.88 $Y2=1.09
r107 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.785 $Y=1.09
+ $X2=8.115 $Y2=1.09
r108 46 69 2.51835 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.84 $Y=0.865
+ $X2=7.84 $Y2=0.95
r109 46 48 9.67736 $w=5.48e-07 $l=4.45e-07 $layer=LI1_cond $X=7.84 $Y=0.865
+ $X2=7.84 $Y2=0.42
r110 45 64 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.965 $Y=0.95
+ $X2=6.835 $Y2=0.95
r111 44 69 6.19161 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=7.565 $Y=0.95
+ $X2=7.84 $Y2=0.95
r112 44 45 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.565 $Y=0.95
+ $X2=6.965 $Y2=0.95
r113 42 65 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=6.8 $Y=0.42
+ $X2=6.8 $Y2=0.865
r114 39 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.035 $Y=1.1
+ $X2=5.94 $Y2=1.1
r115 38 66 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.705 $Y=1.1
+ $X2=6.835 $Y2=1.1
r116 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.705 $Y=1.1
+ $X2=6.035 $Y2=1.1
r117 34 63 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=1.015
+ $X2=5.94 $Y2=1.1
r118 34 36 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=5.94 $Y=1.015
+ $X2=5.94 $Y2=0.42
r119 33 62 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.175 $Y=1.1
+ $X2=5.08 $Y2=1.1
r120 32 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.845 $Y=1.1
+ $X2=5.94 $Y2=1.1
r121 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.845 $Y=1.1
+ $X2=5.175 $Y2=1.1
r122 28 62 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=1.015
+ $X2=5.08 $Y2=1.1
r123 28 30 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=5.08 $Y=1.015
+ $X2=5.08 $Y2=0.76
r124 26 62 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.985 $Y=1.1
+ $X2=5.08 $Y2=1.1
r125 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.985 $Y=1.1
+ $X2=4.315 $Y2=1.1
r126 22 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.185 $Y=1.015
+ $X2=4.315 $Y2=1.1
r127 22 24 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=4.185 $Y=1.015
+ $X2=4.185 $Y2=0.82
r128 7 60 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.6
+ $Y=0.235 $X2=9.74 $Y2=0.42
r129 6 54 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.74
+ $Y=0.235 $X2=8.88 $Y2=0.42
r130 5 69 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=7.52
+ $Y=0.235 $X2=7.66 $Y2=0.95
r131 5 48 60.6667 $w=1.7e-07 $l=5.85235e-07 $layer=licon1_NDIFF $count=3 $X=7.52
+ $Y=0.235 $X2=8.02 $Y2=0.42
r132 4 42 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.66
+ $Y=0.235 $X2=6.8 $Y2=0.42
r133 3 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.8
+ $Y=0.235 $X2=5.94 $Y2=0.42
r134 2 30 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.235 $X2=5.08 $Y2=0.76
r135 1 24 182 $w=1.7e-07 $l=6.44477e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.22 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 47
+ 51 58 59 62 65
r120 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r121 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r122 59 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r123 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r124 56 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=0 $X2=9.31
+ $Y2=0
r125 56 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.475 $Y=0
+ $X2=9.84 $Y2=0
r126 55 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r127 55 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r128 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r129 52 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=0 $X2=8.45
+ $Y2=0
r130 52 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.615 $Y=0
+ $X2=8.88 $Y2=0
r131 51 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=0 $X2=9.31
+ $Y2=0
r132 51 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.145 $Y=0
+ $X2=8.88 $Y2=0
r133 50 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r134 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r135 47 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=0 $X2=8.45
+ $Y2=0
r136 47 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.285 $Y=0
+ $X2=7.92 $Y2=0
r137 46 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r138 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r139 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r140 42 43 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=6 $Y=0 $X2=6
+ $Y2=0
r141 38 42 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=6
+ $Y2=0
r142 38 39 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r143 35 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r144 35 39 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=0.24
+ $Y2=0
r145 33 45 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.065 $Y=0
+ $X2=6.96 $Y2=0
r146 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.065 $Y=0 $X2=7.23
+ $Y2=0
r147 32 49 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.395 $Y=0
+ $X2=7.92 $Y2=0
r148 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.395 $Y=0 $X2=7.23
+ $Y2=0
r149 30 42 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6
+ $Y2=0
r150 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.37
+ $Y2=0
r151 29 45 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.535 $Y=0
+ $X2=6.96 $Y2=0
r152 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=0 $X2=6.37
+ $Y2=0
r153 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=0.085
+ $X2=9.31 $Y2=0
r154 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.31 $Y=0.085
+ $X2=9.31 $Y2=0.38
r155 21 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=0.085
+ $X2=8.45 $Y2=0
r156 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.45 $Y=0.085
+ $X2=8.45 $Y2=0.38
r157 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.23 $Y=0.085
+ $X2=7.23 $Y2=0
r158 17 19 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=7.23 $Y=0.085
+ $X2=7.23 $Y2=0.575
r159 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0
r160 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0.38
r161 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.17
+ $Y=0.235 $X2=9.31 $Y2=0.38
r162 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.31
+ $Y=0.235 $X2=8.45 $Y2=0.38
r163 2 19 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=7.09
+ $Y=0.235 $X2=7.23 $Y2=0.575
r164 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.23
+ $Y=0.235 $X2=6.37 $Y2=0.38
.ends

