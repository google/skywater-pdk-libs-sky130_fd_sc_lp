* File: sky130_fd_sc_lp__a21boi_m.pex.spice
* Created: Wed Sep  2 09:19:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BOI_M%B1_N 3 7 11 12 13 14 15 16 22
r35 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.565
+ $Y=0.97 $X2=0.565 $Y2=0.97
r36 15 16 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.642 $Y=1.665
+ $X2=0.642 $Y2=2.035
r37 14 15 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.642 $Y=1.295
+ $X2=0.642 $Y2=1.665
r38 14 23 11.5244 $w=3.23e-07 $l=3.25e-07 $layer=LI1_cond $X=0.642 $Y=1.295
+ $X2=0.642 $Y2=0.97
r39 13 23 1.59569 $w=3.23e-07 $l=4.5e-08 $layer=LI1_cond $X=0.642 $Y=0.925
+ $X2=0.642 $Y2=0.97
r40 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.565 $Y=1.31
+ $X2=0.565 $Y2=0.97
r41 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.31
+ $X2=0.565 $Y2=1.475
r42 10 22 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=0.805
+ $X2=0.565 $Y2=0.97
r43 7 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=0.615 $Y=0.445
+ $X2=0.615 $Y2=0.805
r44 3 12 723 $w=1.5e-07 $l=1.41e-06 $layer=POLY_cond $X=0.475 $Y=2.885 $X2=0.475
+ $Y2=1.475
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_M%A_27_535# 1 2 8 11 13 15 17 18 20 23 25 29
+ 30 35 37
c65 15 0 7.39264e-20 $X=1.455 $Y=1.865
r66 32 35 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.215 $Y=0.46
+ $X2=0.4 $Y2=0.46
r67 30 38 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.14 $Y=2.9
+ $X2=0.965 $Y2=2.9
r68 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=2.9 $X2=1.14 $Y2=2.9
r69 27 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.14 $Y=2.665
+ $X2=1.14 $Y2=2.9
r70 26 37 1.79375 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.345 $Y=2.58
+ $X2=0.237 $Y2=2.58
r71 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.055 $Y=2.58
+ $X2=1.14 $Y2=2.665
r72 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.055 $Y=2.58
+ $X2=0.345 $Y2=2.58
r73 21 37 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=0.237 $Y=2.665
+ $X2=0.237 $Y2=2.58
r74 21 23 8.30831 $w=2.13e-07 $l=1.55e-07 $layer=LI1_cond $X=0.237 $Y=2.665
+ $X2=0.237 $Y2=2.82
r75 20 37 4.65272 $w=1.92e-07 $l=9.53677e-08 $layer=LI1_cond $X=0.215 $Y=2.495
+ $X2=0.237 $Y2=2.58
r76 19 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=0.625
+ $X2=0.215 $Y2=0.46
r77 19 20 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=0.215 $Y=0.625
+ $X2=0.215 $Y2=2.495
r78 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.455 $Y=1.865
+ $X2=1.455 $Y2=2.185
r79 14 18 5.30422 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.12 $Y=1.79
+ $X2=1.005 $Y2=1.79
r80 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.38 $Y=1.79
+ $X2=1.455 $Y2=1.865
r81 13 14 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.38 $Y=1.79
+ $X2=1.12 $Y2=1.79
r82 9 18 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=1.045 $Y=1.715
+ $X2=1.005 $Y2=1.79
r83 9 11 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=1.045 $Y=1.715
+ $X2=1.045 $Y2=0.445
r84 8 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=2.735
+ $X2=0.965 $Y2=2.9
r85 7 18 20.4101 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=0.965 $Y=1.865
+ $X2=1.005 $Y2=1.79
r86 7 8 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.965 $Y=1.865
+ $X2=0.965 $Y2=2.735
r87 2 23 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.82
r88 1 35 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.235 $X2=0.4 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_M%A1 3 11 13 14 15 16 17 18 19 24
c49 17 0 1.80356e-19 $X=1.68 $Y=0.555
c50 11 0 2.75185e-20 $X=1.885 $Y=2.185
c51 3 0 3.40444e-20 $X=1.475 $Y=0.445
r52 24 26 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.587 $Y=0.97
+ $X2=1.587 $Y2=0.805
r53 18 19 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=0.925
+ $X2=1.645 $Y2=1.295
r54 18 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=0.97 $X2=1.61 $Y2=0.97
r55 17 18 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=0.555
+ $X2=1.645 $Y2=0.925
r56 15 16 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.865 $Y=1.675
+ $X2=1.865 $Y2=1.825
r57 14 15 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.845 $Y=1.475
+ $X2=1.845 $Y2=1.675
r58 13 14 42.9311 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=1.66 $Y=1.325
+ $X2=1.66 $Y2=1.475
r59 11 16 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.885 $Y=2.185
+ $X2=1.885 $Y2=1.825
r60 5 24 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.587 $Y=0.992
+ $X2=1.587 $Y2=0.97
r61 5 13 49.3865 $w=3.75e-07 $l=3.33e-07 $layer=POLY_cond $X=1.587 $Y=0.992
+ $X2=1.587 $Y2=1.325
r62 3 26 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.475 $Y=0.445
+ $X2=1.475 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_M%A2 3 6 9 10 12 13 14 18
c34 13 0 3.40444e-20 $X=2.16 $Y=0.925
c35 6 0 1.80356e-19 $X=2.315 $Y=2.185
r36 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.295
+ $Y=0.93 $X2=2.295 $Y2=0.93
r37 14 19 13.7915 $w=3.03e-07 $l=3.65e-07 $layer=LI1_cond $X=2.227 $Y=1.295
+ $X2=2.227 $Y2=0.93
r38 13 19 0.188925 $w=3.03e-07 $l=5e-09 $layer=LI1_cond $X=2.227 $Y=0.925
+ $X2=2.227 $Y2=0.93
r39 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.295 $Y=1.27
+ $X2=2.295 $Y2=0.93
r40 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.27
+ $X2=2.295 $Y2=1.435
r41 10 18 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.295 $Y=0.915
+ $X2=2.295 $Y2=0.93
r42 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.222 $Y=0.765
+ $X2=2.222 $Y2=0.915
r43 6 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.315 $Y=2.185
+ $X2=2.315 $Y2=1.435
r44 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.06 $Y=0.445 $X2=2.06
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_M%VPWR 1 2 9 13 15 17 22 29 30 33 36
r33 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.1 $Y2=3.33
r38 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r42 23 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.1 $Y2=3.33
r44 22 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r48 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=3.245 $X2=2.1
+ $Y2=3.33
r52 11 13 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=2.1 $Y=3.245
+ $X2=2.1 $Y2=2.25
r53 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r54 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.95
r55 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.975 $X2=2.1 $Y2=2.25
r56 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.675 $X2=0.69 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_M%Y 1 2 7 8 9 10 11 18
c22 18 0 2.75185e-20 $X=1.26 $Y=0.43
r23 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.23 $Y=1.665
+ $X2=1.23 $Y2=2.035
r24 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.23 $Y=1.295
+ $X2=1.23 $Y2=1.665
r25 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.23 $Y=0.925 $X2=1.23
+ $Y2=1.295
r26 7 8 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.23 $Y=0.555 $X2=1.23
+ $Y2=0.925
r27 7 18 6.26328 $w=2.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.23 $Y=0.555
+ $X2=1.23 $Y2=0.43
r28 2 11 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.975 $X2=1.24 $Y2=2.12
r29 1 18 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.235 $X2=1.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_M%A_306_395# 1 2 9 11 12 15
c18 9 0 1.97726e-19 $X=1.67 $Y=2.12
r19 13 15 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.54 $Y=1.965
+ $X2=2.54 $Y2=2.12
r20 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.445 $Y=1.88
+ $X2=2.54 $Y2=1.965
r21 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.445 $Y=1.88
+ $X2=1.755 $Y2=1.88
r22 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.66 $Y=1.965
+ $X2=1.755 $Y2=1.88
r23 7 9 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.66 $Y=1.965
+ $X2=1.66 $Y2=2.12
r24 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.975 $X2=2.53 $Y2=2.12
r25 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.975 $X2=1.67 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_M%VGND 1 2 9 13 16 17 18 24 30 31 34
r38 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r40 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=0 $X2=2.275
+ $Y2=0
r42 28 30 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.44 $Y=0 $X2=2.64
+ $Y2=0
r43 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.275
+ $Y2=0
r45 24 26 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.2
+ $Y2=0
r46 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r47 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 18 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r49 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r50 16 21 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.72
+ $Y2=0
r51 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.83
+ $Y2=0
r52 15 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.2
+ $Y2=0
r53 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.83
+ $Y2=0
r54 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0.085
+ $X2=2.275 $Y2=0
r55 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.275 $Y=0.085
+ $X2=2.275 $Y2=0.38
r56 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0
r57 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0.38
r58 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.235 $X2=2.275 $Y2=0.38
r59 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.235 $X2=0.83 $Y2=0.38
.ends

