* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfstp_lp CLK D SET_B VGND VNB VPB VPWR Q
M1000 VPWR a_1731_99# a_1726_419# VPB phighvt w=1e+06u l=250000u
+  ad=3.06e+12p pd=2.012e+07u as=2.9e+11p ps=2.58e+06u
M1001 a_2374_74# a_1526_125# a_2287_74# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1002 a_1448_125# a_709_419# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=9.72e+11p ps=1.068e+07u
M1003 VGND a_1526_125# a_2374_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Q a_2287_74# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1005 a_135_409# D VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.7e+11p pd=5.14e+06u as=0p ps=0u
M1006 Q a_2287_74# a_2532_74# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1007 VGND SET_B a_1256_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VGND a_943_321# a_904_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 a_1526_125# a_266_409# a_1448_419# VPB phighvt w=1e+06u l=250000u
+  ad=9.35e+11p pd=5.87e+06u as=2.4e+11p ps=2.48e+06u
M1010 a_135_409# D a_110_57# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=8.82e+10p ps=1.26e+06u
M1011 a_479_409# a_266_409# a_531_109# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1012 a_943_321# a_709_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1013 VGND CLK a_373_109# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1014 a_531_109# a_266_409# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_2532_74# a_2287_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_1526_125# a_2287_74# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1017 a_904_125# a_479_409# a_709_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.701e+11p ps=1.65e+06u
M1018 a_479_409# a_266_409# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1019 a_1256_125# a_709_419# a_943_321# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1020 a_1761_125# a_1731_99# a_1683_125# VNB nshort w=420000u l=150000u
+  ad=2.121e+11p pd=1.85e+06u as=1.008e+11p ps=1.32e+06u
M1021 a_709_419# a_479_409# a_135_409# VPB phighvt w=1e+06u l=250000u
+  ad=6.1e+11p pd=3.22e+06u as=0p ps=0u
M1022 a_110_57# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_373_109# CLK a_266_409# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1024 a_1726_419# a_479_409# a_1526_125# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR SET_B a_943_321# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_881_419# a_266_409# a_709_419# VPB phighvt w=1e+06u l=250000u
+  ad=3.1e+11p pd=2.62e+06u as=0p ps=0u
M1027 VPWR a_943_321# a_881_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_709_419# a_266_409# a_135_409# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR CLK a_266_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1030 a_1526_125# a_479_409# a_1448_125# VNB nshort w=420000u l=150000u
+  ad=2.667e+11p pd=2.11e+06u as=0p ps=0u
M1031 a_1448_419# a_709_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1683_125# a_266_409# a_1526_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1526_125# SET_B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_1526_125# a_1731_99# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1035 a_2104_47# a_1526_125# a_1731_99# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1036 VGND SET_B a_1761_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_1526_125# a_2104_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
