* File: sky130_fd_sc_lp__dlxbn_1.pxi.spice
* Created: Wed Sep  2 09:47:51 2020
* 
x_PM_SKY130_FD_SC_LP__DLXBN_1%D N_D_M1012_g N_D_M1015_g N_D_c_145_n N_D_c_146_n
+ N_D_c_151_n D D N_D_c_148_n PM_SKY130_FD_SC_LP__DLXBN_1%D
x_PM_SKY130_FD_SC_LP__DLXBN_1%GATE_N N_GATE_N_c_180_n N_GATE_N_M1008_g
+ N_GATE_N_M1005_g N_GATE_N_c_182_n N_GATE_N_c_183_n N_GATE_N_c_184_n GATE_N
+ GATE_N N_GATE_N_c_186_n PM_SKY130_FD_SC_LP__DLXBN_1%GATE_N
x_PM_SKY130_FD_SC_LP__DLXBN_1%A_219_135# N_A_219_135#_M1008_d
+ N_A_219_135#_M1005_d N_A_219_135#_M1014_g N_A_219_135#_M1010_g
+ N_A_219_135#_M1011_g N_A_219_135#_c_226_n N_A_219_135#_c_227_n
+ N_A_219_135#_M1006_g N_A_219_135#_c_228_n N_A_219_135#_c_239_n
+ N_A_219_135#_c_229_n N_A_219_135#_c_230_n N_A_219_135#_c_231_n
+ N_A_219_135#_c_232_n N_A_219_135#_c_233_n N_A_219_135#_c_234_n
+ PM_SKY130_FD_SC_LP__DLXBN_1%A_219_135#
x_PM_SKY130_FD_SC_LP__DLXBN_1%A_34_407# N_A_34_407#_M1015_s N_A_34_407#_M1012_s
+ N_A_34_407#_c_332_n N_A_34_407#_M1019_g N_A_34_407#_M1021_g
+ N_A_34_407#_c_339_n N_A_34_407#_c_340_n N_A_34_407#_c_334_n
+ N_A_34_407#_c_342_n N_A_34_407#_c_335_n N_A_34_407#_c_336_n
+ N_A_34_407#_c_343_n PM_SKY130_FD_SC_LP__DLXBN_1%A_34_407#
x_PM_SKY130_FD_SC_LP__DLXBN_1%A_363_483# N_A_363_483#_M1010_s
+ N_A_363_483#_M1014_s N_A_363_483#_M1000_g N_A_363_483#_M1002_g
+ N_A_363_483#_c_409_n N_A_363_483#_c_429_n N_A_363_483#_c_410_n
+ N_A_363_483#_c_411_n N_A_363_483#_c_417_n N_A_363_483#_c_412_n
+ N_A_363_483#_c_419_n N_A_363_483#_c_420_n N_A_363_483#_c_421_n
+ N_A_363_483#_c_413_n N_A_363_483#_c_414_n N_A_363_483#_c_415_n
+ PM_SKY130_FD_SC_LP__DLXBN_1%A_363_483#
x_PM_SKY130_FD_SC_LP__DLXBN_1%A_806_385# N_A_806_385#_M1017_d
+ N_A_806_385#_M1020_d N_A_806_385#_M1009_g N_A_806_385#_M1007_g
+ N_A_806_385#_M1004_g N_A_806_385#_M1016_g N_A_806_385#_c_524_n
+ N_A_806_385#_M1003_g N_A_806_385#_M1013_g N_A_806_385#_c_526_n
+ N_A_806_385#_c_542_n N_A_806_385#_c_543_n N_A_806_385#_c_544_n
+ N_A_806_385#_c_527_n N_A_806_385#_c_528_n N_A_806_385#_c_529_n
+ N_A_806_385#_c_530_n N_A_806_385#_c_531_n N_A_806_385#_c_532_n
+ N_A_806_385#_c_634_p N_A_806_385#_c_533_n N_A_806_385#_c_635_p
+ N_A_806_385#_c_534_n N_A_806_385#_c_535_n N_A_806_385#_c_546_n
+ N_A_806_385#_c_536_n N_A_806_385#_c_537_n
+ PM_SKY130_FD_SC_LP__DLXBN_1%A_806_385#
x_PM_SKY130_FD_SC_LP__DLXBN_1%A_626_47# N_A_626_47#_M1011_d N_A_626_47#_M1000_d
+ N_A_626_47#_M1017_g N_A_626_47#_M1020_g N_A_626_47#_c_682_n
+ N_A_626_47#_c_669_n N_A_626_47#_c_670_n N_A_626_47#_c_671_n
+ N_A_626_47#_c_676_n N_A_626_47#_c_677_n N_A_626_47#_c_672_n
+ N_A_626_47#_c_673_n PM_SKY130_FD_SC_LP__DLXBN_1%A_626_47#
x_PM_SKY130_FD_SC_LP__DLXBN_1%A_1069_161# N_A_1069_161#_M1004_s
+ N_A_1069_161#_M1016_s N_A_1069_161#_M1001_g N_A_1069_161#_c_752_n
+ N_A_1069_161#_M1018_g N_A_1069_161#_c_753_n N_A_1069_161#_c_758_n
+ N_A_1069_161#_c_754_n N_A_1069_161#_c_755_n N_A_1069_161#_c_756_n
+ PM_SKY130_FD_SC_LP__DLXBN_1%A_1069_161#
x_PM_SKY130_FD_SC_LP__DLXBN_1%VPWR N_VPWR_M1012_d N_VPWR_M1014_d N_VPWR_M1009_d
+ N_VPWR_M1016_d N_VPWR_M1013_s N_VPWR_c_803_n N_VPWR_c_804_n N_VPWR_c_805_n
+ N_VPWR_c_806_n N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_809_n VPWR
+ N_VPWR_c_810_n N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_802_n
+ N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n
+ PM_SKY130_FD_SC_LP__DLXBN_1%VPWR
x_PM_SKY130_FD_SC_LP__DLXBN_1%Q_N N_Q_N_M1018_d N_Q_N_M1001_d Q_N Q_N Q_N Q_N
+ N_Q_N_c_890_n N_Q_N_c_893_n Q_N PM_SKY130_FD_SC_LP__DLXBN_1%Q_N
x_PM_SKY130_FD_SC_LP__DLXBN_1%Q N_Q_M1003_d N_Q_M1013_d Q Q Q Q Q Q Q
+ N_Q_c_914_n PM_SKY130_FD_SC_LP__DLXBN_1%Q
x_PM_SKY130_FD_SC_LP__DLXBN_1%VGND N_VGND_M1015_d N_VGND_M1010_d N_VGND_M1007_d
+ N_VGND_M1004_d N_VGND_M1003_s N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n
+ N_VGND_c_928_n N_VGND_c_929_n N_VGND_c_930_n N_VGND_c_931_n VGND
+ N_VGND_c_932_n N_VGND_c_933_n N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n
+ N_VGND_c_937_n N_VGND_c_938_n N_VGND_c_939_n N_VGND_c_940_n
+ PM_SKY130_FD_SC_LP__DLXBN_1%VGND
cc_1 VNB N_D_c_145_n 0.0218055f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.205
cc_2 VNB N_D_c_146_n 0.0198777f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.71
cc_3 VNB D 0.00577315f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_D_c_148_n 0.0164827f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_5 VNB N_GATE_N_c_180_n 0.0167393f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.875
cc_6 VNB N_GATE_N_M1005_g 0.011698f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.885
cc_7 VNB N_GATE_N_c_182_n 0.0283204f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_8 VNB N_GATE_N_c_183_n 0.0384846f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.875
cc_9 VNB N_GATE_N_c_184_n 0.00509755f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB GATE_N 0.0150465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_GATE_N_c_186_n 0.0432785f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_12 VNB N_A_219_135#_M1010_g 0.0455083f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_A_219_135#_M1011_g 0.0287021f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_14 VNB N_A_219_135#_c_226_n 0.0202302f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.295
cc_15 VNB N_A_219_135#_c_227_n 0.00520594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_219_135#_c_228_n 0.0242497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_219_135#_c_229_n 0.0253129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_219_135#_c_230_n 0.0217828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_219_135#_c_231_n 0.0166166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_219_135#_c_232_n 0.0231191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_219_135#_c_233_n 0.00288707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_219_135#_c_234_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_34_407#_c_332_n 0.0114334f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.885
cc_24 VNB N_A_34_407#_M1019_g 0.0521059f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.205
cc_25 VNB N_A_34_407#_c_334_n 0.029301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_34_407#_c_335_n 0.00153612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_34_407#_c_336_n 0.0171626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_363_483#_c_409_n 3.37108e-19 $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_29 VNB N_A_363_483#_c_410_n 0.0182094f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.37
cc_30 VNB N_A_363_483#_c_411_n 0.0043111f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.665
cc_31 VNB N_A_363_483#_c_412_n 0.00714088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_363_483#_c_413_n 0.00792841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_363_483#_c_414_n 0.0338754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_363_483#_c_415_n 0.017507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_806_385#_M1007_g 0.0673556f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_36 VNB N_A_806_385#_M1004_g 0.0183619f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_37 VNB N_A_806_385#_M1016_g 0.00835978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_806_385#_c_524_n 0.0222319f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.665
cc_39 VNB N_A_806_385#_M1013_g 0.00904732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_806_385#_c_526_n 0.0289248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_806_385#_c_527_n 0.0116959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_806_385#_c_528_n 0.017012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_806_385#_c_529_n 0.00207371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_806_385#_c_530_n 0.00118507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_806_385#_c_531_n 0.00538939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_806_385#_c_532_n 8.03598e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_806_385#_c_533_n 0.0113152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_806_385#_c_534_n 0.0079729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_806_385#_c_535_n 0.0163178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_806_385#_c_536_n 0.0434513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_806_385#_c_537_n 0.050715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_626_47#_M1017_g 0.0258472f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.205
cc_53 VNB N_A_626_47#_M1020_g 0.00191515f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_54 VNB N_A_626_47#_c_669_n 0.00735507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_626_47#_c_670_n 0.0045176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_626_47#_c_671_n 0.0103892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_626_47#_c_672_n 0.00457452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_626_47#_c_673_n 0.0403072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1069_161#_c_752_n 0.0215208f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.875
cc_60 VNB N_A_1069_161#_c_753_n 0.00349127f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_61 VNB N_A_1069_161#_c_754_n 0.0130947f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.37
cc_62 VNB N_A_1069_161#_c_755_n 0.00563247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1069_161#_c_756_n 0.0370715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VPWR_c_802_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_Q_N_c_890_n 0.00811918f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.37
cc_66 VNB N_Q_c_914_n 0.0616047f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.37
cc_67 VNB N_VGND_c_925_n 0.0234406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_926_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_927_n 0.00854953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_928_n 0.00961787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_929_n 0.0072037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_930_n 0.0349409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_931_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_932_n 0.0349032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_933_n 0.0404774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_934_n 0.0290439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_935_n 0.0153759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_936_n 0.441502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_937_n 0.0261816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_938_n 0.0043639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_939_n 0.00480879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_940_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VPB N_D_M1012_g 0.0249077f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.355
cc_84 VPB N_D_c_146_n 0.00377957f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.71
cc_85 VPB N_D_c_151_n 0.0165315f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.875
cc_86 VPB D 0.00534353f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_87 VPB N_GATE_N_M1005_g 0.0456853f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.885
cc_88 VPB N_A_219_135#_M1014_g 0.0542749f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.205
cc_89 VPB N_A_219_135#_c_226_n 0.013235f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.295
cc_90 VPB N_A_219_135#_c_227_n 0.00940645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_219_135#_M1006_g 0.0439739f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.665
cc_92 VPB N_A_219_135#_c_239_n 0.019132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_219_135#_c_231_n 0.0113881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_219_135#_c_232_n 0.0059416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_219_135#_c_233_n 0.00236334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_34_407#_c_332_n 0.00904671f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.885
cc_97 VPB N_A_34_407#_M1021_g 0.0210351f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_98 VPB N_A_34_407#_c_339_n 0.0280315f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.37
cc_99 VPB N_A_34_407#_c_340_n 0.0294307f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.37
cc_100 VPB N_A_34_407#_c_334_n 0.0184677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_34_407#_c_342_n 0.0318628f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.665
cc_102 VPB N_A_34_407#_c_343_n 0.0308856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_363_483#_M1000_g 0.0210606f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.205
cc_104 VPB N_A_363_483#_c_417_n 0.0019004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_363_483#_c_412_n 0.00482247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_363_483#_c_419_n 0.0195218f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_363_483#_c_420_n 0.030451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_363_483#_c_421_n 0.00664253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_806_385#_M1009_g 0.0211237f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.205
cc_110 VPB N_A_806_385#_M1007_g 0.0173485f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_111 VPB N_A_806_385#_M1016_g 0.0265814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_806_385#_M1013_g 0.0267896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_806_385#_c_542_n 0.00378908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_806_385#_c_543_n 0.0328533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_806_385#_c_544_n 0.0242479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_806_385#_c_527_n 0.00484125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_806_385#_c_546_n 0.00469391f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_626_47#_M1020_g 0.027811f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_119 VPB N_A_626_47#_c_669_n 0.00428973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_626_47#_c_676_n 0.0106156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_626_47#_c_677_n 0.00488352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_1069_161#_M1001_g 0.0255532f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.205
cc_123 VPB N_A_1069_161#_c_758_n 0.0166367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_1069_161#_c_756_n 0.014833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_803_n 0.0307245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_804_n 0.00691608f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_805_n 0.0109642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_806_n 0.0276359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_807_n 0.0196182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_808_n 0.03935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_809_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_810_n 0.0396624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_811_n 0.041233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_812_n 0.0253121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_813_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_802_n 0.142771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_815_n 0.0272595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_816_n 0.00631679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_817_n 0.0115116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_818_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB Q_N 0.0217658f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.37
cc_142 VPB N_Q_N_c_890_n 0.00432459f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.37
cc_143 VPB N_Q_N_c_893_n 0.00712988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_Q_c_914_n 0.0567722f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.37
cc_145 N_D_c_145_n N_GATE_N_c_180_n 0.0104584f $X=0.54 $Y=1.205 $X2=-0.19
+ $Y2=-0.245
cc_146 N_D_M1012_g N_GATE_N_M1005_g 0.0246231f $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_147 N_D_c_146_n N_GATE_N_M1005_g 0.0168341f $X=0.54 $Y=1.71 $X2=0 $Y2=0
cc_148 D N_GATE_N_c_184_n 0.00508695f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_149 N_D_c_148_n N_GATE_N_c_184_n 0.0168341f $X=0.54 $Y=1.37 $X2=0 $Y2=0
cc_150 N_D_M1012_g N_A_219_135#_c_231_n 3.24225e-19 $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_151 N_D_c_145_n N_A_219_135#_c_231_n 8.13037e-19 $X=0.54 $Y=1.205 $X2=0 $Y2=0
cc_152 D N_A_219_135#_c_231_n 0.0574673f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_153 N_D_c_148_n N_A_219_135#_c_231_n 4.95803e-19 $X=0.54 $Y=1.37 $X2=0 $Y2=0
cc_154 N_D_M1012_g N_A_34_407#_c_334_n 0.0056781f $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_155 N_D_c_145_n N_A_34_407#_c_334_n 0.00491281f $X=0.54 $Y=1.205 $X2=0 $Y2=0
cc_156 D N_A_34_407#_c_334_n 0.0492754f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_157 N_D_c_148_n N_A_34_407#_c_334_n 0.0163648f $X=0.54 $Y=1.37 $X2=0 $Y2=0
cc_158 N_D_M1012_g N_A_34_407#_c_342_n 0.0115818f $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_159 N_D_c_151_n N_A_34_407#_c_342_n 6.28752e-19 $X=0.54 $Y=1.875 $X2=0 $Y2=0
cc_160 D N_A_34_407#_c_342_n 0.0250465f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_161 D N_A_34_407#_c_336_n 0.00214036f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_162 N_D_c_148_n N_A_34_407#_c_336_n 0.00382023f $X=0.54 $Y=1.37 $X2=0 $Y2=0
cc_163 N_D_M1012_g N_A_34_407#_c_343_n 0.00956472f $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_164 N_D_c_151_n N_A_34_407#_c_343_n 0.00149883f $X=0.54 $Y=1.875 $X2=0 $Y2=0
cc_165 N_D_M1012_g N_VPWR_c_803_n 0.00441455f $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_166 N_D_M1012_g N_VPWR_c_802_n 0.0046122f $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_167 N_D_M1012_g N_VPWR_c_815_n 0.00385415f $X=0.51 $Y=2.355 $X2=0 $Y2=0
cc_168 N_D_c_145_n N_VGND_c_925_n 0.00341439f $X=0.54 $Y=1.205 $X2=0 $Y2=0
cc_169 D N_VGND_c_925_n 0.0173091f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_170 N_D_c_145_n N_VGND_c_936_n 0.00455831f $X=0.54 $Y=1.205 $X2=0 $Y2=0
cc_171 N_D_c_145_n N_VGND_c_937_n 0.00389919f $X=0.54 $Y=1.205 $X2=0 $Y2=0
cc_172 N_GATE_N_c_183_n N_A_219_135#_M1010_g 0.0102276f $X=1.51 $Y=1.205 $X2=0
+ $Y2=0
cc_173 N_GATE_N_c_186_n N_A_219_135#_M1010_g 0.00456655f $X=1.6 $Y=0.4 $X2=0
+ $Y2=0
cc_174 N_GATE_N_c_183_n N_A_219_135#_c_228_n 0.00354455f $X=1.51 $Y=1.205 $X2=0
+ $Y2=0
cc_175 N_GATE_N_c_180_n N_A_219_135#_c_231_n 0.0070368f $X=1.02 $Y=1.205 $X2=0
+ $Y2=0
cc_176 N_GATE_N_M1005_g N_A_219_135#_c_231_n 0.0213117f $X=1.02 $Y=2.355 $X2=0
+ $Y2=0
cc_177 N_GATE_N_c_182_n N_A_219_135#_c_231_n 0.0233928f $X=1.435 $Y=1.28 $X2=0
+ $Y2=0
cc_178 N_GATE_N_c_183_n N_A_219_135#_c_231_n 0.0180991f $X=1.51 $Y=1.205 $X2=0
+ $Y2=0
cc_179 N_GATE_N_c_184_n N_A_219_135#_c_231_n 0.00152591f $X=1.02 $Y=1.28 $X2=0
+ $Y2=0
cc_180 GATE_N N_A_219_135#_c_231_n 0.0453727f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_181 N_GATE_N_c_186_n N_A_219_135#_c_231_n 9.97905e-19 $X=1.6 $Y=0.4 $X2=0
+ $Y2=0
cc_182 N_GATE_N_c_182_n N_A_219_135#_c_232_n 0.00354455f $X=1.435 $Y=1.28 $X2=0
+ $Y2=0
cc_183 N_GATE_N_M1005_g N_A_34_407#_c_342_n 0.0202871f $X=1.02 $Y=2.355 $X2=0
+ $Y2=0
cc_184 N_GATE_N_M1005_g N_A_34_407#_c_343_n 9.57066e-19 $X=1.02 $Y=2.355 $X2=0
+ $Y2=0
cc_185 N_GATE_N_c_183_n N_A_363_483#_c_409_n 2.78184e-19 $X=1.51 $Y=1.205 $X2=0
+ $Y2=0
cc_186 GATE_N N_A_363_483#_c_409_n 0.0327381f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_187 N_GATE_N_c_186_n N_A_363_483#_c_409_n 9.85879e-19 $X=1.6 $Y=0.4 $X2=0
+ $Y2=0
cc_188 N_GATE_N_c_183_n N_A_363_483#_c_411_n 0.004138f $X=1.51 $Y=1.205 $X2=0
+ $Y2=0
cc_189 N_GATE_N_M1005_g N_A_363_483#_c_419_n 0.00809552f $X=1.02 $Y=2.355 $X2=0
+ $Y2=0
cc_190 N_GATE_N_M1005_g N_VPWR_c_803_n 0.0176491f $X=1.02 $Y=2.355 $X2=0 $Y2=0
cc_191 N_GATE_N_M1005_g N_VPWR_c_810_n 0.00332367f $X=1.02 $Y=2.355 $X2=0 $Y2=0
cc_192 N_GATE_N_M1005_g N_VPWR_c_802_n 0.00387424f $X=1.02 $Y=2.355 $X2=0 $Y2=0
cc_193 N_GATE_N_c_180_n N_VGND_c_925_n 9.23465e-19 $X=1.02 $Y=1.205 $X2=0 $Y2=0
cc_194 GATE_N N_VGND_c_925_n 0.0354346f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_195 N_GATE_N_c_186_n N_VGND_c_925_n 0.00142946f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_196 GATE_N N_VGND_c_926_n 0.00103126f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_197 N_GATE_N_c_180_n N_VGND_c_932_n 0.00310205f $X=1.02 $Y=1.205 $X2=0 $Y2=0
cc_198 GATE_N N_VGND_c_932_n 0.0480349f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_199 N_GATE_N_c_186_n N_VGND_c_932_n 0.00590073f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_200 N_GATE_N_c_180_n N_VGND_c_936_n 0.0034947f $X=1.02 $Y=1.205 $X2=0 $Y2=0
cc_201 GATE_N N_VGND_c_936_n 0.0259334f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_202 N_GATE_N_c_186_n N_VGND_c_936_n 0.00775507f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_203 N_A_219_135#_c_239_n N_A_34_407#_c_332_n 0.0168908f $X=2.05 $Y=1.865
+ $X2=0 $Y2=0
cc_204 N_A_219_135#_c_229_n N_A_34_407#_c_332_n 0.0501107f $X=3.145 $Y=1.535
+ $X2=0 $Y2=0
cc_205 N_A_219_135#_c_230_n N_A_34_407#_c_332_n 0.00179158f $X=2.98 $Y=1.28
+ $X2=0 $Y2=0
cc_206 N_A_219_135#_c_231_n N_A_34_407#_c_332_n 0.00153131f $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_207 N_A_219_135#_c_232_n N_A_34_407#_c_332_n 0.00828664f $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_208 N_A_219_135#_M1010_g N_A_34_407#_M1019_g 0.041211f $X=2.265 $Y=0.445
+ $X2=0 $Y2=0
cc_209 N_A_219_135#_M1011_g N_A_34_407#_M1019_g 0.0501107f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_210 N_A_219_135#_c_230_n N_A_34_407#_M1019_g 0.0112929f $X=2.98 $Y=1.28 $X2=0
+ $Y2=0
cc_211 N_A_219_135#_c_231_n N_A_34_407#_M1019_g 9.52668e-19 $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_212 N_A_219_135#_c_232_n N_A_34_407#_M1019_g 0.00466642f $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_213 N_A_219_135#_c_233_n N_A_34_407#_M1019_g 0.00301844f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_214 N_A_219_135#_M1014_g N_A_34_407#_M1021_g 0.0182715f $X=2.155 $Y=2.735
+ $X2=0 $Y2=0
cc_215 N_A_219_135#_M1014_g N_A_34_407#_c_339_n 0.0168908f $X=2.155 $Y=2.735
+ $X2=0 $Y2=0
cc_216 N_A_219_135#_M1005_d N_A_34_407#_c_342_n 0.0187793f $X=1.095 $Y=2.035
+ $X2=0 $Y2=0
cc_217 N_A_219_135#_M1014_g N_A_34_407#_c_342_n 0.0131154f $X=2.155 $Y=2.735
+ $X2=0 $Y2=0
cc_218 N_A_219_135#_c_239_n N_A_34_407#_c_342_n 0.00118364f $X=2.05 $Y=1.865
+ $X2=0 $Y2=0
cc_219 N_A_219_135#_c_231_n N_A_34_407#_c_342_n 0.0911119f $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_220 N_A_219_135#_c_227_n N_A_34_407#_c_335_n 4.0375e-19 $X=3.31 $Y=1.61 $X2=0
+ $Y2=0
cc_221 N_A_219_135#_c_239_n N_A_34_407#_c_335_n 0.00191206f $X=2.05 $Y=1.865
+ $X2=0 $Y2=0
cc_222 N_A_219_135#_c_230_n N_A_34_407#_c_335_n 0.0210457f $X=2.98 $Y=1.28 $X2=0
+ $Y2=0
cc_223 N_A_219_135#_c_231_n N_A_34_407#_c_335_n 0.0216926f $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_224 N_A_219_135#_c_233_n N_A_34_407#_c_335_n 0.00622369f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_225 N_A_219_135#_M1006_g N_A_363_483#_M1000_g 0.0103849f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_226 N_A_219_135#_M1010_g N_A_363_483#_c_409_n 6.0147e-19 $X=2.265 $Y=0.445
+ $X2=0 $Y2=0
cc_227 N_A_219_135#_M1014_g N_A_363_483#_c_429_n 0.0100494f $X=2.155 $Y=2.735
+ $X2=0 $Y2=0
cc_228 N_A_219_135#_M1010_g N_A_363_483#_c_410_n 0.013217f $X=2.265 $Y=0.445
+ $X2=0 $Y2=0
cc_229 N_A_219_135#_M1011_g N_A_363_483#_c_410_n 0.0116055f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_230 N_A_219_135#_c_226_n N_A_363_483#_c_410_n 0.00199586f $X=3.67 $Y=1.61
+ $X2=0 $Y2=0
cc_231 N_A_219_135#_c_228_n N_A_363_483#_c_410_n 3.25562e-19 $X=2.105 $Y=1.345
+ $X2=0 $Y2=0
cc_232 N_A_219_135#_c_230_n N_A_363_483#_c_410_n 0.0333664f $X=2.98 $Y=1.28
+ $X2=0 $Y2=0
cc_233 N_A_219_135#_c_231_n N_A_363_483#_c_410_n 0.00295622f $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_234 N_A_219_135#_c_233_n N_A_363_483#_c_410_n 0.0201926f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_235 N_A_219_135#_c_234_n N_A_363_483#_c_410_n 0.00364392f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_236 N_A_219_135#_c_228_n N_A_363_483#_c_411_n 0.00131677f $X=2.105 $Y=1.345
+ $X2=0 $Y2=0
cc_237 N_A_219_135#_c_231_n N_A_363_483#_c_411_n 0.00970533f $X=2.035 $Y=1.36
+ $X2=0 $Y2=0
cc_238 N_A_219_135#_M1006_g N_A_363_483#_c_417_n 5.07755e-19 $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_239 N_A_219_135#_c_226_n N_A_363_483#_c_412_n 0.012793f $X=3.67 $Y=1.61 $X2=0
+ $Y2=0
cc_240 N_A_219_135#_M1006_g N_A_363_483#_c_412_n 0.00505762f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_241 N_A_219_135#_c_229_n N_A_363_483#_c_412_n 0.00559514f $X=3.145 $Y=1.535
+ $X2=0 $Y2=0
cc_242 N_A_219_135#_c_233_n N_A_363_483#_c_412_n 0.0229843f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_243 N_A_219_135#_M1014_g N_A_363_483#_c_419_n 0.00856725f $X=2.155 $Y=2.735
+ $X2=0 $Y2=0
cc_244 N_A_219_135#_c_227_n N_A_363_483#_c_420_n 0.0190483f $X=3.31 $Y=1.61
+ $X2=0 $Y2=0
cc_245 N_A_219_135#_M1006_g N_A_363_483#_c_420_n 0.0194394f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_246 N_A_219_135#_c_233_n N_A_363_483#_c_420_n 4.65285e-19 $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_247 N_A_219_135#_c_226_n N_A_363_483#_c_421_n 5.11953e-19 $X=3.67 $Y=1.61
+ $X2=0 $Y2=0
cc_248 N_A_219_135#_c_227_n N_A_363_483#_c_421_n 0.00234508f $X=3.31 $Y=1.61
+ $X2=0 $Y2=0
cc_249 N_A_219_135#_M1006_g N_A_363_483#_c_421_n 0.00198558f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_250 N_A_219_135#_c_233_n N_A_363_483#_c_421_n 0.0161089f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_251 N_A_219_135#_M1011_g N_A_363_483#_c_413_n 0.0039194f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_252 N_A_219_135#_c_226_n N_A_363_483#_c_413_n 0.00121446f $X=3.67 $Y=1.61
+ $X2=0 $Y2=0
cc_253 N_A_219_135#_c_233_n N_A_363_483#_c_413_n 0.0272403f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_254 N_A_219_135#_c_234_n N_A_363_483#_c_413_n 0.00559514f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_255 N_A_219_135#_c_226_n N_A_363_483#_c_414_n 0.00773562f $X=3.67 $Y=1.61
+ $X2=0 $Y2=0
cc_256 N_A_219_135#_c_234_n N_A_363_483#_c_414_n 0.00495669f $X=3.145 $Y=1.18
+ $X2=0 $Y2=0
cc_257 N_A_219_135#_M1011_g N_A_363_483#_c_415_n 0.022272f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_258 N_A_219_135#_c_226_n N_A_806_385#_M1007_g 0.0203684f $X=3.67 $Y=1.61
+ $X2=0 $Y2=0
cc_259 N_A_219_135#_M1006_g N_A_806_385#_c_542_n 2.96759e-19 $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_260 N_A_219_135#_M1006_g N_A_806_385#_c_543_n 0.060933f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_261 N_A_219_135#_c_226_n N_A_626_47#_c_669_n 0.00472317f $X=3.67 $Y=1.61
+ $X2=0 $Y2=0
cc_262 N_A_219_135#_M1006_g N_A_626_47#_c_669_n 0.00139168f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_263 N_A_219_135#_M1006_g N_A_626_47#_c_676_n 0.0207626f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_264 N_A_219_135#_M1006_g N_A_626_47#_c_677_n 0.012942f $X=3.745 $Y=2.625
+ $X2=0 $Y2=0
cc_265 N_A_219_135#_M1014_g N_VPWR_c_804_n 0.00501558f $X=2.155 $Y=2.735 $X2=0
+ $Y2=0
cc_266 N_A_219_135#_M1006_g N_VPWR_c_805_n 0.00118303f $X=3.745 $Y=2.625 $X2=0
+ $Y2=0
cc_267 N_A_219_135#_M1014_g N_VPWR_c_810_n 0.00390623f $X=2.155 $Y=2.735 $X2=0
+ $Y2=0
cc_268 N_A_219_135#_M1006_g N_VPWR_c_811_n 0.00326366f $X=3.745 $Y=2.625 $X2=0
+ $Y2=0
cc_269 N_A_219_135#_M1014_g N_VPWR_c_802_n 0.00700218f $X=2.155 $Y=2.735 $X2=0
+ $Y2=0
cc_270 N_A_219_135#_M1006_g N_VPWR_c_802_n 0.00307505f $X=3.745 $Y=2.625 $X2=0
+ $Y2=0
cc_271 N_A_219_135#_M1010_g N_VGND_c_926_n 0.00836588f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_272 N_A_219_135#_M1011_g N_VGND_c_926_n 0.00202732f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_273 N_A_219_135#_M1010_g N_VGND_c_932_n 0.00358332f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_274 N_A_219_135#_M1011_g N_VGND_c_933_n 0.00430895f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_275 N_A_219_135#_M1010_g N_VGND_c_936_n 0.00559922f $X=2.265 $Y=0.445 $X2=0
+ $Y2=0
cc_276 N_A_219_135#_M1011_g N_VGND_c_936_n 0.00624229f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_277 N_A_34_407#_M1021_g N_A_363_483#_M1000_g 0.0333102f $X=2.845 $Y=2.735
+ $X2=0 $Y2=0
cc_278 N_A_34_407#_M1021_g N_A_363_483#_c_429_n 0.0171269f $X=2.845 $Y=2.735
+ $X2=0 $Y2=0
cc_279 N_A_34_407#_c_340_n N_A_363_483#_c_429_n 0.00199975f $X=2.68 $Y=2.255
+ $X2=0 $Y2=0
cc_280 N_A_34_407#_c_342_n N_A_363_483#_c_429_n 0.0474548f $X=2.44 $Y=2.2 $X2=0
+ $Y2=0
cc_281 N_A_34_407#_M1019_g N_A_363_483#_c_410_n 0.0122077f $X=2.695 $Y=0.445
+ $X2=0 $Y2=0
cc_282 N_A_34_407#_c_340_n N_A_363_483#_c_417_n 0.0035069f $X=2.68 $Y=2.255
+ $X2=0 $Y2=0
cc_283 N_A_34_407#_c_342_n N_A_363_483#_c_417_n 0.00412351f $X=2.44 $Y=2.2 $X2=0
+ $Y2=0
cc_284 N_A_34_407#_c_332_n N_A_363_483#_c_412_n 0.00372265f $X=2.695 $Y=1.535
+ $X2=0 $Y2=0
cc_285 N_A_34_407#_c_335_n N_A_363_483#_c_412_n 0.00655943f $X=2.605 $Y=1.75
+ $X2=0 $Y2=0
cc_286 N_A_34_407#_M1021_g N_A_363_483#_c_419_n 8.62247e-19 $X=2.845 $Y=2.735
+ $X2=0 $Y2=0
cc_287 N_A_34_407#_c_342_n N_A_363_483#_c_419_n 0.0244295f $X=2.44 $Y=2.2 $X2=0
+ $Y2=0
cc_288 N_A_34_407#_c_339_n N_A_363_483#_c_420_n 0.00551314f $X=2.68 $Y=2.105
+ $X2=0 $Y2=0
cc_289 N_A_34_407#_c_340_n N_A_363_483#_c_420_n 0.0333102f $X=2.68 $Y=2.255
+ $X2=0 $Y2=0
cc_290 N_A_34_407#_c_339_n N_A_363_483#_c_421_n 0.00141359f $X=2.68 $Y=2.105
+ $X2=0 $Y2=0
cc_291 N_A_34_407#_c_340_n N_A_363_483#_c_421_n 0.0010274f $X=2.68 $Y=2.255
+ $X2=0 $Y2=0
cc_292 N_A_34_407#_c_342_n N_A_363_483#_c_421_n 0.00835384f $X=2.44 $Y=2.2 $X2=0
+ $Y2=0
cc_293 N_A_34_407#_c_335_n N_A_363_483#_c_421_n 0.0136518f $X=2.605 $Y=1.75
+ $X2=0 $Y2=0
cc_294 N_A_34_407#_c_342_n N_VPWR_M1012_d 0.0055019f $X=2.44 $Y=2.2 $X2=-0.19
+ $Y2=-0.245
cc_295 N_A_34_407#_c_342_n N_VPWR_c_803_n 0.0218003f $X=2.44 $Y=2.2 $X2=0 $Y2=0
cc_296 N_A_34_407#_c_343_n N_VPWR_c_803_n 0.00945783f $X=0.295 $Y=2.18 $X2=0
+ $Y2=0
cc_297 N_A_34_407#_M1021_g N_VPWR_c_804_n 0.00670485f $X=2.845 $Y=2.735 $X2=0
+ $Y2=0
cc_298 N_A_34_407#_M1021_g N_VPWR_c_811_n 0.00400666f $X=2.845 $Y=2.735 $X2=0
+ $Y2=0
cc_299 N_A_34_407#_M1021_g N_VPWR_c_802_n 0.00599185f $X=2.845 $Y=2.735 $X2=0
+ $Y2=0
cc_300 N_A_34_407#_c_343_n N_VPWR_c_802_n 0.0106715f $X=0.295 $Y=2.18 $X2=0
+ $Y2=0
cc_301 N_A_34_407#_c_343_n N_VPWR_c_815_n 0.00708045f $X=0.295 $Y=2.18 $X2=0
+ $Y2=0
cc_302 N_A_34_407#_M1019_g N_VGND_c_926_n 0.00970404f $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_303 N_A_34_407#_M1019_g N_VGND_c_933_n 0.00358332f $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_304 N_A_34_407#_M1019_g N_VGND_c_936_n 0.00410582f $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_305 N_A_34_407#_c_336_n N_VGND_c_936_n 0.0112326f $X=0.375 $Y=0.87 $X2=0
+ $Y2=0
cc_306 N_A_34_407#_c_336_n N_VGND_c_937_n 0.00620969f $X=0.375 $Y=0.87 $X2=0
+ $Y2=0
cc_307 N_A_363_483#_c_412_n N_A_806_385#_M1007_g 0.00226844f $X=3.495 $Y=1.925
+ $X2=0 $Y2=0
cc_308 N_A_363_483#_c_413_n N_A_806_385#_M1007_g 5.70324e-19 $X=3.595 $Y=0.76
+ $X2=0 $Y2=0
cc_309 N_A_363_483#_c_414_n N_A_806_385#_M1007_g 0.0203599f $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_310 N_A_363_483#_c_415_n N_A_806_385#_M1007_g 0.0194147f $X=3.685 $Y=0.765
+ $X2=0 $Y2=0
cc_311 N_A_363_483#_c_410_n N_A_626_47#_c_682_n 0.0152345f $X=3.41 $Y=0.76 $X2=0
+ $Y2=0
cc_312 N_A_363_483#_c_413_n N_A_626_47#_c_682_n 0.0213138f $X=3.595 $Y=0.76
+ $X2=0 $Y2=0
cc_313 N_A_363_483#_c_414_n N_A_626_47#_c_682_n 0.00292019f $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_314 N_A_363_483#_c_415_n N_A_626_47#_c_682_n 0.00963915f $X=3.685 $Y=0.765
+ $X2=0 $Y2=0
cc_315 N_A_363_483#_c_412_n N_A_626_47#_c_669_n 0.025822f $X=3.495 $Y=1.925
+ $X2=0 $Y2=0
cc_316 N_A_363_483#_c_413_n N_A_626_47#_c_669_n 6.63044e-19 $X=3.595 $Y=0.76
+ $X2=0 $Y2=0
cc_317 N_A_363_483#_c_414_n N_A_626_47#_c_669_n 0.00121915f $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_318 N_A_363_483#_c_412_n N_A_626_47#_c_670_n 0.00787314f $X=3.495 $Y=1.925
+ $X2=0 $Y2=0
cc_319 N_A_363_483#_c_413_n N_A_626_47#_c_670_n 0.0322179f $X=3.595 $Y=0.76
+ $X2=0 $Y2=0
cc_320 N_A_363_483#_c_414_n N_A_626_47#_c_670_n 0.00200461f $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_321 N_A_363_483#_c_415_n N_A_626_47#_c_670_n 0.00384121f $X=3.685 $Y=0.765
+ $X2=0 $Y2=0
cc_322 N_A_363_483#_M1000_g N_A_626_47#_c_676_n 0.00217414f $X=3.205 $Y=2.735
+ $X2=0 $Y2=0
cc_323 N_A_363_483#_c_417_n N_A_626_47#_c_676_n 0.00286794f $X=3.06 $Y=2.455
+ $X2=0 $Y2=0
cc_324 N_A_363_483#_c_420_n N_A_626_47#_c_676_n 0.00347058f $X=3.295 $Y=2.09
+ $X2=0 $Y2=0
cc_325 N_A_363_483#_c_421_n N_A_626_47#_c_676_n 0.0225809f $X=3.495 $Y=2.075
+ $X2=0 $Y2=0
cc_326 N_A_363_483#_M1000_g N_A_626_47#_c_677_n 4.59486e-19 $X=3.205 $Y=2.735
+ $X2=0 $Y2=0
cc_327 N_A_363_483#_c_417_n N_A_626_47#_c_677_n 0.00394334f $X=3.06 $Y=2.455
+ $X2=0 $Y2=0
cc_328 N_A_363_483#_c_412_n N_A_626_47#_c_677_n 0.0122994f $X=3.495 $Y=1.925
+ $X2=0 $Y2=0
cc_329 N_A_363_483#_c_420_n N_A_626_47#_c_677_n 3.73897e-19 $X=3.295 $Y=2.09
+ $X2=0 $Y2=0
cc_330 N_A_363_483#_c_421_n N_A_626_47#_c_677_n 0.0227983f $X=3.495 $Y=2.075
+ $X2=0 $Y2=0
cc_331 N_A_363_483#_c_429_n N_VPWR_M1014_d 0.0110532f $X=2.975 $Y=2.545 $X2=0
+ $Y2=0
cc_332 N_A_363_483#_c_429_n N_VPWR_c_804_n 0.023171f $X=2.975 $Y=2.545 $X2=0
+ $Y2=0
cc_333 N_A_363_483#_c_419_n N_VPWR_c_804_n 0.0146934f $X=1.94 $Y=2.57 $X2=0
+ $Y2=0
cc_334 N_A_363_483#_c_429_n N_VPWR_c_810_n 0.00322361f $X=2.975 $Y=2.545 $X2=0
+ $Y2=0
cc_335 N_A_363_483#_c_419_n N_VPWR_c_810_n 0.0232661f $X=1.94 $Y=2.57 $X2=0
+ $Y2=0
cc_336 N_A_363_483#_M1000_g N_VPWR_c_811_n 0.00531047f $X=3.205 $Y=2.735 $X2=0
+ $Y2=0
cc_337 N_A_363_483#_c_429_n N_VPWR_c_811_n 0.00587385f $X=2.975 $Y=2.545 $X2=0
+ $Y2=0
cc_338 N_A_363_483#_M1000_g N_VPWR_c_802_n 0.0109378f $X=3.205 $Y=2.735 $X2=0
+ $Y2=0
cc_339 N_A_363_483#_c_429_n N_VPWR_c_802_n 0.0195693f $X=2.975 $Y=2.545 $X2=0
+ $Y2=0
cc_340 N_A_363_483#_c_419_n N_VPWR_c_802_n 0.0126112f $X=1.94 $Y=2.57 $X2=0
+ $Y2=0
cc_341 N_A_363_483#_c_429_n A_584_483# 0.0018404f $X=2.975 $Y=2.545 $X2=-0.19
+ $Y2=-0.245
cc_342 N_A_363_483#_c_410_n N_VGND_c_926_n 0.02032f $X=3.41 $Y=0.76 $X2=0 $Y2=0
cc_343 N_A_363_483#_c_409_n N_VGND_c_932_n 0.0108936f $X=2.05 $Y=0.45 $X2=0
+ $Y2=0
cc_344 N_A_363_483#_c_410_n N_VGND_c_932_n 0.0027696f $X=3.41 $Y=0.76 $X2=0
+ $Y2=0
cc_345 N_A_363_483#_c_410_n N_VGND_c_933_n 0.00820211f $X=3.41 $Y=0.76 $X2=0
+ $Y2=0
cc_346 N_A_363_483#_c_415_n N_VGND_c_933_n 0.00362032f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_347 N_A_363_483#_M1010_s N_VGND_c_936_n 0.0031135f $X=1.925 $Y=0.235 $X2=0
+ $Y2=0
cc_348 N_A_363_483#_c_409_n N_VGND_c_936_n 0.0071561f $X=2.05 $Y=0.45 $X2=0
+ $Y2=0
cc_349 N_A_363_483#_c_410_n N_VGND_c_936_n 0.0192975f $X=3.41 $Y=0.76 $X2=0
+ $Y2=0
cc_350 N_A_363_483#_c_415_n N_VGND_c_936_n 0.00591116f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_351 N_A_806_385#_M1007_g N_A_626_47#_M1017_g 0.0289199f $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_352 N_A_806_385#_c_527_n N_A_626_47#_M1017_g 0.00548432f $X=5.105 $Y=1.925
+ $X2=0 $Y2=0
cc_353 N_A_806_385#_c_535_n N_A_626_47#_M1017_g 0.00280949f $X=4.875 $Y=0.42
+ $X2=0 $Y2=0
cc_354 N_A_806_385#_M1009_g N_A_626_47#_M1020_g 0.00471091f $X=4.105 $Y=2.625
+ $X2=0 $Y2=0
cc_355 N_A_806_385#_M1007_g N_A_626_47#_M1020_g 0.00753469f $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_356 N_A_806_385#_c_542_n N_A_626_47#_M1020_g 0.0196451f $X=4.925 $Y=2.09
+ $X2=0 $Y2=0
cc_357 N_A_806_385#_c_543_n N_A_626_47#_M1020_g 0.00792564f $X=4.195 $Y=2.09
+ $X2=0 $Y2=0
cc_358 N_A_806_385#_c_544_n N_A_626_47#_M1020_g 0.0157806f $X=5.09 $Y=2.91 $X2=0
+ $Y2=0
cc_359 N_A_806_385#_c_546_n N_A_626_47#_M1020_g 0.00254439f $X=5.09 $Y=2.03
+ $X2=0 $Y2=0
cc_360 N_A_806_385#_M1007_g N_A_626_47#_c_682_n 0.00640465f $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_361 N_A_806_385#_M1007_g N_A_626_47#_c_669_n 0.0162564f $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_362 N_A_806_385#_c_542_n N_A_626_47#_c_669_n 0.00152455f $X=4.925 $Y=2.09
+ $X2=0 $Y2=0
cc_363 N_A_806_385#_c_543_n N_A_626_47#_c_669_n 0.00143597f $X=4.195 $Y=2.09
+ $X2=0 $Y2=0
cc_364 N_A_806_385#_M1007_g N_A_626_47#_c_670_n 0.0183825f $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_365 N_A_806_385#_M1007_g N_A_626_47#_c_671_n 0.00995838f $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_366 N_A_806_385#_c_542_n N_A_626_47#_c_671_n 0.0165143f $X=4.925 $Y=2.09
+ $X2=0 $Y2=0
cc_367 N_A_806_385#_c_543_n N_A_626_47#_c_671_n 0.00266472f $X=4.195 $Y=2.09
+ $X2=0 $Y2=0
cc_368 N_A_806_385#_M1009_g N_A_626_47#_c_676_n 0.00460688f $X=4.105 $Y=2.625
+ $X2=0 $Y2=0
cc_369 N_A_806_385#_M1007_g N_A_626_47#_c_677_n 0.00380466f $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_370 N_A_806_385#_c_542_n N_A_626_47#_c_677_n 0.0262102f $X=4.925 $Y=2.09
+ $X2=0 $Y2=0
cc_371 N_A_806_385#_c_543_n N_A_626_47#_c_677_n 0.00345817f $X=4.195 $Y=2.09
+ $X2=0 $Y2=0
cc_372 N_A_806_385#_M1007_g N_A_626_47#_c_672_n 7.09717e-19 $X=4.135 $Y=0.445
+ $X2=0 $Y2=0
cc_373 N_A_806_385#_c_542_n N_A_626_47#_c_672_n 0.0108164f $X=4.925 $Y=2.09
+ $X2=0 $Y2=0
cc_374 N_A_806_385#_c_527_n N_A_626_47#_c_672_n 0.0244628f $X=5.105 $Y=1.925
+ $X2=0 $Y2=0
cc_375 N_A_806_385#_c_535_n N_A_626_47#_c_672_n 0.00592417f $X=4.875 $Y=0.42
+ $X2=0 $Y2=0
cc_376 N_A_806_385#_M1004_g N_A_626_47#_c_673_n 0.00215537f $X=5.685 $Y=1.015
+ $X2=0 $Y2=0
cc_377 N_A_806_385#_c_542_n N_A_626_47#_c_673_n 0.00121842f $X=4.925 $Y=2.09
+ $X2=0 $Y2=0
cc_378 N_A_806_385#_c_527_n N_A_626_47#_c_673_n 0.0164577f $X=5.105 $Y=1.925
+ $X2=0 $Y2=0
cc_379 N_A_806_385#_c_535_n N_A_626_47#_c_673_n 0.00564324f $X=4.875 $Y=0.42
+ $X2=0 $Y2=0
cc_380 N_A_806_385#_M1016_g N_A_1069_161#_M1001_g 0.0124349f $X=5.97 $Y=2.145
+ $X2=0 $Y2=0
cc_381 N_A_806_385#_c_531_n N_A_1069_161#_c_752_n 0.00337097f $X=6.445 $Y=1.16
+ $X2=0 $Y2=0
cc_382 N_A_806_385#_c_533_n N_A_1069_161#_c_752_n 0.0187587f $X=7.295 $Y=0.74
+ $X2=0 $Y2=0
cc_383 N_A_806_385#_c_534_n N_A_1069_161#_c_752_n 0.0034275f $X=7.46 $Y=1.35
+ $X2=0 $Y2=0
cc_384 N_A_806_385#_c_537_n N_A_1069_161#_c_752_n 0.00604206f $X=7.685 $Y=1.35
+ $X2=0 $Y2=0
cc_385 N_A_806_385#_M1004_g N_A_1069_161#_c_753_n 0.00597696f $X=5.685 $Y=1.015
+ $X2=0 $Y2=0
cc_386 N_A_806_385#_c_528_n N_A_1069_161#_c_753_n 0.0154284f $X=5.725 $Y=0.465
+ $X2=0 $Y2=0
cc_387 N_A_806_385#_c_532_n N_A_1069_161#_c_753_n 0.0078912f $X=5.895 $Y=1.16
+ $X2=0 $Y2=0
cc_388 N_A_806_385#_c_535_n N_A_1069_161#_c_753_n 0.0433966f $X=4.875 $Y=0.42
+ $X2=0 $Y2=0
cc_389 N_A_806_385#_M1016_g N_A_1069_161#_c_758_n 0.0149156f $X=5.97 $Y=2.145
+ $X2=0 $Y2=0
cc_390 N_A_806_385#_c_544_n N_A_1069_161#_c_758_n 0.0115575f $X=5.09 $Y=2.91
+ $X2=0 $Y2=0
cc_391 N_A_806_385#_c_527_n N_A_1069_161#_c_758_n 0.0126854f $X=5.105 $Y=1.925
+ $X2=0 $Y2=0
cc_392 N_A_806_385#_c_546_n N_A_1069_161#_c_758_n 0.0176777f $X=5.09 $Y=2.03
+ $X2=0 $Y2=0
cc_393 N_A_806_385#_M1016_g N_A_1069_161#_c_754_n 0.00361542f $X=5.97 $Y=2.145
+ $X2=0 $Y2=0
cc_394 N_A_806_385#_c_526_n N_A_1069_161#_c_754_n 0.0177845f $X=5.97 $Y=1.41
+ $X2=0 $Y2=0
cc_395 N_A_806_385#_c_527_n N_A_1069_161#_c_754_n 0.0167761f $X=5.105 $Y=1.925
+ $X2=0 $Y2=0
cc_396 N_A_806_385#_c_531_n N_A_1069_161#_c_754_n 0.00195992f $X=6.445 $Y=1.16
+ $X2=0 $Y2=0
cc_397 N_A_806_385#_c_532_n N_A_1069_161#_c_754_n 0.0149974f $X=5.895 $Y=1.16
+ $X2=0 $Y2=0
cc_398 N_A_806_385#_M1016_g N_A_1069_161#_c_755_n 0.00888533f $X=5.97 $Y=2.145
+ $X2=0 $Y2=0
cc_399 N_A_806_385#_c_526_n N_A_1069_161#_c_755_n 0.00242166f $X=5.97 $Y=1.41
+ $X2=0 $Y2=0
cc_400 N_A_806_385#_c_531_n N_A_1069_161#_c_755_n 0.0529146f $X=6.445 $Y=1.16
+ $X2=0 $Y2=0
cc_401 N_A_806_385#_c_526_n N_A_1069_161#_c_756_n 0.0194215f $X=5.97 $Y=1.41
+ $X2=0 $Y2=0
cc_402 N_A_806_385#_c_531_n N_A_1069_161#_c_756_n 0.00892394f $X=6.445 $Y=1.16
+ $X2=0 $Y2=0
cc_403 N_A_806_385#_c_542_n N_VPWR_M1009_d 0.00689532f $X=4.925 $Y=2.09 $X2=0
+ $Y2=0
cc_404 N_A_806_385#_M1009_g N_VPWR_c_805_n 0.0114277f $X=4.105 $Y=2.625 $X2=0
+ $Y2=0
cc_405 N_A_806_385#_c_542_n N_VPWR_c_805_n 0.0470421f $X=4.925 $Y=2.09 $X2=0
+ $Y2=0
cc_406 N_A_806_385#_c_543_n N_VPWR_c_805_n 0.00413786f $X=4.195 $Y=2.09 $X2=0
+ $Y2=0
cc_407 N_A_806_385#_M1016_g N_VPWR_c_806_n 0.00481843f $X=5.97 $Y=2.145 $X2=0
+ $Y2=0
cc_408 N_A_806_385#_M1013_g N_VPWR_c_807_n 0.0259605f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_409 N_A_806_385#_c_534_n N_VPWR_c_807_n 0.0184481f $X=7.46 $Y=1.35 $X2=0
+ $Y2=0
cc_410 N_A_806_385#_c_537_n N_VPWR_c_807_n 0.00224381f $X=7.685 $Y=1.35 $X2=0
+ $Y2=0
cc_411 N_A_806_385#_M1016_g N_VPWR_c_808_n 0.00308674f $X=5.97 $Y=2.145 $X2=0
+ $Y2=0
cc_412 N_A_806_385#_c_544_n N_VPWR_c_808_n 0.0199714f $X=5.09 $Y=2.91 $X2=0
+ $Y2=0
cc_413 N_A_806_385#_M1009_g N_VPWR_c_811_n 0.00407914f $X=4.105 $Y=2.625 $X2=0
+ $Y2=0
cc_414 N_A_806_385#_M1013_g N_VPWR_c_813_n 0.00486043f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_A_806_385#_M1009_g N_VPWR_c_802_n 0.00425776f $X=4.105 $Y=2.625 $X2=0
+ $Y2=0
cc_416 N_A_806_385#_M1016_g N_VPWR_c_802_n 0.00407903f $X=5.97 $Y=2.145 $X2=0
+ $Y2=0
cc_417 N_A_806_385#_M1013_g N_VPWR_c_802_n 0.00917987f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A_806_385#_c_544_n N_VPWR_c_802_n 0.0120489f $X=5.09 $Y=2.91 $X2=0
+ $Y2=0
cc_419 N_A_806_385#_c_533_n N_Q_N_M1018_d 0.00670674f $X=7.295 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_420 N_A_806_385#_c_524_n N_Q_N_c_890_n 7.23838e-19 $X=7.685 $Y=1.185 $X2=0
+ $Y2=0
cc_421 N_A_806_385#_M1013_g N_Q_N_c_890_n 0.00801365f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_806_385#_c_531_n N_Q_N_c_890_n 0.00732422f $X=6.445 $Y=1.16 $X2=0
+ $Y2=0
cc_423 N_A_806_385#_c_533_n N_Q_N_c_890_n 0.0228472f $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_424 N_A_806_385#_c_534_n N_Q_N_c_890_n 0.042035f $X=7.46 $Y=1.35 $X2=0 $Y2=0
cc_425 N_A_806_385#_c_537_n N_Q_N_c_890_n 0.00313813f $X=7.685 $Y=1.35 $X2=0
+ $Y2=0
cc_426 N_A_806_385#_M1013_g N_Q_N_c_893_n 0.0027362f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_427 N_A_806_385#_c_524_n N_Q_c_914_n 0.0298739f $X=7.685 $Y=1.185 $X2=0 $Y2=0
cc_428 N_A_806_385#_c_534_n N_Q_c_914_n 0.0415788f $X=7.46 $Y=1.35 $X2=0 $Y2=0
cc_429 N_A_806_385#_c_530_n N_VGND_M1004_d 0.0040577f $X=5.81 $Y=1.075 $X2=0
+ $Y2=0
cc_430 N_A_806_385#_c_531_n N_VGND_M1004_d 0.0204357f $X=6.445 $Y=1.16 $X2=0
+ $Y2=0
cc_431 N_A_806_385#_c_634_p N_VGND_M1004_d 0.00439601f $X=6.53 $Y=1.075 $X2=0
+ $Y2=0
cc_432 N_A_806_385#_c_635_p N_VGND_M1004_d 0.00501674f $X=6.615 $Y=0.74 $X2=0
+ $Y2=0
cc_433 N_A_806_385#_c_533_n N_VGND_M1003_s 0.00302014f $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_434 N_A_806_385#_c_534_n N_VGND_M1003_s 8.42155e-19 $X=7.46 $Y=1.35 $X2=0
+ $Y2=0
cc_435 N_A_806_385#_M1007_g N_VGND_c_927_n 0.0087931f $X=4.135 $Y=0.445 $X2=0
+ $Y2=0
cc_436 N_A_806_385#_c_535_n N_VGND_c_927_n 0.0320398f $X=4.875 $Y=0.42 $X2=0
+ $Y2=0
cc_437 N_A_806_385#_M1004_g N_VGND_c_928_n 0.00119168f $X=5.685 $Y=1.015 $X2=0
+ $Y2=0
cc_438 N_A_806_385#_c_529_n N_VGND_c_928_n 0.034172f $X=5.81 $Y=0.675 $X2=0
+ $Y2=0
cc_439 N_A_806_385#_c_530_n N_VGND_c_928_n 0.0171101f $X=5.81 $Y=1.075 $X2=0
+ $Y2=0
cc_440 N_A_806_385#_c_531_n N_VGND_c_928_n 0.0169226f $X=6.445 $Y=1.16 $X2=0
+ $Y2=0
cc_441 N_A_806_385#_c_634_p N_VGND_c_928_n 0.00586784f $X=6.53 $Y=1.075 $X2=0
+ $Y2=0
cc_442 N_A_806_385#_c_635_p N_VGND_c_928_n 0.0140305f $X=6.615 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_806_385#_c_536_n N_VGND_c_928_n 0.00751863f $X=5.74 $Y=0.51 $X2=0
+ $Y2=0
cc_444 N_A_806_385#_c_524_n N_VGND_c_929_n 0.00959844f $X=7.685 $Y=1.185 $X2=0
+ $Y2=0
cc_445 N_A_806_385#_c_533_n N_VGND_c_929_n 0.0222084f $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_446 N_A_806_385#_c_537_n N_VGND_c_929_n 7.79959e-19 $X=7.685 $Y=1.35 $X2=0
+ $Y2=0
cc_447 N_A_806_385#_c_528_n N_VGND_c_930_n 0.0363774f $X=5.725 $Y=0.465 $X2=0
+ $Y2=0
cc_448 N_A_806_385#_c_529_n N_VGND_c_930_n 0.0121867f $X=5.81 $Y=0.675 $X2=0
+ $Y2=0
cc_449 N_A_806_385#_c_535_n N_VGND_c_930_n 0.0292773f $X=4.875 $Y=0.42 $X2=0
+ $Y2=0
cc_450 N_A_806_385#_c_536_n N_VGND_c_930_n 0.00193865f $X=5.74 $Y=0.51 $X2=0
+ $Y2=0
cc_451 N_A_806_385#_M1007_g N_VGND_c_933_n 0.00495961f $X=4.135 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_806_385#_c_533_n N_VGND_c_934_n 0.0107873f $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_453 N_A_806_385#_c_635_p N_VGND_c_934_n 0.00299978f $X=6.615 $Y=0.74 $X2=0
+ $Y2=0
cc_454 N_A_806_385#_c_524_n N_VGND_c_935_n 0.00486043f $X=7.685 $Y=1.185 $X2=0
+ $Y2=0
cc_455 N_A_806_385#_M1017_d N_VGND_c_936_n 0.00336915f $X=4.735 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_A_806_385#_M1007_g N_VGND_c_936_n 0.00912493f $X=4.135 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_806_385#_c_524_n N_VGND_c_936_n 0.00917987f $X=7.685 $Y=1.185 $X2=0
+ $Y2=0
cc_458 N_A_806_385#_c_528_n N_VGND_c_936_n 0.0203371f $X=5.725 $Y=0.465 $X2=0
+ $Y2=0
cc_459 N_A_806_385#_c_529_n N_VGND_c_936_n 0.00660921f $X=5.81 $Y=0.675 $X2=0
+ $Y2=0
cc_460 N_A_806_385#_c_533_n N_VGND_c_936_n 0.0208605f $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_461 N_A_806_385#_c_635_p N_VGND_c_936_n 0.00504936f $X=6.615 $Y=0.74 $X2=0
+ $Y2=0
cc_462 N_A_806_385#_c_535_n N_VGND_c_936_n 0.0164453f $X=4.875 $Y=0.42 $X2=0
+ $Y2=0
cc_463 N_A_806_385#_c_536_n N_VGND_c_936_n 3.21278e-19 $X=5.74 $Y=0.51 $X2=0
+ $Y2=0
cc_464 N_A_626_47#_M1020_g N_A_1069_161#_c_758_n 0.00131064f $X=4.875 $Y=2.445
+ $X2=0 $Y2=0
cc_465 N_A_626_47#_c_676_n N_VPWR_c_804_n 0.00371252f $X=3.53 $Y=2.56 $X2=0
+ $Y2=0
cc_466 N_A_626_47#_M1020_g N_VPWR_c_805_n 0.00483061f $X=4.875 $Y=2.445 $X2=0
+ $Y2=0
cc_467 N_A_626_47#_c_676_n N_VPWR_c_805_n 0.0295534f $X=3.53 $Y=2.56 $X2=0 $Y2=0
cc_468 N_A_626_47#_M1020_g N_VPWR_c_808_n 0.00529818f $X=4.875 $Y=2.445 $X2=0
+ $Y2=0
cc_469 N_A_626_47#_c_676_n N_VPWR_c_811_n 0.0278151f $X=3.53 $Y=2.56 $X2=0 $Y2=0
cc_470 N_A_626_47#_M1020_g N_VPWR_c_802_n 0.0121231f $X=4.875 $Y=2.445 $X2=0
+ $Y2=0
cc_471 N_A_626_47#_c_676_n N_VPWR_c_802_n 0.0238643f $X=3.53 $Y=2.56 $X2=0 $Y2=0
cc_472 N_A_626_47#_c_676_n A_764_483# 0.0026185f $X=3.53 $Y=2.56 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_626_47#_M1017_g N_VGND_c_927_n 0.0159552f $X=4.66 $Y=0.655 $X2=0
+ $Y2=0
cc_474 N_A_626_47#_c_682_n N_VGND_c_927_n 0.0172261f $X=3.95 $Y=0.38 $X2=0 $Y2=0
cc_475 N_A_626_47#_c_670_n N_VGND_c_927_n 0.0455282f $X=4.035 $Y=1.275 $X2=0
+ $Y2=0
cc_476 N_A_626_47#_c_671_n N_VGND_c_927_n 0.0238449f $X=4.585 $Y=1.36 $X2=0
+ $Y2=0
cc_477 N_A_626_47#_c_672_n N_VGND_c_927_n 9.95851e-19 $X=4.715 $Y=1.36 $X2=0
+ $Y2=0
cc_478 N_A_626_47#_M1017_g N_VGND_c_930_n 0.00525069f $X=4.66 $Y=0.655 $X2=0
+ $Y2=0
cc_479 N_A_626_47#_c_682_n N_VGND_c_933_n 0.049717f $X=3.95 $Y=0.38 $X2=0 $Y2=0
cc_480 N_A_626_47#_M1011_d N_VGND_c_936_n 0.00328567f $X=3.13 $Y=0.235 $X2=0
+ $Y2=0
cc_481 N_A_626_47#_M1017_g N_VGND_c_936_n 0.0101648f $X=4.66 $Y=0.655 $X2=0
+ $Y2=0
cc_482 N_A_626_47#_c_682_n N_VGND_c_936_n 0.0348026f $X=3.95 $Y=0.38 $X2=0 $Y2=0
cc_483 N_A_626_47#_c_682_n A_734_47# 0.00834986f $X=3.95 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_484 N_A_626_47#_c_670_n A_734_47# 0.00213563f $X=4.035 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_485 N_A_1069_161#_M1001_g N_VPWR_c_806_n 0.00733792f $X=6.46 $Y=2.455 $X2=0
+ $Y2=0
cc_486 N_A_1069_161#_c_758_n N_VPWR_c_806_n 0.0270402f $X=5.755 $Y=1.97 $X2=0
+ $Y2=0
cc_487 N_A_1069_161#_c_755_n N_VPWR_c_806_n 0.02193f $X=6.45 $Y=1.5 $X2=0 $Y2=0
cc_488 N_A_1069_161#_c_756_n N_VPWR_c_806_n 0.00154585f $X=6.735 $Y=1.5 $X2=0
+ $Y2=0
cc_489 N_A_1069_161#_M1001_g N_VPWR_c_812_n 0.00575161f $X=6.46 $Y=2.455 $X2=0
+ $Y2=0
cc_490 N_A_1069_161#_M1001_g N_VPWR_c_802_n 0.0132031f $X=6.46 $Y=2.455 $X2=0
+ $Y2=0
cc_491 N_A_1069_161#_c_758_n N_VPWR_c_802_n 0.0127828f $X=5.755 $Y=1.97 $X2=0
+ $Y2=0
cc_492 N_A_1069_161#_M1001_g N_Q_N_c_890_n 0.00474981f $X=6.46 $Y=2.455 $X2=0
+ $Y2=0
cc_493 N_A_1069_161#_c_752_n N_Q_N_c_890_n 0.00844137f $X=6.735 $Y=1.335 $X2=0
+ $Y2=0
cc_494 N_A_1069_161#_c_755_n N_Q_N_c_890_n 0.0174394f $X=6.45 $Y=1.5 $X2=0 $Y2=0
cc_495 N_A_1069_161#_c_756_n N_Q_N_c_890_n 0.0151361f $X=6.735 $Y=1.5 $X2=0
+ $Y2=0
cc_496 N_A_1069_161#_M1001_g N_Q_N_c_893_n 0.0035417f $X=6.46 $Y=2.455 $X2=0
+ $Y2=0
cc_497 N_A_1069_161#_c_755_n N_Q_N_c_893_n 0.00196937f $X=6.45 $Y=1.5 $X2=0
+ $Y2=0
cc_498 N_A_1069_161#_c_756_n N_Q_N_c_893_n 0.00889361f $X=6.735 $Y=1.5 $X2=0
+ $Y2=0
cc_499 N_A_1069_161#_c_752_n N_VGND_c_928_n 0.0120719f $X=6.735 $Y=1.335 $X2=0
+ $Y2=0
cc_500 N_A_1069_161#_c_752_n N_VGND_c_929_n 0.0060671f $X=6.735 $Y=1.335 $X2=0
+ $Y2=0
cc_501 N_A_1069_161#_c_752_n N_VGND_c_934_n 0.00436648f $X=6.735 $Y=1.335 $X2=0
+ $Y2=0
cc_502 N_A_1069_161#_c_752_n N_VGND_c_936_n 0.0054106f $X=6.735 $Y=1.335 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_802_n N_Q_N_M1001_d 0.00403632f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_504 N_VPWR_c_812_n Q_N 0.037887f $X=7.305 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_c_802_n Q_N 0.0207165f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_c_806_n N_Q_N_c_893_n 0.00126691f $X=6.21 $Y=1.97 $X2=0 $Y2=0
cc_507 N_VPWR_c_807_n N_Q_N_c_893_n 0.104549f $X=7.47 $Y=1.98 $X2=0 $Y2=0
cc_508 N_VPWR_c_802_n N_Q_M1013_d 0.00371702f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_509 N_VPWR_c_807_n N_Q_c_914_n 0.0480407f $X=7.47 $Y=1.98 $X2=0 $Y2=0
cc_510 N_VPWR_c_813_n N_Q_c_914_n 0.0178111f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_511 N_VPWR_c_802_n N_Q_c_914_n 0.0100304f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_512 N_Q_c_914_n N_VGND_c_935_n 0.0178111f $X=7.9 $Y=0.42 $X2=0 $Y2=0
cc_513 N_Q_M1003_d N_VGND_c_936_n 0.00371702f $X=7.76 $Y=0.235 $X2=0 $Y2=0
cc_514 N_Q_c_914_n N_VGND_c_936_n 0.0100304f $X=7.9 $Y=0.42 $X2=0 $Y2=0
cc_515 N_VGND_c_936_n A_554_47# 0.00256433f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_516 N_VGND_c_936_n A_734_47# 0.00315661f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
