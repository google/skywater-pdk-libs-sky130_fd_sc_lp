* File: sky130_fd_sc_lp__o2111a_1.spice
* Created: Wed Sep  2 10:12:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111a_1.pex.spice"
.subckt sky130_fd_sc_lp__o2111a_1  VNB VPB D1 C1 B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 A_337_49# N_D1_M1005_g N_A_80_21#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1002 A_409_49# N_C1_M1002_g A_337_49# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75000.6 SB=75001.9
+ A=0.126 P=1.98 MULT=1
MM1004 N_A_517_49#_M1004_d N_B1_M1004_g A_409_49# VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1638 PD=1.46 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75001.1
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_517_49#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_517_49#_M1009_d N_A1_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_VPWR_M1011_d N_A_80_21#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.57645 AS=0.3339 PD=2.175 PS=3.05 NRD=12.4898 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1010 N_A_80_21#_M1010_d N_D1_M1010_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.57645 PD=1.54 PS=2.175 NRD=0 NRS=37.1148 M=1 R=8.4 SA=75001.3
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_C1_M1006_g N_A_80_21#_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4347 AS=0.1764 PD=1.95 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1001 N_A_80_21#_M1001_d N_B1_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.4347 PD=1.65 PS=1.95 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 A_685_367# N_A2_M1007_g N_A_80_21#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.2457 PD=1.47 PS=1.65 NRD=7.8012 NRS=6.2449 M=1 R=8.4 SA=75003.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_685_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75003.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o2111a_1.pxi.spice"
*
.ends
*
*
