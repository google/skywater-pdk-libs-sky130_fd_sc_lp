* File: sky130_fd_sc_lp__ebufn_4.pxi.spice
* Created: Fri Aug 28 10:31:49 2020
* 
x_PM_SKY130_FD_SC_LP__EBUFN_4%A_84_21# N_A_84_21#_M1019_d N_A_84_21#_M1005_d
+ N_A_84_21#_M1000_g N_A_84_21#_M1001_g N_A_84_21#_M1003_g N_A_84_21#_M1006_g
+ N_A_84_21#_M1004_g N_A_84_21#_M1011_g N_A_84_21#_M1018_g N_A_84_21#_M1015_g
+ N_A_84_21#_c_132_n N_A_84_21#_c_133_n N_A_84_21#_c_134_n N_A_84_21#_c_135_n
+ N_A_84_21#_c_136_n N_A_84_21#_c_222_p N_A_84_21#_c_145_n N_A_84_21#_c_153_p
+ N_A_84_21#_c_198_p N_A_84_21#_c_146_n N_A_84_21#_c_147_n N_A_84_21#_c_137_n
+ N_A_84_21#_c_138_n N_A_84_21#_c_148_n N_A_84_21#_c_149_n N_A_84_21#_c_139_n
+ N_A_84_21#_c_140_n PM_SKY130_FD_SC_LP__EBUFN_4%A_84_21#
x_PM_SKY130_FD_SC_LP__EBUFN_4%A_456_21# N_A_456_21#_M1012_s N_A_456_21#_M1002_s
+ N_A_456_21#_c_286_n N_A_456_21#_M1008_g N_A_456_21#_c_287_n
+ N_A_456_21#_c_288_n N_A_456_21#_c_289_n N_A_456_21#_M1010_g
+ N_A_456_21#_c_290_n N_A_456_21#_c_291_n N_A_456_21#_M1013_g
+ N_A_456_21#_c_292_n N_A_456_21#_c_293_n N_A_456_21#_M1014_g
+ N_A_456_21#_c_294_n N_A_456_21#_c_295_n N_A_456_21#_c_296_n
+ N_A_456_21#_c_297_n N_A_456_21#_c_298_n N_A_456_21#_c_299_n
+ N_A_456_21#_c_303_n N_A_456_21#_c_300_n N_A_456_21#_c_301_n
+ N_A_456_21#_c_302_n PM_SKY130_FD_SC_LP__EBUFN_4%A_456_21#
x_PM_SKY130_FD_SC_LP__EBUFN_4%TE_B N_TE_B_c_410_n N_TE_B_M1007_g N_TE_B_c_395_n
+ N_TE_B_c_396_n N_TE_B_c_413_n N_TE_B_M1009_g N_TE_B_c_397_n N_TE_B_c_415_n
+ N_TE_B_M1016_g N_TE_B_c_398_n N_TE_B_c_417_n N_TE_B_M1017_g N_TE_B_c_399_n
+ N_TE_B_c_400_n N_TE_B_M1012_g N_TE_B_M1002_g N_TE_B_c_403_n N_TE_B_c_404_n
+ N_TE_B_c_405_n N_TE_B_c_406_n TE_B TE_B TE_B N_TE_B_c_408_n N_TE_B_c_409_n
+ PM_SKY130_FD_SC_LP__EBUFN_4%TE_B
x_PM_SKY130_FD_SC_LP__EBUFN_4%A N_A_M1005_g N_A_M1019_g A N_A_c_528_n
+ N_A_c_529_n PM_SKY130_FD_SC_LP__EBUFN_4%A
x_PM_SKY130_FD_SC_LP__EBUFN_4%A_27_367# N_A_27_367#_M1001_s N_A_27_367#_M1006_s
+ N_A_27_367#_M1015_s N_A_27_367#_M1009_d N_A_27_367#_M1017_d
+ N_A_27_367#_c_563_n N_A_27_367#_c_564_n N_A_27_367#_c_574_n
+ N_A_27_367#_c_576_n N_A_27_367#_c_578_n N_A_27_367#_c_580_n
+ N_A_27_367#_c_589_n N_A_27_367#_c_582_n N_A_27_367#_c_565_n
+ N_A_27_367#_c_566_n N_A_27_367#_c_585_n N_A_27_367#_c_586_n
+ N_A_27_367#_c_603_n PM_SKY130_FD_SC_LP__EBUFN_4%A_27_367#
x_PM_SKY130_FD_SC_LP__EBUFN_4%Z N_Z_M1000_d N_Z_M1004_d N_Z_M1001_d N_Z_M1011_d
+ N_Z_c_646_n N_Z_c_639_n N_Z_c_642_n N_Z_c_640_n N_Z_c_643_n N_Z_c_668_n
+ N_Z_c_641_n N_Z_c_644_n N_Z_c_645_n Z PM_SKY130_FD_SC_LP__EBUFN_4%Z
x_PM_SKY130_FD_SC_LP__EBUFN_4%VPWR N_VPWR_M1007_s N_VPWR_M1016_s N_VPWR_M1002_d
+ N_VPWR_c_705_n N_VPWR_c_706_n N_VPWR_c_707_n N_VPWR_c_708_n N_VPWR_c_709_n
+ N_VPWR_c_710_n VPWR N_VPWR_c_711_n N_VPWR_c_712_n N_VPWR_c_704_n
+ N_VPWR_c_714_n N_VPWR_c_715_n PM_SKY130_FD_SC_LP__EBUFN_4%VPWR
x_PM_SKY130_FD_SC_LP__EBUFN_4%A_27_47# N_A_27_47#_M1000_s N_A_27_47#_M1003_s
+ N_A_27_47#_M1018_s N_A_27_47#_M1010_s N_A_27_47#_M1014_s N_A_27_47#_c_785_n
+ N_A_27_47#_c_787_n N_A_27_47#_c_836_p N_A_27_47#_c_778_n N_A_27_47#_c_779_n
+ N_A_27_47#_c_780_n N_A_27_47#_c_833_p N_A_27_47#_c_781_n N_A_27_47#_c_782_n
+ N_A_27_47#_c_783_n N_A_27_47#_c_792_n N_A_27_47#_c_784_n
+ PM_SKY130_FD_SC_LP__EBUFN_4%A_27_47#
x_PM_SKY130_FD_SC_LP__EBUFN_4%VGND N_VGND_M1008_d N_VGND_M1013_d N_VGND_M1012_d
+ N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n N_VGND_c_857_n
+ VGND N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n
+ N_VGND_c_862_n N_VGND_c_863_n PM_SKY130_FD_SC_LP__EBUFN_4%VGND
cc_1 VNB N_A_84_21#_M1000_g 0.0290732f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_A_84_21#_M1001_g 6.86639e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_A_84_21#_M1003_g 0.0231539f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_4 VNB N_A_84_21#_M1006_g 4.80242e-19 $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_5 VNB N_A_84_21#_M1004_g 0.0241745f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.655
cc_6 VNB N_A_84_21#_M1011_g 5.06756e-19 $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.465
cc_7 VNB N_A_84_21#_M1018_g 0.0238926f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.655
cc_8 VNB N_A_84_21#_M1015_g 5.16052e-19 $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.465
cc_9 VNB N_A_84_21#_c_132_n 0.0412411f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.48
cc_10 VNB N_A_84_21#_c_133_n 0.0204046f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.48
cc_11 VNB N_A_84_21#_c_134_n 0.00525339f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.48
cc_12 VNB N_A_84_21#_c_135_n 0.0207548f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.48
cc_13 VNB N_A_84_21#_c_136_n 0.017361f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.48
cc_14 VNB N_A_84_21#_c_137_n 0.0302364f $X=-0.19 $Y=-0.245 $X2=5.945 $Y2=0.42
cc_15 VNB N_A_84_21#_c_138_n 0.0108069f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.48
cc_16 VNB N_A_84_21#_c_139_n 0.0246046f $X=-0.19 $Y=-0.245 $X2=5.927 $Y2=1.95
cc_17 VNB N_A_84_21#_c_140_n 0.014232f $X=-0.19 $Y=-0.245 $X2=5.962 $Y2=1.135
cc_18 VNB N_A_456_21#_c_286_n 0.0157226f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.315
cc_19 VNB N_A_456_21#_c_287_n 0.0123225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_456_21#_c_288_n 0.00866446f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.645
cc_21 VNB N_A_456_21#_c_289_n 0.0155656f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_22 VNB N_A_456_21#_c_290_n 0.0123225f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.315
cc_23 VNB N_A_456_21#_c_291_n 0.0159719f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_24 VNB N_A_456_21#_c_292_n 0.0111217f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_25 VNB N_A_456_21#_c_293_n 0.0190765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_456_21#_c_294_n 0.0217417f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.655
cc_27 VNB N_A_456_21#_c_295_n 0.0142621f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.465
cc_28 VNB N_A_456_21#_c_296_n 0.00514676f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.465
cc_29 VNB N_A_456_21#_c_297_n 0.00514676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_456_21#_c_298_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.315
cc_31 VNB N_A_456_21#_c_299_n 0.0251274f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.655
cc_32 VNB N_A_456_21#_c_300_n 0.00418204f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.48
cc_33 VNB N_A_456_21#_c_301_n 0.0522743f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.48
cc_34 VNB N_A_456_21#_c_302_n 0.0168545f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.48
cc_35 VNB N_TE_B_c_395_n 0.010921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_TE_B_c_396_n 0.00579485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_TE_B_c_397_n 0.0073704f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_38 VNB N_TE_B_c_398_n 0.0119983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_TE_B_c_399_n 0.0106036f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.645
cc_40 VNB N_TE_B_c_400_n 0.0169806f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_41 VNB N_TE_B_M1012_g 0.0242829f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.655
cc_42 VNB N_TE_B_M1002_g 0.0103684f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.465
cc_43 VNB N_TE_B_c_403_n 0.00401367f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.315
cc_44 VNB N_TE_B_c_404_n 0.0040279f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.655
cc_45 VNB N_TE_B_c_405_n 0.00594802f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.655
cc_46 VNB N_TE_B_c_406_n 0.00567891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB TE_B 0.00350142f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.465
cc_48 VNB N_TE_B_c_408_n 0.0332269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_TE_B_c_409_n 0.0191059f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.48
cc_50 VNB N_A_M1019_g 0.0296948f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.315
cc_51 VNB N_A_c_528_n 0.0270868f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_52 VNB N_A_c_529_n 0.00608412f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_53 VNB N_Z_c_639_n 0.00365946f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_54 VNB N_Z_c_640_n 0.00537078f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_55 VNB N_Z_c_641_n 0.0194168f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.655
cc_56 VNB N_VPWR_c_704_n 0.263193f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.48
cc_57 VNB N_A_27_47#_c_778_n 9.63636e-19 $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.655
cc_58 VNB N_A_27_47#_c_779_n 0.00825628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_47#_c_780_n 0.00389025f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.645
cc_60 VNB N_A_27_47#_c_781_n 0.0012126f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.655
cc_61 VNB N_A_27_47#_c_782_n 0.00643864f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.465
cc_62 VNB N_A_27_47#_c_783_n 0.0291024f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.48
cc_63 VNB N_A_27_47#_c_784_n 0.00159014f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.48
cc_64 VNB N_VGND_c_853_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_65 VNB N_VGND_c_854_n 0.00229788f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_66 VNB N_VGND_c_855_n 0.0138211f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_67 VNB N_VGND_c_856_n 0.0131279f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.315
cc_68 VNB N_VGND_c_857_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.655
cc_69 VNB N_VGND_c_858_n 0.0572155f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.645
cc_70 VNB N_VGND_c_859_n 0.0449995f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.48
cc_71 VNB N_VGND_c_860_n 0.0186517f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.48
cc_72 VNB N_VGND_c_861_n 0.326903f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.48
cc_73 VNB N_VGND_c_862_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_863_n 0.00634044f $X=-0.19 $Y=-0.245 $X2=4.325 $Y2=2.1
cc_75 VPB N_A_84_21#_M1001_g 0.0264959f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_76 VPB N_A_84_21#_M1006_g 0.0204154f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_77 VPB N_A_84_21#_M1011_g 0.0212747f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.465
cc_78 VPB N_A_84_21#_M1015_g 0.0216247f $X=-0.19 $Y=1.655 $X2=1.925 $Y2=2.465
cc_79 VPB N_A_84_21#_c_145_n 0.0035164f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.015
cc_80 VPB N_A_84_21#_c_146_n 0.0101516f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=2.27
cc_81 VPB N_A_84_21#_c_147_n 0.0319178f $X=-0.19 $Y=1.655 $X2=5.875 $Y2=2.91
cc_82 VPB N_A_84_21#_c_148_n 0.00811699f $X=-0.19 $Y=1.655 $X2=4.41 $Y2=2.1
cc_83 VPB N_A_84_21#_c_149_n 0.0174703f $X=-0.19 $Y=1.655 $X2=5.875 $Y2=2.115
cc_84 VPB N_A_84_21#_c_139_n 0.0133303f $X=-0.19 $Y=1.655 $X2=5.927 $Y2=1.95
cc_85 VPB N_A_456_21#_c_303_n 0.00897434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_456_21#_c_300_n 0.0032342f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.48
cc_87 VPB N_TE_B_c_410_n 0.0182474f $X=-0.19 $Y=1.655 $X2=5.805 $Y2=0.275
cc_88 VPB N_TE_B_c_395_n 0.00890451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_TE_B_c_396_n 0.00267287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_TE_B_c_413_n 0.017441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_TE_B_c_397_n 0.0044816f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.655
cc_92 VPB N_TE_B_c_415_n 0.0177433f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.645
cc_93 VPB N_TE_B_c_398_n 0.0101682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_TE_B_c_417_n 0.0223919f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_95 VPB N_TE_B_c_399_n 0.0101283f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.645
cc_96 VPB N_TE_B_M1002_g 0.0257193f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.465
cc_97 VPB N_TE_B_c_403_n 0.00111435f $X=-0.19 $Y=1.655 $X2=1.925 $Y2=1.315
cc_98 VPB N_TE_B_c_404_n 0.00111435f $X=-0.19 $Y=1.655 $X2=1.925 $Y2=0.655
cc_99 VPB N_TE_B_c_405_n 0.00277251f $X=-0.19 $Y=1.655 $X2=1.925 $Y2=0.655
cc_100 VPB N_TE_B_c_408_n 0.0141129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_M1005_g 0.0233469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_c_528_n 0.00652972f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_103 VPB N_A_c_529_n 0.00492264f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_104 VPB N_A_27_367#_c_563_n 0.00719502f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_105 VPB N_A_27_367#_c_564_n 0.0438458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_27_367#_c_565_n 0.0032868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_27_367#_c_566_n 0.00649576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_Z_c_642_n 0.00150187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_Z_c_643_n 0.00307912f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.315
cc_110 VPB N_Z_c_644_n 0.00185767f $X=-0.19 $Y=1.655 $X2=1.925 $Y2=1.645
cc_111 VPB N_Z_c_645_n 0.00230938f $X=-0.19 $Y=1.655 $X2=1.925 $Y2=2.465
cc_112 VPB N_VPWR_c_705_n 0.00499451f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_113 VPB N_VPWR_c_706_n 0.0171854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_707_n 0.00505705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_708_n 0.00278884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_709_n 0.037217f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.655
cc_117 VPB N_VPWR_c_710_n 0.00510509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_711_n 0.0611809f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.465
cc_119 VPB N_VPWR_c_712_n 0.020221f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.48
cc_120 VPB N_VPWR_c_704_n 0.0583776f $X=-0.19 $Y=1.655 $X2=1.85 $Y2=1.48
cc_121 VPB N_VPWR_c_714_n 0.00631648f $X=-0.19 $Y=1.655 $X2=1.04 $Y2=1.48
cc_122 VPB N_VPWR_c_715_n 0.0063111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 N_A_84_21#_c_146_n N_A_456_21#_M1002_s 0.0186731f $X=5.71 $Y=2.27 $X2=0
+ $Y2=0
cc_124 N_A_84_21#_M1018_g N_A_456_21#_c_286_n 0.0106815f $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_125 N_A_84_21#_c_153_p N_A_456_21#_c_287_n 0.00133341f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_126 N_A_84_21#_c_136_n N_A_456_21#_c_288_n 0.0106815f $X=1.925 $Y=1.48 $X2=0
+ $Y2=0
cc_127 N_A_84_21#_c_153_p N_A_456_21#_c_288_n 0.00164582f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_128 N_A_84_21#_c_153_p N_A_456_21#_c_290_n 0.00160993f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_129 N_A_84_21#_c_153_p N_A_456_21#_c_292_n 6.97582e-19 $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_130 N_A_84_21#_c_146_n N_A_456_21#_c_303_n 0.0296069f $X=5.71 $Y=2.27 $X2=0
+ $Y2=0
cc_131 N_A_84_21#_c_149_n N_A_456_21#_c_303_n 0.00179975f $X=5.875 $Y=2.115
+ $X2=0 $Y2=0
cc_132 N_A_84_21#_M1015_g N_TE_B_c_410_n 0.0189506f $X=1.925 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_84_21#_c_153_p N_TE_B_c_410_n 0.0122134f $X=4.325 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A_84_21#_c_153_p N_TE_B_c_395_n 0.00722723f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_135 N_A_84_21#_c_136_n N_TE_B_c_396_n 0.0189506f $X=1.925 $Y=1.48 $X2=0 $Y2=0
cc_136 N_A_84_21#_c_145_n N_TE_B_c_396_n 0.00838348f $X=2.13 $Y=2.015 $X2=0
+ $Y2=0
cc_137 N_A_84_21#_c_138_n N_TE_B_c_396_n 0.00219557f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_138 N_A_84_21#_c_153_p N_TE_B_c_413_n 0.012187f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_139 N_A_84_21#_c_153_p N_TE_B_c_397_n 0.00301135f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_140 N_A_84_21#_c_153_p N_TE_B_c_415_n 0.0131687f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_141 N_A_84_21#_c_153_p N_TE_B_c_398_n 0.0056463f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_142 N_A_84_21#_c_153_p N_TE_B_c_417_n 0.0148313f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_143 N_A_84_21#_c_148_n N_TE_B_c_417_n 0.00630378f $X=4.41 $Y=2.1 $X2=0 $Y2=0
cc_144 N_A_84_21#_c_153_p N_TE_B_c_399_n 0.00387648f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_145 N_A_84_21#_c_148_n N_TE_B_c_399_n 0.00354059f $X=4.41 $Y=2.1 $X2=0 $Y2=0
cc_146 N_A_84_21#_c_146_n N_TE_B_M1002_g 0.0203674f $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_147 N_A_84_21#_c_147_n N_TE_B_M1002_g 2.03066e-19 $X=5.875 $Y=2.91 $X2=0
+ $Y2=0
cc_148 N_A_84_21#_c_148_n N_TE_B_M1002_g 0.00412076f $X=4.41 $Y=2.1 $X2=0 $Y2=0
cc_149 N_A_84_21#_c_149_n N_TE_B_M1002_g 0.00188565f $X=5.875 $Y=2.115 $X2=0
+ $Y2=0
cc_150 N_A_84_21#_c_146_n TE_B 0.00506395f $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_151 N_A_84_21#_c_148_n TE_B 0.00218642f $X=4.41 $Y=2.1 $X2=0 $Y2=0
cc_152 N_A_84_21#_c_146_n N_TE_B_c_408_n 0.00336618f $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_153 N_A_84_21#_c_153_p N_TE_B_c_409_n 0.0225286f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_154 N_A_84_21#_c_148_n N_TE_B_c_409_n 0.00368458f $X=4.41 $Y=2.1 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_146_n N_A_M1005_g 0.0131261f $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_156 N_A_84_21#_c_147_n N_A_M1005_g 0.00939097f $X=5.875 $Y=2.91 $X2=0 $Y2=0
cc_157 N_A_84_21#_c_149_n N_A_M1005_g 0.00594566f $X=5.875 $Y=2.115 $X2=0 $Y2=0
cc_158 N_A_84_21#_c_139_n N_A_M1005_g 0.00442969f $X=5.927 $Y=1.95 $X2=0 $Y2=0
cc_159 N_A_84_21#_c_137_n N_A_M1019_g 0.0110938f $X=5.945 $Y=0.42 $X2=0 $Y2=0
cc_160 N_A_84_21#_c_139_n N_A_M1019_g 0.0128598f $X=5.927 $Y=1.95 $X2=0 $Y2=0
cc_161 N_A_84_21#_c_140_n N_A_M1019_g 0.00264415f $X=5.962 $Y=1.135 $X2=0 $Y2=0
cc_162 N_A_84_21#_c_146_n N_A_c_528_n 3.83522e-19 $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_163 N_A_84_21#_c_149_n N_A_c_528_n 2.73982e-19 $X=5.875 $Y=2.115 $X2=0 $Y2=0
cc_164 N_A_84_21#_c_146_n N_A_c_529_n 0.0111644f $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_165 N_A_84_21#_c_149_n N_A_c_529_n 0.00548606f $X=5.875 $Y=2.115 $X2=0 $Y2=0
cc_166 N_A_84_21#_c_139_n N_A_c_529_n 0.0336246f $X=5.927 $Y=1.95 $X2=0 $Y2=0
cc_167 N_A_84_21#_c_140_n N_A_c_529_n 0.00158719f $X=5.962 $Y=1.135 $X2=0 $Y2=0
cc_168 N_A_84_21#_c_145_n N_A_27_367#_M1015_s 0.00315411f $X=2.13 $Y=2.015 $X2=0
+ $Y2=0
cc_169 N_A_84_21#_c_153_p N_A_27_367#_M1015_s 0.00349253f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_170 N_A_84_21#_c_198_p N_A_27_367#_M1015_s 0.00280297f $X=2.215 $Y=2.1 $X2=0
+ $Y2=0
cc_171 N_A_84_21#_c_153_p N_A_27_367#_M1009_d 0.00421743f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_172 N_A_84_21#_c_153_p N_A_27_367#_M1017_d 0.00555623f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_173 N_A_84_21#_c_148_n N_A_27_367#_M1017_d 0.00558334f $X=4.41 $Y=2.1 $X2=0
+ $Y2=0
cc_174 N_A_84_21#_M1001_g N_A_27_367#_c_564_n 0.00331374f $X=0.495 $Y=2.465
+ $X2=0 $Y2=0
cc_175 N_A_84_21#_M1001_g N_A_27_367#_c_574_n 0.0111972f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_84_21#_M1006_g N_A_27_367#_c_574_n 0.0139716f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_84_21#_M1011_g N_A_27_367#_c_576_n 0.00963573f $X=1.425 $Y=2.465
+ $X2=0 $Y2=0
cc_178 N_A_84_21#_M1015_g N_A_27_367#_c_576_n 5.42008e-19 $X=1.925 $Y=2.465
+ $X2=0 $Y2=0
cc_179 N_A_84_21#_M1011_g N_A_27_367#_c_578_n 0.0109138f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_84_21#_M1015_g N_A_27_367#_c_578_n 0.0143041f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_84_21#_c_153_p N_A_27_367#_c_580_n 0.00821038f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_182 N_A_84_21#_c_198_p N_A_27_367#_c_580_n 0.0143066f $X=2.215 $Y=2.1 $X2=0
+ $Y2=0
cc_183 N_A_84_21#_c_153_p N_A_27_367#_c_582_n 0.039137f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_184 N_A_84_21#_c_153_p N_A_27_367#_c_565_n 0.033449f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_185 N_A_84_21#_c_148_n N_A_27_367#_c_565_n 0.00757418f $X=4.41 $Y=2.1 $X2=0
+ $Y2=0
cc_186 N_A_84_21#_M1011_g N_A_27_367#_c_585_n 5.89773e-19 $X=1.425 $Y=2.465
+ $X2=0 $Y2=0
cc_187 N_A_84_21#_c_153_p N_A_27_367#_c_586_n 0.017158f $X=4.325 $Y=2.1 $X2=0
+ $Y2=0
cc_188 N_A_84_21#_M1000_g N_Z_c_646_n 0.00496215f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A_84_21#_M1003_g N_Z_c_646_n 0.0060416f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_190 N_A_84_21#_M1004_g N_Z_c_646_n 2.75157e-19 $X=1.425 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A_84_21#_M1000_g N_Z_c_639_n 0.0116856f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_84_21#_M1003_g N_Z_c_639_n 0.00722618f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A_84_21#_c_132_n N_Z_c_639_n 0.00558967f $X=1 $Y=1.48 $X2=0 $Y2=0
cc_194 N_A_84_21#_c_222_p N_Z_c_639_n 0.00786305f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_195 N_A_84_21#_M1001_g N_Z_c_642_n 0.00809756f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_84_21#_M1006_g N_Z_c_642_n 0.00360365f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_84_21#_c_132_n N_Z_c_642_n 0.0168513f $X=1 $Y=1.48 $X2=0 $Y2=0
cc_198 N_A_84_21#_c_222_p N_Z_c_642_n 0.017791f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_199 N_A_84_21#_M1003_g N_Z_c_640_n 0.00929135f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A_84_21#_M1004_g N_Z_c_640_n 0.012812f $X=1.425 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_84_21#_M1018_g N_Z_c_640_n 0.00418491f $X=1.925 $Y=0.655 $X2=0 $Y2=0
cc_202 N_A_84_21#_c_133_n N_Z_c_640_n 0.00381149f $X=1.35 $Y=1.48 $X2=0 $Y2=0
cc_203 N_A_84_21#_c_135_n N_Z_c_640_n 0.0033142f $X=1.85 $Y=1.48 $X2=0 $Y2=0
cc_204 N_A_84_21#_c_222_p N_Z_c_640_n 0.0636116f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_205 N_A_84_21#_c_138_n N_Z_c_640_n 0.0127632f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_206 N_A_84_21#_M1006_g N_Z_c_643_n 0.0115433f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_84_21#_M1011_g N_Z_c_643_n 0.0151263f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_84_21#_c_133_n N_Z_c_643_n 0.00381149f $X=1.35 $Y=1.48 $X2=0 $Y2=0
cc_209 N_A_84_21#_c_222_p N_Z_c_643_n 0.0491449f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_210 N_A_84_21#_M1018_g N_Z_c_668_n 0.00443774f $X=1.925 $Y=0.655 $X2=0 $Y2=0
cc_211 N_A_84_21#_M1000_g N_Z_c_641_n 0.00931592f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A_84_21#_c_132_n N_Z_c_641_n 0.00811537f $X=1 $Y=1.48 $X2=0 $Y2=0
cc_213 N_A_84_21#_M1001_g N_Z_c_644_n 0.0135322f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A_84_21#_M1006_g N_Z_c_644_n 0.0133609f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_84_21#_M1011_g N_Z_c_644_n 2.75157e-19 $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_84_21#_c_132_n N_Z_c_644_n 0.00165908f $X=1 $Y=1.48 $X2=0 $Y2=0
cc_217 N_A_84_21#_M1015_g N_Z_c_645_n 0.0152686f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_84_21#_c_135_n N_Z_c_645_n 0.00334502f $X=1.85 $Y=1.48 $X2=0 $Y2=0
cc_219 N_A_84_21#_c_222_p N_Z_c_645_n 0.0147215f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_220 N_A_84_21#_c_145_n N_Z_c_645_n 0.00787895f $X=2.13 $Y=2.015 $X2=0 $Y2=0
cc_221 N_A_84_21#_c_138_n N_Z_c_645_n 0.0129867f $X=1.72 $Y=1.48 $X2=0 $Y2=0
cc_222 N_A_84_21#_c_153_p N_VPWR_M1007_s 0.00805614f $X=4.325 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_84_21#_c_153_p N_VPWR_M1016_s 0.011402f $X=4.325 $Y=2.1 $X2=0 $Y2=0
cc_224 N_A_84_21#_c_146_n N_VPWR_M1002_d 0.00870626f $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_225 N_A_84_21#_c_146_n N_VPWR_c_708_n 0.0210288f $X=5.71 $Y=2.27 $X2=0 $Y2=0
cc_226 N_A_84_21#_M1001_g N_VPWR_c_711_n 0.00357877f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_227 N_A_84_21#_M1006_g N_VPWR_c_711_n 0.00357877f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_228 N_A_84_21#_M1011_g N_VPWR_c_711_n 0.00357842f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_229 N_A_84_21#_M1015_g N_VPWR_c_711_n 0.00357877f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_230 N_A_84_21#_c_147_n N_VPWR_c_712_n 0.0285463f $X=5.875 $Y=2.91 $X2=0 $Y2=0
cc_231 N_A_84_21#_M1005_d N_VPWR_c_704_n 0.00231914f $X=5.735 $Y=1.835 $X2=0
+ $Y2=0
cc_232 N_A_84_21#_M1001_g N_VPWR_c_704_n 0.0063022f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_84_21#_M1006_g N_VPWR_c_704_n 0.00560622f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A_84_21#_M1011_g N_VPWR_c_704_n 0.00570659f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A_84_21#_M1015_g N_VPWR_c_704_n 0.00580544f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_236 N_A_84_21#_c_147_n N_VPWR_c_704_n 0.016651f $X=5.875 $Y=2.91 $X2=0 $Y2=0
cc_237 N_A_84_21#_M1000_g N_A_27_47#_c_785_n 0.0111972f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_238 N_A_84_21#_M1003_g N_A_27_47#_c_785_n 0.0116573f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_84_21#_M1004_g N_A_27_47#_c_787_n 0.00866186f $X=1.425 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_84_21#_M1018_g N_A_27_47#_c_787_n 0.0118963f $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_241 N_A_84_21#_M1018_g N_A_27_47#_c_778_n 9.26489e-19 $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_242 N_A_84_21#_M1018_g N_A_27_47#_c_780_n 0.00514561f $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_243 N_A_84_21#_c_138_n N_A_27_47#_c_780_n 0.0150404f $X=1.72 $Y=1.48 $X2=0
+ $Y2=0
cc_244 N_A_84_21#_M1004_g N_A_27_47#_c_792_n 0.00631927f $X=1.425 $Y=0.655 $X2=0
+ $Y2=0
cc_245 N_A_84_21#_M1018_g N_A_27_47#_c_792_n 8.57461e-19 $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_84_21#_M1018_g N_VGND_c_853_n 0.00109254f $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_A_84_21#_c_137_n N_VGND_c_855_n 0.035076f $X=5.945 $Y=0.42 $X2=0 $Y2=0
cc_248 N_A_84_21#_M1000_g N_VGND_c_858_n 0.00357877f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_249 N_A_84_21#_M1003_g N_VGND_c_858_n 0.00357877f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_250 N_A_84_21#_M1004_g N_VGND_c_858_n 0.00357842f $X=1.425 $Y=0.655 $X2=0
+ $Y2=0
cc_251 N_A_84_21#_M1018_g N_VGND_c_858_n 0.00357877f $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_252 N_A_84_21#_c_137_n N_VGND_c_860_n 0.0259379f $X=5.945 $Y=0.42 $X2=0 $Y2=0
cc_253 N_A_84_21#_M1000_g N_VGND_c_861_n 0.0063022f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_254 N_A_84_21#_M1003_g N_VGND_c_861_n 0.00560622f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_255 N_A_84_21#_M1004_g N_VGND_c_861_n 0.00570659f $X=1.425 $Y=0.655 $X2=0
+ $Y2=0
cc_256 N_A_84_21#_M1018_g N_VGND_c_861_n 0.00556082f $X=1.925 $Y=0.655 $X2=0
+ $Y2=0
cc_257 N_A_84_21#_c_137_n N_VGND_c_861_n 0.0140028f $X=5.945 $Y=0.42 $X2=0 $Y2=0
cc_258 N_A_456_21#_c_287_n N_TE_B_c_395_n 0.0156123f $X=2.71 $Y=1.26 $X2=0 $Y2=0
cc_259 N_A_456_21#_c_288_n N_TE_B_c_396_n 0.0156123f $X=2.43 $Y=1.26 $X2=0 $Y2=0
cc_260 N_A_456_21#_c_297_n N_TE_B_c_397_n 0.0156123f $X=3.215 $Y=1.26 $X2=0
+ $Y2=0
cc_261 N_A_456_21#_c_298_n N_TE_B_c_398_n 0.0156123f $X=3.645 $Y=1.26 $X2=0
+ $Y2=0
cc_262 N_A_456_21#_c_303_n N_TE_B_c_417_n 0.00640569f $X=4.94 $Y=1.89 $X2=0
+ $Y2=0
cc_263 N_A_456_21#_c_299_n N_TE_B_c_399_n 0.00319063f $X=4.302 $Y=1.01 $X2=0
+ $Y2=0
cc_264 N_A_456_21#_c_303_n N_TE_B_c_400_n 0.00235249f $X=4.94 $Y=1.89 $X2=0
+ $Y2=0
cc_265 N_A_456_21#_c_300_n N_TE_B_c_400_n 0.00886772f $X=5.025 $Y=1.765 $X2=0
+ $Y2=0
cc_266 N_A_456_21#_c_300_n N_TE_B_M1012_g 0.00759406f $X=5.025 $Y=1.765 $X2=0
+ $Y2=0
cc_267 N_A_456_21#_c_301_n N_TE_B_M1012_g 0.00553782f $X=4.36 $Y=0.505 $X2=0
+ $Y2=0
cc_268 N_A_456_21#_c_302_n N_TE_B_M1012_g 0.00905321f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_269 N_A_456_21#_c_303_n N_TE_B_M1002_g 0.0105615f $X=4.94 $Y=1.89 $X2=0 $Y2=0
cc_270 N_A_456_21#_c_300_n N_TE_B_M1002_g 0.00795932f $X=5.025 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_456_21#_c_296_n N_TE_B_c_403_n 0.0156123f $X=2.785 $Y=1.26 $X2=0
+ $Y2=0
cc_272 N_A_456_21#_c_292_n N_TE_B_c_404_n 0.0156123f $X=3.57 $Y=1.26 $X2=0 $Y2=0
cc_273 N_A_456_21#_c_294_n N_TE_B_c_405_n 0.0169497f $X=4.08 $Y=1.26 $X2=0 $Y2=0
cc_274 N_A_456_21#_c_300_n N_TE_B_c_406_n 0.00243152f $X=5.025 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_A_456_21#_c_295_n TE_B 3.5073e-19 $X=4.155 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A_456_21#_c_299_n TE_B 2.97803e-19 $X=4.302 $Y=1.01 $X2=0 $Y2=0
cc_277 N_A_456_21#_c_303_n TE_B 0.00823012f $X=4.94 $Y=1.89 $X2=0 $Y2=0
cc_278 N_A_456_21#_c_300_n TE_B 0.0309789f $X=5.025 $Y=1.765 $X2=0 $Y2=0
cc_279 N_A_456_21#_c_302_n TE_B 0.0292157f $X=4.945 $Y=0.42 $X2=0 $Y2=0
cc_280 N_A_456_21#_c_294_n N_TE_B_c_408_n 0.00457864f $X=4.08 $Y=1.26 $X2=0
+ $Y2=0
cc_281 N_A_456_21#_c_299_n N_TE_B_c_408_n 0.00436578f $X=4.302 $Y=1.01 $X2=0
+ $Y2=0
cc_282 N_A_456_21#_c_303_n N_TE_B_c_408_n 0.0028411f $X=4.94 $Y=1.89 $X2=0 $Y2=0
cc_283 N_A_456_21#_c_300_n N_TE_B_c_408_n 0.00350132f $X=5.025 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A_456_21#_c_302_n N_TE_B_c_408_n 0.00861956f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_285 N_A_456_21#_c_292_n N_TE_B_c_409_n 0.00587908f $X=3.57 $Y=1.26 $X2=0
+ $Y2=0
cc_286 N_A_456_21#_c_293_n N_TE_B_c_409_n 0.0021218f $X=3.645 $Y=1.185 $X2=0
+ $Y2=0
cc_287 N_A_456_21#_c_294_n N_TE_B_c_409_n 0.0137995f $X=4.08 $Y=1.26 $X2=0 $Y2=0
cc_288 N_A_456_21#_c_295_n N_TE_B_c_409_n 0.0057939f $X=4.155 $Y=1.185 $X2=0
+ $Y2=0
cc_289 N_A_456_21#_c_298_n N_TE_B_c_409_n 0.00277321f $X=3.645 $Y=1.26 $X2=0
+ $Y2=0
cc_290 N_A_456_21#_c_299_n N_TE_B_c_409_n 8.36173e-19 $X=4.302 $Y=1.01 $X2=0
+ $Y2=0
cc_291 N_A_456_21#_c_302_n N_TE_B_c_409_n 0.0198548f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_292 N_A_456_21#_c_303_n N_A_M1005_g 0.00101407f $X=4.94 $Y=1.89 $X2=0 $Y2=0
cc_293 N_A_456_21#_c_300_n N_A_M1019_g 9.86252e-19 $X=5.025 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A_456_21#_c_300_n N_A_c_528_n 3.17777e-19 $X=5.025 $Y=1.765 $X2=0 $Y2=0
cc_295 N_A_456_21#_c_303_n N_A_c_529_n 8.21121e-19 $X=4.94 $Y=1.89 $X2=0 $Y2=0
cc_296 N_A_456_21#_c_300_n N_A_c_529_n 0.0213788f $X=5.025 $Y=1.765 $X2=0 $Y2=0
cc_297 N_A_456_21#_M1002_s N_VPWR_c_704_n 0.0172056f $X=4.685 $Y=1.785 $X2=0
+ $Y2=0
cc_298 N_A_456_21#_c_286_n N_A_27_47#_c_778_n 0.00189764f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_299 N_A_456_21#_c_286_n N_A_27_47#_c_779_n 0.00757398f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_300 N_A_456_21#_c_287_n N_A_27_47#_c_779_n 0.00817193f $X=2.71 $Y=1.26 $X2=0
+ $Y2=0
cc_301 N_A_456_21#_c_288_n N_A_27_47#_c_779_n 0.00636401f $X=2.43 $Y=1.26 $X2=0
+ $Y2=0
cc_302 N_A_456_21#_c_289_n N_A_27_47#_c_779_n 0.00736574f $X=2.785 $Y=1.185
+ $X2=0 $Y2=0
cc_303 N_A_456_21#_c_290_n N_A_27_47#_c_779_n 0.0016711f $X=3.14 $Y=1.26 $X2=0
+ $Y2=0
cc_304 N_A_456_21#_c_296_n N_A_27_47#_c_779_n 0.00359985f $X=2.785 $Y=1.26 $X2=0
+ $Y2=0
cc_305 N_A_456_21#_c_291_n N_A_27_47#_c_781_n 0.0103941f $X=3.215 $Y=1.185 $X2=0
+ $Y2=0
cc_306 N_A_456_21#_c_292_n N_A_27_47#_c_781_n 0.00340523f $X=3.57 $Y=1.26 $X2=0
+ $Y2=0
cc_307 N_A_456_21#_c_293_n N_A_27_47#_c_781_n 0.00925856f $X=3.645 $Y=1.185
+ $X2=0 $Y2=0
cc_308 N_A_456_21#_c_294_n N_A_27_47#_c_781_n 0.00142459f $X=4.08 $Y=1.26 $X2=0
+ $Y2=0
cc_309 N_A_456_21#_c_299_n N_A_27_47#_c_781_n 0.00179468f $X=4.302 $Y=1.01 $X2=0
+ $Y2=0
cc_310 N_A_456_21#_c_302_n N_A_27_47#_c_781_n 0.0151542f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_311 N_A_456_21#_c_291_n N_A_27_47#_c_782_n 6.55694e-19 $X=3.215 $Y=1.185
+ $X2=0 $Y2=0
cc_312 N_A_456_21#_c_293_n N_A_27_47#_c_782_n 0.00807611f $X=3.645 $Y=1.185
+ $X2=0 $Y2=0
cc_313 N_A_456_21#_c_301_n N_A_27_47#_c_782_n 0.00495189f $X=4.36 $Y=0.505 $X2=0
+ $Y2=0
cc_314 N_A_456_21#_c_302_n N_A_27_47#_c_782_n 0.0418682f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_315 N_A_456_21#_c_289_n N_A_27_47#_c_784_n 0.00203628f $X=2.785 $Y=1.185
+ $X2=0 $Y2=0
cc_316 N_A_456_21#_c_290_n N_A_27_47#_c_784_n 0.00983516f $X=3.14 $Y=1.26 $X2=0
+ $Y2=0
cc_317 N_A_456_21#_c_291_n N_A_27_47#_c_784_n 0.00254621f $X=3.215 $Y=1.185
+ $X2=0 $Y2=0
cc_318 N_A_456_21#_c_286_n N_VGND_c_853_n 0.0131769f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_319 N_A_456_21#_c_287_n N_VGND_c_853_n 7.02169e-19 $X=2.71 $Y=1.26 $X2=0
+ $Y2=0
cc_320 N_A_456_21#_c_289_n N_VGND_c_853_n 0.0120044f $X=2.785 $Y=1.185 $X2=0
+ $Y2=0
cc_321 N_A_456_21#_c_291_n N_VGND_c_853_n 6.24795e-19 $X=3.215 $Y=1.185 $X2=0
+ $Y2=0
cc_322 N_A_456_21#_c_289_n N_VGND_c_854_n 5.68397e-19 $X=2.785 $Y=1.185 $X2=0
+ $Y2=0
cc_323 N_A_456_21#_c_291_n N_VGND_c_854_n 0.0086675f $X=3.215 $Y=1.185 $X2=0
+ $Y2=0
cc_324 N_A_456_21#_c_293_n N_VGND_c_854_n 0.00301179f $X=3.645 $Y=1.185 $X2=0
+ $Y2=0
cc_325 N_A_456_21#_c_300_n N_VGND_c_855_n 0.00499288f $X=5.025 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_A_456_21#_c_302_n N_VGND_c_855_n 0.0322245f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_327 N_A_456_21#_c_289_n N_VGND_c_856_n 0.00486043f $X=2.785 $Y=1.185 $X2=0
+ $Y2=0
cc_328 N_A_456_21#_c_291_n N_VGND_c_856_n 0.00486043f $X=3.215 $Y=1.185 $X2=0
+ $Y2=0
cc_329 N_A_456_21#_c_286_n N_VGND_c_858_n 0.00486043f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_330 N_A_456_21#_c_293_n N_VGND_c_859_n 0.0054895f $X=3.645 $Y=1.185 $X2=0
+ $Y2=0
cc_331 N_A_456_21#_c_301_n N_VGND_c_859_n 0.00577334f $X=4.36 $Y=0.505 $X2=0
+ $Y2=0
cc_332 N_A_456_21#_c_302_n N_VGND_c_859_n 0.0497316f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_333 N_A_456_21#_c_286_n N_VGND_c_861_n 0.0082726f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_334 N_A_456_21#_c_289_n N_VGND_c_861_n 0.00824727f $X=2.785 $Y=1.185 $X2=0
+ $Y2=0
cc_335 N_A_456_21#_c_291_n N_VGND_c_861_n 0.00454119f $X=3.215 $Y=1.185 $X2=0
+ $Y2=0
cc_336 N_A_456_21#_c_293_n N_VGND_c_861_n 0.00743132f $X=3.645 $Y=1.185 $X2=0
+ $Y2=0
cc_337 N_A_456_21#_c_301_n N_VGND_c_861_n 0.00394402f $X=4.36 $Y=0.505 $X2=0
+ $Y2=0
cc_338 N_A_456_21#_c_302_n N_VGND_c_861_n 0.0341779f $X=4.945 $Y=0.42 $X2=0
+ $Y2=0
cc_339 N_TE_B_M1002_g N_A_M1005_g 0.0443283f $X=5.16 $Y=2.465 $X2=0 $Y2=0
cc_340 N_TE_B_M1012_g N_A_M1019_g 0.0267001f $X=5.16 $Y=0.695 $X2=0 $Y2=0
cc_341 N_TE_B_c_406_n N_A_c_528_n 0.0168496f $X=5.16 $Y=1.34 $X2=0 $Y2=0
cc_342 N_TE_B_c_406_n N_A_c_529_n 0.00338335f $X=5.16 $Y=1.34 $X2=0 $Y2=0
cc_343 N_TE_B_c_410_n N_A_27_367#_c_578_n 0.00196648f $X=2.425 $Y=1.725 $X2=0
+ $Y2=0
cc_344 N_TE_B_c_410_n N_A_27_367#_c_580_n 7.32954e-19 $X=2.425 $Y=1.725 $X2=0
+ $Y2=0
cc_345 N_TE_B_c_410_n N_A_27_367#_c_589_n 0.00559687f $X=2.425 $Y=1.725 $X2=0
+ $Y2=0
cc_346 N_TE_B_c_413_n N_A_27_367#_c_589_n 5.7298e-19 $X=2.995 $Y=1.725 $X2=0
+ $Y2=0
cc_347 N_TE_B_c_410_n N_A_27_367#_c_582_n 0.0092802f $X=2.425 $Y=1.725 $X2=0
+ $Y2=0
cc_348 N_TE_B_c_413_n N_A_27_367#_c_582_n 0.0103085f $X=2.995 $Y=1.725 $X2=0
+ $Y2=0
cc_349 N_TE_B_c_415_n N_A_27_367#_c_565_n 0.0111934f $X=3.425 $Y=1.725 $X2=0
+ $Y2=0
cc_350 N_TE_B_c_417_n N_A_27_367#_c_565_n 0.0126717f $X=4.035 $Y=1.725 $X2=0
+ $Y2=0
cc_351 N_TE_B_M1002_g N_A_27_367#_c_565_n 0.00417418f $X=5.16 $Y=2.465 $X2=0
+ $Y2=0
cc_352 N_TE_B_c_415_n N_A_27_367#_c_566_n 8.03689e-19 $X=3.425 $Y=1.725 $X2=0
+ $Y2=0
cc_353 N_TE_B_c_417_n N_A_27_367#_c_566_n 0.00775012f $X=4.035 $Y=1.725 $X2=0
+ $Y2=0
cc_354 N_TE_B_M1002_g N_A_27_367#_c_566_n 0.00840863f $X=5.16 $Y=2.465 $X2=0
+ $Y2=0
cc_355 N_TE_B_c_410_n N_A_27_367#_c_586_n 6.89869e-19 $X=2.425 $Y=1.725 $X2=0
+ $Y2=0
cc_356 N_TE_B_c_413_n N_A_27_367#_c_586_n 0.0046808f $X=2.995 $Y=1.725 $X2=0
+ $Y2=0
cc_357 N_TE_B_c_415_n N_A_27_367#_c_586_n 0.00480362f $X=3.425 $Y=1.725 $X2=0
+ $Y2=0
cc_358 N_TE_B_c_417_n N_A_27_367#_c_586_n 0.00164053f $X=4.035 $Y=1.725 $X2=0
+ $Y2=0
cc_359 N_TE_B_c_413_n N_A_27_367#_c_603_n 0.00410591f $X=2.995 $Y=1.725 $X2=0
+ $Y2=0
cc_360 N_TE_B_c_415_n N_A_27_367#_c_603_n 0.00591537f $X=3.425 $Y=1.725 $X2=0
+ $Y2=0
cc_361 N_TE_B_c_410_n N_Z_c_645_n 8.62452e-19 $X=2.425 $Y=1.725 $X2=0 $Y2=0
cc_362 N_TE_B_c_410_n N_VPWR_c_705_n 0.00558836f $X=2.425 $Y=1.725 $X2=0 $Y2=0
cc_363 N_TE_B_c_413_n N_VPWR_c_705_n 0.00422823f $X=2.995 $Y=1.725 $X2=0 $Y2=0
cc_364 N_TE_B_c_413_n N_VPWR_c_706_n 0.0054895f $X=2.995 $Y=1.725 $X2=0 $Y2=0
cc_365 N_TE_B_c_415_n N_VPWR_c_706_n 0.00415375f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_366 N_TE_B_c_415_n N_VPWR_c_707_n 0.00335544f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_367 N_TE_B_c_417_n N_VPWR_c_707_n 0.00544694f $X=4.035 $Y=1.725 $X2=0 $Y2=0
cc_368 N_TE_B_M1002_g N_VPWR_c_708_n 0.0318086f $X=5.16 $Y=2.465 $X2=0 $Y2=0
cc_369 N_TE_B_c_417_n N_VPWR_c_709_n 0.00415375f $X=4.035 $Y=1.725 $X2=0 $Y2=0
cc_370 N_TE_B_M1002_g N_VPWR_c_709_n 0.00486043f $X=5.16 $Y=2.465 $X2=0 $Y2=0
cc_371 N_TE_B_c_410_n N_VPWR_c_711_n 0.00547432f $X=2.425 $Y=1.725 $X2=0 $Y2=0
cc_372 N_TE_B_c_410_n N_VPWR_c_704_n 0.00658744f $X=2.425 $Y=1.725 $X2=0 $Y2=0
cc_373 N_TE_B_c_413_n N_VPWR_c_704_n 0.00639337f $X=2.995 $Y=1.725 $X2=0 $Y2=0
cc_374 N_TE_B_c_415_n N_VPWR_c_704_n 0.0061249f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_375 N_TE_B_c_417_n N_VPWR_c_704_n 0.00770462f $X=4.035 $Y=1.725 $X2=0 $Y2=0
cc_376 N_TE_B_M1002_g N_VPWR_c_704_n 0.00975473f $X=5.16 $Y=2.465 $X2=0 $Y2=0
cc_377 N_TE_B_c_396_n N_A_27_47#_c_779_n 0.00377134f $X=2.5 $Y=1.65 $X2=0 $Y2=0
cc_378 N_TE_B_c_397_n N_A_27_47#_c_781_n 0.00141587f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_379 N_TE_B_c_409_n N_A_27_47#_c_781_n 0.0381494f $X=4.44 $Y=1.295 $X2=0 $Y2=0
cc_380 N_TE_B_c_395_n N_A_27_47#_c_784_n 0.00117276f $X=2.92 $Y=1.65 $X2=0 $Y2=0
cc_381 N_TE_B_c_409_n N_A_27_47#_c_784_n 0.00476161f $X=4.44 $Y=1.295 $X2=0
+ $Y2=0
cc_382 N_TE_B_M1012_g N_VGND_c_855_n 0.0081345f $X=5.16 $Y=0.695 $X2=0 $Y2=0
cc_383 N_TE_B_M1012_g N_VGND_c_859_n 0.00509933f $X=5.16 $Y=0.695 $X2=0 $Y2=0
cc_384 N_TE_B_M1012_g N_VGND_c_861_n 0.0107152f $X=5.16 $Y=0.695 $X2=0 $Y2=0
cc_385 N_A_M1005_g N_VPWR_c_708_n 0.0060347f $X=5.66 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A_M1005_g N_VPWR_c_712_n 0.0054895f $X=5.66 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A_M1005_g N_VPWR_c_704_n 0.0110901f $X=5.66 $Y=2.465 $X2=0 $Y2=0
cc_388 N_A_M1019_g N_VGND_c_855_n 0.00813484f $X=5.73 $Y=0.695 $X2=0 $Y2=0
cc_389 N_A_c_528_n N_VGND_c_855_n 0.00103097f $X=5.64 $Y=1.51 $X2=0 $Y2=0
cc_390 N_A_c_529_n N_VGND_c_855_n 0.0152531f $X=5.64 $Y=1.51 $X2=0 $Y2=0
cc_391 N_A_M1019_g N_VGND_c_860_n 0.00511358f $X=5.73 $Y=0.695 $X2=0 $Y2=0
cc_392 N_A_M1019_g N_VGND_c_861_n 0.0104941f $X=5.73 $Y=0.695 $X2=0 $Y2=0
cc_393 N_A_27_367#_c_574_n N_Z_M1001_d 0.00332344f $X=1.045 $Y=2.99 $X2=0 $Y2=0
cc_394 N_A_27_367#_c_578_n N_Z_M1011_d 0.00472489f $X=2.045 $Y=2.99 $X2=0 $Y2=0
cc_395 N_A_27_367#_M1006_s N_Z_c_643_n 0.00250873f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_396 N_A_27_367#_c_576_n N_Z_c_643_n 0.0209867f $X=1.21 $Y=2.24 $X2=0 $Y2=0
cc_397 N_A_27_367#_c_564_n N_Z_c_641_n 0.0112876f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_398 N_A_27_367#_c_564_n N_Z_c_644_n 0.00792225f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_399 N_A_27_367#_c_574_n N_Z_c_644_n 0.016693f $X=1.045 $Y=2.99 $X2=0 $Y2=0
cc_400 N_A_27_367#_c_578_n N_Z_c_645_n 0.0196355f $X=2.045 $Y=2.99 $X2=0 $Y2=0
cc_401 N_A_27_367#_c_582_n N_VPWR_M1007_s 0.0068165f $X=3.045 $Y=2.44 $X2=-0.19
+ $Y2=1.655
cc_402 N_A_27_367#_c_565_n N_VPWR_M1016_s 0.0097573f $X=4.085 $Y=2.61 $X2=0
+ $Y2=0
cc_403 N_A_27_367#_c_582_n N_VPWR_c_705_n 0.0243897f $X=3.045 $Y=2.44 $X2=0
+ $Y2=0
cc_404 N_A_27_367#_c_565_n N_VPWR_c_706_n 0.00247188f $X=4.085 $Y=2.61 $X2=0
+ $Y2=0
cc_405 N_A_27_367#_c_603_n N_VPWR_c_706_n 0.018986f $X=3.21 $Y=2.61 $X2=0 $Y2=0
cc_406 N_A_27_367#_c_565_n N_VPWR_c_707_n 0.0241666f $X=4.085 $Y=2.61 $X2=0
+ $Y2=0
cc_407 N_A_27_367#_c_566_n N_VPWR_c_707_n 0.0138561f $X=4.25 $Y=2.8 $X2=0 $Y2=0
cc_408 N_A_27_367#_c_565_n N_VPWR_c_709_n 0.00307177f $X=4.085 $Y=2.61 $X2=0
+ $Y2=0
cc_409 N_A_27_367#_c_566_n N_VPWR_c_709_n 0.0207593f $X=4.25 $Y=2.8 $X2=0 $Y2=0
cc_410 N_A_27_367#_c_563_n N_VPWR_c_711_n 0.017536f $X=0.24 $Y=2.905 $X2=0 $Y2=0
cc_411 N_A_27_367#_c_574_n N_VPWR_c_711_n 0.0364961f $X=1.045 $Y=2.99 $X2=0
+ $Y2=0
cc_412 N_A_27_367#_c_578_n N_VPWR_c_711_n 0.0582459f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_413 N_A_27_367#_c_585_n N_VPWR_c_711_n 0.0207136f $X=1.21 $Y=2.95 $X2=0 $Y2=0
cc_414 N_A_27_367#_M1001_s N_VPWR_c_704_n 0.00231918f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_415 N_A_27_367#_M1006_s N_VPWR_c_704_n 0.00280658f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_416 N_A_27_367#_M1015_s N_VPWR_c_704_n 0.00280658f $X=2 $Y=1.835 $X2=0 $Y2=0
cc_417 N_A_27_367#_M1009_d N_VPWR_c_704_n 0.00223559f $X=3.07 $Y=1.835 $X2=0
+ $Y2=0
cc_418 N_A_27_367#_M1017_d N_VPWR_c_704_n 0.00232718f $X=4.11 $Y=1.835 $X2=0
+ $Y2=0
cc_419 N_A_27_367#_c_563_n N_VPWR_c_704_n 0.00970886f $X=0.24 $Y=2.905 $X2=0
+ $Y2=0
cc_420 N_A_27_367#_c_574_n N_VPWR_c_704_n 0.0241226f $X=1.045 $Y=2.99 $X2=0
+ $Y2=0
cc_421 N_A_27_367#_c_578_n N_VPWR_c_704_n 0.0365877f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_422 N_A_27_367#_c_582_n N_VPWR_c_704_n 0.0113978f $X=3.045 $Y=2.44 $X2=0
+ $Y2=0
cc_423 N_A_27_367#_c_565_n N_VPWR_c_704_n 0.011108f $X=4.085 $Y=2.61 $X2=0 $Y2=0
cc_424 N_A_27_367#_c_566_n N_VPWR_c_704_n 0.0125721f $X=4.25 $Y=2.8 $X2=0 $Y2=0
cc_425 N_A_27_367#_c_585_n N_VPWR_c_704_n 0.0126421f $X=1.21 $Y=2.95 $X2=0 $Y2=0
cc_426 N_A_27_367#_c_603_n N_VPWR_c_704_n 0.012405f $X=3.21 $Y=2.61 $X2=0 $Y2=0
cc_427 N_Z_M1001_d N_VPWR_c_704_n 0.00225186f $X=0.57 $Y=1.835 $X2=0 $Y2=0
cc_428 N_Z_M1011_d N_VPWR_c_704_n 0.00281482f $X=1.5 $Y=1.835 $X2=0 $Y2=0
cc_429 N_Z_c_640_n N_A_27_47#_M1003_s 0.00250873f $X=1.545 $Y=1.06 $X2=0 $Y2=0
cc_430 N_Z_M1000_d N_A_27_47#_c_785_n 0.00332344f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_431 N_Z_c_646_n N_A_27_47#_c_785_n 0.016631f $X=0.71 $Y=0.805 $X2=0 $Y2=0
cc_432 N_Z_c_640_n N_A_27_47#_c_785_n 0.00321827f $X=1.545 $Y=1.06 $X2=0 $Y2=0
cc_433 N_Z_M1004_d N_A_27_47#_c_787_n 0.00472489f $X=1.5 $Y=0.235 $X2=0 $Y2=0
cc_434 N_Z_c_640_n N_A_27_47#_c_787_n 0.00321827f $X=1.545 $Y=1.06 $X2=0 $Y2=0
cc_435 N_Z_c_668_n N_A_27_47#_c_787_n 0.0193546f $X=1.71 $Y=0.805 $X2=0 $Y2=0
cc_436 N_Z_c_640_n N_A_27_47#_c_778_n 0.00854023f $X=1.545 $Y=1.06 $X2=0 $Y2=0
cc_437 N_Z_c_640_n N_A_27_47#_c_780_n 8.53482e-19 $X=1.545 $Y=1.06 $X2=0 $Y2=0
cc_438 N_Z_c_641_n N_A_27_47#_c_783_n 0.0201602f $X=0.535 $Y=1.295 $X2=0 $Y2=0
cc_439 N_Z_c_640_n N_A_27_47#_c_792_n 0.0206278f $X=1.545 $Y=1.06 $X2=0 $Y2=0
cc_440 N_Z_M1000_d N_VGND_c_861_n 0.00225186f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_441 N_Z_M1004_d N_VGND_c_861_n 0.00281482f $X=1.5 $Y=0.235 $X2=0 $Y2=0
cc_442 N_A_27_47#_c_781_n N_VGND_M1013_d 0.00379369f $X=3.695 $Y=0.925 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_779_n N_VGND_c_853_n 0.0216086f $X=2.915 $Y=1.22 $X2=0 $Y2=0
cc_444 N_A_27_47#_c_781_n N_VGND_c_854_n 0.0149979f $X=3.695 $Y=0.925 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_833_p N_VGND_c_856_n 0.0117428f $X=3 $Y=0.42 $X2=0 $Y2=0
cc_446 N_A_27_47#_c_785_n N_VGND_c_858_n 0.0364961f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_447 N_A_27_47#_c_787_n N_VGND_c_858_n 0.037782f $X=2.055 $Y=0.34 $X2=0 $Y2=0
cc_448 N_A_27_47#_c_836_p N_VGND_c_858_n 0.0118138f $X=2.14 $Y=0.425 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_783_n N_VGND_c_858_n 0.017536f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_450 N_A_27_47#_c_792_n N_VGND_c_858_n 0.020435f $X=1.21 $Y=0.38 $X2=0 $Y2=0
cc_451 N_A_27_47#_c_782_n N_VGND_c_859_n 0.0210192f $X=3.86 $Y=0.42 $X2=0 $Y2=0
cc_452 N_A_27_47#_M1000_s N_VGND_c_861_n 0.00231918f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_M1003_s N_VGND_c_861_n 0.00280658f $X=1 $Y=0.235 $X2=0 $Y2=0
cc_454 N_A_27_47#_M1018_s N_VGND_c_861_n 0.00411415f $X=2 $Y=0.235 $X2=0 $Y2=0
cc_455 N_A_27_47#_M1010_s N_VGND_c_861_n 0.00449904f $X=2.86 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_M1014_s N_VGND_c_861_n 0.00231914f $X=3.72 $Y=0.235 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_785_n N_VGND_c_861_n 0.0241226f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_458 N_A_27_47#_c_787_n N_VGND_c_861_n 0.024237f $X=2.055 $Y=0.34 $X2=0 $Y2=0
cc_459 N_A_27_47#_c_836_p N_VGND_c_861_n 0.00658808f $X=2.14 $Y=0.425 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_833_p N_VGND_c_861_n 0.00652089f $X=3 $Y=0.42 $X2=0 $Y2=0
cc_461 N_A_27_47#_c_781_n N_VGND_c_861_n 0.0113364f $X=3.695 $Y=0.925 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_782_n N_VGND_c_861_n 0.0125689f $X=3.86 $Y=0.42 $X2=0 $Y2=0
cc_463 N_A_27_47#_c_783_n N_VGND_c_861_n 0.00970886f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_464 N_A_27_47#_c_792_n N_VGND_c_861_n 0.0125725f $X=1.21 $Y=0.38 $X2=0 $Y2=0
