* File: sky130_fd_sc_lp__dfxtp_1.pex.spice
* Created: Fri Aug 28 10:24:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFXTP_1%CLK 2 7 11 13 14 15 16 17 18 19 25
r32 25 27 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.12
+ $X2=0.352 $Y2=0.955
r33 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.12 $X2=0.32 $Y2=1.12
r34 18 19 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r35 17 18 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r36 17 26 5.93169 $w=3.38e-07 $l=1.75e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.12
r37 16 26 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.12
r38 14 15 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=0.442 $Y=1.865
+ $X2=0.442 $Y2=2.015
r39 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.41 $Y=1.625
+ $X2=0.41 $Y2=1.865
r40 11 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.475 $Y=2.66
+ $X2=0.475 $Y2=2.015
r41 7 27 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.955
r42 2 13 42.4059 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.352 $Y=1.428
+ $X2=0.352 $Y2=1.625
r43 1 25 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.352 $Y=1.152
+ $X2=0.352 $Y2=1.12
r44 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.352 $Y=1.152
+ $X2=0.352 $Y2=1.428
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%D 3 5 7 8 9 17
c40 17 0 2.08001e-19 $X=2.195 $Y=1.51
r41 16 17 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.125 $Y=1.51
+ $X2=2.195 $Y2=1.51
r42 13 16 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.99 $Y=1.51
+ $X2=2.125 $Y2=1.51
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.51 $X2=1.99 $Y2=1.51
r44 9 14 3.7453 $w=4.93e-07 $l=1.55e-07 $layer=LI1_cond $X=1.827 $Y=1.665
+ $X2=1.827 $Y2=1.51
r45 8 14 5.19509 $w=4.93e-07 $l=2.15e-07 $layer=LI1_cond $X=1.827 $Y=1.295
+ $X2=1.827 $Y2=1.51
r46 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=1.51
r47 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=1.025
r48 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.125 $Y=1.675
+ $X2=2.125 $Y2=1.51
r49 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.125 $Y=1.675 $X2=2.125
+ $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%A_217_413# 1 2 9 13 17 19 20 23 27 31 33 36
+ 37 38 41 42 44 47 48 49 50 51 52 53
c163 42 0 1.13262e-19 $X=2.69 $Y=1.74
c164 41 0 7.86011e-20 $X=2.69 $Y=1.74
c165 31 0 1.294e-19 $X=1.325 $Y=1.02
r166 56 60 18.0931 $w=3.33e-07 $l=1.25e-07 $layer=POLY_cond $X=4.94 $Y=1.365
+ $X2=4.815 $Y2=1.365
r167 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.94
+ $Y=1.36 $X2=4.94 $Y2=1.36
r168 50 55 13.6938 $w=2.2e-07 $l=2.59702e-07 $layer=LI1_cond $X=4.845 $Y=1.595
+ $X2=4.897 $Y2=1.36
r169 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.845 $Y=1.595
+ $X2=4.845 $Y2=2.285
r170 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.76 $Y=2.37
+ $X2=4.845 $Y2=2.285
r171 48 49 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=4.76 $Y=2.37
+ $X2=3.495 $Y2=2.37
r172 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=2.455
+ $X2=3.495 $Y2=2.37
r173 46 47 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.41 $Y=2.455
+ $X2=3.41 $Y2=2.605
r174 45 53 3.58391 $w=2.75e-07 $l=9e-08 $layer=LI1_cond $X=2.775 $Y=2.742
+ $X2=2.685 $Y2=2.742
r175 44 47 7.32204 $w=2.75e-07 $l=1.74396e-07 $layer=LI1_cond $X=3.325 $Y=2.742
+ $X2=3.41 $Y2=2.605
r176 44 45 23.0489 $w=2.73e-07 $l=5.5e-07 $layer=LI1_cond $X=3.325 $Y=2.742
+ $X2=2.775 $Y2=2.742
r177 42 57 25.7194 $w=2.53e-07 $l=1.35e-07 $layer=POLY_cond $X=2.69 $Y=1.74
+ $X2=2.555 $Y2=1.74
r178 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.74 $X2=2.69 $Y2=1.74
r179 39 53 2.90466 $w=1.8e-07 $l=1.37e-07 $layer=LI1_cond $X=2.685 $Y=2.605
+ $X2=2.685 $Y2=2.742
r180 39 41 53.298 $w=1.78e-07 $l=8.65e-07 $layer=LI1_cond $X=2.685 $Y=2.605
+ $X2=2.685 $Y2=1.74
r181 37 53 3.58391 $w=2.75e-07 $l=9e-08 $layer=LI1_cond $X=2.595 $Y=2.742
+ $X2=2.685 $Y2=2.742
r182 37 38 21.7916 $w=2.73e-07 $l=5.2e-07 $layer=LI1_cond $X=2.595 $Y=2.742
+ $X2=2.075 $Y2=2.742
r183 36 38 7.32204 $w=2.75e-07 $l=1.74396e-07 $layer=LI1_cond $X=1.99 $Y=2.605
+ $X2=2.075 $Y2=2.742
r184 35 36 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.99 $Y=2.13
+ $X2=1.99 $Y2=2.605
r185 34 52 2.9446 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=1.41 $Y=2.045
+ $X2=1.045 $Y2=2.045
r186 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.905 $Y=2.045
+ $X2=1.99 $Y2=2.13
r187 33 34 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.905 $Y=2.045
+ $X2=1.41 $Y2=2.045
r188 29 52 3.55013 $w=2.62e-07 $l=2.89396e-07 $layer=LI1_cond $X=1.295 $Y=1.96
+ $X2=1.045 $Y2=2.045
r189 29 31 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.295 $Y=1.96
+ $X2=1.295 $Y2=1.02
r190 25 52 3.55013 $w=2.62e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.192 $Y=2.13
+ $X2=1.045 $Y2=2.045
r191 25 27 3.12527 $w=2.93e-07 $l=8e-08 $layer=LI1_cond $X=1.192 $Y=2.13
+ $X2=1.192 $Y2=2.21
r192 21 23 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.505 $Y=1.535
+ $X2=5.505 $Y2=2.105
r193 20 56 48.7533 $w=3.33e-07 $l=2.78478e-07 $layer=POLY_cond $X=5.175 $Y=1.46
+ $X2=4.94 $Y2=1.365
r194 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.43 $Y=1.46
+ $X2=5.505 $Y2=1.535
r195 19 20 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.43 $Y=1.46
+ $X2=5.175 $Y2=1.46
r196 15 60 21.4384 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.815 $Y=1.195
+ $X2=4.815 $Y2=1.365
r197 15 17 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.815 $Y=1.195
+ $X2=4.815 $Y2=0.805
r198 11 42 69.5376 $w=2.53e-07 $l=4.39829e-07 $layer=POLY_cond $X=3.055 $Y=1.575
+ $X2=2.69 $Y2=1.74
r199 11 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.055 $Y=1.575
+ $X2=3.055 $Y2=1.025
r200 7 57 14.9957 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.555 $Y=1.905
+ $X2=2.555 $Y2=1.74
r201 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.555 $Y=1.905
+ $X2=2.555 $Y2=2.275
r202 2 27 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.065 $X2=1.21 $Y2=2.21
r203 1 31 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.815 $X2=1.325 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%A_668_137# 1 2 9 13 17 18 20 21 24 29 30
c74 17 0 1.13262e-19 $X=3.535 $Y=1.53
r75 29 32 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.495 $Y=1.855
+ $X2=4.495 $Y2=1.985
r76 29 30 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.495 $Y=1.855
+ $X2=4.495 $Y2=1.245
r77 24 27 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=4.547 $Y=0.74
+ $X2=4.547 $Y2=1.08
r78 22 30 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=4.547 $Y=1.108
+ $X2=4.547 $Y2=1.245
r79 22 27 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=4.547 $Y=1.108
+ $X2=4.547 $Y2=1.08
r80 20 32 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.41 $Y=1.985
+ $X2=4.495 $Y2=1.985
r81 20 21 31.4706 $w=2.58e-07 $l=7.1e-07 $layer=LI1_cond $X=4.41 $Y=1.985
+ $X2=3.7 $Y2=1.985
r82 18 35 12.2413 $w=3.15e-07 $l=8e-08 $layer=POLY_cond $X=3.535 $Y=1.53
+ $X2=3.615 $Y2=1.53
r83 18 33 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=3.535 $Y=1.53
+ $X2=3.415 $Y2=1.53
r84 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.535
+ $Y=1.53 $X2=3.535 $Y2=1.53
r85 15 21 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=3.535 $Y=1.855
+ $X2=3.7 $Y2=1.985
r86 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.535 $Y=1.855
+ $X2=3.535 $Y2=1.53
r87 11 35 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.615 $Y=1.695
+ $X2=3.615 $Y2=1.53
r88 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.615 $Y=1.695
+ $X2=3.615 $Y2=2.275
r89 7 33 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.365
+ $X2=3.415 $Y2=1.53
r90 7 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.415 $Y=1.365
+ $X2=3.415 $Y2=1.025
r91 2 32 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.895 $X2=4.415 $Y2=2.02
r92 1 27 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=4.4
+ $Y=0.595 $X2=4.54 $Y2=1.08
r93 1 24 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=4.4
+ $Y=0.595 $X2=4.57 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%A_526_413# 1 2 9 11 13 16 18 19 22 31
r72 30 31 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=4.2 $Y=1.51
+ $X2=4.325 $Y2=1.51
r73 26 27 7.19663 $w=3.56e-07 $l=2.1e-07 $layer=LI1_cond $X=2.84 $Y=1.067
+ $X2=3.05 $Y2=1.067
r74 23 30 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.145 $Y=1.51
+ $X2=4.2 $Y2=1.51
r75 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=1.51 $X2=4.145 $Y2=1.51
r76 20 22 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=4.11 $Y=1.275
+ $X2=4.11 $Y2=1.51
r77 19 27 6.94352 $w=3.56e-07 $l=1.67463e-07 $layer=LI1_cond $X=3.155 $Y=1.19
+ $X2=3.05 $Y2=1.067
r78 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.98 $Y=1.19
+ $X2=4.11 $Y2=1.275
r79 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.98 $Y=1.19
+ $X2=3.155 $Y2=1.19
r80 14 27 3.82529 $w=2.1e-07 $l=2.08e-07 $layer=LI1_cond $X=3.05 $Y=1.275
+ $X2=3.05 $Y2=1.067
r81 14 16 52.5498 $w=2.08e-07 $l=9.95e-07 $layer=LI1_cond $X=3.05 $Y=1.275
+ $X2=3.05 $Y2=2.27
r82 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.325 $Y=1.345
+ $X2=4.325 $Y2=1.51
r83 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.325 $Y=1.345
+ $X2=4.325 $Y2=0.915
r84 7 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.2 $Y=1.675 $X2=4.2
+ $Y2=1.51
r85 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.2 $Y=1.675 $X2=4.2
+ $Y2=2.315
r86 2 16 600 $w=1.7e-07 $l=4.91935e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=2.065 $X2=3.03 $Y2=2.27
r87 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.815 $X2=2.84 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%A_110_70# 1 2 7 8 12 16 17 18 19 20 23 25 29
+ 31 35 39 43 45 46 49 52 55 58 59 61
c140 16 0 1.84694e-19 $X=1.54 $Y=1.025
r141 58 60 6.18117 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.802 $Y=1.12
+ $X2=0.802 $Y2=0.955
r142 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.12 $X2=0.925 $Y2=1.12
r143 55 61 47.6909 $w=1.98e-07 $l=8.6e-07 $layer=LI1_cond $X=0.695 $Y=2.485
+ $X2=0.695 $Y2=1.625
r144 52 61 8.85186 $w=4.13e-07 $l=2.07e-07 $layer=LI1_cond $X=0.802 $Y=1.418
+ $X2=0.802 $Y2=1.625
r145 51 58 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=0.802 $Y=1.162
+ $X2=0.802 $Y2=1.12
r146 51 52 7.10905 $w=4.13e-07 $l=2.56e-07 $layer=LI1_cond $X=0.802 $Y=1.162
+ $X2=0.802 $Y2=1.418
r147 49 60 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.725 $Y=0.565
+ $X2=0.725 $Y2=0.955
r148 42 43 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.425 $Y=1.55
+ $X2=1.54 $Y2=1.55
r149 41 59 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.925 $Y=1.475
+ $X2=0.925 $Y2=1.12
r150 37 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.505 $Y=0.255
+ $X2=5.505 $Y2=0.805
r151 33 35 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.71 $Y=3.075
+ $X2=4.71 $Y2=2.315
r152 32 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.33 $Y=3.15
+ $X2=3.255 $Y2=3.15
r153 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.635 $Y=3.15
+ $X2=4.71 $Y2=3.075
r154 31 32 669.16 $w=1.5e-07 $l=1.305e-06 $layer=POLY_cond $X=4.635 $Y=3.15
+ $X2=3.33 $Y2=3.15
r155 27 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=3.075
+ $X2=3.255 $Y2=3.15
r156 27 29 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.255 $Y=3.075
+ $X2=3.255 $Y2=2.275
r157 26 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=0.18
+ $X2=2.625 $Y2=0.18
r158 25 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.43 $Y=0.18
+ $X2=5.505 $Y2=0.255
r159 25 26 1399.85 $w=1.5e-07 $l=2.73e-06 $layer=POLY_cond $X=5.43 $Y=0.18
+ $X2=2.7 $Y2=0.18
r160 21 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=0.255
+ $X2=2.625 $Y2=0.18
r161 21 23 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.625 $Y=0.255
+ $X2=2.625 $Y2=1.025
r162 19 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=0.18
+ $X2=2.625 $Y2=0.18
r163 19 20 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=2.55 $Y=0.18
+ $X2=1.615 $Y2=0.18
r164 17 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=3.15
+ $X2=3.255 $Y2=3.15
r165 17 18 861.447 $w=1.5e-07 $l=1.68e-06 $layer=POLY_cond $X=3.18 $Y=3.15
+ $X2=1.5 $Y2=3.15
r166 14 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.54 $Y=1.475
+ $X2=1.54 $Y2=1.55
r167 14 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.54 $Y=1.475
+ $X2=1.54 $Y2=1.025
r168 13 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.54 $Y=0.255
+ $X2=1.615 $Y2=0.18
r169 13 16 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.54 $Y=0.255
+ $X2=1.54 $Y2=1.025
r170 10 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.425 $Y=3.075
+ $X2=1.5 $Y2=3.15
r171 10 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.425 $Y=3.075
+ $X2=1.425 $Y2=2.385
r172 9 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=1.625
+ $X2=1.425 $Y2=1.55
r173 9 12 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.425 $Y=1.625
+ $X2=1.425 $Y2=2.385
r174 8 41 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.09 $Y=1.55
+ $X2=0.925 $Y2=1.475
r175 7 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.35 $Y=1.55
+ $X2=1.425 $Y2=1.55
r176 7 8 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.35 $Y=1.55 $X2=1.09
+ $Y2=1.55
r177 2 55 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.34 $X2=0.69 $Y2=2.485
r178 1 49 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.35 $X2=0.69 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%A_1158_93# 1 2 9 13 15 17 21 23 25 27 32 33
+ 42
r72 42 43 7.03628 $w=4.3e-07 $l=2.48e-07 $layer=LI1_cond $X=6.822 $Y=1.462
+ $X2=6.822 $Y2=1.71
r73 40 42 8.85209 $w=4.3e-07 $l=3.12e-07 $layer=LI1_cond $X=6.822 $Y=1.15
+ $X2=6.822 $Y2=1.462
r74 40 41 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=7.04
+ $Y=1.15 $X2=7.04 $Y2=1.15
r75 38 40 17.8744 $w=4.3e-07 $l=6.3e-07 $layer=LI1_cond $X=6.822 $Y=0.52
+ $X2=6.822 $Y2=1.15
r76 33 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.57
+ $X2=5.955 $Y2=1.735
r77 33 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.57
+ $X2=5.955 $Y2=1.405
r78 32 35 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.955 $Y=1.57
+ $X2=5.955 $Y2=1.71
r79 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.955
+ $Y=1.57 $X2=5.955 $Y2=1.57
r80 25 43 2.51413 $w=4.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.737 $Y=1.795
+ $X2=6.822 $Y2=1.71
r81 25 27 7.14806 $w=3.93e-07 $l=2.45e-07 $layer=LI1_cond $X=6.737 $Y=1.795
+ $X2=6.737 $Y2=2.04
r82 24 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.12 $Y=1.71
+ $X2=5.955 $Y2=1.71
r83 23 43 6.22023 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=6.54 $Y=1.71
+ $X2=6.822 $Y2=1.71
r84 23 24 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6.54 $Y=1.71
+ $X2=6.12 $Y2=1.71
r85 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.685 $Y=1.655
+ $X2=7.685 $Y2=2.465
r86 15 19 32.2548 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.685 $Y=1.32
+ $X2=7.685 $Y2=1.655
r87 15 41 60.1335 $w=5.17e-07 $l=6.45e-07 $layer=POLY_cond $X=7.685 $Y=1.32
+ $X2=7.04 $Y2=1.32
r88 15 17 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=7.685 $Y=1.25
+ $X2=7.685 $Y2=0.655
r89 13 46 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.865 $Y=2.105
+ $X2=5.865 $Y2=1.735
r90 9 45 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.865 $Y=0.805 $X2=5.865
+ $Y2=1.405
r91 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.485
+ $Y=1.895 $X2=6.625 $Y2=2.04
r92 1 38 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=6.445
+ $Y=0.375 $X2=6.64 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%A_957_379# 1 2 7 9 10 12 14 16 21 24 29 31
+ 32 33
c78 24 0 3.01023e-20 $X=6.335 $Y=1.21
r79 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.5
+ $Y=1.29 $X2=6.5 $Y2=1.29
r80 33 36 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=6.465 $Y=1.21
+ $X2=6.465 $Y2=1.29
r81 27 29 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.155 $Y=0.805
+ $X2=5.3 $Y2=0.805
r82 25 32 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.395 $Y=1.21 $X2=5.3
+ $Y2=1.21
r83 24 33 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.335 $Y=1.21
+ $X2=6.465 $Y2=1.21
r84 24 25 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.335 $Y=1.21
+ $X2=5.395 $Y2=1.21
r85 22 32 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=5.29 $Y=1.295
+ $X2=5.3 $Y2=1.21
r86 22 31 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=5.29 $Y=1.295
+ $X2=5.29 $Y2=1.875
r87 21 32 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=1.125 $X2=5.3
+ $Y2=1.21
r88 20 29 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=0.97 $X2=5.3
+ $Y2=0.805
r89 20 21 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=5.3 $Y=0.97 $X2=5.3
+ $Y2=1.125
r90 16 18 23.9186 $w=2.63e-07 $l=5.5e-07 $layer=LI1_cond $X=5.242 $Y=2.04
+ $X2=5.242 $Y2=2.59
r91 14 31 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=5.242 $Y=2.007
+ $X2=5.242 $Y2=1.875
r92 14 16 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=5.242 $Y=2.007
+ $X2=5.242 $Y2=2.04
r93 10 37 38.6889 $w=3.41e-07 $l=1.96914e-07 $layer=POLY_cond $X=6.41 $Y=1.455
+ $X2=6.48 $Y2=1.29
r94 10 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.41 $Y=1.455
+ $X2=6.41 $Y2=2.315
r95 7 37 43.6361 $w=3.41e-07 $l=2.48998e-07 $layer=POLY_cond $X=6.37 $Y=1.09
+ $X2=6.48 $Y2=1.29
r96 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.37 $Y=1.09 $X2=6.37
+ $Y2=0.695
r97 2 18 600 $w=1.7e-07 $l=8.76342e-07 $layer=licon1_PDIFF $count=1 $X=4.785
+ $Y=1.895 $X2=5.195 $Y2=2.59
r98 2 16 600 $w=1.7e-07 $l=4.77022e-07 $layer=licon1_PDIFF $count=1 $X=4.785
+ $Y=1.895 $X2=5.195 $Y2=2.04
r99 1 27 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.595 $X2=5.155 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%VPWR 1 2 3 4 5 16 18 22 26 28 32 38 42 44 49
+ 54 61 62 68 71 74 77
c87 32 0 3.01023e-20 $X=6.145 $Y=2.05
r88 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r89 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r90 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 62 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r93 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r94 59 77 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.605 $Y=3.33
+ $X2=7.455 $Y2=3.33
r95 59 61 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.605 $Y=3.33
+ $X2=7.92 $Y2=3.33
r96 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r97 58 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33 $X2=6
+ $Y2=3.33
r98 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r99 55 74 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.36 $Y=3.33 $X2=6.17
+ $Y2=3.33
r100 55 57 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.36 $Y=3.33 $X2=6.96
+ $Y2=3.33
r101 54 77 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.305 $Y=3.33
+ $X2=7.455 $Y2=3.33
r102 54 57 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.305 $Y=3.33
+ $X2=6.96 $Y2=3.33
r103 53 69 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 50 68 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.622 $Y2=3.33
r106 50 52 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=3.6 $Y2=3.33
r107 49 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.925 $Y2=3.33
r108 49 52 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.6 $Y2=3.33
r109 48 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 48 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r111 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 45 65 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r113 45 47 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 44 68 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.51 $Y=3.33
+ $X2=1.622 $Y2=3.33
r115 44 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.51 $Y=3.33
+ $X2=1.2 $Y2=3.33
r116 42 75 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r117 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r118 42 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r119 38 41 36.8782 $w=2.98e-07 $l=9.6e-07 $layer=LI1_cond $X=7.455 $Y=1.99
+ $X2=7.455 $Y2=2.95
r120 36 77 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.455 $Y=3.245
+ $X2=7.455 $Y2=3.33
r121 36 41 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=7.455 $Y=3.245
+ $X2=7.455 $Y2=2.95
r122 32 35 16.9834 $w=3.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.17 $Y=2.05
+ $X2=6.17 $Y2=2.61
r123 30 74 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=3.245
+ $X2=6.17 $Y2=3.33
r124 30 35 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=6.17 $Y=3.245
+ $X2=6.17 $Y2=2.61
r125 29 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=3.33
+ $X2=3.925 $Y2=3.33
r126 28 74 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=6.17 $Y2=3.33
r127 28 29 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=4.09 $Y2=3.33
r128 24 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=3.245
+ $X2=3.925 $Y2=3.33
r129 24 26 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.925 $Y=3.245
+ $X2=3.925 $Y2=2.72
r130 20 68 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.622 $Y=3.245
+ $X2=1.622 $Y2=3.33
r131 20 22 39.9514 $w=2.23e-07 $l=7.8e-07 $layer=LI1_cond $X=1.622 $Y=3.245
+ $X2=1.622 $Y2=2.465
r132 16 65 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r133 16 18 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.49
r134 5 41 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=7.345
+ $Y=1.835 $X2=7.47 $Y2=2.95
r135 5 38 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=7.345
+ $Y=1.835 $X2=7.47 $Y2=1.99
r136 4 35 600 $w=1.7e-07 $l=8.32797e-07 $layer=licon1_PDIFF $count=1 $X=5.94
+ $Y=1.895 $X2=6.195 $Y2=2.61
r137 4 32 600 $w=1.7e-07 $l=2.71662e-07 $layer=licon1_PDIFF $count=1 $X=5.94
+ $Y=1.895 $X2=6.145 $Y2=2.05
r138 3 26 600 $w=1.7e-07 $l=7.63512e-07 $layer=licon1_PDIFF $count=1 $X=3.69
+ $Y=2.065 $X2=3.925 $Y2=2.72
r139 2 22 600 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=2.065 $X2=1.64 $Y2=2.465
r140 1 18 300 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.34 $X2=0.26 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%A_440_413# 1 2 9 12
c21 9 0 1.84694e-19 $X=2.34 $Y=2.27
r22 12 14 8.12648 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=1.025
+ $X2=2.41 $Y2=1.19
r23 9 14 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=2.335 $Y=2.27
+ $X2=2.335 $Y2=1.19
r24 2 9 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=2.065 $X2=2.34 $Y2=2.27
r25 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.815 $X2=2.41 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%Q 1 2 7 8 9 10 11 12 13 22
r13 13 40 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=2.775
+ $X2=7.92 $Y2=2.91
r14 12 13 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=2.405
+ $X2=7.92 $Y2=2.775
r15 11 12 15.4984 $w=2.88e-07 $l=3.9e-07 $layer=LI1_cond $X=7.92 $Y=2.015
+ $X2=7.92 $Y2=2.405
r16 10 11 13.9088 $w=2.88e-07 $l=3.5e-07 $layer=LI1_cond $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=2.015
r17 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=1.295
+ $X2=7.92 $Y2=1.665
r18 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=0.925 $X2=7.92
+ $Y2=1.295
r19 7 8 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=0.555 $X2=7.92
+ $Y2=0.925
r20 7 22 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=0.555
+ $X2=7.92 $Y2=0.42
r21 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.835 $X2=7.9 $Y2=2.91
r22 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=7.76 $Y=1.835
+ $X2=7.9 $Y2=2.015
r23 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.76
+ $Y=0.235 $X2=7.9 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_1%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 39 48
+ 52 57 64 65 71 76 79
r79 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r80 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r81 71 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r82 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r84 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r85 62 79 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=7.605 $Y=0 $X2=7.472
+ $Y2=0
r86 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.605 $Y=0 $X2=7.92
+ $Y2=0
r87 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r88 61 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6
+ $Y2=0
r89 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r90 58 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6.14
+ $Y2=0
r91 58 60 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6.96
+ $Y2=0
r92 57 79 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.34 $Y=0 $X2=7.472
+ $Y2=0
r93 57 60 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.34 $Y=0 $X2=6.96
+ $Y2=0
r94 56 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r95 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 53 71 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=3.905
+ $Y2=0
r97 53 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.56
+ $Y2=0
r98 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=0 $X2=6.14
+ $Y2=0
r99 52 55 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=5.975 $Y=0
+ $X2=4.56 $Y2=0
r100 51 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r101 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r102 48 71 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.905
+ $Y2=0
r103 48 50 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=3.57 $Y=0 $X2=2.16
+ $Y2=0
r104 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r105 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r106 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r107 44 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r108 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r109 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r110 41 68 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r111 41 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r112 39 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r113 39 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r114 39 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r115 37 46 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.68
+ $Y2=0
r116 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.875
+ $Y2=0
r117 36 50 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.16
+ $Y2=0
r118 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.875
+ $Y2=0
r119 32 79 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.472 $Y=0.085
+ $X2=7.472 $Y2=0
r120 32 34 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=7.472 $Y=0.085
+ $X2=7.472 $Y2=0.38
r121 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=0.085
+ $X2=6.14 $Y2=0
r122 28 30 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.14 $Y=0.085
+ $X2=6.14 $Y2=0.52
r123 24 71 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0
r124 24 26 13.2104 $w=6.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0.825
r125 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0
r126 20 22 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0.94
r127 16 68 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r128 16 18 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.56
r129 5 34 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=7.345
+ $Y=0.235 $X2=7.47 $Y2=0.38
r130 4 30 91 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=2 $X=5.94
+ $Y=0.595 $X2=6.14 $Y2=0.52
r131 3 26 91 $w=1.7e-07 $l=5.89979e-07 $layer=licon1_NDIFF $count=2 $X=3.49
+ $Y=0.815 $X2=4.075 $Y2=0.825
r132 2 22 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=1.615
+ $Y=0.815 $X2=1.875 $Y2=0.94
r133 1 18 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.35 $X2=0.26 $Y2=0.56
.ends

