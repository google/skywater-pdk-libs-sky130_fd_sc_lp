* File: sky130_fd_sc_lp__o22ai_2.pex.spice
* Created: Fri Aug 28 11:10:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22AI_2%B1 1 3 6 8 10 13 17 20 28
r41 24 34 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=0.295 $Y=1.44
+ $X2=0.295 $Y2=1.48
r42 23 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.34 $Y=1.44
+ $X2=0.555 $Y2=1.44
r43 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.44 $X2=0.34 $Y2=1.44
r44 20 24 5.96801 $w=2.78e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=1.295
+ $X2=0.295 $Y2=1.44
r45 18 28 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.77 $Y=1.44
+ $X2=0.985 $Y2=1.44
r46 18 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.77 $Y=1.44
+ $X2=0.555 $Y2=1.44
r47 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.44 $X2=0.77 $Y2=1.44
r48 15 34 1.39851 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=0.435 $Y=1.48
+ $X2=0.295 $Y2=1.48
r49 15 17 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.435 $Y=1.48
+ $X2=0.77 $Y2=1.48
r50 11 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.605
+ $X2=0.985 $Y2=1.44
r51 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.985 $Y=1.605
+ $X2=0.985 $Y2=2.465
r52 8 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.275
+ $X2=0.985 $Y2=1.44
r53 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.985 $Y=1.275
+ $X2=0.985 $Y2=0.745
r54 4 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.605
+ $X2=0.555 $Y2=1.44
r55 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.555 $Y=1.605
+ $X2=0.555 $Y2=2.465
r56 1 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.275
+ $X2=0.555 $Y2=1.44
r57 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.555 $Y=1.275
+ $X2=0.555 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%B2 3 5 7 10 12 14 15 16 24
r51 22 24 53.2078 $w=3.08e-07 $l=3.4e-07 $layer=POLY_cond $X=1.505 $Y=1.44
+ $X2=1.845 $Y2=1.44
r52 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.44 $X2=1.505 $Y2=1.44
r53 20 22 1.56494 $w=3.08e-07 $l=1e-08 $layer=POLY_cond $X=1.495 $Y=1.44
+ $X2=1.505 $Y2=1.44
r54 19 20 12.5195 $w=3.08e-07 $l=8e-08 $layer=POLY_cond $X=1.415 $Y=1.44
+ $X2=1.495 $Y2=1.44
r55 16 23 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=1.68 $Y=1.367
+ $X2=1.505 $Y2=1.367
r56 15 23 11.1586 $w=3.13e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=1.367
+ $X2=1.505 $Y2=1.367
r57 12 24 12.5195 $w=3.08e-07 $l=2.0106e-07 $layer=POLY_cond $X=1.925 $Y=1.275
+ $X2=1.845 $Y2=1.44
r58 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.925 $Y=1.275
+ $X2=1.925 $Y2=0.745
r59 8 24 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.605
+ $X2=1.845 $Y2=1.44
r60 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.845 $Y=1.605
+ $X2=1.845 $Y2=2.465
r61 5 20 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.275
+ $X2=1.495 $Y2=1.44
r62 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.495 $Y=1.275
+ $X2=1.495 $Y2=0.745
r63 1 19 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.605
+ $X2=1.415 $Y2=1.44
r64 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.415 $Y=1.605
+ $X2=1.415 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%A2 1 3 6 8 10 13 15 16 17 31
c54 31 0 1.85774e-19 $X=3.225 $Y=1.44
r55 30 31 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.155 $Y=1.44
+ $X2=3.225 $Y2=1.44
r56 28 30 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.135 $Y=1.44
+ $X2=3.155 $Y2=1.44
r57 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.135
+ $Y=1.44 $X2=3.135 $Y2=1.44
r58 26 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.795 $Y=1.44
+ $X2=3.135 $Y2=1.44
r59 25 26 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.725 $Y=1.44
+ $X2=2.795 $Y2=1.44
r60 22 25 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.705 $Y=1.44
+ $X2=2.725 $Y2=1.44
r61 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.44 $X2=2.705 $Y2=1.44
r62 17 29 17.0123 $w=3.13e-07 $l=4.65e-07 $layer=LI1_cond $X=3.6 $Y=1.367
+ $X2=3.135 $Y2=1.367
r63 16 29 0.548782 $w=3.13e-07 $l=1.5e-08 $layer=LI1_cond $X=3.12 $Y=1.367
+ $X2=3.135 $Y2=1.367
r64 16 23 15.183 $w=3.13e-07 $l=4.15e-07 $layer=LI1_cond $X=3.12 $Y=1.367
+ $X2=2.705 $Y2=1.367
r65 15 23 2.37806 $w=3.13e-07 $l=6.5e-08 $layer=LI1_cond $X=2.64 $Y=1.367
+ $X2=2.705 $Y2=1.367
r66 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=1.605
+ $X2=3.225 $Y2=1.44
r67 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.225 $Y=1.605
+ $X2=3.225 $Y2=2.465
r68 8 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=1.275
+ $X2=3.155 $Y2=1.44
r69 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.155 $Y=1.275
+ $X2=3.155 $Y2=0.745
r70 4 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.605
+ $X2=2.795 $Y2=1.44
r71 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.795 $Y=1.605
+ $X2=2.795 $Y2=2.465
r72 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.275
+ $X2=2.725 $Y2=1.44
r73 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.725 $Y=1.275
+ $X2=2.725 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%A1 1 3 6 8 10 13 15 16 22
c40 22 0 1.52337e-19 $X=4.085 $Y=1.44
c41 16 0 9.19853e-20 $X=4.56 $Y=1.295
c42 6 0 1.09502e-19 $X=3.655 $Y=2.465
r43 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.44 $X2=4.105 $Y2=1.44
r44 22 24 3.07987 $w=3.13e-07 $l=2e-08 $layer=POLY_cond $X=4.085 $Y=1.44
+ $X2=4.105 $Y2=1.44
r45 21 22 10.7796 $w=3.13e-07 $l=7e-08 $layer=POLY_cond $X=4.015 $Y=1.44
+ $X2=4.085 $Y2=1.44
r46 20 21 55.4377 $w=3.13e-07 $l=3.6e-07 $layer=POLY_cond $X=3.655 $Y=1.44
+ $X2=4.015 $Y2=1.44
r47 19 20 10.7796 $w=3.13e-07 $l=7e-08 $layer=POLY_cond $X=3.585 $Y=1.44
+ $X2=3.655 $Y2=1.44
r48 16 25 16.6464 $w=3.13e-07 $l=4.55e-07 $layer=LI1_cond $X=4.56 $Y=1.367
+ $X2=4.105 $Y2=1.367
r49 15 25 0.914637 $w=3.13e-07 $l=2.5e-08 $layer=LI1_cond $X=4.08 $Y=1.367
+ $X2=4.105 $Y2=1.367
r50 11 22 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.085 $Y=1.605
+ $X2=4.085 $Y2=1.44
r51 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.085 $Y=1.605
+ $X2=4.085 $Y2=2.465
r52 8 21 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.275
+ $X2=4.015 $Y2=1.44
r53 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.015 $Y=1.275
+ $X2=4.015 $Y2=0.745
r54 4 20 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.605
+ $X2=3.655 $Y2=1.44
r55 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.655 $Y=1.605
+ $X2=3.655 $Y2=2.465
r56 1 19 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.275
+ $X2=3.585 $Y2=1.44
r57 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.585 $Y=1.275
+ $X2=3.585 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%A_43_367# 1 2 3 12 16 17 19 22 24 26
r37 24 31 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=2.905
+ $X2=2.095 $Y2=2.99
r38 24 26 31.2489 $w=2.58e-07 $l=7.05e-07 $layer=LI1_cond $X=2.095 $Y=2.905
+ $X2=2.095 $Y2=2.2
r39 23 29 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.295 $Y=2.99 $X2=1.2
+ $Y2=2.99
r40 22 31 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.965 $Y=2.99
+ $X2=2.095 $Y2=2.99
r41 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.965 $Y=2.99
+ $X2=1.295 $Y2=2.99
r42 19 29 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.905 $X2=1.2
+ $Y2=2.99
r43 19 21 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=1.2 $Y=2.905
+ $X2=1.2 $Y2=1.98
r44 18 21 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=1.2 $Y=1.945 $X2=1.2
+ $Y2=1.98
r45 16 18 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.105 $Y=1.86
+ $X2=1.2 $Y2=1.945
r46 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=1.86
+ $X2=0.435 $Y2=1.86
r47 12 14 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.305 $Y=1.98
+ $X2=0.305 $Y2=2.91
r48 10 17 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.305 $Y=1.945
+ $X2=0.435 $Y2=1.86
r49 10 12 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.305 $Y=1.945
+ $X2=0.305 $Y2=1.98
r50 3 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.91
r51 3 26 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.2
r52 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=2.91
r53 2 21 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=1.98
r54 1 14 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.91
r55 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%VPWR 1 2 9 15 20 21 22 24 37 38 41
r59 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r62 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r63 32 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 31 34 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r65 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.77 $Y2=3.33
r67 29 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 27 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.77 $Y2=3.33
r71 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 22 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 22 32 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r74 20 34 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.6 $Y2=3.33
r75 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.87 $Y2=3.33
r76 19 37 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.87 $Y2=3.33
r78 15 18 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=3.87 $Y=2.12
+ $X2=3.87 $Y2=2.97
r79 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=3.33
r80 13 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=2.97
r81 9 12 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.77 $Y=2.2 $X2=0.77
+ $Y2=2.95
r82 7 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245 $X2=0.77
+ $Y2=3.33
r83 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=2.95
r84 2 18 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.835 $X2=3.87 $Y2=2.97
r85 2 15 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.835 $X2=3.87 $Y2=2.12
r86 1 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=2.95
r87 1 9 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%Y 1 2 3 4 13 19 21 22 23 27 30 34 35 36 41
+ 47
c67 23 0 1.09502e-19 $X=2.845 $Y=1.78
r68 42 47 1.35582 $w=2.53e-07 $l=3e-08 $layer=LI1_cond $X=2.127 $Y=1.695
+ $X2=2.127 $Y2=1.665
r69 36 42 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.127 $Y=1.78
+ $X2=2.127 $Y2=1.695
r70 36 47 1.26543 $w=2.53e-07 $l=2.8e-08 $layer=LI1_cond $X=2.127 $Y=1.637
+ $X2=2.127 $Y2=1.665
r71 35 36 15.4563 $w=2.53e-07 $l=3.42e-07 $layer=LI1_cond $X=2.127 $Y=1.295
+ $X2=2.127 $Y2=1.637
r72 35 41 11.9764 $w=2.53e-07 $l=2.65e-07 $layer=LI1_cond $X=2.127 $Y=1.295
+ $X2=2.127 $Y2=1.03
r73 34 41 3.12278 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=2.127 $Y=0.925
+ $X2=2.127 $Y2=1.03
r74 30 32 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.77 $Y=0.68
+ $X2=0.77 $Y2=0.925
r75 25 27 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.01 $Y=1.865
+ $X2=3.01 $Y2=1.98
r76 24 36 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.255 $Y=1.78
+ $X2=2.127 $Y2=1.78
r77 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.845 $Y=1.78
+ $X2=3.01 $Y2=1.865
r78 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.845 $Y=1.78
+ $X2=2.255 $Y2=1.78
r79 21 36 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2 $Y=1.78 $X2=2.127
+ $Y2=1.78
r80 21 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2 $Y=1.78 $X2=1.795
+ $Y2=1.78
r81 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.63 $Y=1.865
+ $X2=1.795 $Y2=1.78
r82 17 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.63 $Y=1.865
+ $X2=1.63 $Y2=1.98
r83 14 32 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.925
+ $X2=0.77 $Y2=0.925
r84 14 16 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=0.935 $Y=0.925
+ $X2=1.71 $Y2=0.925
r85 13 34 3.77708 $w=2.1e-07 $l=1.27e-07 $layer=LI1_cond $X=2 $Y=0.925 $X2=2.127
+ $Y2=0.925
r86 13 16 15.316 $w=2.08e-07 $l=2.9e-07 $layer=LI1_cond $X=2 $Y=0.925 $X2=1.71
+ $Y2=0.925
r87 4 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=1.98
r88 3 19 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.49
+ $Y=1.835 $X2=1.63 $Y2=1.98
r89 2 16 182 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.325 $X2=1.71 $Y2=0.925
r90 1 30 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.325 $X2=0.77 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%A_491_367# 1 2 3 10 12 14 17 20 21 24
c35 21 0 1.52337e-19 $X=3.535 $Y=1.78
r36 24 26 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=4.335 $Y=1.98
+ $X2=4.335 $Y2=2.91
r37 22 24 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.335 $Y=1.865
+ $X2=4.335 $Y2=1.98
r38 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.205 $Y=1.78
+ $X2=4.335 $Y2=1.865
r39 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.205 $Y=1.78
+ $X2=3.535 $Y2=1.78
r40 17 31 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=2.905
+ $X2=3.44 $Y2=2.99
r41 17 19 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=3.44 $Y=2.905
+ $X2=3.44 $Y2=1.98
r42 16 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.44 $Y=1.865
+ $X2=3.535 $Y2=1.78
r43 16 19 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=3.44 $Y=1.865
+ $X2=3.44 $Y2=1.98
r44 15 29 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.675 $Y=2.99
+ $X2=2.545 $Y2=2.99
r45 14 31 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=3.44 $Y2=2.99
r46 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=2.675 $Y2=2.99
r47 10 29 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=2.905
+ $X2=2.545 $Y2=2.99
r48 10 12 31.2489 $w=2.58e-07 $l=7.05e-07 $layer=LI1_cond $X=2.545 $Y=2.905
+ $X2=2.545 $Y2=2.2
r49 3 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.835 $X2=4.3 $Y2=2.91
r50 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.835 $X2=4.3 $Y2=1.98
r51 2 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.835 $X2=3.44 $Y2=2.91
r52 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.835 $X2=3.44 $Y2=1.98
r53 1 29 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.835 $X2=2.58 $Y2=2.91
r54 1 12 400 $w=1.7e-07 $l=4.22907e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.835 $X2=2.58 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%A_43_65# 1 2 3 4 5 18 21 22 23 26 27 28 32
+ 34 36 38 42 48
c65 48 0 9.37886e-20 $X=3.37 $Y=0.955
r66 41 42 7.16841 $w=3.93e-07 $l=1.15e-07 $layer=LI1_cond $X=1.22 $Y=0.452
+ $X2=1.105 $Y2=0.452
r67 36 50 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.265 $Y=0.87
+ $X2=4.265 $Y2=0.955
r68 36 38 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=4.265 $Y=0.87
+ $X2=4.265 $Y2=0.48
r69 35 48 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.465 $Y=0.955
+ $X2=3.375 $Y2=0.955
r70 34 50 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.135 $Y=0.955
+ $X2=4.265 $Y2=0.955
r71 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.135 $Y=0.955
+ $X2=3.465 $Y2=0.955
r72 30 48 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=0.87
+ $X2=3.375 $Y2=0.955
r73 30 32 24.0303 $w=1.78e-07 $l=3.9e-07 $layer=LI1_cond $X=3.375 $Y=0.87
+ $X2=3.375 $Y2=0.48
r74 29 46 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.605 $Y=0.955
+ $X2=2.515 $Y2=0.955
r75 28 48 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.285 $Y=0.955
+ $X2=3.375 $Y2=0.955
r76 28 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.285 $Y=0.955
+ $X2=2.605 $Y2=0.955
r77 27 46 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.87
+ $X2=2.515 $Y2=0.955
r78 26 44 5.59371 $w=1.8e-07 $l=1.98e-07 $layer=LI1_cond $X=2.515 $Y=0.65
+ $X2=2.515 $Y2=0.452
r79 26 27 13.5556 $w=1.78e-07 $l=2.2e-07 $layer=LI1_cond $X=2.515 $Y=0.65
+ $X2=2.515 $Y2=0.87
r80 23 41 2.39241 $w=3.93e-07 $l=8.2e-08 $layer=LI1_cond $X=1.302 $Y=0.452
+ $X2=1.22 $Y2=0.452
r81 23 25 24.4493 $w=3.93e-07 $l=8.38e-07 $layer=LI1_cond $X=1.302 $Y=0.452
+ $X2=2.14 $Y2=0.452
r82 22 44 2.54259 $w=3.95e-07 $l=9e-08 $layer=LI1_cond $X=2.425 $Y=0.452
+ $X2=2.515 $Y2=0.452
r83 22 25 8.31509 $w=3.93e-07 $l=2.85e-07 $layer=LI1_cond $X=2.425 $Y=0.452
+ $X2=2.14 $Y2=0.452
r84 21 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.435 $Y=0.34
+ $X2=1.105 $Y2=0.34
r85 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.305 $Y=0.425
+ $X2=0.435 $Y2=0.34
r86 16 18 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.305 $Y=0.425
+ $X2=0.305 $Y2=0.47
r87 5 50 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.325 $X2=4.23 $Y2=0.955
r88 5 38 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.325 $X2=4.23 $Y2=0.48
r89 4 48 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=3.23
+ $Y=0.325 $X2=3.37 $Y2=0.955
r90 4 32 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.23
+ $Y=0.325 $X2=3.37 $Y2=0.48
r91 3 46 182 $w=1.7e-07 $l=7.63544e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.325 $X2=2.51 $Y2=0.875
r92 3 44 182 $w=1.7e-07 $l=5.77971e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.325 $X2=2.51 $Y2=0.47
r93 3 25 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.325 $X2=2.14 $Y2=0.525
r94 2 41 182 $w=1.7e-07 $l=2.26274e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.325 $X2=1.22 $Y2=0.485
r95 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.325 $X2=0.34 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_2%VGND 1 2 9 13 16 17 19 20 21 34 35
r48 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r49 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r50 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r52 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r53 24 28 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r54 24 25 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 21 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r56 21 25 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=0.24
+ $Y2=0
r57 19 31 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.6
+ $Y2=0
r58 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.8
+ $Y2=0
r59 18 34 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=4.56
+ $Y2=0
r60 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=3.8
+ $Y2=0
r61 16 28 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.64
+ $Y2=0
r62 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.94
+ $Y2=0
r63 15 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.6
+ $Y2=0
r64 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.94
+ $Y2=0
r65 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=0.085 $X2=3.8
+ $Y2=0
r66 11 13 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=3.8 $Y=0.085 $X2=3.8
+ $Y2=0.575
r67 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085 $X2=2.94
+ $Y2=0
r68 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.94 $Y=0.085 $X2=2.94
+ $Y2=0.575
r69 2 13 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.66
+ $Y=0.325 $X2=3.8 $Y2=0.575
r70 1 9 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.325 $X2=2.94 $Y2=0.575
.ends

