* File: sky130_fd_sc_lp__clkinv_lp.pxi.spice
* Created: Fri Aug 28 10:18:25 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINV_LP%A N_A_M1000_g N_A_M1001_g N_A_c_29_n N_A_M1002_g
+ N_A_M1003_g N_A_c_32_n N_A_c_38_n N_A_c_33_n A A A N_A_c_35_n
+ PM_SKY130_FD_SC_LP__CLKINV_LP%A
x_PM_SKY130_FD_SC_LP__CLKINV_LP%VPWR N_VPWR_M1001_s N_VPWR_c_65_n N_VPWR_c_66_n
+ VPWR N_VPWR_c_67_n N_VPWR_c_64_n PM_SKY130_FD_SC_LP__CLKINV_LP%VPWR
x_PM_SKY130_FD_SC_LP__CLKINV_LP%Y N_Y_M1002_d N_Y_M1003_d Y Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__CLKINV_LP%Y
x_PM_SKY130_FD_SC_LP__CLKINV_LP%VGND N_VGND_M1000_s N_VGND_c_98_n N_VGND_c_99_n
+ VGND N_VGND_c_100_n N_VGND_c_101_n PM_SKY130_FD_SC_LP__CLKINV_LP%VGND
cc_1 VNB N_A_M1000_g 0.0350701f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.67
cc_2 VNB N_A_c_29_n 0.00722552f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.255
cc_3 VNB N_A_M1002_g 0.0299316f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_4 VNB N_A_M1003_g 0.0171175f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.66
cc_5 VNB N_A_c_32_n 0.0146721f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.255
cc_6 VNB N_A_c_33_n 0.00615289f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.255
cc_7 VNB A 0.029322f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_c_35_n 0.024341f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.345
cc_9 VNB N_VPWR_c_64_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_10 VNB Y 0.0235589f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.66
cc_11 VNB Y 0.038341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_98_n 0.0138117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_99_n 0.0370466f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.66
cc_14 VNB N_VGND_c_100_n 0.0300679f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_15 VNB N_VGND_c_101_n 0.128946f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.67
cc_16 VPB N_A_M1001_g 0.0439711f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.66
cc_17 VPB N_A_M1003_g 0.0508495f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.66
cc_18 VPB N_A_c_38_n 0.0175337f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.85
cc_19 VPB A 0.0381088f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_20 VPB N_A_c_35_n 0.00217867f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.345
cc_21 VPB N_VPWR_c_65_n 0.0134446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_66_n 0.0364925f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.66
cc_23 VPB N_VPWR_c_67_n 0.0292607f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.67
cc_24 VPB N_VPWR_c_64_n 0.0594858f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.67
cc_25 VPB Y 0.0093975f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.67
cc_26 VPB Y 0.022107f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.67
cc_27 VPB Y 0.0334624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 N_A_M1001_g N_VPWR_c_66_n 0.0171482f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_29 N_A_M1003_g N_VPWR_c_66_n 0.0025492f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_30 N_A_c_38_n N_VPWR_c_66_n 7.38037e-19 $X=0.455 $Y=1.85 $X2=0 $Y2=0
cc_31 A N_VPWR_c_66_n 0.0305155f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_32 N_A_M1001_g N_VPWR_c_67_n 0.00396895f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_33 N_A_M1003_g N_VPWR_c_67_n 0.00449508f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_34 N_A_M1001_g N_VPWR_c_64_n 0.0076915f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_35 N_A_M1003_g N_VPWR_c_64_n 0.00873509f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_36 N_A_M1000_g Y 0.00130204f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_37 N_A_M1002_g Y 0.0105259f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_38 N_A_M1001_g Y 0.00192394f $X=0.545 $Y=2.66 $X2=0 $Y2=0
cc_39 N_A_M1003_g Y 0.00436693f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_40 N_A_M1003_g Y 0.00913196f $X=0.935 $Y=2.66 $X2=0 $Y2=0
cc_41 N_A_M1002_g Y 0.0409418f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_42 A Y 0.0630741f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_43 N_A_M1000_g N_VGND_c_99_n 0.0141994f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_44 N_A_M1002_g N_VGND_c_99_n 0.0018473f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_45 N_A_c_32_n N_VGND_c_99_n 0.00132932f $X=0.455 $Y=1.255 $X2=0 $Y2=0
cc_46 A N_VGND_c_99_n 0.0205783f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A_M1000_g N_VGND_c_100_n 0.00426961f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_48 N_A_M1002_g N_VGND_c_100_n 0.00491683f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_VGND_c_101_n 0.00434697f $X=0.545 $Y=0.67 $X2=0 $Y2=0
cc_50 N_A_M1002_g N_VGND_c_101_n 0.00517496f $X=0.935 $Y=0.67 $X2=0 $Y2=0
cc_51 N_VPWR_c_66_n Y 0.021527f $X=0.33 $Y=2.485 $X2=0 $Y2=0
cc_52 N_VPWR_c_67_n Y 0.0158357f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_53 N_VPWR_c_64_n Y 0.0121432f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_54 Y N_VGND_c_99_n 0.0145731f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_55 Y N_VGND_c_100_n 0.0105762f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_56 Y N_VGND_c_101_n 0.011362f $X=1.115 $Y=0.47 $X2=0 $Y2=0
