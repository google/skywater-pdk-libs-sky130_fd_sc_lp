* File: sky130_fd_sc_lp__o21ba_2.spice
* Created: Wed Sep  2 10:16:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ba_2.pex.spice"
.subckt sky130_fd_sc_lp__o21ba_2  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_B1_N_M1008_g N_A_28_131#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_186_21#_M1001_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_X_M1001_d N_A_186_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_492_47#_M1007_d N_A_28_131#_M1007_g N_A_186_21#_M1007_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_492_47#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1003 N_A_492_47#_M1003_d N_A1_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1512 PD=2.25 PS=1.2 NRD=0 NRS=1.428 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_B1_N_M1010_g N_A_28_131#_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.107625 AS=0.1113 PD=0.8775 PS=1.37 NRD=94.3827 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1010_d N_A_186_21#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.322875 AS=0.1764 PD=2.6325 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_186_21#_M1011_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.27405 AS=0.1764 PD=1.695 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1000 N_A_186_21#_M1000_d N_A_28_131#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1827 AS=0.27405 PD=1.55 PS=1.695 NRD=0 NRS=13.2778 M=1 R=8.4
+ SA=75001.4 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1006 A_564_367# N_A2_M1006_g N_A_186_21#_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1827 PD=1.685 PS=1.55 NRD=24.6053 NRS=1.5563 M=1 R=8.4
+ SA=75001.9 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_564_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.26775 PD=3.05 PS=1.685 NRD=0 NRS=24.6053 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_40 VNB 0 2.74051e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o21ba_2.pxi.spice"
*
.ends
*
*
