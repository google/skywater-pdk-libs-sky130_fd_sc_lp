* File: sky130_fd_sc_lp__sleep_pargate_plv_28.pxi.spice
* Created: Fri Aug 28 11:32:16 2020
* 
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_28%SLEEP N_SLEEP_c_42_n N_SLEEP_M1000_g
+ N_SLEEP_c_43_n N_SLEEP_M1001_g N_SLEEP_c_44_n N_SLEEP_M1002_g N_SLEEP_c_45_n
+ N_SLEEP_M1003_g N_SLEEP_c_38_n N_SLEEP_c_47_n N_SLEEP_c_39_n N_SLEEP_c_49_n
+ N_SLEEP_c_50_n SLEEP SLEEP SLEEP SLEEP SLEEP N_SLEEP_c_41_n N_SLEEP_c_53_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_28%SLEEP
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_28%VIRTPWR N_VIRTPWR_M1000_d
+ N_VIRTPWR_M1001_d N_VIRTPWR_M1003_d N_VIRTPWR_c_120_n N_VIRTPWR_c_121_n
+ VIRTPWR N_VIRTPWR_c_122_n N_VIRTPWR_c_131_n N_VIRTPWR_c_135_n
+ N_VIRTPWR_c_139_n N_VIRTPWR_c_143_n N_VIRTPWR_c_123_n N_VIRTPWR_c_124_n
+ N_VIRTPWR_c_125_n N_VIRTPWR_c_115_n N_VIRTPWR_c_127_n N_VIRTPWR_c_116_n
+ N_VIRTPWR_c_117_n N_VIRTPWR_c_118_n VIRTPWR N_VIRTPWR_c_119_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_28%VIRTPWR
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_28%VPWR N_VPWR_M1000_s N_VPWR_M1002_s
+ VPWR N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_246_n
+ N_VPWR_c_248_n N_VPWR_c_250_n N_VPWR_c_252_n N_VPWR_c_229_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_28%VPWR
cc_1 noxref_1 N_SLEEP_c_38_n 0.00748887f $X=-0.19 $Y=-0.002 $X2=8.377 $Y2=1.82
cc_2 noxref_1 N_SLEEP_c_39_n 0.00985261f $X=-0.19 $Y=-0.002 $X2=8.377 $Y2=1.465
cc_3 noxref_1 SLEEP 0.0275283f $X=-0.19 $Y=-0.002 $X2=8.315 $Y2=0.84
cc_4 noxref_1 N_SLEEP_c_41_n 0.0520945f $X=-0.19 $Y=-0.002 $X2=8.42 $Y2=0.965
cc_5 noxref_1 VIRTPWR 0.105802f $X=-0.19 $Y=-0.002 $X2=8.377 $Y2=1.97
cc_6 noxref_1 N_VIRTPWR_c_115_n 0.0836651f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_7 noxref_1 N_VIRTPWR_c_116_n 0.0786895f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_8 noxref_1 N_VIRTPWR_c_117_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_9 noxref_1 N_VIRTPWR_c_118_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_10 noxref_1 N_VIRTPWR_c_119_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_11 noxref_1 N_VPWR_c_229_n 0.56571f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_12 VPB N_SLEEP_c_42_n 0.0222395f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=1.465
cc_13 VPB N_SLEEP_c_43_n 0.0164013f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=1.895
cc_14 VPB N_SLEEP_c_44_n 0.0164013f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.325
cc_15 VPB N_SLEEP_c_45_n 0.045835f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.755
cc_16 VPB N_SLEEP_c_38_n 0.0165207f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=1.82
cc_17 VPB N_SLEEP_c_47_n 0.0240095f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=2.25
cc_18 VPB N_SLEEP_c_39_n 0.00103476f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=1.465
cc_19 VPB N_SLEEP_c_49_n 0.0108874f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=1.895
cc_20 VPB N_SLEEP_c_50_n 0.0108874f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=2.325
cc_21 VPB SLEEP 0.0277668f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=0.84
cc_22 VPB N_SLEEP_c_41_n 0.0259328f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=0.965
cc_23 VPB N_SLEEP_c_53_n 0.0240095f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=2.665
cc_24 VPB N_VIRTPWR_c_120_n 0.0130323f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.755
cc_25 VPB N_VIRTPWR_c_121_n 0.0357155f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=1.82
cc_26 VPB N_VIRTPWR_c_122_n 0.15875f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=0.965
cc_27 VPB N_VIRTPWR_c_123_n 0.00413698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VIRTPWR_c_124_n 0.00214921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_VIRTPWR_c_125_n 0.0329627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VIRTPWR_c_115_n 0.0405705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VIRTPWR_c_127_n 0.0130323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VIRTPWR_c_116_n 0.0404102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_230_n 0.00214921f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=1.58
cc_34 VPB N_VPWR_c_231_n 0.00214921f $X=-0.19 $Y=1.655 $X2=8.52 $Y2=1.665
cc_35 VPB N_VPWR_c_232_n 0.00677224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_229_n 0.122603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 N_SLEEP_c_45_n N_VIRTPWR_c_120_n 0.0158929f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_38 N_SLEEP_c_45_n N_VIRTPWR_c_121_n 0.00259154f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_39 N_SLEEP_c_42_n N_VIRTPWR_c_131_n 0.00539584f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_40 N_SLEEP_c_43_n N_VIRTPWR_c_131_n 0.00101539f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_41 N_SLEEP_c_44_n N_VIRTPWR_c_131_n 0.00101539f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_42 N_SLEEP_c_45_n N_VIRTPWR_c_131_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_43 N_SLEEP_c_42_n N_VIRTPWR_c_135_n 0.00539584f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_44 N_SLEEP_c_43_n N_VIRTPWR_c_135_n 0.00101539f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_45 N_SLEEP_c_44_n N_VIRTPWR_c_135_n 0.00101539f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_46 N_SLEEP_c_45_n N_VIRTPWR_c_135_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_47 N_SLEEP_c_42_n N_VIRTPWR_c_139_n 0.00539584f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_48 N_SLEEP_c_43_n N_VIRTPWR_c_139_n 0.00101539f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_49 N_SLEEP_c_44_n N_VIRTPWR_c_139_n 0.00101539f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_50 N_SLEEP_c_45_n N_VIRTPWR_c_139_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_51 N_SLEEP_c_42_n N_VIRTPWR_c_143_n 0.00539734f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_52 N_SLEEP_c_43_n N_VIRTPWR_c_143_n 0.00101545f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_53 N_SLEEP_c_44_n N_VIRTPWR_c_143_n 0.00101545f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_54 N_SLEEP_c_45_n N_VIRTPWR_c_143_n 0.00539734f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_55 N_SLEEP_c_42_n N_VIRTPWR_c_123_n 0.0119829f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_56 SLEEP N_VIRTPWR_c_123_n 0.0112238f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_57 N_SLEEP_c_41_n N_VIRTPWR_c_123_n 0.00525497f $X=8.42 $Y=0.965 $X2=0 $Y2=0
cc_58 N_SLEEP_c_43_n N_VIRTPWR_c_124_n 0.0102402f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_59 N_SLEEP_c_44_n N_VIRTPWR_c_124_n 0.0102402f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_60 N_SLEEP_c_47_n N_VIRTPWR_c_124_n 0.00207026f $X=8.377 $Y=2.25 $X2=0 $Y2=0
cc_61 SLEEP N_VIRTPWR_c_124_n 0.0107074f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_62 N_SLEEP_c_45_n N_VIRTPWR_c_125_n 0.00576677f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_63 SLEEP N_VIRTPWR_c_125_n 0.0165417f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_64 N_SLEEP_c_45_n N_VIRTPWR_c_115_n 0.0037323f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_65 SLEEP N_VIRTPWR_c_115_n 0.0123629f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_66 N_SLEEP_c_45_n N_VIRTPWR_c_116_n 0.00224979f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_67 N_SLEEP_c_42_n N_VPWR_c_230_n 0.010275f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_68 N_SLEEP_c_43_n N_VPWR_c_230_n 0.0102402f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_69 N_SLEEP_c_38_n N_VPWR_c_230_n 0.00207026f $X=8.377 $Y=1.82 $X2=0 $Y2=0
cc_70 SLEEP N_VPWR_c_230_n 0.0107074f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_71 N_SLEEP_c_44_n N_VPWR_c_231_n 0.0102402f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_72 N_SLEEP_c_45_n N_VPWR_c_231_n 0.010275f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_73 SLEEP N_VPWR_c_231_n 0.0107074f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_74 N_SLEEP_c_53_n N_VPWR_c_231_n 0.00207026f $X=8.42 $Y=2.665 $X2=0 $Y2=0
cc_75 N_SLEEP_c_42_n N_VPWR_c_232_n 0.00908402f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_76 N_SLEEP_c_43_n N_VPWR_c_232_n 0.00343818f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_77 N_SLEEP_c_44_n N_VPWR_c_232_n 0.00343818f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_78 N_SLEEP_c_45_n N_VPWR_c_232_n 0.00303147f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_79 N_SLEEP_c_43_n N_VPWR_c_246_n 0.00101546f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_80 N_SLEEP_c_44_n N_VPWR_c_246_n 0.00101546f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_81 N_SLEEP_c_43_n N_VPWR_c_248_n 0.00101546f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_82 N_SLEEP_c_44_n N_VPWR_c_248_n 0.00101546f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_83 N_SLEEP_c_43_n N_VPWR_c_250_n 0.00101546f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_84 N_SLEEP_c_44_n N_VPWR_c_250_n 0.00101546f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_85 N_SLEEP_c_43_n N_VPWR_c_252_n 0.00320659f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_86 N_SLEEP_c_44_n N_VPWR_c_252_n 0.00320659f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_87 SLEEP N_VPWR_c_252_n 0.0203545f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_88 N_SLEEP_c_42_n N_VPWR_c_229_n 0.00722775f $X=8.17 $Y=1.465 $X2=0 $Y2=0
cc_89 N_SLEEP_c_43_n N_VPWR_c_229_n 0.00392683f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_90 N_SLEEP_c_44_n N_VPWR_c_229_n 0.00392683f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_91 N_SLEEP_c_45_n N_VPWR_c_229_n 0.00984441f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_92 N_SLEEP_c_38_n N_VPWR_c_229_n 0.00118998f $X=8.377 $Y=1.82 $X2=0 $Y2=0
cc_93 N_SLEEP_c_47_n N_VPWR_c_229_n 0.00118998f $X=8.377 $Y=2.25 $X2=0 $Y2=0
cc_94 SLEEP N_VPWR_c_229_n 0.0916633f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_95 N_SLEEP_c_41_n N_VPWR_c_229_n 0.0121961f $X=8.42 $Y=0.965 $X2=0 $Y2=0
cc_96 N_SLEEP_c_53_n N_VPWR_c_229_n 0.00118998f $X=8.42 $Y=2.665 $X2=0 $Y2=0
cc_97 N_VIRTPWR_c_131_n N_VPWR_M1000_s 2.87738e-19 $X=2.34 $Y=1.25 $X2=-0.19
+ $Y2=-0.002
cc_98 N_VIRTPWR_c_135_n N_VPWR_M1000_s 2.87738e-19 $X=3.895 $Y=1.25 $X2=-0.19
+ $Y2=-0.002
cc_99 N_VIRTPWR_c_139_n N_VPWR_M1000_s 2.87738e-19 $X=5.45 $Y=1.25 $X2=-0.19
+ $Y2=-0.002
cc_100 N_VIRTPWR_c_143_n N_VPWR_M1000_s 2.8786e-19 $X=7.005 $Y=1.25 $X2=-0.19
+ $Y2=-0.002
cc_101 N_VIRTPWR_c_131_n N_VPWR_M1002_s 2.87738e-19 $X=2.34 $Y=1.25 $X2=0 $Y2=0
cc_102 N_VIRTPWR_c_135_n N_VPWR_M1002_s 2.87738e-19 $X=3.895 $Y=1.25 $X2=0 $Y2=0
cc_103 N_VIRTPWR_c_139_n N_VPWR_M1002_s 2.87738e-19 $X=5.45 $Y=1.25 $X2=0 $Y2=0
cc_104 N_VIRTPWR_c_143_n N_VPWR_M1002_s 2.8786e-19 $X=7.005 $Y=1.25 $X2=0 $Y2=0
cc_105 N_VIRTPWR_c_131_n N_VPWR_c_230_n 0.0346616f $X=2.34 $Y=1.25 $X2=0 $Y2=0
cc_106 N_VIRTPWR_c_135_n N_VPWR_c_230_n 0.0346616f $X=3.895 $Y=1.25 $X2=0 $Y2=0
cc_107 N_VIRTPWR_c_139_n N_VPWR_c_230_n 0.0346616f $X=5.45 $Y=1.25 $X2=0 $Y2=0
cc_108 N_VIRTPWR_c_143_n N_VPWR_c_230_n 0.0356496f $X=7.005 $Y=1.25 $X2=0 $Y2=0
cc_109 N_VIRTPWR_c_123_n N_VPWR_c_230_n 0.258116f $X=7.785 $Y=1.25 $X2=0 $Y2=0
cc_110 N_VIRTPWR_c_124_n N_VPWR_c_230_n 0.251237f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_111 N_VIRTPWR_c_120_n N_VPWR_c_231_n 0.262559f $X=1.342 $Y=3.127 $X2=0 $Y2=0
cc_112 N_VIRTPWR_c_131_n N_VPWR_c_231_n 0.0346616f $X=2.34 $Y=1.25 $X2=0 $Y2=0
cc_113 N_VIRTPWR_c_135_n N_VPWR_c_231_n 0.0346616f $X=3.895 $Y=1.25 $X2=0 $Y2=0
cc_114 N_VIRTPWR_c_139_n N_VPWR_c_231_n 0.0346616f $X=5.45 $Y=1.25 $X2=0 $Y2=0
cc_115 N_VIRTPWR_c_143_n N_VPWR_c_231_n 0.0356496f $X=7.005 $Y=1.25 $X2=0 $Y2=0
cc_116 N_VIRTPWR_c_124_n N_VPWR_c_231_n 0.251237f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_117 N_VIRTPWR_c_115_n N_VPWR_c_231_n 0.00290716f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_118 N_VIRTPWR_c_116_n N_VPWR_c_231_n 0.00285709f $X=1.845 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VIRTPWR_c_117_n N_VPWR_c_231_n 0.0012824f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_120 N_VIRTPWR_c_118_n N_VPWR_c_231_n 0.0012824f $X=4.955 $Y=3.33 $X2=0 $Y2=0
cc_121 N_VIRTPWR_c_119_n N_VPWR_c_231_n 0.0012824f $X=6.51 $Y=3.33 $X2=0 $Y2=0
cc_122 N_VIRTPWR_M1001_d N_VPWR_c_232_n 3.18208e-19 $X=1.055 $Y=1.97 $X2=0 $Y2=0
cc_123 N_VIRTPWR_c_120_n N_VPWR_c_232_n 0.00580238f $X=1.342 $Y=3.127 $X2=0
+ $Y2=0
cc_124 N_VIRTPWR_c_131_n N_VPWR_c_232_n 0.0970367f $X=2.34 $Y=1.25 $X2=0 $Y2=0
cc_125 N_VIRTPWR_c_123_n N_VPWR_c_232_n 0.0160547f $X=7.785 $Y=1.25 $X2=0 $Y2=0
cc_126 N_VIRTPWR_c_124_n N_VPWR_c_232_n 0.0377876f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_127 N_VIRTPWR_c_116_n N_VPWR_c_232_n 0.026124f $X=1.845 $Y=3.33 $X2=0 $Y2=0
cc_128 N_VIRTPWR_c_122_n N_VPWR_c_246_n 0.00708574f $X=7.768 $Y=3.127 $X2=0
+ $Y2=0
cc_129 N_VIRTPWR_c_131_n N_VPWR_c_246_n 0.0970367f $X=2.34 $Y=1.25 $X2=0 $Y2=0
cc_130 N_VIRTPWR_c_135_n N_VPWR_c_246_n 0.0970367f $X=3.895 $Y=1.25 $X2=0 $Y2=0
cc_131 N_VIRTPWR_c_123_n N_VPWR_c_246_n 0.0160547f $X=7.785 $Y=1.25 $X2=0 $Y2=0
cc_132 N_VIRTPWR_c_124_n N_VPWR_c_246_n 0.0358966f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_133 N_VIRTPWR_c_117_n N_VPWR_c_246_n 0.0229031f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_134 N_VIRTPWR_c_122_n N_VPWR_c_248_n 0.00708574f $X=7.768 $Y=3.127 $X2=0
+ $Y2=0
cc_135 N_VIRTPWR_c_135_n N_VPWR_c_248_n 0.0970367f $X=3.895 $Y=1.25 $X2=0 $Y2=0
cc_136 N_VIRTPWR_c_139_n N_VPWR_c_248_n 0.0970367f $X=5.45 $Y=1.25 $X2=0 $Y2=0
cc_137 N_VIRTPWR_c_123_n N_VPWR_c_248_n 0.0160547f $X=7.785 $Y=1.25 $X2=0 $Y2=0
cc_138 N_VIRTPWR_c_124_n N_VPWR_c_248_n 0.0358966f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_139 N_VIRTPWR_c_118_n N_VPWR_c_248_n 0.0229031f $X=4.955 $Y=3.33 $X2=0 $Y2=0
cc_140 N_VIRTPWR_c_122_n N_VPWR_c_250_n 0.00708574f $X=7.768 $Y=3.127 $X2=0
+ $Y2=0
cc_141 N_VIRTPWR_c_139_n N_VPWR_c_250_n 0.0970367f $X=5.45 $Y=1.25 $X2=0 $Y2=0
cc_142 N_VIRTPWR_c_143_n N_VPWR_c_250_n 0.0970546f $X=7.005 $Y=1.25 $X2=0 $Y2=0
cc_143 N_VIRTPWR_c_123_n N_VPWR_c_250_n 0.0160547f $X=7.785 $Y=1.25 $X2=0 $Y2=0
cc_144 N_VIRTPWR_c_124_n N_VPWR_c_250_n 0.0358966f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_145 N_VIRTPWR_c_119_n N_VPWR_c_250_n 0.0229031f $X=6.51 $Y=3.33 $X2=0 $Y2=0
cc_146 N_VIRTPWR_M1001_d N_VPWR_c_252_n 2.87889e-19 $X=1.055 $Y=1.97 $X2=0 $Y2=0
cc_147 N_VIRTPWR_c_122_n N_VPWR_c_252_n 0.00580238f $X=7.768 $Y=3.127 $X2=0
+ $Y2=0
cc_148 N_VIRTPWR_c_143_n N_VPWR_c_252_n 0.0970546f $X=7.005 $Y=1.25 $X2=0 $Y2=0
cc_149 N_VIRTPWR_c_123_n N_VPWR_c_252_n 0.0160547f $X=7.785 $Y=1.25 $X2=0 $Y2=0
cc_150 N_VIRTPWR_c_124_n N_VPWR_c_252_n 0.0393669f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_151 N_VIRTPWR_c_115_n N_VPWR_c_252_n 0.026124f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_152 N_VIRTPWR_c_120_n N_VPWR_c_229_n 0.00611837f $X=1.342 $Y=3.127 $X2=0
+ $Y2=0
cc_153 VIRTPWR N_VPWR_c_229_n 0.224849f $X=0 $Y=3.085 $X2=0 $Y2=0
cc_154 N_VIRTPWR_c_122_n N_VPWR_c_229_n 0.0186573f $X=7.768 $Y=3.127 $X2=0 $Y2=0
cc_155 N_VIRTPWR_c_131_n N_VPWR_c_229_n 0.291337f $X=2.34 $Y=1.25 $X2=0 $Y2=0
cc_156 N_VIRTPWR_c_135_n N_VPWR_c_229_n 0.291337f $X=3.895 $Y=1.25 $X2=0 $Y2=0
cc_157 N_VIRTPWR_c_139_n N_VPWR_c_229_n 0.291337f $X=5.45 $Y=1.25 $X2=0 $Y2=0
cc_158 N_VIRTPWR_c_143_n N_VPWR_c_229_n 0.29811f $X=7.005 $Y=1.25 $X2=0 $Y2=0
cc_159 N_VIRTPWR_c_123_n N_VPWR_c_229_n 0.107316f $X=7.785 $Y=1.25 $X2=0 $Y2=0
cc_160 N_VIRTPWR_c_124_n N_VPWR_c_229_n 0.0173287f $X=7.785 $Y=2.11 $X2=0 $Y2=0
cc_161 N_VIRTPWR_c_115_n N_VPWR_c_229_n 0.227442f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VIRTPWR_c_127_n N_VPWR_c_229_n 0.00787277f $X=8.055 $Y=3.127 $X2=0
+ $Y2=0
cc_163 N_VIRTPWR_c_116_n N_VPWR_c_229_n 0.212348f $X=1.845 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VIRTPWR_c_117_n N_VPWR_c_229_n 0.0980574f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VIRTPWR_c_118_n N_VPWR_c_229_n 0.0980574f $X=4.955 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VIRTPWR_c_119_n N_VPWR_c_229_n 0.0980574f $X=6.51 $Y=3.33 $X2=0 $Y2=0
