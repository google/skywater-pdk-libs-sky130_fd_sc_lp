* File: sky130_fd_sc_lp__dlclkp_1.pex.spice
* Created: Wed Sep  2 09:45:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%A_80_269# 1 2 9 13 18 19 21 24 25 27 30 31
+ 36 37
c92 27 0 1.98194e-19 $X=1.895 $Y=0.7
r93 35 37 16.6364 $w=1.78e-07 $l=2.7e-07 $layer=LI1_cond $X=1.4 $Y=1.65 $X2=1.67
+ $Y2=1.65
r94 35 36 5.28416 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=1.65
+ $X2=1.315 $Y2=1.65
r95 31 41 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.51
+ $X2=0.597 $Y2=1.675
r96 31 40 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.51
+ $X2=0.597 $Y2=1.345
r97 30 33 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.665 $Y=1.51
+ $X2=0.665 $Y2=1.645
r98 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.51 $X2=0.63 $Y2=1.51
r99 25 27 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=1.755 $Y=0.695
+ $X2=1.895 $Y2=0.695
r100 24 37 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.67 $Y=1.56 $X2=1.67
+ $Y2=1.65
r101 23 25 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.67 $Y=0.795
+ $X2=1.755 $Y2=0.695
r102 23 24 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.67 $Y=0.795
+ $X2=1.67 $Y2=1.56
r103 19 21 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.485 $Y=2.61
+ $X2=1.905 $Y2=2.61
r104 18 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.4 $Y=2.485
+ $X2=1.485 $Y2=2.61
r105 17 35 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.4 $Y=1.74 $X2=1.4
+ $Y2=1.65
r106 17 18 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.4 $Y=1.74
+ $X2=1.4 $Y2=2.485
r107 16 33 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.795 $Y=1.645
+ $X2=0.665 $Y2=1.645
r108 16 36 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.795 $Y=1.645
+ $X2=1.315 $Y2=1.645
r109 13 40 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.63 $Y=0.655
+ $X2=0.63 $Y2=1.345
r110 9 41 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.675
r111 2 21 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=2.4 $X2=1.905 $Y2=2.61
r112 1 27 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.755
+ $Y=0.405 $X2=1.895 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%GATE 3 7 9 12
r48 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.295
+ $X2=1.23 $Y2=1.46
r49 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.295
+ $X2=1.23 $Y2=1.13
r50 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.295 $X2=1.23 $Y2=1.295
r51 7 14 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.32 $Y=0.615
+ $X2=1.32 $Y2=1.13
r52 3 15 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=1.29 $Y=2.72
+ $X2=1.29 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%A_315_382# 1 2 9 13 16 17 19 21 24 27 30 34
+ 35 38 42
c129 35 0 1.59082e-19 $X=2.13 $Y=1.13
c130 30 0 1.11739e-19 $X=2.095 $Y=2.075
r131 45 46 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=3.695 $Y=2.12
+ $X2=3.695 $Y2=2.31
r132 42 45 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=3.695 $Y=2.02
+ $X2=3.695 $Y2=2.12
r133 38 40 6.35831 $w=2.88e-07 $l=1.6e-07 $layer=LI1_cond $X=3.355 $Y=0.61
+ $X2=3.355 $Y2=0.77
r134 35 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.13
+ $X2=2.13 $Y2=0.965
r135 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.13 $X2=2.13 $Y2=1.13
r136 31 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.01 $Y=1.13
+ $X2=2.13 $Y2=1.13
r137 29 30 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=2.075
+ $X2=2.095 $Y2=2.075
r138 27 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=2.075
+ $X2=1.74 $Y2=2.24
r139 26 29 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.74 $Y=2.075
+ $X2=2.01 $Y2=2.075
r140 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=2.075 $X2=1.74 $Y2=2.075
r141 23 24 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=4.67 $Y=0.855
+ $X2=4.67 $Y2=2.225
r142 22 46 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.825 $Y=2.31
+ $X2=3.695 $Y2=2.31
r143 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.585 $Y=2.31
+ $X2=4.67 $Y2=2.225
r144 21 22 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.585 $Y=2.31
+ $X2=3.825 $Y2=2.31
r145 20 40 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.5 $Y=0.77
+ $X2=3.355 $Y2=0.77
r146 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.585 $Y=0.77
+ $X2=4.67 $Y2=0.855
r147 19 20 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=4.585 $Y=0.77
+ $X2=3.5 $Y2=0.77
r148 17 42 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.565 $Y=2.02
+ $X2=3.695 $Y2=2.02
r149 17 30 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=3.565 $Y=2.02
+ $X2=2.095 $Y2=2.02
r150 16 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=1.91
+ $X2=2.01 $Y2=2.075
r151 15 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=1.295
+ $X2=2.01 $Y2=1.13
r152 15 16 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.01 $Y=1.295
+ $X2=2.01 $Y2=1.91
r153 13 52 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.11 $Y=0.615
+ $X2=2.11 $Y2=0.965
r154 9 50 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.65 $Y=2.72
+ $X2=1.65 $Y2=2.24
r155 2 45 600 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.975 $X2=3.65 $Y2=2.12
r156 1 38 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.405 $X2=3.335 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%A_27_367# 1 2 9 13 14 15 18 22 26 29 32 34
+ 36 39 40 41 43 44 45 47 48 49 51 52 54 57 58 60 61 63 65 69 70 72 76 81 84
c231 84 0 1.98194e-19 $X=2.67 $Y=0.935
c232 76 0 9.55795e-20 $X=3.75 $Y=2.65
c233 70 0 1.71081e-20 $X=2.67 $Y=1.1
c234 69 0 4.87977e-20 $X=2.67 $Y=1.1
c235 63 0 1.46981e-19 $X=0.337 $Y=0.957
c236 18 0 1.18845e-19 $X=5.295 $Y=0.605
r237 81 88 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.75 $Y=2.94
+ $X2=3.75 $Y2=3.115
r238 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.75
+ $Y=2.94 $X2=3.75 $Y2=2.94
r239 78 80 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.75 $Y=2.655
+ $X2=3.75 $Y2=2.94
r240 76 78 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.75 $Y=2.65
+ $X2=3.75 $Y2=2.655
r241 72 74 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.31 $Y=2.36
+ $X2=3.31 $Y2=2.655
r242 70 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.1
+ $X2=2.67 $Y2=0.935
r243 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.1 $X2=2.67 $Y2=1.1
r244 61 92 12.9107 $w=2.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.51 $Y=1.17
+ $X2=5.585 $Y2=1.17
r245 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.51
+ $Y=1.17 $X2=5.51 $Y2=1.17
r246 58 60 14.9457 $w=3.18e-07 $l=4.15e-07 $layer=LI1_cond $X=5.095 $Y=1.165
+ $X2=5.51 $Y2=1.165
r247 56 58 7.68211 $w=3.2e-07 $l=1.9799e-07 $layer=LI1_cond $X=5.01 $Y=1.325
+ $X2=5.095 $Y2=1.165
r248 56 57 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=5.01 $Y=1.325
+ $X2=5.01 $Y2=2.565
r249 55 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=2.65
+ $X2=3.75 $Y2=2.65
r250 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.925 $Y=2.65
+ $X2=5.01 $Y2=2.565
r251 54 55 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.925 $Y=2.65
+ $X2=3.915 $Y2=2.65
r252 53 74 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=2.655
+ $X2=3.31 $Y2=2.655
r253 52 78 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=2.655
+ $X2=3.75 $Y2=2.655
r254 52 53 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=3.585 $Y=2.655
+ $X2=3.395 $Y2=2.655
r255 51 69 4.93904 $w=3.13e-07 $l=1.35e-07 $layer=LI1_cond $X=2.535 $Y=1.107
+ $X2=2.67 $Y2=1.107
r256 50 51 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.535 $Y=0.425
+ $X2=2.535 $Y2=0.95
r257 48 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=2.36
+ $X2=3.31 $Y2=2.36
r258 48 49 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.225 $Y=2.36
+ $X2=2.445 $Y2=2.36
r259 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=2.445
+ $X2=2.445 $Y2=2.36
r260 46 47 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.36 $Y=2.445
+ $X2=2.36 $Y2=2.905
r261 44 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.45 $Y=0.34
+ $X2=2.535 $Y2=0.425
r262 44 45 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.45 $Y=0.34
+ $X2=1.415 $Y2=0.34
r263 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.33 $Y=0.425
+ $X2=1.415 $Y2=0.34
r264 42 43 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.33 $Y=0.425
+ $X2=1.33 $Y2=0.82
r265 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.275 $Y=2.99
+ $X2=2.36 $Y2=2.905
r266 40 41 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.275 $Y=2.99
+ $X2=1.145 $Y2=2.99
r267 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.905
+ $X2=1.145 $Y2=2.99
r268 38 39 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.06 $Y=2.07
+ $X2=1.06 $Y2=2.905
r269 37 63 4.29663 $w=1.7e-07 $l=2.67741e-07 $layer=LI1_cond $X=0.58 $Y=0.905
+ $X2=0.337 $Y2=0.957
r270 36 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.245 $Y=0.905
+ $X2=1.33 $Y2=0.82
r271 36 37 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.245 $Y=0.905
+ $X2=0.58 $Y2=0.905
r272 35 65 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.985
+ $X2=0.26 $Y2=1.985
r273 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=1.985
+ $X2=1.06 $Y2=2.07
r274 34 35 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.975 $Y=1.985
+ $X2=0.425 $Y2=1.985
r275 30 65 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.07 $X2=0.26
+ $Y2=1.985
r276 30 32 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=0.26 $Y=2.07
+ $X2=0.26 $Y2=2.91
r277 29 65 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.23 $Y=1.9
+ $X2=0.26 $Y2=1.985
r278 28 63 2.56749 $w=3.75e-07 $l=1.83875e-07 $layer=LI1_cond $X=0.23 $Y=1.095
+ $X2=0.337 $Y2=0.957
r279 28 29 34.3599 $w=2.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.23 $Y=1.095
+ $X2=0.23 $Y2=1.9
r280 24 63 2.56749 $w=3.75e-07 $l=1.37996e-07 $layer=LI1_cond $X=0.335 $Y=0.82
+ $X2=0.337 $Y2=0.957
r281 24 26 9.96732 $w=4.78e-07 $l=4e-07 $layer=LI1_cond $X=0.335 $Y=0.82
+ $X2=0.335 $Y2=0.42
r282 20 92 17.3521 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=1.335
+ $X2=5.585 $Y2=1.17
r283 20 22 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.585 $Y=1.335
+ $X2=5.585 $Y2=2.155
r284 16 61 37.0107 $w=2.8e-07 $l=2.85832e-07 $layer=POLY_cond $X=5.295 $Y=1.005
+ $X2=5.51 $Y2=1.17
r285 16 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.295 $Y=1.005
+ $X2=5.295 $Y2=0.605
r286 14 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=3.115
+ $X2=3.75 $Y2=3.115
r287 14 15 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=3.585 $Y=3.115
+ $X2=2.625 $Y2=3.115
r288 13 84 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.58 $Y=0.615
+ $X2=2.58 $Y2=0.935
r289 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=3.04
+ $X2=2.625 $Y2=3.115
r290 7 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.55 $Y=3.04 $X2=2.55
+ $Y2=2.61
r291 2 65 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r292 2 32 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r293 1 26 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.29
+ $Y=0.235 $X2=0.415 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%A_321_55# 1 2 9 11 12 15 19 21 23 25 28 29
+ 30 31 36 37 38 40 42 46
c107 37 0 8.84298e-20 $X=3.17 $Y=1.505
c108 31 0 1.59082e-19 $X=3.045 $Y=1.635
c109 28 0 4.87977e-20 $X=3.21 $Y=1.505
c110 21 0 2.06425e-19 $X=3.27 $Y=1.865
c111 12 0 1.11739e-19 $X=1.755 $Y=1.595
r112 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.21
+ $Y=1.2 $X2=3.21 $Y2=1.2
r113 40 48 2.9017 $w=3.3e-07 $l=1.13e-07 $layer=LI1_cond $X=4.25 $Y=1.25
+ $X2=4.25 $Y2=1.137
r114 40 42 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.25 $Y=1.25
+ $X2=4.25 $Y2=1.96
r115 39 45 3.593 $w=2.25e-07 $l=1.25e-07 $layer=LI1_cond $X=3.295 $Y=1.137
+ $X2=3.17 $Y2=1.137
r116 38 48 4.237 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=1.137
+ $X2=4.25 $Y2=1.137
r117 38 39 40.4636 $w=2.23e-07 $l=7.9e-07 $layer=LI1_cond $X=4.085 $Y=1.137
+ $X2=3.295 $Y2=1.137
r118 36 45 3.24808 $w=2.5e-07 $l=1.13e-07 $layer=LI1_cond $X=3.17 $Y=1.25
+ $X2=3.17 $Y2=1.137
r119 36 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.17 $Y=1.25
+ $X2=3.17 $Y2=1.505
r120 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=1.68 $X2=2.43 $Y2=1.68
r121 31 37 6.8199 $w=2.6e-07 $l=1.82071e-07 $layer=LI1_cond $X=3.045 $Y=1.635
+ $X2=3.17 $Y2=1.505
r122 31 33 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=3.045 $Y=1.635
+ $X2=2.43 $Y2=1.635
r123 29 34 98.578 $w=3.6e-07 $l=6.15e-07 $layer=POLY_cond $X=3.045 $Y=1.685
+ $X2=2.43 $Y2=1.685
r124 29 30 0.267992 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=3.045 $Y=1.685
+ $X2=3.045 $Y2=1.505
r125 28 46 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=3.21 $Y=1.505
+ $X2=3.21 $Y2=1.2
r126 28 30 28.1878 $w=2.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.505
+ $X2=3.045 $Y2=1.505
r127 27 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.035
+ $X2=3.21 $Y2=1.2
r128 24 34 26.4478 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.685
+ $X2=2.43 $Y2=1.685
r129 24 25 12.2198 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.265 $Y=1.685
+ $X2=2.19 $Y2=1.685
r130 21 30 28.1878 $w=2.4e-07 $l=4.58912e-07 $layer=POLY_cond $X=3.27 $Y=1.865
+ $X2=3.045 $Y2=1.505
r131 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.27 $Y=1.865
+ $X2=3.27 $Y2=2.295
r132 19 27 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.12 $Y=0.615
+ $X2=3.12 $Y2=1.035
r133 13 25 13.9189 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.19 $Y=1.865
+ $X2=2.19 $Y2=1.685
r134 13 15 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.19 $Y=1.865
+ $X2=2.19 $Y2=2.61
r135 11 25 12.2198 $w=2.7e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.115 $Y=1.595
+ $X2=2.19 $Y2=1.685
r136 11 12 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=2.115 $Y=1.595
+ $X2=1.755 $Y2=1.595
r137 7 12 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.68 $Y=1.505
+ $X2=1.755 $Y2=1.595
r138 7 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.68 $Y=1.505
+ $X2=1.68 $Y2=0.615
r139 2 42 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.835 $X2=4.25 $Y2=1.96
r140 1 48 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.825 $X2=4.095 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%CLK 1 5 7 9 10 11 14 16 18 22 24 28 30
c75 30 0 7.13217e-20 $X=3.945 $Y=1.585
c76 7 0 8.01478e-20 $X=4.565 $Y=1.725
r77 27 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.585
+ $X2=3.945 $Y2=1.585
r78 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.585 $X2=3.78 $Y2=1.585
r79 24 28 6.01275 $w=3.43e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=1.592
+ $X2=3.78 $Y2=1.592
r80 21 22 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.935 $Y=1.65
+ $X2=5.155 $Y2=1.65
r81 19 20 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=4.31 $Y=1.65
+ $X2=4.565 $Y2=1.65
r82 16 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.155 $Y=1.725
+ $X2=5.155 $Y2=1.65
r83 16 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.155 $Y=1.725
+ $X2=5.155 $Y2=2.155
r84 12 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.935 $Y=1.575
+ $X2=4.935 $Y2=1.65
r85 12 14 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=4.935 $Y=1.575
+ $X2=4.935 $Y2=0.605
r86 11 20 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.64 $Y=1.65
+ $X2=4.565 $Y2=1.65
r87 10 21 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.86 $Y=1.65
+ $X2=4.935 $Y2=1.65
r88 10 11 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.86 $Y=1.65
+ $X2=4.64 $Y2=1.65
r89 7 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.565 $Y=1.725
+ $X2=4.565 $Y2=1.65
r90 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.565 $Y=1.725
+ $X2=4.565 $Y2=2.155
r91 3 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.31 $Y=1.575
+ $X2=4.31 $Y2=1.65
r92 3 5 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.31 $Y=1.575 $X2=4.31
+ $Y2=1.035
r93 1 19 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.235 $Y=1.65
+ $X2=4.31 $Y2=1.65
r94 1 30 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.235 $Y=1.65
+ $X2=3.945 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%A_1046_367# 1 2 9 13 17 19 20 21 24 26 32
c58 21 0 1.18845e-19 $X=5.945 $Y=0.75
c59 20 0 7.97162e-20 $X=5.465 $Y=1.58
r60 32 35 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.132 $Y=1.5
+ $X2=6.132 $Y2=1.665
r61 32 34 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.132 $Y=1.5
+ $X2=6.132 $Y2=1.335
r62 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.5 $X2=6.11 $Y2=1.5
r63 26 28 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.51 $Y=0.605
+ $X2=5.51 $Y2=0.75
r64 24 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=1.495
+ $X2=6.07 $Y2=1.58
r65 23 24 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=6.07 $Y=0.835
+ $X2=6.07 $Y2=1.495
r66 22 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=0.75
+ $X2=5.51 $Y2=0.75
r67 21 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.945 $Y=0.75
+ $X2=6.07 $Y2=0.835
r68 21 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.945 $Y=0.75
+ $X2=5.675 $Y2=0.75
r69 19 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=1.58
+ $X2=6.07 $Y2=1.58
r70 19 20 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.945 $Y=1.58
+ $X2=5.465 $Y2=1.58
r71 15 20 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.365 $Y=1.665
+ $X2=5.465 $Y2=1.58
r72 15 17 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.365 $Y=1.665
+ $X2=5.365 $Y2=1.96
r73 13 35 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=6.245 $Y=2.465
+ $X2=6.245 $Y2=1.665
r74 9 34 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.245 $Y=0.655
+ $X2=6.245 $Y2=1.335
r75 2 17 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.23
+ $Y=1.835 $X2=5.37 $Y2=1.96
r76 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.395 $X2=5.51 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%VPWR 1 2 3 4 15 19 23 27 32 33 35 36 37 39
+ 57 63 64 67 70
c88 64 0 1.90993e-19 $X=6.48 $Y=3.33
r89 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 64 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r92 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r93 61 70 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=5.915 $Y2=3.33
r94 61 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6.48 $Y2=3.33
r95 60 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r96 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 57 70 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=5.635 $Y=3.33
+ $X2=5.915 $Y2=3.33
r98 57 59 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.635 $Y=3.33
+ $X2=5.52 $Y2=3.33
r99 56 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r100 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r101 52 55 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r102 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 50 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r104 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 47 50 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 46 49 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 44 67 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.705 $Y2=3.33
r110 44 46 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 39 67 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.705 $Y2=3.33
r114 39 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r115 37 56 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 37 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 35 55 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.86 $Y2=3.33
r119 34 59 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.025 $Y=3.33
+ $X2=5.52 $Y2=3.33
r120 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=3.33
+ $X2=4.86 $Y2=3.33
r121 32 49 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.715 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=3.33
+ $X2=2.88 $Y2=3.33
r123 31 52 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.045 $Y=3.33
+ $X2=3.12 $Y2=3.33
r124 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=3.33
+ $X2=2.88 $Y2=3.33
r125 27 30 14.3102 $w=5.58e-07 $l=6.7e-07 $layer=LI1_cond $X=5.915 $Y=1.96
+ $X2=5.915 $Y2=2.63
r126 25 70 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=3.245
+ $X2=5.915 $Y2=3.33
r127 25 30 13.1355 $w=5.58e-07 $l=6.15e-07 $layer=LI1_cond $X=5.915 $Y=3.245
+ $X2=5.915 $Y2=2.63
r128 21 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.86 $Y=3.245
+ $X2=4.86 $Y2=3.33
r129 21 23 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.86 $Y=3.245
+ $X2=4.86 $Y2=3.01
r130 17 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=3.33
r131 17 19 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=2.745
r132 13 67 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=3.245
+ $X2=0.705 $Y2=3.33
r133 13 15 46.5818 $w=1.98e-07 $l=8.4e-07 $layer=LI1_cond $X=0.705 $Y=3.245
+ $X2=0.705 $Y2=2.405
r134 4 30 300 $w=1.7e-07 $l=9.6238e-07 $layer=licon1_PDIFF $count=2 $X=5.66
+ $Y=1.835 $X2=6.03 $Y2=2.63
r135 4 27 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.66
+ $Y=1.835 $X2=5.8 $Y2=1.96
r136 3 23 600 $w=1.7e-07 $l=1.28028e-06 $layer=licon1_PDIFF $count=1 $X=4.64
+ $Y=1.835 $X2=4.86 $Y2=3.01
r137 2 19 600 $w=1.7e-07 $l=4.54973e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=2.4 $X2=2.88 $Y2=2.745
r138 1 15 300 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%GCLK 1 2 7 8 9 10 11 18
r10 11 32 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=6.495 $Y=2.775
+ $X2=6.495 $Y2=2.91
r11 10 11 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=6.495 $Y=2.405
+ $X2=6.495 $Y2=2.775
r12 9 10 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=6.495 $Y=1.98
+ $X2=6.495 $Y2=2.405
r13 8 9 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=6.495 $Y=1.665
+ $X2=6.495 $Y2=1.98
r14 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=6.495 $Y=1.295
+ $X2=6.495 $Y2=1.665
r15 7 18 38.7841 $w=2.58e-07 $l=8.75e-07 $layer=LI1_cond $X=6.495 $Y=1.295
+ $X2=6.495 $Y2=0.42
r16 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.91
r17 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=1.98
r18 1 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.235 $X2=6.46 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_1%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 47
+ 54 61 62 65 68
c72 62 0 1.46981e-19 $X=6.48 $Y=0
r73 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r74 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r75 62 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r76 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r77 59 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.03
+ $Y2=0
r78 59 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.48
+ $Y2=0
r79 58 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r80 58 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r81 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r82 55 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.77 $Y=0 $X2=4.605
+ $Y2=0
r83 55 57 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.77 $Y=0 $X2=5.52
+ $Y2=0
r84 54 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=6.03
+ $Y2=0
r85 54 57 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=5.52
+ $Y2=0
r86 53 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r87 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r88 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r89 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r90 47 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.605
+ $Y2=0
r91 47 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.08
+ $Y2=0
r92 46 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r93 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r94 43 46 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r95 42 45 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r96 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r97 39 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r98 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r99 35 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r100 35 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r101 33 45 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r102 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.915
+ $Y2=0
r103 32 49 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.12
+ $Y2=0
r104 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.915
+ $Y2=0
r105 30 38 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.72
+ $Y2=0
r106 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.91
+ $Y2=0
r107 29 42 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.2
+ $Y2=0
r108 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.91
+ $Y2=0
r109 25 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0
r110 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0.38
r111 21 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.605 $Y=0.085
+ $X2=4.605 $Y2=0
r112 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.605 $Y=0.085
+ $X2=4.605 $Y2=0.42
r113 17 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r114 17 19 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.615
r115 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=0.085
+ $X2=0.91 $Y2=0
r116 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.91 $Y=0.085
+ $X2=0.91 $Y2=0.535
r117 4 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.235 $X2=6.03 $Y2=0.38
r118 3 23 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.825 $X2=4.605 $Y2=0.42
r119 2 19 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2.655
+ $Y=0.405 $X2=2.88 $Y2=0.615
r120 1 15 182 $w=1.7e-07 $l=3.8923e-07 $layer=licon1_NDIFF $count=1 $X=0.705
+ $Y=0.235 $X2=0.91 $Y2=0.535
.ends

