* File: sky130_fd_sc_lp__buflp_1.spice
* Created: Wed Sep  2 09:36:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buflp_1.pex.spice"
.subckt sky130_fd_sc_lp__buflp_1  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1003 A_116_47# N_A_86_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2394 PD=1.08 PS=2.25 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A_86_21#_M1000_g A_116_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1974 AS=0.1008 PD=1.68 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1006 A_308_131# N_A_M1006_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0987 PD=0.66 PS=0.84 NRD=18.564 NRS=51.42 M=1 R=2.8 SA=75001.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_86_21#_M1004_d N_A_M1004_g A_308_131# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_116_367# N_A_86_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3591 PD=1.5 PS=3.09 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_86_21#_M1005_g A_116_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.295437 AS=0.1512 PD=2.22821 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1007 A_308_403# N_A_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.150063 PD=0.88 PS=1.13179 NRD=19.9955 NRS=43.8522 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_86_21#_M1001_d N_A_M1001_g A_308_403# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__buflp_1.pxi.spice"
*
.ends
*
*
