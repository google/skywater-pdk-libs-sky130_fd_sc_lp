* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 COUT a_80_27# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_417_457# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_1212_411# B a_1290_411# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR A a_231_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR A a_854_411# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_818_83# a_80_27# a_1118_411# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_854_411# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_431_137# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1290_411# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_231_457# B a_80_27# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VGND A a_267_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1118_411# CIN a_1212_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND B a_431_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 COUT a_80_27# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_1118_411# CIN a_1212_411# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VPWR B a_854_411# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_854_411# a_80_27# a_1118_411# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_267_137# B a_80_27# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1212_125# B a_1290_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_818_83# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR B a_417_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_1290_125# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_80_27# CIN a_417_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VPWR a_1118_411# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VGND A a_818_83# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_1118_411# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_80_27# CIN a_431_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VGND B a_818_83# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
