* File: sky130_fd_sc_lp__a22oi_m.spice
* Created: Wed Sep  2 09:23:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a22oi_m  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1007 A_133_47# N_B2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1239 PD=0.63 PS=1.43 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g A_133_47# VNB NSHORT L=0.15 W=0.42 AD=0.08295
+ AS=0.0441 PD=0.815 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1002 A_314_47# N_A1_M1002_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.08295 PD=0.63 PS=0.815 NRD=14.28 NRS=32.856 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g A_314_47# VNB NSHORT L=0.15 W=0.42 AD=0.1281
+ AS=0.0441 PD=1.45 PS=0.63 NRD=11.424 NRS=14.28 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g N_A_39_496#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=37.5088 M=1 R=2.8 SA=75000.3
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_A_39_496#_M1006_d N_B1_M1006_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_39_496#_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_39_496#_M1000_d N_A2_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__a22oi_m.pxi.spice"
*
.ends
*
*
