* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and3_4 A B C VGND VNB VPB VPWR X
X0 X a_77_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_77_47# A a_160_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR a_77_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_77_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_77_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_77_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR a_77_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 X a_77_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_160_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND a_77_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_77_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR B a_77_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 X a_77_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
