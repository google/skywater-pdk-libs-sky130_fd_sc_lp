* File: sky130_fd_sc_lp__a31o_0.pex.spice
* Created: Wed Sep  2 09:26:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31O_0%A_86_241# 1 2 9 13 18 19 23 24 25 26 27 28 29
+ 31 35 37 43
r97 35 43 7.04571 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.775 $Y=2.545
+ $X2=2.775 $Y2=2.395
r98 35 37 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.775 $Y=2.545
+ $X2=2.775 $Y2=2.56
r99 33 43 28.8364 $w=1.98e-07 $l=5.2e-07 $layer=LI1_cond $X=2.725 $Y=1.875
+ $X2=2.725 $Y2=2.395
r100 29 41 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.32 $Y=0.46
+ $X2=1.32 $Y2=0.755
r101 29 31 36.1448 $w=3.28e-07 $l=1.035e-06 $layer=LI1_cond $X=1.405 $Y=0.46
+ $X2=2.44 $Y2=0.46
r102 27 33 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.625 $Y=1.79
+ $X2=2.725 $Y2=1.875
r103 27 28 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=2.625 $Y=1.79
+ $X2=0.76 $Y2=1.79
r104 25 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.755
+ $X2=1.32 $Y2=0.755
r105 25 26 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.235 $Y=0.755
+ $X2=0.76 $Y2=0.755
r106 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.595
+ $Y=1.37 $X2=0.595 $Y2=1.37
r107 21 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.635 $Y=1.705
+ $X2=0.76 $Y2=1.79
r108 21 23 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.635 $Y=1.705
+ $X2=0.635 $Y2=1.37
r109 20 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.635 $Y=0.84
+ $X2=0.76 $Y2=0.755
r110 20 23 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=0.635 $Y=0.84
+ $X2=0.635 $Y2=1.37
r111 18 24 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=0.595 $Y=1.84
+ $X2=0.595 $Y2=1.37
r112 18 19 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.665 $Y=1.84
+ $X2=0.665 $Y2=1.99
r113 16 24 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.205
+ $X2=0.595 $Y2=1.37
r114 13 19 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.825 $Y=2.735
+ $X2=0.825 $Y2=1.99
r115 9 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.605 $Y=0.46
+ $X2=0.605 $Y2=1.205
r116 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.62
+ $Y=2.415 $X2=2.76 $Y2=2.56
r117 1 31 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.26
+ $Y=0.25 $X2=2.44 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%A3 2 5 9 11 12 15
c47 12 0 5.5274e-20 $X=1.2 $Y=1.295
r48 15 17 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.095
+ $X2=1.18 $Y2=0.93
r49 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.165
+ $Y=1.095 $X2=1.165 $Y2=1.095
r50 12 16 0.820838 $w=5.08e-07 $l=3.5e-08 $layer=LI1_cond $X=1.2 $Y=1.265
+ $X2=1.165 $Y2=1.265
r51 9 17 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.285 $Y=0.46 $X2=1.285
+ $Y2=0.93
r52 5 11 581.989 $w=1.5e-07 $l=1.135e-06 $layer=POLY_cond $X=1.255 $Y=2.735
+ $X2=1.255 $Y2=1.6
r53 2 11 44.5126 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.18 $Y=1.42 $X2=1.18
+ $Y2=1.6
r54 1 15 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.18 $Y=1.11 $X2=1.18
+ $Y2=1.095
r55 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.18 $Y=1.11 $X2=1.18
+ $Y2=1.42
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%A2 3 7 11 12 13 14 18
c41 13 0 1.22151e-19 $X=1.68 $Y=0.925
c42 7 0 1.51277e-19 $X=1.73 $Y=0.46
c43 3 0 5.5274e-20 $X=1.685 $Y=2.735
r44 13 14 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.707 $Y=0.925
+ $X2=1.707 $Y2=1.295
r45 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.735
+ $Y=1.005 $X2=1.735 $Y2=1.005
r46 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.735 $Y=1.345
+ $X2=1.735 $Y2=1.005
r47 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.735 $Y=1.345
+ $X2=1.735 $Y2=1.51
r48 10 18 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.735 $Y=0.84
+ $X2=1.735 $Y2=1.005
r49 7 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.73 $Y=0.46 $X2=1.73
+ $Y2=0.84
r50 3 12 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=1.685 $Y=2.735
+ $X2=1.685 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%A1 3 7 11 12 15 16 17 18 22
c44 17 0 1.51277e-19 $X=2.16 $Y=0.925
c45 7 0 1.22151e-19 $X=2.185 $Y=0.46
r46 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.275
+ $Y=1.005 $X2=2.275 $Y2=1.005
r47 18 23 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=2.2 $Y=1.295 $X2=2.2
+ $Y2=1.005
r48 17 23 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=2.2 $Y=0.925 $X2=2.2
+ $Y2=1.005
r49 15 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.275 $Y=1.345
+ $X2=2.275 $Y2=1.005
r50 15 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.345
+ $X2=2.275 $Y2=1.51
r51 14 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.84
+ $X2=2.275 $Y2=1.005
r52 11 12 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.165 $Y=1.75
+ $X2=2.165 $Y2=1.9
r53 11 16 93.2903 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=2.2 $Y=1.75 $X2=2.2
+ $Y2=1.51
r54 7 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.185 $Y=0.46
+ $X2=2.185 $Y2=0.84
r55 3 12 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=2.115 $Y=2.735
+ $X2=2.115 $Y2=1.9
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%B1 1 3 6 9 14 15 16 21
r30 21 24 68.9276 $w=6.05e-07 $l=5.05e-07 $layer=POLY_cond $X=2.952 $Y=1.005
+ $X2=2.952 $Y2=1.51
r31 21 23 49.6377 $w=6.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.952 $Y=1.005
+ $X2=2.952 $Y2=0.84
r32 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.135 $Y=1.295
+ $X2=3.135 $Y2=1.665
r33 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.135 $Y=0.925
+ $X2=3.135 $Y2=1.295
r34 14 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.005 $X2=3.09 $Y2=1.005
r35 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.755 $Y=2.215
+ $X2=2.545 $Y2=2.215
r36 9 24 198.946 $w=2.1e-07 $l=6.3e-07 $layer=POLY_cond $X=2.755 $Y=2.14
+ $X2=2.755 $Y2=1.51
r37 6 23 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.725 $Y=0.46
+ $X2=2.725 $Y2=0.84
r38 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.545 $Y=2.29
+ $X2=2.545 $Y2=2.215
r39 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.545 $Y=2.29
+ $X2=2.545 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%X 1 2 7 8 9 10 11 12 13 26 41 44
r21 44 45 4.81525 $w=6.53e-07 $l=1e-08 $layer=LI1_cond $X=0.412 $Y=2.405
+ $X2=0.412 $Y2=2.395
r22 23 37 0.103554 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=0.212 $Y=0.5
+ $X2=0.212 $Y2=0.385
r23 23 26 2.48566 $w=2.53e-07 $l=5.5e-08 $layer=LI1_cond $X=0.212 $Y=0.5
+ $X2=0.212 $Y2=0.555
r24 13 48 3.92606 $w=6.53e-07 $l=2.15e-07 $layer=LI1_cond $X=0.412 $Y=2.775
+ $X2=0.412 $Y2=2.56
r25 12 48 2.15477 $w=6.53e-07 $l=1.18e-07 $layer=LI1_cond $X=0.412 $Y=2.442
+ $X2=0.412 $Y2=2.56
r26 12 44 0.675647 $w=6.53e-07 $l=3.7e-08 $layer=LI1_cond $X=0.412 $Y=2.442
+ $X2=0.412 $Y2=2.405
r27 12 45 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=0.212 $Y=2.357
+ $X2=0.212 $Y2=2.395
r28 11 12 14.5524 $w=2.53e-07 $l=3.22e-07 $layer=LI1_cond $X=0.212 $Y=2.035
+ $X2=0.212 $Y2=2.357
r29 10 11 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.665
+ $X2=0.212 $Y2=2.035
r30 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.295
+ $X2=0.212 $Y2=1.665
r31 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=0.925
+ $X2=0.212 $Y2=1.295
r32 7 41 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=0.385
+ $X2=0.39 $Y2=0.385
r33 7 37 1.40297 $w=2.28e-07 $l=2.8e-08 $layer=LI1_cond $X=0.24 $Y=0.385
+ $X2=0.212 $Y2=0.385
r34 7 8 16.0438 $w=2.53e-07 $l=3.55e-07 $layer=LI1_cond $X=0.212 $Y=0.57
+ $X2=0.212 $Y2=0.925
r35 7 26 0.677908 $w=2.53e-07 $l=1.5e-08 $layer=LI1_cond $X=0.212 $Y=0.57
+ $X2=0.212 $Y2=0.555
r36 2 48 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.485
+ $Y=2.415 $X2=0.61 $Y2=2.56
r37 1 41 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.25 $X2=0.39 $Y2=0.375
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%VPWR 1 2 9 13 16 17 19 20 21 34 35
r37 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r40 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 21 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 19 28 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.775 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 19 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.775 $Y=3.33
+ $X2=1.9 $Y2=3.33
r47 18 31 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 18 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.9 $Y2=3.33
r49 16 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 16 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.91 $Y=3.33 $X2=1.04
+ $Y2=3.33
r51 15 28 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.17 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 15 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.17 $Y=3.33 $X2=1.04
+ $Y2=3.33
r53 11 20 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.9 $Y=3.245
+ $X2=1.9 $Y2=3.33
r54 11 13 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=1.9 $Y=3.245
+ $X2=1.9 $Y2=2.56
r55 7 17 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.04 $Y=3.245
+ $X2=1.04 $Y2=3.33
r56 7 9 30.3624 $w=2.58e-07 $l=6.85e-07 $layer=LI1_cond $X=1.04 $Y=3.245
+ $X2=1.04 $Y2=2.56
r57 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.76
+ $Y=2.415 $X2=1.9 $Y2=2.56
r58 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.9
+ $Y=2.415 $X2=1.04 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%A_266_483# 1 2 9 11 12 15
r25 13 15 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.325 $Y=2.225
+ $X2=2.325 $Y2=2.56
r26 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.195 $Y=2.14
+ $X2=2.325 $Y2=2.225
r27 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.195 $Y=2.14
+ $X2=1.605 $Y2=2.14
r28 7 12 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.472 $Y=2.225
+ $X2=1.605 $Y2=2.14
r29 7 9 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=1.472 $Y=2.225
+ $X2=1.472 $Y2=2.56
r30 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.19
+ $Y=2.415 $X2=2.33 $Y2=2.56
r31 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.33
+ $Y=2.415 $X2=1.47 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_0%VGND 1 2 9 11 13 16 17 18 24 33
r38 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r40 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r42 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 24 32 4.49945 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=3.067
+ $Y2=0
r44 24 29 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.64
+ $Y2=0
r45 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r46 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 18 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r48 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 16 21 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.72
+ $Y2=0
r50 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.9
+ $Y2=0
r51 15 26 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.2
+ $Y2=0
r52 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.9
+ $Y2=0
r53 11 32 3.26672 $w=3.3e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=3.067 $Y2=0
r54 11 13 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.46
r55 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0
r56 7 9 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0.375
r57 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.25 $X2=2.94 $Y2=0.46
r58 1 9 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.68 $Y=0.25
+ $X2=0.9 $Y2=0.375
.ends

