* File: sky130_fd_sc_lp__o21bai_lp.pex.spice
* Created: Fri Aug 28 11:07:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%A1 3 5 8 9 10 11 12 17 20
r30 19 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.485 $Y=1.435
+ $X2=0.5 $Y2=1.435
r31 16 19 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.29 $Y=1.435
+ $X2=0.485 $Y2=1.435
r32 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.435 $X2=0.29 $Y2=1.435
r33 11 12 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=2.035
r34 11 17 8.55038 $w=3.08e-07 $l=2.3e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=1.435
r35 9 10 42.2382 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.547 $Y=1.84
+ $X2=0.547 $Y2=1.99
r36 8 10 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.575 $Y=2.565
+ $X2=0.575 $Y2=1.99
r37 3 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.27 $X2=0.5
+ $Y2=1.435
r38 3 5 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.5 $Y=1.27 $X2=0.5
+ $Y2=0.76
r39 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.6
+ $X2=0.485 $Y2=1.435
r40 1 9 93.2903 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=0.485 $Y=1.6 $X2=0.485
+ $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%A2 3 7 8 9 17 18 19
r40 17 20 30.6647 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.972 $Y=1.435
+ $X2=0.972 $Y2=1.6
r41 17 19 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.972 $Y=1.435
+ $X2=0.972 $Y2=1.27
r42 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.435 $X2=0.95 $Y2=1.435
r43 8 9 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.96 $Y=1.665 $X2=0.96
+ $Y2=2.035
r44 8 18 3.87462 $w=7.08e-07 $l=2.3e-07 $layer=LI1_cond $X=0.96 $Y=1.665
+ $X2=0.96 $Y2=1.435
r45 7 19 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.085 $Y=0.76
+ $X2=1.085 $Y2=1.27
r46 3 20 239.758 $w=2.5e-07 $l=9.65e-07 $layer=POLY_cond $X=1.035 $Y=2.565
+ $X2=1.035 $Y2=1.6
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%A_288_21# 1 2 7 9 12 16 19 24 27 29 32 36
c69 29 0 1.49081e-20 $X=3.16 $Y=1.495
c70 24 0 7.80858e-20 $X=3.16 $Y=1.33
c71 7 0 8.16745e-20 $X=1.515 $Y=1.36
r72 32 34 9.68446 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.08 $Y=0.41 $X2=3.08
+ $Y2=0.61
r73 27 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.495
+ $X2=2.455 $Y2=1.495
r74 26 29 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.62 $Y=1.495
+ $X2=3.16 $Y2=1.495
r75 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.495 $X2=2.62 $Y2=1.495
r76 24 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=1.33
+ $X2=3.16 $Y2=1.495
r77 24 34 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.16 $Y=1.33
+ $X2=3.16 $Y2=0.61
r78 19 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.62 $Y=2.145
+ $X2=2.62 $Y2=2.855
r79 17 26 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=1.66
+ $X2=2.62 $Y2=1.495
r80 17 19 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.62 $Y=1.66
+ $X2=2.62 $Y2=2.145
r81 15 16 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.69 $Y=1.435
+ $X2=1.565 $Y2=1.435
r82 15 36 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.69 $Y=1.435
+ $X2=2.455 $Y2=1.435
r83 10 16 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.565 $Y=1.51
+ $X2=1.565 $Y2=1.435
r84 10 12 262.119 $w=2.5e-07 $l=1.055e-06 $layer=POLY_cond $X=1.565 $Y=1.51
+ $X2=1.565 $Y2=2.565
r85 7 16 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=1.515 $Y=1.36
+ $X2=1.565 $Y2=1.435
r86 7 9 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.515 $Y=1.36 $X2=1.515
+ $Y2=0.76
r87 2 21 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.48 $Y=2
+ $X2=2.62 $Y2=2.855
r88 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48 $Y=2
+ $X2=2.62 $Y2=2.145
r89 1 32 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%B1_N 1 3 6 8 9 10 14 17 19 21 24
c54 24 0 7.80858e-20 $X=2.415 $Y=0.955
c55 1 0 1.49081e-20 $X=2.355 $Y=3.075
r56 24 27 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.415 $Y=0.955
+ $X2=2.415 $Y2=1.015
r57 24 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=0.955
+ $X2=2.415 $Y2=0.79
r58 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=0.955 $X2=2.415 $Y2=0.955
r59 21 25 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.64 $Y=0.955
+ $X2=2.415 $Y2=0.955
r60 18 19 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.865 $Y=1.015
+ $X2=3.1 $Y2=1.015
r61 16 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=1.09 $X2=3.1
+ $Y2=1.015
r62 16 17 1017.84 $w=1.5e-07 $l=1.985e-06 $layer=POLY_cond $X=3.1 $Y=1.09
+ $X2=3.1 $Y2=3.075
r63 12 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=0.94
+ $X2=2.865 $Y2=1.015
r64 12 14 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.865 $Y=0.94
+ $X2=2.865 $Y2=0.445
r65 11 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.015
+ $X2=2.415 $Y2=1.015
r66 10 18 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.79 $Y=1.015
+ $X2=2.865 $Y2=1.015
r67 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.79 $Y=1.015
+ $X2=2.58 $Y2=1.015
r68 8 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.025 $Y=3.15
+ $X2=3.1 $Y2=3.075
r69 8 9 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.025 $Y=3.15
+ $X2=2.48 $Y2=3.15
r70 6 26 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.505 $Y=0.445
+ $X2=2.505 $Y2=0.79
r71 1 9 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=2.355 $Y=3.075
+ $X2=2.48 $Y2=3.15
r72 1 3 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.355 $Y=3.075
+ $X2=2.355 $Y2=2.5
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%VPWR 1 2 7 9 13 15 17 27 28 34
r35 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 25 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r39 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.83 $Y2=3.33
r41 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 18 31 4.66755 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.237 $Y2=3.33
r45 18 20 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=1.83 $Y2=3.33
r47 17 20 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 15 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 15 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=3.245
+ $X2=1.83 $Y2=3.33
r52 11 13 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.83 $Y=3.245
+ $X2=1.83 $Y2=2.87
r53 7 31 3.09863 $w=3.3e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.237 $Y2=3.33
r54 7 9 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.31 $Y=3.245 $X2=0.31
+ $Y2=2.475
r55 2 13 600 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=2.065 $X2=1.83 $Y2=2.87
r56 1 9 300 $w=1.7e-07 $l=4.77022e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.065 $X2=0.31 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%Y 1 2 9 13 16 18 19
r46 19 22 3.22751 $w=6.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.96 $Y=2.035
+ $X2=1.96 $Y2=1.865
r47 18 22 3.79707 $w=6.28e-07 $l=2e-07 $layer=LI1_cond $X=1.96 $Y=1.665 $X2=1.96
+ $Y2=1.865
r48 18 26 6.68592 $w=6.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=1.55
r49 17 19 5.22098 $w=6.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.96 $Y=2.31
+ $X2=1.96 $Y2=2.035
r50 13 26 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.77 $Y=0.76
+ $X2=1.77 $Y2=1.55
r51 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.395
+ $X2=1.3 $Y2=2.395
r52 9 17 10.2785 $w=1.7e-07 $l=3.54965e-07 $layer=LI1_cond $X=1.645 $Y=2.395
+ $X2=1.96 $Y2=2.31
r53 9 10 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.645 $Y=2.395
+ $X2=1.465 $Y2=2.395
r54 2 16 300 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=2.065 $X2=1.3 $Y2=2.475
r55 1 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.55 $X2=1.73 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%A_28_110# 1 2 7 10 15
c23 7 0 8.16745e-20 $X=1.135 $Y=1.015
r24 15 17 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.3 $Y=0.77 $X2=1.3
+ $Y2=1.015
r25 10 12 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.285 $Y=0.77
+ $X2=0.285 $Y2=1.015
r26 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=1.015
+ $X2=0.285 $Y2=1.015
r27 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=1.015
+ $X2=1.3 $Y2=1.015
r28 7 8 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.135 $Y=1.015
+ $X2=0.45 $Y2=1.015
r29 2 15 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.55 $X2=1.3 $Y2=0.77
r30 1 10 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.55 $X2=0.285 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r41 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.29
+ $Y2=0
r46 27 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=3.12
+ $Y2=0
r47 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.8
+ $Y2=0
r50 23 25 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.2
+ $Y2=0
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.29
+ $Y2=0
r52 22 25 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.2
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.8
+ $Y2=0
r56 17 19 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r60 11 13 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.41
r61 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r62 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0.675
r63 2 13 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.235 $X2=2.29 $Y2=0.41
r64 1 9 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.55 $X2=0.8 $Y2=0.675
.ends

