* File: sky130_fd_sc_lp__or4b_1.pex.spice
* Created: Wed Sep  2 10:32:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4B_1%D_N 3 7 9 10 14
r26 14 17 82.2934 $w=5.15e-07 $l=5.05e-07 $layer=POLY_cond $X=0.477 $Y=1.73
+ $X2=0.477 $Y2=2.235
r27 14 16 46.971 $w=5.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.477 $Y=1.73
+ $X2=0.477 $Y2=1.565
r28 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.73 $X2=0.385 $Y2=1.73
r29 10 15 8.89861 $w=3.93e-07 $l=3.05e-07 $layer=LI1_cond $X=0.282 $Y=2.035
+ $X2=0.282 $Y2=1.73
r30 9 15 1.89643 $w=3.93e-07 $l=6.5e-08 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=1.73
r31 7 17 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.66 $Y=2.865
+ $X2=0.66 $Y2=2.235
r32 3 16 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.66 $Y=0.865 $X2=0.66
+ $Y2=1.565
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%A_64_131# 1 2 9 11 13 16 20 23 25
c49 25 0 1.76279e-19 $X=0.77 $Y=1.38
c50 11 0 1.52115e-19 $X=1.44 $Y=1.725
r51 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.38 $X2=1.11 $Y2=1.38
r52 25 27 15.6528 $w=2.65e-07 $l=3.4e-07 $layer=LI1_cond $X=0.77 $Y=1.38
+ $X2=1.11 $Y2=1.38
r53 22 25 1.31371 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.545
+ $X2=0.77 $Y2=1.38
r54 22 23 41.2959 $w=2.38e-07 $l=8.6e-07 $layer=LI1_cond $X=0.77 $Y=1.545
+ $X2=0.77 $Y2=2.405
r55 18 23 22.3775 $w=1.68e-07 $l=3.43e-07 $layer=LI1_cond $X=0.427 $Y=2.49
+ $X2=0.77 $Y2=2.49
r56 18 20 11.3291 $w=2.93e-07 $l=2.9e-07 $layer=LI1_cond $X=0.427 $Y=2.575
+ $X2=0.427 $Y2=2.865
r57 14 25 14.9623 $w=2.65e-07 $l=3.25e-07 $layer=LI1_cond $X=0.445 $Y=1.38
+ $X2=0.77 $Y2=1.38
r58 14 16 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.445 $Y=1.215
+ $X2=0.445 $Y2=0.865
r59 11 28 64.3978 $w=3.37e-07 $l=4.37579e-07 $layer=POLY_cond $X=1.44 $Y=1.725
+ $X2=1.23 $Y2=1.38
r60 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.44 $Y=1.725
+ $X2=1.44 $Y2=2.045
r61 7 28 38.6529 $w=3.37e-07 $l=2.09105e-07 $layer=POLY_cond $X=1.13 $Y=1.215
+ $X2=1.23 $Y2=1.38
r62 7 9 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.13 $Y=1.215 $X2=1.13
+ $Y2=0.865
r63 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.32
+ $Y=2.655 $X2=0.445 $Y2=2.865
r64 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.32
+ $Y=0.655 $X2=0.445 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%C 1 3 4 5 9 12 13 14 15 21
c51 9 0 7.08837e-20 $X=1.91 $Y=2.045
c52 5 0 1.1344e-19 $X=1.635 $Y=1.26
r53 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.89
+ $Y=2.58 $X2=1.89 $Y2=2.58
r54 15 22 4.0213 $w=5.78e-07 $l=1.95e-07 $layer=LI1_cond $X=2.015 $Y=2.775
+ $X2=2.015 $Y2=2.58
r55 14 22 3.60886 $w=5.78e-07 $l=1.75e-07 $layer=LI1_cond $X=2.015 $Y=2.405
+ $X2=2.015 $Y2=2.58
r56 13 14 7.63016 $w=5.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=2.015 $Y2=2.405
r57 12 13 7.63016 $w=5.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.015 $Y=1.665
+ $X2=2.015 $Y2=2.035
r58 11 21 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=2.415
+ $X2=1.89 $Y2=2.58
r59 9 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.91 $Y=2.045
+ $X2=1.91 $Y2=2.415
r60 6 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.91 $Y=1.335 $X2=1.91
+ $Y2=2.045
r61 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.835 $Y=1.26
+ $X2=1.91 $Y2=1.335
r62 4 5 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.835 $Y=1.26 $X2=1.635
+ $Y2=1.26
r63 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.56 $Y=1.185
+ $X2=1.635 $Y2=1.26
r64 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.56 $Y=1.185 $X2=1.56
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%B 4 7 10 11 12 16
c38 12 0 7.25772e-20 $X=2.64 $Y=0.555
c39 4 0 5.93855e-20 $X=2.27 $Y=0.865
r40 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=0.38
+ $X2=2.24 $Y2=0.545
r41 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=0.38 $X2=2.24 $Y2=0.38
r42 12 17 12.8049 $w=3.58e-07 $l=4e-07 $layer=LI1_cond $X=2.64 $Y=0.475 $X2=2.24
+ $Y2=0.475
r43 11 17 2.56098 $w=3.58e-07 $l=8e-08 $layer=LI1_cond $X=2.16 $Y=0.475 $X2=2.24
+ $Y2=0.475
r44 9 10 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.305 $Y=1.555
+ $X2=2.305 $Y2=1.705
r45 7 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.34 $Y=2.045 $X2=2.34
+ $Y2=1.705
r46 4 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.27 $Y=0.865 $X2=2.27
+ $Y2=1.555
r47 4 19 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.27 $Y=0.865
+ $X2=2.27 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%A 3 6 7 8 9 17
r36 14 17 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.56 $Y=2.79 $X2=2.7
+ $Y2=2.79
r37 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=2.79 $X2=2.56 $Y2=2.79
r38 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.605 $Y=2.405
+ $X2=2.605 $Y2=2.775
r39 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.605 $Y=2.035
+ $X2=2.605 $Y2=2.405
r40 3 6 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=2.7 $Y=0.865 $X2=2.7
+ $Y2=2.045
r41 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=2.625 $X2=2.7
+ $Y2=2.79
r42 1 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.7 $Y=2.625 $X2=2.7
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%A_220_367# 1 2 3 10 12 15 18 20 21 25 27 32
+ 37 39 40
c77 32 0 8.04481e-21 $X=1.455 $Y=2.045
c78 27 0 5.93855e-20 $X=2.96 $Y=1.325
c79 18 0 1.52115e-19 $X=1.45 $Y=1.24
c80 15 0 7.25772e-20 $X=3.285 $Y=0.655
r81 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.46 $X2=3.15 $Y2=1.46
r82 35 37 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.345 $Y=0.865
+ $X2=1.45 $Y2=0.865
r83 30 32 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.225 $Y=2.045
+ $X2=1.455 $Y2=2.045
r84 28 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=1.325
+ $X2=2.485 $Y2=1.325
r85 27 44 4.38253 $w=3.53e-07 $l=1.35e-07 $layer=LI1_cond $X=3.137 $Y=1.325
+ $X2=3.137 $Y2=1.46
r86 27 28 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.96 $Y=1.325
+ $X2=2.65 $Y2=1.325
r87 23 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=1.24
+ $X2=2.485 $Y2=1.325
r88 23 25 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.485 $Y=1.24
+ $X2=2.485 $Y2=0.93
r89 22 39 1.44715 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.545 $Y=1.325
+ $X2=1.455 $Y2=1.325
r90 21 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=1.325
+ $X2=2.485 $Y2=1.325
r91 21 22 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.32 $Y=1.325
+ $X2=1.545 $Y2=1.325
r92 20 32 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=1.88
+ $X2=1.455 $Y2=2.045
r93 19 39 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.325
r94 19 20 28.9596 $w=1.78e-07 $l=4.7e-07 $layer=LI1_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.88
r95 18 39 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.45 $Y=1.24
+ $X2=1.455 $Y2=1.325
r96 17 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=1.03
+ $X2=1.45 $Y2=0.865
r97 17 18 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.45 $Y=1.03
+ $X2=1.45 $Y2=1.24
r98 13 45 38.7956 $w=3.51e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.285 $Y=1.295
+ $X2=3.19 $Y2=1.46
r99 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.285 $Y=1.295
+ $X2=3.285 $Y2=0.655
r100 10 45 57.3341 $w=3.51e-07 $l=3.17017e-07 $layer=POLY_cond $X=3.225 $Y=1.76
+ $X2=3.19 $Y2=1.46
r101 10 12 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.225 $Y=1.76
+ $X2=3.225 $Y2=2.465
r102 3 30 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.835 $X2=1.225 $Y2=2.045
r103 2 25 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.655 $X2=2.485 $Y2=0.93
r104 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.205
+ $Y=0.655 $X2=1.345 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%VPWR 1 2 9 13 18 19 21 22 23 36 37
r37 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r38 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 30 33 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 27 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 23 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 23 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 21 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 21 22 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=3.035 $Y2=3.33
r48 20 36 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 20 22 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.035 $Y2=3.33
r50 18 26 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 18 19 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.892 $Y2=3.33
r52 17 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.04 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 17 19 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.892 $Y2=3.33
r54 13 16 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=3.035 $Y=1.98
+ $X2=3.035 $Y2=2.95
r55 11 22 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=3.245
+ $X2=3.035 $Y2=3.33
r56 11 16 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.035 $Y=3.245
+ $X2=3.035 $Y2=2.95
r57 7 19 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.892 $Y=3.245
+ $X2=0.892 $Y2=3.33
r58 7 9 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=0.892 $Y=3.245
+ $X2=0.892 $Y2=2.91
r59 2 16 400 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=3.01 $Y2=2.95
r60 2 13 400 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=3.01 $Y2=1.98
r61 1 9 600 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=2.655 $X2=0.875 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%X 1 2 7 8 9 10 11 12 13 25 38 48 52
r18 52 53 5.99337 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=1.98
+ $X2=3.545 $Y2=1.815
r19 36 38 0.274391 $w=4.18e-07 $l=1e-08 $layer=LI1_cond $X=3.545 $Y=2.025
+ $X2=3.545 $Y2=2.035
r20 23 48 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=3.58 $Y=0.92 $X2=3.58
+ $Y2=0.925
r21 13 45 3.70428 $w=4.18e-07 $l=1.35e-07 $layer=LI1_cond $X=3.545 $Y=2.775
+ $X2=3.545 $Y2=2.91
r22 12 13 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.545 $Y=2.405
+ $X2=3.545 $Y2=2.775
r23 11 36 1.04269 $w=4.18e-07 $l=3.8e-08 $layer=LI1_cond $X=3.545 $Y=1.987
+ $X2=3.545 $Y2=2.025
r24 11 52 0.192074 $w=4.18e-07 $l=7e-09 $layer=LI1_cond $X=3.545 $Y=1.987
+ $X2=3.545 $Y2=1.98
r25 11 12 9.13723 $w=4.18e-07 $l=3.33e-07 $layer=LI1_cond $X=3.545 $Y=2.072
+ $X2=3.545 $Y2=2.405
r26 11 38 1.01525 $w=4.18e-07 $l=3.7e-08 $layer=LI1_cond $X=3.545 $Y=2.072
+ $X2=3.545 $Y2=2.035
r27 10 53 6.40246 $w=2.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.62 $Y=1.665
+ $X2=3.62 $Y2=1.815
r28 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.62 $Y=1.295
+ $X2=3.62 $Y2=1.665
r29 9 50 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=3.62 $Y=1.295 $X2=3.62
+ $Y2=1.095
r30 8 50 4.91241 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=3.58 $Y=0.965
+ $X2=3.58 $Y2=1.095
r31 8 48 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=3.58 $Y=0.965 $X2=3.58
+ $Y2=0.925
r32 8 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=3.58 $Y=0.88 $X2=3.58
+ $Y2=0.92
r33 7 8 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=3.58 $Y=0.555
+ $X2=3.58 $Y2=0.88
r34 7 25 4.44514 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.58 $Y=0.555
+ $X2=3.58 $Y2=0.42
r35 2 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.835 $X2=3.44 $Y2=1.98
r36 2 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.835 $X2=3.44 $Y2=2.91
r37 1 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.36
+ $Y=0.235 $X2=3.5 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_1%VGND 1 2 3 12 16 20 25 26 28 29 30 39 45 46
+ 49
r51 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 46 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r53 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r54 43 49 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.065
+ $Y2=0
r55 43 45 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.6
+ $Y2=0
r56 42 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r57 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r58 39 49 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=3.065
+ $Y2=0
r59 39 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=2.64
+ $Y2=0
r60 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r61 34 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r62 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r63 30 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r64 30 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r65 28 37 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.68
+ $Y2=0
r66 28 29 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.805
+ $Y2=0
r67 27 41 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.64
+ $Y2=0
r68 27 29 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.805
+ $Y2=0
r69 25 33 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.78 $Y=0 $X2=0.72
+ $Y2=0
r70 25 26 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.78 $Y=0 $X2=0.895
+ $Y2=0
r71 24 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.68
+ $Y2=0
r72 24 26 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.895
+ $Y2=0
r73 20 22 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=3.065 $Y=0.38
+ $X2=3.065 $Y2=0.905
r74 18 49 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0
r75 18 20 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0.38
r76 14 29 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0.085
+ $X2=1.805 $Y2=0
r77 14 16 43.2545 $w=1.98e-07 $l=7.8e-07 $layer=LI1_cond $X=1.805 $Y=0.085
+ $X2=1.805 $Y2=0.865
r78 10 26 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0
r79 10 12 39.0829 $w=2.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0.865
r80 3 22 182 $w=1.7e-07 $l=3.4821e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.655 $X2=3.01 $Y2=0.905
r81 3 20 182 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.655 $X2=3.07 $Y2=0.38
r82 2 16 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.655 $X2=1.79 $Y2=0.865
r83 1 12 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.735
+ $Y=0.655 $X2=0.895 $Y2=0.865
.ends

