* File: sky130_fd_sc_lp__nor4bb_2.pex.spice
* Created: Fri Aug 28 10:59:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%C_N 3 6 9 11 12 13 17
r33 17 19 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.687 $Y=1.745
+ $X2=0.687 $Y2=1.58
r34 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.745 $Y2=2.035
r35 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.72
+ $Y=1.745 $X2=0.72 $Y2=1.745
r36 9 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.585 $Y=2.77
+ $X2=0.585 $Y2=2.25
r37 6 11 46.9352 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.687 $Y=2.053
+ $X2=0.687 $Y2=2.25
r38 5 17 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.687 $Y=1.777
+ $X2=0.687 $Y2=1.745
r39 5 6 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.687 $Y=1.777
+ $X2=0.687 $Y2=2.053
r40 3 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.565 $Y=1.03
+ $X2=0.565 $Y2=1.58
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%D_N 3 7 11 12 13 14 15 20
c38 13 0 2.06186e-20 $X=1.2 $Y=1.665
r39 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.335
+ $Y=1.745 $X2=1.335 $Y2=1.745
r40 14 15 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.237 $Y=2.035
+ $X2=1.237 $Y2=2.405
r41 14 21 9.1564 $w=3.63e-07 $l=2.9e-07 $layer=LI1_cond $X=1.237 $Y=2.035
+ $X2=1.237 $Y2=1.745
r42 13 21 2.5259 $w=3.63e-07 $l=8e-08 $layer=LI1_cond $X=1.237 $Y=1.665
+ $X2=1.237 $Y2=1.745
r43 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.335 $Y=2.085
+ $X2=1.335 $Y2=1.745
r44 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=2.085
+ $X2=1.335 $Y2=2.25
r45 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.58
+ $X2=1.335 $Y2=1.745
r46 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.425 $Y=1.03
+ $X2=1.425 $Y2=1.58
r47 3 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.355 $Y=2.77
+ $X2=1.355 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%A_286_512# 1 2 7 9 11 14 16 18 20 23 25 26
+ 27 32 36 39 40
c77 40 0 2.06186e-20 $X=2.04 $Y=1.095
c78 23 0 6.06445e-20 $X=3.085 $Y=2.405
r79 42 43 17.435 $w=3.98e-07 $l=4.7e-07 $layer=LI1_cond $X=2.005 $Y=1.13
+ $X2=2.005 $Y2=1.6
r80 40 46 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.095
+ $X2=2.04 $Y2=1.26
r81 39 42 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=2.005 $Y=1.095
+ $X2=2.005 $Y2=1.13
r82 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.04
+ $Y=1.095 $X2=2.04 $Y2=1.095
r83 34 36 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.57 $Y=2.835
+ $X2=1.89 $Y2=2.835
r84 32 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=2.67
+ $X2=1.89 $Y2=2.835
r85 32 43 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=1.89 $Y=2.67
+ $X2=1.89 $Y2=1.6
r86 27 42 3.25816 $w=2.6e-07 $l=2e-07 $layer=LI1_cond $X=1.805 $Y=1.13 $X2=2.005
+ $Y2=1.13
r87 27 29 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=1.13
+ $X2=1.64 $Y2=1.13
r88 21 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.085 $Y=1.335
+ $X2=3.085 $Y2=1.26
r89 21 23 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=3.085 $Y=1.335
+ $X2=3.085 $Y2=2.405
r90 18 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.085 $Y=1.185
+ $X2=3.085 $Y2=1.26
r91 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.085 $Y=1.185
+ $X2=3.085 $Y2=0.655
r92 17 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.73 $Y=1.26 $X2=2.655
+ $Y2=1.26
r93 16 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.01 $Y=1.26
+ $X2=3.085 $Y2=1.26
r94 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.01 $Y=1.26
+ $X2=2.73 $Y2=1.26
r95 12 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.335
+ $X2=2.655 $Y2=1.26
r96 12 14 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.655 $Y=1.335
+ $X2=2.655 $Y2=2.405
r97 9 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.185 $X2=2.655
+ $Y2=1.26
r98 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.655 $Y=1.185
+ $X2=2.655 $Y2=0.655
r99 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.26
+ $X2=2.04 $Y2=1.26
r100 7 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.26 $X2=2.655
+ $Y2=1.26
r101 7 8 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.58 $Y=1.26
+ $X2=2.205 $Y2=1.26
r102 2 34 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=2.56 $X2=1.57 $Y2=2.835
r103 1 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.82 $X2=1.64 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%A_45_164# 1 2 9 13 17 21 25 29 32 33 34 36
+ 37 39 42 44 45 51
c111 34 0 1.23009e-19 $X=1.295 $Y=0.745
c112 17 0 1.65947e-19 $X=3.945 $Y=0.655
r113 50 51 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.945 $Y=1.42
+ $X2=3.985 $Y2=1.42
r114 44 45 6.95017 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.325 $Y=2.77
+ $X2=0.325 $Y2=2.605
r115 40 50 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.66 $Y=1.42
+ $X2=3.945 $Y2=1.42
r116 40 47 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.66 $Y=1.42
+ $X2=3.515 $Y2=1.42
r117 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.42 $X2=3.66 $Y2=1.42
r118 37 39 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.555 $Y=1.42
+ $X2=3.66 $Y2=1.42
r119 36 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.47 $Y=1.335
+ $X2=2.555 $Y2=1.42
r120 35 36 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.47 $Y=0.83
+ $X2=2.47 $Y2=1.335
r121 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.385 $Y=0.745
+ $X2=2.47 $Y2=0.83
r122 33 34 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=2.385 $Y=0.745
+ $X2=1.295 $Y2=0.745
r123 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=0.83
+ $X2=1.295 $Y2=0.745
r124 31 32 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.21 $Y=0.83
+ $X2=1.21 $Y2=1.24
r125 30 42 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.435 $Y=1.325
+ $X2=0.31 $Y2=1.325
r126 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.125 $Y=1.325
+ $X2=1.21 $Y2=1.24
r127 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.125 $Y=1.325
+ $X2=0.435 $Y2=1.325
r128 27 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=1.41
+ $X2=0.31 $Y2=1.325
r129 27 45 55.0868 $w=2.48e-07 $l=1.195e-06 $layer=LI1_cond $X=0.31 $Y=1.41
+ $X2=0.31 $Y2=2.605
r130 23 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=1.24
+ $X2=0.31 $Y2=1.325
r131 23 25 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=0.31 $Y=1.24
+ $X2=0.31 $Y2=1.03
r132 19 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.585
+ $X2=3.985 $Y2=1.42
r133 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.985 $Y=1.585
+ $X2=3.985 $Y2=2.405
r134 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.255
+ $X2=3.945 $Y2=1.42
r135 15 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.945 $Y=1.255
+ $X2=3.945 $Y2=0.655
r136 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.585
+ $X2=3.515 $Y2=1.42
r137 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.515 $Y=1.585
+ $X2=3.515 $Y2=2.405
r138 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.255
+ $X2=3.515 $Y2=1.42
r139 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.515 $Y=1.255 $X2=3.515
+ $Y2=0.655
r140 2 44 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=2.56 $X2=0.37 $Y2=2.77
r141 1 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.82 $X2=0.35 $Y2=1.03
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%B 1 3 4 6 7 9 10 12 13 20
c52 13 0 1.65947e-19 $X=4.56 $Y=1.295
c53 1 0 8.51735e-20 $X=4.855 $Y=1.185
r54 20 21 8.6264 $w=4.47e-07 $l=8e-08 $layer=POLY_cond $X=5.285 $Y=1.455
+ $X2=5.365 $Y2=1.455
r55 19 20 37.7405 $w=4.47e-07 $l=3.5e-07 $layer=POLY_cond $X=4.935 $Y=1.455
+ $X2=5.285 $Y2=1.455
r56 18 19 8.6264 $w=4.47e-07 $l=8e-08 $layer=POLY_cond $X=4.855 $Y=1.455
+ $X2=4.935 $Y2=1.455
r57 16 18 25.34 $w=4.47e-07 $l=2.35e-07 $layer=POLY_cond $X=4.62 $Y=1.455
+ $X2=4.855 $Y2=1.455
r58 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.62
+ $Y=1.35 $X2=4.62 $Y2=1.35
r59 10 21 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.365 $Y=1.725
+ $X2=5.365 $Y2=1.455
r60 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.365 $Y=1.725
+ $X2=5.365 $Y2=2.465
r61 7 20 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.285 $Y=1.185
+ $X2=5.285 $Y2=1.455
r62 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.285 $Y=1.185
+ $X2=5.285 $Y2=0.655
r63 4 19 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.935 $Y=1.725
+ $X2=4.935 $Y2=1.455
r64 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.935 $Y=1.725
+ $X2=4.935 $Y2=2.465
r65 1 18 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.855 $Y=1.185
+ $X2=4.855 $Y2=1.455
r66 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.855 $Y=1.185
+ $X2=4.855 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%A 1 3 6 8 10 13 15 20
c36 20 0 1.37468e-20 $X=6.225 $Y=1.35
r37 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.315
+ $Y=1.35 $X2=6.315 $Y2=1.35
r38 20 22 13.9038 $w=3.12e-07 $l=9e-08 $layer=POLY_cond $X=6.225 $Y=1.35
+ $X2=6.315 $Y2=1.35
r39 19 20 12.359 $w=3.12e-07 $l=8e-08 $layer=POLY_cond $X=6.145 $Y=1.35
+ $X2=6.225 $Y2=1.35
r40 18 19 54.0705 $w=3.12e-07 $l=3.5e-07 $layer=POLY_cond $X=5.795 $Y=1.35
+ $X2=6.145 $Y2=1.35
r41 15 23 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=1.35
+ $X2=6.315 $Y2=1.35
r42 11 20 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.515
+ $X2=6.225 $Y2=1.35
r43 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.225 $Y=1.515
+ $X2=6.225 $Y2=2.465
r44 8 19 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.145 $Y=1.185
+ $X2=6.145 $Y2=1.35
r45 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.145 $Y=1.185
+ $X2=6.145 $Y2=0.655
r46 4 18 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=1.515
+ $X2=5.795 $Y2=1.35
r47 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.795 $Y=1.515
+ $X2=5.795 $Y2=2.465
r48 1 18 12.359 $w=3.12e-07 $l=2.0106e-07 $layer=POLY_cond $X=5.715 $Y=1.185
+ $X2=5.795 $Y2=1.35
r49 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.715 $Y=1.185
+ $X2=5.715 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%VPWR 1 2 9 13 15 20 30 31 34 41
r63 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r64 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r65 34 37 9.72929 $w=6.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.97 $Y=2.785
+ $X2=0.97 $Y2=3.33
r66 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r67 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r68 28 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.01 $Y2=3.33
r69 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.48 $Y2=3.33
r70 27 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r71 26 27 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r72 24 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 23 26 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=5.52 $Y2=3.33
r74 23 24 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 21 37 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=0.97 $Y2=3.33
r76 21 23 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 20 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6.01 $Y2=3.33
r78 20 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 18 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r80 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 15 37 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.97 $Y2=3.33
r82 15 17 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r83 13 27 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=5.52 $Y2=3.33
r84 13 24 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 9 12 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=6.01 $Y=2.11 $X2=6.01
+ $Y2=2.95
r86 7 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245 $X2=6.01
+ $Y2=3.33
r87 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.95
r88 2 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=1.835 $X2=6.01 $Y2=2.95
r89 2 9 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=1.835 $X2=6.01 $Y2=2.11
r90 1 34 300 $w=1.7e-07 $l=5.81722e-07 $layer=licon1_PDIFF $count=2 $X=0.66
+ $Y=2.56 $X2=1.14 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%A_463_355# 1 2 3 12 16 17 18 22 29
r34 23 27 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.415 $Y=2.1
+ $X2=3.31 $Y2=2.1
r35 22 29 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.085 $Y=2.1
+ $X2=4.225 $Y2=2.1
r36 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.085 $Y=2.1
+ $X2=3.415 $Y2=2.1
r37 19 21 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=3.31 $Y=2.905
+ $X2=3.31 $Y2=2.88
r38 18 27 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.185
+ $X2=3.31 $Y2=2.1
r39 18 21 36.7056 $w=2.08e-07 $l=6.95e-07 $layer=LI1_cond $X=3.31 $Y=2.185
+ $X2=3.31 $Y2=2.88
r40 16 19 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.205 $Y=2.99
+ $X2=3.31 $Y2=2.905
r41 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.205 $Y=2.99
+ $X2=2.535 $Y2=2.99
r42 12 15 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=2.405 $Y=1.92
+ $X2=2.405 $Y2=2.89
r43 10 17 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.405 $Y=2.905
+ $X2=2.535 $Y2=2.99
r44 10 15 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=2.405 $Y=2.905
+ $X2=2.405 $Y2=2.89
r45 3 29 300 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=2 $X=4.06
+ $Y=1.775 $X2=4.2 $Y2=2.18
r46 2 27 400 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.775 $X2=3.3 $Y2=2.18
r47 2 21 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.775 $X2=3.3 $Y2=2.88
r48 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.775 $X2=2.44 $Y2=2.89
r49 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.775 $X2=2.44 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%Y 1 2 3 4 5 18 24 27 30 32 36 38 42 44 45
+ 51 52 53 60 65 69 74
c96 45 0 1.37468e-20 $X=5.025 $Y=0.927
c97 38 0 8.51735e-20 $X=5.835 $Y=1.15
r98 73 74 6.6234 $w=3.23e-07 $l=1.18e-07 $layer=LI1_cond $X=4.112 $Y=1.002
+ $X2=4.23 $Y2=1.002
r99 60 65 0.490401 $w=2.33e-07 $l=1e-08 $layer=LI1_cond $X=4.112 $Y=1.675
+ $X2=4.112 $Y2=1.665
r100 59 73 2.65601 $w=2.35e-07 $l=1.63e-07 $layer=LI1_cond $X=4.112 $Y=1.165
+ $X2=4.112 $Y2=1.002
r101 53 60 2.96548 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.112 $Y=1.76
+ $X2=4.112 $Y2=1.675
r102 53 65 1.86352 $w=2.33e-07 $l=3.8e-08 $layer=LI1_cond $X=4.112 $Y=1.627
+ $X2=4.112 $Y2=1.665
r103 52 53 16.2813 $w=2.33e-07 $l=3.32e-07 $layer=LI1_cond $X=4.112 $Y=1.295
+ $X2=4.112 $Y2=1.627
r104 52 59 6.37522 $w=2.33e-07 $l=1.3e-07 $layer=LI1_cond $X=4.112 $Y=1.295
+ $X2=4.112 $Y2=1.165
r105 51 73 1.13471 $w=3.23e-07 $l=3.2e-08 $layer=LI1_cond $X=4.08 $Y=1.002
+ $X2=4.112 $Y2=1.002
r106 48 49 9.05491 $w=2.78e-07 $l=2.2e-07 $layer=LI1_cond $X=5.025 $Y=0.93
+ $X2=5.025 $Y2=1.15
r107 45 48 0.123476 $w=2.78e-07 $l=3e-09 $layer=LI1_cond $X=5.025 $Y=0.927
+ $X2=5.025 $Y2=0.93
r108 45 46 4.77808 $w=2.78e-07 $l=8.7e-08 $layer=LI1_cond $X=5.025 $Y=0.927
+ $X2=5.025 $Y2=0.84
r109 44 53 46.2481 $w=2.43e-07 $l=9.6e-07 $layer=LI1_cond $X=3.035 $Y=1.76
+ $X2=3.995 $Y2=1.76
r110 40 42 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=5.93 $Y=1.065
+ $X2=5.93 $Y2=0.42
r111 39 49 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.165 $Y=1.15
+ $X2=5.025 $Y2=1.15
r112 38 40 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.835 $Y=1.15
+ $X2=5.93 $Y2=1.065
r113 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.835 $Y=1.15
+ $X2=5.165 $Y2=1.15
r114 36 46 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=5.07 $Y=0.42
+ $X2=5.07 $Y2=0.84
r115 32 45 3.50883 $w=1.75e-07 $l=1.4e-07 $layer=LI1_cond $X=4.885 $Y=0.927
+ $X2=5.025 $Y2=0.927
r116 32 74 41.5117 $w=1.73e-07 $l=6.55e-07 $layer=LI1_cond $X=4.885 $Y=0.927
+ $X2=4.23 $Y2=0.927
r117 28 51 12.4109 $w=3.23e-07 $l=3.5e-07 $layer=LI1_cond $X=3.73 $Y=1.002
+ $X2=4.08 $Y2=1.002
r118 28 69 5.97798 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=3.73 $Y=1.002
+ $X2=3.635 $Y2=1.002
r119 28 30 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=3.73 $Y=0.84
+ $X2=3.73 $Y2=0.42
r120 27 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.965 $Y=1.08
+ $X2=3.635 $Y2=1.08
r121 22 27 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.87 $Y=0.995
+ $X2=2.965 $Y2=1.08
r122 22 24 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.42
r123 18 20 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=2.87 $Y=1.92
+ $X2=2.87 $Y2=2.65
r124 16 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.87 $Y=1.845
+ $X2=3.035 $Y2=1.76
r125 16 18 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.87 $Y=1.845
+ $X2=2.87 $Y2=1.92
r126 5 20 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.775 $X2=2.87 $Y2=2.65
r127 5 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.775 $X2=2.87 $Y2=1.92
r128 4 42 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.79
+ $Y=0.235 $X2=5.93 $Y2=0.42
r129 3 48 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.235 $X2=5.07 $Y2=0.93
r130 3 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.235 $X2=5.07 $Y2=0.42
r131 2 28 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.235 $X2=3.73 $Y2=0.93
r132 2 30 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.235 $X2=3.73 $Y2=0.42
r133 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.73
+ $Y=0.235 $X2=2.87 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%A_718_355# 1 2 9 11 12 13 15
c29 12 0 6.06445e-20 $X=3.915 $Y=2.99
r30 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=2.905 $X2=5.15
+ $Y2=2.99
r31 13 15 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=5.15 $Y=2.905
+ $X2=5.15 $Y2=2.11
r32 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=2.99
+ $X2=5.15 $Y2=2.99
r33 11 12 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.985 $Y=2.99
+ $X2=3.915 $Y2=2.99
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.75 $Y=2.905
+ $X2=3.915 $Y2=2.99
r35 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.75 $Y=2.905
+ $X2=3.75 $Y2=2.46
r36 2 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.835 $X2=5.15 $Y2=2.91
r37 2 15 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.835 $X2=5.15 $Y2=2.11
r38 1 9 300 $w=1.7e-07 $l=7.60805e-07 $layer=licon1_PDIFF $count=2 $X=3.59
+ $Y=1.775 $X2=3.75 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%A_919_367# 1 2 3 12 14 15 18 22 26 30
r39 26 28 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=6.475 $Y=1.98
+ $X2=6.475 $Y2=2.91
r40 24 26 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=6.475 $Y=1.855
+ $X2=6.475 $Y2=1.98
r41 23 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.675 $Y=1.77
+ $X2=5.58 $Y2=1.77
r42 22 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.345 $Y=1.77
+ $X2=6.475 $Y2=1.855
r43 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.345 $Y=1.77
+ $X2=5.675 $Y2=1.77
r44 18 20 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=5.58 $Y=1.98
+ $X2=5.58 $Y2=2.91
r45 16 30 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=1.855
+ $X2=5.58 $Y2=1.77
r46 16 18 7.29665 $w=1.88e-07 $l=1.25e-07 $layer=LI1_cond $X=5.58 $Y=1.855
+ $X2=5.58 $Y2=1.98
r47 14 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.485 $Y=1.77
+ $X2=5.58 $Y2=1.77
r48 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.485 $Y=1.77
+ $X2=4.815 $Y2=1.77
r49 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.685 $Y=1.855
+ $X2=4.815 $Y2=1.77
r50 10 12 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=4.685 $Y=1.855
+ $X2=4.685 $Y2=1.98
r51 3 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.835 $X2=6.44 $Y2=2.91
r52 3 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.835 $X2=6.44 $Y2=1.98
r53 2 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.44
+ $Y=1.835 $X2=5.58 $Y2=2.91
r54 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.44
+ $Y=1.835 $X2=5.58 $Y2=1.98
r55 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.595
+ $Y=1.835 $X2=4.72 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_2%VGND 1 2 3 4 5 6 21 25 29 33 35 37 40 41 43
+ 44 45 47 66 71 77 82 88 90 94
c93 1 0 1.23009e-19 $X=0.64 $Y=0.82
r94 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r95 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r96 87 88 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=0.292
+ $X2=4.805 $Y2=0.292
r97 84 87 1.26737 $w=7.53e-07 $l=8e-08 $layer=LI1_cond $X=4.56 $Y=0.292 $X2=4.64
+ $Y2=0.292
r98 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r99 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r100 80 84 7.60421 $w=7.53e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=0.292
+ $X2=4.56 $Y2=0.292
r101 80 82 9.88706 $w=7.53e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=0.292
+ $X2=3.995 $Y2=0.292
r102 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r103 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r104 75 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r105 75 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r106 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r107 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.5
+ $Y2=0
r108 72 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=6
+ $Y2=0
r109 71 93 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=6.195 $Y=0
+ $X2=6.457 $Y2=0
r110 71 74 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6
+ $Y2=0
r111 70 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r112 70 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r113 69 88 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.04 $Y=0
+ $X2=4.805 $Y2=0
r114 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r115 66 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.5
+ $Y2=0
r116 66 69 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.04
+ $Y2=0
r117 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r118 64 82 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.995
+ $Y2=0
r119 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r120 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r121 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r122 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r123 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r124 55 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r125 54 57 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r126 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r127 52 77 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.785
+ $Y2=0
r128 52 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r129 50 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r130 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r131 47 77 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.785
+ $Y2=0
r132 47 49 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r133 45 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r134 45 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r135 43 60 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.12
+ $Y2=0
r136 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.3
+ $Y2=0
r137 42 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.6
+ $Y2=0
r138 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.3
+ $Y2=0
r139 40 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.275 $Y=0
+ $X2=2.16 $Y2=0
r140 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.44
+ $Y2=0
r141 39 60 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.605 $Y=0
+ $X2=3.12 $Y2=0
r142 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=2.44
+ $Y2=0
r143 35 93 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.457 $Y2=0
r144 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.36 $Y2=0.38
r145 31 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r146 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.38
r147 27 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.085 $X2=3.3
+ $Y2=0
r148 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0.36
r149 23 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.085
+ $X2=2.44 $Y2=0
r150 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.44 $Y=0.085
+ $X2=2.44 $Y2=0.38
r151 19 77 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r152 19 21 29.6585 $w=3.38e-07 $l=8.75e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.96
r153 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.22
+ $Y=0.235 $X2=6.36 $Y2=0.38
r154 5 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.235 $X2=5.5 $Y2=0.38
r155 4 87 91 $w=1.7e-07 $l=7.59342e-07 $layer=licon1_NDIFF $count=2 $X=4.02
+ $Y=0.235 $X2=4.64 $Y2=0.545
r156 3 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.16
+ $Y=0.235 $X2=3.3 $Y2=0.36
r157 2 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.235 $X2=2.44 $Y2=0.38
r158 1 21 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.82 $X2=0.79 $Y2=0.96
.ends

