* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a311oi_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_158_473# A3 VPWR VPB phighvt w=640000u l=150000u
+  ad=4.096e+11p pd=3.84e+06u as=3.488e+11p ps=3.65e+06u
M1001 a_158_473# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_432_473# B1 a_158_473# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1003 Y A1 a_252_47# VNB nshort w=420000u l=150000u
+  ad=2.415e+11p pd=2.83e+06u as=8.82e+10p ps=1.26e+06u
M1004 Y C1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=5.145e+11p ps=4.13e+06u
M1005 VPWR A2 a_158_473# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_180_47# A3 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_252_47# A2 a_180_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y C1 a_432_473# VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1009 VGND B1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
