* File: sky130_fd_sc_lp__sdfrtp_ov2.spice
* Created: Fri Aug 28 11:28:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrtp_ov2.pex.spice"
.subckt sky130_fd_sc_lp__sdfrtp_ov2  VNB VPB SCE D SCD RESET_B CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_SCE_M1024_g N_A_35_74#_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 noxref_25 N_A_35_74#_M1005_g N_noxref_24_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1034 N_A_380_50#_M1034_d N_D_M1034_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.129575 AS=0.0441 PD=1.085 PS=0.63 NRD=34.284 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1038 noxref_26 N_SCE_M1038_g N_A_380_50#_M1034_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.129575 PD=0.63 PS=1.085 NRD=14.28 NRS=32.856 M=1 R=2.8
+ SA=75000.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_noxref_24_M1000_d N_SCD_M1000_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.0441 PD=0.745 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_RESET_B_M1026_g N_noxref_24_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.126 AS=0.06825 PD=1.44 PS=0.745 NRD=9.996 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 N_A_809_463#_M1033_d N_A_865_255#_M1033_g N_A_380_50#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1554 PD=0.7 PS=1.58 NRD=0 NRS=30 M=1 R=2.8
+ SA=75000.3 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1035 A_991_119# N_A_757_317#_M1035_g N_A_809_463#_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1009 A_1085_119# N_A_937_333#_M1009_g A_991_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0672 PD=0.81 PS=0.74 NRD=37.14 NRS=30 M=1 R=2.8 SA=75001.2
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_RESET_B_M1036_g A_1085_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.10815 AS=0.0777 PD=0.935 PS=0.81 NRD=67.14 NRS=37.14 M=1 R=2.8 SA=75001.6
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_937_333#_M1010_d N_A_809_463#_M1010_g N_VGND_M1036_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.09975 AS=0.10815 PD=0.895 PS=0.935 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75003 A=0.063 P=1.14 MULT=1
MM1028 N_A_1445_113#_M1028_d N_A_757_317#_M1028_g N_A_937_333#_M1010_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.1302 AS=0.09975 PD=1.04 PS=0.895 NRD=0 NRS=55.704
+ M=1 R=2.8 SA=75002.9 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1011 A_1599_113# N_A_865_255#_M1011_g N_A_1445_113#_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1302 PD=0.63 PS=1.04 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75003.7 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1641_21#_M1020_g A_1599_113# VNB NSHORT L=0.15 W=0.42
+ AD=0.1266 AS=0.0441 PD=1.035 PS=0.63 NRD=45.708 NRS=14.28 M=1 R=2.8 SA=75004
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 A_1818_119# N_RESET_B_M1004_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1266 PD=0.63 PS=1.035 NRD=14.28 NRS=41.424 M=1 R=2.8 SA=75004.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_1641_21#_M1008_d N_A_1445_113#_M1008_g A_1818_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_A_865_255#_M1030_g N_A_757_317#_M1030_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1766 AS=0.1197 PD=1.425 PS=1.41 NRD=104.412 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1018 N_A_865_255#_M1018_d N_CLK_M1018_g N_VGND_M1030_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.1766 PD=1.41 PS=1.425 NRD=0 NRS=104.412 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_A_1445_113#_M1039_g N_A_2408_367#_M1039_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0854 AS=0.1113 PD=0.8 PS=1.37 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_Q_M1016_d N_A_2408_367#_M1016_g N_VGND_M1039_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1708 PD=2.21 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.4 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_SCE_M1012_g N_A_35_74#_M1012_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.115623 AS=0.3872 PD=1.16528 PS=2.49 NRD=13.8491 NRS=0 M=1 R=4.26667
+ SA=75000.5 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1001 A_355_463# N_SCE_M1001_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0758774 PD=0.63 PS=0.764717 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001
+ SB=75003.8 A=0.063 P=1.14 MULT=1
MM1027 N_A_380_50#_M1027_d N_D_M1027_g A_355_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.4
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1015 A_513_463# N_A_35_74#_M1015_g N_A_380_50#_M1027_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=49.25 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_SCD_M1006_g A_513_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1178 AS=0.0672 PD=1.07 PS=0.74 NRD=30.4759 NRS=49.25 M=1 R=2.8 SA=75002.3
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1025 N_A_380_50#_M1025_d N_RESET_B_M1025_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1178 PD=0.7 PS=1.07 NRD=0 NRS=105.75 M=1 R=2.8
+ SA=75002.8 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1019 N_A_809_463#_M1019_d N_A_757_317#_M1019_g N_A_380_50#_M1025_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.3 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1037 A_895_463# N_A_865_255#_M1037_g N_A_809_463#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75003.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_937_333#_M1002_g A_895_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=25.7873 NRS=23.443 M=1 R=2.8
+ SA=75004.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_809_463#_M1013_d N_RESET_B_M1013_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=25.7873 M=1 R=2.8
+ SA=75004.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_A_937_333#_M1029_d N_A_809_463#_M1029_g N_VPWR_M1029_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.33185 PD=0.7 PS=2.77 NRD=0 NRS=344.789 M=1 R=2.8
+ SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_1445_113#_M1017_d N_A_865_255#_M1017_g N_A_937_333#_M1029_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.208425 AS=0.0588 PD=1.66 PS=0.7 NRD=0 NRS=0 M=1
+ R=2.8 SA=75000.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1021 A_1578_533# N_A_757_317#_M1021_g N_A_1445_113#_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.208425 PD=0.86 PS=1.66 NRD=77.3816 NRS=206.948 M=1 R=2.8
+ SA=75000.3 SB=75002 A=0.063 P=1.14 MULT=1
MM1031 N_VPWR_M1031_d N_A_1641_21#_M1031_g A_1578_533# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.14385 AS=0.0924 PD=1.105 PS=0.86 NRD=0 NRS=77.3816 M=1 R=2.8 SA=75000.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1022 N_A_1641_21#_M1022_d N_RESET_B_M1022_g N_VPWR_M1031_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.14385 PD=0.7 PS=1.105 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_1445_113#_M1014_g N_A_1641_21#_M1022_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_865_255#_M1032_g N_A_757_317#_M1032_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.2394 AS=0.1113 PD=1.74 PS=1.37 NRD=241.542 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_865_255#_M1007_d N_CLK_M1007_g N_VPWR_M1032_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.2394 PD=1.37 PS=1.74 NRD=0 NRS=53.9386 M=1 R=2.8
+ SA=75000.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_1445_113#_M1003_g N_A_2408_367#_M1003_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.14912 AS=0.1696 PD=1.14189 PS=1.81 NRD=24.625 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1023 N_Q_M1023_d N_A_2408_367#_M1023_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.29358 PD=3.05 PS=2.24811 NRD=0 NRS=8.077 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.7743 P=31.37
c_145 VNB 0 8.87678e-20 $X=0 $Y=0
c_269 VPB 0 4.76477e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfrtp_ov2.pxi.spice"
*
.ends
*
*
