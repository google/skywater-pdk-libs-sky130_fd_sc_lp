* File: sky130_fd_sc_lp__and3_0.pex.spice
* Created: Wed Sep  2 09:31:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3_0%A 2 7 10 11 12 13 14 15 16 21 23
r42 21 23 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.02
+ $X2=0.605 $Y2=0.855
r43 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.02 $X2=0.59 $Y2=1.02
r44 15 16 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.677 $Y=1.295
+ $X2=0.677 $Y2=1.665
r45 15 22 8.68279 $w=3.63e-07 $l=2.75e-07 $layer=LI1_cond $X=0.677 $Y=1.295
+ $X2=0.677 $Y2=1.02
r46 14 22 2.99951 $w=3.63e-07 $l=9.5e-08 $layer=LI1_cond $X=0.677 $Y=0.925
+ $X2=0.677 $Y2=1.02
r47 12 13 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.697 $Y=2.155
+ $X2=0.697 $Y2=2.305
r48 11 12 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.695 $Y=1.525
+ $X2=0.695 $Y2=2.155
r49 10 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.715 $Y=2.625
+ $X2=0.715 $Y2=2.305
r50 7 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.71 $Y=0.535
+ $X2=0.71 $Y2=0.855
r51 2 11 43.2685 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.605 $Y=1.345
+ $X2=0.605 $Y2=1.525
r52 1 21 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=0.605 $Y=1.035
+ $X2=0.605 $Y2=1.02
r53 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=0.605 $Y=1.035
+ $X2=0.605 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_0%B 3 7 11 12 13 14 18
c49 7 0 1.10891e-19 $X=1.145 $Y=2.625
c50 3 0 1.7829e-19 $X=1.07 $Y=0.535
r51 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.41 $X2=1.16 $Y2=1.41
r52 14 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.195 $Y=1.665
+ $X2=1.195 $Y2=1.41
r53 13 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.41
r54 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.75
+ $X2=1.16 $Y2=1.41
r55 11 12 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.75
+ $X2=1.16 $Y2=1.915
r56 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.245
+ $X2=1.16 $Y2=1.41
r57 7 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.145 $Y=2.625
+ $X2=1.145 $Y2=1.915
r58 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.07 $Y=0.535
+ $X2=1.07 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_0%C 1 3 6 8 11 18 19 20 21 22 23 29 31 38
c62 31 0 3.91566e-20 $X=1.715 $Y=1.21
c63 21 0 1.7829e-19 $X=1.68 $Y=1.295
r64 32 38 2.46275 $w=3.63e-07 $l=7.8e-08 $layer=LI1_cond $X=1.712 $Y=1.743
+ $X2=1.712 $Y2=1.665
r65 29 31 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.375
+ $X2=1.715 $Y2=1.21
r66 22 23 10.6199 $w=3.32e-07 $l=2.89e-07 $layer=LI1_cond $X=1.712 $Y=1.746
+ $X2=1.712 $Y2=2.035
r67 22 32 0.224154 $w=3.65e-07 $l=3e-09 $layer=LI1_cond $X=1.712 $Y=1.746
+ $X2=1.712 $Y2=1.743
r68 22 38 0.126295 $w=3.63e-07 $l=4e-09 $layer=LI1_cond $X=1.712 $Y=1.661
+ $X2=1.712 $Y2=1.665
r69 21 22 11.556 $w=3.63e-07 $l=3.66e-07 $layer=LI1_cond $X=1.712 $Y=1.295
+ $X2=1.712 $Y2=1.661
r70 21 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.375 $X2=1.73 $Y2=1.375
r71 18 19 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=1.592 $Y=2.125
+ $X2=1.592 $Y2=2.275
r72 18 20 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.61 $Y=2.125
+ $X2=1.61 $Y2=1.88
r73 11 20 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.715 $Y=1.7
+ $X2=1.715 $Y2=1.88
r74 10 29 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.715 $Y=1.39
+ $X2=1.715 $Y2=1.375
r75 10 11 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.715 $Y=1.39
+ $X2=1.715 $Y2=1.7
r76 8 14 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.625 $Y=0.93
+ $X2=1.43 $Y2=0.93
r77 8 31 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.005
+ $X2=1.625 $Y2=1.21
r78 6 19 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.575 $Y=2.625
+ $X2=1.575 $Y2=2.275
r79 1 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.43 $Y=0.855
+ $X2=1.43 $Y2=0.93
r80 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.43 $Y=0.855 $X2=1.43
+ $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_0%A_68_65# 1 2 3 11 14 18 20 22 25 27 28 31 34
+ 37 38 41 42 44 46 47
c100 41 0 3.91566e-20 $X=2.27 $Y=1.12
c101 25 0 1.10891e-19 $X=0.5 $Y=2.625
r102 46 47 8.17035 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.625
+ $X2=1.355 $Y2=2.46
r103 42 50 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.292 $Y=1.12
+ $X2=2.292 $Y2=0.955
r104 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27
+ $Y=1.12 $X2=2.27 $Y2=1.12
r105 39 41 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=2.23 $Y=1 $X2=2.23
+ $Y2=1.12
r106 37 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.105 $Y=0.915
+ $X2=2.23 $Y2=1
r107 37 38 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.105 $Y=0.915
+ $X2=1.26 $Y2=0.915
r108 35 47 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.32 $Y=2.265
+ $X2=1.32 $Y2=2.46
r109 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.175 $Y=0.83
+ $X2=1.26 $Y2=0.915
r110 33 34 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.175 $Y=0.67
+ $X2=1.175 $Y2=0.83
r111 32 44 3.69268 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.625 $Y=2.18
+ $X2=0.39 $Y2=2.18
r112 31 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.225 $Y=2.18
+ $X2=1.32 $Y2=2.265
r113 31 32 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.225 $Y=2.18
+ $X2=0.625 $Y2=2.18
r114 28 30 5.37807 $w=2.98e-07 $l=1.4e-07 $layer=LI1_cond $X=0.325 $Y=0.52
+ $X2=0.465 $Y2=0.52
r115 27 33 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.09 $Y=0.52
+ $X2=1.175 $Y2=0.67
r116 27 30 24.0092 $w=2.98e-07 $l=6.25e-07 $layer=LI1_cond $X=1.09 $Y=0.52
+ $X2=0.465 $Y2=0.52
r117 23 44 2.96976 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.39 $Y=2.265
+ $X2=0.39 $Y2=2.18
r118 23 25 9.16145 $w=4.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.39 $Y=2.265
+ $X2=0.39 $Y2=2.625
r119 22 44 2.96976 $w=3.2e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.24 $Y=2.095
+ $X2=0.39 $Y2=2.18
r120 21 28 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.24 $Y=0.67
+ $X2=0.325 $Y2=0.52
r121 21 22 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=0.24 $Y=0.67
+ $X2=0.24 $Y2=2.095
r122 18 50 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.405 $Y=0.535
+ $X2=2.405 $Y2=0.955
r123 14 20 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=2.345 $Y=2.735
+ $X2=2.345 $Y2=1.625
r124 11 20 41.3024 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=2.292 $Y=1.438
+ $X2=2.292 $Y2=1.625
r125 10 42 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=2.292 $Y=1.142
+ $X2=2.292 $Y2=1.12
r126 10 11 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=2.292 $Y=1.142
+ $X2=2.292 $Y2=1.438
r127 3 46 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.415 $X2=1.36 $Y2=2.625
r128 2 25 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.375
+ $Y=2.415 $X2=0.5 $Y2=2.625
r129 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.325 $X2=0.465 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_0%VPWR 1 2 9 11 15 18 19 20 28 29 32
r33 33 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 32 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 29 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 26 32 12.6176 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=1.957 $Y2=3.33
r39 26 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 20 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 20 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 18 23 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 18 19 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.925 $Y2=3.33
r45 13 32 2.53987 $w=6.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.957 $Y=3.245
+ $X2=1.957 $Y2=3.33
r46 13 15 13.5424 $w=6.03e-07 $l=6.85e-07 $layer=LI1_cond $X=1.957 $Y=3.245
+ $X2=1.957 $Y2=2.56
r47 12 19 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.925 $Y2=3.33
r48 11 32 12.6176 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=1.655 $Y=3.33
+ $X2=1.957 $Y2=3.33
r49 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.655 $Y=3.33
+ $X2=1.055 $Y2=3.33
r50 7 19 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=3.33
r51 7 9 27.4813 $w=2.58e-07 $l=6.2e-07 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=2.625
r52 2 15 400 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=2.415 $X2=2.13 $Y2=2.56
r53 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=2.415 $X2=1.79 $Y2=2.56
r54 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.79
+ $Y=2.415 $X2=0.93 $Y2=2.625
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_0%X 1 2 7 8 9 10 11 12 13 41
r16 41 42 1.12001 $w=3.63e-07 $l=1e-08 $layer=LI1_cond $X=2.612 $Y=2.405
+ $X2=2.612 $Y2=2.395
r17 36 45 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=2.612 $Y=2.577
+ $X2=2.612 $Y2=2.56
r18 13 36 6.25161 $w=3.63e-07 $l=1.98e-07 $layer=LI1_cond $X=2.612 $Y=2.775
+ $X2=2.612 $Y2=2.577
r19 12 45 3.72571 $w=3.63e-07 $l=1.18e-07 $layer=LI1_cond $X=2.612 $Y=2.442
+ $X2=2.612 $Y2=2.56
r20 12 41 1.16823 $w=3.63e-07 $l=3.7e-08 $layer=LI1_cond $X=2.612 $Y=2.442
+ $X2=2.612 $Y2=2.405
r21 12 42 1.62196 $w=2.68e-07 $l=3.8e-08 $layer=LI1_cond $X=2.66 $Y=2.357
+ $X2=2.66 $Y2=2.395
r22 11 12 13.7439 $w=2.68e-07 $l=3.22e-07 $layer=LI1_cond $X=2.66 $Y=2.035
+ $X2=2.66 $Y2=2.357
r23 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=1.665
+ $X2=2.66 $Y2=2.035
r24 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=1.295
+ $X2=2.66 $Y2=1.665
r25 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=0.925 $X2=2.66
+ $Y2=1.295
r26 7 8 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.66 $Y=0.535 $X2=2.66
+ $Y2=0.925
r27 2 45 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.42
+ $Y=2.415 $X2=2.56 $Y2=2.56
r28 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.325 $X2=2.62 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_0%VGND 1 4 16 17 22 28
r26 27 28 11.0915 $w=7.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0.287
+ $X2=2.355 $Y2=0.287
r27 24 27 0.481642 $w=7.43e-07 $l=3e-08 $layer=LI1_cond $X=2.16 $Y=0.287
+ $X2=2.19 $Y2=0.287
r28 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r29 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r30 20 24 7.70628 $w=7.43e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.287
+ $X2=2.16 $Y2=0.287
r31 20 22 11.6534 $w=7.43e-07 $l=2e-07 $layer=LI1_cond $X=1.68 $Y=0.287 $X2=1.48
+ $Y2=0.287
r32 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r33 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r34 16 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.355
+ $Y2=0
r35 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r36 12 22 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.48
+ $Y2=0
r37 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 9 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r39 8 12 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r40 8 9 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 4 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r42 4 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r43 1 27 91 $w=1.7e-07 $l=7.82991e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.325 $X2=2.19 $Y2=0.535
.ends

