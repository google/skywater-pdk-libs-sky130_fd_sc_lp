* File: sky130_fd_sc_lp__dfrbp_2.pex.spice
* Created: Wed Sep  2 09:43:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFRBP_2%CLK 3 5 7 9 10
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=1.805 $X2=0.635 $Y2=1.805
r36 10 15 6.97531 $w=3.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.715 $Y=2.035
+ $X2=0.715 $Y2=1.805
r37 9 15 4.24584 $w=3.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.715 $Y=1.665
+ $X2=0.715 $Y2=1.805
r38 5 14 38.7751 $w=2.77e-07 $l=2.09105e-07 $layer=POLY_cond $X=0.5 $Y=1.97
+ $X2=0.6 $Y2=1.805
r39 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.5 $Y=1.97 $X2=0.5
+ $Y2=2.68
r40 1 14 89.2372 $w=2.77e-07 $l=5.13712e-07 $layer=POLY_cond $X=0.475 $Y=1.35
+ $X2=0.6 $Y2=1.805
r41 1 3 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.475 $Y=1.35
+ $X2=0.475 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%D 3 6 9 10 11 12 13 17
c51 12 0 9.92892e-20 $X=2.16 $Y=1.295
r52 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.51
+ $Y=1.65 $X2=2.51 $Y2=1.65
r53 13 18 0.309331 $w=5.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.35 $Y=1.665
+ $X2=2.35 $Y2=1.65
r54 12 18 7.32082 $w=5.78e-07 $l=3.55e-07 $layer=LI1_cond $X=2.35 $Y=1.295
+ $X2=2.35 $Y2=1.65
r55 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.51 $Y=1.99
+ $X2=2.51 $Y2=1.65
r56 10 11 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.99
+ $X2=2.51 $Y2=2.155
r57 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.485
+ $X2=2.51 $Y2=1.65
r58 6 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.45 $Y=2.525
+ $X2=2.45 $Y2=2.155
r59 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.42 $Y=1.165 $X2=2.42
+ $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_196_79# 1 2 9 11 13 14 16 17 21 25 28 29
+ 31 33 36 37 39 43 49 50 51 55 59 60 72
c187 60 0 1.05865e-20 $X=3.54 $Y=1.78
c188 59 0 5.60296e-20 $X=3.54 $Y=1.78
r189 60 66 12.479 $w=3.09e-07 $l=8e-08 $layer=POLY_cond $X=3.54 $Y=1.697
+ $X2=3.46 $Y2=1.697
r190 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.54
+ $Y=1.78 $X2=3.54 $Y2=1.78
r191 56 59 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.29 $Y=1.78
+ $X2=3.54 $Y2=1.78
r192 51 53 11.5244 $w=2.38e-07 $l=2.4e-07 $layer=LI1_cond $X=2.195 $Y=0.715
+ $X2=2.195 $Y2=0.955
r193 49 50 13.6023 $w=1.78e-07 $l=2.2e-07 $layer=LI1_cond $X=1.312 $Y=1.935
+ $X2=1.312 $Y2=2.155
r194 44 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.385 $Y=1.555
+ $X2=6.55 $Y2=1.555
r195 44 69 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.385 $Y=1.555
+ $X2=6.285 $Y2=1.555
r196 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.385
+ $Y=1.555 $X2=6.385 $Y2=1.555
r197 41 43 40.9747 $w=1.78e-07 $l=6.65e-07 $layer=LI1_cond $X=6.38 $Y=0.89
+ $X2=6.38 $Y2=1.555
r198 40 64 2.11506 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=4.775 $Y=0.805
+ $X2=4.667 $Y2=0.805
r199 39 41 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.29 $Y=0.805
+ $X2=6.38 $Y2=0.89
r200 39 40 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=6.29 $Y=0.805
+ $X2=4.775 $Y2=0.805
r201 38 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=0.715
+ $X2=3.29 $Y2=0.715
r202 37 64 4.82418 $w=2.13e-07 $l=9e-08 $layer=LI1_cond $X=4.667 $Y=0.715
+ $X2=4.667 $Y2=0.805
r203 37 38 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=4.56 $Y=0.715
+ $X2=3.375 $Y2=0.715
r204 36 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=1.615
+ $X2=3.29 $Y2=1.78
r205 35 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.8 $X2=3.29
+ $Y2=0.715
r206 35 36 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.29 $Y=0.8
+ $X2=3.29 $Y2=1.615
r207 34 51 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.315 $Y=0.715
+ $X2=2.195 $Y2=0.715
r208 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=0.715
+ $X2=3.29 $Y2=0.715
r209 33 34 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.205 $Y=0.715
+ $X2=2.315 $Y2=0.715
r210 32 47 14.6964 $w=3.03e-07 $l=4.57324e-07 $layer=LI1_cond $X=1.415 $Y=0.955
+ $X2=1.207 $Y2=0.59
r211 31 53 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.075 $Y=0.955
+ $X2=2.195 $Y2=0.955
r212 31 32 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.075 $Y=0.955
+ $X2=1.415 $Y2=0.955
r213 29 32 5.41666 $w=3.03e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.325 $Y=1.04
+ $X2=1.415 $Y2=0.955
r214 29 49 55.1465 $w=1.78e-07 $l=8.95e-07 $layer=LI1_cond $X=1.325 $Y=1.04
+ $X2=1.325 $Y2=1.935
r215 28 50 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.295 $Y=2.305
+ $X2=1.295 $Y2=2.155
r216 23 28 7.43437 $w=3.2e-07 $l=2.31571e-07 $layer=LI1_cond $X=1.215 $Y=2.5
+ $X2=1.295 $Y2=2.305
r217 23 25 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.215 $Y=2.5
+ $X2=1.215 $Y2=2.515
r218 19 21 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=6.935 $Y=1.72
+ $X2=6.935 $Y2=2.69
r219 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.86 $Y=1.645
+ $X2=6.935 $Y2=1.72
r220 17 72 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.86 $Y=1.645
+ $X2=6.55 $Y2=1.645
r221 14 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.285 $Y=1.39
+ $X2=6.285 $Y2=1.555
r222 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.285 $Y=1.39
+ $X2=6.285 $Y2=0.96
r223 11 60 47.5761 $w=3.09e-07 $l=4.10317e-07 $layer=POLY_cond $X=3.845 $Y=1.45
+ $X2=3.54 $Y2=1.697
r224 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.845 $Y=1.45
+ $X2=3.845 $Y2=1.165
r225 7 66 19.6649 $w=1.5e-07 $l=2.48e-07 $layer=POLY_cond $X=3.46 $Y=1.945
+ $X2=3.46 $Y2=1.697
r226 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.46 $Y=1.945
+ $X2=3.46 $Y2=2.525
r227 2 25 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.005
+ $Y=2.36 $X2=1.145 $Y2=2.515
r228 1 47 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.395 $X2=1.12 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_811_341# 1 2 9 11 13 17 20 21 23 24 25 27
+ 30 33 37
c112 17 0 1.05865e-20 $X=4.22 $Y=1.82
r113 33 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.955 $Y=1.155
+ $X2=5.955 $Y2=1.32
r114 28 37 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=6.057 $Y=2.07
+ $X2=6.057 $Y2=1.985
r115 28 30 36.1814 $w=2.13e-07 $l=6.75e-07 $layer=LI1_cond $X=6.057 $Y=2.07
+ $X2=6.057 $Y2=2.745
r116 27 37 4.65272 $w=1.92e-07 $l=9.53677e-08 $layer=LI1_cond $X=6.035 $Y=1.9
+ $X2=6.057 $Y2=1.985
r117 27 35 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.035 $Y=1.9
+ $X2=6.035 $Y2=1.32
r118 24 37 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.95 $Y=1.985
+ $X2=6.057 $Y2=1.985
r119 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.95 $Y=1.985
+ $X2=5.26 $Y2=1.985
r120 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.175 $Y=1.9
+ $X2=5.26 $Y2=1.985
r121 22 23 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.175 $Y=1.61
+ $X2=5.175 $Y2=1.9
r122 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.09 $Y=1.525
+ $X2=5.175 $Y2=1.61
r123 20 21 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=5.09 $Y=1.525
+ $X2=4.305 $Y2=1.525
r124 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=1.82 $X2=4.22 $Y2=1.82
r125 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.22 $Y=1.61
+ $X2=4.305 $Y2=1.525
r126 15 17 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.22 $Y=1.61
+ $X2=4.22 $Y2=1.82
r127 11 18 38.5818 $w=3.27e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.25 $Y=1.985
+ $X2=4.22 $Y2=1.82
r128 11 13 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.25 $Y=1.985
+ $X2=4.25 $Y2=2.525
r129 7 18 38.5818 $w=3.27e-07 $l=1.69926e-07 $layer=POLY_cond $X=4.23 $Y=1.655
+ $X2=4.22 $Y2=1.82
r130 7 9 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=4.23 $Y=1.655
+ $X2=4.23 $Y2=1.165
r131 2 37 400 $w=1.7e-07 $l=3.08504e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.895 $X2=6.06 $Y2=2.065
r132 2 30 400 $w=1.7e-07 $l=9.60339e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.895 $X2=6.06 $Y2=2.745
r133 1 33 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.64 $X2=5.955 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%RESET_B 3 8 9 10 14 19 23 27 32 35 37 38 39
+ 40 41 48 49 52 53 55 57 64 71
c194 71 0 5.49373e-20 $X=7.92 $Y=2.035
c195 57 0 2.01996e-20 $X=4.807 $Y=1.79
c196 49 0 1.63892e-19 $X=7.92 $Y=2.035
c197 38 0 2.9381e-20 $X=4.415 $Y=2.035
c198 37 0 1.00911e-19 $X=4.677 $Y=1.56
c199 9 0 9.92892e-20 $X=4.58 $Y=0.54
r200 62 64 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=7.925 $Y=2.115
+ $X2=8.11 $Y2=2.115
r201 62 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.925
+ $Y=2.115 $X2=7.925 $Y2=2.115
r202 59 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.835 $Y=2.115
+ $X2=7.925 $Y2=2.115
r203 55 58 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.807 $Y=1.955
+ $X2=4.807 $Y2=2.12
r204 55 57 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.807 $Y=1.955
+ $X2=4.807 $Y2=1.79
r205 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.825
+ $Y=1.955 $X2=4.825 $Y2=1.955
r206 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.795
+ $Y=1.65 $X2=1.795 $Y2=1.65
r207 49 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r208 48 56 10.0404 $w=3.22e-07 $l=2.65e-07 $layer=LI1_cond $X=4.56 $Y=1.955
+ $X2=4.825 $Y2=1.955
r209 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.035
+ $X2=4.56 $Y2=2.035
r210 44 53 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=1.737 $Y=2.035
+ $X2=1.737 $Y2=1.65
r211 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.035
r212 41 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.035
+ $X2=4.56 $Y2=2.035
r213 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r214 40 41 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.705 $Y2=2.035
r215 39 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=2.035
+ $X2=1.68 $Y2=2.035
r216 38 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=4.56 $Y2=2.035
r217 38 39 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=1.825 $Y2=2.035
r218 37 57 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.7 $Y=1.56 $X2=4.7
+ $Y2=1.79
r219 36 37 37.4087 $w=1.95e-07 $l=1.1e-07 $layer=POLY_cond $X=4.677 $Y=1.45
+ $X2=4.677 $Y2=1.56
r220 34 52 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.795 $Y=1.99
+ $X2=1.795 $Y2=1.65
r221 34 35 45.2978 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.99
+ $X2=1.795 $Y2=2.155
r222 30 52 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.795 $Y=1.635
+ $X2=1.795 $Y2=1.65
r223 30 32 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.795 $Y=1.56
+ $X2=2.06 $Y2=1.56
r224 25 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.11 $Y=2.28
+ $X2=8.11 $Y2=2.115
r225 25 27 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.11 $Y=2.28
+ $X2=8.11 $Y2=2.69
r226 21 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.835 $Y=1.95
+ $X2=7.835 $Y2=2.115
r227 21 23 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=7.835 $Y=1.95
+ $X2=7.835 $Y2=0.85
r228 19 58 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.8 $Y=2.525
+ $X2=4.8 $Y2=2.12
r229 14 36 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.655 $Y=1.165
+ $X2=4.655 $Y2=1.45
r230 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.655 $Y=0.615
+ $X2=4.655 $Y2=1.165
r231 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.58 $Y=0.54
+ $X2=4.655 $Y2=0.615
r232 9 10 1253.71 $w=1.5e-07 $l=2.445e-06 $layer=POLY_cond $X=4.58 $Y=0.54
+ $X2=2.135 $Y2=0.54
r233 6 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=1.485
+ $X2=2.06 $Y2=1.56
r234 6 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.06 $Y=1.485
+ $X2=2.06 $Y2=1.165
r235 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.06 $Y=0.615
+ $X2=2.135 $Y2=0.54
r236 5 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.06 $Y=0.615
+ $X2=2.06 $Y2=1.165
r237 3 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.88 $Y=2.525
+ $X2=1.88 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_637_191# 1 2 3 10 12 15 18 19 20 21 22 25
+ 42
c104 25 0 1.2111e-19 $X=5.525 $Y=1.555
c105 20 0 1.60894e-19 $X=3.985 $Y=2.385
r106 41 42 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.74 $Y=1.555
+ $X2=5.75 $Y2=1.555
r107 32 33 9.71338 $w=3.14e-07 $l=2.5e-07 $layer=LI1_cond $X=3.63 $Y=1.135
+ $X2=3.88 $Y2=1.135
r108 29 30 6.34772 $w=3.94e-07 $l=2.05e-07 $layer=LI1_cond $X=3.675 $Y=2.517
+ $X2=3.88 $Y2=2.517
r109 26 41 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.525 $Y=1.555
+ $X2=5.74 $Y2=1.555
r110 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.525
+ $Y=1.555 $X2=5.525 $Y2=1.555
r111 23 25 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=5.525 $Y=1.26
+ $X2=5.525 $Y2=1.555
r112 22 33 15.3951 $w=3.14e-07 $l=3.67287e-07 $layer=LI1_cond $X=4.235 $Y=1.16
+ $X2=3.88 $Y2=1.135
r113 21 23 6.82232 $w=2e-07 $l=1.39642e-07 $layer=LI1_cond $X=5.43 $Y=1.16
+ $X2=5.525 $Y2=1.26
r114 21 22 66.2682 $w=1.98e-07 $l=1.195e-06 $layer=LI1_cond $X=5.43 $Y=1.16
+ $X2=4.235 $Y2=1.16
r115 20 30 7.27085 $w=3.94e-07 $l=1.76873e-07 $layer=LI1_cond $X=3.985 $Y=2.385
+ $X2=3.88 $Y2=2.517
r116 19 37 6.82058 $w=2.43e-07 $l=1.45e-07 $layer=LI1_cond $X=4.992 $Y=2.385
+ $X2=4.992 $Y2=2.53
r117 19 20 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.87 $Y=2.385
+ $X2=3.985 $Y2=2.385
r118 18 30 5.68665 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.88 $Y=2.3
+ $X2=3.88 $Y2=2.517
r119 17 33 4.32966 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=1.3
+ $X2=3.88 $Y2=1.135
r120 17 18 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.88 $Y=1.3 $X2=3.88
+ $Y2=2.3
r121 13 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.75 $Y=1.72
+ $X2=5.75 $Y2=1.555
r122 13 15 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.75 $Y=1.72
+ $X2=5.75 $Y2=2.315
r123 10 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=1.39
+ $X2=5.74 $Y2=1.555
r124 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.74 $Y=1.39
+ $X2=5.74 $Y2=0.96
r125 3 37 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=4.875
+ $Y=2.315 $X2=5.015 $Y2=2.53
r126 2 29 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=3.535
+ $Y=2.315 $X2=3.675 $Y2=2.535
r127 1 32 182 $w=1.7e-07 $l=5.27376e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.955 $X2=3.63 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_27_79# 1 2 10 14 15 16 17 18 20 22 24 25
+ 27 28 32 34 38 42 44 48 50 51 54 58 60 64 65 67 68
c164 32 0 2.9381e-20 $X=3.89 $Y=2.525
c165 25 0 1.57615e-19 $X=3.11 $Y=1.45
c166 22 0 2.16924e-19 $X=2.96 $Y=3.075
r167 65 71 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.972 $Y=1.09
+ $X2=0.972 $Y2=1.255
r168 65 70 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.972 $Y=1.09
+ $X2=0.972 $Y2=0.925
r169 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.09 $X2=0.95 $Y2=1.09
r170 62 67 0.466467 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=0.4 $Y=1.09
+ $X2=0.26 $Y2=1.09
r171 62 64 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.4 $Y=1.09
+ $X2=0.95 $Y2=1.09
r172 58 68 5.89299 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.25 $Y=2.465
+ $X2=0.25 $Y2=2.335
r173 58 60 2.21624 $w=2.58e-07 $l=5e-08 $layer=LI1_cond $X=0.25 $Y=2.465
+ $X2=0.25 $Y2=2.515
r174 56 67 6.31733 $w=2.57e-07 $l=1.76125e-07 $layer=LI1_cond $X=0.237 $Y=1.255
+ $X2=0.26 $Y2=1.09
r175 56 68 52.9633 $w=2.33e-07 $l=1.08e-06 $layer=LI1_cond $X=0.237 $Y=1.255
+ $X2=0.237 $Y2=2.335
r176 52 67 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=0.925
+ $X2=0.26 $Y2=1.09
r177 52 54 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.925
+ $X2=0.26 $Y2=0.59
r178 46 48 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=2.96 $Y=1.86
+ $X2=3.09 $Y2=1.86
r179 44 45 49.1513 $w=1.52e-07 $l=1.55e-07 $layer=POLY_cond $X=0.93 $Y=2.202
+ $X2=1.085 $Y2=2.202
r180 40 42 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=7.045 $Y=0.255
+ $X2=7.045 $Y2=0.85
r181 36 38 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=6.41 $Y=3.075
+ $X2=6.41 $Y2=2.48
r182 35 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.965 $Y=3.15
+ $X2=3.89 $Y2=3.15
r183 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.335 $Y=3.15
+ $X2=6.41 $Y2=3.075
r184 34 35 1215.26 $w=1.5e-07 $l=2.37e-06 $layer=POLY_cond $X=6.335 $Y=3.15
+ $X2=3.965 $Y2=3.15
r185 30 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.89 $Y=3.075
+ $X2=3.89 $Y2=3.15
r186 30 32 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.89 $Y=3.075
+ $X2=3.89 $Y2=2.525
r187 29 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.035 $Y=3.15
+ $X2=2.96 $Y2=3.15
r188 28 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.89 $Y2=3.15
r189 28 29 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.035 $Y2=3.15
r190 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.11 $Y=1.45
+ $X2=3.11 $Y2=1.165
r191 24 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.09 $Y=1.785
+ $X2=3.09 $Y2=1.86
r192 23 25 28.8623 $w=1.67e-07 $l=1.09545e-07 $layer=POLY_cond $X=3.09 $Y=1.55
+ $X2=3.11 $Y2=1.45
r193 23 24 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.09 $Y=1.55
+ $X2=3.09 $Y2=1.785
r194 22 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.96 $Y=3.075
+ $X2=2.96 $Y2=3.15
r195 21 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.96 $Y=1.935
+ $X2=2.96 $Y2=1.86
r196 21 22 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.96 $Y=1.935
+ $X2=2.96 $Y2=3.075
r197 20 45 3.14937 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=1.085 $Y=2.12
+ $X2=1.085 $Y2=2.202
r198 20 71 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=1.085 $Y=2.12
+ $X2=1.085 $Y2=1.255
r199 17 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=3.15
+ $X2=2.96 $Y2=3.15
r200 17 18 964 $w=1.5e-07 $l=1.88e-06 $layer=POLY_cond $X=2.885 $Y=3.15
+ $X2=1.005 $Y2=3.15
r201 15 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.97 $Y=0.18
+ $X2=7.045 $Y2=0.255
r202 15 16 3071.47 $w=1.5e-07 $l=5.99e-06 $layer=POLY_cond $X=6.97 $Y=0.18
+ $X2=0.98 $Y2=0.18
r203 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=3.075
+ $X2=1.005 $Y2=3.15
r204 12 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.93 $Y=3.075
+ $X2=0.93 $Y2=2.68
r205 11 44 3.14937 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=0.93 $Y=2.285
+ $X2=0.93 $Y2=2.202
r206 11 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.93 $Y=2.285
+ $X2=0.93 $Y2=2.68
r207 10 70 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=0.605
+ $X2=0.905 $Y2=0.925
r208 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=0.255
+ $X2=0.98 $Y2=0.18
r209 7 10 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.905 $Y=0.255
+ $X2=0.905 $Y2=0.605
r210 2 60 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.36 $X2=0.285 $Y2=2.515
r211 1 54 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.395 $X2=0.26 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_1444_320# 1 2 9 13 17 18 21 25 27 31 34 36
+ 37 38
c90 38 0 4.6324e-20 $X=8.355 $Y=1.69
c91 37 0 1.20202e-19 $X=7.385 $Y=1.765
c92 34 0 7.47908e-20 $X=8.885 $Y=1.6
c93 31 0 6.70338e-20 $X=8.745 $Y=1.685
c94 17 0 1.63892e-19 $X=7.385 $Y=2.105
c95 9 0 5.49373e-20 $X=7.295 $Y=2.69
r96 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.385
+ $Y=1.765 $X2=7.385 $Y2=1.765
r97 33 34 21.8141 $w=2.78e-07 $l=5.3e-07 $layer=LI1_cond $X=8.885 $Y=1.07
+ $X2=8.885 $Y2=1.6
r98 32 38 7.28786 $w=1.75e-07 $l=1.37477e-07 $layer=LI1_cond $X=8.49 $Y=1.685
+ $X2=8.355 $Y2=1.69
r99 31 34 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=8.745 $Y=1.685
+ $X2=8.885 $Y2=1.6
r100 31 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.745 $Y=1.685
+ $X2=8.49 $Y2=1.685
r101 27 33 6.84494 $w=2.5e-07 $l=1.92614e-07 $layer=LI1_cond $X=8.745 $Y=0.945
+ $X2=8.885 $Y2=1.07
r102 27 29 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.745 $Y=0.945
+ $X2=8.41 $Y2=0.945
r103 23 38 0.161356 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=8.355 $Y=1.78
+ $X2=8.355 $Y2=1.69
r104 23 25 38.8416 $w=2.68e-07 $l=9.1e-07 $layer=LI1_cond $X=8.355 $Y=1.78
+ $X2=8.355 $Y2=2.69
r105 22 36 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.55 $Y=1.69
+ $X2=7.385 $Y2=1.69
r106 21 38 7.28786 $w=1.75e-07 $l=1.35e-07 $layer=LI1_cond $X=8.22 $Y=1.69
+ $X2=8.355 $Y2=1.69
r107 21 22 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=8.22 $Y=1.69
+ $X2=7.55 $Y2=1.69
r108 17 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.385 $Y=2.105
+ $X2=7.385 $Y2=1.765
r109 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.385 $Y=2.105
+ $X2=7.385 $Y2=2.27
r110 16 37 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.385 $Y=1.6
+ $X2=7.385 $Y2=1.765
r111 13 16 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=7.405 $Y=0.85
+ $X2=7.405 $Y2=1.6
r112 9 18 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=7.295 $Y=2.69
+ $X2=7.295 $Y2=2.27
r113 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=2.48 $X2=8.325 $Y2=2.69
r114 1 29 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.64 $X2=8.41 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_1272_128# 1 2 7 9 12 14 15 18 22 24 28 32
+ 34 37 40 44 46 47 50 52 53 55 61 67 70 71
c164 70 0 1.20202e-19 $X=6.68 $Y=2.04
c165 52 0 5.41964e-20 $X=10.465 $Y=1.425
c166 28 0 1.41825e-19 $X=9.495 $Y=2.27
c167 18 0 4.6324e-20 $X=9.065 $Y=2.27
r168 68 74 23.4306 $w=2.88e-07 $l=1.4e-07 $layer=POLY_cond $X=8.4 $Y=1.335
+ $X2=8.54 $Y2=1.335
r169 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.4
+ $Y=1.335 $X2=8.4 $Y2=1.335
r170 65 71 1.5279 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=6.84 $Y=1.335 $X2=6.74
+ $Y2=1.335
r171 65 67 91.0622 $w=1.88e-07 $l=1.56e-06 $layer=LI1_cond $X=6.84 $Y=1.335
+ $X2=8.4 $Y2=1.335
r172 63 71 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=6.74 $Y=1.43 $X2=6.74
+ $Y2=1.335
r173 63 70 33.8273 $w=1.98e-07 $l=6.1e-07 $layer=LI1_cond $X=6.74 $Y=1.43
+ $X2=6.74 $Y2=2.04
r174 59 71 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=6.74 $Y=1.24 $X2=6.74
+ $Y2=1.335
r175 59 61 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.74 $Y=1.24
+ $X2=6.74 $Y2=0.905
r176 55 57 19.4475 $w=3.18e-07 $l=5.4e-07 $layer=LI1_cond $X=6.68 $Y=2.205
+ $X2=6.68 $Y2=2.745
r177 53 70 7.37399 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=6.68 $Y=2.2
+ $X2=6.68 $Y2=2.04
r178 53 55 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=6.68 $Y=2.2 $X2=6.68
+ $Y2=2.205
r179 48 50 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.45 $Y=0.98
+ $X2=10.54 $Y2=0.98
r180 42 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.54 $Y=0.905
+ $X2=10.54 $Y2=0.98
r181 42 44 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=10.54 $Y=0.905
+ $X2=10.54 $Y2=0.555
r182 38 52 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=10.48 $Y=1.5
+ $X2=10.465 $Y2=1.425
r183 38 40 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=10.48 $Y=1.5
+ $X2=10.48 $Y2=2.155
r184 37 52 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=10.45 $Y=1.35
+ $X2=10.465 $Y2=1.425
r185 36 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.45 $Y=1.055
+ $X2=10.45 $Y2=0.98
r186 36 37 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=10.45 $Y=1.055
+ $X2=10.45 $Y2=1.35
r187 35 47 12.05 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=9.65 $Y=1.425
+ $X2=9.535 $Y2=1.425
r188 34 52 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.375 $Y=1.425
+ $X2=10.465 $Y2=1.425
r189 34 35 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=10.375 $Y=1.425
+ $X2=9.65 $Y2=1.425
r190 30 47 12.05 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=9.575 $Y=1.35
+ $X2=9.535 $Y2=1.425
r191 30 32 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.575 $Y=1.35
+ $X2=9.575 $Y2=0.67
r192 26 47 12.05 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=9.495 $Y=1.5
+ $X2=9.535 $Y2=1.425
r193 26 28 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=9.495 $Y=1.5
+ $X2=9.495 $Y2=2.27
r194 25 46 12.05 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=9.22 $Y=1.425
+ $X2=9.105 $Y2=1.425
r195 24 47 12.05 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=9.42 $Y=1.425
+ $X2=9.535 $Y2=1.425
r196 24 25 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=9.42 $Y=1.425
+ $X2=9.22 $Y2=1.425
r197 20 46 12.05 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=9.145 $Y=1.35
+ $X2=9.105 $Y2=1.425
r198 20 22 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.145 $Y=1.35
+ $X2=9.145 $Y2=0.67
r199 16 46 12.05 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=9.065 $Y=1.5
+ $X2=9.105 $Y2=1.425
r200 16 18 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=9.065 $Y=1.5
+ $X2=9.065 $Y2=2.27
r201 15 74 23.5717 $w=2.88e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.615 $Y=1.425
+ $X2=8.54 $Y2=1.335
r202 14 46 12.05 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=8.99 $Y=1.425
+ $X2=9.105 $Y2=1.425
r203 14 15 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=8.99 $Y=1.425
+ $X2=8.615 $Y2=1.425
r204 10 74 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.54 $Y=1.5
+ $X2=8.54 $Y2=1.335
r205 10 12 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=8.54 $Y=1.5
+ $X2=8.54 $Y2=2.69
r206 7 68 34.309 $w=2.88e-07 $l=2.75409e-07 $layer=POLY_cond $X=8.195 $Y=1.17
+ $X2=8.4 $Y2=1.335
r207 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.195 $Y=1.17
+ $X2=8.195 $Y2=0.85
r208 2 57 600 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=1 $X=6.485
+ $Y=2.06 $X2=6.625 $Y2=2.745
r209 2 55 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.485
+ $Y=2.06 $X2=6.625 $Y2=2.205
r210 1 61 182 $w=1.7e-07 $l=4.89898e-07 $layer=licon1_NDIFF $count=1 $X=6.36
+ $Y=0.64 $X2=6.735 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_2028_367# 1 2 9 12 14 18 22 24 27 31 35 36
+ 38 40
r67 41 42 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=10.952 $Y=1.55
+ $X2=10.952 $Y2=1.625
r68 36 41 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=10.952 $Y=1.46
+ $X2=10.952 $Y2=1.55
r69 36 40 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=10.952 $Y=1.46
+ $X2=10.952 $Y2=1.295
r70 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.93
+ $Y=1.46 $X2=10.93 $Y2=1.46
r71 33 38 1.39677 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=10.49 $Y=1.46
+ $X2=10.307 $Y2=1.46
r72 33 35 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=10.49 $Y=1.46
+ $X2=10.93 $Y2=1.46
r73 29 38 5.10169 $w=3.35e-07 $l=1.79374e-07 $layer=LI1_cond $X=10.277 $Y=1.625
+ $X2=10.307 $Y2=1.46
r74 29 31 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=10.277 $Y=1.625
+ $X2=10.277 $Y2=1.98
r75 25 38 5.10169 $w=3.35e-07 $l=1.65e-07 $layer=LI1_cond $X=10.307 $Y=1.295
+ $X2=10.307 $Y2=1.46
r76 25 27 23.5225 $w=3.63e-07 $l=7.45e-07 $layer=LI1_cond $X=10.307 $Y=1.295
+ $X2=10.307 $Y2=0.55
r77 20 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.495 $Y=1.625
+ $X2=11.495 $Y2=1.55
r78 20 22 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=11.495 $Y=1.625
+ $X2=11.495 $Y2=2.465
r79 16 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.495 $Y=1.475
+ $X2=11.495 $Y2=1.55
r80 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=11.495 $Y=1.475
+ $X2=11.495 $Y2=0.765
r81 15 41 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=11.14 $Y=1.55
+ $X2=10.952 $Y2=1.55
r82 14 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.42 $Y=1.55
+ $X2=11.495 $Y2=1.55
r83 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=11.42 $Y=1.55
+ $X2=11.14 $Y2=1.55
r84 12 42 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=11.065 $Y=2.465
+ $X2=11.065 $Y2=1.625
r85 9 40 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.065 $Y=0.765
+ $X2=11.065 $Y2=1.295
r86 2 31 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.14
+ $Y=1.835 $X2=10.265 $Y2=1.98
r87 1 27 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=10.2
+ $Y=0.345 $X2=10.325 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 56
+ 62 66 68 73 74 75 77 82 87 95 100 108 117 121 127 130 133 136 139 142 145 149
r155 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r156 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r157 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r159 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r160 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r161 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r162 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r163 125 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r164 125 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r165 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r166 122 145 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=10.955 $Y=3.33
+ $X2=10.777 $Y2=3.33
r167 122 124 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.955 $Y=3.33
+ $X2=11.28 $Y2=3.33
r168 121 148 4.38626 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=11.58 $Y=3.33
+ $X2=11.79 $Y2=3.33
r169 121 124 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=11.58 $Y=3.33
+ $X2=11.28 $Y2=3.33
r170 120 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r171 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r172 117 145 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=10.6 $Y=3.33
+ $X2=10.777 $Y2=3.33
r173 117 119 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.6 $Y=3.33
+ $X2=10.32 $Y2=3.33
r174 116 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r175 116 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r176 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r177 113 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=3.33
+ $X2=8.85 $Y2=3.33
r178 113 115 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.015 $Y=3.33
+ $X2=9.36 $Y2=3.33
r179 112 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r180 112 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r181 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r182 109 139 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.685 $Y2=3.33
r183 109 111 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r184 108 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.85 $Y2=3.33
r185 108 111 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.4 $Y2=3.33
r186 107 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r187 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r188 103 106 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r189 101 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.535 $Y2=3.33
r190 101 103 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.7 $Y=3.33 $X2=6
+ $Y2=3.33
r191 100 139 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=7.345 $Y=3.33
+ $X2=7.685 $Y2=3.33
r192 100 106 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.345 $Y=3.33
+ $X2=6.96 $Y2=3.33
r193 99 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r194 99 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r195 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r196 96 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.69 $Y=3.33
+ $X2=4.525 $Y2=3.33
r197 96 98 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.69 $Y=3.33
+ $X2=5.04 $Y2=3.33
r198 95 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.535 $Y2=3.33
r199 95 98 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.04 $Y2=3.33
r200 94 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r201 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r202 91 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r203 91 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r204 90 93 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r205 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r206 88 130 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.165 $Y2=3.33
r207 88 90 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=3.33 $X2=2.64
+ $Y2=3.33
r208 87 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.36 $Y=3.33
+ $X2=4.525 $Y2=3.33
r209 87 93 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r210 86 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r211 86 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r212 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r213 83 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=3.33
+ $X2=0.715 $Y2=3.33
r214 83 85 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.88 $Y=3.33 $X2=1.68
+ $Y2=3.33
r215 82 130 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.99 $Y=3.33
+ $X2=2.165 $Y2=3.33
r216 82 85 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.99 $Y=3.33
+ $X2=1.68 $Y2=3.33
r217 80 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r218 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r219 77 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.715 $Y2=3.33
r220 77 79 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.24 $Y2=3.33
r221 75 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r222 75 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r223 75 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r224 73 115 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.625 $Y=3.33
+ $X2=9.36 $Y2=3.33
r225 73 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.625 $Y=3.33
+ $X2=9.75 $Y2=3.33
r226 72 119 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.875 $Y=3.33
+ $X2=10.32 $Y2=3.33
r227 72 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.875 $Y=3.33
+ $X2=9.75 $Y2=3.33
r228 68 71 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=11.727 $Y=1.98
+ $X2=11.727 $Y2=2.95
r229 66 148 3.09127 $w=2.95e-07 $l=1.12161e-07 $layer=LI1_cond $X=11.727
+ $Y=3.245 $X2=11.79 $Y2=3.33
r230 66 71 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=11.727 $Y=3.245
+ $X2=11.727 $Y2=2.95
r231 62 65 15.907 $w=3.53e-07 $l=4.9e-07 $layer=LI1_cond $X=10.777 $Y=1.98
+ $X2=10.777 $Y2=2.47
r232 60 145 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=10.777 $Y=3.245
+ $X2=10.777 $Y2=3.33
r233 60 65 25.159 $w=3.53e-07 $l=7.75e-07 $layer=LI1_cond $X=10.777 $Y=3.245
+ $X2=10.777 $Y2=2.47
r234 56 59 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=9.75 $Y=1.785
+ $X2=9.75 $Y2=2.755
r235 54 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.75 $Y=3.245
+ $X2=9.75 $Y2=3.33
r236 54 59 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=9.75 $Y=3.245
+ $X2=9.75 $Y2=2.755
r237 50 53 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.85 $Y=2.025
+ $X2=8.85 $Y2=2.755
r238 48 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=3.245
+ $X2=8.85 $Y2=3.33
r239 48 53 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=8.85 $Y=3.245
+ $X2=8.85 $Y2=2.755
r240 44 139 2.80049 $w=6.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=3.245
+ $X2=7.685 $Y2=3.33
r241 44 46 9.76211 $w=6.78e-07 $l=5.55e-07 $layer=LI1_cond $X=7.685 $Y=3.245
+ $X2=7.685 $Y2=2.69
r242 40 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=3.33
r243 40 42 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=2.38
r244 36 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=3.245
+ $X2=4.525 $Y2=3.33
r245 36 38 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.525 $Y=3.245
+ $X2=4.525 $Y2=2.75
r246 32 130 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=3.33
r247 32 34 16.2988 $w=3.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=2.75
r248 28 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=3.33
r249 28 30 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=2.515
r250 9 71 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.835 $X2=11.71 $Y2=2.95
r251 9 68 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.835 $X2=11.71 $Y2=1.98
r252 8 65 300 $w=1.7e-07 $l=7.68473e-07 $layer=licon1_PDIFF $count=2 $X=10.555
+ $Y=1.835 $X2=10.85 $Y2=2.47
r253 8 62 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.555
+ $Y=1.835 $X2=10.695 $Y2=1.98
r254 7 59 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.57
+ $Y=1.64 $X2=9.71 $Y2=2.755
r255 7 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.57
+ $Y=1.64 $X2=9.71 $Y2=1.785
r256 6 53 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=8.615
+ $Y=2.48 $X2=8.85 $Y2=2.755
r257 6 50 300 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_PDIFF $count=2 $X=8.615
+ $Y=2.48 $X2=8.85 $Y2=2.025
r258 5 46 300 $w=1.7e-07 $l=6.21188e-07 $layer=licon1_PDIFF $count=2 $X=7.37
+ $Y=2.48 $X2=7.895 $Y2=2.69
r259 4 42 600 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.895 $X2=5.535 $Y2=2.38
r260 3 38 600 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=2.315 $X2=4.525 $Y2=2.75
r261 2 34 600 $w=1.7e-07 $l=5.29693e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=2.315 $X2=2.165 $Y2=2.75
r262 1 30 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.36 $X2=0.715 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%A_308_463# 1 2 3 4 13 17 21 25
c51 25 0 1.57615e-19 $X=2.922 $Y=2.425
r52 25 27 7.74185 $w=5.09e-07 $l=3.23e-07 $layer=LI1_cond $X=2.922 $Y=2.425
+ $X2=3.245 $Y2=2.425
r53 24 25 6.15992 $w=5.09e-07 $l=2.57e-07 $layer=LI1_cond $X=2.665 $Y=2.425
+ $X2=2.922 $Y2=2.425
r54 15 25 5.55206 $w=2.25e-07 $l=3.1e-07 $layer=LI1_cond $X=2.922 $Y=2.115
+ $X2=2.922 $Y2=2.425
r55 15 17 49.1709 $w=2.23e-07 $l=9.6e-07 $layer=LI1_cond $X=2.922 $Y=2.115
+ $X2=2.922 $Y2=1.155
r56 14 21 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.75 $Y=2.41 $X2=1.65
+ $Y2=2.41
r57 13 24 8.32598 $w=5.09e-07 $l=1.1225e-07 $layer=LI1_cond $X=2.56 $Y=2.41
+ $X2=2.665 $Y2=2.425
r58 13 14 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.56 $Y=2.41
+ $X2=1.75 $Y2=2.41
r59 4 27 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.315 $X2=3.245 $Y2=2.52
r60 3 24 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=2.315 $X2=2.665 $Y2=2.52
r61 2 21 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=2.315 $X2=1.665 $Y2=2.49
r62 1 17 182 $w=1.7e-07 $l=4.89898e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.955 $X2=2.895 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%Q_N 1 2 7 8 9 10 11 12 13 24 48
r21 28 48 1.10812 $w=2.58e-07 $l=2.5e-08 $layer=LI1_cond $X=9.325 $Y=0.95
+ $X2=9.325 $Y2=0.925
r22 12 13 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=9.325 $Y=2.405
+ $X2=9.325 $Y2=2.755
r23 11 12 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=9.325 $Y=2.035
+ $X2=9.325 $Y2=2.405
r24 11 36 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=9.325 $Y=2.035
+ $X2=9.325 $Y2=1.785
r25 10 36 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=9.325 $Y=1.665
+ $X2=9.325 $Y2=1.785
r26 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=9.325 $Y=1.295
+ $X2=9.325 $Y2=1.665
r27 8 48 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=9.325 $Y=0.895
+ $X2=9.325 $Y2=0.925
r28 8 46 4.18113 $w=2.58e-07 $l=7.5e-08 $layer=LI1_cond $X=9.325 $Y=0.895
+ $X2=9.325 $Y2=0.82
r29 8 9 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=9.325 $Y=0.965
+ $X2=9.325 $Y2=1.295
r30 8 28 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=9.325 $Y=0.965
+ $X2=9.325 $Y2=0.95
r31 7 46 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=9.36 $Y=0.555
+ $X2=9.36 $Y2=0.82
r32 7 24 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=9.36 $Y=0.555
+ $X2=9.36 $Y2=0.42
r33 2 13 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=1.64 $X2=9.28 $Y2=2.755
r34 2 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=1.64 $X2=9.28 $Y2=1.785
r35 1 8 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=9.22
+ $Y=0.25 $X2=9.36 $Y2=0.965
r36 1 24 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=9.22
+ $Y=0.25 $X2=9.36 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%Q 1 2 7 8 9 10 11 12 13
c17 7 0 5.41964e-20 $X=11.28 $Y=0.555
r18 13 39 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=11.297 $Y=2.775
+ $X2=11.297 $Y2=2.91
r19 12 13 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=11.297 $Y=2.405
+ $X2=11.297 $Y2=2.775
r20 11 12 21.7684 $w=2.23e-07 $l=4.25e-07 $layer=LI1_cond $X=11.297 $Y=1.98
+ $X2=11.297 $Y2=2.405
r21 10 11 16.1342 $w=2.23e-07 $l=3.15e-07 $layer=LI1_cond $X=11.297 $Y=1.665
+ $X2=11.297 $Y2=1.98
r22 9 10 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=11.297 $Y=1.295
+ $X2=11.297 $Y2=1.665
r23 8 9 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=11.297 $Y=0.925
+ $X2=11.297 $Y2=1.295
r24 7 8 21.7684 $w=2.23e-07 $l=4.25e-07 $layer=LI1_cond $X=11.297 $Y=0.5
+ $X2=11.297 $Y2=0.925
r25 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.14
+ $Y=1.835 $X2=11.28 $Y2=2.91
r26 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.14
+ $Y=1.835 $X2=11.28 $Y2=1.98
r27 1 7 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=11.14
+ $Y=0.345 $X2=11.28 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__DFRBP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 55
+ 57 60 61 62 64 69 74 86 90 95 100 106 109 112 115 118 121 125
r127 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r128 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r129 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r130 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r131 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r132 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r133 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r134 104 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r135 104 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r136 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r137 101 121 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=11.015 $Y=0
+ $X2=10.837 $Y2=0
r138 101 103 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.015 $Y=0
+ $X2=11.28 $Y2=0
r139 100 124 4.38626 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=11.58 $Y=0
+ $X2=11.79 $Y2=0
r140 100 103 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=11.58 $Y=0
+ $X2=11.28 $Y2=0
r141 99 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r142 99 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r143 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r144 96 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.955 $Y=0
+ $X2=9.79 $Y2=0
r145 96 98 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.955 $Y=0
+ $X2=10.32 $Y2=0
r146 95 121 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=10.66 $Y=0
+ $X2=10.837 $Y2=0
r147 95 98 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.66 $Y=0
+ $X2=10.32 $Y2=0
r148 94 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r149 94 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r150 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r151 91 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.095 $Y=0
+ $X2=8.93 $Y2=0
r152 91 93 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.095 $Y=0
+ $X2=9.36 $Y2=0
r153 90 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.625 $Y=0
+ $X2=9.79 $Y2=0
r154 90 93 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.625 $Y=0
+ $X2=9.36 $Y2=0
r155 89 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r156 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r157 86 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.765 $Y=0
+ $X2=8.93 $Y2=0
r158 86 88 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.765 $Y=0 $X2=8.4
+ $Y2=0
r159 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r160 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r161 82 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.575 $Y=0
+ $X2=5.41 $Y2=0
r162 82 84 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=5.575 $Y=0
+ $X2=7.44 $Y2=0
r163 81 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r164 80 81 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r165 78 81 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=5.04 $Y2=0
r166 78 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r167 77 80 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=5.04
+ $Y2=0
r168 77 78 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r169 75 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0
+ $X2=1.74 $Y2=0
r170 75 77 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=0
+ $X2=2.16 $Y2=0
r171 74 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.245 $Y=0
+ $X2=5.41 $Y2=0
r172 74 80 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.245 $Y=0
+ $X2=5.04 $Y2=0
r173 73 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r174 73 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r175 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r176 70 106 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.7
+ $Y2=0
r177 70 72 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.2
+ $Y2=0
r178 69 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=0
+ $X2=1.74 $Y2=0
r179 69 72 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.2
+ $Y2=0
r180 67 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r181 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r182 64 106 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.7
+ $Y2=0
r183 64 66 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.24
+ $Y2=0
r184 62 85 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=0 $X2=7.44
+ $Y2=0
r185 62 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r186 60 84 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.455 $Y=0 $X2=7.44
+ $Y2=0
r187 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=0 $X2=7.62
+ $Y2=0
r188 59 88 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.785 $Y=0 $X2=8.4
+ $Y2=0
r189 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.785 $Y=0 $X2=7.62
+ $Y2=0
r190 55 124 3.09127 $w=2.95e-07 $l=1.12161e-07 $layer=LI1_cond $X=11.727
+ $Y=0.085 $X2=11.79 $Y2=0
r191 55 57 15.8217 $w=2.93e-07 $l=4.05e-07 $layer=LI1_cond $X=11.727 $Y=0.085
+ $X2=11.727 $Y2=0.49
r192 51 53 17.2055 $w=3.53e-07 $l=5.3e-07 $layer=LI1_cond $X=10.837 $Y=0.49
+ $X2=10.837 $Y2=1.02
r193 49 121 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=10.837 $Y=0.085
+ $X2=10.837 $Y2=0
r194 49 51 13.1476 $w=3.53e-07 $l=4.05e-07 $layer=LI1_cond $X=10.837 $Y=0.085
+ $X2=10.837 $Y2=0.49
r195 45 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=0.085
+ $X2=9.79 $Y2=0
r196 45 47 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=9.79 $Y=0.085
+ $X2=9.79 $Y2=0.395
r197 41 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.93 $Y=0.085
+ $X2=8.93 $Y2=0
r198 41 43 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=8.93 $Y=0.085
+ $X2=8.93 $Y2=0.52
r199 37 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.62 $Y=0.085
+ $X2=7.62 $Y2=0
r200 37 39 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=7.62 $Y=0.085
+ $X2=7.62 $Y2=0.85
r201 33 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=0.085
+ $X2=5.41 $Y2=0
r202 33 35 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=0.085
+ $X2=5.41 $Y2=0.455
r203 29 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0
r204 29 31 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0.59
r205 25 106 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0
r206 25 27 22.384 $w=2.58e-07 $l=5.05e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.59
r207 8 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.57
+ $Y=0.345 $X2=11.71 $Y2=0.49
r208 7 53 182 $w=1.7e-07 $l=7.83741e-07 $layer=licon1_NDIFF $count=1 $X=10.615
+ $Y=0.345 $X2=10.85 $Y2=1.02
r209 7 51 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=10.615
+ $Y=0.345 $X2=10.755 $Y2=0.49
r210 6 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.65
+ $Y=0.25 $X2=9.79 $Y2=0.395
r211 5 43 182 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_NDIFF $count=1 $X=8.805
+ $Y=0.25 $X2=8.93 $Y2=0.52
r212 4 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.48
+ $Y=0.64 $X2=7.62 $Y2=0.85
r213 3 35 182 $w=1.7e-07 $l=8.95768e-07 $layer=licon1_NDIFF $count=1 $X=4.73
+ $Y=0.955 $X2=5.41 $Y2=0.455
r214 2 31 182 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.43 $X2=1.74 $Y2=0.59
r215 1 27 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.395 $X2=0.69 $Y2=0.59
.ends

