* File: sky130_fd_sc_lp__a22o_m.pex.spice
* Created: Fri Aug 28 09:54:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22O_M%A_85_317# 1 2 9 13 17 19 20 21 22 24 27 30 35
+ 37
c80 9 0 1.59309e-19 $X=0.66 $Y=2.715
r81 37 40 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.01 $Y=2.41
+ $X2=2.01 $Y2=2.63
r82 32 35 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.71 $Y=0.81
+ $X2=1.825 $Y2=0.81
r83 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.75 $X2=0.59 $Y2=1.75
r84 26 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0.975
+ $X2=1.71 $Y2=0.81
r85 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.71 $Y=0.975
+ $X2=1.71 $Y2=1.585
r86 24 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.41
+ $X2=2.01 $Y2=2.41
r87 24 25 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.845 $Y=2.41
+ $X2=0.935 $Y2=2.41
r88 23 29 6.18617 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=1.67
+ $X2=0.72 $Y2=1.67
r89 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.625 $Y=1.67
+ $X2=1.71 $Y2=1.585
r90 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.625 $Y=1.67
+ $X2=0.935 $Y2=1.67
r91 21 25 11.7614 $w=4.3e-07 $l=4.65242e-07 $layer=LI1_cond $X=0.72 $Y=2.04
+ $X2=0.935 $Y2=2.41
r92 20 29 2.44569 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.755
+ $X2=0.72 $Y2=1.67
r93 20 21 7.63829 $w=4.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=1.755
+ $X2=0.72 $Y2=2.04
r94 18 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=2.09
+ $X2=0.59 $Y2=1.75
r95 18 19 43.0552 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=2.09
+ $X2=0.59 $Y2=2.255
r96 17 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.59 $Y=1.735
+ $X2=0.59 $Y2=1.75
r97 16 17 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.605 $Y=1.585
+ $X2=0.605 $Y2=1.735
r98 13 16 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.71 $Y=0.835
+ $X2=0.71 $Y2=1.585
r99 9 19 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.66 $Y=2.715
+ $X2=0.66 $Y2=2.255
r100 2 40 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=1.755
+ $Y=2.505 $X2=2.01 $Y2=2.63
r101 1 35 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.625 $X2=1.825 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%A2 3 6 8 9 13 15
c38 6 0 7.92268e-20 $X=1.25 $Y=2.715
r39 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.32
+ $X2=1.16 $Y2=1.485
r40 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.32
+ $X2=1.16 $Y2=1.155
r41 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.32 $X2=1.16 $Y2=1.32
r42 8 9 25.0256 $w=1.93e-07 $l=4.4e-07 $layer=LI1_cond $X=0.72 $Y=1.307 $X2=1.16
+ $Y2=1.307
r43 6 16 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.25 $Y=2.715
+ $X2=1.25 $Y2=1.485
r44 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.25 $Y=0.835
+ $X2=1.25 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%A1 3 6 10 11 14 18 19 20 21 28 33 45
c58 33 0 1.81351e-20 $X=1.7 $Y=0.515
c59 28 0 1.61987e-19 $X=2.96 $Y=1.775
r60 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.96
+ $Y=1.775 $X2=2.96 $Y2=1.775
r61 20 21 7.50083 $w=5.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.91 $Y=2.035
+ $X2=2.91 $Y2=2.405
r62 20 29 5.27085 $w=5.88e-07 $l=2.6e-07 $layer=LI1_cond $X=2.91 $Y=2.035
+ $X2=2.91 $Y2=1.775
r63 19 29 2.22998 $w=5.88e-07 $l=1.1e-07 $layer=LI1_cond $X=2.91 $Y=1.665
+ $X2=2.91 $Y2=1.775
r64 18 45 9.92676 $w=7.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.825 $Y=1.295
+ $X2=2.825 $Y2=1.21
r65 18 19 5.11545 $w=7.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.91 $Y=1.38
+ $X2=2.91 $Y2=1.665
r66 16 45 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.53 $Y=0.435
+ $X2=2.53 $Y2=1.21
r67 14 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=0.35 $X2=1.7
+ $Y2=0.515
r68 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=0.35 $X2=1.7 $Y2=0.35
r69 11 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=0.35
+ $X2=2.53 $Y2=0.435
r70 11 13 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.445 $Y=0.35
+ $X2=1.7 $Y2=0.35
r71 9 28 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.96 $Y=2.13
+ $X2=2.96 $Y2=1.775
r72 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.91 $Y=2.13 $X2=2.91
+ $Y2=2.28
r73 6 10 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=2.77 $Y=2.755
+ $X2=2.77 $Y2=2.28
r74 3 33 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.61 $Y=0.835
+ $X2=1.61 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%B1 3 5 7 8 9 14
c40 8 0 1.81351e-20 $X=2.16 $Y=1.295
c41 3 0 3.56444e-20 $X=1.68 $Y=2.715
r42 14 16 16.3698 $w=2.65e-07 $l=9e-08 $layer=POLY_cond $X=2.06 $Y=1.36 $X2=2.15
+ $Y2=1.36
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.32 $X2=2.06 $Y2=1.32
r44 9 15 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.11 $Y=1.665
+ $X2=2.11 $Y2=1.32
r45 8 15 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.11 $Y=1.295
+ $X2=2.11 $Y2=1.32
r46 5 16 16.0701 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.15 $Y=1.155
+ $X2=2.15 $Y2=1.36
r47 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.15 $Y=1.155 $X2=2.15
+ $Y2=0.835
r48 1 14 69.117 $w=2.65e-07 $l=4.71487e-07 $layer=POLY_cond $X=1.68 $Y=1.565
+ $X2=2.06 $Y2=1.36
r49 1 3 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=1.68 $Y=1.565
+ $X2=1.68 $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%B2 1 3 7 9 10 11 17
c44 17 0 1.61987e-19 $X=2.27 $Y=2.035
c45 3 0 1.70555e-19 $X=2.34 $Y=2.755
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.27
+ $Y=2.035 $X2=2.27 $Y2=2.035
r47 11 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.27 $Y2=2.035
r48 10 11 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=2.16 $Y2=2.035
r49 9 10 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.035 $X2=1.68
+ $Y2=2.035
r50 5 16 65.5678 $w=3.12e-07 $l=4.14367e-07 $layer=POLY_cond $X=2.51 $Y=1.695
+ $X2=2.345 $Y2=2.035
r51 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.51 $Y=1.695 $X2=2.51
+ $Y2=0.835
r52 1 16 38.5325 $w=3.12e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.34 $Y=2.2
+ $X2=2.345 $Y2=2.035
r53 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.34 $Y=2.2 $X2=2.34
+ $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%X 1 2 7 9 12 13 14 15 16 35
r22 16 35 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.24 $Y=2.695
+ $X2=0.445 $Y2=2.695
r23 16 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=2.695
+ $X2=0.24 $Y2=2.53
r24 15 22 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.53
r25 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r26 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r27 12 13 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r28 11 12 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.24 $Y=1.005
+ $X2=0.24 $Y2=1.295
r29 7 11 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.325 $Y=0.9
+ $X2=0.24 $Y2=1.005
r30 7 9 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.325 $Y=0.9 $X2=0.475
+ $Y2=0.9
r31 2 35 600 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=1 $X=0.32
+ $Y=2.505 $X2=0.445 $Y2=2.695
r32 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.35
+ $Y=0.625 $X2=0.475 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%VPWR 1 2 9 11 13 16 17 18 24 33
c37 33 0 3.56444e-20 $X=3.12 $Y=3.33
c38 13 0 1.70555e-19 $X=3.005 $Y=2.82
r39 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 24 32 4.5891 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.84 $Y=3.33 $X2=3.1
+ $Y2=3.33
r45 24 29 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.84 $Y=3.33 $X2=2.64
+ $Y2=3.33
r46 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 18 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 16 21 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.73 $Y=3.33 $X2=0.72
+ $Y2=3.33
r51 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=3.33
+ $X2=0.895 $Y2=3.33
r52 15 26 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.06 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.895 $Y2=3.33
r54 11 32 3.17707 $w=3.3e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.005 $Y=3.245
+ $X2=3.1 $Y2=3.33
r55 11 13 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=3.005 $Y=3.245
+ $X2=3.005 $Y2=2.82
r56 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=3.33
r57 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=2.78
r58 2 13 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=2.545 $X2=3.005 $Y2=2.82
r59 1 9 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=2.505 $X2=0.895 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%A_265_501# 1 2 7 10 15
c25 10 0 1.59309e-19 $X=1.465 $Y=2.78
c26 7 0 7.92268e-20 $X=2.45 $Y=2.98
r27 15 17 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=2.555 $Y=2.84
+ $X2=2.555 $Y2=2.98
r28 10 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.465 $Y=2.78 $X2=1.465
+ $Y2=2.98
r29 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=2.98
+ $X2=1.465 $Y2=2.98
r30 7 17 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.45 $Y=2.98 $X2=2.555
+ $Y2=2.98
r31 7 8 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.45 $Y=2.98 $X2=1.63
+ $Y2=2.98
r32 2 15 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.545 $X2=2.555 $Y2=2.84
r33 1 10 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=2.505 $X2=1.465 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_M%VGND 1 2 9 13 16 17 19 20 21 34 35
r30 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r31 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r32 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r33 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r34 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r36 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 21 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r38 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r39 19 31 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.64
+ $Y2=0
r40 19 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.89
+ $Y2=0
r41 18 34 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=3.12
+ $Y2=0
r42 18 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.89
+ $Y2=0
r43 16 24 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.72
+ $Y2=0
r44 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.985
+ $Y2=0
r45 15 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.2
+ $Y2=0
r46 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=0.985
+ $Y2=0
r47 11 20 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0
r48 11 13 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0.77
r49 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0
r50 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0.77
r51 2 13 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.625 $X2=2.88 $Y2=0.77
r52 1 9 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.785
+ $Y=0.625 $X2=0.985 $Y2=0.77
.ends

