* NGSPICE file created from sky130_fd_sc_lp__clkinv_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__clkinv_lp A VGND VNB VPB VPWR Y
M1000 a_124_92# A VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_124_468# A VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.824e+11p ps=1.85e+06u
M1002 Y A a_124_92# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 Y A a_124_468# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
.ends

