* File: sky130_fd_sc_lp__o2bb2a_4.pex.spice
* Created: Wed Sep  2 10:21:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%B1 3 7 11 15 17 20 23 25 27 28 31 32 33 34
c89 23 0 5.31934e-20 $X=0.72 $Y=2.31
c90 11 0 1.10714e-19 $X=1.875 $Y=2.465
c91 7 0 1.91137e-19 $X=0.585 $Y=2.465
r92 33 34 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.405
+ $X2=1.68 $Y2=2.405
r93 33 44 22.4737 $w=1.88e-07 $l=3.85e-07 $layer=LI1_cond $X=1.2 $Y=2.405
+ $X2=0.815 $Y2=2.405
r94 32 44 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.815 $Y2=2.405
r95 31 34 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.405
+ $X2=1.68 $Y2=2.405
r96 28 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=1.51
+ $X2=1.93 $Y2=1.675
r97 28 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=1.51
+ $X2=1.93 $Y2=1.345
r98 27 30 7.37583 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.97 $Y=1.51
+ $X2=1.97 $Y2=1.65
r99 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.51 $X2=1.93 $Y2=1.51
r100 25 31 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=1.935 $Y=2.31
+ $X2=1.845 $Y2=2.405
r101 25 30 40.6667 $w=1.78e-07 $l=6.6e-07 $layer=LI1_cond $X=1.935 $Y=2.31
+ $X2=1.935 $Y2=1.65
r102 23 32 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=2.31
+ $X2=0.72 $Y2=2.405
r103 22 23 38.8182 $w=1.88e-07 $l=6.65e-07 $layer=LI1_cond $X=0.72 $Y=1.645
+ $X2=0.72 $Y2=2.31
r104 20 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.495 $Y2=1.675
r105 20 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.495 $Y2=1.345
r106 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.495
+ $Y=1.51 $X2=0.495 $Y2=1.51
r107 17 22 6.93705 $w=2.4e-07 $l=1.60624e-07 $layer=LI1_cond $X=0.625 $Y=1.525
+ $X2=0.72 $Y2=1.645
r108 17 19 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.625 $Y=1.525
+ $X2=0.495 $Y2=1.525
r109 15 42 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.955 $Y=0.655
+ $X2=1.955 $Y2=1.345
r110 11 43 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.875 $Y=2.465
+ $X2=1.875 $Y2=1.675
r111 7 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.585 $Y=2.465
+ $X2=0.585 $Y2=1.675
r112 3 39 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.585 $Y=0.655
+ $X2=0.585 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%B2 3 7 11 15 17 23 24
c54 3 0 7.75885e-20 $X=1.015 $Y=0.655
r55 22 24 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.15 $Y=1.51
+ $X2=1.445 $Y2=1.51
r56 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.51 $X2=1.15 $Y2=1.51
r57 19 22 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.015 $Y=1.51
+ $X2=1.15 $Y2=1.51
r58 17 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.51
r59 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=1.51
r60 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=2.465
r61 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.345
+ $X2=1.445 $Y2=1.51
r62 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.445 $Y=1.345
+ $X2=1.445 $Y2=0.655
r63 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=1.51
r64 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=2.465
r65 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.345
+ $X2=1.015 $Y2=1.51
r66 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.015 $Y=1.345
+ $X2=1.015 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%A_462_21# 1 2 3 10 12 15 17 19 22 24 27 30
+ 32 34 35 39 41 43 44
c116 17 0 1.99532e-19 $X=2.815 $Y=1.185
c117 10 0 1.95499e-19 $X=2.385 $Y=1.185
r118 49 50 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.35
+ $X2=2.98 $Y2=1.35
r119 48 49 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=2.55 $Y=1.35
+ $X2=2.815 $Y2=1.35
r120 46 48 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.35
+ $X2=2.55 $Y2=1.35
r121 43 44 8.17035 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=0.785
+ $X2=4.245 $Y2=0.785
r122 37 39 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=3.965 $Y=2.095
+ $X2=4.84 $Y2=2.095
r123 35 37 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=3.475 $Y=2.095
+ $X2=3.965 $Y2=2.095
r124 34 44 44.9474 $w=1.88e-07 $l=7.7e-07 $layer=LI1_cond $X=3.475 $Y=0.82
+ $X2=4.245 $Y2=0.82
r125 32 35 7.61292 $w=3.3e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.385 $Y=1.93
+ $X2=3.475 $Y2=2.095
r126 31 41 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=1.515
+ $X2=3.385 $Y2=1.35
r127 31 32 25.5707 $w=1.78e-07 $l=4.15e-07 $layer=LI1_cond $X=3.385 $Y=1.515
+ $X2=3.385 $Y2=1.93
r128 30 41 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=1.185
+ $X2=3.385 $Y2=1.35
r129 29 34 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.385 $Y=0.915
+ $X2=3.475 $Y2=0.82
r130 29 30 16.6364 $w=1.78e-07 $l=2.7e-07 $layer=LI1_cond $X=3.385 $Y=0.915
+ $X2=3.385 $Y2=1.185
r131 27 50 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.015 $Y=1.35
+ $X2=2.98 $Y2=1.35
r132 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.015
+ $Y=1.35 $X2=3.015 $Y2=1.35
r133 24 41 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.295 $Y=1.35
+ $X2=3.385 $Y2=1.35
r134 24 26 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.295 $Y=1.35
+ $X2=3.015 $Y2=1.35
r135 20 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=2.98 $Y2=1.35
r136 20 22 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.98 $Y=1.515
+ $X2=2.98 $Y2=2.465
r137 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.185
+ $X2=2.815 $Y2=1.35
r138 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.815 $Y=1.185
+ $X2=2.815 $Y2=0.655
r139 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.55 $Y2=1.35
r140 13 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.55 $Y=1.515
+ $X2=2.55 $Y2=2.465
r141 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.185
+ $X2=2.385 $Y2=1.35
r142 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.385 $Y=1.185
+ $X2=2.385 $Y2=0.655
r143 3 39 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=4.7
+ $Y=1.835 $X2=4.84 $Y2=2.095
r144 2 37 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=1.835 $X2=3.965 $Y2=2.095
r145 1 43 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.235 $X2=4.41 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%A1_N 3 7 10 13 15 17 21 23 26 28 31 37
c84 26 0 5.09057e-20 $X=3.73 $Y=1.35
c85 17 0 8.01762e-20 $X=5.045 $Y=1.17
r86 26 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.35
+ $X2=3.73 $Y2=1.515
r87 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.35
+ $X2=3.73 $Y2=1.185
r88 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.35 $X2=3.73 $Y2=1.35
r89 23 37 6.90882 $w=4.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.08 $Y=1.3
+ $X2=4.175 $Y2=1.3
r90 23 27 9.38035 $w=4.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.08 $Y=1.3 $X2=3.73
+ $Y2=1.3
r91 21 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.075 $Y=1.35
+ $X2=5.075 $Y2=1.515
r92 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.075 $Y=1.35
+ $X2=5.075 $Y2=1.185
r93 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.075
+ $Y=1.35 $X2=5.075 $Y2=1.35
r94 17 20 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=5.045 $Y=1.17
+ $X2=5.045 $Y2=1.35
r95 15 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.92 $Y=1.17
+ $X2=5.045 $Y2=1.17
r96 15 37 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.92 $Y=1.17
+ $X2=4.175 $Y2=1.17
r97 13 32 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.055 $Y=2.465
+ $X2=5.055 $Y2=1.515
r98 10 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.055 $Y=0.655
+ $X2=5.055 $Y2=1.185
r99 7 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.765 $Y=0.655
+ $X2=3.765 $Y2=1.185
r100 3 29 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.75 $Y=2.465
+ $X2=3.75 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%A2_N 1 3 4 6 7 9 10 12 13 19 20
c52 19 0 5.09057e-20 $X=4.51 $Y=1.51
c53 7 0 8.01762e-20 $X=4.625 $Y=1.185
r54 18 20 10.4585 $w=5.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.51 $Y=1.455
+ $X2=4.625 $Y2=1.455
r55 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.51 $X2=4.51 $Y2=1.51
r56 16 18 28.6472 $w=5.3e-07 $l=3.15e-07 $layer=POLY_cond $X=4.195 $Y=1.455
+ $X2=4.51 $Y2=1.455
r57 15 16 1.36415 $w=5.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.18 $Y=1.455
+ $X2=4.195 $Y2=1.455
r58 13 19 4.41058 $w=4.03e-07 $l=1.55e-07 $layer=LI1_cond $X=4.547 $Y=1.665
+ $X2=4.547 $Y2=1.51
r59 10 20 32.8864 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.625 $Y=1.725
+ $X2=4.625 $Y2=1.455
r60 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.625 $Y=1.725
+ $X2=4.625 $Y2=2.465
r61 7 20 32.8864 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.625 $Y=1.185
+ $X2=4.625 $Y2=1.455
r62 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.625 $Y=1.185
+ $X2=4.625 $Y2=0.655
r63 4 16 32.8864 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.195 $Y=1.185
+ $X2=4.195 $Y2=1.455
r64 4 6 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.195 $Y=1.185
+ $X2=4.195 $Y2=0.655
r65 1 15 32.8864 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.18 $Y=1.725
+ $X2=4.18 $Y2=1.455
r66 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.18 $Y=1.725 $X2=4.18
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%A_218_367# 1 2 3 12 16 20 24 28 32 36 40 42
+ 47 48 49 52 56 59 62 64 67 68 73 76 77 78 89
c186 77 0 3.95031e-19 $X=2.76 $Y=1.73
c187 62 0 1.10714e-19 $X=2.765 $Y=2.91
c188 49 0 7.75885e-20 $X=1.665 $Y=1.085
c189 42 0 1.91137e-19 $X=1.485 $Y=2.035
r190 86 87 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.685 $Y=1.49
+ $X2=6.85 $Y2=1.49
r191 85 86 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.42 $Y=1.49
+ $X2=6.685 $Y2=1.49
r192 84 85 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.49
+ $X2=6.42 $Y2=1.49
r193 83 84 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=5.99 $Y=1.49
+ $X2=6.255 $Y2=1.49
r194 82 83 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.49
+ $X2=5.99 $Y2=1.49
r195 74 89 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=7.01 $Y=1.49
+ $X2=7.115 $Y2=1.49
r196 74 87 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=7.01 $Y=1.49
+ $X2=6.85 $Y2=1.49
r197 73 74 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.01
+ $Y=1.49 $X2=7.01 $Y2=1.49
r198 71 82 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.65 $Y=1.49
+ $X2=5.825 $Y2=1.49
r199 71 79 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.65 $Y=1.49 $X2=5.56
+ $Y2=1.49
r200 70 73 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=5.65 $Y=1.49
+ $X2=7.01 $Y2=1.49
r201 70 71 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.65
+ $Y=1.49 $X2=5.65 $Y2=1.49
r202 68 70 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.51 $Y=1.49
+ $X2=5.65 $Y2=1.49
r203 66 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.425 $Y=1.575
+ $X2=5.51 $Y2=1.49
r204 66 67 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=5.425 $Y=1.575
+ $X2=5.425 $Y2=2.43
r205 65 78 3.29449 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=2.93 $Y=2.52
+ $X2=2.76 $Y2=2.52
r206 64 67 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.34 $Y=2.52
+ $X2=5.425 $Y2=2.43
r207 64 65 148.495 $w=1.78e-07 $l=2.41e-06 $layer=LI1_cond $X=5.34 $Y=2.52
+ $X2=2.93 $Y2=2.52
r208 60 78 3.2666 $w=3.05e-07 $l=1.06066e-07 $layer=LI1_cond $X=2.725 $Y=2.61
+ $X2=2.76 $Y2=2.52
r209 60 62 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=2.725 $Y=2.61
+ $X2=2.725 $Y2=2.91
r210 57 78 3.2666 $w=3.05e-07 $l=9e-08 $layer=LI1_cond $X=2.76 $Y=2.43 $X2=2.76
+ $Y2=2.52
r211 57 59 15.2529 $w=3.38e-07 $l=4.5e-07 $layer=LI1_cond $X=2.76 $Y=2.43
+ $X2=2.76 $Y2=1.98
r212 56 77 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.76 $Y=1.9
+ $X2=2.76 $Y2=1.73
r213 56 59 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=2.76 $Y=1.9 $X2=2.76
+ $Y2=1.98
r214 54 76 4.48993 $w=2.12e-07 $l=1.09407e-07 $layer=LI1_cond $X=2.675 $Y=1.175
+ $X2=2.632 $Y2=1.085
r215 54 77 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.675 $Y=1.175
+ $X2=2.675 $Y2=1.73
r216 50 76 4.48993 $w=2.12e-07 $l=9e-08 $layer=LI1_cond $X=2.632 $Y=0.995
+ $X2=2.632 $Y2=1.085
r217 50 52 10.1686 $w=2.53e-07 $l=2.25e-07 $layer=LI1_cond $X=2.632 $Y=0.995
+ $X2=2.632 $Y2=0.77
r218 48 76 1.94654 $w=1.8e-07 $l=1.27e-07 $layer=LI1_cond $X=2.505 $Y=1.085
+ $X2=2.632 $Y2=1.085
r219 48 49 51.7576 $w=1.78e-07 $l=8.4e-07 $layer=LI1_cond $X=2.505 $Y=1.085
+ $X2=1.665 $Y2=1.085
r220 46 49 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=1.575 $Y=1.175
+ $X2=1.665 $Y2=1.085
r221 46 47 46.5202 $w=1.78e-07 $l=7.55e-07 $layer=LI1_cond $X=1.575 $Y=1.175
+ $X2=1.575 $Y2=1.93
r222 42 47 6.86909 $w=2.1e-07 $l=1.43091e-07 $layer=LI1_cond $X=1.485 $Y=2.035
+ $X2=1.575 $Y2=1.93
r223 42 44 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=1.485 $Y=2.035
+ $X2=1.23 $Y2=2.035
r224 38 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.115 $Y=1.325
+ $X2=7.115 $Y2=1.49
r225 38 40 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.115 $Y=1.325
+ $X2=7.115 $Y2=0.655
r226 34 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.85 $Y=1.655
+ $X2=6.85 $Y2=1.49
r227 34 36 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.85 $Y=1.655
+ $X2=6.85 $Y2=2.465
r228 30 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.685 $Y=1.325
+ $X2=6.685 $Y2=1.49
r229 30 32 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.685 $Y=1.325
+ $X2=6.685 $Y2=0.655
r230 26 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.42 $Y=1.655
+ $X2=6.42 $Y2=1.49
r231 26 28 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.42 $Y=1.655
+ $X2=6.42 $Y2=2.465
r232 22 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.325
+ $X2=6.255 $Y2=1.49
r233 22 24 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.255 $Y=1.325
+ $X2=6.255 $Y2=0.655
r234 18 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.99 $Y=1.655
+ $X2=5.99 $Y2=1.49
r235 18 20 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.99 $Y=1.655
+ $X2=5.99 $Y2=2.465
r236 14 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=1.49
r237 14 16 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=0.655
r238 10 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=1.655
+ $X2=5.56 $Y2=1.49
r239 10 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.56 $Y=1.655
+ $X2=5.56 $Y2=2.465
r240 3 62 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=1.835 $X2=2.765 $Y2=2.91
r241 3 59 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.625
+ $Y=1.835 $X2=2.765 $Y2=1.98
r242 2 44 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.835 $X2=1.23 $Y2=2.035
r243 1 52 182 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.235 $X2=2.6 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%VPWR 1 2 3 4 5 6 7 22 24 28 31 34 40 44 48
+ 52 56 62 63 65 66 67 68 69 71 96 97 103 107 111 113
r125 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 109 111 9.15996 $w=6.33e-07 $l=1e-07 $layer=LI1_cond $X=3.6 $Y=3.097
+ $X2=3.7 $Y2=3.097
r127 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r128 106 109 1.22433 $w=6.33e-07 $l=6.5e-08 $layer=LI1_cond $X=3.535 $Y=3.097
+ $X2=3.6 $Y2=3.097
r129 106 107 16.7885 $w=6.33e-07 $l=5.05e-07 $layer=LI1_cond $X=3.535 $Y=3.097
+ $X2=3.03 $Y2=3.097
r130 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r131 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 97 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r133 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r134 94 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=3.33
+ $X2=7.065 $Y2=3.33
r135 94 96 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.23 $Y=3.33
+ $X2=7.44 $Y2=3.33
r136 93 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r137 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r138 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r139 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r140 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r141 86 111 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.7 $Y2=3.33
r142 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 83 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r144 83 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 82 107 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=3.03 $Y2=3.33
r146 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r147 80 103 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.177 $Y2=3.33
r148 80 82 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.64 $Y2=3.33
r149 78 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r150 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r152 75 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 74 77 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r154 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r155 72 100 3.915 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r156 72 74 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.72 $Y2=3.33
r157 71 103 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.177 $Y2=3.33
r158 71 77 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r159 69 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r160 69 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 67 92 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.04 $Y=3.33 $X2=6
+ $Y2=3.33
r162 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.04 $Y=3.33
+ $X2=6.205 $Y2=3.33
r163 65 89 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.105 $Y=3.33
+ $X2=5.04 $Y2=3.33
r164 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=3.33
+ $X2=5.27 $Y2=3.33
r165 64 92 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.435 $Y=3.33 $X2=6
+ $Y2=3.33
r166 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.27 $Y2=3.33
r167 62 86 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.23 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=3.33
+ $X2=4.395 $Y2=3.33
r169 61 89 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r170 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=4.395 $Y2=3.33
r171 56 59 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=7.065 $Y=2.18
+ $X2=7.065 $Y2=2.95
r172 54 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=3.245
+ $X2=7.065 $Y2=3.33
r173 54 59 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.065 $Y=3.245
+ $X2=7.065 $Y2=2.95
r174 53 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.37 $Y=3.33
+ $X2=6.205 $Y2=3.33
r175 52 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.9 $Y=3.33
+ $X2=7.065 $Y2=3.33
r176 52 53 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.9 $Y=3.33
+ $X2=6.37 $Y2=3.33
r177 48 51 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.205 $Y=2.18
+ $X2=6.205 $Y2=2.95
r178 46 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.205 $Y=3.245
+ $X2=6.205 $Y2=3.33
r179 46 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.205 $Y=3.245
+ $X2=6.205 $Y2=2.95
r180 42 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=3.245
+ $X2=5.27 $Y2=3.33
r181 42 44 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.27 $Y=3.245
+ $X2=5.27 $Y2=2.89
r182 38 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.395 $Y=3.245
+ $X2=4.395 $Y2=3.33
r183 38 40 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.395 $Y=3.245
+ $X2=4.395 $Y2=2.89
r184 37 60 1.53659 $w=2.23e-07 $l=3e-08 $layer=LI1_cond $X=2.307 $Y=2.64
+ $X2=2.307 $Y2=2.67
r185 34 37 34.8294 $w=2.23e-07 $l=6.8e-07 $layer=LI1_cond $X=2.307 $Y=1.96
+ $X2=2.307 $Y2=2.64
r186 29 103 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.177 $Y=3.245
+ $X2=2.177 $Y2=3.33
r187 29 31 6.90519 $w=4.83e-07 $l=2.8e-07 $layer=LI1_cond $X=2.177 $Y=3.245
+ $X2=2.177 $Y2=2.965
r188 28 60 9.43373 $w=4.83e-07 $l=2.42e-07 $layer=LI1_cond $X=2.177 $Y=2.912
+ $X2=2.177 $Y2=2.67
r189 28 31 1.30705 $w=4.83e-07 $l=5.3e-08 $layer=LI1_cond $X=2.177 $Y=2.912
+ $X2=2.177 $Y2=2.965
r190 24 27 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=0.33 $Y=1.98
+ $X2=0.33 $Y2=2.95
r191 22 100 3.22816 $w=2.5e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.227 $Y2=3.33
r192 22 27 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.33 $Y2=2.95
r193 7 59 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.925
+ $Y=1.835 $X2=7.065 $Y2=2.95
r194 7 56 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=6.925
+ $Y=1.835 $X2=7.065 $Y2=2.18
r195 6 51 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.065
+ $Y=1.835 $X2=6.205 $Y2=2.95
r196 6 48 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=6.065
+ $Y=1.835 $X2=6.205 $Y2=2.18
r197 5 44 600 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=5.13
+ $Y=1.835 $X2=5.27 $Y2=2.89
r198 4 40 600 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.835 $X2=4.395 $Y2=2.89
r199 3 106 300 $w=1.7e-07 $l=1.27257e-06 $layer=licon1_PDIFF $count=2 $X=3.055
+ $Y=1.835 $X2=3.535 $Y2=2.89
r200 2 37 400 $w=1.7e-07 $l=9.78749e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.335 $Y2=2.64
r201 2 34 400 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.335 $Y2=1.96
r202 2 31 600 $w=1.7e-07 $l=1.19796e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.09 $Y2=2.965
r203 1 27 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.95
r204 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%A_132_367# 1 2 11
r15 8 11 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=0.8 $Y=2.835 $X2=1.66
+ $Y2=2.835
r16 2 11 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.835 $X2=1.66 $Y2=2.835
r17 1 8 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%X 1 2 3 4 15 19 20 23 25 26 29 33 37 39 41
+ 42 43 44 49 50 52 56
r63 50 56 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=7.47 $Y=1.745 $X2=7.47
+ $Y2=1.665
r64 49 52 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=7.47 $Y=1.235 $X2=7.47
+ $Y2=1.295
r65 44 50 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=7.47 $Y=1.835 $X2=7.47
+ $Y2=1.745
r66 44 56 0.138293 $w=2.48e-07 $l=3e-09 $layer=LI1_cond $X=7.47 $Y=1.662
+ $X2=7.47 $Y2=1.665
r67 43 49 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=7.47 $Y=1.14 $X2=7.47
+ $Y2=1.235
r68 43 44 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=7.47 $Y=1.307
+ $X2=7.47 $Y2=1.662
r69 43 52 0.553173 $w=2.48e-07 $l=1.2e-08 $layer=LI1_cond $X=7.47 $Y=1.307
+ $X2=7.47 $Y2=1.295
r70 40 42 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=6.995 $Y=1.14 $X2=6.9
+ $Y2=1.14
r71 39 43 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=7.345 $Y=1.14
+ $X2=7.47 $Y2=1.14
r72 39 40 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=7.345 $Y=1.14
+ $X2=6.995 $Y2=1.14
r73 35 42 1.34256 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=6.9 $Y=1.045 $X2=6.9
+ $Y2=1.14
r74 35 37 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=6.9 $Y=1.045
+ $X2=6.9 $Y2=0.42
r75 34 41 5.16603 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=6.72 $Y=1.835 $X2=6.63
+ $Y2=1.835
r76 33 44 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=7.345 $Y=1.835
+ $X2=7.47 $Y2=1.835
r77 33 34 38.5101 $w=1.78e-07 $l=6.25e-07 $layer=LI1_cond $X=7.345 $Y=1.835
+ $X2=6.72 $Y2=1.835
r78 29 31 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=6.63 $Y=1.98 $X2=6.63
+ $Y2=2.91
r79 27 41 1.34256 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=6.63 $Y=1.925 $X2=6.63
+ $Y2=1.835
r80 27 29 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=6.63 $Y=1.925
+ $X2=6.63 $Y2=1.98
r81 25 42 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=6.805 $Y=1.14 $X2=6.9
+ $Y2=1.14
r82 25 26 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=6.805 $Y=1.14
+ $X2=6.135 $Y2=1.14
r83 21 26 7.03324 $w=1.9e-07 $l=1.71026e-07 $layer=LI1_cond $X=6.005 $Y=1.045
+ $X2=6.135 $Y2=1.14
r84 21 23 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=6.005 $Y=1.045
+ $X2=6.005 $Y2=0.42
r85 19 41 5.16603 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=6.54 $Y=1.835 $X2=6.63
+ $Y2=1.835
r86 19 20 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=6.54 $Y=1.835
+ $X2=5.87 $Y2=1.835
r87 15 17 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=5.775 $Y=1.98
+ $X2=5.775 $Y2=2.91
r88 13 20 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=5.775 $Y=1.925
+ $X2=5.87 $Y2=1.835
r89 13 15 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=5.775 $Y=1.925
+ $X2=5.775 $Y2=1.98
r90 4 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.495
+ $Y=1.835 $X2=6.635 $Y2=2.91
r91 4 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.495
+ $Y=1.835 $X2=6.635 $Y2=1.98
r92 3 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.635
+ $Y=1.835 $X2=5.775 $Y2=2.91
r93 3 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.635
+ $Y=1.835 $X2=5.775 $Y2=1.98
r94 2 37 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.76
+ $Y=0.235 $X2=6.9 $Y2=0.42
r95 1 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.9
+ $Y=0.235 $X2=6.04 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%A_49_47# 1 2 3 4 15 17 18 21 27 29 30 31 39
r59 32 37 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0.345
+ $X2=2.17 $Y2=0.345
r60 31 39 3.54319 $w=1.8e-07 $l=9.7e-08 $layer=LI1_cond $X=2.93 $Y=0.345
+ $X2=3.027 $Y2=0.345
r61 31 32 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=2.93 $Y=0.345
+ $X2=2.335 $Y2=0.345
r62 29 37 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.17 $Y=0.435 $X2=2.17
+ $Y2=0.345
r63 29 30 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.17 $Y=0.435
+ $X2=2.17 $Y2=0.655
r64 28 35 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.325 $Y=0.74
+ $X2=1.23 $Y2=0.74
r65 27 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.005 $Y=0.74
+ $X2=2.17 $Y2=0.655
r66 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.005 $Y=0.74
+ $X2=1.325 $Y2=0.74
r67 24 26 8.31818 $w=1.78e-07 $l=1.35e-07 $layer=LI1_cond $X=1.225 $Y=1.065
+ $X2=1.225 $Y2=0.93
r68 23 35 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.225 $Y=0.825
+ $X2=1.23 $Y2=0.74
r69 23 26 6.4697 $w=1.78e-07 $l=1.05e-07 $layer=LI1_cond $X=1.225 $Y=0.825
+ $X2=1.225 $Y2=0.93
r70 19 35 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.655
+ $X2=1.23 $Y2=0.74
r71 19 21 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.23 $Y=0.655
+ $X2=1.23 $Y2=0.42
r72 17 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.135 $Y=1.15
+ $X2=1.225 $Y2=1.065
r73 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.135 $Y=1.15
+ $X2=0.465 $Y2=1.15
r74 13 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.335 $Y=1.065
+ $X2=0.465 $Y2=1.15
r75 13 15 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=0.335 $Y=1.065
+ $X2=0.335 $Y2=0.42
r76 4 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.89
+ $Y=0.235 $X2=3.03 $Y2=0.42
r77 3 37 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.03
+ $Y=0.235 $X2=2.17 $Y2=0.37
r78 2 26 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.93
r79 2 21 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.42
r80 1 15 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 43 45
+ 50 55 63 68 73 79 82 85 88 91 95
r120 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r121 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r122 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r123 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r124 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r125 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 77 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r127 77 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r128 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r129 74 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.635 $Y=0 $X2=6.47
+ $Y2=0
r130 74 76 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.635 $Y=0
+ $X2=6.96 $Y2=0
r131 73 94 4.59886 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=7.165 $Y=0
+ $X2=7.422 $Y2=0
r132 73 76 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.165 $Y=0
+ $X2=6.96 $Y2=0
r133 72 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r134 72 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r135 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r136 69 88 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=5.705 $Y=0 $X2=5.44
+ $Y2=0
r137 69 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.705 $Y=0 $X2=6
+ $Y2=0
r138 68 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6.47
+ $Y2=0
r139 68 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6
+ $Y2=0
r140 67 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r141 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r142 64 85 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.515
+ $Y2=0
r143 64 66 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=3.645 $Y=0
+ $X2=5.04 $Y2=0
r144 63 88 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.44
+ $Y2=0
r145 63 66 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.175 $Y=0
+ $X2=5.04 $Y2=0
r146 62 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r147 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r148 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r149 59 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r150 58 61 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r151 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r152 56 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.66
+ $Y2=0
r153 56 58 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=2.16 $Y2=0
r154 55 85 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.515
+ $Y2=0
r155 55 61 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=3.12 $Y2=0
r156 54 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r157 54 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r158 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r159 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.8
+ $Y2=0
r160 51 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.2
+ $Y2=0
r161 50 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.66
+ $Y2=0
r162 50 53 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.2
+ $Y2=0
r163 48 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r164 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r165 45 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.8
+ $Y2=0
r166 45 47 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0
+ $X2=0.24 $Y2=0
r167 43 67 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=5.04
+ $Y2=0
r168 43 86 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r169 39 94 3.16731 $w=3.3e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.33 $Y=0.085
+ $X2=7.422 $Y2=0
r170 39 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.33 $Y=0.085
+ $X2=7.33 $Y2=0.38
r171 35 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0
r172 35 37 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0.36
r173 31 88 2.222 $w=5.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=0.085 $X2=5.44
+ $Y2=0
r174 31 33 6.65742 $w=5.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.44 $Y=0.085
+ $X2=5.44 $Y2=0.38
r175 27 85 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=0.085
+ $X2=3.515 $Y2=0
r176 27 29 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=3.515 $Y=0.085
+ $X2=3.515 $Y2=0.39
r177 23 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0
r178 23 25 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0.375
r179 19 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r180 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.8 $Y=0.085
+ $X2=0.8 $Y2=0.38
r181 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.19
+ $Y=0.235 $X2=7.33 $Y2=0.38
r182 5 37 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.33
+ $Y=0.235 $X2=6.47 $Y2=0.36
r183 4 33 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=5.13
+ $Y=0.235 $X2=5.61 $Y2=0.38
r184 3 29 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=3.425
+ $Y=0.235 $X2=3.55 $Y2=0.39
r185 2 25 182 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.235 $X2=1.66 $Y2=0.375
r186 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.235 $X2=0.8 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_4%A_768_47# 1 2 7 11 13
r19 11 16 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=4.875 $Y=0.485
+ $X2=4.875 $Y2=0.37
r20 11 13 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=4.875 $Y=0.485
+ $X2=4.875 $Y2=0.75
r21 7 16 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=4.745 $Y=0.37
+ $X2=4.875 $Y2=0.37
r22 7 9 38.3313 $w=2.28e-07 $l=7.65e-07 $layer=LI1_cond $X=4.745 $Y=0.37
+ $X2=3.98 $Y2=0.37
r23 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.7
+ $Y=0.235 $X2=4.84 $Y2=0.38
r24 2 13 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=4.7
+ $Y=0.235 $X2=4.84 $Y2=0.75
r25 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.84
+ $Y=0.235 $X2=3.98 $Y2=0.38
.ends

