* File: sky130_fd_sc_lp__and2_4.spice
* Created: Wed Sep  2 09:30:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2_4.pex.spice"
.subckt sky130_fd_sc_lp__and2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_110_47# N_A_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g A_110_47# VNB NSHORT L=0.15 W=0.84 AD=0.1785
+ AS=0.0882 PD=1.265 PS=1.05 NRD=9.996 NRS=7.14 M=1 R=5.6 SA=75000.6 SB=75002.1
+ A=0.126 P=1.98 MULT=1
MM1002 N_X_M1002_d N_A_27_47#_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1785 PD=1.12 PS=1.265 NRD=0 NRS=10.704 M=1 R=5.6 SA=75001.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1002_d N_A_27_47#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1007_d N_A_27_47#_M1007_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1009 N_X_M1007_d N_A_27_47#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_A_27_47#_M1011_d N_A_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_A_27_47#_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.22365 AS=0.1764 PD=1.615 PS=1.54 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1005_d N_A_27_47#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.22365 AS=0.1764 PD=1.615 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_47#_M1006_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1006_d N_A_27_47#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_47#_M1010_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__and2_4.pxi.spice"
*
.ends
*
*
