* NGSPICE file created from sky130_fd_sc_lp__buflp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__buflp_4 A VGND VNB VPB VPWR X
M1000 VPWR a_84_21# a_114_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.2411e+12p pd=9.53e+06u as=1.5876e+12p ps=1.26e+07u
M1001 X a_84_21# a_114_47# VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=9.408e+11p ps=8.96e+06u
M1002 X a_84_21# a_114_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_84_21# a_114_47# VNB nshort w=840000u l=150000u
+  ad=1.0626e+12p pd=7.57e+06u as=0p ps=0u
M1004 a_114_47# a_84_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_886_47# A VGND VNB nshort w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=0p ps=0u
M1006 a_84_21# A a_886_47# VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1007 X a_84_21# a_114_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.82e+11p pd=6.44e+06u as=0p ps=0u
M1008 a_84_21# A a_886_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=3.024e+11p ps=3e+06u
M1009 a_114_47# a_84_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_114_367# a_84_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_114_367# a_84_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_114_367# a_84_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_84_21# a_114_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_84_21# a_114_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_114_47# a_84_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_114_47# a_84_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_114_367# a_84_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_886_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_84_21# a_114_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

