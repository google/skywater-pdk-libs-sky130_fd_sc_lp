* File: sky130_fd_sc_lp__o2111a_0.spice
* Created: Wed Sep  2 10:12:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111a_0.pex.spice"
.subckt sky130_fd_sc_lp__o2111a_0  VNB VPB D1 C1 B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_315_47# N_D1_M1001_g N_A_80_21#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 A_387_47# N_C1_M1004_g A_315_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_459_47#_M1005_d N_B1_M1005_g A_387_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_459_47#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=9.996 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_459_47#_M1009_d N_A1_M1009_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0735 PD=1.37 PS=0.77 NRD=0 NRS=9.996 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.112 AS=0.1696 PD=0.99 PS=1.81 NRD=10.7562 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1008 N_A_80_21#_M1008_d N_D1_M1008_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=10.7562 M=1 R=4.26667 SA=75000.7
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_A_80_21#_M1008_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1984 AS=0.0896 PD=1.26 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1011 N_A_80_21#_M1011_d N_B1_M1011_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1984 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1006 A_585_481# N_A2_M1006_g N_A_80_21#_M1011_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g A_585_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75002.7
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_88 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o2111a_0.pxi.spice"
*
.ends
*
*
