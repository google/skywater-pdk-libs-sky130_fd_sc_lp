# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__einvn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.425000 1.765000 1.750000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.071000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.470000 1.745000 4.725000 2.860000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.512000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.825000 0.595000 1.155000 1.075000 ;
        RECT 0.825000 1.075000 2.245000 1.245000 ;
        RECT 0.905000 1.920000 2.175000 2.090000 ;
        RECT 0.905000 2.090000 1.235000 2.735000 ;
        RECT 1.845000 0.595000 2.245000 1.075000 ;
        RECT 1.845000 2.090000 2.175000 2.735000 ;
        RECT 1.945000 1.245000 2.245000 1.500000 ;
        RECT 1.945000 1.500000 2.175000 1.920000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.375000  0.255000 2.675000 0.425000 ;
      RECT 0.375000  0.425000 0.645000 1.205000 ;
      RECT 0.395000  1.920000 0.665000 2.905000 ;
      RECT 0.395000  2.905000 2.535000 3.075000 ;
      RECT 1.335000  0.425000 1.665000 0.895000 ;
      RECT 1.405000  2.260000 1.675000 2.905000 ;
      RECT 2.345000  1.755000 4.300000 1.925000 ;
      RECT 2.345000  1.925000 2.535000 2.905000 ;
      RECT 2.415000  0.425000 2.675000 0.725000 ;
      RECT 2.415000  0.725000 3.865000 0.895000 ;
      RECT 2.415000  0.895000 2.605000 1.265000 ;
      RECT 2.705000  2.095000 3.035000 3.245000 ;
      RECT 2.775000  1.065000 3.105000 1.395000 ;
      RECT 2.775000  1.395000 5.655000 1.575000 ;
      RECT 3.175000  0.085000 3.505000 0.555000 ;
      RECT 3.205000  1.925000 3.395000 3.075000 ;
      RECT 3.565000  2.095000 3.895000 3.245000 ;
      RECT 3.605000  0.895000 3.865000 1.055000 ;
      RECT 3.605000  1.055000 4.725000 1.225000 ;
      RECT 3.675000  0.255000 3.865000 0.725000 ;
      RECT 4.035000  0.085000 4.365000 0.885000 ;
      RECT 4.065000  1.925000 4.300000 3.075000 ;
      RECT 4.535000  0.255000 4.725000 1.055000 ;
      RECT 4.895000  0.085000 5.225000 1.115000 ;
      RECT 4.895000  1.815000 5.180000 3.245000 ;
      RECT 5.350000  1.575000 5.655000 3.075000 ;
      RECT 5.395000  0.255000 5.655000 1.395000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__einvn_4
END LIBRARY
