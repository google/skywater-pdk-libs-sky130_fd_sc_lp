* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_778_399# a_733_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 VPWR SCE a_204_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_182_120# D a_268_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1102_93# a_1188_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_2008_122# a_2122_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_204_489# D a_182_120# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_182_120# a_1102_93# a_733_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 Q a_2122_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_1102_93# a_1188_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_2097_122# a_2122_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_2122_329# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND SCE a_332_94# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1060_119# a_1102_93# a_733_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_110_120# SCE a_182_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_182_120# a_332_94# a_27_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 VGND CLK a_1188_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_2008_122# a_1188_93# a_2097_122# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_2122_329# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VGND a_2122_329# a_2710_56# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_733_21# a_1188_93# a_993_425# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND SCD a_110_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_268_120# a_332_94# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VGND a_778_399# a_1060_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 Q a_2122_329# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VPWR a_2008_122# a_2122_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 VGND a_2710_56# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_733_21# a_1188_93# a_182_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_778_399# a_733_21# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 Q_N a_2710_56# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 a_27_489# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 VPWR CLK a_1188_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_2008_122# a_1102_93# a_2116_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VPWR a_2710_56# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_2116_463# a_2122_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 a_332_94# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 a_778_399# a_1188_93# a_2008_122# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X36 VPWR a_778_399# a_993_425# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 Q_N a_2710_56# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 a_778_399# a_1102_93# a_2008_122# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VPWR a_2122_329# a_2710_56# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
