* File: sky130_fd_sc_lp__srdlxtp_1.pex.spice
* Created: Fri Aug 28 11:33:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%A_84_153# 1 2 9 13 15 19 23 25 27 29 31 35
+ 36 39 40 41 44 47 50 52 53 55 58 60 61 67 73 75 79 81 90
c234 67 0 1.99017e-20 $X=2.475 $Y=1.71
c235 27 0 5.10977e-20 $X=3.84 $Y=0.445
r236 81 83 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=6.155 $Y=0.465
+ $X2=6.155 $Y2=0.59
r237 75 78 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.21 $Y=1.35
+ $X2=4.21 $Y2=1.515
r238 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.35 $X2=4.21 $Y2=1.35
r239 70 72 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=1.79
+ $X2=2.475 $Y2=1.955
r240 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.79 $X2=2.48 $Y2=1.79
r241 67 70 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.475 $Y=1.71
+ $X2=2.475 $Y2=1.79
r242 65 90 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.04 $Y=1.79 $X2=1.04
+ $Y2=1.7
r243 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.79 $X2=1.04 $Y2=1.79
r244 61 64 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.04 $Y=1.71 $X2=1.04
+ $Y2=1.79
r245 58 86 3.09537 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=6.705 $Y=2.075
+ $X2=6.705 $Y2=2.205
r246 58 60 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.705 $Y=2.075
+ $X2=6.705 $Y2=1.82
r247 57 60 52.7819 $w=2.48e-07 $l=1.145e-06 $layer=LI1_cond $X=6.705 $Y=0.675
+ $X2=6.705 $Y2=1.82
r248 56 83 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=0.59
+ $X2=6.155 $Y2=0.59
r249 55 57 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.58 $Y=0.59
+ $X2=6.705 $Y2=0.675
r250 55 56 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.58 $Y=0.59
+ $X2=6.32 $Y2=0.59
r251 54 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=2.16
+ $X2=4.29 $Y2=2.16
r252 53 86 4.04779 $w=1.7e-07 $l=1.45774e-07 $layer=LI1_cond $X=6.58 $Y=2.16
+ $X2=6.705 $Y2=2.205
r253 53 54 143.856 $w=1.68e-07 $l=2.205e-06 $layer=LI1_cond $X=6.58 $Y=2.16
+ $X2=4.375 $Y2=2.16
r254 51 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=2.245
+ $X2=4.29 $Y2=2.16
r255 51 52 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.29 $Y=2.245
+ $X2=4.29 $Y2=2.905
r256 50 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=2.075
+ $X2=4.29 $Y2=2.16
r257 50 78 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.29 $Y=2.075
+ $X2=4.29 $Y2=1.515
r258 48 73 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=3.475 $Y=2.99
+ $X2=3.312 $Y2=2.99
r259 47 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.205 $Y=2.99
+ $X2=4.29 $Y2=2.905
r260 47 48 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.205 $Y=2.99
+ $X2=3.475 $Y2=2.99
r261 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.31
+ $Y=2.13 $X2=3.31 $Y2=2.13
r262 42 73 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.312 $Y=2.905
+ $X2=3.312 $Y2=2.99
r263 42 44 27.4813 $w=3.23e-07 $l=7.75e-07 $layer=LI1_cond $X=3.312 $Y=2.905
+ $X2=3.312 $Y2=2.13
r264 40 73 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=3.15 $Y=2.99
+ $X2=3.312 $Y2=2.99
r265 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.15 $Y=2.99
+ $X2=2.48 $Y2=2.99
r266 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.395 $Y=2.905
+ $X2=2.48 $Y2=2.99
r267 39 72 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.395 $Y=2.905
+ $X2=2.395 $Y2=1.955
r268 37 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=1.71
+ $X2=1.04 $Y2=1.71
r269 36 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=1.71
+ $X2=2.475 $Y2=1.71
r270 36 37 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.31 $Y=1.71
+ $X2=1.205 $Y2=1.71
r271 35 45 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.45 $Y=2.13
+ $X2=3.31 $Y2=2.13
r272 34 45 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.105 $Y=2.13
+ $X2=3.31 $Y2=2.13
r273 31 71 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=2.955 $Y=1.79
+ $X2=2.48 $Y2=1.79
r274 31 34 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.03 $Y=1.79
+ $X2=3.03 $Y2=2.13
r275 25 76 72.2024 $w=2.47e-07 $l=4.44916e-07 $layer=POLY_cond $X=3.84 $Y=1.185
+ $X2=4.21 $Y2=1.35
r276 25 27 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.84 $Y=1.185
+ $X2=3.84 $Y2=0.445
r277 21 35 26.8146 $w=2.88e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.525 $Y=2.295
+ $X2=3.45 $Y2=2.13
r278 21 23 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.525 $Y=2.295
+ $X2=3.525 $Y2=2.775
r279 17 34 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.03 $Y=2.295
+ $X2=3.03 $Y2=2.13
r280 17 19 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.03 $Y=2.295
+ $X2=3.03 $Y2=2.775
r281 16 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=1.7
+ $X2=0.495 $Y2=1.7
r282 15 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.875 $Y=1.7
+ $X2=1.04 $Y2=1.7
r283 15 16 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=0.875 $Y=1.7
+ $X2=0.57 $Y2=1.7
r284 11 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.775
+ $X2=0.495 $Y2=1.7
r285 11 13 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=0.495 $Y=1.775
+ $X2=0.495 $Y2=2.735
r286 7 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.625
+ $X2=0.495 $Y2=1.7
r287 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.495 $Y=1.625
+ $X2=0.495 $Y2=1.105
r288 2 86 600 $w=1.7e-07 $l=6.19375e-07 $layer=licon1_PDIFF $count=1 $X=6.385
+ $Y=1.675 $X2=6.665 $Y2=2.17
r289 2 60 600 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=6.385
+ $Y=1.675 $X2=6.665 $Y2=1.82
r290 1 81 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=6.01
+ $Y=0.235 $X2=6.155 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%D 3 7 9 10 11
r47 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=0.95 $X2=1.15 $Y2=0.95
r48 9 14 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.415 $Y=0.95
+ $X2=1.15 $Y2=0.95
r49 9 10 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=0.95
+ $X2=1.415 $Y2=0.785
r50 5 10 37.0704 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=1.545 $Y=0.785
+ $X2=1.415 $Y2=0.785
r51 5 7 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.545 $Y=0.785
+ $X2=1.545 $Y2=0.445
r52 1 10 37.0704 $w=1.5e-07 $l=3.65582e-07 $layer=POLY_cond $X=1.49 $Y=1.115
+ $X2=1.415 $Y2=0.785
r53 1 3 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=1.49 $Y=1.115
+ $X2=1.49 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%A_226_491# 1 2 9 11 13 14 16 19 21 22 23
+ 27 28 31 33 37 40
c104 37 0 1.69905e-19 $X=2.025 $Y=0.93
c105 33 0 1.69905e-19 $X=2.025 $Y=0.7
c106 11 0 1.85752e-20 $X=2.305 $Y=0.765
r107 37 43 16.4318 $w=2.64e-07 $l=9e-08 $layer=POLY_cond $X=2.025 $Y=0.93
+ $X2=1.935 $Y2=0.93
r108 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.025
+ $Y=0.93 $X2=2.025 $Y2=0.93
r109 33 36 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.025 $Y=0.7
+ $X2=2.025 $Y2=0.93
r110 28 41 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.94 $Y=2.13
+ $X2=1.94 $Y2=2.27
r111 28 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.94 $Y=2.13
+ $X2=1.94 $Y2=1.965
r112 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.13 $X2=1.94 $Y2=2.13
r113 25 27 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.94 $Y=2.435
+ $X2=1.94 $Y2=2.13
r114 24 31 8.354 $w=3.87e-07 $l=3.67628e-07 $layer=LI1_cond $X=1.655 $Y=0.7
+ $X2=1.41 $Y2=0.435
r115 23 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0.7
+ $X2=2.025 $Y2=0.7
r116 23 24 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.86 $Y=0.7
+ $X2=1.655 $Y2=0.7
r117 21 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.775 $Y=2.52
+ $X2=1.94 $Y2=2.435
r118 21 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.775 $Y=2.52
+ $X2=1.44 $Y2=2.52
r119 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.275 $Y=2.605
+ $X2=1.44 $Y2=2.52
r120 17 19 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.275 $Y=2.605
+ $X2=1.275 $Y2=2.755
r121 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.6 $Y=2.345
+ $X2=2.6 $Y2=2.775
r122 11 37 51.1212 $w=2.64e-07 $l=3.52987e-07 $layer=POLY_cond $X=2.305 $Y=0.765
+ $X2=2.025 $Y2=0.93
r123 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.305 $Y=0.765
+ $X2=2.305 $Y2=0.445
r124 10 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.105 $Y=2.27
+ $X2=1.94 $Y2=2.27
r125 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.525 $Y=2.27
+ $X2=2.6 $Y2=2.345
r126 9 10 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.525 $Y=2.27
+ $X2=2.105 $Y2=2.27
r127 7 43 15.9823 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.095
+ $X2=1.935 $Y2=0.93
r128 7 40 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.935 $Y=1.095
+ $X2=1.935 $Y2=1.965
r129 2 19 600 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=2.455 $X2=1.275 $Y2=2.755
r130 1 31 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.235 $X2=1.33 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%A_114_179# 1 2 9 11 15 18 19 20 21 25 28
+ 30 36 42 44 46 47 49 50
c131 50 0 1.89807e-19 $X=2.785 $Y=1.22
c132 49 0 1.69905e-19 $X=2.785 $Y=1.22
c133 21 0 1.59492e-19 $X=3.995 $Y=1.8
c134 15 0 6.47033e-20 $X=3.235 $Y=0.445
r135 50 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.785 $Y=1.22
+ $X2=2.785 $Y2=1.31
r136 50 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.22
+ $X2=2.785 $Y2=1.055
r137 49 52 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.785 $Y=1.22
+ $X2=2.785 $Y2=1.37
r138 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=1.22 $X2=2.785 $Y2=1.22
r139 46 47 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=2.56
+ $X2=0.705 $Y2=2.395
r140 43 44 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.795 $Y=1.37
+ $X2=0.665 $Y2=1.37
r141 42 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=1.37
+ $X2=2.785 $Y2=1.37
r142 42 43 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=2.62 $Y=1.37
+ $X2=0.795 $Y2=1.37
r143 38 44 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.62 $Y=1.455
+ $X2=0.665 $Y2=1.37
r144 38 47 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.62 $Y=1.455
+ $X2=0.62 $Y2=2.395
r145 34 44 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=1.285
+ $X2=0.665 $Y2=1.37
r146 34 36 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.665 $Y=1.285
+ $X2=0.665 $Y2=1.105
r147 30 32 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.76 $Y=1.65
+ $X2=3.76 $Y2=1.8
r148 27 28 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=3.235 $Y=1.31
+ $X2=3.42 $Y2=1.31
r149 23 25 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=4.12 $Y=1.875
+ $X2=4.12 $Y2=2.595
r150 22 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=1.8
+ $X2=3.76 $Y2=1.8
r151 21 23 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.995 $Y=1.8
+ $X2=4.12 $Y2=1.875
r152 21 22 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=3.995 $Y=1.8
+ $X2=3.835 $Y2=1.8
r153 19 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.685 $Y=1.65
+ $X2=3.76 $Y2=1.65
r154 19 20 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.685 $Y=1.65
+ $X2=3.495 $Y2=1.65
r155 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.42 $Y=1.575
+ $X2=3.495 $Y2=1.65
r156 17 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.42 $Y=1.385
+ $X2=3.42 $Y2=1.31
r157 17 18 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.42 $Y=1.385
+ $X2=3.42 $Y2=1.575
r158 13 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.235 $Y=1.235
+ $X2=3.235 $Y2=1.31
r159 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.235 $Y=1.235
+ $X2=3.235 $Y2=0.445
r160 12 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.31
+ $X2=2.785 $Y2=1.31
r161 11 27 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.16 $Y=1.31
+ $X2=3.235 $Y2=1.31
r162 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.16 $Y=1.31
+ $X2=2.95 $Y2=1.31
r163 9 55 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.875 $Y=0.445
+ $X2=2.875 $Y2=1.055
r164 2 46 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.415 $X2=0.71 $Y2=2.56
r165 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.895 $X2=0.71 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%A_831_21# 1 2 9 11 12 15 19 22 23 24 30 32
+ 38
c77 24 0 1.59492e-19 $X=5.445 $Y=1.74
c78 23 0 1.05754e-19 $X=4.625 $Y=0.87
c79 15 0 2.50468e-19 $X=4.61 $Y=2.595
r80 37 38 8.36806 $w=2.88e-07 $l=5e-08 $layer=POLY_cond $X=4.61 $Y=1.74 $X2=4.66
+ $Y2=1.74
r81 32 34 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.595 $Y=0.465
+ $X2=5.595 $Y2=0.675
r82 30 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=1.575
+ $X2=5.53 $Y2=1.74
r83 30 34 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.53 $Y=1.575 $X2=5.53
+ $Y2=0.675
r84 27 38 15.0625 $w=2.88e-07 $l=9e-08 $layer=POLY_cond $X=4.75 $Y=1.74 $X2=4.66
+ $Y2=1.74
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.75
+ $Y=1.74 $X2=4.75 $Y2=1.74
r86 24 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=1.74 $X2=5.53
+ $Y2=1.74
r87 24 26 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.445 $Y=1.74
+ $X2=4.75 $Y2=1.74
r88 22 38 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.575
+ $X2=4.66 $Y2=1.74
r89 21 23 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=4.66 $Y=0.945
+ $X2=4.625 $Y2=0.87
r90 21 22 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.66 $Y=0.945
+ $X2=4.66 $Y2=1.575
r91 17 23 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=4.59 $Y=0.795
+ $X2=4.625 $Y2=0.87
r92 17 19 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.59 $Y=0.795
+ $X2=4.59 $Y2=0.445
r93 13 37 6.18571 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.61 $Y=1.905
+ $X2=4.61 $Y2=1.74
r94 13 15 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.61 $Y=1.905
+ $X2=4.61 $Y2=2.595
r95 11 23 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=4.515 $Y=0.87
+ $X2=4.625 $Y2=0.87
r96 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.515 $Y=0.87
+ $X2=4.305 $Y2=0.87
r97 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.23 $Y=0.795
+ $X2=4.305 $Y2=0.87
r98 7 9 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.23 $Y=0.795 $X2=4.23
+ $Y2=0.445
r99 2 36 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.305
+ $Y=1.675 $X2=5.45 $Y2=1.82
r100 1 32 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=5.455
+ $Y=0.235 $X2=5.595 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%GATE 2 5 9 11 12 13 17 18
r42 17 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.262 $Y=1.01
+ $X2=6.262 $Y2=0.845
r43 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.245
+ $Y=1.01 $X2=6.245 $Y2=1.01
r44 12 13 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=6.147 $Y=1.295
+ $X2=6.147 $Y2=1.665
r45 12 18 6.493 $w=5.23e-07 $l=2.85e-07 $layer=LI1_cond $X=6.147 $Y=1.295
+ $X2=6.147 $Y2=1.01
r46 9 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.37 $Y=0.445 $X2=6.37
+ $Y2=0.845
r47 5 11 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.31 $Y=1.995
+ $X2=6.31 $Y2=1.515
r48 2 11 42.0615 $w=3.65e-07 $l=1.82e-07 $layer=POLY_cond $X=6.262 $Y=1.333
+ $X2=6.262 $Y2=1.515
r49 1 17 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=6.262 $Y=1.027
+ $X2=6.262 $Y2=1.01
r50 1 2 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=6.262 $Y=1.027
+ $X2=6.262 $Y2=1.333
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%SLEEP_B 3 7 9 11 12 13 18
r46 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.18
+ $Y=0.94 $X2=7.18 $Y2=0.94
r47 18 20 18.3814 $w=2.36e-07 $l=9e-08 $layer=POLY_cond $X=7.09 $Y=0.955
+ $X2=7.18 $Y2=0.955
r48 17 18 42.8898 $w=2.36e-07 $l=2.1e-07 $layer=POLY_cond $X=6.88 $Y=0.955
+ $X2=7.09 $Y2=0.955
r49 13 21 7.86311 $w=5.38e-07 $l=3.55e-07 $layer=LI1_cond $X=7.285 $Y=1.295
+ $X2=7.285 $Y2=0.94
r50 12 21 0.332244 $w=5.38e-07 $l=1.5e-08 $layer=LI1_cond $X=7.285 $Y=0.925
+ $X2=7.285 $Y2=0.94
r51 9 18 13.389 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.09 $Y=0.775 $X2=7.09
+ $Y2=0.955
r52 9 11 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=7.09 $Y=0.775 $X2=7.09
+ $Y2=0.445
r53 5 17 13.389 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.88 $Y=1.105 $X2=6.88
+ $Y2=0.955
r54 5 7 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=6.88 $Y=1.105 $X2=6.88
+ $Y2=1.995
r55 1 17 30.6356 $w=2.36e-07 $l=1.5e-07 $layer=POLY_cond $X=6.73 $Y=0.955
+ $X2=6.88 $Y2=0.955
r56 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.73 $Y=0.955 $X2=6.73
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%A_662_47# 1 2 9 13 18 19 20 22 23 26 27 28
+ 31 35 39 41 44 48 50 52 54 55 56 64
c159 56 0 1.05754e-19 $X=5.11 $Y=0.93
c160 50 0 1.51059e-19 $X=3.855 $Y=2.405
c161 48 0 9.9409e-20 $X=3.855 $Y=2.24
c162 18 0 6.66559e-20 $X=5.715 $Y=2.175
r163 60 64 51.6429 $w=2.52e-07 $l=2.7e-07 $layer=POLY_cond $X=5.11 $Y=1.01
+ $X2=5.38 $Y2=1.01
r164 60 62 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=5.11 $Y=1.01
+ $X2=5.02 $Y2=1.01
r165 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.11
+ $Y=1.01 $X2=5.11 $Y2=1.01
r166 56 59 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.11 $Y=0.93 $X2=5.11
+ $Y2=1.01
r167 53 54 2.76166 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.86 $Y=0.93 $X2=3.66
+ $Y2=0.93
r168 52 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.945 $Y=0.93
+ $X2=5.11 $Y2=0.93
r169 52 53 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=4.945 $Y=0.93
+ $X2=3.86 $Y2=0.93
r170 48 55 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.24
+ $X2=3.855 $Y2=2.075
r171 48 50 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.24
+ $X2=3.855 $Y2=2.405
r172 46 54 3.70735 $w=2.5e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.775 $Y=1.015
+ $X2=3.66 $Y2=0.93
r173 46 55 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.775 $Y=1.015
+ $X2=3.775 $Y2=2.075
r174 42 54 3.70735 $w=2.5e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.625 $Y=0.845
+ $X2=3.66 $Y2=0.93
r175 42 44 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=3.625 $Y=0.845
+ $X2=3.625 $Y2=0.465
r176 37 39 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.5 $Y=1.42
+ $X2=7.66 $Y2=1.42
r177 33 35 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.08 $Y=0.925
+ $X2=8.08 $Y2=0.485
r178 29 31 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=8.01 $Y=2.785
+ $X2=8.01 $Y2=2.155
r179 27 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.005 $Y=1
+ $X2=8.08 $Y2=0.925
r180 27 28 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.005 $Y=1
+ $X2=7.735 $Y2=1
r181 26 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.66 $Y=1.345
+ $X2=7.66 $Y2=1.42
r182 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.66 $Y=1.075
+ $X2=7.735 $Y2=1
r183 25 26 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.66 $Y=1.075
+ $X2=7.66 $Y2=1.345
r184 24 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.575 $Y=2.86
+ $X2=7.5 $Y2=2.86
r185 23 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.935 $Y=2.86
+ $X2=8.01 $Y2=2.785
r186 23 24 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.935 $Y=2.86
+ $X2=7.575 $Y2=2.86
r187 22 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.5 $Y=2.785
+ $X2=7.5 $Y2=2.86
r188 21 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.5 $Y=1.495
+ $X2=7.5 $Y2=1.42
r189 21 22 661.468 $w=1.5e-07 $l=1.29e-06 $layer=POLY_cond $X=7.5 $Y=1.495
+ $X2=7.5 $Y2=2.785
r190 19 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.425 $Y=2.86
+ $X2=7.5 $Y2=2.86
r191 19 20 812.734 $w=1.5e-07 $l=1.585e-06 $layer=POLY_cond $X=7.425 $Y=2.86
+ $X2=5.84 $Y2=2.86
r192 16 20 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=5.715 $Y=2.785
+ $X2=5.84 $Y2=2.86
r193 16 18 151.557 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.715 $Y=2.785
+ $X2=5.715 $Y2=2.175
r194 15 64 64.0754 $w=2.52e-07 $l=4.09268e-07 $layer=POLY_cond $X=5.715 $Y=1.175
+ $X2=5.38 $Y2=1.01
r195 15 18 248.454 $w=2.5e-07 $l=1e-06 $layer=POLY_cond $X=5.715 $Y=1.175
+ $X2=5.715 $Y2=2.175
r196 11 64 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=0.845
+ $X2=5.38 $Y2=1.01
r197 11 13 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.38 $Y=0.845
+ $X2=5.38 $Y2=0.445
r198 7 62 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.02 $Y=0.845
+ $X2=5.02 $Y2=1.01
r199 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.02 $Y=0.845 $X2=5.02
+ $Y2=0.445
r200 2 50 600 $w=1.7e-07 $l=2.78882e-07 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=2.455 $X2=3.855 $Y2=2.405
r201 1 44 182 $w=1.7e-07 $l=4.14337e-07 $layer=licon1_NDIFF $count=1 $X=3.31
+ $Y=0.235 $X2=3.625 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%A_1530_367# 1 2 9 13 17 20 25 26 28 30 33
r59 30 32 6.98917 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.865 $Y=0.43
+ $X2=7.865 $Y2=0.605
r60 26 36 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.517 $Y=1.48
+ $X2=8.517 $Y2=1.645
r61 26 35 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.517 $Y=1.48
+ $X2=8.517 $Y2=1.315
r62 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.5
+ $Y=1.48 $X2=8.5 $Y2=1.48
r63 23 33 0.30096 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=8.03 $Y=1.48 $X2=7.91
+ $Y2=1.48
r64 23 25 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=8.03 $Y=1.48 $X2=8.5
+ $Y2=1.48
r65 21 33 7.52254 $w=2.05e-07 $l=1.81659e-07 $layer=LI1_cond $X=7.875 $Y=1.645
+ $X2=7.91 $Y2=1.48
r66 21 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.875 $Y=1.645
+ $X2=7.875 $Y2=1.815
r67 20 33 7.52254 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=7.91 $Y=1.315
+ $X2=7.91 $Y2=1.48
r68 20 32 34.0931 $w=2.38e-07 $l=7.1e-07 $layer=LI1_cond $X=7.91 $Y=1.315
+ $X2=7.91 $Y2=0.605
r69 17 28 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=1.98
+ $X2=7.795 $Y2=1.815
r70 13 36 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.625 $Y=2.465
+ $X2=8.625 $Y2=1.645
r71 9 35 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.625 $Y=0.695
+ $X2=8.625 $Y2=1.315
r72 2 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.65
+ $Y=1.835 $X2=7.795 $Y2=1.98
r73 1 30 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=7.72
+ $Y=0.275 $X2=7.865 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%VPWR 1 2 3 10 12 16 20 24 26 31 41 42 48
+ 51
r89 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r90 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r93 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r94 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.34 $Y2=3.33
r95 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.88 $Y2=3.33
r96 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r97 37 38 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r98 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 34 37 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=7.92 $Y2=3.33
r100 34 35 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.775 $Y2=3.33
r102 32 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 31 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.175 $Y=3.33
+ $X2=8.34 $Y2=3.33
r104 31 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.175 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 30 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r107 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 27 45 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r109 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.775 $Y2=3.33
r111 26 29 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 24 38 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 24 35 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=2.16 $Y2=3.33
r114 20 23 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=8.34 $Y=1.98
+ $X2=8.34 $Y2=2.465
r115 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.34 $Y=3.245
+ $X2=8.34 $Y2=3.33
r116 18 23 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=8.34 $Y=3.245
+ $X2=8.34 $Y2=2.465
r117 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.33
r118 14 16 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=2.945
r119 10 45 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r120 10 12 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.56
r121 3 23 300 $w=1.7e-07 $l=7.46693e-07 $layer=licon1_PDIFF $count=2 $X=8.085
+ $Y=1.835 $X2=8.34 $Y2=2.465
r122 3 20 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=8.085
+ $Y=1.835 $X2=8.34 $Y2=1.98
r123 2 16 600 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=2.455 $X2=1.775 $Y2=2.945
r124 1 12 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.415 $X2=0.28 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%A_476_47# 1 2 7 12 14 19 20 24
c61 14 0 6.47033e-20 $X=2.525 $Y=0.465
c62 7 0 6.96729e-20 $X=3.12 $Y=0.59
r63 22 24 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.895 $Y=1.71
+ $X2=3.205 $Y2=1.71
r64 19 20 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.61
+ $X2=2.815 $Y2=2.445
r65 14 16 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.525 $Y=0.465
+ $X2=2.525 $Y2=0.59
r66 12 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=1.625
+ $X2=3.205 $Y2=1.71
r67 11 12 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.205 $Y=0.675
+ $X2=3.205 $Y2=1.625
r68 9 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=1.795
+ $X2=2.895 $Y2=1.71
r69 9 20 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.895 $Y=1.795
+ $X2=2.895 $Y2=2.445
r70 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0.59
+ $X2=2.525 $Y2=0.59
r71 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.12 $Y=0.59
+ $X2=3.205 $Y2=0.675
r72 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=0.59 $X2=2.69
+ $Y2=0.59
r73 2 19 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=2.455 $X2=2.815 $Y2=2.61
r74 1 14 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.525 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%KAPWR 1 2 3 10 12 16 19 24 30 31
c94 12 0 6.66559e-20 $X=7 $Y=2.61
r95 27 31 12.631 $w=6.58e-07 $l=2.8e-07 $layer=LI1_cond $X=4.875 $Y=2.745
+ $X2=5.155 $Y2=2.745
r96 27 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.82
+ $X2=5.04 $Y2=2.82
r97 24 30 0.262345 $w=2.7e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=2.81
+ $X2=5.04 $Y2=2.81
r98 21 22 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.98 $Y=2.61
+ $X2=5.98 $Y2=2.805
r99 19 21 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.98 $Y=2.515
+ $X2=5.98 $Y2=2.61
r100 14 16 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=7.165 $Y=2.525
+ $X2=7.165 $Y2=1.82
r101 13 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=2.61
+ $X2=5.98 $Y2=2.61
r102 12 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7 $Y=2.61
+ $X2=7.165 $Y2=2.525
r103 12 13 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=7 $Y=2.61
+ $X2=6.145 $Y2=2.61
r104 10 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=2.805
+ $X2=5.98 $Y2=2.805
r105 10 31 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.815 $Y=2.805
+ $X2=5.155 $Y2=2.805
r106 3 16 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=6.955
+ $Y=1.675 $X2=7.165 $Y2=1.82
r107 2 19 600 $w=1.7e-07 $l=9.07304e-07 $layer=licon1_PDIFF $count=1 $X=5.84
+ $Y=1.675 $X2=5.98 $Y2=2.515
r108 1 27 600 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=1 $X=4.735
+ $Y=2.095 $X2=4.875 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%Q 1 2 9 11 15 16 17 23 29
r20 21 29 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.84 $Y=0.97
+ $X2=8.84 $Y2=0.925
r21 17 31 7.76373 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.84 $Y=0.99
+ $X2=8.84 $Y2=1.135
r22 17 21 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=8.84 $Y=0.99 $X2=8.84
+ $Y2=0.97
r23 17 29 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=8.84 $Y=0.905 $X2=8.84
+ $Y2=0.925
r24 16 17 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.84 $Y=0.555
+ $X2=8.84 $Y2=0.905
r25 16 23 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.84 $Y=0.555
+ $X2=8.84 $Y2=0.42
r26 15 31 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.92 $Y=1.815
+ $X2=8.92 $Y2=1.135
r27 9 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.84 $Y=1.98
+ $X2=8.84 $Y2=1.815
r28 9 11 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=8.84 $Y=1.98 $X2=8.84
+ $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.835 $X2=8.84 $Y2=2.91
r30 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.835 $X2=8.84 $Y2=1.98
r31 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.275 $X2=8.84 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLXTP_1%VGND 1 2 3 4 5 16 18 22 26 30 34 39 40 42
+ 43 45 46 47 68 74 75 81
r121 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r122 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 75 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r124 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r125 72 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.495 $Y=0 $X2=8.37
+ $Y2=0
r126 72 74 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.495 $Y=0
+ $X2=8.88 $Y2=0
r127 71 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r128 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r129 68 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=8.37
+ $Y2=0
r130 68 70 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.245 $Y=0
+ $X2=7.92 $Y2=0
r131 67 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r132 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r133 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r134 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r135 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r136 57 60 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r137 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r138 55 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r139 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r140 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r141 52 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r142 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r143 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r144 49 78 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r145 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r146 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r147 47 58 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=2.16
+ $Y2=0
r148 47 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r149 45 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=6.96
+ $Y2=0
r150 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=7.305
+ $Y2=0
r151 44 70 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=7.92
+ $Y2=0
r152 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=7.305
+ $Y2=0
r153 42 60 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.56
+ $Y2=0
r154 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.805
+ $Y2=0
r155 41 63 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.97 $Y=0 $X2=5.04
+ $Y2=0
r156 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=0 $X2=4.805
+ $Y2=0
r157 39 54 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=1.68 $Y2=0
r158 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.99
+ $Y2=0
r159 38 57 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.155 $Y=0 $X2=2.16
+ $Y2=0
r160 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=1.99
+ $Y2=0
r161 34 36 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=8.37 $Y=0.42
+ $X2=8.37 $Y2=0.97
r162 32 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0
r163 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0.42
r164 28 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0
r165 28 30 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0.41
r166 24 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.805 $Y=0.085
+ $X2=4.805 $Y2=0
r167 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.805 $Y=0.085
+ $X2=4.805 $Y2=0.445
r168 20 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0
r169 20 22 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0.28
r170 16 78 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r171 16 18 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=1.105
r172 5 36 182 $w=1.7e-07 $l=8.12558e-07 $layer=licon1_NDIFF $count=1 $X=8.155
+ $Y=0.275 $X2=8.41 $Y2=0.97
r173 5 34 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=8.155
+ $Y=0.275 $X2=8.41 $Y2=0.42
r174 4 30 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=7.165
+ $Y=0.235 $X2=7.305 $Y2=0.41
r175 3 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.665
+ $Y=0.235 $X2=4.805 $Y2=0.445
r176 2 22 182 $w=1.7e-07 $l=3.91855e-07 $layer=licon1_NDIFF $count=1 $X=1.62
+ $Y=0.235 $X2=1.99 $Y2=0.28
r177 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.895 $X2=0.28 $Y2=1.105
.ends

