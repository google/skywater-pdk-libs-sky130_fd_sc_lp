* File: sky130_fd_sc_lp__o22ai_m.pex.spice
* Created: Wed Sep  2 10:21:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22AI_M%B1 2 3 4 5 6 7 9 12 16 17 18 19 20 21 22 30
r43 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.105 $X2=0.27 $Y2=1.105
r44 21 22 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.405
+ $X2=0.255 $Y2=2.775
r45 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r46 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r47 18 19 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r48 18 31 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.105
r49 17 31 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.105
r50 15 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.445
+ $X2=0.27 $Y2=1.105
r51 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.445
+ $X2=0.27 $Y2=1.61
r52 14 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.09
+ $X2=0.27 $Y2=1.105
r53 10 12 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.915 $Y=2.39
+ $X2=0.915 $Y2=2.885
r54 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.845 $Y=0.94
+ $X2=0.845 $Y2=0.62
r55 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.84 $Y=2.315
+ $X2=0.915 $Y2=2.39
r56 5 6 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.84 $Y=2.315
+ $X2=0.435 $Y2=2.315
r57 4 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=1.015
+ $X2=0.27 $Y2=1.09
r58 3 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.77 $Y=1.015
+ $X2=0.845 $Y2=0.94
r59 3 4 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.77 $Y=1.015
+ $X2=0.435 $Y2=1.015
r60 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.36 $Y=2.24
+ $X2=0.435 $Y2=2.315
r61 2 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.24 $X2=0.36
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_M%B2 3 7 11 12 13 14 15 20
c43 3 0 1.60235e-19 $X=1.275 $Y=0.62
r44 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.185
+ $Y=1.495 $X2=1.185 $Y2=1.495
r45 14 15 22.1818 $w=1.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.192 $Y=1.665
+ $X2=1.192 $Y2=2.035
r46 14 21 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=1.192 $Y=1.665
+ $X2=1.192 $Y2=1.495
r47 13 21 11.9902 $w=1.83e-07 $l=2e-07 $layer=LI1_cond $X=1.192 $Y=1.295
+ $X2=1.192 $Y2=1.495
r48 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.185 $Y=1.835
+ $X2=1.185 $Y2=1.495
r49 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.835
+ $X2=1.185 $Y2=2
r50 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.33
+ $X2=1.185 $Y2=1.495
r51 7 12 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=1.275 $Y=2.885
+ $X2=1.275 $Y2=2
r52 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.275 $Y=0.62
+ $X2=1.275 $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_M%A2 3 7 11 12 13 14 15 20
r46 14 15 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.665
+ $X2=1.717 $Y2=2.035
r47 13 14 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.295
+ $X2=1.717 $Y2=1.665
r48 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.755
+ $Y=1.375 $X2=1.755 $Y2=1.375
r49 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.755 $Y=1.715
+ $X2=1.755 $Y2=1.375
r50 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.715
+ $X2=1.755 $Y2=1.88
r51 10 20 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.21
+ $X2=1.755 $Y2=1.375
r52 7 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.785 $Y=0.62
+ $X2=1.785 $Y2=1.21
r53 3 12 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.705 $Y=2.885
+ $X2=1.705 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_M%A1 3 7 12 16 17 18 19 25
r31 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.325
+ $Y=1.765 $X2=2.325 $Y2=1.765
r32 18 19 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.242 $Y=2.035
+ $X2=2.242 $Y2=2.405
r33 18 26 9.28835 $w=3.33e-07 $l=2.7e-07 $layer=LI1_cond $X=2.242 $Y=2.035
+ $X2=2.242 $Y2=1.765
r34 17 26 3.44013 $w=3.33e-07 $l=1e-07 $layer=LI1_cond $X=2.242 $Y=1.665
+ $X2=2.242 $Y2=1.765
r35 16 17 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.242 $Y=1.295
+ $X2=2.242 $Y2=1.665
r36 15 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.6
+ $X2=2.325 $Y2=1.765
r37 12 25 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.325 $Y=2.12
+ $X2=2.325 $Y2=1.765
r38 9 12 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.065 $Y=2.195
+ $X2=2.325 $Y2=2.195
r39 7 15 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.235 $Y=0.62
+ $X2=2.235 $Y2=1.6
r40 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.065 $Y=2.27
+ $X2=2.065 $Y2=2.195
r41 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.065 $Y=2.27
+ $X2=2.065 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_M%VPWR 1 2 9 13 15 17 22 29 30 33 36
r40 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.28 $Y2=3.33
r45 27 29 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=0.7 $Y2=3.33
r49 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.28 $Y2=3.33
r51 22 25 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.7 $Y2=3.33
r55 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=3.33
r59 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=2.95
r60 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=3.33
r61 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=2.95
r62 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=2.675 $X2=2.28 $Y2=2.95
r63 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.675 $X2=0.7 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_M%Y 1 2 7 8 9 11 16 17 18
r55 17 18 9.06605 $w=3.38e-07 $l=2.25e-07 $layer=LI1_cond $X=1.2 $Y=2.715
+ $X2=1.2 $Y2=2.49
r56 16 18 8.04919 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=0.92 $Y=2.405
+ $X2=1.115 $Y2=2.405
r57 9 17 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.285 $Y=2.82
+ $X2=1.2 $Y2=2.715
r58 9 11 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=1.285 $Y=2.82
+ $X2=1.49 $Y2=2.82
r59 8 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.835 $Y=2.32
+ $X2=0.92 $Y2=2.405
r60 7 15 8.52485 $w=3.22e-07 $l=3.07409e-07 $layer=LI1_cond $X=0.835 $Y=1.01
+ $X2=1.06 $Y2=0.815
r61 7 8 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=0.835 $Y=1.01
+ $X2=0.835 $Y2=2.32
r62 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.35
+ $Y=2.675 $X2=1.49 $Y2=2.82
r63 1 15 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=0.92
+ $Y=0.41 $X2=1.06 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_M%A_85_82# 1 2 3 10 15 16 17 20 22
c35 15 0 1.54761e-19 $X=1.57 $Y=0.555
r36 22 25 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.55 $Y=0.355 $X2=0.55
+ $Y2=0.555
r37 18 20 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.46 $Y=0.84
+ $X2=2.46 $Y2=0.685
r38 16 18 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.365 $Y=0.925
+ $X2=2.46 $Y2=0.84
r39 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.365 $Y=0.925
+ $X2=1.675 $Y2=0.925
r40 13 17 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.57 $Y=0.84
+ $X2=1.675 $Y2=0.925
r41 13 15 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=1.57 $Y=0.84
+ $X2=1.57 $Y2=0.555
r42 12 15 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.57 $Y=0.44
+ $X2=1.57 $Y2=0.555
r43 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=0.355
+ $X2=0.55 $Y2=0.355
r44 10 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.465 $Y=0.355
+ $X2=1.57 $Y2=0.44
r45 10 11 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.465 $Y=0.355
+ $X2=0.715 $Y2=0.355
r46 3 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.41 $X2=2.45 $Y2=0.685
r47 2 15 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.35
+ $Y=0.41 $X2=1.57 $Y2=0.555
r48 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.425
+ $Y=0.41 $X2=0.55 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_M%VGND 1 6 9 10 11 21 22
c23 6 0 1.60235e-19 $X=2.02 $Y=0.555
r24 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r25 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r26 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r27 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r28 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r30 11 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.24
+ $Y2=0
r31 9 18 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.68
+ $Y2=0
r32 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.02
+ $Y2=0
r33 8 21 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.64
+ $Y2=0
r34 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.02
+ $Y2=0
r35 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085 $X2=2.02
+ $Y2=0
r36 4 6 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.02 $Y=0.085 $X2=2.02
+ $Y2=0.555
r37 1 6 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.41 $X2=2.02 $Y2=0.555
.ends

