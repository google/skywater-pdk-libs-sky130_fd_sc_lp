# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.840000 1.365000 1.760000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.150000 1.850000 7.595000 3.075000 ;
        RECT 7.325000 0.255000 7.595000 1.850000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.465000 2.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.640000 0.805000 6.195000 1.390000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.095000  2.660000 0.425000 3.245000 ;
      RECT 0.290000  0.085000 0.540000 0.670000 ;
      RECT 0.710000  0.390000 1.075000 0.670000 ;
      RECT 0.710000  0.670000 0.880000 1.930000 ;
      RECT 0.710000  1.930000 2.055000 2.100000 ;
      RECT 0.710000  2.100000 1.215000 2.990000 ;
      RECT 1.245000  0.085000 1.475000 0.670000 ;
      RECT 1.455000  2.270000 1.715000 3.245000 ;
      RECT 1.645000  0.390000 1.975000 1.555000 ;
      RECT 1.645000  1.555000 2.630000 1.760000 ;
      RECT 1.885000  2.100000 2.055000 2.875000 ;
      RECT 1.885000  2.875000 3.085000 3.045000 ;
      RECT 2.145000  0.370000 3.850000 0.525000 ;
      RECT 2.145000  0.525000 5.355000 0.540000 ;
      RECT 2.145000  0.540000 2.405000 1.345000 ;
      RECT 2.225000  1.760000 2.630000 1.885000 ;
      RECT 2.225000  1.885000 2.475000 2.695000 ;
      RECT 2.640000  0.710000 2.970000 1.040000 ;
      RECT 2.800000  1.040000 2.970000 1.500000 ;
      RECT 2.800000  1.500000 3.085000 2.875000 ;
      RECT 3.140000  0.710000 3.495000 1.275000 ;
      RECT 3.140000  1.275000 4.580000 1.330000 ;
      RECT 3.255000  1.330000 4.580000 1.475000 ;
      RECT 3.255000  1.475000 3.495000 2.690000 ;
      RECT 3.680000  0.540000 5.355000 0.695000 ;
      RECT 3.685000  1.645000 4.930000 1.815000 ;
      RECT 3.685000  1.815000 3.965000 1.975000 ;
      RECT 4.020000  0.085000 4.350000 0.355000 ;
      RECT 4.135000  1.985000 4.465000 3.245000 ;
      RECT 4.530000  0.865000 4.930000 1.105000 ;
      RECT 4.635000  1.815000 4.930000 2.225000 ;
      RECT 4.635000  2.225000 5.790000 2.395000 ;
      RECT 4.635000  2.395000 4.930000 3.075000 ;
      RECT 4.760000  1.105000 4.930000 1.645000 ;
      RECT 5.085000  0.305000 5.355000 0.525000 ;
      RECT 5.110000  0.695000 5.355000 1.795000 ;
      RECT 5.110000  1.795000 5.440000 2.055000 ;
      RECT 5.575000  0.085000 5.785000 0.635000 ;
      RECT 5.620000  1.560000 6.630000 1.730000 ;
      RECT 5.620000  1.730000 5.790000 2.225000 ;
      RECT 5.620000  2.565000 5.950000 3.245000 ;
      RECT 6.130000  1.910000 6.970000 2.080000 ;
      RECT 6.130000  2.080000 6.460000 2.440000 ;
      RECT 6.365000  0.305000 6.635000 0.985000 ;
      RECT 6.365000  0.985000 6.970000 1.155000 ;
      RECT 6.365000  1.345000 6.630000 1.560000 ;
      RECT 6.640000  2.250000 6.970000 3.245000 ;
      RECT 6.800000  1.155000 6.970000 1.185000 ;
      RECT 6.800000  1.185000 7.155000 1.515000 ;
      RECT 6.800000  1.515000 6.970000 1.910000 ;
      RECT 6.825000  0.085000 7.155000 0.815000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__sdlclkp_1
END LIBRARY
