* File: sky130_fd_sc_lp__dlybuf4s50kapwr_1.pxi.spice
* Created: Wed Sep  2 09:49:45 2020
* 
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A N_A_M1004_g N_A_M1007_g A A N_A_c_56_n
+ PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A_27_52# N_A_27_52#_M1004_s
+ N_A_27_52#_M1007_s N_A_27_52#_M1000_g N_A_27_52#_c_89_n N_A_27_52#_c_96_n
+ N_A_27_52#_c_97_n N_A_27_52#_c_90_n N_A_27_52#_c_91_n N_A_27_52#_c_98_n
+ N_A_27_52#_c_115_n N_A_27_52#_c_92_n N_A_27_52#_c_93_n N_A_27_52#_M1003_g
+ PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A_27_52#
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A_282_52# N_A_282_52#_M1003_d
+ N_A_282_52#_M1000_d N_A_282_52#_M1006_g N_A_282_52#_M1002_g
+ N_A_282_52#_c_158_n N_A_282_52#_c_159_n N_A_282_52#_c_164_n
+ N_A_282_52#_c_160_n N_A_282_52#_c_161_n N_A_282_52#_c_166_n
+ N_A_282_52#_c_162_n PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A_282_52#
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A_394_52# N_A_394_52#_M1006_s
+ N_A_394_52#_M1002_s N_A_394_52#_M1005_g N_A_394_52#_M1001_g
+ N_A_394_52#_c_231_n N_A_394_52#_c_233_n N_A_394_52#_c_235_n
+ N_A_394_52#_c_226_n N_A_394_52#_c_227_n N_A_394_52#_c_222_n
+ N_A_394_52#_c_223_n N_A_394_52#_c_251_n N_A_394_52#_c_224_n
+ PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%A_394_52#
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%KAPWR N_KAPWR_M1007_d N_KAPWR_M1002_d
+ KAPWR N_KAPWR_c_294_n N_KAPWR_c_306_n N_KAPWR_c_293_n KAPWR
+ PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%KAPWR
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%X N_X_M1005_d N_X_M1001_d X X X X X X X
+ N_X_c_330_n N_X_c_333_n X PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%X
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%VGND N_VGND_M1004_d N_VGND_M1006_d
+ N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n N_VGND_c_359_n VGND
+ N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n
+ PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%VGND
x_PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%VPWR VPWR N_VPWR_c_394_n VPWR
+ PM_SKY130_FD_SC_LP__DLYBUF4S50KAPWR_1%VPWR
cc_1 VNB N_A_M1004_g 0.0594522f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.47
cc_2 VNB A 0.0208018f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_56_n 0.0326678f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_4 VNB N_A_27_52#_c_89_n 0.0205357f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_5 VNB N_A_27_52#_c_90_n 0.0050785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_52#_c_91_n 0.0115829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_52#_c_92_n 0.00219081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_52#_c_93_n 0.0108849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_52#_M1003_g 0.0660704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_282_52#_c_158_n 0.011676f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_11 VNB N_A_282_52#_c_159_n 0.0150178f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.295
cc_12 VNB N_A_282_52#_c_160_n 0.0124045f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.665
cc_13 VNB N_A_282_52#_c_161_n 0.0396892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_282_52#_c_162_n 0.0419838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_394_52#_M1005_g 0.0517917f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A_394_52#_M1001_g 0.00175473f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_17 VNB N_A_394_52#_c_222_n 0.0138107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_394_52#_c_223_n 4.4684e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_394_52#_c_224_n 0.0349986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB X 0.0542411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_330_n 0.0186904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_356_n 0.00643581f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_VGND_c_357_n 0.0035061f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_24 VNB N_VGND_c_358_n 0.0503863f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_25 VNB N_VGND_c_359_n 0.00532387f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.665
cc_26 VNB N_VGND_c_360_n 0.0179296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_361_n 0.0230432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_362_n 0.22942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_363_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB VPWR 0.163682f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.335
cc_31 VPB N_A_M1007_g 0.0249089f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_32 VPB A 0.00827303f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_33 VPB N_A_c_56_n 0.00600603f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_34 VPB N_A_27_52#_M1000_g 0.046205f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_35 VPB N_A_27_52#_c_96_n 0.00794922f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_36 VPB N_A_27_52#_c_97_n 0.0273368f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.665
cc_37 VPB N_A_27_52#_c_98_n 0.00375793f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.5
cc_38 VPB N_A_27_52#_c_92_n 0.00495942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_52#_c_93_n 0.0365622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_282_52#_M1002_g 0.0711035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_282_52#_c_164_n 0.0102217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_282_52#_c_161_n 0.011742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_282_52#_c_166_n 0.0129165f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_394_52#_M1001_g 0.0248382f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_45 VPB N_A_394_52#_c_226_n 0.00281615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_394_52#_c_227_n 0.0023233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_394_52#_c_223_n 0.00305928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_KAPWR_c_293_n 0.0292908f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.5
cc_49 VPB X 0.00848832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB X 0.0427819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_X_c_333_n 0.0178335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB VPWR 0.045888f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.335
cc_53 VPB N_VPWR_c_394_n 0.105044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 A N_A_27_52#_M1007_s 0.00237131f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A_M1007_g N_A_27_52#_M1000_g 0.0257545f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_M1004_g N_A_27_52#_c_89_n 0.00946431f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_57 N_A_M1007_g N_A_27_52#_c_96_n 7.4234e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_58 A N_A_27_52#_c_96_n 0.0239868f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_59 N_A_c_56_n N_A_27_52#_c_96_n 7.87914e-19 $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_60 N_A_M1007_g N_A_27_52#_c_97_n 0.00978853f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_A_27_52#_c_90_n 0.0106533f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_62 A N_A_27_52#_c_90_n 0.0106601f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A_M1004_g N_A_27_52#_c_91_n 0.00435937f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_64 A N_A_27_52#_c_91_n 0.0289379f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_c_56_n N_A_27_52#_c_91_n 0.00100334f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_66 N_A_M1007_g N_A_27_52#_c_98_n 0.00881033f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_67 A N_A_27_52#_c_98_n 0.00941865f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_M1004_g N_A_27_52#_c_115_n 0.00261224f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_69 A N_A_27_52#_c_115_n 0.017308f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 A N_A_27_52#_c_92_n 0.0114464f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_c_56_n N_A_27_52#_c_92_n 0.00196087f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_72 A N_A_27_52#_c_93_n 3.24068e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_c_56_n N_A_27_52#_c_93_n 0.0257545f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_74 N_A_M1004_g N_A_27_52#_M1003_g 0.0257545f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_75 A N_A_27_52#_M1003_g 0.00183643f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_M1007_g N_KAPWR_c_294_n 0.00387353f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_M1007_g N_KAPWR_c_293_n 0.00453799f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_VGND_c_356_n 0.00322874f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_79 N_A_M1004_g N_VGND_c_360_n 0.00547602f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_80 N_A_M1004_g N_VGND_c_362_n 0.00694827f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_81 N_A_M1007_g VPWR 0.00638975f $X=0.475 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_82 N_A_M1007_g N_VPWR_c_394_n 0.0054895f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_27_52#_c_93_n N_A_282_52#_M1002_g 0.00287905f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_84 N_A_27_52#_c_115_n N_A_282_52#_c_159_n 0.0221959f $X=1.085 $Y=1.535 $X2=0
+ $Y2=0
cc_85 N_A_27_52#_c_92_n N_A_282_52#_c_159_n 0.00828764f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_86 N_A_27_52#_c_93_n N_A_282_52#_c_159_n 0.00414437f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_87 N_A_27_52#_M1003_g N_A_282_52#_c_159_n 0.00567511f $X=1.16 $Y=0.76 $X2=0
+ $Y2=0
cc_88 N_A_27_52#_M1000_g N_A_282_52#_c_164_n 0.00398828f $X=1.16 $Y=2.595 $X2=0
+ $Y2=0
cc_89 N_A_27_52#_c_92_n N_A_282_52#_c_164_n 0.0285056f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_90 N_A_27_52#_c_93_n N_A_282_52#_c_164_n 0.00361912f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_91 N_A_27_52#_c_93_n N_A_282_52#_c_161_n 0.00235448f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_92 N_A_27_52#_M1003_g N_A_282_52#_c_161_n 0.00316492f $X=1.16 $Y=0.76 $X2=0
+ $Y2=0
cc_93 N_A_27_52#_M1000_g N_A_282_52#_c_166_n 0.0170195f $X=1.16 $Y=2.595 $X2=0
+ $Y2=0
cc_94 N_A_27_52#_c_92_n N_A_282_52#_c_166_n 0.00501863f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_95 N_A_27_52#_c_93_n N_A_282_52#_c_166_n 0.00392394f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_96 N_A_27_52#_c_98_n N_KAPWR_M1007_d 0.00996866f $X=0.91 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_27_52#_M1000_g N_KAPWR_c_294_n 0.0160858f $X=1.16 $Y=2.595 $X2=0 $Y2=0
cc_98 N_A_27_52#_c_97_n N_KAPWR_c_294_n 0.0296181f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_99 N_A_27_52#_c_98_n N_KAPWR_c_294_n 0.0189214f $X=0.91 $Y=2.117 $X2=0 $Y2=0
cc_100 N_A_27_52#_c_92_n N_KAPWR_c_294_n 0.00107017f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_101 N_A_27_52#_M1000_g N_KAPWR_c_293_n 0.0157963f $X=1.16 $Y=2.595 $X2=0
+ $Y2=0
cc_102 N_A_27_52#_c_97_n N_KAPWR_c_293_n 0.0387447f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_103 N_A_27_52#_c_98_n N_KAPWR_c_293_n 0.0065323f $X=0.91 $Y=2.117 $X2=0 $Y2=0
cc_104 N_A_27_52#_c_92_n N_KAPWR_c_293_n 0.0116844f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A_27_52#_c_90_n N_VGND_M1004_d 0.00954115f $X=0.91 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_106 N_A_27_52#_c_90_n N_VGND_c_356_n 0.0207743f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_107 N_A_27_52#_M1003_g N_VGND_c_356_n 0.00356758f $X=1.16 $Y=0.76 $X2=0 $Y2=0
cc_108 N_A_27_52#_M1003_g N_VGND_c_358_n 0.0186549f $X=1.16 $Y=0.76 $X2=0 $Y2=0
cc_109 N_A_27_52#_c_89_n N_VGND_c_360_n 0.0152237f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_110 N_A_27_52#_c_89_n N_VGND_c_362_n 0.0118277f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_111 N_A_27_52#_c_90_n N_VGND_c_362_n 0.01767f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_112 N_A_27_52#_M1003_g N_VGND_c_362_n 0.0228755f $X=1.16 $Y=0.76 $X2=0 $Y2=0
cc_113 N_A_27_52#_M1007_s VPWR 0.00110569f $X=0.135 $Y=1.835 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_27_52#_M1000_g VPWR 0.0153579f $X=1.16 $Y=2.595 $X2=-0.19 $Y2=-0.245
cc_115 N_A_27_52#_c_97_n VPWR 0.00303861f $X=0.26 $Y=2.915 $X2=-0.19 $Y2=-0.245
cc_116 N_A_27_52#_M1000_g N_VPWR_c_394_n 0.0189208f $X=1.16 $Y=2.595 $X2=0 $Y2=0
cc_117 N_A_27_52#_c_97_n N_VPWR_c_394_n 0.0210467f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_118 N_A_282_52#_c_162_n N_A_394_52#_M1005_g 0.0251716f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_119 N_A_282_52#_M1002_g N_A_394_52#_M1001_g 0.0251716f $X=2.485 $Y=2.595
+ $X2=0 $Y2=0
cc_120 N_A_282_52#_c_158_n N_A_394_52#_c_231_n 0.0577683f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_121 N_A_282_52#_c_162_n N_A_394_52#_c_231_n 0.0289245f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_122 N_A_282_52#_c_160_n N_A_394_52#_c_233_n 0.0305669f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_123 N_A_282_52#_c_162_n N_A_394_52#_c_233_n 0.0415495f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_124 N_A_282_52#_c_158_n N_A_394_52#_c_235_n 0.00858119f $X=1.55 $Y=0.435
+ $X2=0 $Y2=0
cc_125 N_A_282_52#_c_159_n N_A_394_52#_c_235_n 0.0121129f $X=1.755 $Y=1.655
+ $X2=0 $Y2=0
cc_126 N_A_282_52#_c_160_n N_A_394_52#_c_235_n 0.0177106f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_127 N_A_282_52#_c_161_n N_A_394_52#_c_235_n 0.00503939f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_128 N_A_282_52#_c_162_n N_A_394_52#_c_235_n 8.78991e-19 $X=2.375 $Y=1.37
+ $X2=0 $Y2=0
cc_129 N_A_282_52#_M1002_g N_A_394_52#_c_226_n 0.0162472f $X=2.485 $Y=2.595
+ $X2=0 $Y2=0
cc_130 N_A_282_52#_c_160_n N_A_394_52#_c_226_n 0.0101562f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_131 N_A_282_52#_M1002_g N_A_394_52#_c_227_n 0.029647f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_132 N_A_282_52#_c_164_n N_A_394_52#_c_227_n 0.00990869f $X=1.755 $Y=2.1 $X2=0
+ $Y2=0
cc_133 N_A_282_52#_c_160_n N_A_394_52#_c_227_n 0.0270017f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_134 N_A_282_52#_c_161_n N_A_394_52#_c_227_n 0.00459953f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_135 N_A_282_52#_c_166_n N_A_394_52#_c_227_n 0.0129926f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_136 N_A_282_52#_c_160_n N_A_394_52#_c_222_n 0.0207685f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_137 N_A_282_52#_c_162_n N_A_394_52#_c_222_n 0.00694396f $X=2.375 $Y=1.37
+ $X2=0 $Y2=0
cc_138 N_A_282_52#_c_160_n N_A_394_52#_c_223_n 0.00227963f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_139 N_A_282_52#_c_161_n N_A_394_52#_c_223_n 0.00442182f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_140 N_A_282_52#_M1002_g N_A_394_52#_c_251_n 0.0248611f $X=2.485 $Y=2.595
+ $X2=0 $Y2=0
cc_141 N_A_282_52#_c_166_n N_A_394_52#_c_251_n 0.0649556f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_142 N_A_282_52#_c_161_n N_A_394_52#_c_224_n 0.0251716f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_143 N_A_282_52#_c_166_n N_KAPWR_c_294_n 0.0189978f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_144 N_A_282_52#_M1002_g N_KAPWR_c_306_n 0.0215549f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_145 N_A_282_52#_M1002_g N_KAPWR_c_293_n 0.0168329f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_146 N_A_282_52#_c_166_n N_KAPWR_c_293_n 0.0507826f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_147 N_A_282_52#_M1002_g N_X_c_333_n 8.17318e-19 $X=2.485 $Y=2.595 $X2=0 $Y2=0
cc_148 N_A_282_52#_c_162_n N_VGND_c_357_n 0.0176721f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_149 N_A_282_52#_c_158_n N_VGND_c_358_n 0.0250858f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_150 N_A_282_52#_c_162_n N_VGND_c_358_n 0.0173758f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_151 N_A_282_52#_c_158_n N_VGND_c_362_n 0.0155553f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_152 N_A_282_52#_c_162_n N_VGND_c_362_n 0.030234f $X=2.375 $Y=1.37 $X2=0 $Y2=0
cc_153 N_A_282_52#_M1000_d VPWR 0.00110569f $X=1.41 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_282_52#_M1002_g VPWR 0.0152399f $X=2.485 $Y=2.595 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_282_52#_c_166_n VPWR 0.00423096f $X=1.55 $Y=2.265 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_282_52#_M1002_g N_VPWR_c_394_n 0.0187841f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_157 N_A_282_52#_c_166_n N_VPWR_c_394_n 0.0301474f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_158 N_A_394_52#_c_226_n N_KAPWR_M1002_d 0.00441005f $X=2.855 $Y=1.91 $X2=0
+ $Y2=0
cc_159 N_A_394_52#_M1001_g N_KAPWR_c_306_n 0.00494635f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_394_52#_c_226_n N_KAPWR_c_306_n 0.0244283f $X=2.855 $Y=1.91 $X2=0
+ $Y2=0
cc_161 N_A_394_52#_c_227_n N_KAPWR_c_306_n 0.00665185f $X=2.54 $Y=1.91 $X2=0
+ $Y2=0
cc_162 N_A_394_52#_c_222_n N_KAPWR_c_306_n 5.09408e-19 $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_163 N_A_394_52#_c_251_n N_KAPWR_c_306_n 0.0235724f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_164 N_A_394_52#_M1002_s N_KAPWR_c_293_n 0.00186053f $X=1.97 $Y=2.095 $X2=0
+ $Y2=0
cc_165 N_A_394_52#_M1001_g N_KAPWR_c_293_n 0.00883115f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_394_52#_c_227_n N_KAPWR_c_293_n 0.00913551f $X=2.54 $Y=1.91 $X2=0
+ $Y2=0
cc_167 N_A_394_52#_c_251_n N_KAPWR_c_293_n 0.0312924f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_168 N_A_394_52#_M1005_g X 0.0163897f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_169 N_A_394_52#_M1001_g X 0.00381153f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_394_52#_c_222_n X 0.0389414f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_171 N_A_394_52#_c_223_n X 0.00696747f $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_172 N_A_394_52#_c_224_n X 0.00819462f $X=3.26 $Y=1.46 $X2=0 $Y2=0
cc_173 N_A_394_52#_M1001_g X 0.0134471f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_394_52#_M1005_g N_X_c_330_n 0.00495371f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A_394_52#_c_222_n N_X_c_330_n 0.00268942f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_176 N_A_394_52#_c_224_n N_X_c_330_n 0.00229273f $X=3.26 $Y=1.46 $X2=0 $Y2=0
cc_177 N_A_394_52#_M1001_g N_X_c_333_n 0.00406351f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_394_52#_c_226_n N_X_c_333_n 0.012527f $X=2.855 $Y=1.91 $X2=0 $Y2=0
cc_179 N_A_394_52#_c_222_n N_X_c_333_n 0.00881742f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_180 N_A_394_52#_c_223_n N_X_c_333_n 6.43138e-19 $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_181 N_A_394_52#_c_224_n N_X_c_333_n 0.00425967f $X=3.26 $Y=1.46 $X2=0 $Y2=0
cc_182 N_A_394_52#_c_233_n N_VGND_M1006_d 0.00205184f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_183 N_A_394_52#_c_222_n N_VGND_M1006_d 0.00293623f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_184 N_A_394_52#_M1005_g N_VGND_c_357_n 0.00514775f $X=3.17 $Y=0.47 $X2=0
+ $Y2=0
cc_185 N_A_394_52#_c_231_n N_VGND_c_357_n 0.0133572f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_186 N_A_394_52#_c_233_n N_VGND_c_357_n 0.00446569f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_187 N_A_394_52#_c_222_n N_VGND_c_357_n 0.0103475f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_188 N_A_394_52#_c_231_n N_VGND_c_358_n 0.0140261f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_189 N_A_394_52#_M1005_g N_VGND_c_361_n 0.0051159f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_190 N_A_394_52#_M1005_g N_VGND_c_362_n 0.0104241f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_191 N_A_394_52#_c_231_n N_VGND_c_362_n 0.00945114f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_192 N_A_394_52#_M1002_s VPWR 0.00127104f $X=1.97 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_394_52#_M1001_g VPWR 0.00656747f $X=3.17 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_394_52#_c_251_n VPWR 0.00228685f $X=2.095 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_394_52#_M1001_g N_VPWR_c_394_n 0.00564131f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A_394_52#_c_251_n N_VPWR_c_394_n 0.0153681f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_197 N_KAPWR_c_306_n X 0.0357183f $X=2.875 $Y=2.27 $X2=0 $Y2=0
cc_198 N_KAPWR_c_293_n X 0.056983f $X=2.875 $Y=2.81 $X2=0 $Y2=0
cc_199 N_KAPWR_M1007_d VPWR 0.0016543f $X=0.55 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_200 N_KAPWR_M1002_d VPWR 0.00169056f $X=2.735 $Y=2.095 $X2=-0.19 $Y2=1.655
cc_201 N_KAPWR_c_294_n VPWR 0.00306447f $X=0.76 $Y=2.49 $X2=-0.19 $Y2=1.655
cc_202 N_KAPWR_c_306_n VPWR 0.00303333f $X=2.875 $Y=2.27 $X2=-0.19 $Y2=1.655
cc_203 N_KAPWR_c_293_n VPWR 0.38781f $X=2.875 $Y=2.81 $X2=-0.19 $Y2=1.655
cc_204 N_KAPWR_c_294_n N_VPWR_c_394_n 0.0206605f $X=0.76 $Y=2.49 $X2=0 $Y2=0
cc_205 N_KAPWR_c_306_n N_VPWR_c_394_n 0.0209582f $X=2.875 $Y=2.27 $X2=0 $Y2=0
cc_206 N_KAPWR_c_293_n N_VPWR_c_394_n 0.00908252f $X=2.875 $Y=2.81 $X2=0 $Y2=0
cc_207 N_X_c_330_n N_VGND_c_361_n 0.0254f $X=3.632 $Y=0.475 $X2=0 $Y2=0
cc_208 N_X_c_330_n N_VGND_c_362_n 0.0197894f $X=3.632 $Y=0.475 $X2=0 $Y2=0
cc_209 N_X_M1001_d VPWR 0.00110569f $X=3.245 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_210 X VPWR 0.00483484f $X=3.515 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_211 X N_VPWR_c_394_n 0.0347023f $X=3.515 $Y=1.95 $X2=0 $Y2=0
