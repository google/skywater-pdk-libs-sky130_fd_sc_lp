* File: sky130_fd_sc_lp__or3b_4.pxi.spice
* Created: Wed Sep  2 10:31:19 2020
* 
x_PM_SKY130_FD_SC_LP__OR3B_4%C_N N_C_N_M1015_g N_C_N_M1014_g C_N C_N C_N C_N C_N
+ N_C_N_c_87_n N_C_N_c_88_n PM_SKY130_FD_SC_LP__OR3B_4%C_N
x_PM_SKY130_FD_SC_LP__OR3B_4%A_253_23# N_A_253_23#_M1004_d N_A_253_23#_M1006_d
+ N_A_253_23#_M1000_d N_A_253_23#_M1003_g N_A_253_23#_M1001_g
+ N_A_253_23#_M1009_g N_A_253_23#_M1002_g N_A_253_23#_M1011_g
+ N_A_253_23#_M1008_g N_A_253_23#_M1012_g N_A_253_23#_M1013_g
+ N_A_253_23#_c_119_n N_A_253_23#_c_120_n N_A_253_23#_c_121_n
+ N_A_253_23#_c_217_p N_A_253_23#_c_159_p N_A_253_23#_c_122_n
+ N_A_253_23#_c_123_n N_A_253_23#_c_124_n N_A_253_23#_c_132_n
+ N_A_253_23#_c_133_n N_A_253_23#_c_125_n N_A_253_23#_c_134_n
+ N_A_253_23#_c_126_n N_A_253_23#_c_127_n PM_SKY130_FD_SC_LP__OR3B_4%A_253_23#
x_PM_SKY130_FD_SC_LP__OR3B_4%A N_A_M1004_g N_A_M1010_g A A N_A_c_254_n
+ N_A_c_255_n PM_SKY130_FD_SC_LP__OR3B_4%A
x_PM_SKY130_FD_SC_LP__OR3B_4%B N_B_M1005_g N_B_M1007_g B B N_B_c_293_n
+ N_B_c_294_n PM_SKY130_FD_SC_LP__OR3B_4%B
x_PM_SKY130_FD_SC_LP__OR3B_4%A_49_133# N_A_49_133#_M1015_s N_A_49_133#_M1014_s
+ N_A_49_133#_M1006_g N_A_49_133#_M1000_g N_A_49_133#_c_331_n
+ N_A_49_133#_c_337_n N_A_49_133#_c_338_n N_A_49_133#_c_332_n
+ N_A_49_133#_c_333_n N_A_49_133#_c_334_n PM_SKY130_FD_SC_LP__OR3B_4%A_49_133#
x_PM_SKY130_FD_SC_LP__OR3B_4%VPWR N_VPWR_M1014_d N_VPWR_M1002_s N_VPWR_M1013_s
+ N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n
+ N_VPWR_c_411_n N_VPWR_c_412_n VPWR N_VPWR_c_413_n N_VPWR_c_414_n
+ N_VPWR_c_405_n N_VPWR_c_416_n PM_SKY130_FD_SC_LP__OR3B_4%VPWR
x_PM_SKY130_FD_SC_LP__OR3B_4%X N_X_M1003_s N_X_M1011_s N_X_M1001_d N_X_M1008_d
+ N_X_c_459_n N_X_c_460_n N_X_c_461_n N_X_c_509_p N_X_c_462_n N_X_c_510_p
+ N_X_c_463_n X X X X X PM_SKY130_FD_SC_LP__OR3B_4%X
x_PM_SKY130_FD_SC_LP__OR3B_4%VGND N_VGND_M1015_d N_VGND_M1009_d N_VGND_M1012_d
+ N_VGND_M1007_d N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n
+ N_VGND_c_525_n N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n
+ N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n VGND N_VGND_c_533_n
+ N_VGND_c_534_n PM_SKY130_FD_SC_LP__OR3B_4%VGND
cc_1 VNB N_C_N_M1014_g 0.00775418f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.045
cc_2 VNB C_N 0.00750026f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_3 VNB N_C_N_c_87_n 0.0435522f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_4 VNB N_C_N_c_88_n 0.0222097f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.195
cc_5 VNB N_A_253_23#_M1003_g 0.0267214f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_6 VNB N_A_253_23#_M1009_g 0.0222417f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_7 VNB N_A_253_23#_M1011_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.295
cc_8 VNB N_A_253_23#_M1012_g 0.0238888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_253_23#_c_119_n 0.00328096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_253_23#_c_120_n 0.00208003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_253_23#_c_121_n 0.00434633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_253_23#_c_122_n 0.00585184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_253_23#_c_123_n 0.0388491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_253_23#_c_124_n 0.00760296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_253_23#_c_125_n 0.0124234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_253_23#_c_126_n 0.0230885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_253_23#_c_127_n 0.0684616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_M1004_g 0.0247972f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.875
cc_19 VNB N_A_c_254_n 0.0259056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_255_n 9.66218e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_M1007_g 0.0251986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_293_n 0.0238929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_294_n 0.00321801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_49_133#_M1006_g 0.031278f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_25 VNB N_A_49_133#_c_331_n 0.0435214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_49_133#_c_332_n 3.70724e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_49_133#_c_333_n 0.00590888f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.295
cc_28 VNB N_A_49_133#_c_334_n 0.0271237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_405_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_459_n 0.00731156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_460_n 0.00121166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_461_n 0.00146247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_462_n 0.00567396f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.195
cc_34 VNB N_X_c_463_n 0.00172486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_521_n 0.00485741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_522_n 4.90414e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.36
cc_37 VNB N_VGND_c_523_n 0.004684f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.555
cc_38 VNB N_VGND_c_524_n 0.0052823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_525_n 0.0318901f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.665
cc_40 VNB N_VGND_c_526_n 0.00490486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_527_n 0.0146736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_528_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_529_n 0.0153253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_530_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_531_n 0.0170436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_532_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_533_n 0.0222964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_534_n 0.270565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VPB N_C_N_M1014_g 0.0238168f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.045
cc_50 VPB C_N 0.0012647f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_51 VPB N_A_253_23#_M1001_g 0.0220117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_253_23#_M1002_g 0.0183264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_253_23#_M1008_g 0.0183478f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.035
cc_54 VPB N_A_253_23#_M1013_g 0.0200463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_253_23#_c_132_n 0.0168454f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_253_23#_c_133_n 0.0338754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_253_23#_c_134_n 0.0139053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_253_23#_c_126_n 0.00780318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_253_23#_c_127_n 0.0113369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_M1010_g 0.018717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_c_254_n 0.00686048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_c_255_n 0.00169877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_B_M1005_g 0.0177506f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.875
cc_64 VPB N_B_c_293_n 0.00678108f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B_c_294_n 0.0021342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_49_133#_M1000_g 0.0241645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_49_133#_c_331_n 0.0278078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_49_133#_c_337_n 0.0205679f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.195
cc_69 VPB N_A_49_133#_c_338_n 0.0127947f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.525
cc_70 VPB N_A_49_133#_c_332_n 0.00115408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_49_133#_c_334_n 0.00787462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_406_n 0.0199016f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_73 VPB N_VPWR_c_407_n 3.18512e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_408_n 0.00498793f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.36
cc_75 VPB N_VPWR_c_409_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.555
cc_76 VPB N_VPWR_c_410_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_411_n 0.0175054f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.925
cc_78 VPB N_VPWR_c_412_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_413_n 0.0338062f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.665
cc_80 VPB N_VPWR_c_414_n 0.0509108f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_405_n 0.0617843f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_416_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_X_c_459_n 0.003413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB X 0.00821584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 C_N N_A_253_23#_M1003_g 0.00230001f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_86 N_C_N_c_87_n N_A_253_23#_M1003_g 0.00786953f $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_87 N_C_N_c_88_n N_A_253_23#_M1003_g 0.00611836f $X=0.697 $Y=1.195 $X2=0 $Y2=0
cc_88 C_N N_A_253_23#_M1001_g 0.00103663f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_89 N_C_N_M1014_g N_A_253_23#_c_127_n 0.0120606f $X=0.585 $Y=2.045 $X2=0 $Y2=0
cc_90 N_C_N_c_87_n N_A_253_23#_c_127_n 7.14624e-19 $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_91 C_N N_A_49_133#_c_331_n 0.0791337f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_92 N_C_N_c_88_n N_A_49_133#_c_331_n 0.0213263f $X=0.697 $Y=1.195 $X2=0 $Y2=0
cc_93 N_C_N_M1014_g N_A_49_133#_c_337_n 0.0118035f $X=0.585 $Y=2.045 $X2=0 $Y2=0
cc_94 C_N N_A_49_133#_c_337_n 0.0130299f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_95 C_N N_VPWR_M1014_d 0.00405642f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_96 N_C_N_M1014_g N_X_c_459_n 0.00205359f $X=0.585 $Y=2.045 $X2=0 $Y2=0
cc_97 C_N N_X_c_459_n 0.067878f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_98 N_C_N_c_87_n N_X_c_459_n 0.00235976f $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_99 C_N N_X_c_461_n 0.0143412f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_100 N_C_N_c_87_n N_X_c_461_n 4.65549e-19 $X=0.72 $Y=1.36 $X2=0 $Y2=0
cc_101 N_C_N_c_88_n N_X_c_461_n 3.86395e-19 $X=0.697 $Y=1.195 $X2=0 $Y2=0
cc_102 C_N N_VGND_M1015_d 0.00505218f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_103 C_N N_VGND_c_521_n 0.0333643f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_104 N_C_N_c_88_n N_VGND_c_521_n 0.00102461f $X=0.697 $Y=1.195 $X2=0 $Y2=0
cc_105 C_N N_VGND_c_525_n 0.00623633f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_106 N_C_N_c_88_n N_VGND_c_525_n 0.00319672f $X=0.697 $Y=1.195 $X2=0 $Y2=0
cc_107 C_N N_VGND_c_534_n 0.00710559f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_108 N_C_N_c_88_n N_VGND_c_534_n 0.00354586f $X=0.697 $Y=1.195 $X2=0 $Y2=0
cc_109 N_A_253_23#_M1012_g N_A_M1004_g 0.0171601f $X=2.63 $Y=0.665 $X2=0 $Y2=0
cc_110 N_A_253_23#_c_120_n N_A_M1004_g 0.00343808f $X=2.765 $Y=1.415 $X2=0 $Y2=0
cc_111 N_A_253_23#_c_121_n N_A_M1004_g 0.0144173f $X=3.22 $Y=1.09 $X2=0 $Y2=0
cc_112 N_A_253_23#_M1013_g N_A_M1010_g 0.0345181f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_253_23#_c_119_n N_A_c_254_n 0.00162512f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_114 N_A_253_23#_c_120_n N_A_c_254_n 4.22693e-19 $X=2.765 $Y=1.415 $X2=0 $Y2=0
cc_115 N_A_253_23#_c_121_n N_A_c_254_n 0.00300998f $X=3.22 $Y=1.09 $X2=0 $Y2=0
cc_116 N_A_253_23#_c_124_n N_A_c_254_n 7.12607e-19 $X=3.362 $Y=1.09 $X2=0 $Y2=0
cc_117 N_A_253_23#_c_127_n N_A_c_254_n 0.0208365f $X=2.63 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A_253_23#_M1013_g N_A_c_255_n 0.00515946f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_253_23#_c_119_n N_A_c_255_n 0.0190588f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_120 N_A_253_23#_c_120_n N_A_c_255_n 0.00512111f $X=2.765 $Y=1.415 $X2=0 $Y2=0
cc_121 N_A_253_23#_c_121_n N_A_c_255_n 0.0153044f $X=3.22 $Y=1.09 $X2=0 $Y2=0
cc_122 N_A_253_23#_c_124_n N_A_c_255_n 0.00481434f $X=3.362 $Y=1.09 $X2=0 $Y2=0
cc_123 N_A_253_23#_c_127_n N_A_c_255_n 4.67307e-19 $X=2.63 $Y=1.51 $X2=0 $Y2=0
cc_124 N_A_253_23#_c_132_n N_B_M1005_g 0.00145067f $X=4.32 $Y=2.91 $X2=0 $Y2=0
cc_125 N_A_253_23#_c_159_p N_B_M1007_g 0.00996904f $X=3.355 $Y=0.42 $X2=0 $Y2=0
cc_126 N_A_253_23#_c_122_n N_B_M1007_g 0.012748f $X=4.175 $Y=1.09 $X2=0 $Y2=0
cc_127 N_A_253_23#_c_123_n N_B_M1007_g 3.74669e-19 $X=4.32 $Y=0.42 $X2=0 $Y2=0
cc_128 N_A_253_23#_c_124_n N_B_M1007_g 0.00133542f $X=3.362 $Y=1.09 $X2=0 $Y2=0
cc_129 N_A_253_23#_c_122_n N_B_c_293_n 0.00370552f $X=4.175 $Y=1.09 $X2=0 $Y2=0
cc_130 N_A_253_23#_c_122_n N_B_c_294_n 0.0181426f $X=4.175 $Y=1.09 $X2=0 $Y2=0
cc_131 N_A_253_23#_c_124_n N_B_c_294_n 0.00541498f $X=3.362 $Y=1.09 $X2=0 $Y2=0
cc_132 N_A_253_23#_c_159_p N_A_49_133#_M1006_g 3.82399e-19 $X=3.355 $Y=0.42
+ $X2=0 $Y2=0
cc_133 N_A_253_23#_c_122_n N_A_49_133#_M1006_g 0.0131224f $X=4.175 $Y=1.09 $X2=0
+ $Y2=0
cc_134 N_A_253_23#_c_123_n N_A_49_133#_M1006_g 0.0113063f $X=4.32 $Y=0.42 $X2=0
+ $Y2=0
cc_135 N_A_253_23#_c_125_n N_A_49_133#_M1006_g 0.00217175f $X=4.442 $Y=1.09
+ $X2=0 $Y2=0
cc_136 N_A_253_23#_c_126_n N_A_49_133#_M1006_g 0.00340142f $X=4.485 $Y=1.815
+ $X2=0 $Y2=0
cc_137 N_A_253_23#_c_132_n N_A_49_133#_M1000_g 0.00791029f $X=4.32 $Y=2.91 $X2=0
+ $Y2=0
cc_138 N_A_253_23#_c_134_n N_A_49_133#_M1000_g 0.0119249f $X=4.345 $Y=1.98 $X2=0
+ $Y2=0
cc_139 N_A_253_23#_c_126_n N_A_49_133#_M1000_g 0.001576f $X=4.485 $Y=1.815 $X2=0
+ $Y2=0
cc_140 N_A_253_23#_M1001_g N_A_49_133#_c_337_n 0.0135613f $X=1.375 $Y=2.465
+ $X2=0 $Y2=0
cc_141 N_A_253_23#_M1002_g N_A_49_133#_c_337_n 0.0118101f $X=1.805 $Y=2.465
+ $X2=0 $Y2=0
cc_142 N_A_253_23#_M1008_g N_A_49_133#_c_337_n 0.0118101f $X=2.235 $Y=2.465
+ $X2=0 $Y2=0
cc_143 N_A_253_23#_M1013_g N_A_49_133#_c_337_n 0.0128109f $X=2.665 $Y=2.465
+ $X2=0 $Y2=0
cc_144 N_A_253_23#_c_119_n N_A_49_133#_c_337_n 0.00299097f $X=2.68 $Y=1.53 $X2=0
+ $Y2=0
cc_145 N_A_253_23#_c_133_n N_A_49_133#_c_337_n 0.0143326f $X=4.432 $Y=2.76 $X2=0
+ $Y2=0
cc_146 N_A_253_23#_c_134_n N_A_49_133#_c_332_n 0.0379014f $X=4.345 $Y=1.98 $X2=0
+ $Y2=0
cc_147 N_A_253_23#_c_126_n N_A_49_133#_c_332_n 0.00422426f $X=4.485 $Y=1.815
+ $X2=0 $Y2=0
cc_148 N_A_253_23#_c_122_n N_A_49_133#_c_333_n 0.0188979f $X=4.175 $Y=1.09 $X2=0
+ $Y2=0
cc_149 N_A_253_23#_c_125_n N_A_49_133#_c_333_n 0.0154781f $X=4.442 $Y=1.09 $X2=0
+ $Y2=0
cc_150 N_A_253_23#_c_134_n N_A_49_133#_c_333_n 0.00829455f $X=4.345 $Y=1.98
+ $X2=0 $Y2=0
cc_151 N_A_253_23#_c_126_n N_A_49_133#_c_333_n 0.0231087f $X=4.485 $Y=1.815
+ $X2=0 $Y2=0
cc_152 N_A_253_23#_c_125_n N_A_49_133#_c_334_n 0.00419322f $X=4.442 $Y=1.09
+ $X2=0 $Y2=0
cc_153 N_A_253_23#_c_134_n N_A_49_133#_c_334_n 0.00239124f $X=4.345 $Y=1.98
+ $X2=0 $Y2=0
cc_154 N_A_253_23#_c_126_n N_A_49_133#_c_334_n 0.00290875f $X=4.485 $Y=1.815
+ $X2=0 $Y2=0
cc_155 N_A_253_23#_M1001_g N_VPWR_c_406_n 0.0151619f $X=1.375 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_253_23#_M1002_g N_VPWR_c_406_n 0.00172252f $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_253_23#_M1001_g N_VPWR_c_407_n 0.00172252f $X=1.375 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_253_23#_M1002_g N_VPWR_c_407_n 0.0131009f $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_253_23#_M1008_g N_VPWR_c_407_n 0.0135932f $X=2.235 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_253_23#_M1013_g N_VPWR_c_407_n 0.00177278f $X=2.665 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_253_23#_M1013_g N_VPWR_c_408_n 0.00242503f $X=2.665 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_253_23#_M1001_g N_VPWR_c_409_n 0.00486043f $X=1.375 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_253_23#_M1002_g N_VPWR_c_409_n 0.00486043f $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_253_23#_M1008_g N_VPWR_c_411_n 0.00486043f $X=2.235 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_253_23#_M1013_g N_VPWR_c_411_n 0.00585385f $X=2.665 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_253_23#_c_132_n N_VPWR_c_414_n 0.0369586f $X=4.32 $Y=2.91 $X2=0 $Y2=0
cc_167 N_A_253_23#_M1000_d N_VPWR_c_405_n 0.00244481f $X=4.18 $Y=1.835 $X2=0
+ $Y2=0
cc_168 N_A_253_23#_M1001_g N_VPWR_c_405_n 0.00462979f $X=1.375 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_253_23#_M1002_g N_VPWR_c_405_n 0.00462979f $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_253_23#_M1008_g N_VPWR_c_405_n 0.00462979f $X=2.235 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_253_23#_M1013_g N_VPWR_c_405_n 0.00664543f $X=2.665 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_253_23#_c_132_n N_VPWR_c_405_n 0.0212417f $X=4.32 $Y=2.91 $X2=0 $Y2=0
cc_173 N_A_253_23#_M1003_g N_X_c_459_n 0.00513677f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A_253_23#_c_119_n N_X_c_459_n 0.0182946f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_175 N_A_253_23#_c_127_n N_X_c_459_n 0.00637925f $X=2.63 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A_253_23#_M1003_g N_X_c_460_n 0.0162165f $X=1.34 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A_253_23#_c_119_n N_X_c_460_n 0.00522319f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_178 N_A_253_23#_M1009_g N_X_c_462_n 0.0140849f $X=1.77 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_253_23#_M1011_g N_X_c_462_n 0.0137525f $X=2.2 $Y=0.665 $X2=0 $Y2=0
cc_180 N_A_253_23#_M1012_g N_X_c_462_n 0.00131397f $X=2.63 $Y=0.665 $X2=0 $Y2=0
cc_181 N_A_253_23#_c_119_n N_X_c_462_n 0.0634453f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_182 N_A_253_23#_c_120_n N_X_c_462_n 0.00561291f $X=2.765 $Y=1.415 $X2=0 $Y2=0
cc_183 N_A_253_23#_c_217_p N_X_c_462_n 0.00839918f $X=2.85 $Y=1.09 $X2=0 $Y2=0
cc_184 N_A_253_23#_c_127_n N_X_c_462_n 0.00526937f $X=2.63 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A_253_23#_c_119_n N_X_c_463_n 0.0181083f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_186 N_A_253_23#_c_127_n N_X_c_463_n 0.00268515f $X=2.63 $Y=1.51 $X2=0 $Y2=0
cc_187 N_A_253_23#_M1001_g X 0.0149999f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_253_23#_M1002_g X 0.0129491f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_253_23#_M1008_g X 0.0129491f $X=2.235 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_253_23#_M1013_g X 0.0106999f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_253_23#_c_119_n X 0.103703f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_192 N_A_253_23#_c_127_n X 0.00842638f $X=2.63 $Y=1.51 $X2=0 $Y2=0
cc_193 N_A_253_23#_c_121_n N_VGND_M1012_d 0.00166894f $X=3.22 $Y=1.09 $X2=0
+ $Y2=0
cc_194 N_A_253_23#_c_217_p N_VGND_M1012_d 9.7203e-19 $X=2.85 $Y=1.09 $X2=0 $Y2=0
cc_195 N_A_253_23#_c_122_n N_VGND_M1007_d 0.0029901f $X=4.175 $Y=1.09 $X2=0
+ $Y2=0
cc_196 N_A_253_23#_M1003_g N_VGND_c_521_n 0.00335739f $X=1.34 $Y=0.665 $X2=0
+ $Y2=0
cc_197 N_A_253_23#_M1003_g N_VGND_c_522_n 6.27137e-19 $X=1.34 $Y=0.665 $X2=0
+ $Y2=0
cc_198 N_A_253_23#_M1009_g N_VGND_c_522_n 0.0113053f $X=1.77 $Y=0.665 $X2=0
+ $Y2=0
cc_199 N_A_253_23#_M1011_g N_VGND_c_522_n 0.0113264f $X=2.2 $Y=0.665 $X2=0 $Y2=0
cc_200 N_A_253_23#_M1012_g N_VGND_c_522_n 6.30876e-19 $X=2.63 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_253_23#_M1012_g N_VGND_c_523_n 0.00168948f $X=2.63 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_253_23#_c_121_n N_VGND_c_523_n 0.0128182f $X=3.22 $Y=1.09 $X2=0 $Y2=0
cc_203 N_A_253_23#_c_217_p N_VGND_c_523_n 0.00789872f $X=2.85 $Y=1.09 $X2=0
+ $Y2=0
cc_204 N_A_253_23#_c_122_n N_VGND_c_524_n 0.0220482f $X=4.175 $Y=1.09 $X2=0
+ $Y2=0
cc_205 N_A_253_23#_M1003_g N_VGND_c_527_n 0.00575161f $X=1.34 $Y=0.665 $X2=0
+ $Y2=0
cc_206 N_A_253_23#_M1009_g N_VGND_c_527_n 0.00477554f $X=1.77 $Y=0.665 $X2=0
+ $Y2=0
cc_207 N_A_253_23#_M1011_g N_VGND_c_529_n 0.00477554f $X=2.2 $Y=0.665 $X2=0
+ $Y2=0
cc_208 N_A_253_23#_M1012_g N_VGND_c_529_n 0.00575161f $X=2.63 $Y=0.665 $X2=0
+ $Y2=0
cc_209 N_A_253_23#_c_159_p N_VGND_c_531_n 0.0160847f $X=3.355 $Y=0.42 $X2=0
+ $Y2=0
cc_210 N_A_253_23#_c_123_n N_VGND_c_533_n 0.0358127f $X=4.32 $Y=0.42 $X2=0 $Y2=0
cc_211 N_A_253_23#_M1004_d N_VGND_c_534_n 0.00240953f $X=3.215 $Y=0.245 $X2=0
+ $Y2=0
cc_212 N_A_253_23#_M1006_d N_VGND_c_534_n 0.00212301f $X=4.18 $Y=0.245 $X2=0
+ $Y2=0
cc_213 N_A_253_23#_M1003_g N_VGND_c_534_n 0.0118214f $X=1.34 $Y=0.665 $X2=0
+ $Y2=0
cc_214 N_A_253_23#_M1009_g N_VGND_c_534_n 0.00825815f $X=1.77 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_253_23#_M1011_g N_VGND_c_534_n 0.00825815f $X=2.2 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_253_23#_M1012_g N_VGND_c_534_n 0.0107552f $X=2.63 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_253_23#_c_159_p N_VGND_c_534_n 0.010888f $X=3.355 $Y=0.42 $X2=0 $Y2=0
cc_218 N_A_253_23#_c_123_n N_VGND_c_534_n 0.0206303f $X=4.32 $Y=0.42 $X2=0 $Y2=0
cc_219 N_A_M1010_g N_B_M1005_g 0.0587523f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A_M1004_g N_B_M1007_g 0.0238362f $X=3.14 $Y=0.665 $X2=0 $Y2=0
cc_221 N_A_c_254_n N_B_c_293_n 0.0587523f $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_222 N_A_c_255_n N_B_c_293_n 9.12849e-19 $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_223 N_A_c_254_n N_B_c_294_n 0.00347495f $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_224 N_A_c_255_n N_B_c_294_n 0.048827f $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_225 N_A_M1010_g N_A_49_133#_c_337_n 0.0122589f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_c_254_n N_A_49_133#_c_337_n 0.00188461f $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_227 N_A_c_255_n N_A_49_133#_c_337_n 0.0151999f $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_c_255_n N_VPWR_M1013_s 0.0039973f $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_229 N_A_M1010_g N_VPWR_c_408_n 0.00391869f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_M1010_g N_VPWR_c_414_n 0.00585385f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_M1010_g N_VPWR_c_405_n 0.00647749f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_M1010_g X 3.52111e-19 $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A_c_255_n X 0.0173638f $X=3.115 $Y=1.51 $X2=0 $Y2=0
cc_234 N_A_M1004_g N_VGND_c_523_n 0.00176321f $X=3.14 $Y=0.665 $X2=0 $Y2=0
cc_235 N_A_M1004_g N_VGND_c_531_n 0.00575161f $X=3.14 $Y=0.665 $X2=0 $Y2=0
cc_236 N_A_M1004_g N_VGND_c_534_n 0.0107806f $X=3.14 $Y=0.665 $X2=0 $Y2=0
cc_237 N_B_M1007_g N_A_49_133#_M1006_g 0.0176694f $X=3.57 $Y=0.665 $X2=0 $Y2=0
cc_238 N_B_M1005_g N_A_49_133#_M1000_g 0.0473992f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B_c_294_n N_A_49_133#_M1000_g 0.00137748f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_240 N_B_M1005_g N_A_49_133#_c_337_n 0.0120754f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B_c_293_n N_A_49_133#_c_337_n 0.00209032f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_242 N_B_c_294_n N_A_49_133#_c_337_n 0.0148433f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_243 N_B_M1005_g N_A_49_133#_c_332_n 0.00451271f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B_c_294_n N_A_49_133#_c_332_n 0.0367228f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_245 N_B_c_293_n N_A_49_133#_c_333_n 0.00204499f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_246 N_B_c_294_n N_A_49_133#_c_333_n 0.0230416f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_247 N_B_c_293_n N_A_49_133#_c_334_n 0.0204692f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_248 N_B_c_294_n N_A_49_133#_c_334_n 2.93344e-19 $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_249 N_B_M1005_g N_VPWR_c_414_n 0.00585385f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_250 N_B_M1005_g N_VPWR_c_405_n 0.00666612f $X=3.565 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B_c_294_n A_728_367# 0.00328939f $X=3.655 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_252 N_B_M1007_g N_VGND_c_524_n 0.00173081f $X=3.57 $Y=0.665 $X2=0 $Y2=0
cc_253 N_B_M1007_g N_VGND_c_531_n 0.00561712f $X=3.57 $Y=0.665 $X2=0 $Y2=0
cc_254 N_B_M1007_g N_VGND_c_534_n 0.0105764f $X=3.57 $Y=0.665 $X2=0 $Y2=0
cc_255 N_A_49_133#_c_337_n N_VPWR_M1014_d 0.0051849f $X=3.92 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_256 N_A_49_133#_c_337_n N_VPWR_M1002_s 0.00342847f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A_49_133#_c_337_n N_VPWR_M1013_s 0.0098468f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A_49_133#_c_337_n N_VPWR_c_406_n 0.021529f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_259 N_A_49_133#_c_337_n N_VPWR_c_407_n 0.016709f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_49_133#_c_337_n N_VPWR_c_408_n 0.0219723f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A_49_133#_M1000_g N_VPWR_c_414_n 0.0054895f $X=4.105 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_A_49_133#_M1000_g N_VPWR_c_405_n 0.00961856f $X=4.105 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_A_49_133#_c_337_n N_VPWR_c_405_n 0.088613f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_49_133#_c_338_n N_VPWR_c_405_n 0.00977402f $X=0.455 $Y=2.4 $X2=0
+ $Y2=0
cc_265 N_A_49_133#_c_337_n N_X_M1001_d 0.00503872f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_266 N_A_49_133#_c_337_n N_X_M1008_d 0.00503872f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_267 N_A_49_133#_c_337_n N_X_c_459_n 0.0146845f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_268 N_A_49_133#_c_337_n X 0.0840767f $X=3.92 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A_49_133#_c_337_n A_656_367# 0.0056012f $X=3.92 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_270 N_A_49_133#_c_337_n A_728_367# 0.0115932f $X=3.92 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_271 N_A_49_133#_c_332_n A_728_367# 0.00490017f $X=4.005 $Y=2.315 $X2=-0.19
+ $Y2=-0.245
cc_272 N_A_49_133#_M1006_g N_VGND_c_524_n 0.00314823f $X=4.105 $Y=0.665 $X2=0
+ $Y2=0
cc_273 N_A_49_133#_c_331_n N_VGND_c_525_n 0.00412163f $X=0.37 $Y=0.875 $X2=0
+ $Y2=0
cc_274 N_A_49_133#_M1006_g N_VGND_c_533_n 0.00569184f $X=4.105 $Y=0.665 $X2=0
+ $Y2=0
cc_275 N_A_49_133#_M1006_g N_VGND_c_534_n 0.0117802f $X=4.105 $Y=0.665 $X2=0
+ $Y2=0
cc_276 N_A_49_133#_c_331_n N_VGND_c_534_n 0.00711232f $X=0.37 $Y=0.875 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_405_n N_X_M1001_d 0.00412982f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_278 N_VPWR_c_405_n N_X_M1008_d 0.00412982f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_M1014_d N_X_c_459_n 0.0070153f $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_280 N_VPWR_M1014_d X 6.19929e-19 $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_281 N_VPWR_M1002_s X 0.00180541f $X=1.88 $Y=1.835 $X2=0 $Y2=0
cc_282 N_VPWR_c_405_n A_656_367# 0.00309736f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_283 N_VPWR_c_405_n A_728_367# 0.00576069f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_284 N_X_c_460_n N_VGND_M1015_d 2.33864e-19 $X=1.43 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_285 N_X_c_461_n N_VGND_M1015_d 0.00211337f $X=1.185 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_286 N_X_c_462_n N_VGND_M1009_d 0.00176461f $X=2.32 $Y=1.16 $X2=0 $Y2=0
cc_287 N_X_c_460_n N_VGND_c_521_n 0.00183477f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_288 N_X_c_461_n N_VGND_c_521_n 0.016139f $X=1.185 $Y=1.16 $X2=0 $Y2=0
cc_289 N_X_c_462_n N_VGND_c_522_n 0.0170777f $X=2.32 $Y=1.16 $X2=0 $Y2=0
cc_290 N_X_c_509_p N_VGND_c_527_n 0.0135169f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_291 N_X_c_510_p N_VGND_c_529_n 0.0124525f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_292 N_X_M1003_s N_VGND_c_534_n 0.00432284f $X=1.415 $Y=0.245 $X2=0 $Y2=0
cc_293 N_X_M1011_s N_VGND_c_534_n 0.00536646f $X=2.275 $Y=0.245 $X2=0 $Y2=0
cc_294 N_X_c_509_p N_VGND_c_534_n 0.00847534f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_295 N_X_c_510_p N_VGND_c_534_n 0.00730901f $X=2.415 $Y=0.42 $X2=0 $Y2=0
