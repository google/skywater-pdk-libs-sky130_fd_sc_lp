* File: sky130_fd_sc_lp__or2b_m.spice
* Created: Wed Sep  2 10:30:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2b_m.pex.spice"
.subckt sky130_fd_sc_lp__or2b_m  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B_N_M1002_g N_A_27_496#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_224_378#_M1000_d N_A_27_496#_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_224_378#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.09975 AS=0.0588 PD=0.895 PS=0.7 NRD=32.856 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_224_378#_M1006_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.09975 PD=1.37 PS=0.895 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B_N_M1005_g N_A_27_496#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_307_378# N_A_27_496#_M1001_g N_A_224_378#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_307_378# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07455 AS=0.0441 PD=0.775 PS=0.63 NRD=35.1645 NRS=23.443 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_224_378#_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.07455 PD=1.41 PS=0.775 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__or2b_m.pxi.spice"
*
.ends
*
*
