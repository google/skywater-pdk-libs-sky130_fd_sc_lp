* File: sky130_fd_sc_lp__a22o_lp.spice
* Created: Wed Sep  2 09:22:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22o_lp.pex.spice"
.subckt sky130_fd_sc_lp__a22o_lp  VNB VPB A1 B2 B1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* B1	B1
* B2	B2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 A_225_47# N_B2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_243_409#_M1004_d N_B1_M1004_g A_225_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1008 A_389_47# N_A1_M1008_g N_A_243_409#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0588 PD=0.84 PS=0.7 NRD=44.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_389_47# VNB NSHORT L=0.15 W=0.42 AD=0.07665
+ AS=0.0882 PD=0.785 PS=0.84 NRD=24.276 NRS=44.28 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_606_47# N_A_243_409#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.07665 PD=0.66 PS=0.785 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_243_409#_M1003_g A_606_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_137_409#_M1009_d N_A1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1006 N_A_243_409#_M1006_d N_B2_M1006_g N_A_137_409#_M1009_d VPB PHIGHVT L=0.25
+ W=1 AD=0.2925 AS=0.14 PD=1.585 PS=1.28 NRD=60.0653 NRS=0 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1000 N_A_137_409#_M1000_d N_B1_M1000_g N_A_243_409#_M1006_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.2925 PD=1.28 PS=1.585 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_137_409#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.255 AS=0.14 PD=1.51 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1010 N_X_M1010_d N_A_243_409#_M1010_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.255 PD=2.57 PS=1.51 NRD=0 NRS=45.2903 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a22o_lp.pxi.spice"
*
.ends
*
*
