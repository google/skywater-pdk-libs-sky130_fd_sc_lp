# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux2_m
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__mux2_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.445000 1.765000 1.775000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 0.265000 2.465000 0.435000 ;
        RECT 2.295000 0.435000 2.465000 1.835000 ;
        RECT 2.295000 1.835000 2.725000 2.165000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.365000 2.015000 1.620000 2.345000 ;
        RECT 1.450000 2.345000 1.620000 2.895000 ;
        RECT 1.450000 2.895000 2.660000 3.065000 ;
        RECT 2.490000 2.345000 3.365000 2.490000 ;
        RECT 2.490000 2.490000 3.205000 2.515000 ;
        RECT 2.490000 2.515000 2.660000 2.895000 ;
        RECT 3.035000 1.580000 3.365000 2.345000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.231000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.585000 0.610000 0.915000 ;
        RECT 0.155000 0.915000 0.325000 2.530000 ;
        RECT 0.155000 2.530000 0.760000 2.860000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.695000  1.095000 2.115000 1.265000 ;
      RECT 0.695000  1.265000 0.865000 2.015000 ;
      RECT 0.790000  0.085000 1.120000 0.875000 ;
      RECT 0.940000  2.675000 1.270000 3.245000 ;
      RECT 1.640000  0.795000 1.970000 1.095000 ;
      RECT 1.945000  1.265000 2.115000 2.525000 ;
      RECT 1.945000  2.525000 2.310000 2.715000 ;
      RECT 2.645000  0.085000 2.975000 0.875000 ;
      RECT 2.655000  1.155000 3.720000 1.325000 ;
      RECT 2.655000  1.325000 2.825000 1.485000 ;
      RECT 2.880000  2.695000 3.210000 3.245000 ;
      RECT 3.240000  0.795000 3.570000 1.155000 ;
      RECT 3.390000  2.670000 3.720000 2.880000 ;
      RECT 3.550000  1.325000 3.720000 2.670000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2_m
END LIBRARY
