* File: sky130_fd_sc_lp__and2b_lp.pex.spice
* Created: Wed Sep  2 09:31:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2B_LP%A_108_127# 1 2 7 9 12 14 16 20 22 23 24 25
+ 30 33 38
c69 38 0 8.07371e-20 $X=1.005 $Y=1.46
r70 34 36 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.615 $Y=1.46
+ $X2=0.75 $Y2=1.46
r71 28 30 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.18 $Y=1.255
+ $X2=2.18 $Y2=1.135
r72 24 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=2.415
+ $X2=1.75 $Y2=2.415
r73 24 25 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.585 $Y=2.415
+ $X2=1.08 $Y2=2.415
r74 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=1.34
+ $X2=2.18 $Y2=1.255
r75 22 23 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.015 $Y=1.34 $X2=1.08
+ $Y2=1.34
r76 21 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.915 $Y=1.46
+ $X2=1.005 $Y2=1.46
r77 21 36 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.46
+ $X2=0.75 $Y2=1.46
r78 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=1.46 $X2=0.915 $Y2=1.46
r79 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.915 $Y=2.33
+ $X2=1.08 $Y2=2.415
r80 18 20 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.915 $Y=2.33
+ $X2=0.915 $Y2=1.46
r81 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.915 $Y=1.425
+ $X2=1.08 $Y2=1.34
r82 17 20 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.915 $Y=1.425
+ $X2=0.915 $Y2=1.46
r83 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.295
+ $X2=1.005 $Y2=1.46
r84 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=1.295
+ $X2=1.005 $Y2=0.975
r85 10 36 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.75 $Y=1.625
+ $X2=0.75 $Y2=1.46
r86 10 12 241 $w=2.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.75 $Y=1.625 $X2=0.75
+ $Y2=2.595
r87 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.46
r88 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=0.975
r89 2 33 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=1.61
+ $Y=2.095 $X2=1.75 $Y2=2.495
r90 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.925 $X2=2.18 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_LP%B 3 7 9 12 13
c39 13 0 8.07371e-20 $X=1.485 $Y=1.77
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.77
+ $X2=1.485 $Y2=1.605
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.485
+ $Y=1.77 $X2=1.485 $Y2=1.77
r42 9 13 6.67286 $w=4.73e-07 $l=2.65e-07 $layer=LI1_cond $X=1.557 $Y=2.035
+ $X2=1.557 $Y2=1.77
r43 7 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.49 $Y=0.975
+ $X2=1.49 $Y2=1.605
r44 1 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.935
+ $X2=1.485 $Y2=1.77
r45 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.485 $Y=1.935
+ $X2=1.485 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_LP%A_378_159# 1 2 9 13 15 18 22 25 26 28
c52 9 0 1.91655e-19 $X=1.965 $Y=1.135
r53 31 33 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.965 $Y=1.77
+ $X2=2.015 $Y2=1.77
r54 28 30 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.08 $Y=0.445
+ $X2=3.08 $Y2=0.675
r55 25 26 6.46576 $w=2.5e-07 $l=2.29063e-07 $layer=LI1_cond $X=3.16 $Y=1.605
+ $X2=3.007 $Y2=1.77
r56 25 30 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.16 $Y=1.605
+ $X2=3.16 $Y2=0.675
r57 20 26 6.46576 $w=2.5e-07 $l=1.9775e-07 $layer=LI1_cond $X=2.935 $Y=1.935
+ $X2=3.007 $Y2=1.77
r58 20 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.935 $Y=1.935
+ $X2=2.935 $Y2=2.24
r59 18 33 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.14 $Y=1.77
+ $X2=2.015 $Y2=1.77
r60 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.77 $X2=2.14 $Y2=1.77
r61 15 26 0.364692 $w=3.3e-07 $l=2.37e-07 $layer=LI1_cond $X=2.77 $Y=1.77
+ $X2=3.007 $Y2=1.77
r62 15 17 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.77 $Y=1.77
+ $X2=2.14 $Y2=1.77
r63 11 33 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=1.935
+ $X2=2.015 $Y2=1.77
r64 11 13 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.015 $Y=1.935
+ $X2=2.015 $Y2=2.595
r65 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.605
+ $X2=1.965 $Y2=1.77
r66 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.965 $Y=1.605 $X2=1.965
+ $Y2=1.135
r67 2 22 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.795
+ $Y=2.095 $X2=2.935 $Y2=2.24
r68 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_LP%A_N 3 7 11 13 20 21
c36 20 0 1.91655e-19 $X=2.69 $Y=1.2
r37 19 21 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.69 $Y=1.2
+ $X2=2.865 $Y2=1.2
r38 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.2 $X2=2.69 $Y2=1.2
r39 17 19 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.67 $Y=1.2 $X2=2.69
+ $Y2=1.2
r40 15 17 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.475 $Y=1.2
+ $X2=2.67 $Y2=1.2
r41 13 20 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.69 $Y=1.295
+ $X2=2.69 $Y2=1.2
r42 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.035
+ $X2=2.865 $Y2=1.2
r43 9 11 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.865 $Y=1.035
+ $X2=2.865 $Y2=0.445
r44 5 17 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.365
+ $X2=2.67 $Y2=1.2
r45 5 7 305.598 $w=2.5e-07 $l=1.23e-06 $layer=POLY_cond $X=2.67 $Y=1.365
+ $X2=2.67 $Y2=2.595
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.475 $Y=1.035
+ $X2=2.475 $Y2=1.2
r47 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.475 $Y=1.035
+ $X2=2.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_LP%X 1 2 7 8 9 10 11 12 13
r14 12 13 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.347 $Y=2.405
+ $X2=0.347 $Y2=2.775
r15 12 35 4.2731 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.347 $Y=2.405
+ $X2=0.347 $Y2=2.24
r16 11 35 5.30901 $w=4.43e-07 $l=2.05e-07 $layer=LI1_cond $X=0.347 $Y=2.035
+ $X2=0.347 $Y2=2.24
r17 10 11 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.347 $Y=1.665
+ $X2=0.347 $Y2=2.035
r18 9 10 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.347 $Y=1.295
+ $X2=0.347 $Y2=1.665
r19 9 27 8.28723 $w=4.43e-07 $l=3.2e-07 $layer=LI1_cond $X=0.347 $Y=1.295
+ $X2=0.347 $Y2=0.975
r20 8 27 1.29488 $w=4.43e-07 $l=5e-08 $layer=LI1_cond $X=0.347 $Y=0.925
+ $X2=0.347 $Y2=0.975
r21 7 8 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.347 $Y=0.555
+ $X2=0.347 $Y2=0.925
r22 2 35 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.34
+ $Y=2.095 $X2=0.485 $Y2=2.24
r23 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.765 $X2=0.4 $Y2=0.975
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_LP%VPWR 1 2 9 13 16 17 18 24 30 31 34
r44 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.28 $Y2=3.33
r48 28 30 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.28 $Y2=3.33
r51 24 26 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 16 21 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=1.015 $Y2=3.33
r58 15 26 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.18 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=3.33
+ $X2=1.015 $Y2=3.33
r60 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=3.33
r61 11 13 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=2.28
r62 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=3.245
+ $X2=1.015 $Y2=3.33
r63 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.015 $Y=3.245
+ $X2=1.015 $Y2=2.895
r64 2 13 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=2.14
+ $Y=2.095 $X2=2.28 $Y2=2.28
r65 1 9 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=0.875
+ $Y=2.095 $X2=1.015 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_LP%VGND 1 2 9 11 15 17 19 26 27 30 33
r36 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r37 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r39 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.26
+ $Y2=0
r41 24 26 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=3.12
+ $Y2=0
r42 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r43 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r45 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.72
+ $Y2=0
r46 17 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r47 17 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r48 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0
r49 13 15 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0.445
r50 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r51 11 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.26
+ $Y2=0
r52 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=1.385
+ $Y2=0
r53 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085 $X2=1.22
+ $Y2=0
r54 7 9 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.91
r55 2 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.26 $Y2=0.445
r56 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.765 $X2=1.22 $Y2=0.91
.ends

