* File: sky130_fd_sc_lp__o32a_m.pxi.spice
* Created: Fri Aug 28 11:17:51 2020
* 
x_PM_SKY130_FD_SC_LP__O32A_M%A1 N_A1_c_77_n N_A1_M1009_g N_A1_M1000_g
+ N_A1_c_79_n A1 A1 A1 N_A1_c_81_n N_A1_c_82_n PM_SKY130_FD_SC_LP__O32A_M%A1
x_PM_SKY130_FD_SC_LP__O32A_M%A2 N_A2_M1006_g N_A2_M1002_g N_A2_c_113_n
+ N_A2_c_118_n A2 A2 A2 A2 N_A2_c_115_n PM_SKY130_FD_SC_LP__O32A_M%A2
x_PM_SKY130_FD_SC_LP__O32A_M%A_86_55# N_A_86_55#_M1008_d N_A_86_55#_M1001_d
+ N_A_86_55#_M1005_g N_A_86_55#_M1011_g N_A_86_55#_c_156_n N_A_86_55#_c_157_n
+ N_A_86_55#_c_158_n N_A_86_55#_c_159_n N_A_86_55#_c_160_n N_A_86_55#_c_161_n
+ N_A_86_55#_c_162_n N_A_86_55#_c_153_n N_A_86_55#_c_154_n
+ PM_SKY130_FD_SC_LP__O32A_M%A_86_55#
x_PM_SKY130_FD_SC_LP__O32A_M%A3 N_A3_M1001_g N_A3_M1004_g N_A3_c_224_n
+ N_A3_c_229_n A3 A3 A3 A3 N_A3_c_226_n PM_SKY130_FD_SC_LP__O32A_M%A3
x_PM_SKY130_FD_SC_LP__O32A_M%B2 N_B2_M1008_g N_B2_M1010_g N_B2_c_271_n
+ N_B2_c_272_n B2 N_B2_c_273_n PM_SKY130_FD_SC_LP__O32A_M%B2
x_PM_SKY130_FD_SC_LP__O32A_M%B1 N_B1_M1007_g N_B1_M1003_g B1 B1 B1 N_B1_c_315_n
+ N_B1_c_316_n PM_SKY130_FD_SC_LP__O32A_M%B1
x_PM_SKY130_FD_SC_LP__O32A_M%X N_X_M1005_s N_X_M1011_s N_X_c_344_n X X X X X X X
+ N_X_c_346_n PM_SKY130_FD_SC_LP__O32A_M%X
x_PM_SKY130_FD_SC_LP__O32A_M%VPWR N_VPWR_M1011_d N_VPWR_M1003_d N_VPWR_c_356_n
+ N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n VPWR N_VPWR_c_360_n
+ N_VPWR_c_361_n N_VPWR_c_355_n N_VPWR_c_363_n PM_SKY130_FD_SC_LP__O32A_M%VPWR
x_PM_SKY130_FD_SC_LP__O32A_M%VGND N_VGND_M1005_d N_VGND_M1002_d N_VGND_c_398_n
+ N_VGND_c_399_n N_VGND_c_400_n VGND N_VGND_c_401_n N_VGND_c_402_n
+ N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n PM_SKY130_FD_SC_LP__O32A_M%VGND
x_PM_SKY130_FD_SC_LP__O32A_M%A_249_81# N_A_249_81#_M1009_d N_A_249_81#_M1004_d
+ N_A_249_81#_M1007_d N_A_249_81#_c_443_n N_A_249_81#_c_438_n
+ N_A_249_81#_c_439_n N_A_249_81#_c_452_n N_A_249_81#_c_440_n
+ N_A_249_81#_c_441_n N_A_249_81#_c_442_n PM_SKY130_FD_SC_LP__O32A_M%A_249_81#
cc_1 VNB N_A1_c_77_n 0.0208333f $X=-0.19 $Y=-0.245 $X2=1.057 $Y2=1.418
cc_2 VNB N_A1_M1000_g 0.0025853f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=2.225
cc_3 VNB N_A1_c_79_n 0.0195561f $X=-0.19 $Y=-0.245 $X2=1.057 $Y2=1.605
cc_4 VNB A1 0.0138653f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_5 VNB N_A1_c_81_n 0.0200875f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.1
cc_6 VNB N_A1_c_82_n 0.0180293f $X=-0.19 $Y=-0.245 $X2=1.057 $Y2=0.935
cc_7 VNB N_A2_M1002_g 0.0309669f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=2.225
cc_8 VNB N_A2_c_113_n 0.0207732f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_9 VNB A2 8.52225e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_A2_c_115_n 0.0162062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_86_55#_M1005_g 0.0628108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_86_55#_c_153_n 0.00470503f $X=-0.19 $Y=-0.245 $X2=0.877 $Y2=1.665
cc_13 VNB N_A_86_55#_c_154_n 0.00778131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A3_M1004_g 0.031622f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=2.225
cc_15 VNB N_A3_c_224_n 0.0207436f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_16 VNB A3 9.47981e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_A3_c_226_n 0.0162166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B2_M1008_g 0.0244024f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.935
cc_19 VNB N_B2_c_271_n 0.0230023f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_20 VNB N_B2_c_272_n 0.00307126f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_21 VNB N_B2_c_273_n 0.0164398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_M1003_g 0.0023723f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.605
cc_23 VNB B1 0.0347228f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=2.225
cc_24 VNB N_B1_c_315_n 0.0923772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_316_n 0.0181703f $X=-0.19 $Y=-0.245 $X2=1.057 $Y2=1.1
cc_26 VNB X 0.0120316f $X=-0.19 $Y=-0.245 $X2=1.057 $Y2=1.605
cc_27 VNB X 0.0404818f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_28 VNB N_VPWR_c_355_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_398_n 0.00946249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_399_n 0.0232186f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_31 VNB N_VGND_c_400_n 0.00886846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_401_n 0.0189723f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.1
cc_33 VNB N_VGND_c_402_n 0.0495508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_403_n 0.247564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_404_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_405_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_249_81#_c_438_n 0.0272967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_249_81#_c_439_n 0.0077309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_249_81#_c_440_n 0.00538595f $X=-0.19 $Y=-0.245 $X2=1.057 $Y2=0.935
cc_40 VNB N_A_249_81#_c_441_n 0.00285871f $X=-0.19 $Y=-0.245 $X2=0.877 $Y2=0.925
cc_41 VNB N_A_249_81#_c_442_n 0.0186746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A1_M1000_g 0.0318731f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.225
cc_43 VPB A1 0.0123809f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_44 VPB N_A2_M1006_g 0.0183328f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=0.935
cc_45 VPB N_A2_c_113_n 0.00232332f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_46 VPB N_A2_c_118_n 0.0169723f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_47 VPB A2 0.00281222f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_48 VPB N_A_86_55#_M1005_g 0.0585746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_86_55#_c_156_n 0.127187f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_50 VPB N_A_86_55#_c_157_n 0.0151863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_86_55#_c_158_n 0.00820249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_86_55#_c_159_n 0.0536747f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=1.1
cc_53 VPB N_A_86_55#_c_160_n 0.00464443f $X=-0.19 $Y=1.655 $X2=1.057 $Y2=0.935
cc_54 VPB N_A_86_55#_c_161_n 0.0155586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_86_55#_c_162_n 0.0066127f $X=-0.19 $Y=1.655 $X2=0.877 $Y2=1.1
cc_56 VPB N_A_86_55#_c_153_n 0.00200071f $X=-0.19 $Y=1.655 $X2=0.877 $Y2=1.665
cc_57 VPB N_A3_M1001_g 0.0209964f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=0.935
cc_58 VPB N_A3_c_224_n 0.00232001f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_59 VPB N_A3_c_229_n 0.019037f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_60 VPB A3 0.002464f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_61 VPB N_B2_M1010_g 0.0257111f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.225
cc_62 VPB N_B2_c_272_n 0.0127254f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_63 VPB N_B1_M1003_g 0.037758f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.605
cc_64 VPB B1 0.0123155f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.225
cc_65 VPB N_X_c_344_n 0.00434092f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.225
cc_66 VPB X 0.0215161f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_67 VPB N_X_c_346_n 0.0308029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_356_n 0.0212619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_357_n 0.0534117f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_70 VPB N_VPWR_c_358_n 0.0682373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_359_n 0.00632158f $X=-0.19 $Y=1.655 $X2=1.057 $Y2=1.1
cc_72 VPB N_VPWR_c_360_n 0.0187155f $X=-0.19 $Y=1.655 $X2=1.057 $Y2=0.935
cc_73 VPB N_VPWR_c_361_n 0.0120081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_355_n 0.0772566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_363_n 0.00583335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 A1 N_A2_M1002_g 9.93013e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_77 N_A1_c_82_n N_A2_M1002_g 0.02507f $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_78 N_A1_c_79_n N_A2_c_113_n 0.0282323f $X=1.057 $Y=1.605 $X2=0 $Y2=0
cc_79 N_A1_M1000_g N_A2_c_118_n 0.0282323f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_80 N_A1_c_77_n A2 0.00526781f $X=1.057 $Y=1.418 $X2=0 $Y2=0
cc_81 A1 A2 0.0206266f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_82 N_A1_c_77_n N_A2_c_115_n 0.0282323f $X=1.057 $Y=1.418 $X2=0 $Y2=0
cc_83 A1 N_A2_c_115_n 0.00169671f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A1_M1000_g N_A_86_55#_M1005_g 0.0176019f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_85 A1 N_A_86_55#_M1005_g 0.0100897f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A1_c_81_n N_A_86_55#_M1005_g 0.0256483f $X=1.035 $Y=1.1 $X2=0 $Y2=0
cc_87 N_A1_c_82_n N_A_86_55#_M1005_g 0.00952063f $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_88 N_A1_M1000_g N_A_86_55#_c_156_n 0.00564446f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_89 A1 X 0.0489424f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A1_M1000_g N_VPWR_c_356_n 0.00586908f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_91 A1 N_VPWR_c_356_n 0.0125156f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A1_M1000_g N_VPWR_c_355_n 8.50146e-19 $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_93 A1 N_VGND_c_398_n 0.0223879f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_94 N_A1_c_81_n N_VGND_c_398_n 2.09235e-19 $X=1.035 $Y=1.1 $X2=0 $Y2=0
cc_95 N_A1_c_82_n N_VGND_c_398_n 0.0075344f $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_96 N_A1_c_82_n N_VGND_c_399_n 0.00552345f $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_97 N_A1_c_82_n N_VGND_c_400_n 0.00110481f $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_98 A1 N_VGND_c_403_n 0.0094001f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_99 N_A1_c_82_n N_VGND_c_403_n 0.00534666f $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_100 N_A1_c_82_n N_A_249_81#_c_443_n 2.03427e-19 $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_101 A1 N_A_249_81#_c_439_n 0.0136485f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 N_A1_c_82_n N_A_249_81#_c_439_n 0.00158972f $X=1.057 $Y=0.935 $X2=0 $Y2=0
cc_103 N_A2_M1006_g N_A_86_55#_c_156_n 0.00526169f $X=1.53 $Y=2.225 $X2=0 $Y2=0
cc_104 A2 N_A_86_55#_c_156_n 0.00513767f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A2_M1006_g N_A3_M1001_g 0.0192051f $X=1.53 $Y=2.225 $X2=0 $Y2=0
cc_106 A2 N_A3_M1001_g 0.00481612f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A2_M1002_g N_A3_M1004_g 0.0156078f $X=1.6 $Y=0.615 $X2=0 $Y2=0
cc_108 N_A2_c_113_n N_A3_c_224_n 0.0138171f $X=1.62 $Y=1.69 $X2=0 $Y2=0
cc_109 N_A2_c_118_n N_A3_c_229_n 0.0138171f $X=1.62 $Y=1.855 $X2=0 $Y2=0
cc_110 N_A2_M1006_g A3 5.96081e-19 $X=1.53 $Y=2.225 $X2=0 $Y2=0
cc_111 A2 A3 0.0577896f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_112 N_A2_c_115_n A3 0.00209845f $X=1.62 $Y=1.35 $X2=0 $Y2=0
cc_113 A2 N_A3_c_226_n 0.00239472f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_114 N_A2_c_115_n N_A3_c_226_n 0.0138171f $X=1.62 $Y=1.35 $X2=0 $Y2=0
cc_115 A2 N_VPWR_c_356_n 0.00827328f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A2_M1006_g N_VPWR_c_355_n 8.50146e-19 $X=1.53 $Y=2.225 $X2=0 $Y2=0
cc_117 A2 N_VPWR_c_355_n 0.00785601f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_118 A2 A_321_403# 0.00464229f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_119 N_A2_M1002_g N_VGND_c_399_n 0.00532616f $X=1.6 $Y=0.615 $X2=0 $Y2=0
cc_120 N_A2_M1002_g N_VGND_c_400_n 0.00721488f $X=1.6 $Y=0.615 $X2=0 $Y2=0
cc_121 N_A2_M1002_g N_VGND_c_403_n 0.00520409f $X=1.6 $Y=0.615 $X2=0 $Y2=0
cc_122 N_A2_M1002_g N_A_249_81#_c_443_n 2.08812e-19 $X=1.6 $Y=0.615 $X2=0 $Y2=0
cc_123 N_A2_M1002_g N_A_249_81#_c_438_n 0.0125344f $X=1.6 $Y=0.615 $X2=0 $Y2=0
cc_124 A2 N_A_249_81#_c_438_n 0.0169211f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A2_c_115_n N_A_249_81#_c_438_n 0.00288634f $X=1.62 $Y=1.35 $X2=0 $Y2=0
cc_126 N_A2_c_115_n N_A_249_81#_c_439_n 0.00160691f $X=1.62 $Y=1.35 $X2=0 $Y2=0
cc_127 N_A_86_55#_c_156_n N_A3_M1001_g 0.00412554f $X=2.11 $Y=3.03 $X2=0 $Y2=0
cc_128 N_A_86_55#_c_159_n N_A3_M1001_g 0.00233074f $X=2.275 $Y=2.94 $X2=0 $Y2=0
cc_129 N_A_86_55#_c_160_n N_A3_M1001_g 0.00124165f $X=2.53 $Y=2.23 $X2=0 $Y2=0
cc_130 N_A_86_55#_c_161_n N_A3_M1001_g 0.00237626f $X=2.53 $Y=2.29 $X2=0 $Y2=0
cc_131 N_A_86_55#_M1001_d A3 0.00406328f $X=2.145 $Y=2.015 $X2=0 $Y2=0
cc_132 N_A_86_55#_c_158_n A3 0.00511521f $X=2.425 $Y=2.94 $X2=0 $Y2=0
cc_133 N_A_86_55#_c_159_n A3 0.00236986f $X=2.275 $Y=2.94 $X2=0 $Y2=0
cc_134 N_A_86_55#_c_160_n A3 0.0241621f $X=2.53 $Y=2.23 $X2=0 $Y2=0
cc_135 N_A_86_55#_c_161_n A3 0.0185063f $X=2.53 $Y=2.29 $X2=0 $Y2=0
cc_136 N_A_86_55#_c_153_n N_B2_M1008_g 0.00180664f $X=3.13 $Y=1.875 $X2=0 $Y2=0
cc_137 N_A_86_55#_c_154_n N_B2_M1008_g 0.00706699f $X=2.895 $Y=0.7 $X2=0 $Y2=0
cc_138 N_A_86_55#_c_161_n N_B2_M1010_g 0.00203086f $X=2.53 $Y=2.29 $X2=0 $Y2=0
cc_139 N_A_86_55#_c_162_n N_B2_M1010_g 0.0147797f $X=3.045 $Y=1.96 $X2=0 $Y2=0
cc_140 N_A_86_55#_c_153_n N_B2_M1010_g 0.00190405f $X=3.13 $Y=1.875 $X2=0 $Y2=0
cc_141 N_A_86_55#_c_160_n N_B2_c_272_n 0.00297157f $X=2.53 $Y=2.23 $X2=0 $Y2=0
cc_142 N_A_86_55#_c_162_n N_B2_c_272_n 0.00229679f $X=3.045 $Y=1.96 $X2=0 $Y2=0
cc_143 N_A_86_55#_c_160_n B2 0.00827856f $X=2.53 $Y=2.23 $X2=0 $Y2=0
cc_144 N_A_86_55#_c_162_n B2 0.0165246f $X=3.045 $Y=1.96 $X2=0 $Y2=0
cc_145 N_A_86_55#_c_153_n B2 0.0366424f $X=3.13 $Y=1.875 $X2=0 $Y2=0
cc_146 N_A_86_55#_c_154_n B2 0.010617f $X=2.895 $Y=0.7 $X2=0 $Y2=0
cc_147 N_A_86_55#_c_153_n N_B2_c_273_n 0.00591755f $X=3.13 $Y=1.875 $X2=0 $Y2=0
cc_148 N_A_86_55#_c_154_n N_B2_c_273_n 0.00322853f $X=2.895 $Y=0.7 $X2=0 $Y2=0
cc_149 N_A_86_55#_c_162_n N_B1_M1003_g 0.0176949f $X=3.045 $Y=1.96 $X2=0 $Y2=0
cc_150 N_A_86_55#_c_153_n N_B1_M1003_g 0.00947143f $X=3.13 $Y=1.875 $X2=0 $Y2=0
cc_151 N_A_86_55#_c_153_n B1 0.0508193f $X=3.13 $Y=1.875 $X2=0 $Y2=0
cc_152 N_A_86_55#_c_154_n B1 0.0124755f $X=2.895 $Y=0.7 $X2=0 $Y2=0
cc_153 N_A_86_55#_c_153_n N_B1_c_315_n 0.0178117f $X=3.13 $Y=1.875 $X2=0 $Y2=0
cc_154 N_A_86_55#_c_154_n N_B1_c_315_n 0.00288281f $X=2.895 $Y=0.7 $X2=0 $Y2=0
cc_155 N_A_86_55#_c_154_n N_B1_c_316_n 0.00679195f $X=2.895 $Y=0.7 $X2=0 $Y2=0
cc_156 N_A_86_55#_M1005_g X 0.0346178f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_157 N_A_86_55#_M1005_g N_X_c_346_n 0.00972466f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_158 N_A_86_55#_M1005_g N_VPWR_c_356_n 0.0203197f $X=0.505 $Y=0.615 $X2=0
+ $Y2=0
cc_159 N_A_86_55#_c_156_n N_VPWR_c_356_n 0.0255805f $X=2.11 $Y=3.03 $X2=0 $Y2=0
cc_160 N_A_86_55#_c_157_n N_VPWR_c_356_n 0.00583501f $X=0.58 $Y=3.03 $X2=0 $Y2=0
cc_161 N_A_86_55#_c_158_n N_VPWR_c_357_n 0.00638735f $X=2.425 $Y=2.94 $X2=0
+ $Y2=0
cc_162 N_A_86_55#_c_161_n N_VPWR_c_357_n 0.0169548f $X=2.53 $Y=2.29 $X2=0 $Y2=0
cc_163 N_A_86_55#_c_162_n N_VPWR_c_357_n 0.00105058f $X=3.045 $Y=1.96 $X2=0
+ $Y2=0
cc_164 N_A_86_55#_c_156_n N_VPWR_c_358_n 0.0403394f $X=2.11 $Y=3.03 $X2=0 $Y2=0
cc_165 N_A_86_55#_c_158_n N_VPWR_c_358_n 0.0259503f $X=2.425 $Y=2.94 $X2=0 $Y2=0
cc_166 N_A_86_55#_c_157_n N_VPWR_c_360_n 0.0045659f $X=0.58 $Y=3.03 $X2=0 $Y2=0
cc_167 N_A_86_55#_c_156_n N_VPWR_c_355_n 0.0521462f $X=2.11 $Y=3.03 $X2=0 $Y2=0
cc_168 N_A_86_55#_c_157_n N_VPWR_c_355_n 0.00904332f $X=0.58 $Y=3.03 $X2=0 $Y2=0
cc_169 N_A_86_55#_c_158_n N_VPWR_c_355_n 0.017886f $X=2.425 $Y=2.94 $X2=0 $Y2=0
cc_170 N_A_86_55#_c_159_n N_VPWR_c_355_n 0.00783053f $X=2.275 $Y=2.94 $X2=0
+ $Y2=0
cc_171 N_A_86_55#_c_162_n A_566_403# 0.00499838f $X=3.045 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_86_55#_M1005_g N_VGND_c_398_n 0.0118585f $X=0.505 $Y=0.615 $X2=0
+ $Y2=0
cc_173 N_A_86_55#_M1005_g N_VGND_c_401_n 0.00532616f $X=0.505 $Y=0.615 $X2=0
+ $Y2=0
cc_174 N_A_86_55#_M1005_g N_VGND_c_403_n 0.00520409f $X=0.505 $Y=0.615 $X2=0
+ $Y2=0
cc_175 N_A_86_55#_c_154_n N_A_249_81#_c_438_n 0.0141649f $X=2.895 $Y=0.7 $X2=0
+ $Y2=0
cc_176 N_A_86_55#_c_154_n N_A_249_81#_c_452_n 0.00822286f $X=2.895 $Y=0.7 $X2=0
+ $Y2=0
cc_177 N_A_86_55#_M1008_d N_A_249_81#_c_440_n 0.0022017f $X=2.755 $Y=0.405 $X2=0
+ $Y2=0
cc_178 N_A_86_55#_c_154_n N_A_249_81#_c_440_n 0.0207309f $X=2.895 $Y=0.7 $X2=0
+ $Y2=0
cc_179 N_A3_M1004_g N_B2_M1008_g 0.020186f $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_180 N_A3_M1001_g N_B2_M1010_g 0.00868461f $X=2.07 $Y=2.225 $X2=0 $Y2=0
cc_181 N_A3_c_229_n N_B2_M1010_g 0.00302414f $X=2.16 $Y=1.855 $X2=0 $Y2=0
cc_182 A3 N_B2_M1010_g 0.00181231f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A3_c_226_n N_B2_c_271_n 0.0141576f $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_184 N_A3_c_224_n N_B2_c_272_n 0.0141576f $X=2.16 $Y=1.69 $X2=0 $Y2=0
cc_185 A3 B2 0.0236701f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A3_c_226_n B2 0.00187834f $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_187 N_A3_M1004_g N_B2_c_273_n 0.0141576f $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_188 A3 N_B2_c_273_n 0.00205361f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A3_M1001_g N_VPWR_c_355_n 6.49005e-19 $X=2.07 $Y=2.225 $X2=0 $Y2=0
cc_190 A3 N_VPWR_c_355_n 0.00154013f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A3_M1004_g N_VGND_c_400_n 0.00394976f $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_192 N_A3_M1004_g N_VGND_c_402_n 0.00552345f $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_193 N_A3_M1004_g N_VGND_c_403_n 0.00534666f $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_194 N_A3_M1004_g N_A_249_81#_c_438_n 0.0148305f $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_195 A3 N_A_249_81#_c_438_n 0.0125942f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A3_c_226_n N_A_249_81#_c_438_n 0.0040064f $X=2.16 $Y=1.35 $X2=0 $Y2=0
cc_197 N_A3_M1004_g N_A_249_81#_c_452_n 5.59817e-19 $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_198 N_A3_M1004_g N_A_249_81#_c_441_n 0.00158151f $X=2.25 $Y=0.615 $X2=0 $Y2=0
cc_199 N_B2_M1010_g N_B1_M1003_g 0.0397523f $X=2.755 $Y=2.225 $X2=0 $Y2=0
cc_200 N_B2_c_271_n N_B1_M1003_g 0.0209512f $X=2.7 $Y=1.61 $X2=0 $Y2=0
cc_201 B2 N_B1_c_315_n 5.98591e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_202 N_B2_c_273_n N_B1_c_315_n 0.0209512f $X=2.7 $Y=1.27 $X2=0 $Y2=0
cc_203 N_B2_M1008_g N_B1_c_316_n 0.0188218f $X=2.68 $Y=0.615 $X2=0 $Y2=0
cc_204 N_B2_M1010_g N_VPWR_c_357_n 9.99969e-19 $X=2.755 $Y=2.225 $X2=0 $Y2=0
cc_205 N_B2_M1010_g N_VPWR_c_358_n 0.00297774f $X=2.755 $Y=2.225 $X2=0 $Y2=0
cc_206 N_B2_M1010_g N_VPWR_c_355_n 0.00400849f $X=2.755 $Y=2.225 $X2=0 $Y2=0
cc_207 N_B2_M1008_g N_VGND_c_402_n 9.29198e-19 $X=2.68 $Y=0.615 $X2=0 $Y2=0
cc_208 N_B2_M1008_g N_A_249_81#_c_438_n 0.00140499f $X=2.68 $Y=0.615 $X2=0 $Y2=0
cc_209 B2 N_A_249_81#_c_438_n 0.00117071f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_210 N_B2_c_273_n N_A_249_81#_c_438_n 4.62881e-19 $X=2.7 $Y=1.27 $X2=0 $Y2=0
cc_211 N_B2_M1008_g N_A_249_81#_c_452_n 4.02684e-19 $X=2.68 $Y=0.615 $X2=0 $Y2=0
cc_212 N_B2_M1008_g N_A_249_81#_c_440_n 0.0134613f $X=2.68 $Y=0.615 $X2=0 $Y2=0
cc_213 N_B1_M1003_g N_VPWR_c_357_n 0.00993911f $X=3.15 $Y=2.225 $X2=0 $Y2=0
cc_214 B1 N_VPWR_c_357_n 0.00587178f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_215 N_B1_c_315_n N_VPWR_c_357_n 0.00498931f $X=3.48 $Y=1.1 $X2=0 $Y2=0
cc_216 N_B1_M1003_g N_VPWR_c_358_n 0.00247589f $X=3.15 $Y=2.225 $X2=0 $Y2=0
cc_217 N_B1_M1003_g N_VPWR_c_355_n 0.00336713f $X=3.15 $Y=2.225 $X2=0 $Y2=0
cc_218 N_B1_c_316_n N_VGND_c_402_n 9.29198e-19 $X=3.36 $Y=0.935 $X2=0 $Y2=0
cc_219 B1 N_VGND_c_403_n 0.0048785f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_220 N_B1_c_316_n N_A_249_81#_c_440_n 0.0116853f $X=3.36 $Y=0.935 $X2=0 $Y2=0
cc_221 B1 N_A_249_81#_c_442_n 0.0139625f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_222 N_B1_c_315_n N_A_249_81#_c_442_n 0.00641544f $X=3.48 $Y=1.1 $X2=0 $Y2=0
cc_223 N_B1_c_316_n N_A_249_81#_c_442_n 0.00208142f $X=3.36 $Y=0.935 $X2=0 $Y2=0
cc_224 N_X_c_346_n N_VPWR_c_356_n 0.0403375f $X=0.29 $Y=2.29 $X2=0 $Y2=0
cc_225 N_X_c_346_n N_VPWR_c_360_n 0.0071358f $X=0.29 $Y=2.29 $X2=0 $Y2=0
cc_226 N_X_c_346_n N_VPWR_c_355_n 0.00813043f $X=0.29 $Y=2.29 $X2=0 $Y2=0
cc_227 X N_VGND_c_401_n 0.00654658f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_228 X N_VGND_c_403_n 0.00806527f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_229 N_VGND_c_399_n N_A_249_81#_c_443_n 0.00445248f $X=1.67 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_403_n N_A_249_81#_c_443_n 0.00613177f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_c_400_n N_A_249_81#_c_438_n 0.0227966f $X=1.835 $Y=0.55 $X2=0
+ $Y2=0
cc_232 N_VGND_c_403_n N_A_249_81#_c_438_n 0.0188632f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_402_n N_A_249_81#_c_440_n 0.0418106f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_403_n N_A_249_81#_c_440_n 0.0257833f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_400_n N_A_249_81#_c_441_n 0.00799668f $X=1.835 $Y=0.55 $X2=0
+ $Y2=0
cc_236 N_VGND_c_402_n N_A_249_81#_c_441_n 0.0128106f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_403_n N_A_249_81#_c_441_n 0.0073517f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_402_n N_A_249_81#_c_442_n 0.021223f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_403_n N_A_249_81#_c_442_n 0.0125082f $X=3.6 $Y=0 $X2=0 $Y2=0
