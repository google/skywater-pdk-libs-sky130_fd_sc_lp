* File: sky130_fd_sc_lp__o21a_1.pex.spice
* Created: Fri Aug 28 11:03:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21A_1%A_80_21# 1 2 7 9 12 14 15 16 17 20 22 24 36
r53 28 36 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.61 $Y=1.35
+ $X2=0.665 $Y2=1.35
r54 28 33 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.61 $Y=1.35
+ $X2=0.475 $Y2=1.35
r55 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.35 $X2=0.61 $Y2=1.35
r56 22 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=2.1 $X2=1.77
+ $Y2=2.015
r57 22 24 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.77 $Y=2.1 $X2=1.77
+ $Y2=2.49
r58 18 20 25.5458 $w=2.98e-07 $l=6.65e-07 $layer=LI1_cond $X=1.195 $Y=1.085
+ $X2=1.195 $Y2=0.42
r59 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=2.015
+ $X2=1.77 $Y2=2.015
r60 16 17 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.605 $Y=2.015
+ $X2=0.905 $Y2=2.015
r61 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.82 $Y=1.93
+ $X2=0.905 $Y2=2.015
r62 14 18 15.7759 $w=2.9e-07 $l=5.03115e-07 $layer=LI1_cond $X=0.82 $Y=1.385
+ $X2=1.195 $Y2=1.085
r63 14 27 8.83448 $w=2.9e-07 $l=2.1e-07 $layer=LI1_cond $X=0.82 $Y=1.385
+ $X2=0.61 $Y2=1.385
r64 14 15 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.82 $Y=1.515
+ $X2=0.82 $Y2=1.93
r65 10 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.515
+ $X2=0.665 $Y2=1.35
r66 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.665 $Y=1.515
+ $X2=0.665 $Y2=2.465
r67 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=1.35
r68 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
r69 2 32 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.835 $X2=1.77 $Y2=2.015
r70 2 24 300 $w=1.7e-07 $l=7.52712e-07 $layer=licon1_PDIFF $count=2 $X=1.56
+ $Y=1.835 $X2=1.77 $Y2=2.49
r71 1 20 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.255 $X2=1.21 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_1%B1 3 7 9 13 14
c34 13 0 2.31702e-19 $X=1.25 $Y=1.51
r35 14 15 9.06583 $w=3.19e-07 $l=6e-08 $layer=POLY_cond $X=1.425 $Y=1.51
+ $X2=1.485 $Y2=1.51
r36 12 14 26.442 $w=3.19e-07 $l=1.75e-07 $layer=POLY_cond $X=1.25 $Y=1.51
+ $X2=1.425 $Y2=1.51
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.51 $X2=1.25 $Y2=1.51
r38 9 13 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.245 $Y=1.665
+ $X2=1.245 $Y2=1.51
r39 5 15 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.675
+ $X2=1.485 $Y2=1.51
r40 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.485 $Y=1.675
+ $X2=1.485 $Y2=2.465
r41 1 14 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.51
r42 1 3 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_1%A2 3 7 9 10 14
c34 14 0 1.78149e-19 $X=1.935 $Y=1.51
c35 7 0 5.35535e-20 $X=2.025 $Y=2.465
r36 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.51
+ $X2=1.935 $Y2=1.675
r37 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.51
+ $X2=1.935 $Y2=1.345
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.51 $X2=1.935 $Y2=1.51
r39 10 15 7.74029 $w=3.33e-07 $l=2.25e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=1.935 $Y2=1.592
r40 9 15 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.935 $Y2=1.592
r41 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.025 $Y=2.465
+ $X2=2.025 $Y2=1.675
r42 3 16 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.855 $Y=0.675
+ $X2=1.855 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_1%A1 3 7 9 14 15
r25 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.46 $X2=2.59 $Y2=1.46
r26 11 14 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.385 $Y=1.46
+ $X2=2.59 $Y2=1.46
r27 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.46
r28 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.625
+ $X2=2.385 $Y2=1.46
r29 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.385 $Y=1.625
+ $X2=2.385 $Y2=2.465
r30 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.295
+ $X2=2.385 $Y2=1.46
r31 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.385 $Y=1.295
+ $X2=2.385 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_1%X 1 2 7 8 9 10 11 12 13 24 34 37
r18 35 37 1.43009 $w=4.58e-07 $l=5.5e-08 $layer=LI1_cond $X=0.315 $Y=1.925
+ $X2=0.315 $Y2=1.98
r19 34 48 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=1.665 $X2=0.22
+ $Y2=1.695
r20 13 45 3.51023 $w=4.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.315 $Y=2.775
+ $X2=0.315 $Y2=2.91
r21 12 13 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=2.405
+ $X2=0.315 $Y2=2.775
r22 11 12 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=2.035
+ $X2=0.315 $Y2=2.405
r23 11 37 1.43009 $w=4.58e-07 $l=5.5e-08 $layer=LI1_cond $X=0.315 $Y=2.035
+ $X2=0.315 $Y2=1.98
r24 10 35 5.27835 $w=4.58e-07 $l=2.03e-07 $layer=LI1_cond $X=0.315 $Y=1.722
+ $X2=0.315 $Y2=1.925
r25 10 48 2.7257 $w=4.58e-07 $l=2.7e-08 $layer=LI1_cond $X=0.315 $Y=1.722
+ $X2=0.315 $Y2=1.695
r26 10 34 1.19513 $w=2.68e-07 $l=2.8e-08 $layer=LI1_cond $X=0.22 $Y=1.637
+ $X2=0.22 $Y2=1.665
r27 9 10 14.5976 $w=2.68e-07 $l=3.42e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.637
r28 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.925 $X2=0.22
+ $Y2=1.295
r29 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.555 $X2=0.22
+ $Y2=0.925
r30 7 24 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=0.555
+ $X2=0.22 $Y2=0.42
r31 2 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.45 $Y2=2.91
r32 2 37 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.45 $Y2=1.98
r33 1 24 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_1%VPWR 1 2 11 13 15 19 21 27 33
r34 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 28 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 27 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 25 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 22 27 13.8654 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.075 $Y2=3.33
r41 22 24 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 21 32 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.657 $Y2=3.33
r43 21 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 19 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 19 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 15 18 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=2.6 $Y=2.015
+ $X2=2.6 $Y2=2.95
r47 13 32 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.657 $Y2=3.33
r48 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.6 $Y2=2.95
r49 9 27 2.92113 $w=7.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.075 $Y=3.245
+ $X2=1.075 $Y2=3.33
r50 9 11 14.1204 $w=7.18e-07 $l=8.5e-07 $layer=LI1_cond $X=1.075 $Y=3.245
+ $X2=1.075 $Y2=2.395
r51 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.835 $X2=2.6 $Y2=2.95
r52 2 15 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=2.46 $Y=1.835
+ $X2=2.6 $Y2=2.015
r53 1 11 150 $w=1.7e-07 $l=7.81281e-07 $layer=licon1_PDIFF $count=4 $X=0.74
+ $Y=1.835 $X2=1.27 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.12
+ $Y2=0
r39 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.64
+ $Y2=0
r40 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r42 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r43 23 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.68
+ $Y2=0
r44 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=2.12
+ $Y2=0
r45 22 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.68
+ $Y2=0
r46 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r49 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r50 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r51 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r52 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0
r53 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0.4
r54 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r55 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r56 2 13 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.255 $X2=2.12 $Y2=0.4
r57 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_1%A_300_51# 1 2 9 11 12 15
r26 13 15 22.4912 $w=3.08e-07 $l=6.05e-07 $layer=LI1_cond $X=2.61 $Y=1.025
+ $X2=2.61 $Y2=0.42
r27 11 13 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.455 $Y=1.11
+ $X2=2.61 $Y2=1.025
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.455 $Y=1.11
+ $X2=1.785 $Y2=1.11
r29 7 12 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.65 $Y=1.025
+ $X2=1.785 $Y2=1.11
r30 7 9 25.8233 $w=2.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.65 $Y=1.025
+ $X2=1.65 $Y2=0.42
r31 2 15 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.46
+ $Y=0.255 $X2=2.6 $Y2=0.42
r32 1 9 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.255 $X2=1.64 $Y2=0.42
.ends

