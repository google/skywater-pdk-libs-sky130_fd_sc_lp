* File: sky130_fd_sc_lp__nand3b_1.pex.spice
* Created: Fri Aug 28 10:49:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3B_1%A_N 3 7 9 12 13
c28 13 0 1.92174e-19 $X=0.67 $Y=1.51
r29 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=1.51
+ $X2=0.67 $Y2=1.675
r30 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=1.51
+ $X2=0.67 $Y2=1.345
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.51 $X2=0.67 $Y2=1.51
r32 9 13 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.69 $Y=1.665
+ $X2=0.69 $Y2=1.51
r33 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.76 $Y=2.045
+ $X2=0.76 $Y2=1.675
r34 3 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.76 $Y=0.865
+ $X2=0.76 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_1%C 3 7 9 12 13
c32 13 0 7.87058e-20 $X=1.21 $Y=1.51
c33 7 0 1.92174e-19 $X=1.3 $Y=2.465
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.21 $Y=1.51
+ $X2=1.21 $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.21 $Y=1.51
+ $X2=1.21 $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.51 $X2=1.21 $Y2=1.51
r37 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.21 $Y=1.665
+ $X2=1.21 $Y2=1.51
r38 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.3 $Y=2.465 $X2=1.3
+ $Y2=1.675
r39 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.3 $Y=0.655 $X2=1.3
+ $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_1%B 3 7 9 12 13
c35 3 0 7.87058e-20 $X=1.73 $Y=2.465
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.675
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.345
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.51 $X2=1.75 $Y2=1.51
r39 9 13 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.73 $Y=1.665
+ $X2=1.73 $Y2=1.51
r40 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.755 $Y=0.655
+ $X2=1.755 $Y2=1.345
r41 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.73 $Y=2.465
+ $X2=1.73 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_1%A_84_131# 1 2 9 12 15 16 22 26 28 32 35
r56 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.35
+ $X2=2.29 $Y2=1.515
r57 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.35
+ $X2=2.29 $Y2=1.185
r58 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.35 $X2=2.29 $Y2=1.35
r59 28 31 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=1.17
+ $X2=2.25 $Y2=1.35
r60 23 26 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=0.24 $Y=2.065
+ $X2=0.545 $Y2=2.065
r61 21 22 7.99165 $w=4.88e-07 $l=1.05e-07 $layer=LI1_cond $X=0.545 $Y=1.01
+ $X2=0.65 $Y2=1.01
r62 18 21 7.44498 $w=4.88e-07 $l=3.05e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.545 $Y2=1.01
r63 16 28 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=1.17
+ $X2=2.25 $Y2=1.17
r64 16 22 96.2299 $w=1.68e-07 $l=1.475e-06 $layer=LI1_cond $X=2.125 $Y=1.17
+ $X2=0.65 $Y2=1.17
r65 15 23 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.92
+ $X2=0.24 $Y2=2.065
r66 14 18 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.24 $Y=1.255
+ $X2=0.24 $Y2=1.01
r67 14 15 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=0.24 $Y=1.255
+ $X2=0.24 $Y2=1.92
r68 12 36 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.2 $Y=2.465 $X2=2.2
+ $Y2=1.515
r69 9 35 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.2 $Y=0.655 $X2=2.2
+ $Y2=1.185
r70 2 26 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.42
+ $Y=1.835 $X2=0.545 $Y2=2.045
r71 1 21 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.42
+ $Y=0.655 $X2=0.545 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_1%VPWR 1 2 9 15 18 19 21 22 23 33 34
r30 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r33 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 23 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 23 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 21 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.97 $Y2=3.33
r38 20 33 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=1.97 $Y2=3.33
r40 18 26 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.88 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 18 19 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.88 $Y=3.33 $X2=1.03
+ $Y2=3.33
r42 17 30 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.18 $Y=3.33 $X2=1.68
+ $Y2=3.33
r43 17 19 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.18 $Y=3.33 $X2=1.03
+ $Y2=3.33
r44 13 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=3.245
+ $X2=1.97 $Y2=3.33
r45 13 15 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=1.97 $Y=3.245
+ $X2=1.97 $Y2=2.365
r46 9 12 16.7104 $w=2.98e-07 $l=4.35e-07 $layer=LI1_cond $X=1.03 $Y=2.085
+ $X2=1.03 $Y2=2.52
r47 7 19 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=3.245 $X2=1.03
+ $Y2=3.33
r48 7 12 27.8507 $w=2.98e-07 $l=7.25e-07 $layer=LI1_cond $X=1.03 $Y=3.245
+ $X2=1.03 $Y2=2.52
r49 2 15 300 $w=1.7e-07 $l=6.06918e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.835 $X2=1.97 $Y2=2.365
r50 1 12 300 $w=1.7e-07 $l=8.00297e-07 $layer=licon1_PDIFF $count=2 $X=0.835
+ $Y=1.835 $X2=1.085 $Y2=2.52
r51 1 9 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.835
+ $Y=1.835 $X2=0.975 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_1%Y 1 2 3 10 12 14 18 19 20 21 22 23 24 37 53
r38 37 58 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=2.67 $Y=0.925
+ $X2=2.67 $Y2=0.915
r39 24 48 7.64504 $w=4.83e-07 $l=3.1e-07 $layer=LI1_cond $X=2.552 $Y=2.775
+ $X2=2.552 $Y2=2.465
r40 23 48 1.47968 $w=4.83e-07 $l=6e-08 $layer=LI1_cond $X=2.552 $Y=2.405
+ $X2=2.552 $Y2=2.465
r41 22 35 2.61584 $w=3.67e-07 $l=1.54771e-07 $layer=LI1_cond $X=2.552 $Y=2.005
+ $X2=2.67 $Y2=1.92
r42 22 43 2.61584 $w=3.67e-07 $l=8.5e-08 $layer=LI1_cond $X=2.552 $Y=2.005
+ $X2=2.552 $Y2=2.09
r43 22 23 7.39842 $w=4.83e-07 $l=3e-07 $layer=LI1_cond $X=2.552 $Y=2.105
+ $X2=2.552 $Y2=2.405
r44 22 43 0.369921 $w=4.83e-07 $l=1.5e-08 $layer=LI1_cond $X=2.552 $Y=2.105
+ $X2=2.552 $Y2=2.09
r45 21 35 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=1.92
r46 20 21 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.665
r47 19 58 4.83154 $w=5.88e-07 $l=3.8e-08 $layer=LI1_cond $X=2.5 $Y=0.877 $X2=2.5
+ $Y2=0.915
r48 19 20 15.3505 $w=2.48e-07 $l=3.33e-07 $layer=LI1_cond $X=2.67 $Y=0.962
+ $X2=2.67 $Y2=1.295
r49 19 37 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=2.67 $Y=0.962
+ $X2=2.67 $Y2=0.925
r50 18 19 6.52775 $w=5.88e-07 $l=3.22e-07 $layer=LI1_cond $X=2.5 $Y=0.555
+ $X2=2.5 $Y2=0.877
r51 18 53 3.54769 $w=5.88e-07 $l=1.75e-07 $layer=LI1_cond $X=2.5 $Y=0.555
+ $X2=2.5 $Y2=0.38
r52 15 17 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.635 $Y=2.005
+ $X2=1.492 $Y2=2.005
r53 14 22 4.2195 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=2.31 $Y=2.005
+ $X2=2.552 $Y2=2.005
r54 14 15 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.31 $Y=2.005
+ $X2=1.635 $Y2=2.005
r55 10 17 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.492 $Y=2.09
+ $X2=1.492 $Y2=2.005
r56 10 12 15.1637 $w=2.83e-07 $l=3.75e-07 $layer=LI1_cond $X=1.492 $Y=2.09
+ $X2=1.492 $Y2=2.465
r57 3 22 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=2.005
r58 3 48 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.835 $X2=2.415 $Y2=2.465
r59 2 17 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=1.375
+ $Y=1.835 $X2=1.515 $Y2=2.005
r60 2 12 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=1.375
+ $Y=1.835 $X2=1.515 $Y2=2.465
r61 1 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.275
+ $Y=0.235 $X2=2.415 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_1%VGND 1 6 11 12 13 23 24
r22 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r23 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r24 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r25 17 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r26 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r27 13 24 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r28 13 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r29 11 16 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.72
+ $Y2=0
r30 11 12 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.005
+ $Y2=0
r31 10 20 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.19 $Y=0 $X2=1.2
+ $Y2=0
r32 10 12 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=1.005
+ $Y2=0
r33 6 8 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.005 $Y=0.38
+ $X2=1.005 $Y2=0.83
r34 4 12 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.005 $Y=0.085
+ $X2=1.005 $Y2=0
r35 4 6 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.005 $Y=0.085
+ $X2=1.005 $Y2=0.38
r36 1 8 182 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_NDIFF $count=1 $X=0.835
+ $Y=0.655 $X2=0.985 $Y2=0.83
r37 1 6 182 $w=1.7e-07 $l=3.79967e-07 $layer=licon1_NDIFF $count=1 $X=0.835
+ $Y=0.655 $X2=1.085 $Y2=0.38
.ends

