* File: sky130_fd_sc_lp__clkbuf_16.pex.spice
* Created: Wed Sep  2 09:38:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUF_16%A 3 7 11 15 19 23 27 31 33 34 35 49
r74 47 49 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.695 $Y=1.29
+ $X2=1.795 $Y2=1.29
r75 45 47 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.365 $Y=1.29
+ $X2=1.695 $Y2=1.29
r76 44 45 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.935 $Y=1.29
+ $X2=1.365 $Y2=1.29
r77 42 44 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=0.675 $Y=1.29
+ $X2=0.935 $Y2=1.29
r78 39 42 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.505 $Y=1.29
+ $X2=0.675 $Y2=1.29
r79 35 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.695
+ $Y=1.29 $X2=1.695 $Y2=1.29
r80 34 35 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.29 $X2=1.68
+ $Y2=1.29
r81 33 34 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.675 $Y=1.29
+ $X2=1.2 $Y2=1.29
r82 33 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.675
+ $Y=1.29 $X2=0.675 $Y2=1.29
r83 29 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.455
+ $X2=1.795 $Y2=1.29
r84 29 31 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.795 $Y=1.455
+ $X2=1.795 $Y2=2.465
r85 25 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.125
+ $X2=1.795 $Y2=1.29
r86 25 27 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.795 $Y=1.125
+ $X2=1.795 $Y2=0.445
r87 21 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.455
+ $X2=1.365 $Y2=1.29
r88 21 23 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.365 $Y=1.455
+ $X2=1.365 $Y2=2.465
r89 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.125
+ $X2=1.365 $Y2=1.29
r90 17 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.365 $Y=1.125
+ $X2=1.365 $Y2=0.445
r91 13 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.455
+ $X2=0.935 $Y2=1.29
r92 13 15 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.935 $Y=1.455
+ $X2=0.935 $Y2=2.465
r93 9 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.125
+ $X2=0.935 $Y2=1.29
r94 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.935 $Y=1.125
+ $X2=0.935 $Y2=0.445
r95 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.455
+ $X2=0.505 $Y2=1.29
r96 5 7 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.505 $Y=1.455
+ $X2=0.505 $Y2=2.465
r97 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.125
+ $X2=0.505 $Y2=1.29
r98 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.505 $Y=1.125
+ $X2=0.505 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_16%A_116_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131 133
+ 135 139 143 147 151 152 153 154 157 161 165 167 172 175 176 177 180 184 187
+ 190 193 196 199 201 202
r392 202 238 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.425
+ $Y=1.37 $X2=8.425 $Y2=1.37
r393 201 202 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.425 $Y=1.295
+ $X2=8.425 $Y2=1.295
r394 199 233 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.565
+ $Y=1.37 $X2=7.565 $Y2=1.37
r395 198 201 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.565 $Y=1.295
+ $X2=8.425 $Y2=1.295
r396 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.565 $Y=1.295
+ $X2=7.565 $Y2=1.295
r397 196 228 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=1.37 $X2=6.7 $Y2=1.37
r398 195 198 0.554988 $w=2.3e-07 $l=8.65e-07 $layer=MET1_cond $X=6.7 $Y=1.295
+ $X2=7.565 $Y2=1.295
r399 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.7 $Y=1.295
+ $X2=6.7 $Y2=1.295
r400 193 223 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.845
+ $Y=1.37 $X2=5.845 $Y2=1.37
r401 192 195 0.548572 $w=2.3e-07 $l=8.55e-07 $layer=MET1_cond $X=5.845 $Y=1.295
+ $X2=6.7 $Y2=1.295
r402 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.845 $Y=1.295
+ $X2=5.845 $Y2=1.295
r403 190 218 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=1.37 $X2=4.985 $Y2=1.37
r404 189 192 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.985 $Y=1.295
+ $X2=5.845 $Y2=1.295
r405 189 190 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.985 $Y=1.295
+ $X2=4.985 $Y2=1.295
r406 187 213 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.125
+ $Y=1.37 $X2=4.125 $Y2=1.37
r407 186 189 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.125 $Y=1.295
+ $X2=4.985 $Y2=1.295
r408 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.125 $Y=1.295
+ $X2=4.125 $Y2=1.295
r409 184 208 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.265
+ $Y=1.37 $X2=3.265 $Y2=1.37
r410 183 186 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=3.265 $Y=1.295
+ $X2=4.125 $Y2=1.295
r411 183 184 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.265 $Y=1.295
+ $X2=3.265 $Y2=1.295
r412 180 264 9.86936 $w=5.63e-07 $l=2.4e-07 $layer=LI1_cond $X=2.267 $Y=1.295
+ $X2=2.267 $Y2=1.535
r413 179 183 0.513283 $w=2.3e-07 $l=8e-07 $layer=MET1_cond $X=2.465 $Y=1.295
+ $X2=3.265 $Y2=1.295
r414 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.465 $Y=1.295
+ $X2=2.465 $Y2=1.295
r415 175 264 8.0403 $w=2.13e-07 $l=1.5e-07 $layer=LI1_cond $X=2.092 $Y=1.685
+ $X2=2.092 $Y2=1.535
r416 173 205 45.2297 $w=3.57e-07 $l=3.35e-07 $layer=POLY_cond $X=2.28 $Y=1.205
+ $X2=2.615 $Y2=1.205
r417 172 173 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.28
+ $Y=1.03 $X2=2.28 $Y2=1.03
r418 170 180 0.88912 $w=5.63e-07 $l=4.2e-08 $layer=LI1_cond $X=2.267 $Y=1.253
+ $X2=2.267 $Y2=1.295
r419 170 172 4.72081 $w=5.63e-07 $l=2.23e-07 $layer=LI1_cond $X=2.267 $Y=1.253
+ $X2=2.267 $Y2=1.03
r420 169 172 1.79941 $w=5.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.267 $Y=0.945
+ $X2=2.267 $Y2=1.03
r421 168 177 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.71 $Y=1.77
+ $X2=1.585 $Y2=1.77
r422 167 175 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.985 $Y=1.77
+ $X2=2.092 $Y2=1.685
r423 167 168 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.985 $Y=1.77
+ $X2=1.71 $Y2=1.77
r424 166 176 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.705 $Y=0.86
+ $X2=1.582 $Y2=0.86
r425 165 169 9.76632 $w=1.7e-07 $l=3.21705e-07 $layer=LI1_cond $X=1.985 $Y=0.86
+ $X2=2.267 $Y2=0.945
r426 165 166 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.985 $Y=0.86
+ $X2=1.705 $Y2=0.86
r427 161 163 39.1831 $w=2.48e-07 $l=8.5e-07 $layer=LI1_cond $X=1.585 $Y=2.04
+ $X2=1.585 $Y2=2.89
r428 159 177 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=1.855
+ $X2=1.585 $Y2=1.77
r429 159 161 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=1.585 $Y=1.855
+ $X2=1.585 $Y2=2.04
r430 155 176 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.582 $Y=0.775
+ $X2=1.582 $Y2=0.86
r431 155 157 15.5227 $w=2.43e-07 $l=3.3e-07 $layer=LI1_cond $X=1.582 $Y=0.775
+ $X2=1.582 $Y2=0.445
r432 153 177 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.46 $Y=1.77
+ $X2=1.585 $Y2=1.77
r433 153 154 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.46 $Y=1.77
+ $X2=0.855 $Y2=1.77
r434 151 176 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.46 $Y=0.86
+ $X2=1.582 $Y2=0.86
r435 151 152 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.46 $Y=0.86
+ $X2=0.84 $Y2=0.86
r436 147 149 36.9652 $w=2.63e-07 $l=8.5e-07 $layer=LI1_cond $X=0.722 $Y=2.04
+ $X2=0.722 $Y2=2.89
r437 145 154 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.722 $Y=1.855
+ $X2=0.855 $Y2=1.77
r438 145 147 8.04536 $w=2.63e-07 $l=1.85e-07 $layer=LI1_cond $X=0.722 $Y=1.855
+ $X2=0.722 $Y2=2.04
r439 141 152 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.715 $Y=0.775
+ $X2=0.84 $Y2=0.86
r440 141 143 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=0.715 $Y=0.775
+ $X2=0.715 $Y2=0.445
r441 137 139 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=9.065 $Y=1.535
+ $X2=9.065 $Y2=2.465
r442 133 137 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=9.065 $Y=1.205
+ $X2=9.065 $Y2=1.535
r443 133 135 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.065 $Y=1.205
+ $X2=9.065 $Y2=0.445
r444 129 131 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=8.635 $Y=1.535
+ $X2=8.635 $Y2=2.465
r445 125 133 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=8.635 $Y=1.205
+ $X2=9.065 $Y2=1.205
r446 125 129 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=8.635 $Y=1.205
+ $X2=8.635 $Y2=1.535
r447 125 238 28.3529 $w=3.57e-07 $l=2.1e-07 $layer=POLY_cond $X=8.635 $Y=1.205
+ $X2=8.425 $Y2=1.205
r448 125 127 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.635 $Y=1.205
+ $X2=8.635 $Y2=0.445
r449 121 123 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=8.205 $Y=1.535
+ $X2=8.205 $Y2=2.465
r450 117 238 29.7031 $w=3.57e-07 $l=2.2e-07 $layer=POLY_cond $X=8.205 $Y=1.205
+ $X2=8.425 $Y2=1.205
r451 117 121 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=8.205 $Y=1.205
+ $X2=8.205 $Y2=1.535
r452 117 119 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.205 $Y=1.205
+ $X2=8.205 $Y2=0.445
r453 113 115 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=7.775 $Y=1.535
+ $X2=7.775 $Y2=2.465
r454 109 117 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=7.775 $Y=1.205
+ $X2=8.205 $Y2=1.205
r455 109 113 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=7.775 $Y=1.205
+ $X2=7.775 $Y2=1.535
r456 109 233 28.3529 $w=3.57e-07 $l=2.1e-07 $layer=POLY_cond $X=7.775 $Y=1.205
+ $X2=7.565 $Y2=1.205
r457 109 111 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.775 $Y=1.205
+ $X2=7.775 $Y2=0.445
r458 105 107 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=7.345 $Y=1.535
+ $X2=7.345 $Y2=2.465
r459 101 233 29.7031 $w=3.57e-07 $l=2.2e-07 $layer=POLY_cond $X=7.345 $Y=1.205
+ $X2=7.565 $Y2=1.205
r460 101 105 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=7.345 $Y=1.205
+ $X2=7.345 $Y2=1.535
r461 101 103 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.345 $Y=1.205
+ $X2=7.345 $Y2=0.445
r462 97 99 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=6.915 $Y=1.535
+ $X2=6.915 $Y2=2.465
r463 93 101 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=6.915 $Y=1.205
+ $X2=7.345 $Y2=1.205
r464 93 97 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.915 $Y=1.205
+ $X2=6.915 $Y2=1.535
r465 93 228 29.028 $w=3.57e-07 $l=2.15e-07 $layer=POLY_cond $X=6.915 $Y=1.205
+ $X2=6.7 $Y2=1.205
r466 93 95 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.915 $Y=1.205
+ $X2=6.915 $Y2=0.445
r467 89 91 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=6.485 $Y=1.535
+ $X2=6.485 $Y2=2.465
r468 85 228 29.028 $w=3.57e-07 $l=2.15e-07 $layer=POLY_cond $X=6.485 $Y=1.205
+ $X2=6.7 $Y2=1.205
r469 85 89 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.485 $Y=1.205
+ $X2=6.485 $Y2=1.535
r470 85 87 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.485 $Y=1.205
+ $X2=6.485 $Y2=0.445
r471 81 83 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=6.055 $Y=1.535
+ $X2=6.055 $Y2=2.465
r472 77 85 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=6.055 $Y=1.205
+ $X2=6.485 $Y2=1.205
r473 77 81 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.055 $Y=1.205
+ $X2=6.055 $Y2=1.535
r474 77 223 28.3529 $w=3.57e-07 $l=2.1e-07 $layer=POLY_cond $X=6.055 $Y=1.205
+ $X2=5.845 $Y2=1.205
r475 77 79 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.055 $Y=1.205
+ $X2=6.055 $Y2=0.445
r476 73 75 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=5.625 $Y=1.535
+ $X2=5.625 $Y2=2.465
r477 69 223 29.7031 $w=3.57e-07 $l=2.2e-07 $layer=POLY_cond $X=5.625 $Y=1.205
+ $X2=5.845 $Y2=1.205
r478 69 73 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.625 $Y=1.205
+ $X2=5.625 $Y2=1.535
r479 69 71 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.625 $Y=1.205
+ $X2=5.625 $Y2=0.445
r480 65 67 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=5.195 $Y=1.535
+ $X2=5.195 $Y2=2.465
r481 61 69 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=5.195 $Y=1.205
+ $X2=5.625 $Y2=1.205
r482 61 65 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.195 $Y=1.205
+ $X2=5.195 $Y2=1.535
r483 61 218 28.3529 $w=3.57e-07 $l=2.1e-07 $layer=POLY_cond $X=5.195 $Y=1.205
+ $X2=4.985 $Y2=1.205
r484 61 63 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.195 $Y=1.205
+ $X2=5.195 $Y2=0.445
r485 57 59 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=4.765 $Y=1.535
+ $X2=4.765 $Y2=2.465
r486 53 218 29.7031 $w=3.57e-07 $l=2.2e-07 $layer=POLY_cond $X=4.765 $Y=1.205
+ $X2=4.985 $Y2=1.205
r487 53 57 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.765 $Y=1.205
+ $X2=4.765 $Y2=1.535
r488 53 55 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.765 $Y=1.205
+ $X2=4.765 $Y2=0.445
r489 49 51 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=4.335 $Y=1.535
+ $X2=4.335 $Y2=2.465
r490 45 53 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=4.335 $Y=1.205
+ $X2=4.765 $Y2=1.205
r491 45 49 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.335 $Y=1.205
+ $X2=4.335 $Y2=1.535
r492 45 213 28.3529 $w=3.57e-07 $l=2.1e-07 $layer=POLY_cond $X=4.335 $Y=1.205
+ $X2=4.125 $Y2=1.205
r493 45 47 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.335 $Y=1.205
+ $X2=4.335 $Y2=0.445
r494 41 43 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=3.905 $Y=1.535
+ $X2=3.905 $Y2=2.465
r495 37 213 29.7031 $w=3.57e-07 $l=2.2e-07 $layer=POLY_cond $X=3.905 $Y=1.205
+ $X2=4.125 $Y2=1.205
r496 37 41 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.905 $Y=1.205
+ $X2=3.905 $Y2=1.535
r497 37 39 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.905 $Y=1.205
+ $X2=3.905 $Y2=0.445
r498 33 35 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=3.475 $Y=1.535
+ $X2=3.475 $Y2=2.465
r499 29 37 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=3.475 $Y=1.205
+ $X2=3.905 $Y2=1.205
r500 29 33 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.475 $Y=1.205
+ $X2=3.475 $Y2=1.535
r501 29 208 28.3529 $w=3.57e-07 $l=2.1e-07 $layer=POLY_cond $X=3.475 $Y=1.205
+ $X2=3.265 $Y2=1.205
r502 29 31 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.475 $Y=1.205
+ $X2=3.475 $Y2=0.445
r503 25 27 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=3.045 $Y=1.535
+ $X2=3.045 $Y2=2.465
r504 21 208 29.7031 $w=3.57e-07 $l=2.2e-07 $layer=POLY_cond $X=3.045 $Y=1.205
+ $X2=3.265 $Y2=1.205
r505 21 25 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.045 $Y=1.205
+ $X2=3.045 $Y2=1.535
r506 21 205 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=3.045 $Y=1.205
+ $X2=2.615 $Y2=1.205
r507 21 23 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.045 $Y=1.205
+ $X2=3.045 $Y2=0.445
r508 17 205 23.1043 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.615 $Y=1.535
+ $X2=2.615 $Y2=1.205
r509 17 19 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.615 $Y=1.535
+ $X2=2.615 $Y2=2.465
r510 13 205 23.1043 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.615 $Y=0.865
+ $X2=2.615 $Y2=1.205
r511 13 15 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.615 $Y=0.865
+ $X2=2.615 $Y2=0.445
r512 4 163 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.835 $X2=1.58 $Y2=2.89
r513 4 161 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.835 $X2=1.58 $Y2=2.04
r514 3 149 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.89
r515 3 147 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.04
r516 2 157 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.58 $Y2=0.445
r517 1 143 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.235 $X2=0.72 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 34 36 42 48
+ 52 56 62 68 74 80 84 88 94 98 100 105 106 107 108 109 111 116 121 126 138 143
+ 152 155 158 161 164 167 170 174 184
r193 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r194 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r195 167 168 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r196 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r197 162 184 0.0432039 $w=4.9e-07 $l=1.55e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.925 $Y2=3.33
r198 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r199 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r200 156 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r201 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r202 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r204 147 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r205 147 171 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r206 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r207 144 170 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.42 $Y2=3.33
r208 144 146 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.88 $Y2=3.33
r209 143 173 4.56306 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=9.362 $Y2=3.33
r210 143 146 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=8.88 $Y2=3.33
r211 142 171 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r212 142 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r213 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 139 167 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.56 $Y2=3.33
r215 139 141 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.92 $Y2=3.33
r216 138 170 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.265 $Y=3.33
+ $X2=8.42 $Y2=3.33
r217 138 141 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.265 $Y=3.33
+ $X2=7.92 $Y2=3.33
r218 137 168 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r219 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r220 134 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r221 134 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r222 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r223 131 164 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.135 $Y=3.33
+ $X2=4.98 $Y2=3.33
r224 131 133 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.135 $Y=3.33
+ $X2=5.52 $Y2=3.33
r225 130 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r226 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r227 127 161 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.12 $Y2=3.33
r228 127 129 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.56 $Y2=3.33
r229 126 164 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.825 $Y=3.33
+ $X2=4.98 $Y2=3.33
r230 126 129 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.825 $Y=3.33
+ $X2=4.56 $Y2=3.33
r231 125 184 0.0905888 $w=4.9e-07 $l=3.25e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.925 $Y2=3.33
r232 125 159 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r233 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r234 122 158 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.26 $Y2=3.33
r235 122 124 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.6 $Y2=3.33
r236 121 161 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=4.12 $Y2=3.33
r237 121 124 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.6 $Y2=3.33
r238 120 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r239 120 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r240 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r241 117 152 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.157 $Y2=3.33
r242 117 119 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.68 $Y2=3.33
r243 116 155 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.88 $Y=3.33
+ $X2=2.215 $Y2=3.33
r244 116 119 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=3.33
+ $X2=1.68 $Y2=3.33
r245 115 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r246 115 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r247 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r248 112 149 4.39854 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=3.33
+ $X2=0.21 $Y2=3.33
r249 112 114 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.42 $Y=3.33
+ $X2=0.72 $Y2=3.33
r250 111 152 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.157 $Y2=3.33
r251 111 114 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.72 $Y2=3.33
r252 109 165 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r253 109 130 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r254 107 136 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.48 $Y2=3.33
r255 107 108 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.697 $Y2=3.33
r256 105 133 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=3.33
+ $X2=5.52 $Y2=3.33
r257 105 106 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.685 $Y=3.33
+ $X2=5.84 $Y2=3.33
r258 104 136 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.995 $Y=3.33
+ $X2=6.48 $Y2=3.33
r259 104 106 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.995 $Y=3.33
+ $X2=5.84 $Y2=3.33
r260 100 103 30.6118 $w=3.18e-07 $l=8.5e-07 $layer=LI1_cond $X=9.285 $Y=2.04
+ $X2=9.285 $Y2=2.89
r261 98 173 3.11905 $w=3.2e-07 $l=1.17346e-07 $layer=LI1_cond $X=9.285 $Y=3.245
+ $X2=9.362 $Y2=3.33
r262 98 103 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=9.285 $Y=3.245
+ $X2=9.285 $Y2=2.89
r263 94 97 31.5992 $w=3.08e-07 $l=8.5e-07 $layer=LI1_cond $X=8.42 $Y=2.04
+ $X2=8.42 $Y2=2.89
r264 92 170 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=3.33
r265 92 97 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=2.89
r266 88 91 31.5992 $w=3.08e-07 $l=8.5e-07 $layer=LI1_cond $X=7.56 $Y=2.04
+ $X2=7.56 $Y2=2.89
r267 86 167 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=3.245
+ $X2=7.56 $Y2=3.33
r268 86 91 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=7.56 $Y=3.245
+ $X2=7.56 $Y2=2.89
r269 85 108 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.85 $Y=3.33
+ $X2=6.697 $Y2=3.33
r270 84 167 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.405 $Y=3.33
+ $X2=7.56 $Y2=3.33
r271 84 85 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.405 $Y=3.33
+ $X2=6.85 $Y2=3.33
r272 80 83 32.1173 $w=3.03e-07 $l=8.5e-07 $layer=LI1_cond $X=6.697 $Y=2.04
+ $X2=6.697 $Y2=2.89
r273 78 108 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.697 $Y=3.245
+ $X2=6.697 $Y2=3.33
r274 78 83 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=6.697 $Y=3.245
+ $X2=6.697 $Y2=2.89
r275 74 77 31.5992 $w=3.08e-07 $l=8.5e-07 $layer=LI1_cond $X=5.84 $Y=2.04
+ $X2=5.84 $Y2=2.89
r276 72 106 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.84 $Y=3.245
+ $X2=5.84 $Y2=3.33
r277 72 77 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=5.84 $Y=3.245
+ $X2=5.84 $Y2=2.89
r278 68 71 31.5992 $w=3.08e-07 $l=8.5e-07 $layer=LI1_cond $X=4.98 $Y=2.04
+ $X2=4.98 $Y2=2.89
r279 66 164 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=3.245
+ $X2=4.98 $Y2=3.33
r280 66 71 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=4.98 $Y=3.245
+ $X2=4.98 $Y2=2.89
r281 62 65 31.5992 $w=3.08e-07 $l=8.5e-07 $layer=LI1_cond $X=4.12 $Y=2.04
+ $X2=4.12 $Y2=2.89
r282 60 161 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=3.245
+ $X2=4.12 $Y2=3.33
r283 60 65 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=4.12 $Y=3.245
+ $X2=4.12 $Y2=2.89
r284 56 59 31.5992 $w=3.08e-07 $l=8.5e-07 $layer=LI1_cond $X=3.26 $Y=2.04
+ $X2=3.26 $Y2=2.89
r285 54 158 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r286 54 59 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.89
r287 53 155 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.215 $Y2=3.33
r288 52 158 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=3.26 $Y2=3.33
r289 52 53 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=2.55 $Y2=3.33
r290 48 51 13.2104 $w=6.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.215 $Y=2.19
+ $X2=2.215 $Y2=2.93
r291 46 155 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=3.245
+ $X2=2.215 $Y2=3.33
r292 46 51 5.62335 $w=6.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.215 $Y=3.245
+ $X2=2.215 $Y2=2.93
r293 42 45 32.1814 $w=2.63e-07 $l=7.4e-07 $layer=LI1_cond $X=1.157 $Y=2.19
+ $X2=1.157 $Y2=2.93
r294 40 152 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.157 $Y=3.245
+ $X2=1.157 $Y2=3.33
r295 40 45 13.6989 $w=2.63e-07 $l=3.15e-07 $layer=LI1_cond $X=1.157 $Y=3.245
+ $X2=1.157 $Y2=2.93
r296 36 39 33.206 $w=2.93e-07 $l=8.5e-07 $layer=LI1_cond $X=0.272 $Y=2.04
+ $X2=0.272 $Y2=2.89
r297 34 149 3.07898 $w=2.95e-07 $l=1.11781e-07 $layer=LI1_cond $X=0.272 $Y=3.245
+ $X2=0.21 $Y2=3.33
r298 34 39 13.8684 $w=2.93e-07 $l=3.55e-07 $layer=LI1_cond $X=0.272 $Y=3.245
+ $X2=0.272 $Y2=2.89
r299 11 103 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=1.835 $X2=9.28 $Y2=2.89
r300 11 100 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=1.835 $X2=9.28 $Y2=2.04
r301 10 97 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=8.28
+ $Y=1.835 $X2=8.42 $Y2=2.89
r302 10 94 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=8.28
+ $Y=1.835 $X2=8.42 $Y2=2.04
r303 9 91 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=7.42
+ $Y=1.835 $X2=7.56 $Y2=2.89
r304 9 88 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.42
+ $Y=1.835 $X2=7.56 $Y2=2.04
r305 8 83 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=6.56
+ $Y=1.835 $X2=6.7 $Y2=2.89
r306 8 80 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=6.56
+ $Y=1.835 $X2=6.7 $Y2=2.04
r307 7 77 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.835 $X2=5.84 $Y2=2.89
r308 7 74 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.835 $X2=5.84 $Y2=2.04
r309 6 71 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.835 $X2=4.98 $Y2=2.89
r310 6 68 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.835 $X2=4.98 $Y2=2.04
r311 5 65 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.835 $X2=4.12 $Y2=2.89
r312 5 62 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.835 $X2=4.12 $Y2=2.04
r313 4 59 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=1.835 $X2=3.26 $Y2=2.89
r314 4 56 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=1.835 $X2=3.26 $Y2=2.04
r315 3 51 200 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=3 $X=1.87
+ $Y=1.835 $X2=2.01 $Y2=2.93
r316 3 48 200 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=3 $X=1.87
+ $Y=1.835 $X2=2.01 $Y2=2.19
r317 2 45 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=2.93
r318 2 42 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=2.19
r319 1 39 400 $w=1.7e-07 $l=1.12985e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.29 $Y2=2.89
r320 1 36 400 $w=1.7e-07 $l=2.71662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.29 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 49 52 62 72 82 92 102 112 122 126
r179 125 129 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=8.85 $Y=2.035
+ $X2=8.85 $Y2=2.89
r180 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.85 $Y=2.035
+ $X2=8.85 $Y2=2.035
r181 122 125 84.2381 $w=2.08e-07 $l=1.595e-06 $layer=LI1_cond $X=8.85 $Y=0.44
+ $X2=8.85 $Y2=2.035
r182 116 126 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.99 $Y=2.035
+ $X2=8.85 $Y2=2.035
r183 115 119 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=7.99 $Y=2.035
+ $X2=7.99 $Y2=2.89
r184 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.99 $Y=2.035
+ $X2=7.99 $Y2=2.035
r185 112 115 84.2381 $w=2.08e-07 $l=1.595e-06 $layer=LI1_cond $X=7.99 $Y=0.44
+ $X2=7.99 $Y2=2.035
r186 106 116 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.13 $Y=2.035
+ $X2=7.99 $Y2=2.035
r187 105 109 45.8297 $w=2.13e-07 $l=8.55e-07 $layer=LI1_cond $X=7.127 $Y=2.035
+ $X2=7.127 $Y2=2.89
r188 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.035
+ $X2=7.13 $Y2=2.035
r189 102 105 85.4952 $w=2.13e-07 $l=1.595e-06 $layer=LI1_cond $X=7.127 $Y=0.44
+ $X2=7.127 $Y2=2.035
r190 96 106 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.27 $Y=2.035
+ $X2=7.13 $Y2=2.035
r191 95 99 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=6.27 $Y=2.035
+ $X2=6.27 $Y2=2.89
r192 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.27 $Y=2.035
+ $X2=6.27 $Y2=2.035
r193 92 95 84.2381 $w=2.08e-07 $l=1.595e-06 $layer=LI1_cond $X=6.27 $Y=0.44
+ $X2=6.27 $Y2=2.035
r194 85 89 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=5.41 $Y=2.035
+ $X2=5.41 $Y2=2.89
r195 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.41 $Y=2.035
+ $X2=5.41 $Y2=2.035
r196 82 85 84.2381 $w=2.08e-07 $l=1.595e-06 $layer=LI1_cond $X=5.41 $Y=0.44
+ $X2=5.41 $Y2=2.035
r197 76 86 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.55 $Y=2.035
+ $X2=5.41 $Y2=2.035
r198 75 79 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=4.55 $Y=2.035
+ $X2=4.55 $Y2=2.89
r199 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.55 $Y=2.035
+ $X2=4.55 $Y2=2.035
r200 72 75 84.2381 $w=2.08e-07 $l=1.595e-06 $layer=LI1_cond $X=4.55 $Y=0.44
+ $X2=4.55 $Y2=2.035
r201 66 76 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=3.69 $Y=2.035
+ $X2=4.55 $Y2=2.035
r202 65 69 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=3.69 $Y=2.035
+ $X2=3.69 $Y2=2.89
r203 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.69 $Y=2.035
+ $X2=3.69 $Y2=2.035
r204 62 65 84.2381 $w=2.08e-07 $l=1.595e-06 $layer=LI1_cond $X=3.69 $Y=0.44
+ $X2=3.69 $Y2=2.035
r205 56 66 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=2.83 $Y=2.035
+ $X2=3.69 $Y2=2.035
r206 55 59 45.8297 $w=2.13e-07 $l=8.55e-07 $layer=LI1_cond $X=2.827 $Y=2.035
+ $X2=2.827 $Y2=2.89
r207 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.83 $Y=2.035
+ $X2=2.83 $Y2=2.035
r208 52 55 85.4952 $w=2.13e-07 $l=1.595e-06 $layer=LI1_cond $X=2.827 $Y=0.44
+ $X2=2.827 $Y2=2.035
r209 49 96 0.263058 $w=2.3e-07 $l=4.1e-07 $layer=MET1_cond $X=5.86 $Y=2.035
+ $X2=6.27 $Y2=2.035
r210 49 86 0.288722 $w=2.3e-07 $l=4.5e-07 $layer=MET1_cond $X=5.86 $Y=2.035
+ $X2=5.41 $Y2=2.035
r211 16 129 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=8.71
+ $Y=1.835 $X2=8.85 $Y2=2.89
r212 16 125 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=8.71
+ $Y=1.835 $X2=8.85 $Y2=2.04
r213 15 119 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=7.85
+ $Y=1.835 $X2=7.99 $Y2=2.89
r214 15 115 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.85
+ $Y=1.835 $X2=7.99 $Y2=2.04
r215 14 109 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=6.99
+ $Y=1.835 $X2=7.13 $Y2=2.89
r216 14 105 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=6.99
+ $Y=1.835 $X2=7.13 $Y2=2.04
r217 13 99 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=6.13
+ $Y=1.835 $X2=6.27 $Y2=2.89
r218 13 95 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=6.13
+ $Y=1.835 $X2=6.27 $Y2=2.04
r219 12 89 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.835 $X2=5.41 $Y2=2.89
r220 12 85 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.835 $X2=5.41 $Y2=2.04
r221 11 79 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.835 $X2=4.55 $Y2=2.89
r222 11 75 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.835 $X2=4.55 $Y2=2.04
r223 10 69 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.835 $X2=3.69 $Y2=2.89
r224 10 65 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.835 $X2=3.69 $Y2=2.04
r225 9 59 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=2.69
+ $Y=1.835 $X2=2.83 $Y2=2.89
r226 9 55 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.69
+ $Y=1.835 $X2=2.83 $Y2=2.04
r227 8 122 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=8.71
+ $Y=0.235 $X2=8.85 $Y2=0.44
r228 7 112 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=7.85
+ $Y=0.235 $X2=7.99 $Y2=0.44
r229 6 102 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=6.99
+ $Y=0.235 $X2=7.13 $Y2=0.44
r230 5 92 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=6.13
+ $Y=0.235 $X2=6.27 $Y2=0.44
r231 4 82 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.27
+ $Y=0.235 $X2=5.41 $Y2=0.44
r232 3 72 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.235 $X2=4.55 $Y2=0.44
r233 2 62 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.235 $X2=3.69 $Y2=0.44
r234 1 52 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.69
+ $Y=0.235 $X2=2.83 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 34 36 40 42
+ 46 50 54 58 62 64 68 72 74 76 79 80 81 82 83 85 95 100 112 117 126 131 134 136
+ 139 142 145 148 152 162
r165 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r166 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r167 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r168 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r169 140 162 0.0432039 $w=4.9e-07 $l=1.55e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=3.925 $Y2=0
r170 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r171 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r172 133 134 10.4808 $w=6.88e-07 $l=1.5e-07 $layer=LI1_cond $X=2.4 $Y=0.26
+ $X2=2.55 $Y2=0.26
r173 130 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.12 $Y2=0
r174 129 133 4.16027 $w=6.88e-07 $l=2.4e-07 $layer=LI1_cond $X=2.16 $Y=0.26
+ $X2=2.4 $Y2=0.26
r175 129 131 12.821 $w=6.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.16 $Y=0.26
+ $X2=1.875 $Y2=0.26
r176 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r177 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r178 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r179 121 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r180 121 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r181 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r182 118 148 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.575 $Y=0
+ $X2=8.42 $Y2=0
r183 118 120 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.575 $Y=0
+ $X2=8.88 $Y2=0
r184 117 151 4.56306 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=9.362 $Y2=0
r185 117 120 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=8.88 $Y2=0
r186 116 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r187 116 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r188 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r189 113 145 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.56 $Y2=0
r190 113 115 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.92 $Y2=0
r191 112 148 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.265 $Y=0
+ $X2=8.42 $Y2=0
r192 112 115 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.265 $Y=0
+ $X2=7.92 $Y2=0
r193 111 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r194 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r195 108 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.48 $Y2=0
r196 108 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r197 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r198 105 142 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.135 $Y=0
+ $X2=4.98 $Y2=0
r199 105 107 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.135 $Y=0
+ $X2=5.52 $Y2=0
r200 104 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r201 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r202 101 139 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=4.12 $Y2=0
r203 101 103 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=4.56 $Y2=0
r204 100 142 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.98 $Y2=0
r205 100 103 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.56 $Y2=0
r206 99 162 0.0905888 $w=4.9e-07 $l=3.25e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=3.925 $Y2=0
r207 99 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r208 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r209 96 136 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=3.26 $Y2=0
r210 96 98 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.6
+ $Y2=0
r211 95 139 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.965 $Y=0
+ $X2=4.12 $Y2=0
r212 95 98 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=3.6
+ $Y2=0
r213 94 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r214 94 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r215 93 131 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.68 $Y=0
+ $X2=1.875 $Y2=0
r216 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r217 91 126 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.15
+ $Y2=0
r218 91 93 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.68
+ $Y2=0
r219 89 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r220 89 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r221 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r222 86 123 4.39854 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.21
+ $Y2=0
r223 86 88 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.72
+ $Y2=0
r224 85 126 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.15
+ $Y2=0
r225 85 88 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.72
+ $Y2=0
r226 83 143 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=5.04 $Y2=0
r227 83 104 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=4.56 $Y2=0
r228 81 110 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.48 $Y2=0
r229 81 82 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.697 $Y2=0
r230 79 107 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=0
+ $X2=5.52 $Y2=0
r231 79 80 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.685 $Y=0 $X2=5.84
+ $Y2=0
r232 78 110 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.995 $Y=0
+ $X2=6.48 $Y2=0
r233 78 80 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.995 $Y=0 $X2=5.84
+ $Y2=0
r234 74 151 3.11905 $w=3.2e-07 $l=1.17346e-07 $layer=LI1_cond $X=9.285 $Y=0.085
+ $X2=9.362 $Y2=0
r235 74 76 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=9.285 $Y=0.085
+ $X2=9.285 $Y2=0.44
r236 70 148 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0
r237 70 72 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0.44
r238 66 145 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=0.085
+ $X2=7.56 $Y2=0
r239 66 68 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=7.56 $Y=0.085
+ $X2=7.56 $Y2=0.44
r240 65 82 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.85 $Y=0 $X2=6.697
+ $Y2=0
r241 64 145 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.405 $Y=0
+ $X2=7.56 $Y2=0
r242 64 65 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.405 $Y=0
+ $X2=6.85 $Y2=0
r243 60 82 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.697 $Y=0.085
+ $X2=6.697 $Y2=0
r244 60 62 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=6.697 $Y=0.085
+ $X2=6.697 $Y2=0.44
r245 56 80 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.84 $Y=0.085
+ $X2=5.84 $Y2=0
r246 56 58 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=5.84 $Y=0.085
+ $X2=5.84 $Y2=0.44
r247 52 142 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r248 52 54 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.44
r249 48 139 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=0.085
+ $X2=4.12 $Y2=0
r250 48 50 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=4.12 $Y=0.085
+ $X2=4.12 $Y2=0.44
r251 44 136 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=0.085
+ $X2=3.26 $Y2=0
r252 44 46 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=3.26 $Y=0.085
+ $X2=3.26 $Y2=0.44
r253 42 136 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.105 $Y=0
+ $X2=3.26 $Y2=0
r254 42 134 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.105 $Y=0
+ $X2=2.55 $Y2=0
r255 38 126 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r256 38 40 14.6113 $w=2.78e-07 $l=3.55e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.44
r257 34 123 3.07898 $w=2.95e-07 $l=1.11781e-07 $layer=LI1_cond $X=0.272 $Y=0.085
+ $X2=0.21 $Y2=0
r258 34 36 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=0.272 $Y=0.085
+ $X2=0.272 $Y2=0.445
r259 11 76 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.235 $X2=9.28 $Y2=0.44
r260 10 72 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=8.28
+ $Y=0.235 $X2=8.42 $Y2=0.44
r261 9 68 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=7.42
+ $Y=0.235 $X2=7.56 $Y2=0.44
r262 8 62 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=6.56
+ $Y=0.235 $X2=6.7 $Y2=0.44
r263 7 58 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.7
+ $Y=0.235 $X2=5.84 $Y2=0.44
r264 6 54 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.235 $X2=4.98 $Y2=0.44
r265 5 50 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.98
+ $Y=0.235 $X2=4.12 $Y2=0.44
r266 4 46 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.12
+ $Y=0.235 $X2=3.26 $Y2=0.44
r267 3 133 91 $w=1.7e-07 $l=6.24139e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.235 $X2=2.4 $Y2=0.44
r268 2 40 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.44
r269 1 36 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.29 $Y2=0.445
.ends

