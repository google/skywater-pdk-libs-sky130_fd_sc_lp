* File: sky130_fd_sc_lp__clkbuflp_8.pxi.spice
* Created: Wed Sep  2 09:39:13 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUFLP_8%A N_A_M1009_g N_A_M1007_g N_A_M1001_g
+ N_A_M1015_g N_A_M1017_g N_A_M1021_g N_A_M1011_g N_A_M1022_g A A N_A_c_101_n
+ N_A_c_102_n PM_SKY130_FD_SC_LP__CLKBUFLP_8%A
x_PM_SKY130_FD_SC_LP__CLKBUFLP_8%A_130_417# N_A_130_417#_M1001_s
+ N_A_130_417#_M1007_s N_A_130_417#_M1021_s N_A_130_417#_M1005_g
+ N_A_130_417#_M1003_g N_A_130_417#_M1000_g N_A_130_417#_M1004_g
+ N_A_130_417#_M1002_g N_A_130_417#_M1008_g N_A_130_417#_M1016_g
+ N_A_130_417#_M1010_g N_A_130_417#_M1013_g N_A_130_417#_M1006_g
+ N_A_130_417#_M1014_g N_A_130_417#_M1012_g N_A_130_417#_M1018_g
+ N_A_130_417#_M1019_g N_A_130_417#_M1020_g N_A_130_417#_M1023_g
+ N_A_130_417#_c_199_n N_A_130_417#_c_202_n N_A_130_417#_c_184_n
+ N_A_130_417#_c_209_n N_A_130_417#_c_185_n N_A_130_417#_c_186_n
+ N_A_130_417#_c_187_n N_A_130_417#_c_188_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_8%A_130_417#
x_PM_SKY130_FD_SC_LP__CLKBUFLP_8%VPWR N_VPWR_M1007_d N_VPWR_M1015_d
+ N_VPWR_M1022_d N_VPWR_M1004_d N_VPWR_M1013_d N_VPWR_M1018_d N_VPWR_M1023_d
+ N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n
+ N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n
+ N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n VPWR
+ N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_360_n N_VPWR_c_379_n
+ N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_8%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUFLP_8%X N_X_M1000_d N_X_M1006_d N_X_M1003_s
+ N_X_M1008_s N_X_M1014_s N_X_M1020_s N_X_c_482_n N_X_c_487_n N_X_c_471_n
+ N_X_c_478_n N_X_c_472_n N_X_c_506_n N_X_c_510_n N_X_c_514_n N_X_c_518_n X X X
+ X X N_X_c_475_n N_X_c_476_n PM_SKY130_FD_SC_LP__CLKBUFLP_8%X
x_PM_SKY130_FD_SC_LP__CLKBUFLP_8%VGND N_VGND_M1009_d N_VGND_M1011_d
+ N_VGND_M1016_s N_VGND_M1019_s N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n
+ N_VGND_c_590_n VGND N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n
+ N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_596_n N_VGND_c_597_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_8%VGND
cc_1 VNB N_A_M1009_g 0.0373938f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_2 VNB N_A_M1007_g 0.00645022f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.585
cc_3 VNB N_A_M1001_g 0.0268495f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.555
cc_4 VNB N_A_M1015_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.585
cc_5 VNB N_A_M1017_g 0.0257506f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.555
cc_6 VNB N_A_M1021_g 0.00472655f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.585
cc_7 VNB N_A_M1011_g 0.0391041f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.555
cc_8 VNB N_A_M1022_g 0.00527519f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.585
cc_9 VNB A 0.00441045f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A_c_101_n 0.0291071f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.4
cc_11 VNB N_A_c_102_n 0.106768f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.4
cc_12 VNB N_A_130_417#_M1005_g 0.0427486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_130_417#_M1003_g 0.00691238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_130_417#_M1000_g 0.0292254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_130_417#_M1004_g 0.00670015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_130_417#_M1002_g 0.0281162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_130_417#_M1008_g 0.00668281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_130_417#_M1016_g 0.0279039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_130_417#_M1010_g 0.0264533f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.4
cc_20 VNB N_A_130_417#_M1013_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.4
cc_21 VNB N_A_130_417#_M1006_g 0.0266657f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.4
cc_22 VNB N_A_130_417#_M1014_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_130_417#_M1012_g 0.0283706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_130_417#_M1018_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_130_417#_M1019_g 0.0361899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_130_417#_M1020_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_130_417#_M1023_g 0.00745847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_130_417#_c_184_n 0.00189921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_130_417#_c_185_n 0.0123493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_130_417#_c_186_n 0.0106271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_130_417#_c_187_n 0.00183274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_130_417#_c_188_n 0.21953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_360_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_471_n 0.00516499f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.565
cc_35 VNB N_X_c_472_n 0.00230484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB X 0.0780035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB X 0.0210982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_475_n 0.0135209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_476_n 0.00915451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_587_n 0.0107456f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.565
cc_41 VNB N_VGND_c_588_n 0.0298018f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.585
cc_42 VNB N_VGND_c_589_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.555
cc_43 VNB N_VGND_c_590_n 0.00859961f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.585
cc_44 VNB N_VGND_c_591_n 0.0604399f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.555
cc_45 VNB N_VGND_c_592_n 0.0348996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_593_n 0.0346777f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.4
cc_47 VNB N_VGND_c_594_n 0.0418016f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.565
cc_48 VNB N_VGND_c_595_n 0.378178f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.665
cc_49 VNB N_VGND_c_596_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_597_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_A_M1007_g 0.05162f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.585
cc_52 VPB N_A_M1015_g 0.03966f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.585
cc_53 VPB N_A_M1021_g 0.0391819f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.585
cc_54 VPB N_A_M1022_g 0.041206f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.585
cc_55 VPB A 0.0116793f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_56 VPB N_A_130_417#_M1003_g 0.0414132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_130_417#_M1004_g 0.0398013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_130_417#_M1008_g 0.0398013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_130_417#_M1013_g 0.0394337f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=1.4
cc_60 VPB N_A_130_417#_M1014_g 0.0394337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_130_417#_M1018_g 0.0397726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_130_417#_M1020_g 0.0397726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_130_417#_M1023_g 0.0534437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_130_417#_c_185_n 0.00912597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_361_n 0.0103398f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.585
cc_66 VPB N_VPWR_c_362_n 0.0463936f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_363_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_364_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_365_n 0.00308897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_366_n 0.00193185f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=1.4
cc_71 VPB N_VPWR_c_367_n 0.00195444f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.565
cc_72 VPB N_VPWR_c_368_n 0.00216196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_369_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_370_n 0.0460249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_371_n 0.0178027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_372_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_373_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_374_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_375_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_376_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_377_n 0.0153494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_360_n 0.0573115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_379_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_380_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_381_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_382_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_X_c_471_n 0.00497325f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=1.565
cc_88 VPB N_X_c_478_n 0.00230158f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.585
cc_89 VPB X 0.0088319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_X_c_475_n 0.00324829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_X_c_476_n 0.00607059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 N_A_M1022_g N_A_130_417#_M1003_g 0.0230805f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_93 N_A_M1007_g N_A_130_417#_c_199_n 0.0251227f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_94 N_A_M1015_g N_A_130_417#_c_199_n 0.0215039f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_95 N_A_M1021_g N_A_130_417#_c_199_n 6.78081e-19 $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_96 N_A_M1009_g N_A_130_417#_c_202_n 0.00220307f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_97 N_A_M1001_g N_A_130_417#_c_202_n 0.00906401f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_98 N_A_M1017_g N_A_130_417#_c_202_n 0.00961145f $X=1.265 $Y=0.555 $X2=0 $Y2=0
cc_99 N_A_M1011_g N_A_130_417#_c_202_n 0.00343067f $X=1.625 $Y=0.555 $X2=0 $Y2=0
cc_100 N_A_M1001_g N_A_130_417#_c_184_n 0.00465827f $X=0.835 $Y=0.555 $X2=0
+ $Y2=0
cc_101 N_A_M1017_g N_A_130_417#_c_184_n 0.0059863f $X=1.265 $Y=0.555 $X2=0 $Y2=0
cc_102 N_A_c_101_n N_A_130_417#_c_184_n 0.00429998f $X=0.565 $Y=1.4 $X2=0 $Y2=0
cc_103 N_A_M1015_g N_A_130_417#_c_209_n 7.07986e-19 $X=1.055 $Y=2.585 $X2=0
+ $Y2=0
cc_104 N_A_M1021_g N_A_130_417#_c_209_n 0.023344f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_105 N_A_M1022_g N_A_130_417#_c_209_n 0.019934f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_106 N_A_M1007_g N_A_130_417#_c_185_n 0.00813507f $X=0.525 $Y=2.585 $X2=0
+ $Y2=0
cc_107 N_A_M1001_g N_A_130_417#_c_185_n 2.85983e-19 $X=0.835 $Y=0.555 $X2=0
+ $Y2=0
cc_108 N_A_M1015_g N_A_130_417#_c_185_n 0.0268832f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_109 N_A_M1017_g N_A_130_417#_c_185_n 0.00665352f $X=1.265 $Y=0.555 $X2=0
+ $Y2=0
cc_110 N_A_M1021_g N_A_130_417#_c_185_n 0.0246786f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_111 N_A_M1011_g N_A_130_417#_c_185_n 0.00840909f $X=1.625 $Y=0.555 $X2=0
+ $Y2=0
cc_112 N_A_M1022_g N_A_130_417#_c_185_n 0.012166f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_113 A N_A_130_417#_c_185_n 0.0140032f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_c_101_n N_A_130_417#_c_185_n 0.0296324f $X=0.565 $Y=1.4 $X2=0 $Y2=0
cc_115 N_A_c_102_n N_A_130_417#_c_185_n 0.0551147f $X=2.115 $Y=1.4 $X2=0 $Y2=0
cc_116 N_A_c_102_n N_A_130_417#_c_186_n 0.0251311f $X=2.115 $Y=1.4 $X2=0 $Y2=0
cc_117 N_A_M1001_g N_A_130_417#_c_187_n 0.00543401f $X=0.835 $Y=0.555 $X2=0
+ $Y2=0
cc_118 N_A_M1017_g N_A_130_417#_c_187_n 0.00438181f $X=1.265 $Y=0.555 $X2=0
+ $Y2=0
cc_119 N_A_c_102_n N_A_130_417#_c_188_n 0.0230805f $X=2.115 $Y=1.4 $X2=0 $Y2=0
cc_120 N_A_M1007_g N_VPWR_c_362_n 0.0243287f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_121 N_A_M1015_g N_VPWR_c_362_n 0.00118975f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_122 A N_VPWR_c_362_n 0.0246433f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A_M1007_g N_VPWR_c_363_n 0.00839865f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_124 N_A_M1015_g N_VPWR_c_363_n 0.00839865f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_125 N_A_M1007_g N_VPWR_c_364_n 9.25377e-19 $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_126 N_A_M1015_g N_VPWR_c_364_n 0.0220137f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_127 N_A_M1021_g N_VPWR_c_364_n 0.0211007f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_128 N_A_M1022_g N_VPWR_c_364_n 9.25377e-19 $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_129 N_A_c_102_n N_VPWR_c_364_n 3.59803e-19 $X=2.115 $Y=1.4 $X2=0 $Y2=0
cc_130 N_A_M1021_g N_VPWR_c_365_n 9.25377e-19 $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_131 N_A_M1022_g N_VPWR_c_365_n 0.0234356f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_132 N_A_M1021_g N_VPWR_c_371_n 0.00801912f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_133 N_A_M1022_g N_VPWR_c_371_n 0.00870227f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_134 N_A_M1007_g N_VPWR_c_360_n 0.0136348f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_135 N_A_M1015_g N_VPWR_c_360_n 0.0136348f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_136 N_A_M1021_g N_VPWR_c_360_n 0.0127083f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_137 N_A_M1022_g N_VPWR_c_360_n 0.0143487f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_138 N_A_M1022_g N_X_c_482_n 8.56186e-19 $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_139 N_A_M1022_g N_X_c_478_n 7.6783e-19 $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_140 N_A_M1009_g N_VGND_c_588_n 0.0169797f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_VGND_c_588_n 0.002953f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_142 N_A_c_101_n N_VGND_c_588_n 0.0202745f $X=0.565 $Y=1.4 $X2=0 $Y2=0
cc_143 N_A_M1009_g N_VGND_c_591_n 0.00486043f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_144 N_A_M1001_g N_VGND_c_591_n 0.0054895f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_145 N_A_M1017_g N_VGND_c_591_n 0.00823051f $X=1.265 $Y=0.555 $X2=0 $Y2=0
cc_146 N_A_M1011_g N_VGND_c_591_n 0.0218118f $X=1.625 $Y=0.555 $X2=0 $Y2=0
cc_147 N_A_c_102_n N_VGND_c_591_n 0.00348157f $X=2.115 $Y=1.4 $X2=0 $Y2=0
cc_148 N_A_M1009_g N_VGND_c_595_n 0.00814425f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_149 N_A_M1001_g N_VGND_c_595_n 0.00980985f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_150 N_A_M1017_g N_VGND_c_595_n 0.00925395f $X=1.265 $Y=0.555 $X2=0 $Y2=0
cc_151 N_A_M1011_g N_VGND_c_595_n 0.0081443f $X=1.625 $Y=0.555 $X2=0 $Y2=0
cc_152 N_A_130_417#_c_199_n N_VPWR_c_362_n 0.0665496f $X=0.79 $Y=2.23 $X2=0
+ $Y2=0
cc_153 N_A_130_417#_c_199_n N_VPWR_c_363_n 0.0189236f $X=0.79 $Y=2.23 $X2=0
+ $Y2=0
cc_154 N_A_130_417#_c_199_n N_VPWR_c_364_n 0.0635845f $X=0.79 $Y=2.23 $X2=0
+ $Y2=0
cc_155 N_A_130_417#_c_209_n N_VPWR_c_364_n 0.0708348f $X=1.85 $Y=2.23 $X2=0
+ $Y2=0
cc_156 N_A_130_417#_c_185_n N_VPWR_c_364_n 0.0245797f $X=1.995 $Y=1.37 $X2=0
+ $Y2=0
cc_157 N_A_130_417#_M1003_g N_VPWR_c_365_n 0.022713f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_158 N_A_130_417#_M1004_g N_VPWR_c_365_n 9.25377e-19 $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_159 N_A_130_417#_c_209_n N_VPWR_c_365_n 0.0605246f $X=1.85 $Y=2.23 $X2=0
+ $Y2=0
cc_160 N_A_130_417#_c_186_n N_VPWR_c_365_n 0.00969843f $X=3.705 $Y=1.37 $X2=0
+ $Y2=0
cc_161 N_A_130_417#_M1003_g N_VPWR_c_366_n 9.25377e-19 $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_162 N_A_130_417#_M1004_g N_VPWR_c_366_n 0.0224631f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_163 N_A_130_417#_M1008_g N_VPWR_c_366_n 0.0224631f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_164 N_A_130_417#_M1013_g N_VPWR_c_366_n 9.25377e-19 $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_165 N_A_130_417#_M1008_g N_VPWR_c_367_n 9.25377e-19 $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_166 N_A_130_417#_M1013_g N_VPWR_c_367_n 0.0224718f $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_167 N_A_130_417#_M1014_g N_VPWR_c_367_n 0.0224718f $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_168 N_A_130_417#_M1018_g N_VPWR_c_367_n 9.25377e-19 $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_169 N_A_130_417#_c_188_n N_VPWR_c_367_n 3.969e-19 $X=6.355 $Y=1.375 $X2=0
+ $Y2=0
cc_170 N_A_130_417#_M1014_g N_VPWR_c_368_n 9.25377e-19 $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_171 N_A_130_417#_M1018_g N_VPWR_c_368_n 0.0225501f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_172 N_A_130_417#_M1020_g N_VPWR_c_368_n 0.0225501f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_173 N_A_130_417#_M1023_g N_VPWR_c_368_n 9.25377e-19 $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_174 N_A_130_417#_c_188_n N_VPWR_c_368_n 4.71465e-19 $X=6.355 $Y=1.375 $X2=0
+ $Y2=0
cc_175 N_A_130_417#_M1020_g N_VPWR_c_369_n 0.00839865f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_176 N_A_130_417#_M1023_g N_VPWR_c_369_n 0.00839865f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_177 N_A_130_417#_M1020_g N_VPWR_c_370_n 9.25377e-19 $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_178 N_A_130_417#_M1023_g N_VPWR_c_370_n 0.0236952f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_179 N_A_130_417#_c_209_n N_VPWR_c_371_n 0.0192645f $X=1.85 $Y=2.23 $X2=0
+ $Y2=0
cc_180 N_A_130_417#_M1003_g N_VPWR_c_373_n 0.00839865f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_181 N_A_130_417#_M1004_g N_VPWR_c_373_n 0.00839865f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_182 N_A_130_417#_M1008_g N_VPWR_c_375_n 0.00839865f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_183 N_A_130_417#_M1013_g N_VPWR_c_375_n 0.00839865f $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_184 N_A_130_417#_M1014_g N_VPWR_c_376_n 0.00839865f $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_185 N_A_130_417#_M1018_g N_VPWR_c_376_n 0.00839865f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_186 N_A_130_417#_M1007_s N_VPWR_c_360_n 0.00223559f $X=0.65 $Y=2.085 $X2=0
+ $Y2=0
cc_187 N_A_130_417#_M1021_s N_VPWR_c_360_n 0.00223559f $X=1.71 $Y=2.085 $X2=0
+ $Y2=0
cc_188 N_A_130_417#_M1003_g N_VPWR_c_360_n 0.0136348f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_189 N_A_130_417#_M1004_g N_VPWR_c_360_n 0.0136348f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_190 N_A_130_417#_M1008_g N_VPWR_c_360_n 0.0136348f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_191 N_A_130_417#_M1013_g N_VPWR_c_360_n 0.0136348f $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_192 N_A_130_417#_M1014_g N_VPWR_c_360_n 0.0136348f $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_193 N_A_130_417#_M1018_g N_VPWR_c_360_n 0.0136348f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_194 N_A_130_417#_M1020_g N_VPWR_c_360_n 0.0136348f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_195 N_A_130_417#_M1023_g N_VPWR_c_360_n 0.0136348f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_196 N_A_130_417#_c_199_n N_VPWR_c_360_n 0.0123859f $X=0.79 $Y=2.23 $X2=0
+ $Y2=0
cc_197 N_A_130_417#_c_209_n N_VPWR_c_360_n 0.0125574f $X=1.85 $Y=2.23 $X2=0
+ $Y2=0
cc_198 N_A_130_417#_M1003_g N_X_c_482_n 0.0231928f $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_199 N_A_130_417#_M1004_g N_X_c_482_n 0.0231928f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_200 N_A_130_417#_M1008_g N_X_c_482_n 8.56186e-19 $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_201 N_A_130_417#_M1005_g N_X_c_487_n 0.00116621f $X=2.595 $Y=0.51 $X2=0 $Y2=0
cc_202 N_A_130_417#_M1000_g N_X_c_487_n 0.00790997f $X=2.955 $Y=0.51 $X2=0 $Y2=0
cc_203 N_A_130_417#_M1002_g N_X_c_487_n 0.00817908f $X=3.385 $Y=0.51 $X2=0 $Y2=0
cc_204 N_A_130_417#_M1016_g N_X_c_487_n 0.0015572f $X=3.745 $Y=0.51 $X2=0 $Y2=0
cc_205 N_A_130_417#_M1004_g N_X_c_471_n 0.0182166f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_206 N_A_130_417#_M1002_g N_X_c_471_n 0.00995807f $X=3.385 $Y=0.51 $X2=0 $Y2=0
cc_207 N_A_130_417#_M1008_g N_X_c_471_n 0.0182166f $X=3.705 $Y=2.585 $X2=0 $Y2=0
cc_208 N_A_130_417#_M1016_g N_X_c_471_n 0.0144122f $X=3.745 $Y=0.51 $X2=0 $Y2=0
cc_209 N_A_130_417#_c_186_n N_X_c_471_n 0.0937684f $X=3.705 $Y=1.37 $X2=0 $Y2=0
cc_210 N_A_130_417#_c_188_n N_X_c_471_n 0.00632593f $X=6.355 $Y=1.375 $X2=0
+ $Y2=0
cc_211 N_A_130_417#_M1003_g N_X_c_478_n 0.00647735f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_212 N_A_130_417#_M1004_g N_X_c_478_n 0.00293606f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_213 N_A_130_417#_c_186_n N_X_c_478_n 0.027608f $X=3.705 $Y=1.37 $X2=0 $Y2=0
cc_214 N_A_130_417#_c_188_n N_X_c_478_n 0.00275645f $X=6.355 $Y=1.375 $X2=0
+ $Y2=0
cc_215 N_A_130_417#_M1005_g N_X_c_472_n 0.00106455f $X=2.595 $Y=0.51 $X2=0 $Y2=0
cc_216 N_A_130_417#_M1000_g N_X_c_472_n 0.00805932f $X=2.955 $Y=0.51 $X2=0 $Y2=0
cc_217 N_A_130_417#_M1002_g N_X_c_472_n 0.00406564f $X=3.385 $Y=0.51 $X2=0 $Y2=0
cc_218 N_A_130_417#_c_186_n N_X_c_472_n 0.0276413f $X=3.705 $Y=1.37 $X2=0 $Y2=0
cc_219 N_A_130_417#_c_188_n N_X_c_472_n 0.00272104f $X=6.355 $Y=1.375 $X2=0
+ $Y2=0
cc_220 N_A_130_417#_M1004_g N_X_c_506_n 8.56186e-19 $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_221 N_A_130_417#_M1008_g N_X_c_506_n 0.0231928f $X=3.705 $Y=2.585 $X2=0 $Y2=0
cc_222 N_A_130_417#_M1013_g N_X_c_506_n 0.0231928f $X=4.235 $Y=2.585 $X2=0 $Y2=0
cc_223 N_A_130_417#_M1014_g N_X_c_506_n 8.56186e-19 $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_224 N_A_130_417#_M1010_g N_X_c_510_n 0.00155479f $X=4.175 $Y=0.51 $X2=0 $Y2=0
cc_225 N_A_130_417#_M1006_g N_X_c_510_n 0.00821758f $X=4.535 $Y=0.51 $X2=0 $Y2=0
cc_226 N_A_130_417#_M1012_g N_X_c_510_n 0.0097387f $X=4.965 $Y=0.51 $X2=0 $Y2=0
cc_227 N_A_130_417#_M1019_g N_X_c_510_n 0.00151175f $X=5.325 $Y=0.51 $X2=0 $Y2=0
cc_228 N_A_130_417#_M1013_g N_X_c_514_n 8.9921e-19 $X=4.235 $Y=2.585 $X2=0 $Y2=0
cc_229 N_A_130_417#_M1014_g N_X_c_514_n 0.0235159f $X=4.765 $Y=2.585 $X2=0 $Y2=0
cc_230 N_A_130_417#_M1018_g N_X_c_514_n 0.0235159f $X=5.295 $Y=2.585 $X2=0 $Y2=0
cc_231 N_A_130_417#_M1020_g N_X_c_514_n 8.9921e-19 $X=5.825 $Y=2.585 $X2=0 $Y2=0
cc_232 N_A_130_417#_M1018_g N_X_c_518_n 0.00126492f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_233 N_A_130_417#_M1020_g N_X_c_518_n 0.0262623f $X=5.825 $Y=2.585 $X2=0 $Y2=0
cc_234 N_A_130_417#_M1023_g N_X_c_518_n 0.0341532f $X=6.355 $Y=2.585 $X2=0 $Y2=0
cc_235 N_A_130_417#_M1019_g X 0.0151991f $X=5.325 $Y=0.51 $X2=0 $Y2=0
cc_236 N_A_130_417#_M1020_g X 0.00723331f $X=5.825 $Y=2.585 $X2=0 $Y2=0
cc_237 N_A_130_417#_M1023_g X 0.0242936f $X=6.355 $Y=2.585 $X2=0 $Y2=0
cc_238 N_A_130_417#_c_188_n X 0.0435831f $X=6.355 $Y=1.375 $X2=0 $Y2=0
cc_239 N_A_130_417#_M1018_g N_X_c_475_n 0.0187657f $X=5.295 $Y=2.585 $X2=0 $Y2=0
cc_240 N_A_130_417#_M1019_g N_X_c_475_n 0.0086584f $X=5.325 $Y=0.51 $X2=0 $Y2=0
cc_241 N_A_130_417#_M1020_g N_X_c_475_n 0.0150541f $X=5.825 $Y=2.585 $X2=0 $Y2=0
cc_242 N_A_130_417#_c_188_n N_X_c_475_n 0.030556f $X=6.355 $Y=1.375 $X2=0 $Y2=0
cc_243 N_A_130_417#_M1008_g N_X_c_476_n 0.00566544f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_244 N_A_130_417#_M1016_g N_X_c_476_n 7.45367e-19 $X=3.745 $Y=0.51 $X2=0 $Y2=0
cc_245 N_A_130_417#_M1010_g N_X_c_476_n 0.0178431f $X=4.175 $Y=0.51 $X2=0 $Y2=0
cc_246 N_A_130_417#_M1013_g N_X_c_476_n 0.0258114f $X=4.235 $Y=2.585 $X2=0 $Y2=0
cc_247 N_A_130_417#_M1006_g N_X_c_476_n 0.0183041f $X=4.535 $Y=0.51 $X2=0 $Y2=0
cc_248 N_A_130_417#_M1014_g N_X_c_476_n 0.0264499f $X=4.765 $Y=2.585 $X2=0 $Y2=0
cc_249 N_A_130_417#_M1012_g N_X_c_476_n 0.018827f $X=4.965 $Y=0.51 $X2=0 $Y2=0
cc_250 N_A_130_417#_M1018_g N_X_c_476_n 0.00637636f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_251 N_A_130_417#_M1019_g N_X_c_476_n 0.00215701f $X=5.325 $Y=0.51 $X2=0 $Y2=0
cc_252 N_A_130_417#_M1020_g N_X_c_476_n 3.62586e-19 $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_253 N_A_130_417#_c_186_n N_X_c_476_n 0.027121f $X=3.705 $Y=1.37 $X2=0 $Y2=0
cc_254 N_A_130_417#_c_188_n N_X_c_476_n 0.0524917f $X=6.355 $Y=1.375 $X2=0 $Y2=0
cc_255 N_A_130_417#_c_202_n N_VGND_c_588_n 0.0211472f $X=1.05 $Y=0.385 $X2=0
+ $Y2=0
cc_256 N_A_130_417#_M1002_g N_VGND_c_589_n 0.00239092f $X=3.385 $Y=0.51 $X2=0
+ $Y2=0
cc_257 N_A_130_417#_M1016_g N_VGND_c_589_n 0.0113267f $X=3.745 $Y=0.51 $X2=0
+ $Y2=0
cc_258 N_A_130_417#_M1010_g N_VGND_c_589_n 0.0113256f $X=4.175 $Y=0.51 $X2=0
+ $Y2=0
cc_259 N_A_130_417#_M1006_g N_VGND_c_589_n 0.00239092f $X=4.535 $Y=0.51 $X2=0
+ $Y2=0
cc_260 N_A_130_417#_M1012_g N_VGND_c_590_n 0.00255802f $X=4.965 $Y=0.51 $X2=0
+ $Y2=0
cc_261 N_A_130_417#_M1019_g N_VGND_c_590_n 0.0150176f $X=5.325 $Y=0.51 $X2=0
+ $Y2=0
cc_262 N_A_130_417#_c_188_n N_VGND_c_590_n 0.00167892f $X=6.355 $Y=1.375 $X2=0
+ $Y2=0
cc_263 N_A_130_417#_M1005_g N_VGND_c_591_n 0.0238513f $X=2.595 $Y=0.51 $X2=0
+ $Y2=0
cc_264 N_A_130_417#_M1000_g N_VGND_c_591_n 0.00321414f $X=2.955 $Y=0.51 $X2=0
+ $Y2=0
cc_265 N_A_130_417#_c_202_n N_VGND_c_591_n 0.0425937f $X=1.05 $Y=0.385 $X2=0
+ $Y2=0
cc_266 N_A_130_417#_c_185_n N_VGND_c_591_n 0.0164775f $X=1.995 $Y=1.37 $X2=0
+ $Y2=0
cc_267 N_A_130_417#_c_186_n N_VGND_c_591_n 0.0306117f $X=3.705 $Y=1.37 $X2=0
+ $Y2=0
cc_268 N_A_130_417#_M1005_g N_VGND_c_592_n 0.00468308f $X=2.595 $Y=0.51 $X2=0
+ $Y2=0
cc_269 N_A_130_417#_M1000_g N_VGND_c_592_n 0.0055185f $X=2.955 $Y=0.51 $X2=0
+ $Y2=0
cc_270 N_A_130_417#_M1002_g N_VGND_c_592_n 0.0055185f $X=3.385 $Y=0.51 $X2=0
+ $Y2=0
cc_271 N_A_130_417#_M1016_g N_VGND_c_592_n 0.00486043f $X=3.745 $Y=0.51 $X2=0
+ $Y2=0
cc_272 N_A_130_417#_M1010_g N_VGND_c_593_n 0.00486043f $X=4.175 $Y=0.51 $X2=0
+ $Y2=0
cc_273 N_A_130_417#_M1006_g N_VGND_c_593_n 0.0055185f $X=4.535 $Y=0.51 $X2=0
+ $Y2=0
cc_274 N_A_130_417#_M1012_g N_VGND_c_593_n 0.00488972f $X=4.965 $Y=0.51 $X2=0
+ $Y2=0
cc_275 N_A_130_417#_M1019_g N_VGND_c_593_n 0.00486043f $X=5.325 $Y=0.51 $X2=0
+ $Y2=0
cc_276 N_A_130_417#_M1001_s N_VGND_c_595_n 0.00223559f $X=0.91 $Y=0.235 $X2=0
+ $Y2=0
cc_277 N_A_130_417#_M1005_g N_VGND_c_595_n 0.00783538f $X=2.595 $Y=0.51 $X2=0
+ $Y2=0
cc_278 N_A_130_417#_M1000_g N_VGND_c_595_n 0.00988872f $X=2.955 $Y=0.51 $X2=0
+ $Y2=0
cc_279 N_A_130_417#_M1002_g N_VGND_c_595_n 0.00600112f $X=3.385 $Y=0.51 $X2=0
+ $Y2=0
cc_280 N_A_130_417#_M1016_g N_VGND_c_595_n 0.00427207f $X=3.745 $Y=0.51 $X2=0
+ $Y2=0
cc_281 N_A_130_417#_M1010_g N_VGND_c_595_n 0.00426996f $X=4.175 $Y=0.51 $X2=0
+ $Y2=0
cc_282 N_A_130_417#_M1006_g N_VGND_c_595_n 0.00599903f $X=4.535 $Y=0.51 $X2=0
+ $Y2=0
cc_283 N_A_130_417#_M1012_g N_VGND_c_595_n 0.00823628f $X=4.965 $Y=0.51 $X2=0
+ $Y2=0
cc_284 N_A_130_417#_M1019_g N_VGND_c_595_n 0.00814425f $X=5.325 $Y=0.51 $X2=0
+ $Y2=0
cc_285 N_A_130_417#_c_202_n N_VGND_c_595_n 0.0129004f $X=1.05 $Y=0.385 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_360_n N_X_M1003_s 0.00223559f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_287 N_VPWR_c_360_n N_X_M1008_s 0.00223559f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_288 N_VPWR_c_360_n N_X_M1014_s 0.00223559f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_289 N_VPWR_c_360_n N_X_M1020_s 0.00223559f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_290 N_VPWR_c_365_n N_X_c_482_n 0.0652318f $X=2.38 $Y=2.23 $X2=0 $Y2=0
cc_291 N_VPWR_c_366_n N_X_c_482_n 0.0652318f $X=3.44 $Y=2.23 $X2=0 $Y2=0
cc_292 N_VPWR_c_373_n N_X_c_482_n 0.0189236f $X=3.275 $Y=3.33 $X2=0 $Y2=0
cc_293 N_VPWR_c_360_n N_X_c_482_n 0.0123859f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_294 N_VPWR_c_366_n N_X_c_471_n 0.0192682f $X=3.44 $Y=2.23 $X2=0 $Y2=0
cc_295 N_VPWR_c_366_n N_X_c_506_n 0.0652318f $X=3.44 $Y=2.23 $X2=0 $Y2=0
cc_296 N_VPWR_c_367_n N_X_c_506_n 0.0652318f $X=4.5 $Y=2.23 $X2=0 $Y2=0
cc_297 N_VPWR_c_375_n N_X_c_506_n 0.0189236f $X=4.335 $Y=3.33 $X2=0 $Y2=0
cc_298 N_VPWR_c_360_n N_X_c_506_n 0.0123859f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_299 N_VPWR_c_367_n N_X_c_514_n 0.0652318f $X=4.5 $Y=2.23 $X2=0 $Y2=0
cc_300 N_VPWR_c_368_n N_X_c_514_n 0.0652318f $X=5.56 $Y=2.23 $X2=0 $Y2=0
cc_301 N_VPWR_c_376_n N_X_c_514_n 0.0189236f $X=5.395 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_c_360_n N_X_c_514_n 0.0123859f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_c_368_n N_X_c_518_n 0.0652318f $X=5.56 $Y=2.23 $X2=0 $Y2=0
cc_304 N_VPWR_c_369_n N_X_c_518_n 0.0189236f $X=6.455 $Y=3.33 $X2=0 $Y2=0
cc_305 N_VPWR_c_370_n N_X_c_518_n 0.0652318f $X=6.62 $Y=2.23 $X2=0 $Y2=0
cc_306 N_VPWR_c_360_n N_X_c_518_n 0.0123859f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_307 N_VPWR_c_370_n X 0.015325f $X=6.62 $Y=2.23 $X2=0 $Y2=0
cc_308 N_VPWR_c_368_n N_X_c_475_n 0.0162522f $X=5.56 $Y=2.23 $X2=0 $Y2=0
cc_309 N_VPWR_c_367_n N_X_c_476_n 0.0210354f $X=4.5 $Y=2.23 $X2=0 $Y2=0
cc_310 N_X_c_471_n N_VGND_M1016_s 0.00175352f $X=3.805 $Y=1.795 $X2=0 $Y2=0
cc_311 N_X_c_487_n N_VGND_c_589_n 0.00869891f $X=3.17 $Y=0.51 $X2=0 $Y2=0
cc_312 N_X_c_471_n N_VGND_c_589_n 0.0153056f $X=3.805 $Y=1.795 $X2=0 $Y2=0
cc_313 N_X_c_510_n N_VGND_c_589_n 0.00878484f $X=4.75 $Y=0.51 $X2=0 $Y2=0
cc_314 N_X_c_476_n N_VGND_c_589_n 0.00192885f $X=5.195 $Y=1.48 $X2=0 $Y2=0
cc_315 N_X_c_510_n N_VGND_c_590_n 0.0121681f $X=4.75 $Y=0.51 $X2=0 $Y2=0
cc_316 X N_VGND_c_590_n 0.0361179f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_317 N_X_c_475_n N_VGND_c_590_n 0.0125612f $X=5.875 $Y=1.48 $X2=0 $Y2=0
cc_318 N_X_c_487_n N_VGND_c_591_n 0.0153571f $X=3.17 $Y=0.51 $X2=0 $Y2=0
cc_319 N_X_c_472_n N_VGND_c_591_n 0.0037806f $X=3.335 $Y=0.905 $X2=0 $Y2=0
cc_320 N_X_c_487_n N_VGND_c_592_n 0.0120325f $X=3.17 $Y=0.51 $X2=0 $Y2=0
cc_321 N_X_c_510_n N_VGND_c_593_n 0.0139364f $X=4.75 $Y=0.51 $X2=0 $Y2=0
cc_322 X N_VGND_c_594_n 0.0578502f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_323 N_X_M1000_d N_VGND_c_595_n 0.00233619f $X=3.03 $Y=0.235 $X2=0 $Y2=0
cc_324 N_X_M1006_d N_VGND_c_595_n 0.00233619f $X=4.61 $Y=0.235 $X2=0 $Y2=0
cc_325 N_X_c_487_n N_VGND_c_595_n 0.0119011f $X=3.17 $Y=0.51 $X2=0 $Y2=0
cc_326 N_X_c_471_n N_VGND_c_595_n 0.0167568f $X=3.805 $Y=1.795 $X2=0 $Y2=0
cc_327 N_X_c_510_n N_VGND_c_595_n 0.0133456f $X=4.75 $Y=0.51 $X2=0 $Y2=0
cc_328 X N_VGND_c_595_n 0.0331987f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_329 N_X_c_476_n N_VGND_c_595_n 0.0173834f $X=5.195 $Y=1.48 $X2=0 $Y2=0
cc_330 N_X_c_471_n A_1008_47# 0.00191768f $X=3.805 $Y=1.795 $X2=-0.19 $Y2=-0.245
cc_331 N_X_c_476_n A_692_47# 0.00215169f $X=5.195 $Y=1.48 $X2=-0.19 $Y2=-0.245
cc_332 N_VGND_c_595_n A_110_47# 0.00899413f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_333 N_VGND_c_595_n A_268_47# 0.00899413f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_334 N_VGND_c_595_n A_534_47# 0.00899413f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_335 N_VGND_c_595_n A_1008_47# 0.0028771f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_336 N_VGND_c_595_n A_692_47# 0.00287395f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_337 N_VGND_c_595_n A_850_47# 0.00899413f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
