* File: sky130_fd_sc_lp__and2b_2.spice
* Created: Fri Aug 28 10:05:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2b_2.pex.spice"
.subckt sky130_fd_sc_lp__and2b_2  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_N_M1004_g N_A_28_367#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.123333 AS=0.1197 PD=0.926667 PS=1.41 NRD=68.184 NRS=5.712 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1004_d N_A_186_239#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.246667 AS=0.1176 PD=1.85333 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A_186_239#_M1008_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.246667 AS=0.1176 PD=1.85333 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6 SA=75001
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 A_455_133# N_B_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.123333 PD=0.63 PS=0.926667 NRD=14.28 NRS=68.184 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_186_239#_M1005_d N_A_28_367#_M1005_g A_455_133# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_N_M1006_g N_A_28_367#_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1006_d N_A_186_239#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=4.9447 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75001 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A_186_239#_M1001_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.338625 AS=0.1764 PD=2.7075 PS=1.54 NRD=13.8097 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_A_186_239#_M1003_d N_B_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.112875 PD=0.7 PS=0.9025 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_28_367#_M1007_g N_A_186_239#_M1003_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__and2b_2.pxi.spice"
*
.ends
*
*
