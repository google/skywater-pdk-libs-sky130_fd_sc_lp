* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buflp_8 A VGND VNB VPB VPWR X
X0 VGND a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 X a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_644_47# a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_27_47# A a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_27_47# A a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 X a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_114_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_636_367# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_636_367# a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_644_47# a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_636_367# a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_114_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 X a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_114_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND A a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_636_367# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 X a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VGND a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_644_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_644_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_27_47# A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 X a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_636_367# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_644_47# a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_114_367# A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_27_47# A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_114_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 X a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 VPWR a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_636_367# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 VGND a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_644_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 a_636_367# a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 a_636_367# a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 a_644_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 VPWR A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 VPWR a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X40 VGND a_27_47# a_644_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X41 a_114_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X42 a_644_47# a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X43 VPWR a_27_47# a_636_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
