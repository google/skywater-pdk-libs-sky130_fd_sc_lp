* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR a_2227_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_1677_91# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_721_99# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_507_125# a_129_179# a_593_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1533_258# a_1360_451# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_679_125# a_721_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Q_N a_1360_451# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_1533_258# a_1360_451# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_1360_451# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR a_593_125# a_721_99# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_191_21# a_129_179# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_721_99# a_593_125# a_996_169# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 Q_N a_1360_451# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR SET_B a_1360_451# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 Q a_2227_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_1360_451# a_191_21# a_1468_451# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_1468_451# a_1533_258# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VGND a_1360_451# a_2227_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1280_159# a_1533_258# a_1677_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR a_593_125# a_1288_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 VGND CLK a_129_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR a_1360_451# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_1280_159# a_129_179# a_1360_451# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_191_21# a_129_179# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 VGND a_593_125# a_1173_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_996_169# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND a_2227_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_593_125# a_129_179# a_701_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_701_535# a_721_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VPWR a_1360_451# a_2227_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 Q a_2227_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_507_125# a_191_21# a_593_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 a_1288_451# a_129_179# a_1360_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X33 VPWR D a_507_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 VGND D a_507_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_593_125# a_191_21# a_679_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_1360_451# a_191_21# a_1173_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X37 VPWR CLK a_129_179# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
