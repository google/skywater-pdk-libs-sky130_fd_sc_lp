* File: sky130_fd_sc_lp__buf_2.pxi.spice
* Created: Wed Sep  2 09:34:55 2020
* 
x_PM_SKY130_FD_SC_LP__BUF_2%A_90_21# N_A_90_21#_M1004_d N_A_90_21#_M1002_d
+ N_A_90_21#_M1000_g N_A_90_21#_c_44_n N_A_90_21#_M1001_g N_A_90_21#_c_39_n
+ N_A_90_21#_M1003_g N_A_90_21#_M1005_g N_A_90_21#_c_40_n N_A_90_21#_c_53_p
+ N_A_90_21#_c_41_n N_A_90_21#_c_48_n N_A_90_21#_c_67_p N_A_90_21#_c_42_n
+ N_A_90_21#_c_50_n N_A_90_21#_c_51_n N_A_90_21#_c_43_n N_A_90_21#_c_52_n
+ PM_SKY130_FD_SC_LP__BUF_2%A_90_21#
x_PM_SKY130_FD_SC_LP__BUF_2%A N_A_M1004_g N_A_M1002_g A N_A_c_104_n N_A_c_105_n
+ PM_SKY130_FD_SC_LP__BUF_2%A
x_PM_SKY130_FD_SC_LP__BUF_2%VPWR N_VPWR_M1001_s N_VPWR_M1005_s N_VPWR_c_129_n
+ N_VPWR_c_130_n N_VPWR_c_131_n VPWR N_VPWR_c_132_n N_VPWR_c_133_n
+ N_VPWR_c_128_n N_VPWR_c_135_n PM_SKY130_FD_SC_LP__BUF_2%VPWR
x_PM_SKY130_FD_SC_LP__BUF_2%X N_X_M1000_d N_X_M1001_d X X X X X X X N_X_c_157_n
+ X N_X_c_168_n PM_SKY130_FD_SC_LP__BUF_2%X
x_PM_SKY130_FD_SC_LP__BUF_2%VGND N_VGND_M1000_s N_VGND_M1003_s N_VGND_c_177_n
+ N_VGND_c_178_n N_VGND_c_179_n VGND N_VGND_c_180_n N_VGND_c_181_n
+ N_VGND_c_182_n N_VGND_c_183_n PM_SKY130_FD_SC_LP__BUF_2%VGND
cc_1 VNB N_A_90_21#_M1000_g 0.0527848f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_2 VNB N_A_90_21#_c_39_n 0.00488061f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.65
cc_3 VNB N_A_90_21#_c_40_n 0.0060349f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.65
cc_4 VNB N_A_90_21#_c_41_n 0.0416961f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.51
cc_5 VNB N_A_90_21#_c_42_n 0.0446326f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=0.865
cc_6 VNB N_A_90_21#_c_43_n 0.0211803f $X=-0.19 $Y=-0.245 $X2=1.077 $Y2=1.185
cc_7 VNB N_A_M1002_g 0.00403147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A 0.00225867f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_9 VNB N_A_c_104_n 0.0465679f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.725
cc_10 VNB N_A_c_105_n 0.025717f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_11 VNB N_VPWR_c_128_n 0.103974f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.77
cc_12 VNB N_X_c_157_n 0.0109924f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.51
cc_13 VNB N_VGND_c_177_n 0.0125005f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.575
cc_14 VNB N_VGND_c_178_n 0.0496258f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_15 VNB N_VGND_c_179_n 0.0220435f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_16 VNB N_VGND_c_180_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.465
cc_17 VNB N_VGND_c_181_n 0.0207048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_182_n 0.160488f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.77
cc_19 VNB N_VGND_c_183_n 0.01379f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=1.855
cc_20 VPB N_A_90_21#_c_44_n 0.0216091f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.725
cc_21 VPB N_A_90_21#_c_39_n 0.00462802f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=1.65
cc_22 VPB N_A_90_21#_c_40_n 0.0074914f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.65
cc_23 VPB N_A_90_21#_c_41_n 0.0103983f $X=-0.19 $Y=1.655 $X2=1.11 $Y2=1.51
cc_24 VPB N_A_90_21#_c_48_n 0.00759299f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=1.77
cc_25 VPB N_A_90_21#_c_42_n 0.00145951f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=0.865
cc_26 VPB N_A_90_21#_c_50_n 0.0290946f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=1.98
cc_27 VPB N_A_90_21#_c_51_n 0.00764676f $X=-0.19 $Y=1.655 $X2=2.085 $Y2=1.77
cc_28 VPB N_A_90_21#_c_52_n 0.018598f $X=-0.19 $Y=1.655 $X2=1.077 $Y2=1.725
cc_29 VPB N_A_M1002_g 0.0280605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_129_n 0.013741f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.575
cc_31 VPB N_VPWR_c_130_n 0.00423396f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.655
cc_32 VPB N_VPWR_c_131_n 0.0310698f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.65
cc_33 VPB N_VPWR_c_132_n 0.0157625f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=2.465
cc_34 VPB N_VPWR_c_133_n 0.0217138f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=1.77
cc_35 VPB N_VPWR_c_128_n 0.0604633f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.77
cc_36 VPB N_VPWR_c_135_n 0.0129947f $X=-0.19 $Y=1.655 $X2=2.085 $Y2=1.98
cc_37 VPB N_X_c_157_n 6.42864e-19 $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.51
cc_38 N_A_90_21#_c_53_p N_A_M1002_g 5.09752e-19 $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_39 N_A_90_21#_c_41_n N_A_M1002_g 0.00306485f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_40 N_A_90_21#_c_48_n N_A_M1002_g 0.0204409f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_41 N_A_90_21#_c_50_n N_A_M1002_g 2.21843e-19 $X=2.05 $Y=1.98 $X2=0 $Y2=0
cc_42 N_A_90_21#_c_52_n N_A_M1002_g 0.0043113f $X=1.077 $Y=1.725 $X2=0 $Y2=0
cc_43 N_A_90_21#_c_53_p A 0.00939179f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_44 N_A_90_21#_c_41_n A 0.00178835f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_45 N_A_90_21#_c_48_n A 0.0201497f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_46 N_A_90_21#_c_42_n A 0.0252505f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_47 N_A_90_21#_c_53_p N_A_c_104_n 0.00118255f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_48 N_A_90_21#_c_41_n N_A_c_104_n 0.0226462f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_49 N_A_90_21#_c_48_n N_A_c_104_n 0.00626192f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_50 N_A_90_21#_c_42_n N_A_c_105_n 0.0211305f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_51 N_A_90_21#_c_48_n N_VPWR_M1005_s 0.00467055f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_52 N_A_90_21#_c_67_p N_VPWR_M1005_s 0.00161253f $X=1.275 $Y=1.77 $X2=0 $Y2=0
cc_53 N_A_90_21#_c_44_n N_VPWR_c_130_n 0.00312453f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_54 N_A_90_21#_c_44_n N_VPWR_c_131_n 5.32737e-19 $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_55 N_A_90_21#_c_41_n N_VPWR_c_131_n 0.0010375f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_56 N_A_90_21#_c_48_n N_VPWR_c_131_n 0.0365711f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_57 N_A_90_21#_c_67_p N_VPWR_c_131_n 0.0150129f $X=1.275 $Y=1.77 $X2=0 $Y2=0
cc_58 N_A_90_21#_c_50_n N_VPWR_c_131_n 0.0196467f $X=2.05 $Y=1.98 $X2=0 $Y2=0
cc_59 N_A_90_21#_c_52_n N_VPWR_c_131_n 0.0181237f $X=1.077 $Y=1.725 $X2=0 $Y2=0
cc_60 N_A_90_21#_c_44_n N_VPWR_c_132_n 0.00542163f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_61 N_A_90_21#_c_52_n N_VPWR_c_132_n 0.00486043f $X=1.077 $Y=1.725 $X2=0 $Y2=0
cc_62 N_A_90_21#_c_44_n N_VPWR_c_128_n 0.0106638f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_63 N_A_90_21#_c_50_n N_VPWR_c_128_n 0.0101286f $X=2.05 $Y=1.98 $X2=0 $Y2=0
cc_64 N_A_90_21#_c_52_n N_VPWR_c_128_n 0.00830891f $X=1.077 $Y=1.725 $X2=0 $Y2=0
cc_65 N_A_90_21#_c_44_n X 0.0033539f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_66 N_A_90_21#_M1000_g N_X_c_157_n 0.013595f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_67 N_A_90_21#_c_44_n N_X_c_157_n 0.0158034f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_68 N_A_90_21#_c_39_n N_X_c_157_n 0.00969971f $X=0.88 $Y=1.65 $X2=0 $Y2=0
cc_69 N_A_90_21#_c_40_n N_X_c_157_n 0.00638027f $X=0.545 $Y=1.65 $X2=0 $Y2=0
cc_70 N_A_90_21#_c_53_p N_X_c_157_n 0.0252569f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_71 N_A_90_21#_c_67_p N_X_c_157_n 0.0136388f $X=1.275 $Y=1.77 $X2=0 $Y2=0
cc_72 N_A_90_21#_c_43_n N_X_c_157_n 0.00955932f $X=1.077 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A_90_21#_c_52_n N_X_c_157_n 0.00501666f $X=1.077 $Y=1.725 $X2=0 $Y2=0
cc_74 N_A_90_21#_c_44_n N_X_c_168_n 0.00990779f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_75 N_A_90_21#_M1000_g N_VGND_c_178_n 0.00707803f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_76 N_A_90_21#_M1000_g N_VGND_c_179_n 6.94825e-19 $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_77 N_A_90_21#_c_53_p N_VGND_c_179_n 0.0120749f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_78 N_A_90_21#_c_41_n N_VGND_c_179_n 0.00667143f $X=1.11 $Y=1.51 $X2=0 $Y2=0
cc_79 N_A_90_21#_c_48_n N_VGND_c_179_n 0.00730801f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_80 N_A_90_21#_c_43_n N_VGND_c_179_n 0.0176583f $X=1.077 $Y=1.185 $X2=0 $Y2=0
cc_81 N_A_90_21#_M1000_g N_VGND_c_180_n 0.00585385f $X=0.525 $Y=0.655 $X2=0
+ $Y2=0
cc_82 N_A_90_21#_c_43_n N_VGND_c_180_n 0.00486043f $X=1.077 $Y=1.185 $X2=0 $Y2=0
cc_83 N_A_90_21#_c_42_n N_VGND_c_181_n 0.00428705f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_84 N_A_90_21#_M1000_g N_VGND_c_182_n 0.011499f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_85 N_A_90_21#_c_42_n N_VGND_c_182_n 0.00746184f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_86 N_A_90_21#_c_43_n N_VGND_c_182_n 0.00824727f $X=1.077 $Y=1.185 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VPWR_c_131_n 0.0176666f $X=1.835 $Y=2.155 $X2=0 $Y2=0
cc_88 N_A_M1002_g N_VPWR_c_133_n 0.00259749f $X=1.835 $Y=2.155 $X2=0 $Y2=0
cc_89 N_A_M1002_g N_VPWR_c_128_n 0.00344639f $X=1.835 $Y=2.155 $X2=0 $Y2=0
cc_90 A N_VGND_c_179_n 0.0195647f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_c_104_n N_VGND_c_179_n 0.00175237f $X=1.68 $Y=1.35 $X2=0 $Y2=0
cc_92 N_A_c_105_n N_VGND_c_179_n 0.0175507f $X=1.712 $Y=1.185 $X2=0 $Y2=0
cc_93 N_A_c_105_n N_VGND_c_181_n 0.00332367f $X=1.712 $Y=1.185 $X2=0 $Y2=0
cc_94 N_A_c_105_n N_VGND_c_182_n 0.00387424f $X=1.712 $Y=1.185 $X2=0 $Y2=0
cc_95 N_VPWR_c_128_n N_X_M1001_d 0.00380684f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_96 N_VPWR_c_131_n N_X_c_157_n 0.00132345f $X=1.62 $Y=2.11 $X2=0 $Y2=0
cc_97 N_VPWR_c_132_n N_X_c_168_n 0.0142168f $X=1.045 $Y=3.33 $X2=0 $Y2=0
cc_98 N_VPWR_c_128_n N_X_c_168_n 0.00991943f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_99 N_X_c_157_n N_VGND_c_178_n 0.0015231f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_100 N_X_c_157_n N_VGND_c_180_n 0.0136943f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_101 N_X_M1000_d N_VGND_c_182_n 0.0041489f $X=0.6 $Y=0.235 $X2=0 $Y2=0
cc_102 N_X_c_157_n N_VGND_c_182_n 0.00866972f $X=0.74 $Y=0.42 $X2=0 $Y2=0
