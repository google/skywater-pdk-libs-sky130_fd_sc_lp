* NGSPICE file created from sky130_fd_sc_lp__a21o_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_392_367# B1 a_86_269# VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=3.339e+11p ps=3.05e+06u
M1001 X a_86_269# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=7.392e+11p ps=6.8e+06u
M1002 X a_86_269# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.071e+12p ps=9.26e+06u
M1003 a_86_269# B1 VGND VNB nshort w=840000u l=150000u
+  ad=4.2e+11p pd=2.68e+06u as=0p ps=0u
M1004 a_392_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_464_47# A1 a_86_269# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1006 VPWR a_86_269# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_392_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_464_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_86_269# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

