* File: sky130_fd_sc_lp__and2b_1.pxi.spice
* Created: Wed Sep  2 09:30:54 2020
* 
x_PM_SKY130_FD_SC_LP__AND2B_1%A_N N_A_N_c_51_n N_A_N_M1003_g N_A_N_M1007_g A_N
+ N_A_N_c_54_n PM_SKY130_FD_SC_LP__AND2B_1%A_N
x_PM_SKY130_FD_SC_LP__AND2B_1%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1007_s
+ N_A_27_47#_c_83_n N_A_27_47#_M1000_g N_A_27_47#_c_84_n N_A_27_47#_M1006_g
+ N_A_27_47#_c_85_n N_A_27_47#_c_90_n N_A_27_47#_c_86_n N_A_27_47#_c_87_n
+ PM_SKY130_FD_SC_LP__AND2B_1%A_27_47#
x_PM_SKY130_FD_SC_LP__AND2B_1%B N_B_M1004_g N_B_M1001_g B B N_B_c_134_n
+ PM_SKY130_FD_SC_LP__AND2B_1%B
x_PM_SKY130_FD_SC_LP__AND2B_1%A_217_131# N_A_217_131#_M1006_s
+ N_A_217_131#_M1000_d N_A_217_131#_M1002_g N_A_217_131#_M1005_g
+ N_A_217_131#_c_164_n N_A_217_131#_c_165_n N_A_217_131#_c_166_n
+ N_A_217_131#_c_167_n N_A_217_131#_c_168_n N_A_217_131#_c_169_n
+ N_A_217_131#_c_170_n PM_SKY130_FD_SC_LP__AND2B_1%A_217_131#
x_PM_SKY130_FD_SC_LP__AND2B_1%VPWR N_VPWR_M1007_d N_VPWR_M1001_d N_VPWR_c_221_n
+ N_VPWR_c_222_n N_VPWR_c_230_n N_VPWR_c_223_n VPWR N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_220_n N_VPWR_c_227_n N_VPWR_c_228_n
+ PM_SKY130_FD_SC_LP__AND2B_1%VPWR
x_PM_SKY130_FD_SC_LP__AND2B_1%X N_X_M1005_d N_X_M1002_d X X X X X X X
+ N_X_c_257_n X PM_SKY130_FD_SC_LP__AND2B_1%X
x_PM_SKY130_FD_SC_LP__AND2B_1%VGND N_VGND_M1003_d N_VGND_M1004_d N_VGND_c_272_n
+ N_VGND_c_273_n VGND N_VGND_c_274_n N_VGND_c_275_n N_VGND_c_276_n
+ N_VGND_c_277_n N_VGND_c_278_n N_VGND_c_279_n PM_SKY130_FD_SC_LP__AND2B_1%VGND
cc_1 VNB N_A_N_c_51_n 0.0238409f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_2 VNB N_A_N_M1007_g 0.0338299f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.045
cc_3 VNB A_N 0.00314872f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_4 VNB N_A_N_c_54_n 0.0459056f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.93
cc_5 VNB N_A_27_47#_c_83_n 0.0525998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_84_n 0.0197499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_85_n 0.0519319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_86_n 0.00514658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_87_n 0.0186954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_M1004_g 0.039489f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.045
cc_11 VNB N_A_217_131#_M1002_g 0.0084707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_217_131#_c_164_n 0.00380438f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.93
cc_13 VNB N_A_217_131#_c_165_n 0.00103082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_217_131#_c_166_n 0.0028048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_217_131#_c_167_n 0.00537371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_217_131#_c_168_n 0.0361192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_217_131#_c_169_n 0.00595281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_217_131#_c_170_n 0.0218151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_220_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_257_n 0.0654952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_272_n 0.0176076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_273_n 0.0155638f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.93
cc_23 VNB N_VGND_c_274_n 0.017173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_275_n 0.029031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_276_n 0.0160663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_277_n 0.189946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_278_n 0.00574453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_279_n 0.0081157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_A_N_M1007_g 0.0306225f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.045
cc_30 VPB N_A_27_47#_c_83_n 0.00569125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_27_47#_M1000_g 0.022603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_27_47#_c_90_n 0.035376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_A_27_47#_c_86_n 0.00332786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_27_47#_c_87_n 5.12686e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_B_M1004_g 0.0209231f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.045
cc_36 VPB B 0.0238011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_B_c_134_n 0.0768375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_217_131#_M1002_g 0.0256759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_217_131#_c_166_n 0.00489221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_221_n 0.042222f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.93
cc_41 VPB N_VPWR_c_222_n 0.0025173f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.93
cc_42 VPB N_VPWR_c_223_n 0.00461104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_224_n 0.0282768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_225_n 0.0168508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_220_n 0.0871143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_227_n 0.0280771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_228_n 0.00401018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB X 0.0106633f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.93
cc_49 VPB X 0.0508904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_X_c_257_n 0.0022458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 N_A_N_M1007_g N_A_27_47#_c_83_n 0.0207021f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_52 N_A_N_M1007_g N_A_27_47#_M1000_g 0.0151338f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_53 N_A_N_M1007_g N_A_27_47#_c_84_n 0.00170124f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_54 A_N N_A_27_47#_c_84_n 4.11429e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_55 N_A_N_c_54_n N_A_27_47#_c_84_n 0.00366268f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_56 N_A_N_c_51_n N_A_27_47#_c_85_n 0.0138064f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_N_M1007_g N_A_27_47#_c_85_n 0.00867777f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_58 A_N N_A_27_47#_c_85_n 0.0257573f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_59 N_A_N_M1007_g N_A_27_47#_c_90_n 0.00796528f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_60 N_A_N_M1007_g N_A_27_47#_c_86_n 0.0252655f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_61 A_N N_A_27_47#_c_86_n 0.0190348f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_62 N_A_N_c_54_n N_A_27_47#_c_86_n 0.00385311f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_63 N_A_N_c_54_n N_A_27_47#_c_87_n 0.00628325f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_64 N_A_N_c_51_n N_A_217_131#_c_164_n 0.00117895f $X=0.475 $Y=0.765 $X2=0
+ $Y2=0
cc_65 A_N N_A_217_131#_c_164_n 0.0224298f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_66 N_A_N_c_54_n N_A_217_131#_c_164_n 0.00107239f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_67 N_A_N_M1007_g N_A_217_131#_c_165_n 4.04555e-19 $X=0.635 $Y=2.045 $X2=0
+ $Y2=0
cc_68 A_N N_A_217_131#_c_165_n 0.00225336f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_69 N_A_N_M1007_g N_A_217_131#_c_169_n 5.59188e-19 $X=0.635 $Y=2.045 $X2=0
+ $Y2=0
cc_70 N_A_N_M1007_g N_VPWR_c_221_n 0.00435231f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_71 N_A_N_M1007_g N_VPWR_c_230_n 0.00299096f $X=0.635 $Y=2.045 $X2=0 $Y2=0
cc_72 N_A_N_c_51_n N_VGND_c_272_n 0.00497299f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_73 A_N N_VGND_c_272_n 0.0216608f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_74 N_A_N_c_54_n N_VGND_c_272_n 0.00736858f $X=0.69 $Y=0.93 $X2=0 $Y2=0
cc_75 N_A_N_c_51_n N_VGND_c_274_n 0.00585385f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_N_c_51_n N_VGND_c_277_n 0.0129206f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_77 A_N N_VGND_c_277_n 0.00185122f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_83_n N_B_M1004_g 0.0217349f $X=1.23 $Y=1.665 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_84_n N_B_M1004_g 0.048796f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_83_n B 0.00104698f $X=1.23 $Y=1.665 $X2=0 $Y2=0
cc_81 N_A_27_47#_M1000_g B 0.0123391f $X=1.23 $Y=2.045 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_86_n B 0.00362327f $X=1.14 $Y=1.5 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_83_n N_A_217_131#_c_164_n 0.00842275f $X=1.23 $Y=1.665 $X2=0
+ $Y2=0
cc_84 N_A_27_47#_c_84_n N_A_217_131#_c_164_n 0.0104868f $X=1.425 $Y=1.185 $X2=0
+ $Y2=0
cc_85 N_A_27_47#_c_85_n N_A_217_131#_c_164_n 0.00229972f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_86 N_A_27_47#_c_86_n N_A_217_131#_c_164_n 0.00888308f $X=1.14 $Y=1.5 $X2=0
+ $Y2=0
cc_87 N_A_27_47#_c_84_n N_A_217_131#_c_165_n 0.00468445f $X=1.425 $Y=1.185 $X2=0
+ $Y2=0
cc_88 N_A_27_47#_c_83_n N_A_217_131#_c_166_n 0.00984805f $X=1.23 $Y=1.665 $X2=0
+ $Y2=0
cc_89 N_A_27_47#_c_86_n N_A_217_131#_c_166_n 0.0123718f $X=1.14 $Y=1.5 $X2=0
+ $Y2=0
cc_90 N_A_27_47#_c_83_n N_A_217_131#_c_169_n 0.0107311f $X=1.23 $Y=1.665 $X2=0
+ $Y2=0
cc_91 N_A_27_47#_c_86_n N_A_217_131#_c_169_n 0.015957f $X=1.14 $Y=1.5 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_M1000_g N_VPWR_c_221_n 0.00357112f $X=1.23 $Y=2.045 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_83_n N_VPWR_c_230_n 0.00266477f $X=1.23 $Y=1.665 $X2=0 $Y2=0
cc_94 N_A_27_47#_M1000_g N_VPWR_c_230_n 0.00325432f $X=1.23 $Y=2.045 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_86_n N_VPWR_c_230_n 0.0247259f $X=1.14 $Y=1.5 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_84_n N_VGND_c_272_n 0.00182475f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_84_n N_VGND_c_273_n 0.00114427f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_85_n N_VGND_c_274_n 0.0162773f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_84_n N_VGND_c_275_n 0.00312914f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_100 N_A_27_47#_M1003_s N_VGND_c_277_n 0.00272496f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_84_n N_VGND_c_277_n 0.0046122f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_85_n N_VGND_c_277_n 0.0110608f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_103 N_B_M1004_g N_A_217_131#_M1002_g 0.0254754f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_104 B N_A_217_131#_M1002_g 2.75921e-19 $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_105 N_B_M1004_g N_A_217_131#_c_164_n 0.00258553f $X=1.785 $Y=0.865 $X2=0
+ $Y2=0
cc_106 N_B_M1004_g N_A_217_131#_c_165_n 0.00332473f $X=1.785 $Y=0.865 $X2=0
+ $Y2=0
cc_107 N_B_M1004_g N_A_217_131#_c_166_n 0.00809176f $X=1.785 $Y=0.865 $X2=0
+ $Y2=0
cc_108 B N_A_217_131#_c_166_n 0.025437f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_109 N_B_c_134_n N_A_217_131#_c_166_n 0.00100048f $X=1.68 $Y=2.58 $X2=0 $Y2=0
cc_110 N_B_M1004_g N_A_217_131#_c_167_n 0.0245645f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_111 N_B_M1004_g N_A_217_131#_c_168_n 0.0213482f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_112 N_B_M1004_g N_A_217_131#_c_170_n 0.0115485f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_113 B N_VPWR_c_221_n 0.0637237f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_114 N_B_c_134_n N_VPWR_c_221_n 0.00210039f $X=1.68 $Y=2.58 $X2=0 $Y2=0
cc_115 N_B_M1004_g N_VPWR_c_222_n 0.0104506f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_116 B N_VPWR_c_222_n 0.0610708f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_117 B N_VPWR_c_230_n 0.00342368f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_118 N_B_M1004_g N_VPWR_c_223_n 7.05206e-19 $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_119 B N_VPWR_c_224_n 0.0551191f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_120 N_B_c_134_n N_VPWR_c_224_n 0.00649446f $X=1.68 $Y=2.58 $X2=0 $Y2=0
cc_121 B N_VPWR_c_220_n 0.029188f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_122 N_B_c_134_n N_VPWR_c_220_n 0.0124362f $X=1.68 $Y=2.58 $X2=0 $Y2=0
cc_123 N_B_M1004_g N_VGND_c_273_n 0.00987464f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_124 N_B_M1004_g N_VGND_c_275_n 0.00332367f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_125 N_B_M1004_g N_VGND_c_277_n 0.00387424f $X=1.785 $Y=0.865 $X2=0 $Y2=0
cc_126 N_A_217_131#_M1002_g N_VPWR_c_222_n 0.0179999f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_A_217_131#_c_166_n N_VPWR_c_230_n 0.0147857f $X=1.53 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_217_131#_M1002_g N_VPWR_c_223_n 0.00974191f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_217_131#_c_166_n N_VPWR_c_223_n 0.00574876f $X=1.53 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_217_131#_c_167_n N_VPWR_c_223_n 0.0260648f $X=2.235 $Y=1.35 $X2=0
+ $Y2=0
cc_131 N_A_217_131#_c_168_n N_VPWR_c_223_n 0.00435746f $X=2.235 $Y=1.35 $X2=0
+ $Y2=0
cc_132 N_A_217_131#_M1002_g N_VPWR_c_225_n 0.00525069f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_217_131#_M1002_g N_VPWR_c_220_n 0.00984971f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_217_131#_M1002_g X 0.0075822f $X=2.345 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_217_131#_M1002_g N_X_c_257_n 0.0073321f $X=2.345 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_217_131#_c_167_n N_X_c_257_n 0.027358f $X=2.235 $Y=1.35 $X2=0 $Y2=0
cc_137 N_A_217_131#_c_170_n N_X_c_257_n 0.0158951f $X=2.257 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A_217_131#_c_164_n N_VGND_c_273_n 0.019202f $X=1.395 $Y=0.86 $X2=0
+ $Y2=0
cc_139 N_A_217_131#_c_167_n N_VGND_c_273_n 0.0354587f $X=2.235 $Y=1.35 $X2=0
+ $Y2=0
cc_140 N_A_217_131#_c_168_n N_VGND_c_273_n 0.00516644f $X=2.235 $Y=1.35 $X2=0
+ $Y2=0
cc_141 N_A_217_131#_c_170_n N_VGND_c_273_n 0.0223584f $X=2.257 $Y=1.185 $X2=0
+ $Y2=0
cc_142 N_A_217_131#_c_164_n N_VGND_c_275_n 0.00759092f $X=1.395 $Y=0.86 $X2=0
+ $Y2=0
cc_143 N_A_217_131#_c_170_n N_VGND_c_276_n 0.00486043f $X=2.257 $Y=1.185 $X2=0
+ $Y2=0
cc_144 N_A_217_131#_c_164_n N_VGND_c_277_n 0.0148387f $X=1.395 $Y=0.86 $X2=0
+ $Y2=0
cc_145 N_A_217_131#_c_170_n N_VGND_c_277_n 0.00921135f $X=2.257 $Y=1.185 $X2=0
+ $Y2=0
cc_146 N_A_217_131#_c_164_n A_300_131# 0.00370499f $X=1.395 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_217_131#_c_165_n A_300_131# 5.60141e-19 $X=1.485 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_148 N_VPWR_c_220_n N_X_M1002_d 0.00336915f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_149 N_VPWR_c_223_n X 0.0178467f $X=2.15 $Y=1.957 $X2=0 $Y2=0
cc_150 N_VPWR_c_225_n X 0.023184f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_151 N_VPWR_c_220_n X 0.0131407f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_152 N_X_c_257_n N_VGND_c_276_n 0.021037f $X=2.585 $Y=0.42 $X2=0 $Y2=0
cc_153 N_X_M1005_d N_VGND_c_277_n 0.00371702f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_154 N_X_c_257_n N_VGND_c_277_n 0.0117799f $X=2.585 $Y=0.42 $X2=0 $Y2=0
