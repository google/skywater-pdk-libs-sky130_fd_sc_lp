* File: sky130_fd_sc_lp__o221a_m.spice
* Created: Wed Sep  2 10:18:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221a_m.pex.spice"
.subckt sky130_fd_sc_lp__o221a_m  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1001 N_A_110_179#_M1001_d N_C1_M1001_g N_A_27_179#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_196_179#_M1009_d N_B1_M1009_g N_A_110_179#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.10245 AS=0.0588 PD=0.92 PS=0.7 NRD=27.132 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_110_179#_M1005_d N_B2_M1005_g N_A_196_179#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.10245 PD=1.37 PS=0.92 NRD=0 NRS=27.132 M=1 R=2.8
+ SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_196_179#_M1007_d N_A2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_196_179#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_27_179#_M1006_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_C1_M1010_g N_A_27_179#_M1010_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09345 AS=0.1113 PD=0.865 PS=1.37 NRD=37.5088 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1003 A_238_535# N_B1_M1003_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.09345 PD=0.63 PS=0.865 NRD=23.443 NRS=39.8531 M=1 R=2.8
+ SA=75000.8 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 N_A_27_179#_M1011_d N_B2_M1011_g A_238_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 A_396_535# N_A2_M1008_g N_A_27_179#_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=49.25 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_396_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06615 AS=0.0672 PD=0.735 PS=0.74 NRD=16.4101 NRS=49.25 M=1 R=2.8 SA=75002
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_27_179#_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.06615 PD=1.37 PS=0.735 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.93145 P=11.27
c_39 VNB 0 2.94581e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o221a_m.pxi.spice"
*
.ends
*
*
