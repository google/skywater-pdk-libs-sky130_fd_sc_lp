* File: sky130_fd_sc_lp__o221ai_m.pxi.spice
* Created: Fri Aug 28 11:09:04 2020
* 
x_PM_SKY130_FD_SC_LP__O221AI_M%C1 N_C1_M1006_g N_C1_c_73_n N_C1_M1000_g
+ N_C1_c_74_n C1 N_C1_c_78_n N_C1_c_75_n PM_SKY130_FD_SC_LP__O221AI_M%C1
x_PM_SKY130_FD_SC_LP__O221AI_M%B1 N_B1_M1005_g N_B1_M1009_g B1 N_B1_c_120_n
+ PM_SKY130_FD_SC_LP__O221AI_M%B1
x_PM_SKY130_FD_SC_LP__O221AI_M%A2 N_A2_M1008_g N_A2_c_165_n N_A2_c_171_n
+ N_A2_M1007_g N_A2_c_166_n N_A2_c_167_n A2 N_A2_c_169_n
+ PM_SKY130_FD_SC_LP__O221AI_M%A2
x_PM_SKY130_FD_SC_LP__O221AI_M%A1 N_A1_M1003_g N_A1_M1001_g A1 A1 N_A1_c_210_n
+ PM_SKY130_FD_SC_LP__O221AI_M%A1
x_PM_SKY130_FD_SC_LP__O221AI_M%B2 N_B2_M1002_g N_B2_c_251_n N_B2_c_252_n
+ N_B2_M1004_g N_B2_c_243_n N_B2_c_244_n N_B2_c_245_n N_B2_c_246_n N_B2_c_247_n
+ B2 N_B2_c_249_n PM_SKY130_FD_SC_LP__O221AI_M%B2
x_PM_SKY130_FD_SC_LP__O221AI_M%Y N_Y_M1000_s N_Y_M1006_s N_Y_M1002_d N_Y_c_300_n
+ N_Y_c_301_n Y Y Y Y Y Y Y N_Y_c_299_n PM_SKY130_FD_SC_LP__O221AI_M%Y
x_PM_SKY130_FD_SC_LP__O221AI_M%VPWR N_VPWR_M1006_d N_VPWR_M1001_d N_VPWR_c_347_n
+ N_VPWR_c_348_n VPWR N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_346_n
+ N_VPWR_c_352_n N_VPWR_c_353_n PM_SKY130_FD_SC_LP__O221AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O221AI_M%A_148_47# N_A_148_47#_M1000_d N_A_148_47#_M1004_d
+ N_A_148_47#_c_383_n N_A_148_47#_c_384_n N_A_148_47#_c_393_n
+ N_A_148_47#_c_385_n N_A_148_47#_c_386_n N_A_148_47#_c_394_n
+ N_A_148_47#_c_387_n N_A_148_47#_c_388_n N_A_148_47#_c_389_n
+ N_A_148_47#_c_390_n N_A_148_47#_c_391_n PM_SKY130_FD_SC_LP__O221AI_M%A_148_47#
x_PM_SKY130_FD_SC_LP__O221AI_M%A_234_47# N_A_234_47#_M1005_d N_A_234_47#_M1003_d
+ N_A_234_47#_c_482_p N_A_234_47#_c_468_n N_A_234_47#_c_469_n
+ N_A_234_47#_c_485_p PM_SKY130_FD_SC_LP__O221AI_M%A_234_47#
x_PM_SKY130_FD_SC_LP__O221AI_M%VGND N_VGND_M1008_d N_VGND_c_491_n VGND
+ N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n
+ PM_SKY130_FD_SC_LP__O221AI_M%VGND
cc_1 VNB N_C1_c_73_n 0.0196633f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.765
cc_2 VNB N_C1_c_74_n 0.0147535f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.84
cc_3 VNB N_C1_c_75_n 0.0391519f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.87
cc_4 VNB N_B1_M1005_g 0.0385969f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.2
cc_5 VNB N_B1_M1009_g 0.00972295f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.765
cc_6 VNB B1 0.00387835f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.445
cc_7 VNB N_B1_c_120_n 0.0319133f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.84
cc_8 VNB N_A2_M1008_g 0.0247607f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.2
cc_9 VNB N_A2_c_165_n 0.00402642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_166_n 0.0198512f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.84
cc_11 VNB N_A2_c_167_n 0.015813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A2 0.0102391f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.035
cc_13 VNB N_A2_c_169_n 0.0155623f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.87
cc_14 VNB N_A1_M1003_g 0.0584328f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.2
cc_15 VNB N_A1_c_210_n 0.030713f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_16 VNB N_B2_c_243_n 0.0284132f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.84
cc_17 VNB N_B2_c_244_n 0.0144116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B2_c_245_n 0.0160076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B2_c_246_n 0.0200258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_c_247_n 0.0252259f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.035
cc_21 VNB B2 0.00559535f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.035
cc_22 VNB N_B2_c_249_n 0.0281825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB Y 0.0470037f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.035
cc_24 VNB N_Y_c_299_n 0.023968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_346_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_148_47#_c_383_n 0.00507353f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.445
cc_27 VNB N_A_148_47#_c_384_n 0.00334285f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.445
cc_28 VNB N_A_148_47#_c_385_n 0.00639664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_148_47#_c_386_n 0.00419975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_148_47#_c_387_n 0.0144415f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.035
cc_31 VNB N_A_148_47#_c_388_n 0.0251381f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.87
cc_32 VNB N_A_148_47#_c_389_n 0.0323518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_148_47#_c_390_n 5.00661e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_148_47#_c_391_n 0.00337993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_234_47#_c_468_n 0.0186344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_234_47#_c_469_n 0.0078256f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.84
cc_37 VNB N_VGND_c_491_n 0.00295613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_492_n 0.0451014f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.84
cc_39 VNB N_VGND_c_493_n 0.039448f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.2
cc_40 VNB N_VGND_c_494_n 0.195391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_495_n 0.00521963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_C1_M1006_g 0.0266489f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.61
cc_43 VPB C1 0.00343327f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_44 VPB N_C1_c_78_n 0.0336782f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.035
cc_45 VPB N_C1_c_75_n 0.0126965f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.87
cc_46 VPB N_B1_M1009_g 0.0548904f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.765
cc_47 VPB N_A2_c_165_n 0.0622258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_c_171_n 0.0185163f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.765
cc_49 VPB N_A1_M1001_g 0.0199946f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.765
cc_50 VPB A1 0.0101455f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.84
cc_51 VPB N_A1_c_210_n 0.0739956f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_52 VPB N_B2_M1002_g 0.0314433f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.2
cc_53 VPB N_B2_c_251_n 0.129798f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.61
cc_54 VPB N_B2_c_252_n 0.0125602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B2_c_245_n 0.118577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_Y_c_300_n 0.00957889f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.84
cc_57 VPB N_Y_c_301_n 0.00204748f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.84
cc_58 VPB Y 0.0314563f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.035
cc_59 VPB Y 0.034492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_347_n 0.017813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_348_n 0.0185424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_349_n 0.0457835f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.87
cc_63 VPB N_VPWR_c_350_n 0.0166893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_346_n 0.058224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_352_n 0.0289906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_353_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_148_47#_c_384_n 0.00385767f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=0.445
cc_68 VPB N_A_148_47#_c_393_n 3.76099e-19 $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.84
cc_69 VPB N_A_148_47#_c_394_n 0.0215006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_148_47#_c_387_n 0.0048254f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.035
cc_71 VPB N_A_148_47#_c_390_n 0.00215312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_148_47#_c_391_n 0.00395637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 N_C1_c_73_n N_B1_M1005_g 0.0200586f $X=0.665 $Y=0.765 $X2=0 $Y2=0
cc_74 N_C1_c_75_n N_B1_M1005_g 0.00678379f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_75 N_C1_M1006_g N_B1_M1009_g 0.0202885f $X=0.6 $Y=2.61 $X2=0 $Y2=0
cc_76 C1 N_B1_M1009_g 0.00109107f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_77 N_C1_c_78_n N_B1_M1009_g 0.01854f $X=0.67 $Y=2.035 $X2=0 $Y2=0
cc_78 N_C1_c_75_n N_B1_M1009_g 0.009665f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_79 N_C1_c_75_n B1 2.20889e-19 $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_80 N_C1_c_75_n N_B1_c_120_n 0.0177733f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_81 N_C1_M1006_g N_Y_c_300_n 0.0125506f $X=0.6 $Y=2.61 $X2=0 $Y2=0
cc_82 C1 N_Y_c_300_n 0.0220435f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_83 N_C1_c_78_n N_Y_c_300_n 0.00449327f $X=0.67 $Y=2.035 $X2=0 $Y2=0
cc_84 N_C1_M1006_g Y 0.00328159f $X=0.6 $Y=2.61 $X2=0 $Y2=0
cc_85 N_C1_c_73_n Y 0.00174965f $X=0.665 $Y=0.765 $X2=0 $Y2=0
cc_86 N_C1_c_74_n Y 0.0266369f $X=0.665 $Y=0.84 $X2=0 $Y2=0
cc_87 C1 Y 0.0121505f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_88 N_C1_c_78_n Y 0.00417986f $X=0.67 $Y=2.035 $X2=0 $Y2=0
cc_89 N_C1_M1006_g Y 0.00251674f $X=0.6 $Y=2.61 $X2=0 $Y2=0
cc_90 N_C1_c_73_n N_Y_c_299_n 4.52635e-19 $X=0.665 $Y=0.765 $X2=0 $Y2=0
cc_91 N_C1_c_74_n N_Y_c_299_n 0.00223206f $X=0.665 $Y=0.84 $X2=0 $Y2=0
cc_92 N_C1_M1006_g N_VPWR_c_347_n 0.00405893f $X=0.6 $Y=2.61 $X2=0 $Y2=0
cc_93 N_C1_M1006_g N_VPWR_c_346_n 0.00502397f $X=0.6 $Y=2.61 $X2=0 $Y2=0
cc_94 N_C1_M1006_g N_VPWR_c_352_n 0.00481372f $X=0.6 $Y=2.61 $X2=0 $Y2=0
cc_95 N_C1_c_74_n N_A_148_47#_c_383_n 3.52987e-19 $X=0.665 $Y=0.84 $X2=0 $Y2=0
cc_96 N_C1_c_75_n N_A_148_47#_c_383_n 0.013138f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_97 C1 N_A_148_47#_c_384_n 0.00770913f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_98 N_C1_c_78_n N_A_148_47#_c_384_n 0.00290733f $X=0.67 $Y=2.035 $X2=0 $Y2=0
cc_99 C1 N_A_148_47#_c_393_n 0.0118705f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_100 N_C1_c_78_n N_A_148_47#_c_393_n 0.00160526f $X=0.67 $Y=2.035 $X2=0 $Y2=0
cc_101 N_C1_c_75_n N_A_148_47#_c_393_n 0.00708073f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_102 N_C1_c_74_n N_A_148_47#_c_385_n 0.00776884f $X=0.665 $Y=0.84 $X2=0 $Y2=0
cc_103 N_C1_c_75_n N_A_148_47#_c_385_n 0.003777f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_104 N_C1_c_73_n N_A_148_47#_c_386_n 0.00234158f $X=0.665 $Y=0.765 $X2=0 $Y2=0
cc_105 N_C1_c_75_n N_A_148_47#_c_390_n 0.00190797f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_106 N_C1_c_73_n N_VGND_c_492_n 0.00585385f $X=0.665 $Y=0.765 $X2=0 $Y2=0
cc_107 N_C1_c_74_n N_VGND_c_492_n 7.30493e-19 $X=0.665 $Y=0.84 $X2=0 $Y2=0
cc_108 N_C1_c_73_n N_VGND_c_494_n 0.00776234f $X=0.665 $Y=0.765 $X2=0 $Y2=0
cc_109 N_C1_c_74_n N_VGND_c_494_n 9.35314e-19 $X=0.665 $Y=0.84 $X2=0 $Y2=0
cc_110 N_B1_M1005_g N_A2_M1008_g 0.0299292f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_111 N_B1_M1009_g N_A2_c_165_n 0.0184391f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_112 B1 N_A2_c_166_n 6.81367e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B1_c_120_n N_A2_c_166_n 0.0119336f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_114 N_B1_M1009_g N_A2_c_167_n 0.0119336f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_115 N_B1_M1005_g A2 8.99677e-19 $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_116 B1 A2 0.0149667f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_c_120_n A2 0.00129363f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_118 N_B1_M1009_g N_B2_M1002_g 0.0428502f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_119 N_B1_M1009_g N_Y_c_300_n 0.0133584f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_120 N_B1_M1009_g N_VPWR_c_347_n 0.00480551f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_121 N_B1_M1009_g N_VPWR_c_349_n 0.00481372f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_122 N_B1_M1009_g N_VPWR_c_346_n 0.00502397f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_123 N_B1_M1005_g N_A_148_47#_c_383_n 0.00228277f $X=1.095 $Y=0.445 $X2=0
+ $Y2=0
cc_124 N_B1_M1009_g N_A_148_47#_c_383_n 0.00173517f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_125 B1 N_A_148_47#_c_383_n 0.0141376f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B1_c_120_n N_A_148_47#_c_383_n 0.00340759f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_127 N_B1_M1009_g N_A_148_47#_c_384_n 4.53217e-19 $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_128 B1 N_A_148_47#_c_384_n 0.00830414f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B1_c_120_n N_A_148_47#_c_384_n 0.00293883f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_130 N_B1_M1005_g N_A_148_47#_c_385_n 0.00454203f $X=1.095 $Y=0.445 $X2=0
+ $Y2=0
cc_131 B1 N_A_148_47#_c_385_n 0.00622833f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_c_120_n N_A_148_47#_c_385_n 0.0021393f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_133 N_B1_M1005_g N_A_148_47#_c_386_n 0.00249464f $X=1.095 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_B1_M1009_g N_A_148_47#_c_394_n 0.00544601f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_135 B1 N_A_148_47#_c_394_n 0.00506762f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B1_M1009_g N_A_148_47#_c_390_n 0.0110396f $X=1.15 $Y=2.61 $X2=0 $Y2=0
cc_137 B1 N_A_148_47#_c_390_n 0.0116879f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B1_c_120_n N_A_148_47#_c_390_n 0.00169785f $X=1.06 $Y=1.32 $X2=0 $Y2=0
cc_139 N_B1_M1005_g N_A_234_47#_c_469_n 0.00154608f $X=1.095 $Y=0.445 $X2=0
+ $Y2=0
cc_140 B1 N_A_234_47#_c_469_n 0.0029782f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B1_M1005_g N_VGND_c_491_n 0.00145442f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_142 N_B1_M1005_g N_VGND_c_492_n 0.00585385f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_143 N_B1_M1005_g N_VGND_c_494_n 0.0110741f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A2_M1008_g N_A1_M1003_g 0.0173557f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_145 A2 N_A1_M1003_g 0.00329485f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A2_c_169_n N_A1_M1003_g 0.0190056f $X=1.63 $Y=1.08 $X2=0 $Y2=0
cc_147 N_A2_c_171_n N_A1_M1001_g 0.0260663f $X=2.13 $Y=2.195 $X2=0 $Y2=0
cc_148 N_A2_c_165_n A1 0.00117758f $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_149 N_A2_c_165_n N_A1_c_210_n 0.0423429f $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_150 N_A2_c_167_n N_A1_c_210_n 0.0190056f $X=1.63 $Y=1.585 $X2=0 $Y2=0
cc_151 N_A2_c_171_n N_B2_M1002_g 0.0142133f $X=2.13 $Y=2.195 $X2=0 $Y2=0
cc_152 N_A2_c_167_n N_B2_M1002_g 0.00145966f $X=1.63 $Y=1.585 $X2=0 $Y2=0
cc_153 N_A2_c_171_n N_B2_c_251_n 0.0104164f $X=2.13 $Y=2.195 $X2=0 $Y2=0
cc_154 N_A2_c_165_n N_Y_c_300_n 0.00181864f $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_155 N_A2_c_165_n N_Y_c_301_n 0.00576052f $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_156 N_A2_c_171_n N_Y_c_301_n 0.0064698f $X=2.13 $Y=2.195 $X2=0 $Y2=0
cc_157 N_A2_c_171_n N_VPWR_c_348_n 0.00160648f $X=2.13 $Y=2.195 $X2=0 $Y2=0
cc_158 N_A2_c_171_n N_VPWR_c_346_n 9.39239e-19 $X=2.13 $Y=2.195 $X2=0 $Y2=0
cc_159 A2 N_A_148_47#_c_385_n 0.00123049f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_c_165_n N_A_148_47#_c_394_n 0.0173575f $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_161 N_A2_c_167_n N_A_148_47#_c_394_n 0.00340572f $X=1.63 $Y=1.585 $X2=0 $Y2=0
cc_162 A2 N_A_148_47#_c_394_n 0.0240026f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A2_c_165_n N_A_148_47#_c_387_n 8.94941e-19 $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_164 N_A2_c_165_n N_A_148_47#_c_390_n 6.29426e-19 $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_165 N_A2_c_165_n N_A_148_47#_c_391_n 0.00517933f $X=1.72 $Y=1.88 $X2=0 $Y2=0
cc_166 N_A2_c_167_n N_A_148_47#_c_391_n 0.00311607f $X=1.63 $Y=1.585 $X2=0 $Y2=0
cc_167 N_A2_M1008_g N_A_234_47#_c_468_n 0.011968f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_168 A2 N_A_234_47#_c_468_n 0.0240026f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_169 N_A2_c_169_n N_A_234_47#_c_468_n 0.00516074f $X=1.63 $Y=1.08 $X2=0 $Y2=0
cc_170 N_A2_M1008_g N_VGND_c_491_n 0.00733493f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_171 N_A2_M1008_g N_VGND_c_492_n 0.00411627f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_172 N_A2_M1008_g N_VGND_c_494_n 0.00485622f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_173 N_A1_M1001_g N_B2_c_251_n 0.0103107f $X=2.49 $Y=2.525 $X2=0 $Y2=0
cc_174 A1 N_B2_c_243_n 4.13063e-19 $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_175 N_A1_c_210_n N_B2_c_244_n 0.0178838f $X=2.49 $Y=1.812 $X2=0 $Y2=0
cc_176 N_A1_M1001_g N_B2_c_245_n 0.0121916f $X=2.49 $Y=2.525 $X2=0 $Y2=0
cc_177 A1 N_B2_c_245_n 0.020754f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_178 N_A1_c_210_n N_B2_c_245_n 0.0283117f $X=2.49 $Y=1.812 $X2=0 $Y2=0
cc_179 N_A1_M1003_g N_B2_c_246_n 0.0212854f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A1_M1003_g B2 0.00903615f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A1_c_210_n B2 3.62699e-19 $X=2.49 $Y=1.812 $X2=0 $Y2=0
cc_182 N_A1_M1003_g N_B2_c_249_n 0.015258f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A1_M1001_g N_VPWR_c_348_n 0.00941814f $X=2.49 $Y=2.525 $X2=0 $Y2=0
cc_184 A1 N_VPWR_c_348_n 0.0132576f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_185 N_A1_c_210_n N_VPWR_c_348_n 0.00651838f $X=2.49 $Y=1.812 $X2=0 $Y2=0
cc_186 N_A1_M1001_g N_VPWR_c_346_n 7.88961e-19 $X=2.49 $Y=2.525 $X2=0 $Y2=0
cc_187 A1 N_A_148_47#_c_387_n 0.0472861f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_188 N_A1_c_210_n N_A_148_47#_c_387_n 0.0406637f $X=2.49 $Y=1.812 $X2=0 $Y2=0
cc_189 N_A1_c_210_n N_A_148_47#_c_391_n 0.0124151f $X=2.49 $Y=1.812 $X2=0 $Y2=0
cc_190 N_A1_M1003_g N_A_234_47#_c_468_n 0.0163964f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A1_c_210_n N_A_234_47#_c_468_n 0.00369144f $X=2.49 $Y=1.812 $X2=0 $Y2=0
cc_192 N_A1_M1003_g N_VGND_c_491_n 0.00668353f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A1_M1003_g N_VGND_c_493_n 0.00426565f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A1_M1003_g N_VGND_c_494_n 0.00641576f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_195 N_B2_M1002_g N_Y_c_300_n 0.0112432f $X=1.51 $Y=2.61 $X2=0 $Y2=0
cc_196 N_B2_c_251_n N_Y_c_300_n 8.72066e-19 $X=3.105 $Y=3.15 $X2=0 $Y2=0
cc_197 N_B2_M1002_g N_Y_c_301_n 0.00428066f $X=1.51 $Y=2.61 $X2=0 $Y2=0
cc_198 N_B2_c_251_n N_Y_c_301_n 0.00363378f $X=3.105 $Y=3.15 $X2=0 $Y2=0
cc_199 N_B2_M1002_g N_VPWR_c_347_n 0.00742769f $X=1.51 $Y=2.61 $X2=0 $Y2=0
cc_200 N_B2_c_251_n N_VPWR_c_348_n 0.0252552f $X=3.105 $Y=3.15 $X2=0 $Y2=0
cc_201 N_B2_c_245_n N_VPWR_c_348_n 0.0132802f $X=3.18 $Y=3.075 $X2=0 $Y2=0
cc_202 N_B2_c_252_n N_VPWR_c_349_n 0.0377651f $X=1.585 $Y=3.15 $X2=0 $Y2=0
cc_203 N_B2_c_251_n N_VPWR_c_350_n 0.0144454f $X=3.105 $Y=3.15 $X2=0 $Y2=0
cc_204 N_B2_c_251_n N_VPWR_c_346_n 0.0610154f $X=3.105 $Y=3.15 $X2=0 $Y2=0
cc_205 N_B2_c_252_n N_VPWR_c_346_n 0.00720651f $X=1.585 $Y=3.15 $X2=0 $Y2=0
cc_206 N_B2_M1002_g N_A_148_47#_c_394_n 0.00184437f $X=1.51 $Y=2.61 $X2=0 $Y2=0
cc_207 N_B2_c_244_n N_A_148_47#_c_387_n 0.00979365f $X=2.905 $Y=1.36 $X2=0 $Y2=0
cc_208 N_B2_c_245_n N_A_148_47#_c_387_n 0.012322f $X=3.18 $Y=3.075 $X2=0 $Y2=0
cc_209 N_B2_c_247_n N_A_148_47#_c_387_n 0.00242404f $X=2.685 $Y=0.915 $X2=0
+ $Y2=0
cc_210 B2 N_A_148_47#_c_387_n 0.0261287f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_211 N_B2_c_243_n N_A_148_47#_c_388_n 0.00414561f $X=3.105 $Y=1.36 $X2=0 $Y2=0
cc_212 N_B2_c_247_n N_A_148_47#_c_388_n 0.00730375f $X=2.685 $Y=0.915 $X2=0
+ $Y2=0
cc_213 B2 N_A_148_47#_c_388_n 0.0194174f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_214 N_B2_c_243_n N_A_148_47#_c_389_n 0.0166908f $X=3.105 $Y=1.36 $X2=0 $Y2=0
cc_215 N_B2_c_245_n N_A_148_47#_c_389_n 0.00507336f $X=3.18 $Y=3.075 $X2=0 $Y2=0
cc_216 N_B2_c_246_n N_A_148_47#_c_389_n 0.00259723f $X=2.685 $Y=0.765 $X2=0
+ $Y2=0
cc_217 N_B2_c_247_n N_A_148_47#_c_389_n 0.0128638f $X=2.685 $Y=0.915 $X2=0 $Y2=0
cc_218 B2 N_A_148_47#_c_389_n 0.0369045f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_219 N_B2_c_246_n N_A_234_47#_c_468_n 0.00481511f $X=2.685 $Y=0.765 $X2=0
+ $Y2=0
cc_220 N_B2_c_246_n N_VGND_c_493_n 0.00585385f $X=2.685 $Y=0.765 $X2=0 $Y2=0
cc_221 N_B2_c_247_n N_VGND_c_493_n 8.58906e-19 $X=2.685 $Y=0.915 $X2=0 $Y2=0
cc_222 N_B2_c_246_n N_VGND_c_494_n 0.0106575f $X=2.685 $Y=0.765 $X2=0 $Y2=0
cc_223 N_B2_c_247_n N_VGND_c_494_n 9.24424e-19 $X=2.685 $Y=0.915 $X2=0 $Y2=0
cc_224 B2 N_VGND_c_494_n 0.00340038f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_225 N_Y_c_300_n N_VPWR_M1006_d 0.00322761f $X=1.715 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_226 N_Y_c_300_n N_VPWR_c_347_n 0.0217579f $X=1.715 $Y=2.385 $X2=0 $Y2=0
cc_227 Y N_VPWR_c_347_n 0.00271111f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_228 N_Y_c_301_n N_VPWR_c_348_n 0.00392982f $X=1.82 $Y=2.385 $X2=0 $Y2=0
cc_229 N_Y_c_301_n N_VPWR_c_349_n 0.0033189f $X=1.82 $Y=2.385 $X2=0 $Y2=0
cc_230 N_Y_c_300_n N_VPWR_c_346_n 0.0288832f $X=1.715 $Y=2.385 $X2=0 $Y2=0
cc_231 N_Y_c_301_n N_VPWR_c_346_n 0.00500735f $X=1.82 $Y=2.385 $X2=0 $Y2=0
cc_232 Y N_VPWR_c_346_n 0.011332f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_233 Y N_VPWR_c_352_n 0.00991568f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_234 N_Y_c_300_n A_245_480# 0.00196273f $X=1.715 $Y=2.385 $X2=-0.19 $Y2=-0.245
cc_235 Y N_A_148_47#_c_383_n 0.0327119f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_236 N_Y_c_300_n N_A_148_47#_c_384_n 0.00604482f $X=1.715 $Y=2.385 $X2=0 $Y2=0
cc_237 Y N_A_148_47#_c_393_n 0.0108635f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_238 Y N_A_148_47#_c_385_n 0.0106456f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_239 N_Y_c_299_n N_A_148_47#_c_385_n 6.9e-19 $X=0.45 $Y=0.51 $X2=0 $Y2=0
cc_240 Y N_A_148_47#_c_386_n 0.00718018f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_241 N_Y_c_299_n N_A_148_47#_c_386_n 0.00123132f $X=0.45 $Y=0.51 $X2=0 $Y2=0
cc_242 N_Y_c_300_n N_A_148_47#_c_394_n 0.0193744f $X=1.715 $Y=2.385 $X2=0 $Y2=0
cc_243 N_Y_c_301_n N_A_148_47#_c_394_n 0.00815385f $X=1.82 $Y=2.385 $X2=0 $Y2=0
cc_244 N_Y_c_300_n N_A_148_47#_c_390_n 0.0058965f $X=1.715 $Y=2.385 $X2=0 $Y2=0
cc_245 N_Y_c_299_n N_VGND_c_492_n 0.0165677f $X=0.45 $Y=0.51 $X2=0 $Y2=0
cc_246 N_Y_M1000_s N_VGND_c_494_n 0.00247303f $X=0.325 $Y=0.235 $X2=0 $Y2=0
cc_247 N_Y_c_299_n N_VGND_c_494_n 0.014467f $X=0.45 $Y=0.51 $X2=0 $Y2=0
cc_248 N_A_148_47#_c_388_n N_A_234_47#_c_468_n 2.31889e-19 $X=3.085 $Y=0.495
+ $X2=0 $Y2=0
cc_249 N_A_148_47#_c_386_n N_A_234_47#_c_469_n 0.0108396f $X=0.88 $Y=0.51 $X2=0
+ $Y2=0
cc_250 N_A_148_47#_c_386_n N_VGND_c_492_n 0.00819826f $X=0.88 $Y=0.51 $X2=0
+ $Y2=0
cc_251 N_A_148_47#_c_388_n N_VGND_c_493_n 0.0274761f $X=3.085 $Y=0.495 $X2=0
+ $Y2=0
cc_252 N_A_148_47#_M1000_d N_VGND_c_494_n 0.00377351f $X=0.74 $Y=0.235 $X2=0
+ $Y2=0
cc_253 N_A_148_47#_M1004_d N_VGND_c_494_n 0.00244275f $X=2.615 $Y=0.235 $X2=0
+ $Y2=0
cc_254 N_A_148_47#_c_385_n N_VGND_c_494_n 0.00636528f $X=0.88 $Y=0.86 $X2=0
+ $Y2=0
cc_255 N_A_148_47#_c_386_n N_VGND_c_494_n 0.0076345f $X=0.88 $Y=0.51 $X2=0 $Y2=0
cc_256 N_A_148_47#_c_388_n N_VGND_c_494_n 0.0222317f $X=3.085 $Y=0.495 $X2=0
+ $Y2=0
cc_257 N_A_234_47#_c_468_n N_VGND_M1008_d 0.00349577f $X=2.205 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_258 N_A_234_47#_c_468_n N_VGND_c_491_n 0.0196407f $X=2.205 $Y=0.73 $X2=0
+ $Y2=0
cc_259 N_A_234_47#_c_482_p N_VGND_c_492_n 0.00845107f $X=1.325 $Y=0.51 $X2=0
+ $Y2=0
cc_260 N_A_234_47#_c_468_n N_VGND_c_492_n 0.00263146f $X=2.205 $Y=0.73 $X2=0
+ $Y2=0
cc_261 N_A_234_47#_c_468_n N_VGND_c_493_n 0.00376082f $X=2.205 $Y=0.73 $X2=0
+ $Y2=0
cc_262 N_A_234_47#_c_485_p N_VGND_c_493_n 0.00903611f $X=2.325 $Y=0.495 $X2=0
+ $Y2=0
cc_263 N_A_234_47#_M1005_d N_VGND_c_494_n 0.00433181f $X=1.17 $Y=0.235 $X2=0
+ $Y2=0
cc_264 N_A_234_47#_M1003_d N_VGND_c_494_n 0.00361939f $X=2.185 $Y=0.235 $X2=0
+ $Y2=0
cc_265 N_A_234_47#_c_482_p N_VGND_c_494_n 0.00761208f $X=1.325 $Y=0.51 $X2=0
+ $Y2=0
cc_266 N_A_234_47#_c_468_n N_VGND_c_494_n 0.0126592f $X=2.205 $Y=0.73 $X2=0
+ $Y2=0
cc_267 N_A_234_47#_c_485_p N_VGND_c_494_n 0.00822141f $X=2.325 $Y=0.495 $X2=0
+ $Y2=0
