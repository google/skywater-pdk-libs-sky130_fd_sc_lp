* File: sky130_fd_sc_lp__nor4bb_4.spice
* Created: Wed Sep  2 10:11:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4bb_4.pex.spice"
.subckt sky130_fd_sc_lp__nor4bb_4  VNB VPB D_N C_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_D_N_M1015_g N_A_37_51#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1028 N_A_206_51#_M1028_d N_C_N_M1028_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A_37_51#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2814 AS=0.1176 PD=2.35 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.3
+ SB=75007.3 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_37_51#_M1009_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.189 AS=0.1176 PD=1.29 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75006.8 A=0.126 P=1.98 MULT=1
MM1026 N_VGND_M1009_d N_A_37_51#_M1026_g N_Y_M1026_s VNB NSHORT L=0.15 W=0.84
+ AD=0.189 AS=0.1176 PD=1.29 PS=1.12 NRD=12.852 NRS=0 M=1 R=5.6 SA=75001.3
+ SB=75006.2 A=0.126 P=1.98 MULT=1
MM1029 N_VGND_M1029_d N_A_37_51#_M1029_g N_Y_M1026_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75005.8 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A_206_51#_M1000_g N_VGND_M1029_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75002.2 SB=75005.3
+ A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1000_d N_A_206_51#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75004.9 A=0.126 P=1.98 MULT=1
MM1022 N_Y_M1022_d N_A_206_51#_M1022_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1034 N_Y_M1022_d N_A_206_51#_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2793 PD=1.12 PS=1.505 NRD=0 NRS=0 M=1 R=5.6 SA=75003.5 SB=75004
+ A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1034_s N_B_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.84 AD=0.2793
+ AS=0.1176 PD=1.505 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.3 SB=75003.2 A=0.126
+ P=1.98 MULT=1
MM1023 N_VGND_M1023_d N_B_M1023_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.8 SB=75002.8 A=0.126
+ P=1.98 MULT=1
MM1024 N_VGND_M1023_d N_B_M1024_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.2 SB=75002.3 A=0.126
+ P=1.98 MULT=1
MM1035 N_VGND_M1035_d N_B_M1035_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.6 SB=75001.9 A=0.126
+ P=1.98 MULT=1
MM1016 N_Y_M1016_d N_A_M1016_g N_VGND_M1035_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006 SB=75001.5 A=0.126
+ P=1.98 MULT=1
MM1017 N_Y_M1016_d N_A_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.5 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.9 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1031 N_Y_M1018_d N_A_M1031_g N_VGND_M1031_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75007.3 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1032 N_VPWR_M1032_d N_D_N_M1032_g N_A_37_51#_M1032_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_206_51#_M1010_d N_C_N_M1010_g N_VPWR_M1032_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_347_349#_M1005_d N_A_37_51#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1012 N_A_347_349#_M1012_d N_A_37_51#_M1012_g N_Y_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1019 N_A_347_349#_M1012_d N_A_37_51#_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1030 N_A_347_349#_M1030_d N_A_37_51#_M1030_g N_Y_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1001 N_A_774_349#_M1001_d N_A_206_51#_M1001_g N_A_347_349#_M1030_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1007 N_A_774_349#_M1001_d N_A_206_51#_M1007_g N_A_347_349#_M1007_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_A_774_349#_M1013_d N_A_206_51#_M1013_g N_A_347_349#_M1007_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_A_774_349#_M1013_d N_A_206_51#_M1027_g N_A_347_349#_M1027_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1008 N_A_1139_367#_M1008_d N_B_M1008_g N_A_774_349#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1014 N_A_1139_367#_M1014_d N_B_M1014_g N_A_774_349#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1021 N_A_1139_367#_M1014_d N_B_M1021_g N_A_774_349#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1033 N_A_1139_367#_M1033_d N_B_M1033_g N_A_774_349#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.17955 AS=0.1764 PD=1.545 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_1139_367#_M1033_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.17955 PD=1.54 PS=1.545 NRD=0 NRS=0.7683 M=1 R=8.4
+ SA=75001.9 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1003_d N_A_M1011_g N_A_1139_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g N_A_1139_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1020_d N_A_M1025_g N_A_1139_367#_M1025_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref VNB VPB NWDIODE A=18.9772 P=23.87
*
.include "sky130_fd_sc_lp__nor4bb_4.pxi.spice"
*
.ends
*
*
