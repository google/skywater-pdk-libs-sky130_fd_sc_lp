* File: sky130_fd_sc_lp__sdfxbp_1.pex.spice
* Created: Wed Sep  2 10:36:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%SCD 3 7 11 13 14 15 16 21
c26 13 0 1.7997e-19 $X=0.385 $Y=1.88
r27 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.375 $X2=0.385 $Y2=1.375
r28 15 16 9.51718 $w=4.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=2.035
r29 15 22 7.45941 $w=4.63e-07 $l=2.9e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=1.375
r30 14 22 2.05777 $w=4.63e-07 $l=8e-08 $layer=LI1_cond $X=0.317 $Y=1.295
+ $X2=0.317 $Y2=1.375
r31 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.715
+ $X2=0.385 $Y2=1.375
r32 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.715
+ $X2=0.385 $Y2=1.88
r33 11 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.385 $Y=1.36
+ $X2=0.385 $Y2=1.375
r34 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.42 $Y=1.21
+ $X2=0.42 $Y2=1.36
r35 7 10 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.545 $Y=0.805
+ $X2=0.545 $Y2=1.21
r36 3 13 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.475 $Y=2.735
+ $X2=0.475 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%D 3 7 11 12 13 14 18 19
r34 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.355
+ $Y=1.44 $X2=1.355 $Y2=1.44
r35 13 14 8.85098 $w=4.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.27 $Y=1.665
+ $X2=1.27 $Y2=2.035
r36 13 19 5.38235 $w=4.98e-07 $l=2.25e-07 $layer=LI1_cond $X=1.27 $Y=1.665
+ $X2=1.27 $Y2=1.44
r37 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.355 $Y=1.78
+ $X2=1.355 $Y2=1.44
r38 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.78
+ $X2=1.355 $Y2=1.945
r39 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.275
+ $X2=1.355 $Y2=1.44
r40 7 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.445 $Y=0.805 $X2=1.445
+ $Y2=1.275
r41 3 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.265 $Y=2.735
+ $X2=1.265 $Y2=1.945
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_324_431# 1 2 7 9 12 14 20 21 28
c56 28 0 1.86861e-19 $X=2.7 $Y=0.805
r57 26 28 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.45 $Y=0.805
+ $X2=2.7 $Y2=0.805
r58 20 23 43.3074 $w=2.08e-07 $l=8.2e-07 $layer=LI1_cond $X=2.7 $Y=1.74 $X2=2.7
+ $Y2=2.56
r59 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.69
+ $Y=1.74 $X2=2.69 $Y2=1.74
r60 18 28 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=0.97 $X2=2.7
+ $Y2=0.805
r61 18 20 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=2.7 $Y=0.97 $X2=2.7
+ $Y2=1.74
r62 17 21 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=2.69 $Y=2.155
+ $X2=2.69 $Y2=1.74
r63 15 16 13.2911 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.92 $Y=2.23
+ $X2=1.77 $Y2=2.23
r64 14 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.525 $Y=2.23
+ $X2=2.69 $Y2=2.155
r65 14 15 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.525 $Y=2.23
+ $X2=1.92 $Y2=2.23
r66 10 16 64.739 $w=2.35e-07 $l=3.01993e-07 $layer=POLY_cond $X=1.805 $Y=1.945
+ $X2=1.77 $Y2=2.23
r67 10 12 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=1.805 $Y=1.945
+ $X2=1.805 $Y2=0.805
r68 7 16 21.6667 $w=2.35e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.695 $Y=2.305
+ $X2=1.77 $Y2=2.23
r69 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.695 $Y=2.305
+ $X2=1.695 $Y2=2.735
r70 2 23 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=2.405 $X2=2.71 $Y2=2.56
r71 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.595 $X2=2.45 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%SCE 3 5 7 8 11 13 17 19 22 23 24 25 30 31
c75 17 0 1.86861e-19 $X=3.18 $Y=2.725
r76 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=0.43 $X2=3.09 $Y2=0.43
r77 24 25 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.095 $Y=0.925
+ $X2=3.095 $Y2=1.295
r78 23 24 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.095 $Y=0.555
+ $X2=3.095 $Y2=0.925
r79 23 31 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=0.555
+ $X2=3.095 $Y2=0.43
r80 21 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.09 $Y=0.77
+ $X2=3.09 $Y2=0.43
r81 21 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.77
+ $X2=3.09 $Y2=0.935
r82 20 30 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.09 $Y=0.255
+ $X2=3.09 $Y2=0.43
r83 17 22 917.851 $w=1.5e-07 $l=1.79e-06 $layer=POLY_cond $X=3.18 $Y=2.725
+ $X2=3.18 $Y2=0.935
r84 14 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=0.18
+ $X2=2.235 $Y2=0.18
r85 13 20 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.925 $Y=0.18
+ $X2=3.09 $Y2=0.255
r86 13 14 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.925 $Y=0.18
+ $X2=2.31 $Y2=0.18
r87 9 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.235 $Y=0.255
+ $X2=2.235 $Y2=0.18
r88 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.235 $Y=0.255
+ $X2=2.235 $Y2=0.805
r89 7 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=0.18
+ $X2=2.235 $Y2=0.18
r90 7 8 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=2.16 $Y=0.18 $X2=0.98
+ $Y2=0.18
r91 3 5 989.638 $w=1.5e-07 $l=1.93e-06 $layer=POLY_cond $X=0.905 $Y=0.805
+ $X2=0.905 $Y2=2.735
r92 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=0.255
+ $X2=0.98 $Y2=0.18
r93 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.905 $Y=0.255
+ $X2=0.905 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_767_121# 1 2 3 4 15 19 21 23 25 27 30 31
+ 32 34 35 39 45 46 50 52
c135 39 0 1.79277e-19 $X=10.125 $Y=2.04
c136 32 0 1.7373e-19 $X=6.735 $Y=2.43
c137 15 0 1.75353e-19 $X=4.795 $Y=2.335
r138 47 50 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=9.17 $Y=0.835
+ $X2=9.48 $Y2=0.835
r139 45 53 13.8594 $w=3.13e-07 $l=9e-08 $layer=POLY_cond $X=4.885 $Y=1.75
+ $X2=4.795 $Y2=1.75
r140 44 46 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.885 $Y=1.95
+ $X2=5.05 $Y2=1.95
r141 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.77 $X2=4.885 $Y2=1.77
r142 37 39 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=10.135 $Y=2.345
+ $X2=10.135 $Y2=2.04
r143 36 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=2.43
+ $X2=9.17 $Y2=2.43
r144 35 37 6.91519 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=10.02 $Y=2.43
+ $X2=10.135 $Y2=2.345
r145 35 36 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=10.02 $Y=2.43
+ $X2=9.255 $Y2=2.43
r146 34 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.17 $Y=2.345
+ $X2=9.17 $Y2=2.43
r147 33 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.17 $Y=1 $X2=9.17
+ $Y2=0.835
r148 33 34 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=9.17 $Y=1
+ $X2=9.17 $Y2=2.345
r149 31 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.085 $Y=2.43
+ $X2=9.17 $Y2=2.43
r150 31 32 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=9.085 $Y=2.43
+ $X2=6.735 $Y2=2.43
r151 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.65 $Y=2.345
+ $X2=6.735 $Y2=2.43
r152 29 30 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=6.65 $Y=1.855
+ $X2=6.65 $Y2=2.345
r153 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.565 $Y=1.77
+ $X2=6.65 $Y2=1.855
r154 27 46 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=6.565 $Y=1.77
+ $X2=5.05 $Y2=1.77
r155 26 42 2.63167 $w=5.3e-07 $l=1.35e-07 $layer=LI1_cond $X=4.065 $Y=1.95
+ $X2=3.93 $Y2=1.95
r156 25 44 2.25675 $w=5.28e-07 $l=1e-07 $layer=LI1_cond $X=4.785 $Y=1.95
+ $X2=4.885 $Y2=1.95
r157 25 26 16.2486 $w=5.28e-07 $l=7.2e-07 $layer=LI1_cond $X=4.785 $Y=1.95
+ $X2=4.065 $Y2=1.95
r158 21 42 5.16588 $w=2.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.93 $Y=1.685
+ $X2=3.93 $Y2=1.95
r159 21 23 38.6282 $w=2.68e-07 $l=9.05e-07 $layer=LI1_cond $X=3.93 $Y=1.685
+ $X2=3.93 $Y2=0.78
r160 17 45 31.5687 $w=3.13e-07 $l=2.82754e-07 $layer=POLY_cond $X=5.09 $Y=1.565
+ $X2=4.885 $Y2=1.75
r161 17 19 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.09 $Y=1.565
+ $X2=5.09 $Y2=0.815
r162 13 53 19.9686 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.795 $Y=1.935
+ $X2=4.795 $Y2=1.75
r163 13 15 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.795 $Y=1.935
+ $X2=4.795 $Y2=2.335
r164 4 39 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.985
+ $Y=1.895 $X2=10.125 $Y2=2.04
r165 3 42 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.975 $X2=3.96 $Y2=2.12
r166 2 50 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.355
+ $Y=0.625 $X2=9.48 $Y2=0.835
r167 1 23 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=3.835
+ $Y=0.605 $X2=3.98 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_1075_95# 1 2 9 11 12 15 17 18 21 23 24 27
+ 29 32 34 35 38 41 46 47 50 51 53 55 59 61
c164 46 0 2.75459e-19 $X=7 $Y=1.66
c165 41 0 6.43713e-20 $X=11.895 $Y=1.015
c166 34 0 1.84815e-19 $X=11.895 $Y=3.075
c167 15 0 1.81155e-19 $X=6.005 $Y=2.715
r168 57 61 0.94211 $w=3.3e-07 $l=1.88e-07 $layer=LI1_cond $X=7.28 $Y=0.78
+ $X2=7.092 $Y2=0.78
r169 57 59 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=7.28 $Y=0.78
+ $X2=7.515 $Y2=0.78
r170 53 55 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=7.165 $Y=2.07
+ $X2=7.47 $Y2=2.07
r171 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.115
+ $Y=0.35 $X2=7.115 $Y2=0.35
r172 48 61 5.66538 $w=2.95e-07 $l=1.76125e-07 $layer=LI1_cond $X=7.115 $Y=0.615
+ $X2=7.092 $Y2=0.78
r173 48 50 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=7.115 $Y=0.615
+ $X2=7.115 $Y2=0.35
r174 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7 $Y=1.66
+ $X2=7 $Y2=1.66
r175 44 53 7.03324 $w=1.9e-07 $l=1.71026e-07 $layer=LI1_cond $X=7.035 $Y=1.975
+ $X2=7.165 $Y2=2.07
r176 44 46 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=7.035 $Y=1.975
+ $X2=7.035 $Y2=1.66
r177 43 61 5.66538 $w=2.95e-07 $l=1.9139e-07 $layer=LI1_cond $X=7.035 $Y=0.945
+ $X2=7.092 $Y2=0.78
r178 43 46 31.6922 $w=2.58e-07 $l=7.15e-07 $layer=LI1_cond $X=7.035 $Y=0.945
+ $X2=7.035 $Y2=1.66
r179 39 41 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=11.775 $Y=1.015
+ $X2=11.895 $Y2=1.015
r180 37 51 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=7.115 $Y=0.255
+ $X2=7.115 $Y2=0.35
r181 35 47 46.7153 $w=6.7e-07 $l=5.85e-07 $layer=POLY_cond $X=6.415 $Y=1.83
+ $X2=7 $Y2=1.83
r182 35 36 29.4955 $w=6.7e-07 $l=4.1e-07 $layer=POLY_cond $X=6.415 $Y=1.83
+ $X2=6.005 $Y2=1.83
r183 33 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.895 $Y=1.09
+ $X2=11.895 $Y2=1.015
r184 33 34 1017.84 $w=1.5e-07 $l=1.985e-06 $layer=POLY_cond $X=11.895 $Y=1.09
+ $X2=11.895 $Y2=3.075
r185 32 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.775 $Y=0.94
+ $X2=11.775 $Y2=1.015
r186 31 32 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=11.775 $Y=0.255
+ $X2=11.775 $Y2=0.94
r187 30 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.77 $Y=0.18
+ $X2=9.695 $Y2=0.18
r188 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.7 $Y=0.18
+ $X2=11.775 $Y2=0.255
r189 29 30 989.638 $w=1.5e-07 $l=1.93e-06 $layer=POLY_cond $X=11.7 $Y=0.18
+ $X2=9.77 $Y2=0.18
r190 25 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.695 $Y=0.255
+ $X2=9.695 $Y2=0.18
r191 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.695 $Y=0.255
+ $X2=9.695 $Y2=0.835
r192 23 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.82 $Y=3.15
+ $X2=11.895 $Y2=3.075
r193 23 24 1258.84 $w=1.5e-07 $l=2.455e-06 $layer=POLY_cond $X=11.82 $Y=3.15
+ $X2=9.365 $Y2=3.15
r194 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.29 $Y=3.075
+ $X2=9.365 $Y2=3.15
r195 19 21 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.29 $Y=3.075
+ $X2=9.29 $Y2=2.695
r196 18 37 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.28 $Y=0.18
+ $X2=7.115 $Y2=0.255
r197 17 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.62 $Y=0.18
+ $X2=9.695 $Y2=0.18
r198 17 18 1199.87 $w=1.5e-07 $l=2.34e-06 $layer=POLY_cond $X=9.62 $Y=0.18
+ $X2=7.28 $Y2=0.18
r199 13 36 38.5613 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.005 $Y=2.165
+ $X2=6.005 $Y2=1.83
r200 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.005 $Y=2.165
+ $X2=6.005 $Y2=2.715
r201 11 36 39.618 $w=6.6e-07 $l=2.64858e-07 $layer=POLY_cond $X=5.93 $Y=1.6
+ $X2=6.005 $Y2=1.83
r202 11 12 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=5.93 $Y=1.6
+ $X2=5.525 $Y2=1.6
r203 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.45 $Y=1.525
+ $X2=5.525 $Y2=1.6
r204 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.45 $Y=1.525
+ $X2=5.45 $Y2=0.815
r205 2 55 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.325
+ $Y=1.955 $X2=7.47 $Y2=2.08
r206 1 59 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.39
+ $Y=0.595 $X2=7.515 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_722_23# 1 2 8 10 11 12 13 15 16 17 19 20
+ 22 23 26 27 28 30 33 37 39 40 43 48 49
c131 30 0 1.75353e-19 $X=6.055 $Y=2.12
r132 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.545
+ $Y=0.35 $X2=6.545 $Y2=0.35
r133 41 43 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=6.22 $Y=2.215
+ $X2=6.22 $Y2=2.63
r134 39 48 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.38 $Y=0.345
+ $X2=6.545 $Y2=0.345
r135 39 40 36.0455 $w=1.78e-07 $l=5.85e-07 $layer=LI1_cond $X=6.38 $Y=0.345
+ $X2=5.795 $Y2=0.345
r136 35 40 7.34943 $w=1.8e-07 $l=1.87681e-07 $layer=LI1_cond $X=5.647 $Y=0.435
+ $X2=5.795 $Y2=0.345
r137 35 37 14.845 $w=2.93e-07 $l=3.8e-07 $layer=LI1_cond $X=5.647 $Y=0.435
+ $X2=5.647 $Y2=0.815
r138 33 52 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.555 $Y=2.12
+ $X2=5.415 $Y2=2.12
r139 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.555
+ $Y=2.12 $X2=5.555 $Y2=2.12
r140 30 41 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=6.055 $Y=2.12
+ $X2=6.22 $Y2=2.215
r141 30 32 29.1866 $w=1.88e-07 $l=5e-07 $layer=LI1_cond $X=6.055 $Y=2.12
+ $X2=5.555 $Y2=2.12
r142 29 49 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=6.545 $Y=0.265
+ $X2=6.545 $Y2=0.35
r143 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=2.285
+ $X2=5.415 $Y2=2.12
r144 25 26 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.415 $Y=2.285
+ $X2=5.415 $Y2=3.075
r145 24 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.345 $Y=3.15
+ $X2=4.27 $Y2=3.15
r146 23 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.34 $Y=3.15
+ $X2=5.415 $Y2=3.075
r147 23 24 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=5.34 $Y=3.15
+ $X2=4.345 $Y2=3.15
r148 20 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=3.075
+ $X2=4.27 $Y2=3.15
r149 20 22 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.27 $Y=3.075
+ $X2=4.27 $Y2=2.545
r150 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.195 $Y=1.355
+ $X2=4.195 $Y2=0.925
r151 15 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=3.15
+ $X2=4.27 $Y2=3.15
r152 15 16 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.195 $Y=3.15
+ $X2=3.76 $Y2=3.15
r153 14 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.76 $Y=1.43
+ $X2=3.685 $Y2=1.43
r154 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.12 $Y=1.43
+ $X2=4.195 $Y2=1.355
r155 13 14 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.12 $Y=1.43
+ $X2=3.76 $Y2=1.43
r156 11 29 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.38 $Y=0.19
+ $X2=6.545 $Y2=0.265
r157 11 12 1343.45 $w=1.5e-07 $l=2.62e-06 $layer=POLY_cond $X=6.38 $Y=0.19
+ $X2=3.76 $Y2=0.19
r158 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.685 $Y=3.075
+ $X2=3.76 $Y2=3.15
r159 9 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.685 $Y=1.505
+ $X2=3.685 $Y2=1.43
r160 9 10 805.043 $w=1.5e-07 $l=1.57e-06 $layer=POLY_cond $X=3.685 $Y=1.505
+ $X2=3.685 $Y2=3.075
r161 8 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.685 $Y=1.355
+ $X2=3.685 $Y2=1.43
r162 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.685 $Y=0.265
+ $X2=3.76 $Y2=0.19
r163 7 8 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.685 $Y=0.265
+ $X2=3.685 $Y2=1.355
r164 2 43 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.08
+ $Y=2.505 $X2=6.22 $Y2=2.63
r165 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.525
+ $Y=0.605 $X2=5.665 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_1161_95# 1 2 7 9 10 11 12 14 15 16 17 19
+ 21 23 25 26 30 34 37 38 42 46 47 54 55 58 59
c156 42 0 3.22864e-20 $X=7.57 $Y=1.29
c157 30 0 3.52766e-19 $X=9.91 $Y=2.315
r158 57 59 6.89376 $w=5.48e-07 $l=3.17e-07 $layer=LI1_cond $X=8.485 $Y=1.9
+ $X2=8.802 $Y2=1.9
r159 57 58 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.485 $Y=1.9
+ $X2=8.32 $Y2=1.9
r160 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.82
+ $Y=1.06 $X2=8.82 $Y2=1.06
r161 52 59 6.02202 $w=2.25e-07 $l=2.75e-07 $layer=LI1_cond $X=8.802 $Y=1.625
+ $X2=8.802 $Y2=1.9
r162 52 54 28.9391 $w=2.23e-07 $l=5.65e-07 $layer=LI1_cond $X=8.802 $Y=1.625
+ $X2=8.802 $Y2=1.06
r163 51 54 5.89026 $w=2.23e-07 $l=1.15e-07 $layer=LI1_cond $X=8.802 $Y=0.945
+ $X2=8.802 $Y2=1.06
r164 47 51 7.1387 $w=3.3e-07 $l=2.13787e-07 $layer=LI1_cond $X=8.69 $Y=0.78
+ $X2=8.802 $Y2=0.945
r165 47 49 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=8.69 $Y=0.78
+ $X2=8.375 $Y2=0.78
r166 46 58 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.655 $Y=1.71
+ $X2=8.32 $Y2=1.71
r167 43 63 10.2281 $w=3.77e-07 $l=8e-08 $layer=POLY_cond $X=7.605 $Y=1.29
+ $X2=7.605 $Y2=1.21
r168 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.57
+ $Y=1.29 $X2=7.57 $Y2=1.29
r169 40 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.53 $Y=1.625
+ $X2=7.655 $Y2=1.71
r170 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.53 $Y=1.625
+ $X2=7.53 $Y2=1.29
r171 38 39 55.7151 $w=1.86e-07 $l=2.15e-07 $layer=POLY_cond $X=9.91 $Y=1.445
+ $X2=10.125 $Y2=1.445
r172 36 55 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.82 $Y=1.415
+ $X2=8.82 $Y2=1.06
r173 36 37 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=8.82 $Y=1.415
+ $X2=8.82 $Y2=1.49
r174 32 39 7.89931 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=10.125 $Y=1.325
+ $X2=10.125 $Y2=1.445
r175 32 34 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=10.125 $Y=1.325
+ $X2=10.125 $Y2=0.835
r176 28 38 7.89931 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=9.91 $Y=1.565
+ $X2=9.91 $Y2=1.445
r177 28 30 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=9.91 $Y=1.565
+ $X2=9.91 $Y2=2.315
r178 27 37 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.985 $Y=1.49
+ $X2=8.82 $Y2=1.49
r179 26 38 21.3816 $w=1.86e-07 $l=9.48683e-08 $layer=POLY_cond $X=9.835 $Y=1.49
+ $X2=9.91 $Y2=1.445
r180 26 27 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=9.835 $Y=1.49
+ $X2=8.985 $Y2=1.49
r181 24 37 13.5877 $w=2.4e-07 $l=9.28709e-08 $layer=POLY_cond $X=8.78 $Y=1.565
+ $X2=8.82 $Y2=1.49
r182 24 25 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=8.78 $Y=1.565
+ $X2=8.78 $Y2=3.035
r183 21 63 28.9397 $w=3.77e-07 $l=1.62019e-07 $layer=POLY_cond $X=7.73 $Y=1.125
+ $X2=7.605 $Y2=1.21
r184 21 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.73 $Y=1.125
+ $X2=7.73 $Y2=0.805
r185 17 43 82.6373 $w=3.77e-07 $l=5.4353e-07 $layer=POLY_cond $X=7.685 $Y=1.795
+ $X2=7.605 $Y2=1.29
r186 17 19 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.685 $Y=1.795
+ $X2=7.685 $Y2=2.275
r187 15 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.705 $Y=3.11
+ $X2=8.78 $Y2=3.035
r188 15 16 1125.52 $w=1.5e-07 $l=2.195e-06 $layer=POLY_cond $X=8.705 $Y=3.11
+ $X2=6.51 $Y2=3.11
r189 12 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.435 $Y=3.035
+ $X2=6.51 $Y2=3.11
r190 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.435 $Y=3.035
+ $X2=6.435 $Y2=2.715
r191 10 63 24.4204 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.405 $Y=1.21
+ $X2=7.605 $Y2=1.21
r192 10 11 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=7.405 $Y=1.21
+ $X2=5.955 $Y2=1.21
r193 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.88 $Y=1.135
+ $X2=5.955 $Y2=1.21
r194 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.88 $Y=1.135
+ $X2=5.88 $Y2=0.815
r195 2 57 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.345
+ $Y=1.955 $X2=8.485 $Y2=2.08
r196 1 49 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=8.235
+ $Y=0.595 $X2=8.375 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%CLK 3 6 8 9 13 15
c37 13 0 3.22864e-20 $X=8.25 $Y=1.295
c38 9 0 1.33087e-19 $X=8.4 $Y=1.295
r39 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.25 $Y=1.295
+ $X2=8.25 $Y2=1.46
r40 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.25 $Y=1.295
+ $X2=8.25 $Y2=1.13
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.25
+ $Y=1.295 $X2=8.25 $Y2=1.295
r42 9 14 5.16019 $w=3.33e-07 $l=1.5e-07 $layer=LI1_cond $X=8.4 $Y=1.287 $X2=8.25
+ $Y2=1.287
r43 8 14 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=7.92 $Y=1.287
+ $X2=8.25 $Y2=1.287
r44 6 16 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=8.27 $Y=2.275
+ $X2=8.27 $Y2=1.46
r45 3 15 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=8.16 $Y=0.805
+ $X2=8.16 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_2082_99# 1 2 9 11 13 16 19 21 25 27 31 34
+ 35 36 37 38 40 41 44 48 49 53 55 59
c125 55 0 9.69379e-20 $X=10.74 $Y=1.88
c126 53 0 1.10201e-19 $X=10.575 $Y=1.88
c127 41 0 1.73242e-19 $X=11.645 $Y=1.805
c128 9 0 1.05913e-19 $X=10.485 $Y=0.835
r129 53 61 14.7551 $w=2.94e-07 $l=9e-08 $layer=POLY_cond $X=10.575 $Y=1.905
+ $X2=10.485 $Y2=1.905
r130 52 55 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=10.575 $Y=1.88
+ $X2=10.74 $Y2=1.88
r131 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.575
+ $Y=1.88 $X2=10.575 $Y2=1.88
r132 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.375
+ $Y=1.14 $X2=12.375 $Y2=1.14
r133 46 57 14.878 $w=4.51e-07 $l=6.84945e-07 $layer=LI1_cond $X=11.785 $Y=1.31
+ $X2=11.482 $Y2=0.76
r134 46 48 10.5326 $w=6.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.785 $Y=1.31
+ $X2=12.375 $Y2=1.31
r135 42 59 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.645 $Y=1.975
+ $X2=11.645 $Y2=1.89
r136 42 44 2.67531 $w=2.78e-07 $l=6.5e-08 $layer=LI1_cond $X=11.645 $Y=1.975
+ $X2=11.645 $Y2=2.04
r137 41 59 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.645 $Y=1.805
+ $X2=11.645 $Y2=1.89
r138 40 46 10.8055 $w=4.51e-07 $l=3.98905e-07 $layer=LI1_cond $X=11.645 $Y=1.645
+ $X2=11.785 $Y2=1.31
r139 40 41 6.58539 $w=2.78e-07 $l=1.6e-07 $layer=LI1_cond $X=11.645 $Y=1.645
+ $X2=11.645 $Y2=1.805
r140 38 59 3.18746 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=11.505 $Y=1.89
+ $X2=11.645 $Y2=1.89
r141 38 55 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=11.505 $Y=1.89
+ $X2=10.74 $Y2=1.89
r142 35 49 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=12.375 $Y=1.495
+ $X2=12.375 $Y2=1.14
r143 35 36 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=12.375 $Y=1.495
+ $X2=12.375 $Y2=1.57
r144 34 49 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.375 $Y=0.975
+ $X2=12.375 $Y2=1.14
r145 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=13.31 $Y=1.495
+ $X2=13.31 $Y2=0.815
r146 28 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.985 $Y=1.57
+ $X2=12.91 $Y2=1.57
r147 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.235 $Y=1.57
+ $X2=13.31 $Y2=1.495
r148 27 28 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=13.235 $Y=1.57
+ $X2=12.985 $Y2=1.57
r149 23 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.91 $Y=1.645
+ $X2=12.91 $Y2=1.57
r150 23 25 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=12.91 $Y=1.645
+ $X2=12.91 $Y2=2.465
r151 22 36 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.54 $Y=1.57
+ $X2=12.375 $Y2=1.57
r152 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.835 $Y=1.57
+ $X2=12.91 $Y2=1.57
r153 21 22 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=12.835 $Y=1.57
+ $X2=12.54 $Y2=1.57
r154 17 36 13.5877 $w=2.4e-07 $l=7.98436e-08 $layer=POLY_cond $X=12.385 $Y=1.645
+ $X2=12.375 $Y2=1.57
r155 17 19 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=12.385 $Y=1.645
+ $X2=12.385 $Y2=2.155
r156 16 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.36 $Y=0.655
+ $X2=12.36 $Y2=0.975
r157 11 53 46.7245 $w=2.94e-07 $l=3.67933e-07 $layer=POLY_cond $X=10.86 $Y=2.095
+ $X2=10.575 $Y2=1.905
r158 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.86 $Y=2.095
+ $X2=10.86 $Y2=2.415
r159 7 61 18.4939 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.485 $Y=1.715
+ $X2=10.485 $Y2=1.905
r160 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=10.485 $Y=1.715
+ $X2=10.485 $Y2=0.835
r161 2 44 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=11.46
+ $Y=1.895 $X2=11.62 $Y2=2.04
r162 1 57 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=11.155
+ $Y=0.625 $X2=11.295 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_1873_497# 1 2 7 9 12 16 20 24 26 28 33
c61 26 0 2.3558e-19 $X=11.17 $Y=1.54
c62 16 0 1.10201e-19 $X=9.695 $Y=2.05
c63 12 0 9.69379e-20 $X=11.385 $Y=2.315
r64 27 33 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.17 $Y=1.54
+ $X2=11.385 $Y2=1.54
r65 27 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.17 $Y=1.54
+ $X2=11.08 $Y2=1.54
r66 26 28 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=11.17 $Y=1.54
+ $X2=11.005 $Y2=1.54
r67 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.17
+ $Y=1.54 $X2=11.17 $Y2=1.54
r68 23 24 3.80956 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=10.075 $Y=1.53
+ $X2=9.802 $Y2=1.53
r69 23 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=10.075 $Y=1.53
+ $X2=11.005 $Y2=1.53
r70 18 24 2.88756 $w=3.3e-07 $l=1.44375e-07 $layer=LI1_cond $X=9.91 $Y=1.445
+ $X2=9.802 $Y2=1.53
r71 18 20 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=9.91 $Y=1.445
+ $X2=9.91 $Y2=0.9
r72 14 24 2.88756 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=9.695 $Y=1.615
+ $X2=9.802 $Y2=1.53
r73 14 16 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=9.695 $Y=1.615
+ $X2=9.695 $Y2=2.05
r74 10 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.385 $Y=1.705
+ $X2=11.385 $Y2=1.54
r75 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=11.385 $Y=1.705
+ $X2=11.385 $Y2=2.315
r76 7 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.08 $Y=1.375
+ $X2=11.08 $Y2=1.54
r77 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.08 $Y=1.375
+ $X2=11.08 $Y2=0.945
r78 2 16 600 $w=1.7e-07 $l=5.76867e-07 $layer=licon1_PDIFF $count=1 $X=9.365
+ $Y=2.485 $X2=9.695 $Y2=2.05
r79 1 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.77
+ $Y=0.625 $X2=9.91 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_2409_367# 1 2 9 12 15 16 20 21 27 31 34
c65 15 0 5.51483e-20 $X=12.725 $Y=1.815
r66 29 31 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=12.575 $Y=0.64
+ $X2=12.725 $Y2=0.64
r67 26 27 9.26921 $w=6.78e-07 $l=8.5e-08 $layer=LI1_cond $X=12.725 $Y=2.155
+ $X2=12.81 $Y2=2.155
r68 24 26 9.76211 $w=6.78e-07 $l=5.55e-07 $layer=LI1_cond $X=12.17 $Y=2.155
+ $X2=12.725 $Y2=2.155
r69 21 35 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=13.812 $Y=1.51
+ $X2=13.812 $Y2=1.675
r70 21 34 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=13.812 $Y=1.51
+ $X2=13.812 $Y2=1.345
r71 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.79
+ $Y=1.51 $X2=13.79 $Y2=1.51
r72 18 20 37.5696 $w=2.48e-07 $l=8.15e-07 $layer=LI1_cond $X=13.75 $Y=2.325
+ $X2=13.75 $Y2=1.51
r73 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.625 $Y=2.41
+ $X2=13.75 $Y2=2.325
r74 16 27 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=13.625 $Y=2.41
+ $X2=12.81 $Y2=2.41
r75 15 26 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=12.725 $Y=1.815
+ $X2=12.725 $Y2=2.155
r76 14 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.725 $Y=0.805
+ $X2=12.725 $Y2=0.64
r77 14 15 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=12.725 $Y=0.805
+ $X2=12.725 $Y2=1.815
r78 12 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=13.925 $Y=2.465
+ $X2=13.925 $Y2=1.675
r79 9 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.755 $Y=0.815
+ $X2=13.755 $Y2=1.345
r80 2 24 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.045
+ $Y=1.835 $X2=12.17 $Y2=1.98
r81 1 29 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=12.435
+ $Y=0.445 $X2=12.575 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_27_483# 1 2 9 11 12 13
c28 11 0 1.7997e-19 $X=1.745 $Y=2.375
r29 13 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.91 $Y=2.375
+ $X2=1.91 $Y2=2.56
r30 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=2.375
+ $X2=1.91 $Y2=2.375
r31 11 12 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.745 $Y=2.375
+ $X2=0.355 $Y2=2.375
r32 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=2.46
+ $X2=0.355 $Y2=2.375
r33 7 9 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=0.225 $Y=2.46 $X2=0.225
+ $Y2=2.56
r34 2 16 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=2.415 $X2=1.91 $Y2=2.56
r35 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.415 $X2=0.26 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48 51
+ 52 53 55 67 71 79 87 92 99 100 103 106 109 112 115 118
r135 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r136 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r137 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r138 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r139 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r141 100 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r142 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r143 97 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=13.71 $Y2=3.33
r144 97 99 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=14.16 $Y2=3.33
r145 96 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r146 96 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r147 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r148 93 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.86 $Y=3.33
+ $X2=12.695 $Y2=3.33
r149 93 95 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=12.86 $Y=3.33
+ $X2=13.2 $Y2=3.33
r150 92 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.71 $Y2=3.33
r151 92 95 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.2 $Y2=3.33
r152 91 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r153 91 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r154 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r155 88 112 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=11.335 $Y=3.33
+ $X2=11.157 $Y2=3.33
r156 88 90 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=11.335 $Y=3.33
+ $X2=12.24 $Y2=3.33
r157 87 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.53 $Y=3.33
+ $X2=12.695 $Y2=3.33
r158 87 90 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=12.53 $Y=3.33
+ $X2=12.24 $Y2=3.33
r159 86 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r160 85 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r161 83 86 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r162 83 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r163 82 85 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r164 82 83 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r165 80 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.16 $Y=3.33
+ $X2=7.995 $Y2=3.33
r166 80 82 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.16 $Y=3.33
+ $X2=8.4 $Y2=3.33
r167 79 112 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=10.98 $Y=3.33
+ $X2=11.157 $Y2=3.33
r168 79 85 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.98 $Y=3.33
+ $X2=10.8 $Y2=3.33
r169 78 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r170 77 78 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r171 75 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r172 74 77 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r173 74 75 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r174 72 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=4.485 $Y2=3.33
r175 72 74 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=5.04 $Y2=3.33
r176 71 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.83 $Y=3.33
+ $X2=7.995 $Y2=3.33
r177 71 77 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.83 $Y=3.33
+ $X2=7.44 $Y2=3.33
r178 70 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r179 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r180 67 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.485 $Y2=3.33
r181 67 69 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r182 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r183 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r184 63 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r185 63 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r186 62 65 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r187 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r188 60 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r189 60 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r190 58 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r191 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r192 55 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r193 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r194 53 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r195 53 75 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r196 51 65 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.12 $Y2=3.33
r197 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.445 $Y2=3.33
r198 50 69 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=4.08 $Y2=3.33
r199 50 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=3.445 $Y2=3.33
r200 46 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=3.33
r201 46 48 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=2.77
r202 42 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.695 $Y=3.245
+ $X2=12.695 $Y2=3.33
r203 42 44 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=12.695 $Y=3.245
+ $X2=12.695 $Y2=2.77
r204 38 112 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.157 $Y=3.245
+ $X2=11.157 $Y2=3.33
r205 38 40 32.9501 $w=3.53e-07 $l=1.015e-06 $layer=LI1_cond $X=11.157 $Y=3.245
+ $X2=11.157 $Y2=2.23
r206 34 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.995 $Y=3.245
+ $X2=7.995 $Y2=3.33
r207 34 36 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.995 $Y=3.245
+ $X2=7.995 $Y2=2.78
r208 30 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=3.33
r209 30 32 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=2.82
r210 26 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=3.245
+ $X2=3.445 $Y2=3.33
r211 26 28 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=3.445 $Y=3.245
+ $X2=3.445 $Y2=2.89
r212 22 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r213 22 24 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.755
r214 7 48 600 $w=1.7e-07 $l=9.9554e-07 $layer=licon1_PDIFF $count=1 $X=13.585
+ $Y=1.835 $X2=13.71 $Y2=2.77
r215 6 44 600 $w=1.7e-07 $l=1.04592e-06 $layer=licon1_PDIFF $count=1 $X=12.46
+ $Y=1.835 $X2=12.695 $Y2=2.77
r216 5 40 300 $w=1.7e-07 $l=2.47184e-07 $layer=licon1_PDIFF $count=2 $X=10.935
+ $Y=2.205 $X2=11.17 $Y2=2.23
r217 4 36 600 $w=1.7e-07 $l=9.35147e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.955 $X2=7.995 $Y2=2.78
r218 3 32 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=2.125 $X2=4.485 $Y2=2.82
r219 2 28 600 $w=1.7e-07 $l=5.57136e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=2.405 $X2=3.41 $Y2=2.89
r220 1 24 600 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.415 $X2=0.69 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_196_119# 1 2 3 4 15 17 21 22 23 26 27 30
+ 32 33 34 35 38 39 40 42 43 44 47 49 53 54 55
c170 54 0 1.8781e-19 $X=3.06 $Y=2.47
r171 55 58 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.71 $Y=2.47
+ $X2=5.71 $Y2=2.63
r172 45 47 25.5009 $w=2.33e-07 $l=5.2e-07 $layer=LI1_cond $X=6.082 $Y=1.335
+ $X2=6.082 $Y2=0.815
r173 43 45 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=5.965 $Y=1.42
+ $X2=6.082 $Y2=1.335
r174 43 44 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=5.965 $Y=1.42
+ $X2=4.405 $Y2=1.42
r175 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.32 $Y=1.335
+ $X2=4.405 $Y2=1.42
r176 41 42 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=4.32 $Y=0.435
+ $X2=4.32 $Y2=1.335
r177 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.235 $Y=0.35
+ $X2=4.32 $Y2=0.435
r178 39 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.235 $Y=0.35
+ $X2=3.555 $Y2=0.35
r179 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=0.435
+ $X2=3.555 $Y2=0.35
r180 37 38 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=3.47 $Y=0.435
+ $X2=3.47 $Y2=1.56
r181 36 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=2.47
+ $X2=3.06 $Y2=2.47
r182 35 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.545 $Y=2.47
+ $X2=5.71 $Y2=2.47
r183 35 36 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.545 $Y=2.47
+ $X2=3.145 $Y2=2.47
r184 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.385 $Y=1.645
+ $X2=3.47 $Y2=1.56
r185 33 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.385 $Y=1.645
+ $X2=3.145 $Y2=1.645
r186 31 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=2.555
+ $X2=3.06 $Y2=2.47
r187 31 32 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.06 $Y=2.555
+ $X2=3.06 $Y2=2.895
r188 30 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=2.385
+ $X2=3.06 $Y2=2.47
r189 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=1.73
+ $X2=3.145 $Y2=1.645
r190 29 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.06 $Y=1.73
+ $X2=3.06 $Y2=2.385
r191 28 53 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=2.425 $Y=2.98
+ $X2=2.34 $Y2=2.95
r192 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.975 $Y=2.98
+ $X2=3.06 $Y2=2.895
r193 27 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.975 $Y=2.98
+ $X2=2.425 $Y2=2.98
r194 26 53 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.34 $Y=2.835
+ $X2=2.34 $Y2=2.95
r195 25 26 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=2.34 $Y=1.415
+ $X2=2.34 $Y2=2.835
r196 24 49 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.785 $Y=1.31
+ $X2=1.785 $Y2=1.09
r197 23 25 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.255 $Y=1.31
+ $X2=2.34 $Y2=1.415
r198 23 24 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=2.255 $Y=1.31
+ $X2=1.87 $Y2=1.31
r199 21 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=1.09
+ $X2=1.785 $Y2=1.09
r200 21 22 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.7 $Y=1.09
+ $X2=1.34 $Y2=1.09
r201 17 53 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=2.95 $X2=2.34
+ $Y2=2.95
r202 17 19 38.8323 $w=2.28e-07 $l=7.75e-07 $layer=LI1_cond $X=2.255 $Y=2.95
+ $X2=1.48 $Y2=2.95
r203 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.175 $Y=1.005
+ $X2=1.34 $Y2=1.09
r204 13 15 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.175 $Y=1.005
+ $X2=1.175 $Y2=0.805
r205 4 58 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.505 $X2=5.71 $Y2=2.63
r206 3 19 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.415 $X2=1.48 $Y2=2.93
r207 2 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.955
+ $Y=0.605 $X2=6.095 $Y2=0.815
r208 1 15 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.595 $X2=1.175 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_974_425# 1 2 7 10 15
c34 15 0 7.42513e-21 $X=6.73 $Y=2.78
r35 15 17 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6.73 $Y=2.78 $X2=6.73
+ $Y2=2.98
r36 10 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.105 $Y=2.82
+ $X2=5.105 $Y2=2.98
r37 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=2.98
+ $X2=5.105 $Y2=2.98
r38 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.565 $Y=2.98
+ $X2=6.73 $Y2=2.98
r39 7 8 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=6.565 $Y=2.98
+ $X2=5.27 $Y2=2.98
r40 2 15 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=6.51
+ $Y=2.505 $X2=6.73 $Y2=2.78
r41 1 10 600 $w=1.7e-07 $l=8.03959e-07 $layer=licon1_PDIFF $count=1 $X=4.87
+ $Y=2.125 $X2=5.105 $Y2=2.82
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%A_1786_497# 1 2 7 11 16
c31 16 0 1.73489e-19 $X=9.24 $Y=2.815
r32 14 16 7.61969 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=2.815
+ $X2=9.24 $Y2=2.815
r33 9 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=10.645 $Y=2.725
+ $X2=10.645 $Y2=2.41
r34 7 9 7.17723 $w=2.2e-07 $l=2.13014e-07 $layer=LI1_cond $X=10.48 $Y=2.835
+ $X2=10.645 $Y2=2.725
r35 7 16 64.9559 $w=2.18e-07 $l=1.24e-06 $layer=LI1_cond $X=10.48 $Y=2.835
+ $X2=9.24 $Y2=2.835
r36 2 11 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=10.52
+ $Y=2.205 $X2=10.645 $Y2=2.41
r37 1 14 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=8.93
+ $Y=2.485 $X2=9.075 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%Q 1 2 7 8 9 10 11 20 28
r23 28 37 1.95329 $w=2.93e-07 $l=5e-08 $layer=LI1_cond $X=13.137 $Y=1.295
+ $X2=13.137 $Y2=1.345
r24 10 11 8.74746 $w=4.13e-07 $l=3.15e-07 $layer=LI1_cond $X=13.197 $Y=1.665
+ $X2=13.197 $Y2=1.98
r25 10 29 3.13798 $w=4.13e-07 $l=1.13e-07 $layer=LI1_cond $X=13.197 $Y=1.665
+ $X2=13.197 $Y2=1.552
r26 9 29 5.27625 $w=4.13e-07 $l=1.9e-07 $layer=LI1_cond $X=13.197 $Y=1.362
+ $X2=13.197 $Y2=1.552
r27 9 37 1.45179 $w=4.13e-07 $l=1.7e-08 $layer=LI1_cond $X=13.197 $Y=1.362
+ $X2=13.197 $Y2=1.345
r28 9 28 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=13.137 $Y=1.277
+ $X2=13.137 $Y2=1.295
r29 8 9 13.7512 $w=2.93e-07 $l=3.52e-07 $layer=LI1_cond $X=13.137 $Y=0.925
+ $X2=13.137 $Y2=1.277
r30 7 8 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=13.137 $Y=0.555
+ $X2=13.137 $Y2=0.925
r31 7 20 0.585988 $w=2.93e-07 $l=1.5e-08 $layer=LI1_cond $X=13.137 $Y=0.555
+ $X2=13.137 $Y2=0.54
r32 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.985
+ $Y=1.835 $X2=13.125 $Y2=1.98
r33 1 20 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=12.97
+ $Y=0.395 $X2=13.095 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%Q_N 1 2 7 8 9 10 11 12 13 24 30
r15 22 30 0.381727 $w=4.68e-07 $l=1.5e-08 $layer=LI1_cond $X=14.08 $Y=0.94
+ $X2=14.08 $Y2=0.925
r16 13 44 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=14.18 $Y=2.775
+ $X2=14.18 $Y2=2.91
r17 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=14.18 $Y=2.405
+ $X2=14.18 $Y2=2.775
r18 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=14.18 $Y=1.98
+ $X2=14.18 $Y2=2.405
r19 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=14.18 $Y=1.665
+ $X2=14.18 $Y2=1.98
r20 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=14.18 $Y=1.295
+ $X2=14.18 $Y2=1.665
r21 9 47 5.12197 $w=2.68e-07 $l=1.2e-07 $layer=LI1_cond $X=14.18 $Y=1.295
+ $X2=14.18 $Y2=1.175
r22 8 47 7.23736 $w=4.68e-07 $l=2e-07 $layer=LI1_cond $X=14.08 $Y=0.975
+ $X2=14.08 $Y2=1.175
r23 8 22 0.890697 $w=4.68e-07 $l=3.5e-08 $layer=LI1_cond $X=14.08 $Y=0.975
+ $X2=14.08 $Y2=0.94
r24 8 30 0.890697 $w=4.68e-07 $l=3.5e-08 $layer=LI1_cond $X=14.08 $Y=0.89
+ $X2=14.08 $Y2=0.925
r25 7 8 8.52524 $w=4.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.08 $Y=0.555
+ $X2=14.08 $Y2=0.89
r26 7 24 0.381727 $w=4.68e-07 $l=1.5e-08 $layer=LI1_cond $X=14.08 $Y=0.555
+ $X2=14.08 $Y2=0.54
r27 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14
+ $Y=1.835 $X2=14.14 $Y2=2.91
r28 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14
+ $Y=1.835 $X2=14.14 $Y2=1.98
r29 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.83
+ $Y=0.395 $X2=13.97 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_1%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48
+ 51 52 54 55 56 58 70 77 85 95 96 102 105 108 111
c134 40 0 6.43713e-20 $X=10.845 $Y=0.77
c135 36 0 1.42371e-19 $X=7.945 $Y=0.785
r136 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r137 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r138 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r139 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r140 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r141 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r142 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r143 93 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.24 $Y2=0
r144 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r145 90 111 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.27 $Y=0
+ $X2=12.125 $Y2=0
r146 90 92 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=12.27 $Y=0 $X2=13.2
+ $Y2=0
r147 89 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r148 89 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r149 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r150 86 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.01 $Y=0
+ $X2=10.845 $Y2=0
r151 86 88 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=11.01 $Y=0
+ $X2=11.76 $Y2=0
r152 85 111 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.98 $Y=0
+ $X2=12.125 $Y2=0
r153 85 88 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=11.98 $Y=0
+ $X2=11.76 $Y2=0
r154 84 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r155 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r156 81 84 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r157 81 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r158 80 83 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.32
+ $Y2=0
r159 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r160 78 105 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=8.08 $Y=0
+ $X2=7.942 $Y2=0
r161 78 80 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.08 $Y=0 $X2=8.4
+ $Y2=0
r162 77 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.68 $Y=0
+ $X2=10.845 $Y2=0
r163 77 83 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=10.68 $Y=0
+ $X2=10.32 $Y2=0
r164 76 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r165 75 76 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r166 72 75 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.44
+ $Y2=0
r167 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r168 70 105 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.942 $Y2=0
r169 70 75 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.44 $Y2=0
r170 69 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r171 69 103 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=2.16 $Y2=0
r172 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r173 66 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.02 $Y2=0
r174 66 68 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=4.56 $Y2=0
r175 65 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r176 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r177 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r178 62 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r179 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r180 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r181 59 99 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=0
+ $X2=0.247 $Y2=0
r182 59 61 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.495 $Y=0
+ $X2=0.72 $Y2=0
r183 58 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=2.02 $Y2=0
r184 58 64 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.68 $Y2=0
r185 56 76 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=7.44
+ $Y2=0
r186 56 73 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=5.04
+ $Y2=0
r187 54 92 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.2 $Y2=0
r188 54 55 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.565 $Y2=0
r189 53 95 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=13.675 $Y=0
+ $X2=14.16 $Y2=0
r190 53 55 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=13.675 $Y=0
+ $X2=13.565 $Y2=0
r191 51 68 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.575 $Y=0 $X2=4.56
+ $Y2=0
r192 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.575 $Y=0 $X2=4.74
+ $Y2=0
r193 50 72 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.905 $Y=0
+ $X2=5.04 $Y2=0
r194 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=0 $X2=4.74
+ $Y2=0
r195 46 55 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=13.565 $Y=0.085
+ $X2=13.565 $Y2=0
r196 46 48 23.8346 $w=2.18e-07 $l=4.55e-07 $layer=LI1_cond $X=13.565 $Y=0.085
+ $X2=13.565 $Y2=0.54
r197 42 111 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.125 $Y=0.085
+ $X2=12.125 $Y2=0
r198 42 44 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=12.125 $Y=0.085
+ $X2=12.125 $Y2=0.64
r199 38 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.845 $Y=0.085
+ $X2=10.845 $Y2=0
r200 38 40 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=10.845 $Y=0.085
+ $X2=10.845 $Y2=0.77
r201 34 105 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.942 $Y=0.085
+ $X2=7.942 $Y2=0
r202 34 36 29.3349 $w=2.73e-07 $l=7e-07 $layer=LI1_cond $X=7.942 $Y=0.085
+ $X2=7.942 $Y2=0.785
r203 30 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=0.085
+ $X2=4.74 $Y2=0
r204 30 32 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=4.74 $Y=0.085
+ $X2=4.74 $Y2=0.73
r205 26 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r206 26 28 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.73
r207 22 99 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.247 $Y2=0
r208 22 24 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.33 $Y2=0.805
r209 7 48 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=13.385
+ $Y=0.395 $X2=13.54 $Y2=0.54
r210 6 44 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=12.02
+ $Y=0.445 $X2=12.145 $Y2=0.64
r211 5 40 91 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=2 $X=10.56
+ $Y=0.625 $X2=10.845 $Y2=0.77
r212 4 36 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=7.805
+ $Y=0.595 $X2=7.945 $Y2=0.785
r213 3 32 91 $w=1.7e-07 $l=5.28819e-07 $layer=licon1_NDIFF $count=2 $X=4.27
+ $Y=0.605 $X2=4.74 $Y2=0.73
r214 2 28 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.595 $X2=2.02 $Y2=0.73
r215 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.595 $X2=0.33 $Y2=0.805
.ends

