* File: sky130_fd_sc_lp__dfxbp_2.spice
* Created: Fri Aug 28 10:23:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfxbp_2.pex.spice"
.subckt sky130_fd_sc_lp__dfxbp_2  VNB VPB CLK D VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1008 N_A_110_70#_M1008_d N_CLK_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_110_70#_M1028_g N_A_236_463#_M1028_s VNB NSHORT L=0.15
+ W=0.42 AD=0.06825 AS=0.1113 PD=0.745 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75005.2 A=0.063 P=1.14 MULT=1
MM1024 N_A_429_119#_M1024_d N_D_M1024_g N_VGND_M1028_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.06825 PD=0.81 PS=0.745 NRD=17.136 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_537_119#_M1001_d N_A_110_70#_M1001_g N_A_429_119#_M1024_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.06405 AS=0.0819 PD=0.725 PS=0.81 NRD=7.14 NRS=14.28 M=1
+ R=2.8 SA=75001.2 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1000 A_628_119# N_A_236_463#_M1000_g N_A_537_119#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.06405 PD=0.63 PS=0.725 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_670_93#_M1006_g A_628_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.168198 AS=0.0441 PD=1.16491 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1022 N_A_670_93#_M1022_d N_A_537_119#_M1022_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.64 AD=0.130294 AS=0.256302 PD=1.22566 PS=1.77509 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1025 N_A_982_369#_M1025_d N_A_236_463#_M1025_g N_A_670_93#_M1022_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0987 AS=0.0855057 PD=0.89 PS=0.80434 NRD=27.132 NRS=27.852
+ M=1 R=2.8 SA=75003.5 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1026 A_1125_119# N_A_110_70#_M1026_g N_A_982_369#_M1025_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0462 AS=0.0987 PD=0.64 PS=0.89 NRD=15.708 NRS=27.132 M=1 R=2.8
+ SA=75004.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_1169_93#_M1004_g A_1125_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.119938 AS=0.0462 PD=0.935094 PS=0.64 NRD=37.848 NRS=15.708 M=1 R=2.8
+ SA=75004.5 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1005 N_A_1169_93#_M1005_d N_A_982_369#_M1005_g N_VGND_M1004_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.182762 PD=1.81 PS=1.42491 NRD=0 NRS=24.372 M=1
+ R=4.26667 SA=75003.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_A_1169_93#_M1018_g N_A_1513_137#_M1018_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.138733 AS=0.1197 PD=0.976667 PS=1.41 NRD=78.66 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1020 N_Q_N_M1020_d N_A_1513_137#_M1020_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.277467 PD=1.12 PS=1.95333 NRD=0 NRS=17.136 M=1 R=5.6
+ SA=75000.6 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1029 N_Q_N_M1020_d N_A_1513_137#_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75001 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1013 N_Q_M1013_d N_A_1169_93#_M1013_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6 SA=75001.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_Q_M1013_d N_A_1169_93#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1002 N_A_110_70#_M1002_d N_CLK_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VPWR_M1015_d N_A_110_70#_M1015_g N_A_236_463#_M1015_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.177328 AS=0.1696 PD=1.43698 PS=1.81 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1027 N_A_429_119#_M1027_d N_D_M1027_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.116372 PD=0.7 PS=0.943019 NRD=0 NRS=104.154 M=1 R=2.8
+ SA=75000.9 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_537_119#_M1016_d N_A_236_463#_M1016_g N_A_429_119#_M1027_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1212 AS=0.0588 PD=1.07 PS=0.7 NRD=44.5417 NRS=0 M=1
+ R=2.8 SA=75001.3 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1017 A_669_499# N_A_110_70#_M1017_g N_A_537_119#_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0882 AS=0.1212 PD=0.96 PS=1.07 NRD=72.693 NRS=46.886 M=1 R=2.8
+ SA=75001.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_670_93#_M1007_g A_669_499# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.128233 AS=0.0882 PD=0.95 PS=0.96 NRD=56.2829 NRS=72.693 M=1 R=2.8
+ SA=75001.5 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_670_93#_M1009_d N_A_537_119#_M1009_g N_VPWR_M1007_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.256467 PD=1.12 PS=1.9 NRD=0 NRS=19.9167 M=1 R=5.6
+ SA=75001 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1023 N_A_982_369#_M1023_d N_A_110_70#_M1023_g N_A_670_93#_M1009_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.3752 AS=0.1176 PD=2.08667 PS=1.12 NRD=82.0702 NRS=0 M=1
+ R=5.6 SA=75001.5 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1019 A_1157_453# N_A_236_463#_M1019_g N_A_982_369#_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0763 AS=0.1876 PD=0.79 PS=1.04333 NRD=59.3955 NRS=44.5417 M=1
+ R=2.8 SA=75003.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_1169_93#_M1010_g A_1157_453# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0959 AS=0.0763 PD=0.84 PS=0.79 NRD=0 NRS=59.3955 M=1 R=2.8 SA=75003.5
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1030 N_A_1169_93#_M1030_d N_A_982_369#_M1030_g N_VPWR_M1010_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1918 PD=2.21 PS=1.68 NRD=0 NRS=16.4101 M=1 R=5.6
+ SA=75002.1 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_VPWR_M1021_d N_A_1169_93#_M1021_g N_A_1513_137#_M1021_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.17472 AS=0.1696 PD=1.19579 PS=1.81 NRD=36.9178 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1021_d N_A_1513_137#_M1011_g N_Q_N_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.34398 AS=0.1764 PD=2.35421 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1031 N_VPWR_M1031_d N_A_1513_137#_M1031_g N_Q_N_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.27405 AS=0.1764 PD=1.695 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75001 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1003 N_Q_M1003_d N_A_1169_93#_M1003_g N_VPWR_M1031_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.27405 PD=1.54 PS=1.695 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75001.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1012 N_Q_M1003_d N_A_1169_93#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.4031 P=25.61
c_106 VNB 0 1.27355e-19 $X=0 $Y=0
c_1163 A_669_499# 0 1.82964e-19 $X=3.345 $Y=2.495
*
.include "sky130_fd_sc_lp__dfxbp_2.pxi.spice"
*
.ends
*
*
