* File: sky130_fd_sc_lp__clkbuf_1.pex.spice
* Created: Wed Sep  2 09:38:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUF_1%A_69_161# 1 2 9 13 15 18 22 26 31 32 33
r52 31 32 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=2.085
+ $X2=1.175 $Y2=1.92
r53 28 33 6.67463 $w=2.4e-07 $l=1.96914e-07 $layer=LI1_cond $X=1.27 $Y=1.135
+ $X2=1.2 $Y2=0.97
r54 28 32 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.27 $Y=1.135
+ $X2=1.27 $Y2=1.92
r55 24 33 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=0.805 $X2=1.2
+ $Y2=0.97
r56 24 26 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.2 $Y=0.805 $X2=1.2
+ $Y2=0.465
r57 20 31 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.175 $Y=2.1
+ $X2=1.175 $Y2=2.085
r58 20 22 25.7699 $w=3.58e-07 $l=8.05e-07 $layer=LI1_cond $X=1.175 $Y=2.1
+ $X2=1.175 $Y2=2.905
r59 18 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.97
+ $X2=0.51 $Y2=1.135
r60 18 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.97
+ $X2=0.51 $Y2=0.805
r61 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=0.97 $X2=0.51 $Y2=0.97
r62 15 33 0.225187 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=0.97
+ $X2=1.2 $Y2=0.97
r63 15 17 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=1.045 $Y=0.97
+ $X2=0.51 $Y2=0.97
r64 13 36 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.48 $Y=2.465
+ $X2=0.48 $Y2=1.135
r65 9 35 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.48 $Y=0.465 $X2=0.48
+ $Y2=0.805
r66 2 31 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.085
r67 2 22 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.905
r68 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.255 $X2=1.175 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_1%A 3 7 9 12 13 17
r33 12 15 49.7087 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.93 $Y=1.51
+ $X2=0.93 $Y2=1.695
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.51
+ $X2=0.93 $Y2=1.345
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=1.51 $X2=0.93 $Y2=1.51
r36 9 13 5.97563 $w=4.03e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=1.547
+ $X2=0.93 $Y2=1.547
r37 9 17 0.569108 $w=4.03e-07 $l=2e-08 $layer=LI1_cond $X=0.72 $Y=1.547 $X2=0.7
+ $Y2=1.547
r38 7 14 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.96 $Y=0.465
+ $X2=0.96 $Y2=1.345
r39 3 15 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.91 $Y=2.465 $X2=0.91
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_1%X 1 2 12 14 15 16 17 36 38
r20 23 38 0.557634 $w=3.08e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=1.68
+ $X2=0.24 $Y2=1.665
r21 17 33 5.0187 $w=3.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=2.775
+ $X2=0.24 $Y2=2.91
r22 16 17 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.775
r23 15 16 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r24 14 38 1.30115 $w=3.08e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.63
+ $X2=0.24 $Y2=1.665
r25 14 36 6.23675 $w=3.08e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=1.63
+ $X2=0.24 $Y2=1.525
r26 14 15 11.8962 $w=3.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.24 $Y=1.715
+ $X2=0.24 $Y2=2.035
r27 14 23 1.30115 $w=3.08e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.715
+ $X2=0.24 $Y2=1.68
r28 9 12 3.26812 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=0.17 $Y=0.467
+ $X2=0.265 $Y2=0.467
r29 7 9 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.17 $Y=0.635 $X2=0.17
+ $Y2=0.467
r30 7 36 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=0.17 $Y=0.635
+ $X2=0.17 $Y2=1.525
r31 2 33 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.91
r32 2 15 400 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.05
r33 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.255 $X2=0.265 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_1%VPWR 1 6 10 12 19 20 23
r20 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r21 17 23 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.695 $Y2=3.33
r22 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=1.2 $Y2=3.33
r23 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 12 23 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.695 $Y2=3.33
r25 12 14 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r26 10 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r27 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 10 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 6 9 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.695 $Y=2.085
+ $X2=0.695 $Y2=2.905
r30 4 23 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r31 4 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.905
r32 1 9 400 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.905
r33 1 6 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_1%VGND 1 6 8 10 17 18 21
r19 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r20 15 21 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.737
+ $Y2=0
r21 15 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r22 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r23 10 21 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.737
+ $Y2=0
r24 10 12 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.24
+ $Y2=0
r25 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r26 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r27 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r28 4 21 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0
r29 4 6 15.9247 $w=2.73e-07 $l=3.8e-07 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0.465
r30 1 6 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.255 $X2=0.745 $Y2=0.465
.ends

