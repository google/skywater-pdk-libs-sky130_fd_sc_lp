* File: sky130_fd_sc_lp__dlrbn_1.pex.spice
* Created: Fri Aug 28 10:25:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRBN_1%GATE_N 2 5 9 11 12 13 14 15 21
c31 5 0 9.43755e-20 $X=0.485 $Y=0.56
r32 21 23 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.417 $Y=1.38
+ $X2=0.417 $Y2=1.215
r33 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.395
+ $Y=1.38 $X2=0.395 $Y2=1.38
r34 14 15 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=2.035
r35 14 22 8.31509 $w=3.93e-07 $l=2.85e-07 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=1.38
r36 13 22 2.47994 $w=3.93e-07 $l=8.5e-08 $layer=LI1_cond $X=0.282 $Y=1.295
+ $X2=0.282 $Y2=1.38
r37 12 13 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=0.925
+ $X2=0.282 $Y2=1.295
r38 9 11 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=0.53 $Y=2.685 $X2=0.53
+ $Y2=1.885
r39 5 23 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.485 $Y=0.56
+ $X2=0.485 $Y2=1.215
r40 2 11 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.417 $Y=1.698
+ $X2=0.417 $Y2=1.885
r41 1 21 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.417 $Y=1.402
+ $X2=0.417 $Y2=1.38
r42 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.417 $Y=1.402
+ $X2=0.417 $Y2=1.698
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_112_70# 1 2 7 8 11 15 17 20 22 23 27 29 31
+ 33 36 38 42 44 46 49 50 53 57 58 59 60
c129 53 0 9.43755e-20 $X=0.7 $Y=0.505
c130 38 0 1.81888e-19 $X=2.785 $Y=2.49
c131 27 0 8.4529e-20 $X=3.075 $Y=1.045
r132 57 59 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.862 $Y=1.67
+ $X2=0.862 $Y2=1.505
r133 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.98
+ $Y=1.67 $X2=0.98 $Y2=1.67
r134 55 59 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=0.745 $Y=0.67
+ $X2=0.745 $Y2=1.505
r135 53 55 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.717 $Y=0.505
+ $X2=0.717 $Y2=0.67
r136 50 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.57 $Y=2.94 $X2=1.57
+ $Y2=3.03
r137 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=2.94 $X2=1.57 $Y2=2.94
r138 47 62 2.82016 $w=3e-07 $l=9.5e-08 $layer=LI1_cond $X=0.85 $Y=2.925
+ $X2=0.755 $Y2=2.925
r139 47 49 27.6586 $w=2.98e-07 $l=7.2e-07 $layer=LI1_cond $X=0.85 $Y=2.925
+ $X2=1.57 $Y2=2.925
r140 46 60 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=0.755 $Y=2.52
+ $X2=0.755 $Y2=2.175
r141 44 62 4.45288 $w=1.9e-07 $l=1.5e-07 $layer=LI1_cond $X=0.755 $Y=2.775
+ $X2=0.755 $Y2=2.925
r142 44 46 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=0.755 $Y=2.775
+ $X2=0.755 $Y2=2.52
r143 42 60 9.01764 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=0.862 $Y=1.973
+ $X2=0.862 $Y2=2.175
r144 41 57 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=0.862 $Y=1.707
+ $X2=0.862 $Y2=1.67
r145 41 42 7.56913 $w=4.03e-07 $l=2.66e-07 $layer=LI1_cond $X=0.862 $Y=1.707
+ $X2=0.862 $Y2=1.973
r146 34 36 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.785 $Y=1.735
+ $X2=3.075 $Y2=1.735
r147 32 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.98 $Y=1.655
+ $X2=0.98 $Y2=1.67
r148 29 31 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.465 $Y=2.415
+ $X2=3.465 $Y2=2.095
r149 25 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.075 $Y=1.66
+ $X2=3.075 $Y2=1.735
r150 25 27 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.075 $Y=1.66
+ $X2=3.075 $Y2=1.045
r151 24 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.86 $Y=2.49
+ $X2=2.785 $Y2=2.49
r152 23 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=2.49
+ $X2=3.465 $Y2=2.415
r153 23 24 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.39 $Y=2.49
+ $X2=2.86 $Y2=2.49
r154 21 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=2.565
+ $X2=2.785 $Y2=2.49
r155 21 22 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.785 $Y=2.565
+ $X2=2.785 $Y2=2.955
r156 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=2.415
+ $X2=2.785 $Y2=2.49
r157 19 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=1.81
+ $X2=2.785 $Y2=1.735
r158 19 20 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.785 $Y=1.81
+ $X2=2.785 $Y2=2.415
r159 18 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.735 $Y=3.03
+ $X2=1.57 $Y2=3.03
r160 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.71 $Y=3.03
+ $X2=2.785 $Y2=2.955
r161 17 18 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=2.71 $Y=3.03
+ $X2=1.735 $Y2=3.03
r162 13 33 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.71 $Y=1.655
+ $X2=1.695 $Y2=1.58
r163 13 15 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.71 $Y=1.655
+ $X2=1.71 $Y2=2.115
r164 9 33 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.68 $Y=1.505
+ $X2=1.695 $Y2=1.58
r165 9 11 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.68 $Y=1.505
+ $X2=1.68 $Y2=0.93
r166 8 32 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.145 $Y=1.58
+ $X2=0.98 $Y2=1.655
r167 7 33 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.605 $Y=1.58
+ $X2=1.695 $Y2=1.58
r168 7 8 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.605 $Y=1.58
+ $X2=1.145 $Y2=1.58
r169 2 62 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=2.365 $X2=0.745 $Y2=2.86
r170 2 46 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=2.365 $X2=0.745 $Y2=2.52
r171 1 53 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.35 $X2=0.7 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%D 1 3 6 8 9 17
c37 17 0 3.00579e-20 $X=2.295 $Y=1.415
c38 6 0 1.3134e-20 $X=2.295 $Y=2.115
r39 15 17 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.16 $Y=1.415
+ $X2=2.295 $Y2=1.415
r40 12 15 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.11 $Y=1.415 $X2=2.16
+ $Y2=1.415
r41 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.415 $X2=2.16 $Y2=1.415
r42 8 9 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.395 $X2=2.16
+ $Y2=1.395
r43 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.58
+ $X2=2.295 $Y2=1.415
r44 4 6 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.295 $Y=1.58
+ $X2=2.295 $Y2=2.115
r45 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.25
+ $X2=2.11 $Y2=1.415
r46 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.11 $Y=1.25 $X2=2.11
+ $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_207_40# 1 2 7 12 13 14 17 21 29 33 34 35
c81 34 0 3.00579e-20 $X=1.452 $Y=1.775
c82 33 0 1.3134e-20 $X=1.495 $Y=1.94
r83 33 34 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=1.452 $Y=1.94
+ $X2=1.452 $Y2=1.775
r84 29 31 5.96739 $w=2.76e-07 $l=1.35e-07 $layer=LI1_cond $X=1.33 $Y=0.9
+ $X2=1.465 $Y2=0.9
r85 24 29 3.57235 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.33 $Y=1.04 $X2=1.33
+ $Y2=0.9
r86 24 34 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.33 $Y=1.04
+ $X2=1.33 $Y2=1.775
r87 22 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.2 $Y=0.365 $X2=1.2
+ $Y2=0.275
r88 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=0.365 $X2=1.2 $Y2=0.365
r89 19 29 5.74638 $w=2.76e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=0.9 $X2=1.33
+ $Y2=0.9
r90 19 21 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.2 $Y=0.76 $X2=1.2
+ $Y2=0.365
r91 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.99 $Y=1.515
+ $X2=3.99 $Y2=2.205
r92 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.915 $Y=1.44
+ $X2=3.99 $Y2=1.515
r93 13 14 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.915 $Y=1.44
+ $X2=3.58 $Y2=1.44
r94 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.505 $Y=1.365
+ $X2=3.58 $Y2=1.44
r95 10 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.505 $Y=1.365
+ $X2=3.505 $Y2=1.045
r96 9 12 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.505 $Y=0.35
+ $X2=3.505 $Y2=1.045
r97 8 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.275
+ $X2=1.2 $Y2=0.275
r98 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.43 $Y=0.275
+ $X2=3.505 $Y2=0.35
r99 7 8 1058.86 $w=1.5e-07 $l=2.065e-06 $layer=POLY_cond $X=3.43 $Y=0.275
+ $X2=1.365 $Y2=0.275
r100 2 33 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.37
+ $Y=1.795 $X2=1.495 $Y2=1.94
r101 1 31 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.72 $X2=1.465 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_437_144# 1 2 8 9 10 13 15 17 19 22 25 27
+ 29 31 32 37 39
c92 22 0 2.08516e-20 $X=2.51 $Y=0.71
c93 19 0 2.50734e-20 $X=4.6 $Y=0.95
r94 35 37 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.325 $Y=0.875
+ $X2=2.51 $Y2=0.875
r95 32 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=0.35
+ $X2=3.955 $Y2=0.515
r96 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.955
+ $Y=0.35 $X2=3.955 $Y2=0.35
r97 29 31 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.595 $Y=0.35
+ $X2=3.955 $Y2=0.35
r98 25 39 5.8268 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=2.525 $Y=1.875
+ $X2=2.525 $Y2=1.775
r99 25 27 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.525 $Y=1.875
+ $X2=2.525 $Y2=1.94
r100 23 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.04
+ $X2=2.51 $Y2=0.875
r101 23 39 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.51 $Y=1.04
+ $X2=2.51 $Y2=1.775
r102 22 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=0.71
+ $X2=2.51 $Y2=0.875
r103 21 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.51 $Y=0.435
+ $X2=2.595 $Y2=0.35
r104 21 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.51 $Y=0.435
+ $X2=2.51 $Y2=0.71
r105 18 19 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.35 $Y=0.95
+ $X2=4.6 $Y2=0.95
r106 15 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.6 $Y=0.875
+ $X2=4.6 $Y2=0.95
r107 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.6 $Y=0.875
+ $X2=4.6 $Y2=0.555
r108 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.95
r109 11 13 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=2.205
r110 9 18 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.275 $Y=0.95
+ $X2=4.35 $Y2=0.95
r111 9 10 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=4.275 $Y=0.95
+ $X2=4.12 $Y2=0.95
r112 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.045 $Y=0.875
+ $X2=4.12 $Y2=0.95
r113 8 42 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.045 $Y=0.875
+ $X2=4.045 $Y2=0.515
r114 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.37
+ $Y=1.795 $X2=2.51 $Y2=1.94
r115 1 35 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.185
+ $Y=0.72 $X2=2.325 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_955_271# 1 2 9 13 17 19 21 24 26 28 29 32
+ 35 38 41 42 43 44 46 48 52 53 56 57 58 60 61 63 66 67 70 80
c171 66 0 5.00887e-20 $X=5.58 $Y=1.52
c172 35 0 1.81832e-20 $X=5.58 $Y=1.93
c173 19 0 4.11833e-20 $X=7.105 $Y=1.185
r174 64 80 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=8.745 $Y=1.425
+ $X2=8.905 $Y2=1.425
r175 64 77 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.745 $Y=1.425
+ $X2=8.655 $Y2=1.425
r176 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.745
+ $Y=1.425 $X2=8.745 $Y2=1.425
r177 61 63 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=8.435 $Y=1.425
+ $X2=8.745 $Y2=1.425
r178 60 61 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.35 $Y=1.26
+ $X2=8.435 $Y2=1.425
r179 59 60 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=8.35 $Y=0.425
+ $X2=8.35 $Y2=1.26
r180 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.265 $Y=0.34
+ $X2=8.35 $Y2=0.425
r181 57 58 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=8.265 $Y=0.34
+ $X2=7.08 $Y2=0.34
r182 56 70 4.14756 $w=2.2e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.99 $Y=0.83
+ $X2=6.95 $Y2=0.915
r183 55 58 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.99 $Y=0.425
+ $X2=7.08 $Y2=0.34
r184 55 56 24.9545 $w=1.78e-07 $l=4.05e-07 $layer=LI1_cond $X=6.99 $Y=0.425
+ $X2=6.99 $Y2=0.83
r185 53 76 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=6.985 $Y=1.35
+ $X2=7.105 $Y2=1.35
r186 53 74 13.7714 $w=3.15e-07 $l=9e-08 $layer=POLY_cond $X=6.985 $Y=1.35
+ $X2=6.895 $Y2=1.35
r187 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.985
+ $Y=1.35 $X2=6.985 $Y2=1.35
r188 50 70 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1 $X2=6.95
+ $Y2=0.915
r189 50 52 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=6.95 $Y=1 $X2=6.95
+ $Y2=1.35
r190 46 69 3.0159 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=6.172 $Y=2.1
+ $X2=6.172 $Y2=2.015
r191 46 48 41.4879 $w=2.23e-07 $l=8.1e-07 $layer=LI1_cond $X=6.172 $Y=2.1
+ $X2=6.172 $Y2=2.91
r192 45 67 3.35233 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.93 $Y=0.915
+ $X2=5.735 $Y2=0.915
r193 44 70 2.28545 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.82 $Y=0.915
+ $X2=6.95 $Y2=0.915
r194 44 45 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.82 $Y=0.915
+ $X2=5.93 $Y2=0.915
r195 42 69 3.9739 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=6.06 $Y=2.015
+ $X2=6.172 $Y2=2.015
r196 42 43 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.06 $Y=2.015
+ $X2=5.735 $Y2=2.015
r197 41 66 6.41553 $w=2.52e-07 $l=1.9139e-07 $layer=LI1_cond $X=5.637 $Y=1.355
+ $X2=5.58 $Y2=1.52
r198 40 67 3.22182 $w=2.92e-07 $l=1.33918e-07 $layer=LI1_cond $X=5.637 $Y=1
+ $X2=5.735 $Y2=0.915
r199 40 41 20.1911 $w=1.93e-07 $l=3.55e-07 $layer=LI1_cond $X=5.637 $Y=1
+ $X2=5.637 $Y2=1.355
r200 36 67 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0.83
+ $X2=5.735 $Y2=0.915
r201 36 38 13.0019 $w=3.88e-07 $l=4.4e-07 $layer=LI1_cond $X=5.735 $Y=0.83
+ $X2=5.735 $Y2=0.39
r202 35 43 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.58 $Y=1.93
+ $X2=5.735 $Y2=2.015
r203 34 66 6.41553 $w=2.52e-07 $l=1.65e-07 $layer=LI1_cond $X=5.58 $Y=1.685
+ $X2=5.58 $Y2=1.52
r204 34 35 9.10802 $w=3.08e-07 $l=2.45e-07 $layer=LI1_cond $X=5.58 $Y=1.685
+ $X2=5.58 $Y2=1.93
r205 32 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.94 $Y=1.52
+ $X2=4.94 $Y2=1.685
r206 32 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.94 $Y=1.52
+ $X2=4.94 $Y2=1.355
r207 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.94
+ $Y=1.52 $X2=4.94 $Y2=1.52
r208 29 66 0.398883 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=5.425 $Y=1.52
+ $X2=5.58 $Y2=1.52
r209 29 31 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=5.425 $Y=1.52
+ $X2=4.94 $Y2=1.52
r210 26 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.905 $Y=1.26
+ $X2=8.905 $Y2=1.425
r211 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.905 $Y=1.26
+ $X2=8.905 $Y2=0.73
r212 22 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=1.59
+ $X2=8.655 $Y2=1.425
r213 22 24 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=8.655 $Y=1.59
+ $X2=8.655 $Y2=2.465
r214 19 76 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.105 $Y=1.185
+ $X2=7.105 $Y2=1.35
r215 19 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.105 $Y=1.185
+ $X2=7.105 $Y2=0.865
r216 15 74 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.895 $Y=1.515
+ $X2=6.895 $Y2=1.35
r217 15 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.895 $Y=1.515
+ $X2=6.895 $Y2=2.155
r218 13 72 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.03 $Y=0.555
+ $X2=5.03 $Y2=1.355
r219 9 73 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.875 $Y=2.095
+ $X2=4.875 $Y2=1.685
r220 2 69 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=6.015
+ $Y=1.835 $X2=6.155 $Y2=2.095
r221 2 48 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.015
+ $Y=1.835 $X2=6.155 $Y2=2.91
r222 1 38 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=5.64
+ $Y=0.235 $X2=5.765 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_630_167# 1 2 7 10 11 12 13 15 18 20 22 23
+ 24 25 26 29 33 34 36
c111 22 0 1.81888e-19 $X=2.88 $Y=2.43
c112 12 0 1.19417e-19 $X=5.495 $Y=1.65
c113 10 0 2.80616e-20 $X=5.42 $Y=2.955
r114 36 38 7.92402 $w=4.08e-07 $l=2.65e-07 $layer=LI1_cond $X=3.51 $Y=2.452
+ $X2=3.775 $Y2=2.452
r115 34 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.51 $Y=2.94 $X2=3.51
+ $Y2=3.03
r116 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.51
+ $Y=2.94 $X2=3.51 $Y2=2.94
r117 31 36 1.98218 $w=3.3e-07 $l=2.58e-07 $layer=LI1_cond $X=3.51 $Y=2.71
+ $X2=3.51 $Y2=2.452
r118 31 33 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.51 $Y=2.71
+ $X2=3.51 $Y2=2.94
r119 27 29 20.744 $w=2.23e-07 $l=4.05e-07 $layer=LI1_cond $X=3.272 $Y=1.515
+ $X2=3.272 $Y2=1.11
r120 25 36 6.14407 $w=4.08e-07 $l=2.1609e-07 $layer=LI1_cond $X=3.345 $Y=2.57
+ $X2=3.51 $Y2=2.452
r121 25 26 15.6403 $w=2.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.345 $Y=2.57
+ $X2=2.965 $Y2=2.57
r122 23 27 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.16 $Y=1.6
+ $X2=3.272 $Y2=1.515
r123 23 24 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.16 $Y=1.6
+ $X2=2.965 $Y2=1.6
r124 22 26 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.88 $Y=2.43
+ $X2=2.965 $Y2=2.57
r125 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.88 $Y=1.685
+ $X2=2.965 $Y2=1.6
r126 21 22 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.88 $Y=1.685
+ $X2=2.88 $Y2=2.43
r127 16 20 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=5.98 $Y=1.575
+ $X2=5.96 $Y2=1.65
r128 16 18 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=5.98 $Y=1.575
+ $X2=5.98 $Y2=0.655
r129 13 20 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=5.94 $Y=1.725
+ $X2=5.96 $Y2=1.65
r130 13 15 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.94 $Y=1.725
+ $X2=5.94 $Y2=2.465
r131 11 20 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=5.865 $Y=1.65
+ $X2=5.96 $Y2=1.65
r132 11 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.865 $Y=1.65
+ $X2=5.495 $Y2=1.65
r133 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.42 $Y=1.725
+ $X2=5.495 $Y2=1.65
r134 9 10 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=5.42 $Y=1.725
+ $X2=5.42 $Y2=2.955
r135 8 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.675 $Y=3.03
+ $X2=3.51 $Y2=3.03
r136 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.345 $Y=3.03
+ $X2=5.42 $Y2=2.955
r137 7 8 856.319 $w=1.5e-07 $l=1.67e-06 $layer=POLY_cond $X=5.345 $Y=3.03
+ $X2=3.675 $Y2=3.03
r138 2 38 600 $w=1.7e-07 $l=5.80732e-07 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.885 $X2=3.775 $Y2=2.36
r139 1 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.835 $X2=3.29 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%RESET_B 3 7 9 11 18
c41 11 0 6.92449e-20 $X=6.48 $Y=1.665
c42 7 0 6.82718e-20 $X=6.37 $Y=2.465
r43 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.375
+ $X2=6.43 $Y2=1.54
r44 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.375
+ $X2=6.43 $Y2=1.21
r45 11 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.43
+ $Y=1.375 $X2=6.43 $Y2=1.375
r46 9 11 8.71718 $w=5.88e-07 $l=4.3e-07 $layer=LI1_cond $X=6 $Y=1.465 $X2=6.43
+ $Y2=1.465
r47 7 21 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=6.37 $Y=2.465
+ $X2=6.37 $Y2=1.54
r48 3 20 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.34 $Y=0.655
+ $X2=6.34 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_1394_367# 1 2 7 8 11 13 15 17 21 22 26 31
r47 29 31 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.415 $Y=0.87
+ $X2=7.53 $Y2=0.87
r48 24 26 7.49781 $w=6.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.11 $Y=2.15
+ $X2=7.53 $Y2=2.15
r49 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.56
+ $Y=1.74 $X2=7.56 $Y2=1.74
r50 19 26 6.10292 $w=2.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.53 $Y=1.815
+ $X2=7.53 $Y2=2.15
r51 19 21 3.20123 $w=2.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.53 $Y=1.815
+ $X2=7.53 $Y2=1.74
r52 18 31 1.91462 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.53 $Y=1.035
+ $X2=7.53 $Y2=0.87
r53 18 21 30.0916 $w=2.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.53 $Y=1.035
+ $X2=7.53 $Y2=1.74
r54 16 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.56 $Y=1.725
+ $X2=7.56 $Y2=1.74
r55 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.225 $Y=1.725
+ $X2=8.225 $Y2=1.65
r56 13 15 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.225 $Y=1.725
+ $X2=8.225 $Y2=2.465
r57 9 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.225 $Y=1.575
+ $X2=8.225 $Y2=1.65
r58 9 11 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=8.225 $Y=1.575
+ $X2=8.225 $Y2=0.73
r59 8 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.725 $Y=1.65
+ $X2=7.56 $Y2=1.725
r60 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.15 $Y=1.65
+ $X2=8.225 $Y2=1.65
r61 7 8 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=8.15 $Y=1.65
+ $X2=7.725 $Y2=1.65
r62 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.97
+ $Y=1.835 $X2=7.11 $Y2=1.98
r63 1 29 182 $w=1.7e-07 $l=3.25192e-07 $layer=licon1_NDIFF $count=1 $X=7.18
+ $Y=0.655 $X2=7.415 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%VPWR 1 2 3 4 5 6 19 21 25 28 31 35 37 41 47
+ 52 53 54 55 57 65 77 87 88 94 97 100 103
r119 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r120 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r122 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r123 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 88 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.4 $Y2=3.33
r125 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r126 85 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.545 $Y=3.33
+ $X2=8.415 $Y2=3.33
r127 85 87 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=8.545 $Y=3.33
+ $X2=9.36 $Y2=3.33
r128 84 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r129 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r130 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 81 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r132 80 83 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r134 78 100 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=6.632 $Y2=3.33
r135 78 80 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=6.96 $Y2=3.33
r136 77 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.285 $Y=3.33
+ $X2=8.415 $Y2=3.33
r137 77 83 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.285 $Y=3.33
+ $X2=7.92 $Y2=3.33
r138 76 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r140 73 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.565 $Y2=3.33
r141 73 75 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 72 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r144 69 72 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 69 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r146 68 71 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r147 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r148 66 94 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.075 $Y2=3.33
r149 66 68 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r150 65 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.565 $Y2=3.33
r151 65 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=3.33 $X2=4.08
+ $Y2=3.33
r152 64 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r153 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r154 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r155 61 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r156 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r157 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r158 58 91 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=3.33
+ $X2=0.24 $Y2=3.33
r159 58 60 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=3.33
+ $X2=0.72 $Y2=3.33
r160 57 94 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.075 $Y2=3.33
r161 57 63 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r162 55 76 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r163 55 98 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r164 53 75 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=5.56 $Y=3.33 $X2=5.52
+ $Y2=3.33
r165 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=3.33
+ $X2=5.725 $Y2=3.33
r166 51 52 5.76222 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.04 $Y=2.435
+ $X2=2.04 $Y2=2.605
r167 47 50 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=8.415 $Y=1.98
+ $X2=8.415 $Y2=2.95
r168 45 103 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.415 $Y=3.245
+ $X2=8.415 $Y2=3.33
r169 45 50 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=8.415 $Y=3.245
+ $X2=8.415 $Y2=2.95
r170 41 44 15.42 $w=3.53e-07 $l=4.75e-07 $layer=LI1_cond $X=6.632 $Y=2.015
+ $X2=6.632 $Y2=2.49
r171 39 100 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=6.632 $Y=3.245
+ $X2=6.632 $Y2=3.33
r172 39 44 24.5097 $w=3.53e-07 $l=7.55e-07 $layer=LI1_cond $X=6.632 $Y=3.245
+ $X2=6.632 $Y2=2.49
r173 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=5.725 $Y2=3.33
r174 37 100 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=6.632 $Y2=3.33
r175 37 38 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=5.89 $Y2=3.33
r176 33 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.725 $Y=3.245
+ $X2=5.725 $Y2=3.33
r177 33 35 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=5.725 $Y=3.245
+ $X2=5.725 $Y2=2.375
r178 29 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=3.33
r179 29 31 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=2.31
r180 28 94 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=3.33
r181 28 52 21.693 $w=3.38e-07 $l=6.4e-07 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=2.605
r182 25 51 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2 $Y=1.94 $X2=2
+ $Y2=2.435
r183 19 91 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.315 $Y=3.245
+ $X2=0.24 $Y2=3.33
r184 19 21 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=0.315 $Y=3.245
+ $X2=0.315 $Y2=2.51
r185 6 50 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.3
+ $Y=1.835 $X2=8.44 $Y2=2.95
r186 6 47 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.3
+ $Y=1.835 $X2=8.44 $Y2=1.98
r187 5 44 300 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=2 $X=6.445
+ $Y=1.835 $X2=6.585 $Y2=2.49
r188 5 41 600 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_PDIFF $count=1 $X=6.445
+ $Y=1.835 $X2=6.645 $Y2=2.015
r189 4 35 300 $w=1.7e-07 $l=5.9925e-07 $layer=licon1_PDIFF $count=2 $X=5.6
+ $Y=1.835 $X2=5.725 $Y2=2.375
r190 3 31 600 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.885 $X2=4.565 $Y2=2.31
r191 2 25 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=1.785
+ $Y=1.795 $X2=2 $Y2=1.94
r192 1 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.19
+ $Y=2.365 $X2=0.315 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_625_377# 1 2 7 9 14
r32 14 17 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.09 $Y=1.94
+ $X2=5.09 $Y2=2.095
r33 9 12 8.11948 $w=2.18e-07 $l=1.55e-07 $layer=LI1_cond $X=3.245 $Y=1.94
+ $X2=3.245 $Y2=2.095
r34 8 9 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.355 $Y=1.94 $X2=3.245
+ $Y2=1.94
r35 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=1.94
+ $X2=5.09 $Y2=1.94
r36 7 8 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=4.925 $Y=1.94
+ $X2=3.355 $Y2=1.94
r37 2 17 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.885 $X2=5.09 $Y2=2.095
r38 1 12 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=1.885 $X2=3.25 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%Q_N 1 2 7 8 9 10 11 12 22 32 34
r21 32 34 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=7.975 $Y=2.015
+ $X2=7.975 $Y2=2.035
r22 30 32 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=7.975 $Y=1.99
+ $X2=7.975 $Y2=2.015
r23 12 41 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=7.975 $Y=2.775
+ $X2=7.975 $Y2=2.91
r24 11 12 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=7.975 $Y=2.405
+ $X2=7.975 $Y2=2.775
r25 10 30 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=7.975 $Y=1.97
+ $X2=7.975 $Y2=1.99
r26 10 44 5.01554 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=7.975 $Y=1.97
+ $X2=7.975 $Y2=1.85
r27 10 11 14.4055 $w=2.78e-07 $l=3.5e-07 $layer=LI1_cond $X=7.975 $Y=2.055
+ $X2=7.975 $Y2=2.405
r28 10 34 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=7.975 $Y=2.055
+ $X2=7.975 $Y2=2.035
r29 9 44 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=7.965 $Y=1.665
+ $X2=7.965 $Y2=1.85
r30 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.965 $Y=1.295
+ $X2=7.965 $Y2=1.665
r31 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.965 $Y=0.925
+ $X2=7.965 $Y2=1.295
r32 7 22 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.965 $Y=0.925
+ $X2=7.965 $Y2=0.76
r33 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.835 $X2=8.01 $Y2=2.91
r34 2 32 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.835 $X2=8.01 $Y2=2.015
r35 1 22 182 $w=1.7e-07 $l=5.08675e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.31 $X2=8.01 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%Q 1 2 7 8 9 10 11 12 13 24 44 48
r21 48 49 4.40758 $w=7.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.14 $Y=1.98
+ $X2=9.14 $Y2=1.815
r22 22 44 0.876335 $w=5.03e-07 $l=3.7e-08 $layer=LI1_cond $X=9.262 $Y=0.888
+ $X2=9.262 $Y2=0.925
r23 13 41 2.15294 $w=7.48e-07 $l=1.35e-07 $layer=LI1_cond $X=9.14 $Y=2.775
+ $X2=9.14 $Y2=2.91
r24 12 13 5.90065 $w=7.48e-07 $l=3.7e-07 $layer=LI1_cond $X=9.14 $Y=2.405
+ $X2=9.14 $Y2=2.775
r25 12 35 3.42876 $w=7.48e-07 $l=2.15e-07 $layer=LI1_cond $X=9.14 $Y=2.405
+ $X2=9.14 $Y2=2.19
r26 11 35 2.4719 $w=7.48e-07 $l=1.55e-07 $layer=LI1_cond $X=9.14 $Y=2.035
+ $X2=9.14 $Y2=2.19
r27 11 48 0.877124 $w=7.48e-07 $l=5.5e-08 $layer=LI1_cond $X=9.14 $Y=2.035
+ $X2=9.14 $Y2=1.98
r28 10 49 3.90026 $w=4.58e-07 $l=1.5e-07 $layer=LI1_cond $X=9.285 $Y=1.665
+ $X2=9.285 $Y2=1.815
r29 9 10 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=9.285 $Y=1.295
+ $X2=9.285 $Y2=1.665
r30 9 46 4.03026 $w=4.58e-07 $l=1.55e-07 $layer=LI1_cond $X=9.285 $Y=1.295
+ $X2=9.285 $Y2=1.14
r31 8 46 4.6421 $w=5.03e-07 $l=1.91e-07 $layer=LI1_cond $X=9.262 $Y=0.949
+ $X2=9.262 $Y2=1.14
r32 8 44 0.568433 $w=5.03e-07 $l=2.4e-08 $layer=LI1_cond $X=9.262 $Y=0.949
+ $X2=9.262 $Y2=0.925
r33 8 22 0.568433 $w=5.03e-07 $l=2.4e-08 $layer=LI1_cond $X=9.262 $Y=0.864
+ $X2=9.262 $Y2=0.888
r34 7 8 7.31858 $w=5.03e-07 $l=3.09e-07 $layer=LI1_cond $X=9.262 $Y=0.555
+ $X2=9.262 $Y2=0.864
r35 7 24 2.36847 $w=5.03e-07 $l=1e-07 $layer=LI1_cond $X=9.262 $Y=0.555
+ $X2=9.262 $Y2=0.455
r36 2 48 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.73
+ $Y=1.835 $X2=8.87 $Y2=1.98
r37 2 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.73
+ $Y=1.835 $X2=8.87 $Y2=2.91
r38 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.98
+ $Y=0.31 $X2=9.12 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 45 60 75 76 82
c111 76 0 2.50734e-20 $X=9.36 $Y=0
r112 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r113 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r114 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r115 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r116 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r117 70 73 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r118 70 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r119 69 72 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r120 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r121 67 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.72 $Y=0 $X2=6.555
+ $Y2=0
r122 67 69 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.72 $Y=0 $X2=6.96
+ $Y2=0
r123 66 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r124 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r125 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r126 62 65 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r127 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r128 60 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.39 $Y=0 $X2=6.555
+ $Y2=0
r129 60 65 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.39 $Y=0 $X2=6
+ $Y2=0
r130 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r131 56 59 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r132 55 58 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r133 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r134 53 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r135 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r136 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r137 50 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r138 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r139 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r140 47 79 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0
+ $X2=0.217 $Y2=0
r141 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=0
+ $X2=0.72 $Y2=0
r142 45 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r143 45 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r144 43 72 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.605 $Y=0 $X2=8.4
+ $Y2=0
r145 43 44 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=8.605 $Y=0
+ $X2=8.722 $Y2=0
r146 42 75 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=9.36
+ $Y2=0
r147 42 44 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=8.722
+ $Y2=0
r148 40 58 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.685 $Y=0
+ $X2=4.56 $Y2=0
r149 40 41 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.685 $Y=0
+ $X2=4.802 $Y2=0
r150 39 62 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=5.04
+ $Y2=0
r151 39 41 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=4.802
+ $Y2=0
r152 37 52 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.68
+ $Y2=0
r153 37 38 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.91
+ $Y2=0
r154 36 55 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=2.16
+ $Y2=0
r155 36 38 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=1.91
+ $Y2=0
r156 32 44 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.722 $Y=0.085
+ $X2=8.722 $Y2=0
r157 32 34 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=8.722 $Y=0.085
+ $X2=8.722 $Y2=0.455
r158 28 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=0.085
+ $X2=6.555 $Y2=0
r159 28 30 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6.555 $Y=0.085
+ $X2=6.555 $Y2=0.54
r160 24 41 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.802 $Y=0.085
+ $X2=4.802 $Y2=0
r161 24 26 23.0489 $w=2.33e-07 $l=4.7e-07 $layer=LI1_cond $X=4.802 $Y=0.085
+ $X2=4.802 $Y2=0.555
r162 20 38 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=0.085
+ $X2=1.91 $Y2=0
r163 20 22 41.3832 $w=2.18e-07 $l=7.9e-07 $layer=LI1_cond $X=1.91 $Y=0.085
+ $X2=1.91 $Y2=0.875
r164 16 79 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r165 16 18 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.54
r166 5 34 91 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=2 $X=8.3
+ $Y=0.31 $X2=8.69 $Y2=0.455
r167 4 30 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.415
+ $Y=0.235 $X2=6.555 $Y2=0.54
r168 3 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.675
+ $Y=0.345 $X2=4.815 $Y2=0.555
r169 2 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.755
+ $Y=0.72 $X2=1.895 $Y2=0.875
r170 1 18 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.35 $X2=0.27 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_547_167# 1 2 9 11 12 14
r34 11 14 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=4.402 $Y=0.69
+ $X2=4.402 $Y2=0.555
r35 11 12 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=4.29 $Y=0.69
+ $X2=2.99 $Y2=0.69
r36 7 12 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=2.877 $Y=0.775
+ $X2=2.99 $Y2=0.69
r37 7 9 13.8293 $w=2.23e-07 $l=2.7e-07 $layer=LI1_cond $X=2.877 $Y=0.775
+ $X2=2.877 $Y2=1.045
r38 2 14 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.26
+ $Y=0.345 $X2=4.385 $Y2=0.555
r39 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.835 $X2=2.86 $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_1%A_716_167# 1 2 7 13
c23 7 0 1.19417e-19 $X=5.14 $Y=1.06
r24 11 13 19.5414 $w=2.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.255 $Y=0.945
+ $X2=5.255 $Y2=0.555
r25 7 11 6.81649 $w=2.3e-07 $l=1.62635e-07 $layer=LI1_cond $X=5.14 $Y=1.06
+ $X2=5.255 $Y2=0.945
r26 7 9 71.1508 $w=2.28e-07 $l=1.42e-06 $layer=LI1_cond $X=5.14 $Y=1.06 $X2=3.72
+ $Y2=1.06
r27 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.345 $X2=5.245 $Y2=0.555
r28 1 9 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.58
+ $Y=0.835 $X2=3.72 $Y2=1.05
.ends

