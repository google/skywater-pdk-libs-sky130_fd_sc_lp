* File: sky130_fd_sc_lp__or2_0.pxi.spice
* Created: Fri Aug 28 11:21:02 2020
* 
x_PM_SKY130_FD_SC_LP__OR2_0%B N_B_M1002_g N_B_M1000_g N_B_c_53_n N_B_c_54_n B B
+ B B N_B_c_56_n PM_SKY130_FD_SC_LP__OR2_0%B
x_PM_SKY130_FD_SC_LP__OR2_0%A N_A_M1004_g N_A_M1003_g N_A_c_86_n N_A_c_90_n A A
+ A N_A_c_88_n PM_SKY130_FD_SC_LP__OR2_0%A
x_PM_SKY130_FD_SC_LP__OR2_0%A_76_473# N_A_76_473#_M1002_d N_A_76_473#_M1000_s
+ N_A_76_473#_c_126_n N_A_76_473#_M1005_g N_A_76_473#_c_132_n
+ N_A_76_473#_M1001_g N_A_76_473#_c_127_n N_A_76_473#_c_134_n
+ N_A_76_473#_c_135_n N_A_76_473#_c_128_n N_A_76_473#_c_137_n
+ N_A_76_473#_c_138_n N_A_76_473#_c_129_n N_A_76_473#_c_130_n
+ N_A_76_473#_c_190_p N_A_76_473#_c_148_n N_A_76_473#_c_131_n
+ PM_SKY130_FD_SC_LP__OR2_0%A_76_473#
x_PM_SKY130_FD_SC_LP__OR2_0%VPWR N_VPWR_M1003_d N_VPWR_c_199_n VPWR
+ N_VPWR_c_200_n N_VPWR_c_201_n N_VPWR_c_198_n N_VPWR_c_203_n
+ PM_SKY130_FD_SC_LP__OR2_0%VPWR
x_PM_SKY130_FD_SC_LP__OR2_0%X N_X_M1005_d N_X_M1001_d N_X_c_222_n X X X X X X X
+ N_X_c_224_n X PM_SKY130_FD_SC_LP__OR2_0%X
x_PM_SKY130_FD_SC_LP__OR2_0%VGND N_VGND_M1002_s N_VGND_M1004_d N_VGND_c_246_n
+ N_VGND_c_247_n N_VGND_c_248_n N_VGND_c_249_n N_VGND_c_250_n VGND
+ N_VGND_c_251_n N_VGND_c_252_n N_VGND_c_253_n PM_SKY130_FD_SC_LP__OR2_0%VGND
cc_1 VNB N_B_M1002_g 0.0268875f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.445
cc_2 VNB N_B_M1000_g 0.00703342f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.575
cc_3 VNB N_B_c_53_n 0.028497f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.36
cc_4 VNB N_B_c_54_n 0.0252522f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.51
cc_5 VNB B 0.0444163f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B_c_56_n 0.0272703f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.005
cc_7 VNB N_A_M1004_g 0.0366587f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.84
cc_8 VNB N_A_c_86_n 0.0236732f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.36
cc_9 VNB A 0.00556132f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_10 VNB N_A_c_88_n 0.0170373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_76_473#_c_126_n 0.019992f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_12 VNB N_A_76_473#_c_127_n 0.0227365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_76_473#_c_128_n 0.0138947f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.005
cc_14 VNB N_A_76_473#_c_129_n 0.00524438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_76_473#_c_130_n 0.0211565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_76_473#_c_131_n 0.0354005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_198_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_X_c_222_n 0.0169827f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_19 VNB X 0.0550106f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.51
cc_20 VNB N_X_c_224_n 0.0218245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_246_n 0.0192624f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.575
cc_22 VNB N_VGND_c_247_n 0.0167181f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.36
cc_23 VNB N_VGND_c_248_n 0.00458801f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_VGND_c_249_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_250_n 0.00564902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_251_n 0.0261552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_252_n 0.153356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_253_n 0.00487954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_B_M1000_g 0.054135f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.575
cc_30 VPB B 0.0460389f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_31 VPB N_A_M1003_g 0.0413404f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_32 VPB N_A_c_90_n 0.0167617f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.51
cc_33 VPB A 0.00171403f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_34 VPB N_A_76_473#_c_132_n 0.0249679f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_35 VPB N_A_76_473#_M1001_g 0.0280986f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_36 VPB N_A_76_473#_c_134_n 0.0216669f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.005
cc_37 VPB N_A_76_473#_c_135_n 0.0145309f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.005
cc_38 VPB N_A_76_473#_c_128_n 0.00255257f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=1.005
cc_39 VPB N_A_76_473#_c_137_n 0.00168696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_76_473#_c_138_n 0.02288f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=1.665
cc_41 VPB N_A_76_473#_c_130_n 0.00300411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_199_n 0.0215101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_200_n 0.0361566f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.36
cc_44 VPB N_VPWR_c_201_n 0.0186467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_198_n 0.0698664f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_203_n 0.0119958f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.005
cc_47 VPB X 0.0359757f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.51
cc_48 VPB X 0.0236706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB X 0.0109972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 N_B_M1002_g N_A_M1004_g 0.0114572f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_51 N_B_c_53_n N_A_c_86_n 0.0114572f $X=0.565 $Y=1.36 $X2=0 $Y2=0
cc_52 N_B_c_54_n N_A_c_86_n 0.0396885f $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_53 N_B_M1000_g N_A_c_90_n 0.0396885f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_54 N_B_c_54_n A 4.11571e-19 $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_55 N_B_c_56_n N_A_c_88_n 0.0114572f $X=0.5 $Y=1.005 $X2=0 $Y2=0
cc_56 N_B_M1000_g N_A_76_473#_c_135_n 0.0147617f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_57 B N_A_76_473#_c_135_n 0.017394f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_B_M1002_g N_A_76_473#_c_128_n 0.00838173f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_59 N_B_M1000_g N_A_76_473#_c_128_n 0.00863736f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_60 N_B_c_54_n N_A_76_473#_c_128_n 0.00417902f $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_61 B N_A_76_473#_c_128_n 0.0908998f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_62 N_B_M1000_g N_A_76_473#_c_137_n 0.0106731f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_63 B N_A_76_473#_c_137_n 7.16836e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_64 N_B_M1000_g N_A_76_473#_c_148_n 0.00366679f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_65 B N_A_76_473#_c_148_n 0.0141002f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_B_M1000_g N_VPWR_c_199_n 0.0011934f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_67 N_B_M1000_g N_VPWR_c_200_n 0.00350693f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_68 N_B_M1000_g N_VPWR_c_198_n 0.00492109f $X=0.72 $Y=2.575 $X2=0 $Y2=0
cc_69 N_B_M1002_g N_VGND_c_246_n 0.00371677f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_70 B N_VGND_c_246_n 0.0236961f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_71 N_B_c_56_n N_VGND_c_246_n 0.00156251f $X=0.5 $Y=1.005 $X2=0 $Y2=0
cc_72 N_B_M1002_g N_VGND_c_247_n 0.00585385f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_73 N_B_M1002_g N_VGND_c_252_n 0.011925f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_74 B N_VGND_c_252_n 0.0100677f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_B_c_56_n N_VGND_c_252_n 2.54101e-19 $X=0.5 $Y=1.005 $X2=0 $Y2=0
cc_76 N_A_M1004_g N_A_76_473#_c_126_n 0.0192799f $X=1.11 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_A_76_473#_c_132_n 0.00921928f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_78 N_A_c_90_n N_A_76_473#_c_132_n 0.01176f $X=1.2 $Y=1.825 $X2=0 $Y2=0
cc_79 N_A_M1003_g N_A_76_473#_M1001_g 0.0067385f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_80 A N_A_76_473#_c_127_n 0.00338783f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A_M1003_g N_A_76_473#_c_135_n 0.00254019f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_82 N_A_M1004_g N_A_76_473#_c_128_n 0.0126208f $X=1.11 $Y=0.445 $X2=0 $Y2=0
cc_83 A N_A_76_473#_c_128_n 0.0770165f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A_M1003_g N_A_76_473#_c_137_n 0.00415668f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_A_76_473#_c_138_n 0.0168892f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_86 N_A_c_90_n N_A_76_473#_c_138_n 0.00123144f $X=1.2 $Y=1.825 $X2=0 $Y2=0
cc_87 A N_A_76_473#_c_138_n 0.0194429f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_A_76_473#_c_129_n 7.04645e-19 $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_89 N_A_c_86_n N_A_76_473#_c_129_n 0.00117524f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_90 A N_A_76_473#_c_129_n 0.0176218f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_91 N_A_c_86_n N_A_76_473#_c_130_n 0.01176f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_92 N_A_M1004_g N_A_76_473#_c_131_n 0.00553232f $X=1.11 $Y=0.445 $X2=0 $Y2=0
cc_93 A N_A_76_473#_c_131_n 0.00872714f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_94 N_A_c_88_n N_A_76_473#_c_131_n 0.01176f $X=1.2 $Y=1.32 $X2=0 $Y2=0
cc_95 N_A_M1003_g N_VPWR_c_199_n 0.0130803f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_96 N_A_M1003_g N_VPWR_c_200_n 0.00382362f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_97 N_A_M1003_g N_VPWR_c_198_n 0.00413371f $X=1.11 $Y=2.575 $X2=0 $Y2=0
cc_98 N_A_M1004_g N_VGND_c_247_n 0.00585385f $X=1.11 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_M1004_g N_VGND_c_248_n 0.00169565f $X=1.11 $Y=0.445 $X2=0 $Y2=0
cc_100 A N_VGND_c_248_n 0.0129121f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_101 N_A_c_88_n N_VGND_c_248_n 5.3343e-19 $X=1.2 $Y=1.32 $X2=0 $Y2=0
cc_102 N_A_M1004_g N_VGND_c_252_n 0.00836958f $X=1.11 $Y=0.445 $X2=0 $Y2=0
cc_103 A N_VGND_c_252_n 0.00375588f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_104 N_A_76_473#_c_135_n A_159_473# 0.00453138f $X=0.765 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_105 N_A_76_473#_c_137_n A_159_473# 4.02591e-19 $X=0.85 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_106 N_A_76_473#_M1001_g N_VPWR_c_199_n 0.00910437f $X=1.88 $Y=2.685 $X2=0
+ $Y2=0
cc_107 N_A_76_473#_c_134_n N_VPWR_c_199_n 0.00140008f $X=1.792 $Y=2.175 $X2=0
+ $Y2=0
cc_108 N_A_76_473#_c_135_n N_VPWR_c_199_n 0.0227412f $X=0.765 $Y=2.575 $X2=0
+ $Y2=0
cc_109 N_A_76_473#_c_137_n N_VPWR_c_199_n 0.00406639f $X=0.85 $Y=2.41 $X2=0
+ $Y2=0
cc_110 N_A_76_473#_c_138_n N_VPWR_c_199_n 0.0532054f $X=1.605 $Y=2.09 $X2=0
+ $Y2=0
cc_111 N_A_76_473#_c_135_n N_VPWR_c_200_n 0.0109112f $X=0.765 $Y=2.575 $X2=0
+ $Y2=0
cc_112 N_A_76_473#_M1001_g N_VPWR_c_201_n 0.00499542f $X=1.88 $Y=2.685 $X2=0
+ $Y2=0
cc_113 N_A_76_473#_M1001_g N_VPWR_c_198_n 0.0106025f $X=1.88 $Y=2.685 $X2=0
+ $Y2=0
cc_114 N_A_76_473#_c_135_n N_VPWR_c_198_n 0.0180395f $X=0.765 $Y=2.575 $X2=0
+ $Y2=0
cc_115 N_A_76_473#_c_126_n N_X_c_222_n 0.00120654f $X=1.54 $Y=0.765 $X2=0 $Y2=0
cc_116 N_A_76_473#_c_127_n N_X_c_222_n 0.00665903f $X=1.68 $Y=0.84 $X2=0 $Y2=0
cc_117 N_A_76_473#_c_126_n X 0.00241133f $X=1.54 $Y=0.765 $X2=0 $Y2=0
cc_118 N_A_76_473#_M1001_g X 0.00656841f $X=1.88 $Y=2.685 $X2=0 $Y2=0
cc_119 N_A_76_473#_c_127_n X 0.0235263f $X=1.68 $Y=0.84 $X2=0 $Y2=0
cc_120 N_A_76_473#_c_138_n X 0.0140122f $X=1.605 $Y=2.09 $X2=0 $Y2=0
cc_121 N_A_76_473#_c_129_n X 0.0382513f $X=1.77 $Y=1.67 $X2=0 $Y2=0
cc_122 N_A_76_473#_c_130_n X 0.017393f $X=1.77 $Y=1.67 $X2=0 $Y2=0
cc_123 N_A_76_473#_M1001_g X 9.14762e-19 $X=1.88 $Y=2.685 $X2=0 $Y2=0
cc_124 N_A_76_473#_c_134_n X 0.00114427f $X=1.792 $Y=2.175 $X2=0 $Y2=0
cc_125 N_A_76_473#_c_190_p N_VGND_c_247_n 0.0127695f $X=0.895 $Y=0.445 $X2=0
+ $Y2=0
cc_126 N_A_76_473#_c_126_n N_VGND_c_248_n 0.0031247f $X=1.54 $Y=0.765 $X2=0
+ $Y2=0
cc_127 N_A_76_473#_c_126_n N_VGND_c_251_n 0.00585385f $X=1.54 $Y=0.765 $X2=0
+ $Y2=0
cc_128 N_A_76_473#_M1002_d N_VGND_c_252_n 0.00302605f $X=0.755 $Y=0.235 $X2=0
+ $Y2=0
cc_129 N_A_76_473#_c_126_n N_VGND_c_252_n 0.0121782f $X=1.54 $Y=0.765 $X2=0
+ $Y2=0
cc_130 N_A_76_473#_c_190_p N_VGND_c_252_n 0.0098423f $X=0.895 $Y=0.445 $X2=0
+ $Y2=0
cc_131 N_VPWR_c_201_n X 0.0194758f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_132 N_VPWR_c_198_n X 0.0135686f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_133 N_VPWR_c_199_n X 0.03028f $X=1.325 $Y=2.51 $X2=0 $Y2=0
cc_134 N_X_c_222_n N_VGND_c_251_n 0.0239649f $X=2.055 $Y=0.477 $X2=0 $Y2=0
cc_135 N_X_c_224_n N_VGND_c_251_n 0.0160903f $X=2.185 $Y=0.675 $X2=0 $Y2=0
cc_136 N_X_M1005_d N_VGND_c_252_n 0.00222801f $X=1.615 $Y=0.235 $X2=0 $Y2=0
cc_137 N_X_c_222_n N_VGND_c_252_n 0.0164422f $X=2.055 $Y=0.477 $X2=0 $Y2=0
cc_138 N_X_c_224_n N_VGND_c_252_n 0.00998544f $X=2.185 $Y=0.675 $X2=0 $Y2=0
