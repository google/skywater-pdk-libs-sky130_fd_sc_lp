# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__srdlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__srdlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.785000 1.315000 1.115000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.675000 0.255000 9.005000 1.135000 ;
        RECT 8.675000 1.815000 9.005000 3.075000 ;
        RECT 8.835000 1.135000 9.005000 1.815000 ;
    END
  END Q
  PIN SLEEP_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.015000 0.775000 7.555000 1.410000 ;
    END
  END SLEEP_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.845000 6.410000 1.780000 ;
    END
  END GATE
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 9.050000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 9.120000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 9.310000 3.520000 ;
        RECT  5.125000 1.495000 7.490000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 1.335000 ;
      RECT 0.115000  2.395000 0.365000 3.245000 ;
      RECT 0.535000  0.875000 0.795000 1.285000 ;
      RECT 0.535000  1.285000 2.950000 1.455000 ;
      RECT 0.535000  1.455000 0.705000 2.395000 ;
      RECT 0.535000  2.395000 0.875000 3.075000 ;
      RECT 0.875000  1.625000 2.640000 1.795000 ;
      RECT 0.875000  1.795000 1.205000 1.955000 ;
      RECT 1.110000  2.435000 2.105000 2.605000 ;
      RECT 1.110000  2.605000 1.440000 3.075000 ;
      RECT 1.165000  0.255000 1.655000 0.615000 ;
      RECT 1.485000  0.615000 2.190000 0.785000 ;
      RECT 1.610000  2.775000 1.940000 3.245000 ;
      RECT 1.775000  1.965000 2.105000 2.435000 ;
      RECT 1.825000  0.085000 2.155000 0.445000 ;
      RECT 1.860000  0.785000 2.190000 1.095000 ;
      RECT 2.310000  1.795000 2.640000 1.955000 ;
      RECT 2.310000  1.955000 2.480000 2.905000 ;
      RECT 2.310000  2.905000 4.375000 3.075000 ;
      RECT 2.360000  0.255000 2.690000 0.505000 ;
      RECT 2.360000  0.505000 3.290000 0.675000 ;
      RECT 2.620000  1.055000 2.950000 1.285000 ;
      RECT 2.650000  2.445000 2.980000 2.735000 ;
      RECT 2.810000  1.625000 3.290000 1.795000 ;
      RECT 2.810000  1.795000 2.980000 2.445000 ;
      RECT 3.120000  0.675000 3.290000 1.625000 ;
      RECT 3.150000  1.965000 3.475000 2.905000 ;
      RECT 3.460000  0.255000 3.790000 0.845000 ;
      RECT 3.460000  0.845000 5.275000 1.015000 ;
      RECT 3.690000  1.015000 3.860000 2.075000 ;
      RECT 3.690000  2.075000 4.020000 2.735000 ;
      RECT 4.045000  1.185000 4.375000 1.515000 ;
      RECT 4.205000  1.515000 4.375000 2.075000 ;
      RECT 4.205000  2.075000 6.830000 2.245000 ;
      RECT 4.205000  2.245000 4.375000 2.905000 ;
      RECT 4.585000  1.575000 5.615000 1.905000 ;
      RECT 4.640000  0.085000 4.970000 0.675000 ;
      RECT 4.710000  2.415000 5.155000 2.720000 ;
      RECT 4.710000  2.720000 6.145000 2.890000 ;
      RECT 4.710000  2.890000 5.155000 3.075000 ;
      RECT 4.945000  1.015000 5.275000 1.175000 ;
      RECT 5.430000  0.255000 5.760000 0.675000 ;
      RECT 5.445000  0.675000 5.615000 1.575000 ;
      RECT 5.815000  2.415000 6.145000 2.525000 ;
      RECT 5.815000  2.525000 7.330000 2.695000 ;
      RECT 5.815000  2.695000 6.145000 2.720000 ;
      RECT 5.990000  0.255000 6.320000 0.505000 ;
      RECT 5.990000  0.505000 6.830000 0.675000 ;
      RECT 6.580000  0.675000 6.830000 2.075000 ;
      RECT 6.580000  2.245000 6.830000 2.335000 ;
      RECT 7.000000  1.655000 7.330000 2.525000 ;
      RECT 7.140000  0.085000 7.470000 0.605000 ;
      RECT 7.630000  1.815000 7.960000 2.495000 ;
      RECT 7.700000  0.255000 8.030000 0.605000 ;
      RECT 7.790000  0.605000 8.030000 1.315000 ;
      RECT 7.790000  1.315000 8.665000 1.645000 ;
      RECT 7.790000  1.645000 7.960000 1.815000 ;
      RECT 8.175000  1.815000 8.505000 3.245000 ;
      RECT 8.245000  0.085000 8.495000 1.135000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  2.735000 5.125000 2.905000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__srdlxtp_1
END LIBRARY
