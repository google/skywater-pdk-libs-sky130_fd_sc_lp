* File: sky130_fd_sc_lp__xnor3_lp.pxi.spice
* Created: Wed Sep  2 10:40:48 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A N_A_M1004_g N_A_M1024_g N_A_M1018_g A
+ N_A_c_175_n PM_SKY130_FD_SC_LP__XNOR3_LP%A
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A_27_109# N_A_27_109#_M1004_s N_A_27_109#_M1023_d
+ N_A_27_109#_M1024_s N_A_27_109#_M1006_d N_A_27_109#_c_213_n
+ N_A_27_109#_M1010_g N_A_27_109#_M1020_g N_A_27_109#_M1015_g
+ N_A_27_109#_c_216_n N_A_27_109#_c_236_n N_A_27_109#_c_217_n
+ N_A_27_109#_c_218_n N_A_27_109#_c_219_n N_A_27_109#_c_220_n
+ N_A_27_109#_c_221_n N_A_27_109#_c_222_n N_A_27_109#_c_223_n
+ N_A_27_109#_c_224_n N_A_27_109#_c_225_n N_A_27_109#_c_226_n
+ N_A_27_109#_c_227_n N_A_27_109#_c_228_n N_A_27_109#_c_229_n
+ N_A_27_109#_c_230_n N_A_27_109#_c_271_p N_A_27_109#_c_231_n
+ N_A_27_109#_c_237_n N_A_27_109#_c_232_n N_A_27_109#_c_233_n
+ N_A_27_109#_c_234_n PM_SKY130_FD_SC_LP__XNOR3_LP%A_27_109#
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A_647_367# N_A_647_367#_M1021_d
+ N_A_647_367#_M1003_d N_A_647_367#_c_369_n N_A_647_367#_c_370_n
+ N_A_647_367#_c_371_n N_A_647_367#_M1011_g N_A_647_367#_c_372_n
+ N_A_647_367#_M1008_g N_A_647_367#_c_374_n N_A_647_367#_M1006_g
+ N_A_647_367#_M1023_g N_A_647_367#_c_377_n N_A_647_367#_c_378_n
+ N_A_647_367#_c_388_n N_A_647_367#_c_379_n N_A_647_367#_c_380_n
+ N_A_647_367#_c_381_n N_A_647_367#_c_382_n
+ PM_SKY130_FD_SC_LP__XNOR3_LP%A_647_367#
x_PM_SKY130_FD_SC_LP__XNOR3_LP%B N_B_M1012_g N_B_M1003_g N_B_M1021_g N_B_c_482_n
+ N_B_c_483_n N_B_M1014_g N_B_c_485_n N_B_M1026_g N_B_c_486_n N_B_M1025_g
+ N_B_c_477_n N_B_M1016_g N_B_c_478_n N_B_c_490_n N_B_c_491_n B B N_B_c_479_n
+ N_B_c_480_n PM_SKY130_FD_SC_LP__XNOR3_LP%B
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A_1318_85# N_A_1318_85#_M1017_s
+ N_A_1318_85#_M1000_s N_A_1318_85#_M1002_g N_A_1318_85#_M1007_g
+ N_A_1318_85#_c_600_n N_A_1318_85#_c_601_n N_A_1318_85#_c_602_n
+ N_A_1318_85#_c_595_n N_A_1318_85#_c_596_n N_A_1318_85#_c_604_n
+ N_A_1318_85#_c_597_n N_A_1318_85#_c_598_n
+ PM_SKY130_FD_SC_LP__XNOR3_LP%A_1318_85#
x_PM_SKY130_FD_SC_LP__XNOR3_LP%C N_C_c_683_n N_C_M1005_g N_C_M1022_g N_C_c_685_n
+ N_C_c_686_n N_C_M1017_g N_C_c_687_n N_C_c_688_n N_C_M1009_g N_C_M1000_g
+ N_C_c_690_n C N_C_c_691_n N_C_c_692_n N_C_c_693_n
+ PM_SKY130_FD_SC_LP__XNOR3_LP%C
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A_1348_111# N_A_1348_111#_M1002_d
+ N_A_1348_111#_M1007_d N_A_1348_111#_M1001_g N_A_1348_111#_c_759_n
+ N_A_1348_111#_M1013_g N_A_1348_111#_c_761_n N_A_1348_111#_c_762_n
+ N_A_1348_111#_M1019_g N_A_1348_111#_c_763_n N_A_1348_111#_c_764_n
+ N_A_1348_111#_c_770_n N_A_1348_111#_c_765_n N_A_1348_111#_c_766_n
+ N_A_1348_111#_c_767_n PM_SKY130_FD_SC_LP__XNOR3_LP%A_1348_111#
x_PM_SKY130_FD_SC_LP__XNOR3_LP%VPWR N_VPWR_M1024_d N_VPWR_M1003_s N_VPWR_M1000_d
+ N_VPWR_c_841_n N_VPWR_c_842_n N_VPWR_c_843_n N_VPWR_c_844_n N_VPWR_c_845_n
+ VPWR N_VPWR_c_846_n N_VPWR_c_847_n N_VPWR_c_848_n N_VPWR_c_840_n
+ N_VPWR_c_850_n N_VPWR_c_851_n PM_SKY130_FD_SC_LP__XNOR3_LP%VPWR
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A_265_409# N_A_265_409#_M1015_d
+ N_A_265_409#_M1008_d N_A_265_409#_M1010_d N_A_265_409#_M1011_d
+ N_A_265_409#_c_908_n N_A_265_409#_c_905_n N_A_265_409#_c_910_n
+ N_A_265_409#_c_906_n N_A_265_409#_c_911_n N_A_265_409#_c_912_n
+ N_A_265_409#_c_907_n PM_SKY130_FD_SC_LP__XNOR3_LP%A_265_409#
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A_763_347# N_A_763_347#_M1026_d
+ N_A_763_347#_M1005_d N_A_763_347#_M1011_s N_A_763_347#_M1016_d
+ N_A_763_347#_c_975_n N_A_763_347#_c_976_n N_A_763_347#_c_987_n
+ N_A_763_347#_c_1006_n N_A_763_347#_c_977_n N_A_763_347#_c_972_n
+ N_A_763_347#_c_978_n N_A_763_347#_c_979_n N_A_763_347#_c_973_n
+ N_A_763_347#_c_981_n N_A_763_347#_c_1034_n N_A_763_347#_c_982_n
+ N_A_763_347#_c_983_n N_A_763_347#_c_984_n N_A_763_347#_c_985_n
+ N_A_763_347#_c_974_n PM_SKY130_FD_SC_LP__XNOR3_LP%A_763_347#
x_PM_SKY130_FD_SC_LP__XNOR3_LP%A_803_81# N_A_803_81#_M1008_s N_A_803_81#_M1025_d
+ N_A_803_81#_M1014_d N_A_803_81#_M1022_d N_A_803_81#_c_1112_n
+ N_A_803_81#_c_1105_n N_A_803_81#_c_1106_n N_A_803_81#_c_1127_n
+ N_A_803_81#_c_1119_n N_A_803_81#_c_1129_n N_A_803_81#_c_1107_n
+ N_A_803_81#_c_1144_n N_A_803_81#_c_1146_n N_A_803_81#_c_1140_n
+ N_A_803_81#_c_1141_n N_A_803_81#_c_1109_n
+ PM_SKY130_FD_SC_LP__XNOR3_LP%A_803_81#
x_PM_SKY130_FD_SC_LP__XNOR3_LP%X N_X_M1019_d N_X_M1013_d N_X_c_1186_n X X X X X
+ PM_SKY130_FD_SC_LP__XNOR3_LP%X
x_PM_SKY130_FD_SC_LP__XNOR3_LP%VGND N_VGND_M1018_d N_VGND_M1012_s N_VGND_M1009_d
+ N_VGND_c_1208_n N_VGND_c_1209_n N_VGND_c_1265_n N_VGND_c_1210_n
+ N_VGND_c_1211_n N_VGND_c_1212_n N_VGND_c_1213_n N_VGND_c_1214_n
+ N_VGND_c_1215_n VGND N_VGND_c_1216_n N_VGND_c_1217_n N_VGND_c_1218_n
+ N_VGND_c_1219_n PM_SKY130_FD_SC_LP__XNOR3_LP%VGND
cc_1 VNB N_A_M1004_g 0.0456538f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.755
cc_2 VNB N_A_M1018_g 0.0347404f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.755
cc_3 VNB N_A_c_175_n 0.0143985f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.68
cc_4 VNB N_A_27_109#_c_213_n 0.0520743f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_A_27_109#_M1020_g 0.0191304f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_6 VNB N_A_27_109#_M1015_g 0.0231958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_109#_c_216_n 0.0285726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_109#_c_217_n 0.0181973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_109#_c_218_n 0.00209696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_109#_c_219_n 0.0201529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_109#_c_220_n 0.00269587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_109#_c_221_n 0.0122714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_109#_c_222_n 0.0200151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_109#_c_223_n 0.00406403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_109#_c_224_n 0.00207709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_109#_c_225_n 0.0152717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_109#_c_226_n 0.00270549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_109#_c_227_n 0.0049546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_109#_c_228_n 0.00404134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_109#_c_229_n 0.00264729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_109#_c_230_n 0.0052068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_109#_c_231_n 0.0132078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_109#_c_232_n 0.0150186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_109#_c_233_n 0.00138224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_109#_c_234_n 0.00293524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_647_367#_c_369_n 0.147448f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.515
cc_27 VNB N_A_647_367#_c_370_n 0.0126891f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.755
cc_28 VNB N_A_647_367#_c_371_n 0.0113973f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.755
cc_29 VNB N_A_647_367#_c_372_n 0.0115547f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_30 VNB N_A_647_367#_M1008_g 0.0249254f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_31 VNB N_A_647_367#_c_374_n 0.00963847f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.68
cc_32 VNB N_A_647_367#_M1006_g 0.00832693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_647_367#_M1023_g 0.0322353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_647_367#_c_377_n 0.0107476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_647_367#_c_378_n 0.00691193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_647_367#_c_379_n 0.00238391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_647_367#_c_380_n 0.00547302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_647_367#_c_381_n 0.0303554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_647_367#_c_382_n 0.0631724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B_M1012_g 0.0396506f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.755
cc_41 VNB N_B_M1021_g 0.0335606f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.755
cc_42 VNB N_B_M1026_g 0.0244559f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.68
cc_43 VNB N_B_M1025_g 0.038199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_B_c_477_n 0.00311814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_B_c_478_n 0.0073337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_B_c_479_n 0.0160791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_B_c_480_n 0.0343154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1318_85#_M1002_g 0.0357935f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.515
cc_49 VNB N_A_1318_85#_c_595_n 0.00961179f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=1.515
cc_50 VNB N_A_1318_85#_c_596_n 0.00309805f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_51 VNB N_A_1318_85#_c_597_n 0.00950626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1318_85#_c_598_n 0.0156997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_C_c_683_n 0.0190497f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_54 VNB N_C_M1022_g 0.021026f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.545
cc_55 VNB N_C_c_685_n 0.0263857f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.515
cc_56 VNB N_C_c_686_n 0.0202524f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.755
cc_57 VNB N_C_c_687_n 0.0153648f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_58 VNB N_C_c_688_n 0.0152683f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.68
cc_59 VNB N_C_M1000_g 0.0236262f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.515
cc_60 VNB N_C_c_690_n 0.0243097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_C_c_691_n 0.00920737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_C_c_692_n 0.0212785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_C_c_693_n 0.0417753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1348_111#_M1001_g 0.0264947f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=0.755
cc_65 VNB N_A_1348_111#_c_759_n 0.0125621f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=0.755
cc_66 VNB N_A_1348_111#_M1013_g 0.00588936f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_67 VNB N_A_1348_111#_c_761_n 0.0250795f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.68
cc_68 VNB N_A_1348_111#_c_762_n 0.0185152f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_69 VNB N_A_1348_111#_c_763_n 0.00576752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1348_111#_c_764_n 0.00355529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1348_111#_c_765_n 0.00174851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1348_111#_c_766_n 0.0391384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1348_111#_c_767_n 0.0510707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VPWR_c_840_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_265_409#_c_905_n 0.0110284f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_76 VNB N_A_265_409#_c_906_n 0.0138605f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_77 VNB N_A_265_409#_c_907_n 0.00320884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_763_347#_c_972_n 0.00183185f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.68
cc_79 VNB N_A_763_347#_c_973_n 0.00627459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_763_347#_c_974_n 0.0076588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_803_81#_c_1105_n 0.0222608f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_82 VNB N_A_803_81#_c_1106_n 7.16783e-19 $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_83 VNB N_A_803_81#_c_1107_n 0.0105955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_X_c_1186_n 0.0246849f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.515
cc_85 VNB X 0.0205443f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.755
cc_86 VNB X 0.00970466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1208_n 0.0172597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1209_n 0.0103244f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_89 VNB N_VGND_c_1210_n 0.0122113f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.68
cc_90 VNB N_VGND_c_1211_n 0.0291263f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.68
cc_91 VNB N_VGND_c_1212_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1213_n 0.0110506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1214_n 0.156593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1215_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1216_n 0.0330959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1217_n 0.0183931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1218_n 0.55426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1219_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VPB N_A_M1024_g 0.0335362f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.545
cc_100 VPB A 0.0019293f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_101 VPB N_A_c_175_n 0.0227619f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.68
cc_102 VPB N_A_27_109#_c_213_n 0.0665258f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_103 VPB N_A_27_109#_c_236_n 0.0390561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_27_109#_c_237_n 0.0166013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_27_109#_c_232_n 0.0177563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_27_109#_c_233_n 0.00174692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_647_367#_c_371_n 0.0121847f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.755
cc_108 VPB N_A_647_367#_M1011_g 0.0273564f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.68
cc_109 VPB N_A_647_367#_c_372_n 0.0134281f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.68
cc_110 VPB N_A_647_367#_M1006_g 0.022172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_647_367#_c_377_n 5.30645e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_647_367#_c_388_n 0.00639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_647_367#_c_379_n 0.003848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_647_367#_c_381_n 0.00749467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_B_M1003_g 0.0328758f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_B_c_482_n 0.12741f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_117 VPB N_B_c_483_n 0.0174968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_B_M1014_g 0.00518358f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.68
cc_119 VPB N_B_c_485_n 0.0161004f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.515
cc_120 VPB N_B_c_486_n 0.0750488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_B_c_477_n 0.0078793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_B_M1016_g 0.0294179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_B_c_478_n 0.00771784f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_B_c_490_n 0.0109283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_B_c_491_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_B_c_479_n 0.0164299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_B_c_480_n 0.0104669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_1318_85#_M1007_g 0.0330777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_1318_85#_c_600_n 0.0872756f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.68
cc_130 VPB N_A_1318_85#_c_601_n 0.0151171f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.68
cc_131 VPB N_A_1318_85#_c_602_n 0.074666f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.68
cc_132 VPB N_A_1318_85#_c_595_n 0.0116418f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.515
cc_133 VPB N_A_1318_85#_c_604_n 0.0121225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_1318_85#_c_597_n 0.00228217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_1318_85#_c_598_n 0.0210368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_C_M1022_g 0.0262785f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.545
cc_137 VPB N_C_M1000_g 0.0372662f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.515
cc_138 VPB N_A_1348_111#_M1013_g 0.0446209f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_139 VPB N_A_1348_111#_c_763_n 0.00138308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_1348_111#_c_770_n 0.00435015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_841_n 0.0092266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_842_n 0.0293698f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.68
cc_143 VPB N_VPWR_c_843_n 0.0142099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_844_n 0.0217494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_845_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_846_n 0.0439257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_847_n 0.145582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_848_n 0.0259642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_840_n 0.108939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_850_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_851_n 0.00546719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_265_409#_c_908_n 0.0270547f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.68
cc_153 VPB N_A_265_409#_c_905_n 0.0123131f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.68
cc_154 VPB N_A_265_409#_c_910_n 0.0541261f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.68
cc_155 VPB N_A_265_409#_c_911_n 0.00160975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_265_409#_c_912_n 0.0251117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_763_347#_c_975_n 0.0204265f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_158 VPB N_A_763_347#_c_976_n 0.00264153f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.68
cc_159 VPB N_A_763_347#_c_977_n 0.0179529f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.68
cc_160 VPB N_A_763_347#_c_978_n 0.00228216f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_763_347#_c_979_n 0.0151226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_763_347#_c_973_n 0.00275402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_763_347#_c_981_n 0.00816879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_763_347#_c_982_n 0.00928937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_763_347#_c_983_n 0.014632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_763_347#_c_984_n 8.29094e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_763_347#_c_985_n 0.00224482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_803_81#_c_1107_n 0.00134894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_803_81#_c_1109_n 0.00160028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB X 0.0486214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB X 0.0250801f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.68
cc_172 N_A_M1024_g N_A_27_109#_c_213_n 0.0133515f $X=0.67 $Y=2.545 $X2=0 $Y2=0
cc_173 N_A_M1018_g N_A_27_109#_c_213_n 0.0276911f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_174 A N_A_27_109#_c_213_n 0.00204487f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A_c_175_n N_A_27_109#_c_213_n 0.00787258f $X=0.67 $Y=1.68 $X2=0 $Y2=0
cc_176 N_A_M1018_g N_A_27_109#_M1020_g 0.0153827f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_177 N_A_M1004_g N_A_27_109#_c_216_n 0.0158051f $X=0.495 $Y=0.755 $X2=0 $Y2=0
cc_178 N_A_M1018_g N_A_27_109#_c_216_n 0.00215172f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_179 N_A_M1024_g N_A_27_109#_c_236_n 0.0143689f $X=0.67 $Y=2.545 $X2=0 $Y2=0
cc_180 N_A_M1004_g N_A_27_109#_c_217_n 0.0112534f $X=0.495 $Y=0.755 $X2=0 $Y2=0
cc_181 N_A_M1018_g N_A_27_109#_c_217_n 0.0161382f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_182 A N_A_27_109#_c_217_n 0.0260347f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A_c_175_n N_A_27_109#_c_217_n 7.85225e-19 $X=0.67 $Y=1.68 $X2=0 $Y2=0
cc_184 N_A_M1018_g N_A_27_109#_c_218_n 0.00112248f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_185 N_A_M1004_g N_A_27_109#_c_231_n 0.00505699f $X=0.495 $Y=0.755 $X2=0 $Y2=0
cc_186 N_A_M1024_g N_A_27_109#_c_237_n 0.00462278f $X=0.67 $Y=2.545 $X2=0 $Y2=0
cc_187 A N_A_27_109#_c_237_n 0.0082919f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A_c_175_n N_A_27_109#_c_237_n 0.00432057f $X=0.67 $Y=1.68 $X2=0 $Y2=0
cc_189 N_A_M1004_g N_A_27_109#_c_232_n 0.0128246f $X=0.495 $Y=0.755 $X2=0 $Y2=0
cc_190 N_A_M1024_g N_A_27_109#_c_232_n 0.00427061f $X=0.67 $Y=2.545 $X2=0 $Y2=0
cc_191 A N_A_27_109#_c_232_n 0.0239283f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A_M1018_g N_A_27_109#_c_233_n 0.00179482f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_193 A N_A_27_109#_c_233_n 0.0146256f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A_c_175_n N_A_27_109#_c_233_n 2.02996e-19 $X=0.67 $Y=1.68 $X2=0 $Y2=0
cc_195 N_A_M1024_g N_VPWR_c_841_n 0.0237187f $X=0.67 $Y=2.545 $X2=0 $Y2=0
cc_196 A N_VPWR_c_841_n 0.00522718f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A_c_175_n N_VPWR_c_841_n 0.00396253f $X=0.67 $Y=1.68 $X2=0 $Y2=0
cc_198 N_A_M1024_g N_VPWR_c_844_n 0.00769046f $X=0.67 $Y=2.545 $X2=0 $Y2=0
cc_199 N_A_M1024_g N_VPWR_c_840_n 0.0141493f $X=0.67 $Y=2.545 $X2=0 $Y2=0
cc_200 N_A_M1004_g N_VGND_c_1208_n 0.00180891f $X=0.495 $Y=0.755 $X2=0 $Y2=0
cc_201 N_A_M1018_g N_VGND_c_1208_n 0.0117171f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_202 N_A_M1004_g N_VGND_c_1211_n 0.00441768f $X=0.495 $Y=0.755 $X2=0 $Y2=0
cc_203 N_A_M1018_g N_VGND_c_1211_n 0.00382362f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_204 N_A_M1004_g N_VGND_c_1218_n 0.00492109f $X=0.495 $Y=0.755 $X2=0 $Y2=0
cc_205 N_A_M1018_g N_VGND_c_1218_n 0.00413371f $X=0.855 $Y=0.755 $X2=0 $Y2=0
cc_206 N_A_27_109#_c_225_n N_A_647_367#_c_369_n 0.0018199f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_207 N_A_27_109#_c_228_n N_A_647_367#_c_369_n 0.00494253f $X=4.425 $Y=0.98
+ $X2=0 $Y2=0
cc_208 N_A_27_109#_c_230_n N_A_647_367#_c_369_n 0.00449437f $X=5.795 $Y=0.7
+ $X2=0 $Y2=0
cc_209 N_A_27_109#_c_234_n N_A_647_367#_c_369_n 9.91946e-19 $X=4.51 $Y=0.7 $X2=0
+ $Y2=0
cc_210 N_A_27_109#_c_225_n N_A_647_367#_c_370_n 0.00359071f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_211 N_A_27_109#_c_228_n N_A_647_367#_c_371_n 0.0149132f $X=4.425 $Y=0.98
+ $X2=0 $Y2=0
cc_212 N_A_27_109#_c_230_n N_A_647_367#_M1008_g 0.0100476f $X=5.795 $Y=0.7 $X2=0
+ $Y2=0
cc_213 N_A_27_109#_c_234_n N_A_647_367#_M1008_g 0.00124462f $X=4.51 $Y=0.7 $X2=0
+ $Y2=0
cc_214 N_A_27_109#_c_271_p N_A_647_367#_c_374_n 0.00347468f $X=5.96 $Y=0.805
+ $X2=0 $Y2=0
cc_215 N_A_27_109#_c_271_p N_A_647_367#_M1006_g 0.0134402f $X=5.96 $Y=0.805
+ $X2=0 $Y2=0
cc_216 N_A_27_109#_c_230_n N_A_647_367#_M1023_g 0.0125813f $X=5.795 $Y=0.7 $X2=0
+ $Y2=0
cc_217 N_A_27_109#_c_271_p N_A_647_367#_M1023_g 0.0101102f $X=5.96 $Y=0.805
+ $X2=0 $Y2=0
cc_218 N_A_27_109#_c_234_n N_A_647_367#_c_377_n 6.71745e-19 $X=4.51 $Y=0.7 $X2=0
+ $Y2=0
cc_219 N_A_27_109#_c_222_n N_A_647_367#_c_378_n 0.012284f $X=2.905 $Y=1.08 $X2=0
+ $Y2=0
cc_220 N_A_27_109#_c_224_n N_A_647_367#_c_378_n 0.0044319f $X=2.99 $Y=0.995
+ $X2=0 $Y2=0
cc_221 N_A_27_109#_c_225_n N_A_647_367#_c_378_n 0.0182051f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_222 N_A_27_109#_c_227_n N_A_647_367#_c_378_n 0.0193562f $X=3.81 $Y=0.895
+ $X2=0 $Y2=0
cc_223 N_A_27_109#_c_229_n N_A_647_367#_c_378_n 0.0133652f $X=3.895 $Y=0.98
+ $X2=0 $Y2=0
cc_224 N_A_27_109#_c_229_n N_A_647_367#_c_380_n 0.00800389f $X=3.895 $Y=0.98
+ $X2=0 $Y2=0
cc_225 N_A_27_109#_c_225_n N_A_647_367#_c_382_n 0.00571747f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_226 N_A_27_109#_c_227_n N_A_647_367#_c_382_n 0.0160646f $X=3.81 $Y=0.895
+ $X2=0 $Y2=0
cc_227 N_A_27_109#_c_229_n N_A_647_367#_c_382_n 0.00817912f $X=3.895 $Y=0.98
+ $X2=0 $Y2=0
cc_228 N_A_27_109#_c_234_n N_A_647_367#_c_382_n 0.00134701f $X=4.51 $Y=0.7 $X2=0
+ $Y2=0
cc_229 N_A_27_109#_c_219_n N_B_M1012_g 2.90321e-19 $X=2.125 $Y=0.35 $X2=0 $Y2=0
cc_230 N_A_27_109#_c_221_n N_B_M1012_g 0.00351756f $X=2.21 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_27_109#_c_222_n N_B_M1012_g 0.0154318f $X=2.905 $Y=1.08 $X2=0 $Y2=0
cc_232 N_A_27_109#_c_224_n N_B_M1012_g 0.00281342f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_27_109#_c_226_n N_B_M1012_g 4.64707e-19 $X=3.075 $Y=0.35 $X2=0 $Y2=0
cc_234 N_A_27_109#_c_222_n N_B_M1021_g 0.00158375f $X=2.905 $Y=1.08 $X2=0 $Y2=0
cc_235 N_A_27_109#_c_224_n N_B_M1021_g 0.00312941f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_27_109#_c_225_n N_B_M1021_g 0.0113243f $X=3.725 $Y=0.35 $X2=0 $Y2=0
cc_237 N_A_27_109#_c_227_n N_B_M1021_g 7.14965e-19 $X=3.81 $Y=0.895 $X2=0 $Y2=0
cc_238 N_A_27_109#_c_230_n N_B_M1026_g 0.0125223f $X=5.795 $Y=0.7 $X2=0 $Y2=0
cc_239 N_A_27_109#_c_271_p N_B_M1026_g 9.20918e-19 $X=5.96 $Y=0.805 $X2=0 $Y2=0
cc_240 N_A_27_109#_c_230_n N_B_M1025_g 0.0021353f $X=5.795 $Y=0.7 $X2=0 $Y2=0
cc_241 N_A_27_109#_c_271_p N_B_M1025_g 0.0138149f $X=5.96 $Y=0.805 $X2=0 $Y2=0
cc_242 N_A_27_109#_c_271_p N_B_c_477_n 0.00348048f $X=5.96 $Y=0.805 $X2=0 $Y2=0
cc_243 N_A_27_109#_c_271_p N_B_M1016_g 0.00681903f $X=5.96 $Y=0.805 $X2=0 $Y2=0
cc_244 N_A_27_109#_c_213_n N_B_c_479_n 0.00240723f $X=1.2 $Y=2.03 $X2=0 $Y2=0
cc_245 N_A_27_109#_c_222_n N_B_c_479_n 0.0562636f $X=2.905 $Y=1.08 $X2=0 $Y2=0
cc_246 N_A_27_109#_c_223_n N_B_c_479_n 0.0147321f $X=2.295 $Y=1.08 $X2=0 $Y2=0
cc_247 N_A_27_109#_c_222_n N_B_c_480_n 0.00144938f $X=2.905 $Y=1.08 $X2=0 $Y2=0
cc_248 N_A_27_109#_c_213_n N_VPWR_c_841_n 0.0242976f $X=1.2 $Y=2.03 $X2=0 $Y2=0
cc_249 N_A_27_109#_c_237_n N_VPWR_c_841_n 0.0702172f $X=0.405 $Y=2.19 $X2=0
+ $Y2=0
cc_250 N_A_27_109#_c_236_n N_VPWR_c_844_n 0.0304602f $X=0.405 $Y=2.9 $X2=0 $Y2=0
cc_251 N_A_27_109#_c_213_n N_VPWR_c_846_n 0.00769046f $X=1.2 $Y=2.03 $X2=0 $Y2=0
cc_252 N_A_27_109#_c_213_n N_VPWR_c_840_n 0.0143431f $X=1.2 $Y=2.03 $X2=0 $Y2=0
cc_253 N_A_27_109#_c_236_n N_VPWR_c_840_n 0.0174175f $X=0.405 $Y=2.9 $X2=0 $Y2=0
cc_254 N_A_27_109#_c_230_n N_A_265_409#_M1008_d 0.00267852f $X=5.795 $Y=0.7
+ $X2=0 $Y2=0
cc_255 N_A_27_109#_c_213_n N_A_265_409#_c_908_n 0.0115307f $X=1.2 $Y=2.03 $X2=0
+ $Y2=0
cc_256 N_A_27_109#_c_213_n N_A_265_409#_c_905_n 0.0286691f $X=1.2 $Y=2.03 $X2=0
+ $Y2=0
cc_257 N_A_27_109#_M1015_g N_A_265_409#_c_905_n 0.00493988f $X=1.645 $Y=0.755
+ $X2=0 $Y2=0
cc_258 N_A_27_109#_c_221_n N_A_265_409#_c_905_n 5.042e-19 $X=2.21 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_27_109#_c_223_n N_A_265_409#_c_905_n 0.0106659f $X=2.295 $Y=1.08
+ $X2=0 $Y2=0
cc_260 N_A_27_109#_c_233_n N_A_265_409#_c_905_n 0.0444677f $X=1.34 $Y=1.33 $X2=0
+ $Y2=0
cc_261 N_A_27_109#_c_228_n N_A_265_409#_c_906_n 0.00159498f $X=4.425 $Y=0.98
+ $X2=0 $Y2=0
cc_262 N_A_27_109#_c_230_n N_A_265_409#_c_906_n 0.0256459f $X=5.795 $Y=0.7 $X2=0
+ $Y2=0
cc_263 N_A_27_109#_c_234_n N_A_265_409#_c_906_n 0.0143392f $X=4.51 $Y=0.7 $X2=0
+ $Y2=0
cc_264 N_A_27_109#_c_213_n N_A_265_409#_c_912_n 0.0172295f $X=1.2 $Y=2.03 $X2=0
+ $Y2=0
cc_265 N_A_27_109#_c_233_n N_A_265_409#_c_912_n 0.0158286f $X=1.34 $Y=1.33 $X2=0
+ $Y2=0
cc_266 N_A_27_109#_M1020_g N_A_265_409#_c_907_n 4.44532e-19 $X=1.285 $Y=0.755
+ $X2=0 $Y2=0
cc_267 N_A_27_109#_M1015_g N_A_265_409#_c_907_n 0.00455537f $X=1.645 $Y=0.755
+ $X2=0 $Y2=0
cc_268 N_A_27_109#_c_218_n N_A_265_409#_c_907_n 0.0363139f $X=1.42 $Y=1.165
+ $X2=0 $Y2=0
cc_269 N_A_27_109#_c_219_n N_A_265_409#_c_907_n 0.0157586f $X=2.125 $Y=0.35
+ $X2=0 $Y2=0
cc_270 N_A_27_109#_c_221_n N_A_265_409#_c_907_n 0.0270531f $X=2.21 $Y=0.995
+ $X2=0 $Y2=0
cc_271 N_A_27_109#_c_230_n N_A_763_347#_M1026_d 0.00433523f $X=5.795 $Y=0.7
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_27_109#_c_271_p N_A_763_347#_c_987_n 0.0129889f $X=5.96 $Y=0.805
+ $X2=0 $Y2=0
cc_273 N_A_27_109#_c_230_n N_A_763_347#_c_972_n 0.0208821f $X=5.795 $Y=0.7 $X2=0
+ $Y2=0
cc_274 N_A_27_109#_c_271_p N_A_763_347#_c_972_n 0.0601696f $X=5.96 $Y=0.805
+ $X2=0 $Y2=0
cc_275 N_A_27_109#_c_228_n N_A_803_81#_M1008_s 0.0150303f $X=4.425 $Y=0.98
+ $X2=-0.19 $Y2=-0.245
cc_276 N_A_27_109#_c_234_n N_A_803_81#_M1008_s 0.00529656f $X=4.51 $Y=0.7
+ $X2=-0.19 $Y2=-0.245
cc_277 N_A_27_109#_c_227_n N_A_803_81#_c_1112_n 0.0198003f $X=3.81 $Y=0.895
+ $X2=0 $Y2=0
cc_278 N_A_27_109#_c_228_n N_A_803_81#_c_1112_n 0.0126671f $X=4.425 $Y=0.98
+ $X2=0 $Y2=0
cc_279 N_A_27_109#_c_234_n N_A_803_81#_c_1112_n 0.00709693f $X=4.51 $Y=0.7 $X2=0
+ $Y2=0
cc_280 N_A_27_109#_c_228_n N_A_803_81#_c_1105_n 0.00628123f $X=4.425 $Y=0.98
+ $X2=0 $Y2=0
cc_281 N_A_27_109#_c_230_n N_A_803_81#_c_1105_n 0.0981496f $X=5.795 $Y=0.7 $X2=0
+ $Y2=0
cc_282 N_A_27_109#_c_234_n N_A_803_81#_c_1105_n 0.0122952f $X=4.51 $Y=0.7 $X2=0
+ $Y2=0
cc_283 N_A_27_109#_c_225_n N_A_803_81#_c_1106_n 0.0146441f $X=3.725 $Y=0.35
+ $X2=0 $Y2=0
cc_284 N_A_27_109#_M1006_d N_A_803_81#_c_1119_n 0.0050656f $X=5.82 $Y=1.735
+ $X2=0 $Y2=0
cc_285 N_A_27_109#_c_271_p N_A_803_81#_c_1119_n 0.0156953f $X=5.96 $Y=0.805
+ $X2=0 $Y2=0
cc_286 N_A_27_109#_c_271_p N_A_803_81#_c_1107_n 0.0761782f $X=5.96 $Y=0.805
+ $X2=0 $Y2=0
cc_287 N_A_27_109#_M1020_g N_VGND_c_1208_n 0.00123075f $X=1.285 $Y=0.755 $X2=0
+ $Y2=0
cc_288 N_A_27_109#_c_216_n N_VGND_c_1208_n 0.0150699f $X=0.28 $Y=0.755 $X2=0
+ $Y2=0
cc_289 N_A_27_109#_c_217_n N_VGND_c_1208_n 0.0199134f $X=1.175 $Y=1.25 $X2=0
+ $Y2=0
cc_290 N_A_27_109#_c_218_n N_VGND_c_1208_n 0.0226764f $X=1.42 $Y=1.165 $X2=0
+ $Y2=0
cc_291 N_A_27_109#_c_220_n N_VGND_c_1208_n 0.014068f $X=1.505 $Y=0.35 $X2=0
+ $Y2=0
cc_292 N_A_27_109#_c_219_n N_VGND_c_1209_n 0.0141599f $X=2.125 $Y=0.35 $X2=0
+ $Y2=0
cc_293 N_A_27_109#_c_221_n N_VGND_c_1209_n 0.0278208f $X=2.21 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_27_109#_c_222_n N_VGND_c_1209_n 0.0170197f $X=2.905 $Y=1.08 $X2=0
+ $Y2=0
cc_295 N_A_27_109#_c_224_n N_VGND_c_1209_n 0.0155096f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_27_109#_c_226_n N_VGND_c_1209_n 0.0139184f $X=3.075 $Y=0.35 $X2=0
+ $Y2=0
cc_297 N_A_27_109#_c_216_n N_VGND_c_1211_n 0.00845426f $X=0.28 $Y=0.755 $X2=0
+ $Y2=0
cc_298 N_A_27_109#_c_225_n N_VGND_c_1214_n 0.0500748f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_299 N_A_27_109#_c_226_n N_VGND_c_1214_n 0.0114622f $X=3.075 $Y=0.35 $X2=0
+ $Y2=0
cc_300 N_A_27_109#_M1020_g N_VGND_c_1216_n 0.00394144f $X=1.285 $Y=0.755 $X2=0
+ $Y2=0
cc_301 N_A_27_109#_M1015_g N_VGND_c_1216_n 6.46133e-19 $X=1.645 $Y=0.755 $X2=0
+ $Y2=0
cc_302 N_A_27_109#_c_219_n N_VGND_c_1216_n 0.049001f $X=2.125 $Y=0.35 $X2=0
+ $Y2=0
cc_303 N_A_27_109#_c_220_n N_VGND_c_1216_n 0.0114622f $X=1.505 $Y=0.35 $X2=0
+ $Y2=0
cc_304 N_A_27_109#_M1020_g N_VGND_c_1218_n 0.00410091f $X=1.285 $Y=0.755 $X2=0
+ $Y2=0
cc_305 N_A_27_109#_c_216_n N_VGND_c_1218_n 0.0107549f $X=0.28 $Y=0.755 $X2=0
+ $Y2=0
cc_306 N_A_27_109#_c_219_n N_VGND_c_1218_n 0.0297409f $X=2.125 $Y=0.35 $X2=0
+ $Y2=0
cc_307 N_A_27_109#_c_220_n N_VGND_c_1218_n 0.00657784f $X=1.505 $Y=0.35 $X2=0
+ $Y2=0
cc_308 N_A_27_109#_c_225_n N_VGND_c_1218_n 0.0298395f $X=3.725 $Y=0.35 $X2=0
+ $Y2=0
cc_309 N_A_27_109#_c_226_n N_VGND_c_1218_n 0.00657784f $X=3.075 $Y=0.35 $X2=0
+ $Y2=0
cc_310 N_A_27_109#_c_218_n A_272_109# 0.00389086f $X=1.42 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_311 N_A_27_109#_c_224_n A_570_101# 0.00144497f $X=2.99 $Y=0.995 $X2=-0.19
+ $Y2=-0.245
cc_312 N_A_647_367#_c_388_n N_B_M1003_g 0.0129649f $X=3.375 $Y=1.98 $X2=0 $Y2=0
cc_313 N_A_647_367#_c_379_n N_B_M1003_g 0.00418166f $X=3.375 $Y=1.815 $X2=0
+ $Y2=0
cc_314 N_A_647_367#_c_378_n N_B_M1021_g 0.00652888f $X=3.46 $Y=0.78 $X2=0 $Y2=0
cc_315 N_A_647_367#_c_380_n N_B_M1021_g 0.00538555f $X=3.665 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A_647_367#_c_381_n N_B_M1021_g 0.0156391f $X=3.665 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A_647_367#_c_382_n N_B_M1021_g 0.0169208f $X=3.665 $Y=1.245 $X2=0 $Y2=0
cc_318 N_A_647_367#_M1011_g N_B_c_482_n 0.0146975f $X=4.305 $Y=2.235 $X2=0 $Y2=0
cc_319 N_A_647_367#_M1006_g N_B_M1014_g 0.0384304f $X=5.695 $Y=2.235 $X2=0 $Y2=0
cc_320 N_A_647_367#_c_369_n N_B_M1026_g 0.00584781f $X=5.67 $Y=0.255 $X2=0 $Y2=0
cc_321 N_A_647_367#_M1008_g N_B_M1026_g 0.0208434f $X=4.725 $Y=0.985 $X2=0 $Y2=0
cc_322 N_A_647_367#_c_374_n N_B_M1026_g 0.00964594f $X=5.695 $Y=1.395 $X2=0
+ $Y2=0
cc_323 N_A_647_367#_M1023_g N_B_M1026_g 0.0140914f $X=5.745 $Y=0.765 $X2=0 $Y2=0
cc_324 N_A_647_367#_M1006_g N_B_c_486_n 0.0146975f $X=5.695 $Y=2.235 $X2=0 $Y2=0
cc_325 N_A_647_367#_M1023_g N_B_M1025_g 0.0268752f $X=5.745 $Y=0.765 $X2=0 $Y2=0
cc_326 N_A_647_367#_c_374_n N_B_c_477_n 0.0268752f $X=5.695 $Y=1.395 $X2=0 $Y2=0
cc_327 N_A_647_367#_M1006_g N_B_M1016_g 0.0268752f $X=5.695 $Y=2.235 $X2=0 $Y2=0
cc_328 N_A_647_367#_M1011_g N_B_c_478_n 0.0122963f $X=4.305 $Y=2.235 $X2=0 $Y2=0
cc_329 N_A_647_367#_c_372_n N_B_c_478_n 0.00376957f $X=4.65 $Y=1.5 $X2=0 $Y2=0
cc_330 N_A_647_367#_M1006_g N_B_c_478_n 0.00964594f $X=5.695 $Y=2.235 $X2=0
+ $Y2=0
cc_331 N_A_647_367#_c_379_n N_B_c_479_n 0.0119536f $X=3.375 $Y=1.815 $X2=0 $Y2=0
cc_332 N_A_647_367#_c_380_n N_B_c_479_n 0.0142731f $X=3.665 $Y=1.41 $X2=0 $Y2=0
cc_333 N_A_647_367#_c_388_n N_B_c_480_n 2.23129e-19 $X=3.375 $Y=1.98 $X2=0 $Y2=0
cc_334 N_A_647_367#_c_379_n N_B_c_480_n 0.00301458f $X=3.375 $Y=1.815 $X2=0
+ $Y2=0
cc_335 N_A_647_367#_M1003_d N_A_265_409#_c_910_n 0.00809794f $X=3.235 $Y=1.835
+ $X2=0 $Y2=0
cc_336 N_A_647_367#_M1011_g N_A_265_409#_c_910_n 0.0344536f $X=4.305 $Y=2.235
+ $X2=0 $Y2=0
cc_337 N_A_647_367#_c_388_n N_A_265_409#_c_910_n 0.0203736f $X=3.375 $Y=1.98
+ $X2=0 $Y2=0
cc_338 N_A_647_367#_c_380_n N_A_265_409#_c_910_n 0.00766273f $X=3.665 $Y=1.41
+ $X2=0 $Y2=0
cc_339 N_A_647_367#_c_381_n N_A_265_409#_c_910_n 0.0118082f $X=3.665 $Y=1.41
+ $X2=0 $Y2=0
cc_340 N_A_647_367#_M1008_g N_A_265_409#_c_906_n 0.023305f $X=4.725 $Y=0.985
+ $X2=0 $Y2=0
cc_341 N_A_647_367#_c_380_n N_A_265_409#_c_906_n 0.00590187f $X=3.665 $Y=1.41
+ $X2=0 $Y2=0
cc_342 N_A_647_367#_c_381_n N_A_265_409#_c_906_n 5.676e-19 $X=3.665 $Y=1.41
+ $X2=0 $Y2=0
cc_343 N_A_647_367#_M1011_g N_A_265_409#_c_911_n 0.0350338f $X=4.305 $Y=2.235
+ $X2=0 $Y2=0
cc_344 N_A_647_367#_c_372_n N_A_265_409#_c_911_n 0.0161542f $X=4.65 $Y=1.5 $X2=0
+ $Y2=0
cc_345 N_A_647_367#_M1008_g N_A_265_409#_c_911_n 3.31555e-19 $X=4.725 $Y=0.985
+ $X2=0 $Y2=0
cc_346 N_A_647_367#_c_377_n N_A_265_409#_c_911_n 0.00477776f $X=4.305 $Y=1.5
+ $X2=0 $Y2=0
cc_347 N_A_647_367#_c_380_n N_A_265_409#_c_911_n 0.00457107f $X=3.665 $Y=1.41
+ $X2=0 $Y2=0
cc_348 N_A_647_367#_M1011_g N_A_763_347#_c_975_n 0.00291876f $X=4.305 $Y=2.235
+ $X2=0 $Y2=0
cc_349 N_A_647_367#_M1011_g N_A_763_347#_c_976_n 0.00358298f $X=4.305 $Y=2.235
+ $X2=0 $Y2=0
cc_350 N_A_647_367#_M1006_g N_A_763_347#_c_976_n 0.00168418f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_351 N_A_647_367#_M1006_g N_A_763_347#_c_987_n 0.00579674f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_352 N_A_647_367#_M1006_g N_A_763_347#_c_977_n 0.00316661f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_353 N_A_647_367#_M1008_g N_A_763_347#_c_972_n 7.761e-19 $X=4.725 $Y=0.985
+ $X2=0 $Y2=0
cc_354 N_A_647_367#_c_374_n N_A_763_347#_c_972_n 0.00450774f $X=5.695 $Y=1.395
+ $X2=0 $Y2=0
cc_355 N_A_647_367#_M1006_g N_A_763_347#_c_972_n 0.0116201f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_356 N_A_647_367#_M1023_g N_A_763_347#_c_972_n 0.00259295f $X=5.745 $Y=0.765
+ $X2=0 $Y2=0
cc_357 N_A_647_367#_M1006_g N_A_763_347#_c_978_n 0.00154888f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_358 N_A_647_367#_M1011_g N_A_763_347#_c_983_n 0.00876487f $X=4.305 $Y=2.235
+ $X2=0 $Y2=0
cc_359 N_A_647_367#_c_382_n N_A_803_81#_c_1112_n 0.00167942f $X=3.665 $Y=1.245
+ $X2=0 $Y2=0
cc_360 N_A_647_367#_c_369_n N_A_803_81#_c_1105_n 0.0413428f $X=5.67 $Y=0.255
+ $X2=0 $Y2=0
cc_361 N_A_647_367#_M1008_g N_A_803_81#_c_1105_n 4.54389e-19 $X=4.725 $Y=0.985
+ $X2=0 $Y2=0
cc_362 N_A_647_367#_M1023_g N_A_803_81#_c_1105_n 0.00837143f $X=5.745 $Y=0.765
+ $X2=0 $Y2=0
cc_363 N_A_647_367#_c_369_n N_A_803_81#_c_1106_n 0.00679683f $X=5.67 $Y=0.255
+ $X2=0 $Y2=0
cc_364 N_A_647_367#_M1006_g N_A_803_81#_c_1127_n 0.00915648f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_365 N_A_647_367#_M1006_g N_A_803_81#_c_1119_n 0.0195966f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_366 N_A_647_367#_M1006_g N_A_803_81#_c_1129_n 0.00200935f $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_367 N_A_647_367#_M1006_g N_A_803_81#_c_1107_n 8.13044e-19 $X=5.695 $Y=2.235
+ $X2=0 $Y2=0
cc_368 N_A_647_367#_c_370_n N_VGND_c_1214_n 0.0415614f $X=3.83 $Y=0.255 $X2=0
+ $Y2=0
cc_369 N_A_647_367#_c_369_n N_VGND_c_1218_n 0.0549621f $X=5.67 $Y=0.255 $X2=0
+ $Y2=0
cc_370 N_A_647_367#_c_370_n N_VGND_c_1218_n 0.00488025f $X=3.83 $Y=0.255 $X2=0
+ $Y2=0
cc_371 N_B_M1025_g N_A_1318_85#_M1002_g 0.0237847f $X=6.175 $Y=0.765 $X2=0 $Y2=0
cc_372 N_B_c_477_n N_A_1318_85#_M1007_g 0.0228926f $X=6.225 $Y=1.635 $X2=0 $Y2=0
cc_373 N_B_M1016_g N_A_1318_85#_c_601_n 0.0228926f $X=6.225 $Y=2.235 $X2=0 $Y2=0
cc_374 N_B_c_477_n N_A_1318_85#_c_595_n 0.0042088f $X=6.225 $Y=1.635 $X2=0 $Y2=0
cc_375 N_B_M1016_g N_A_1348_111#_c_770_n 3.47477e-19 $X=6.225 $Y=2.235 $X2=0
+ $Y2=0
cc_376 N_B_M1003_g N_VPWR_c_842_n 0.0216221f $X=3.11 $Y=2.335 $X2=0 $Y2=0
cc_377 N_B_c_483_n N_VPWR_c_847_n 0.0840857f $X=3.235 $Y=3.15 $X2=0 $Y2=0
cc_378 N_B_c_482_n N_VPWR_c_840_n 0.0602437f $X=5.04 $Y=3.15 $X2=0 $Y2=0
cc_379 N_B_c_483_n N_VPWR_c_840_n 0.017662f $X=3.235 $Y=3.15 $X2=0 $Y2=0
cc_380 N_B_c_486_n N_VPWR_c_840_n 0.0290557f $X=6.1 $Y=3.15 $X2=0 $Y2=0
cc_381 N_B_c_491_n N_VPWR_c_840_n 0.00371008f $X=5.115 $Y=3.15 $X2=0 $Y2=0
cc_382 N_B_c_479_n N_A_265_409#_c_905_n 0.0351159f $X=2.865 $Y=1.51 $X2=0 $Y2=0
cc_383 N_B_M1003_g N_A_265_409#_c_910_n 0.0326334f $X=3.11 $Y=2.335 $X2=0 $Y2=0
cc_384 N_B_c_482_n N_A_265_409#_c_910_n 0.0100514f $X=5.04 $Y=3.15 $X2=0 $Y2=0
cc_385 N_B_M1014_g N_A_265_409#_c_910_n 0.00159308f $X=5.165 $Y=2.235 $X2=0
+ $Y2=0
cc_386 N_B_c_479_n N_A_265_409#_c_910_n 0.0379259f $X=2.865 $Y=1.51 $X2=0 $Y2=0
cc_387 N_B_c_480_n N_A_265_409#_c_910_n 0.00117243f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_388 N_B_M1026_g N_A_265_409#_c_906_n 0.00321291f $X=5.235 $Y=0.985 $X2=0
+ $Y2=0
cc_389 N_B_c_478_n N_A_265_409#_c_906_n 0.00212932f $X=5.175 $Y=1.66 $X2=0 $Y2=0
cc_390 N_B_M1014_g N_A_265_409#_c_911_n 0.00146039f $X=5.165 $Y=2.235 $X2=0
+ $Y2=0
cc_391 N_B_M1026_g N_A_265_409#_c_911_n 3.17402e-19 $X=5.235 $Y=0.985 $X2=0
+ $Y2=0
cc_392 N_B_c_478_n N_A_265_409#_c_911_n 0.00271404f $X=5.175 $Y=1.66 $X2=0 $Y2=0
cc_393 N_B_c_482_n N_A_763_347#_c_975_n 0.0143091f $X=5.04 $Y=3.15 $X2=0 $Y2=0
cc_394 N_B_M1014_g N_A_763_347#_c_976_n 0.023692f $X=5.165 $Y=2.235 $X2=0 $Y2=0
cc_395 N_B_c_485_n N_A_763_347#_c_976_n 0.00164607f $X=5.115 $Y=3.075 $X2=0
+ $Y2=0
cc_396 N_B_c_490_n N_A_763_347#_c_976_n 0.00411549f $X=5.165 $Y=2.865 $X2=0
+ $Y2=0
cc_397 N_B_M1014_g N_A_763_347#_c_987_n 0.0214007f $X=5.165 $Y=2.235 $X2=0 $Y2=0
cc_398 N_B_M1014_g N_A_763_347#_c_1006_n 0.00360135f $X=5.165 $Y=2.235 $X2=0
+ $Y2=0
cc_399 N_B_c_485_n N_A_763_347#_c_977_n 0.0112351f $X=5.115 $Y=3.075 $X2=0 $Y2=0
cc_400 N_B_c_486_n N_A_763_347#_c_977_n 0.0127455f $X=6.1 $Y=3.15 $X2=0 $Y2=0
cc_401 N_B_M1016_g N_A_763_347#_c_977_n 0.0156022f $X=6.225 $Y=2.235 $X2=0 $Y2=0
cc_402 N_B_c_490_n N_A_763_347#_c_977_n 0.00419299f $X=5.165 $Y=2.865 $X2=0
+ $Y2=0
cc_403 N_B_M1014_g N_A_763_347#_c_972_n 0.00430917f $X=5.165 $Y=2.235 $X2=0
+ $Y2=0
cc_404 N_B_M1026_g N_A_763_347#_c_972_n 0.0102897f $X=5.235 $Y=0.985 $X2=0 $Y2=0
cc_405 N_B_M1025_g N_A_763_347#_c_972_n 2.9708e-19 $X=6.175 $Y=0.765 $X2=0 $Y2=0
cc_406 N_B_c_478_n N_A_763_347#_c_972_n 0.0053098f $X=5.175 $Y=1.66 $X2=0 $Y2=0
cc_407 N_B_M1016_g N_A_763_347#_c_978_n 0.010873f $X=6.225 $Y=2.235 $X2=0 $Y2=0
cc_408 N_B_M1003_g N_A_763_347#_c_983_n 0.0122651f $X=3.11 $Y=2.335 $X2=0 $Y2=0
cc_409 N_B_c_482_n N_A_763_347#_c_983_n 0.00794352f $X=5.04 $Y=3.15 $X2=0 $Y2=0
cc_410 N_B_c_482_n N_A_763_347#_c_984_n 8.6217e-19 $X=5.04 $Y=3.15 $X2=0 $Y2=0
cc_411 N_B_c_485_n N_A_763_347#_c_984_n 0.00521259f $X=5.115 $Y=3.075 $X2=0
+ $Y2=0
cc_412 N_B_M1016_g N_A_763_347#_c_985_n 0.00305274f $X=6.225 $Y=2.235 $X2=0
+ $Y2=0
cc_413 N_B_M1026_g N_A_803_81#_c_1105_n 4.54389e-19 $X=5.235 $Y=0.985 $X2=0
+ $Y2=0
cc_414 N_B_M1025_g N_A_803_81#_c_1105_n 0.00883889f $X=6.175 $Y=0.765 $X2=0
+ $Y2=0
cc_415 N_B_M1014_g N_A_803_81#_c_1127_n 0.00773366f $X=5.165 $Y=2.235 $X2=0
+ $Y2=0
cc_416 N_B_M1016_g N_A_803_81#_c_1127_n 0.00167569f $X=6.225 $Y=2.235 $X2=0
+ $Y2=0
cc_417 N_B_M1016_g N_A_803_81#_c_1119_n 0.018851f $X=6.225 $Y=2.235 $X2=0 $Y2=0
cc_418 N_B_M1014_g N_A_803_81#_c_1129_n 0.00443852f $X=5.165 $Y=2.235 $X2=0
+ $Y2=0
cc_419 N_B_M1025_g N_A_803_81#_c_1107_n 0.00729079f $X=6.175 $Y=0.765 $X2=0
+ $Y2=0
cc_420 N_B_c_477_n N_A_803_81#_c_1107_n 0.00414138f $X=6.225 $Y=1.635 $X2=0
+ $Y2=0
cc_421 N_B_M1016_g N_A_803_81#_c_1107_n 0.0140321f $X=6.225 $Y=2.235 $X2=0 $Y2=0
cc_422 N_B_M1016_g N_A_803_81#_c_1140_n 0.00405141f $X=6.225 $Y=2.235 $X2=0
+ $Y2=0
cc_423 N_B_M1016_g N_A_803_81#_c_1141_n 6.73389e-19 $X=6.225 $Y=2.235 $X2=0
+ $Y2=0
cc_424 N_B_M1012_g N_VGND_c_1209_n 0.00782186f $X=2.775 $Y=0.715 $X2=0 $Y2=0
cc_425 N_B_M1012_g N_VGND_c_1214_n 0.00402651f $X=2.775 $Y=0.715 $X2=0 $Y2=0
cc_426 N_B_M1021_g N_VGND_c_1214_n 7.10185e-19 $X=3.165 $Y=0.715 $X2=0 $Y2=0
cc_427 N_B_M1025_g N_VGND_c_1214_n 6.31558e-19 $X=6.175 $Y=0.765 $X2=0 $Y2=0
cc_428 N_B_M1012_g N_VGND_c_1218_n 0.00423264f $X=2.775 $Y=0.715 $X2=0 $Y2=0
cc_429 N_A_1318_85#_M1002_g N_C_c_683_n 0.0161346f $X=6.665 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_430 N_A_1318_85#_M1002_g N_C_M1022_g 0.00437032f $X=6.665 $Y=0.765 $X2=0
+ $Y2=0
cc_431 N_A_1318_85#_c_600_n N_C_M1022_g 0.0137569f $X=8.05 $Y=3.11 $X2=0 $Y2=0
cc_432 N_A_1318_85#_c_595_n N_C_M1022_g 0.0465369f $X=6.775 $Y=1.59 $X2=0 $Y2=0
cc_433 N_A_1318_85#_c_597_n N_C_M1022_g 2.52682e-19 $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_434 N_A_1318_85#_c_598_n N_C_M1022_g 0.0174072f $X=8.215 $Y=1.68 $X2=0 $Y2=0
cc_435 N_A_1318_85#_c_596_n N_C_c_686_n 0.0121863f $X=8.475 $Y=0.705 $X2=0 $Y2=0
cc_436 N_A_1318_85#_c_597_n N_C_c_686_n 0.00153623f $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_437 N_A_1318_85#_c_596_n N_C_c_687_n 0.00408401f $X=8.475 $Y=0.705 $X2=0
+ $Y2=0
cc_438 N_A_1318_85#_c_597_n N_C_c_687_n 0.00807686f $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_439 N_A_1318_85#_c_596_n N_C_c_688_n 0.00685048f $X=8.475 $Y=0.705 $X2=0
+ $Y2=0
cc_440 N_A_1318_85#_c_597_n N_C_c_688_n 0.00908074f $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_441 N_A_1318_85#_c_602_n N_C_M1000_g 0.0172274f $X=8.125 $Y=3.035 $X2=0 $Y2=0
cc_442 N_A_1318_85#_c_604_n N_C_M1000_g 0.0244589f $X=8.48 $Y=2.15 $X2=0 $Y2=0
cc_443 N_A_1318_85#_c_597_n N_C_M1000_g 0.0163991f $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_444 N_A_1318_85#_c_598_n N_C_M1000_g 0.0180153f $X=8.215 $Y=1.68 $X2=0 $Y2=0
cc_445 N_A_1318_85#_c_597_n N_C_c_690_n 0.00704409f $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_446 N_A_1318_85#_c_596_n N_C_c_691_n 0.0216234f $X=8.475 $Y=0.705 $X2=0 $Y2=0
cc_447 N_A_1318_85#_c_597_n N_C_c_691_n 0.0138905f $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_448 N_A_1318_85#_c_596_n N_C_c_692_n 4.56525e-19 $X=8.475 $Y=0.705 $X2=0
+ $Y2=0
cc_449 N_A_1318_85#_c_596_n N_C_c_693_n 0.00189048f $X=8.475 $Y=0.705 $X2=0
+ $Y2=0
cc_450 N_A_1318_85#_c_597_n N_C_c_693_n 0.00212142f $X=8.56 $Y=1.56 $X2=0 $Y2=0
cc_451 N_A_1318_85#_c_598_n N_C_c_693_n 0.0234443f $X=8.215 $Y=1.68 $X2=0 $Y2=0
cc_452 N_A_1318_85#_c_596_n N_A_1348_111#_M1001_g 5.78712e-19 $X=8.475 $Y=0.705
+ $X2=0 $Y2=0
cc_453 N_A_1318_85#_c_597_n N_A_1348_111#_M1001_g 0.00207149f $X=8.56 $Y=1.56
+ $X2=0 $Y2=0
cc_454 N_A_1318_85#_c_597_n N_A_1348_111#_c_759_n 9.94341e-19 $X=8.56 $Y=1.56
+ $X2=0 $Y2=0
cc_455 N_A_1318_85#_c_604_n N_A_1348_111#_M1013_g 0.00109644f $X=8.48 $Y=2.15
+ $X2=0 $Y2=0
cc_456 N_A_1318_85#_M1002_g N_A_1348_111#_c_763_n 0.0184621f $X=6.665 $Y=0.765
+ $X2=0 $Y2=0
cc_457 N_A_1318_85#_M1007_g N_A_1348_111#_c_763_n 0.00250149f $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_458 N_A_1318_85#_c_595_n N_A_1348_111#_c_763_n 0.010853f $X=6.775 $Y=1.59
+ $X2=0 $Y2=0
cc_459 N_A_1318_85#_M1002_g N_A_1348_111#_c_764_n 6.66015e-19 $X=6.665 $Y=0.765
+ $X2=0 $Y2=0
cc_460 N_A_1318_85#_M1007_g N_A_1348_111#_c_770_n 0.0139947f $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_461 N_A_1318_85#_c_596_n N_A_1348_111#_c_766_n 0.0587088f $X=8.475 $Y=0.705
+ $X2=0 $Y2=0
cc_462 N_A_1318_85#_c_600_n N_VPWR_c_843_n 6.74052e-19 $X=8.05 $Y=3.11 $X2=0
+ $Y2=0
cc_463 N_A_1318_85#_c_602_n N_VPWR_c_843_n 7.44632e-19 $X=8.125 $Y=3.035 $X2=0
+ $Y2=0
cc_464 N_A_1318_85#_c_604_n N_VPWR_c_843_n 0.0685263f $X=8.48 $Y=2.15 $X2=0
+ $Y2=0
cc_465 N_A_1318_85#_c_601_n N_VPWR_c_847_n 0.0318716f $X=6.96 $Y=3.11 $X2=0
+ $Y2=0
cc_466 N_A_1318_85#_c_604_n N_VPWR_c_847_n 0.0177662f $X=8.48 $Y=2.15 $X2=0
+ $Y2=0
cc_467 N_A_1318_85#_c_600_n N_VPWR_c_840_n 0.0360168f $X=8.05 $Y=3.11 $X2=0
+ $Y2=0
cc_468 N_A_1318_85#_c_601_n N_VPWR_c_840_n 0.00704774f $X=6.96 $Y=3.11 $X2=0
+ $Y2=0
cc_469 N_A_1318_85#_c_604_n N_VPWR_c_840_n 0.0123184f $X=8.48 $Y=2.15 $X2=0
+ $Y2=0
cc_470 N_A_1318_85#_M1007_g N_A_763_347#_c_978_n 0.00751311f $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_471 N_A_1318_85#_M1007_g N_A_763_347#_c_979_n 0.0146017f $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_472 N_A_1318_85#_c_600_n N_A_763_347#_c_979_n 0.0258575f $X=8.05 $Y=3.11
+ $X2=0 $Y2=0
cc_473 N_A_1318_85#_c_601_n N_A_763_347#_c_979_n 0.00313913f $X=6.96 $Y=3.11
+ $X2=0 $Y2=0
cc_474 N_A_1318_85#_c_602_n N_A_763_347#_c_979_n 0.00506013f $X=8.125 $Y=3.035
+ $X2=0 $Y2=0
cc_475 N_A_1318_85#_c_604_n N_A_763_347#_c_979_n 0.00816064f $X=8.48 $Y=2.15
+ $X2=0 $Y2=0
cc_476 N_A_1318_85#_M1002_g N_A_763_347#_c_973_n 2.91784e-19 $X=6.665 $Y=0.765
+ $X2=0 $Y2=0
cc_477 N_A_1318_85#_c_595_n N_A_763_347#_c_973_n 2.19152e-19 $X=6.775 $Y=1.59
+ $X2=0 $Y2=0
cc_478 N_A_1318_85#_c_597_n N_A_763_347#_c_973_n 0.0056778f $X=8.56 $Y=1.56
+ $X2=0 $Y2=0
cc_479 N_A_1318_85#_c_598_n N_A_763_347#_c_973_n 0.00120871f $X=8.215 $Y=1.68
+ $X2=0 $Y2=0
cc_480 N_A_1318_85#_c_602_n N_A_763_347#_c_981_n 0.00537854f $X=8.125 $Y=3.035
+ $X2=0 $Y2=0
cc_481 N_A_1318_85#_c_604_n N_A_763_347#_c_981_n 0.0106948f $X=8.48 $Y=2.15
+ $X2=0 $Y2=0
cc_482 N_A_1318_85#_c_597_n N_A_763_347#_c_981_n 0.00111603f $X=8.56 $Y=1.56
+ $X2=0 $Y2=0
cc_483 N_A_1318_85#_M1007_g N_A_763_347#_c_1034_n 7.94337e-19 $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_484 N_A_1318_85#_c_602_n N_A_763_347#_c_982_n 0.0185318f $X=8.125 $Y=3.035
+ $X2=0 $Y2=0
cc_485 N_A_1318_85#_c_604_n N_A_763_347#_c_982_n 0.0424623f $X=8.48 $Y=2.15
+ $X2=0 $Y2=0
cc_486 N_A_1318_85#_c_596_n N_A_763_347#_c_974_n 0.0153693f $X=8.475 $Y=0.705
+ $X2=0 $Y2=0
cc_487 N_A_1318_85#_M1002_g N_A_803_81#_c_1107_n 0.00900184f $X=6.665 $Y=0.765
+ $X2=0 $Y2=0
cc_488 N_A_1318_85#_M1007_g N_A_803_81#_c_1107_n 0.00627215f $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_489 N_A_1318_85#_M1007_g N_A_803_81#_c_1144_n 0.010085f $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_490 N_A_1318_85#_c_595_n N_A_803_81#_c_1144_n 0.00264559f $X=6.775 $Y=1.59
+ $X2=0 $Y2=0
cc_491 N_A_1318_85#_c_600_n N_A_803_81#_c_1146_n 9.01126e-19 $X=8.05 $Y=3.11
+ $X2=0 $Y2=0
cc_492 N_A_1318_85#_M1007_g N_A_803_81#_c_1141_n 0.0132477f $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_493 N_A_1318_85#_M1007_g N_A_803_81#_c_1109_n 8.22491e-19 $X=6.835 $Y=2.165
+ $X2=0 $Y2=0
cc_494 N_A_1318_85#_c_600_n N_A_803_81#_c_1109_n 0.00121909f $X=8.05 $Y=3.11
+ $X2=0 $Y2=0
cc_495 N_A_1318_85#_c_602_n N_A_803_81#_c_1109_n 0.00102712f $X=8.125 $Y=3.035
+ $X2=0 $Y2=0
cc_496 N_A_1318_85#_c_596_n N_VGND_c_1213_n 0.00472179f $X=8.475 $Y=0.705 $X2=0
+ $Y2=0
cc_497 N_A_1318_85#_c_597_n N_VGND_c_1213_n 0.0199209f $X=8.56 $Y=1.56 $X2=0
+ $Y2=0
cc_498 N_A_1318_85#_M1002_g N_VGND_c_1214_n 0.00388996f $X=6.665 $Y=0.765 $X2=0
+ $Y2=0
cc_499 N_A_1318_85#_M1002_g N_VGND_c_1218_n 0.00407676f $X=6.665 $Y=0.765 $X2=0
+ $Y2=0
cc_500 N_A_1318_85#_c_596_n A_1634_89# 0.00653524f $X=8.475 $Y=0.705 $X2=-0.19
+ $Y2=-0.245
cc_501 N_C_c_688_n N_A_1348_111#_M1001_g 0.00838724f $X=8.57 $Y=1.155 $X2=0
+ $Y2=0
cc_502 N_C_c_690_n N_A_1348_111#_M1001_g 0.0224286f $X=8.682 $Y=1.23 $X2=0 $Y2=0
cc_503 N_C_M1000_g N_A_1348_111#_c_759_n 0.0224286f $X=8.745 $Y=2.505 $X2=0
+ $Y2=0
cc_504 N_C_c_683_n N_A_1348_111#_c_763_n 0.00577913f $X=7.095 $Y=1.05 $X2=0
+ $Y2=0
cc_505 N_C_M1022_g N_A_1348_111#_c_763_n 0.00372482f $X=7.365 $Y=2.165 $X2=0
+ $Y2=0
cc_506 N_C_c_685_n N_A_1348_111#_c_770_n 0.00499286f $X=7.49 $Y=1.125 $X2=0
+ $Y2=0
cc_507 N_C_c_686_n N_A_1348_111#_c_765_n 4.75334e-19 $X=8.095 $Y=0.975 $X2=0
+ $Y2=0
cc_508 N_C_c_683_n N_A_1348_111#_c_766_n 0.00896313f $X=7.095 $Y=1.05 $X2=0
+ $Y2=0
cc_509 N_C_c_686_n N_A_1348_111#_c_766_n 0.0113495f $X=8.095 $Y=0.975 $X2=0
+ $Y2=0
cc_510 N_C_c_688_n N_A_1348_111#_c_766_n 0.00433478f $X=8.57 $Y=1.155 $X2=0
+ $Y2=0
cc_511 N_C_c_692_n N_A_1348_111#_c_766_n 0.00391291f $X=7.73 $Y=1.14 $X2=0 $Y2=0
cc_512 N_C_c_686_n N_A_1348_111#_c_767_n 0.00233917f $X=8.095 $Y=0.975 $X2=0
+ $Y2=0
cc_513 N_C_c_688_n N_A_1348_111#_c_767_n 0.00120986f $X=8.57 $Y=1.155 $X2=0
+ $Y2=0
cc_514 N_C_M1000_g N_VPWR_c_843_n 0.0236984f $X=8.745 $Y=2.505 $X2=0 $Y2=0
cc_515 N_C_M1000_g N_VPWR_c_847_n 0.00717535f $X=8.745 $Y=2.505 $X2=0 $Y2=0
cc_516 N_C_M1000_g N_VPWR_c_840_n 0.0133121f $X=8.745 $Y=2.505 $X2=0 $Y2=0
cc_517 N_C_M1022_g N_A_763_347#_c_979_n 0.00249917f $X=7.365 $Y=2.165 $X2=0
+ $Y2=0
cc_518 N_C_M1000_g N_A_763_347#_c_979_n 2.32496e-19 $X=8.745 $Y=2.505 $X2=0
+ $Y2=0
cc_519 N_C_c_683_n N_A_763_347#_c_973_n 5.56873e-19 $X=7.095 $Y=1.05 $X2=0 $Y2=0
cc_520 N_C_M1022_g N_A_763_347#_c_973_n 0.0254028f $X=7.365 $Y=2.165 $X2=0 $Y2=0
cc_521 N_C_c_685_n N_A_763_347#_c_973_n 0.00627918f $X=7.49 $Y=1.125 $X2=0 $Y2=0
cc_522 N_C_c_691_n N_A_763_347#_c_973_n 0.0258428f $X=7.895 $Y=1.14 $X2=0 $Y2=0
cc_523 N_C_c_692_n N_A_763_347#_c_973_n 0.00449992f $X=7.73 $Y=1.14 $X2=0 $Y2=0
cc_524 N_C_c_693_n N_A_763_347#_c_973_n 0.00119876f $X=8.17 $Y=1.14 $X2=0 $Y2=0
cc_525 N_C_c_691_n N_A_763_347#_c_981_n 0.0112754f $X=7.895 $Y=1.14 $X2=0 $Y2=0
cc_526 N_C_c_693_n N_A_763_347#_c_981_n 0.00161115f $X=8.17 $Y=1.14 $X2=0 $Y2=0
cc_527 N_C_M1022_g N_A_763_347#_c_1034_n 0.0100246f $X=7.365 $Y=2.165 $X2=0
+ $Y2=0
cc_528 N_C_M1022_g N_A_763_347#_c_982_n 0.00568497f $X=7.365 $Y=2.165 $X2=0
+ $Y2=0
cc_529 N_C_c_683_n N_A_763_347#_c_974_n 0.00510171f $X=7.095 $Y=1.05 $X2=0 $Y2=0
cc_530 N_C_c_685_n N_A_763_347#_c_974_n 0.0106827f $X=7.49 $Y=1.125 $X2=0 $Y2=0
cc_531 N_C_c_686_n N_A_763_347#_c_974_n 0.00405931f $X=8.095 $Y=0.975 $X2=0
+ $Y2=0
cc_532 N_C_c_691_n N_A_763_347#_c_974_n 0.00138097f $X=7.895 $Y=1.14 $X2=0 $Y2=0
cc_533 N_C_M1022_g N_A_803_81#_c_1146_n 0.016282f $X=7.365 $Y=2.165 $X2=0 $Y2=0
cc_534 N_C_M1022_g N_A_803_81#_c_1109_n 0.00542421f $X=7.365 $Y=2.165 $X2=0
+ $Y2=0
cc_535 N_C_M1000_g X 0.00227982f $X=8.745 $Y=2.505 $X2=0 $Y2=0
cc_536 N_C_c_688_n N_VGND_c_1213_n 0.00272516f $X=8.57 $Y=1.155 $X2=0 $Y2=0
cc_537 N_C_c_690_n N_VGND_c_1213_n 9.8317e-19 $X=8.682 $Y=1.23 $X2=0 $Y2=0
cc_538 N_C_c_683_n N_VGND_c_1214_n 6.31558e-19 $X=7.095 $Y=1.05 $X2=0 $Y2=0
cc_539 N_C_c_686_n N_VGND_c_1214_n 8.28597e-19 $X=8.095 $Y=0.975 $X2=0 $Y2=0
cc_540 N_A_1348_111#_M1013_g N_VPWR_c_843_n 0.0254822f $X=9.275 $Y=2.505 $X2=0
+ $Y2=0
cc_541 N_A_1348_111#_M1013_g N_VPWR_c_848_n 0.00716274f $X=9.275 $Y=2.505 $X2=0
+ $Y2=0
cc_542 N_A_1348_111#_M1013_g N_VPWR_c_840_n 0.0135748f $X=9.275 $Y=2.505 $X2=0
+ $Y2=0
cc_543 N_A_1348_111#_c_763_n N_A_763_347#_c_973_n 0.0255648f $X=6.88 $Y=0.765
+ $X2=0 $Y2=0
cc_544 N_A_1348_111#_c_770_n N_A_763_347#_c_973_n 0.0114277f $X=7.1 $Y=1.81
+ $X2=0 $Y2=0
cc_545 N_A_1348_111#_c_763_n N_A_763_347#_c_974_n 0.0146643f $X=6.88 $Y=0.765
+ $X2=0 $Y2=0
cc_546 N_A_1348_111#_c_770_n N_A_763_347#_c_974_n 0.00120987f $X=7.1 $Y=1.81
+ $X2=0 $Y2=0
cc_547 N_A_1348_111#_c_766_n N_A_763_347#_c_974_n 0.0254701f $X=8.855 $Y=0.407
+ $X2=0 $Y2=0
cc_548 N_A_1348_111#_c_764_n N_A_803_81#_c_1105_n 0.0124434f $X=6.965 $Y=0.35
+ $X2=0 $Y2=0
cc_549 N_A_1348_111#_c_763_n N_A_803_81#_c_1107_n 0.0681003f $X=6.88 $Y=0.765
+ $X2=0 $Y2=0
cc_550 N_A_1348_111#_c_770_n N_A_803_81#_c_1107_n 0.0191929f $X=7.1 $Y=1.81
+ $X2=0 $Y2=0
cc_551 N_A_1348_111#_c_770_n N_A_803_81#_c_1144_n 0.00811737f $X=7.1 $Y=1.81
+ $X2=0 $Y2=0
cc_552 N_A_1348_111#_M1007_d N_A_803_81#_c_1146_n 0.00480382f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_A_1348_111#_c_770_n N_A_803_81#_c_1146_n 0.00746126f $X=7.1 $Y=1.81
+ $X2=0 $Y2=0
cc_554 N_A_1348_111#_c_770_n N_A_803_81#_c_1141_n 0.00891688f $X=7.1 $Y=1.81
+ $X2=0 $Y2=0
cc_555 N_A_1348_111#_c_762_n N_X_c_1186_n 0.00478687f $X=9.585 $Y=0.55 $X2=0
+ $Y2=0
cc_556 N_A_1348_111#_M1001_g X 0.0114815f $X=9.225 $Y=0.87 $X2=0 $Y2=0
cc_557 N_A_1348_111#_c_759_n X 0.00158787f $X=9.275 $Y=1.575 $X2=0 $Y2=0
cc_558 N_A_1348_111#_c_762_n X 0.0119024f $X=9.585 $Y=0.55 $X2=0 $Y2=0
cc_559 N_A_1348_111#_c_759_n X 0.00442094f $X=9.275 $Y=1.575 $X2=0 $Y2=0
cc_560 N_A_1348_111#_M1013_g X 0.0291294f $X=9.275 $Y=2.505 $X2=0 $Y2=0
cc_561 N_A_1348_111#_M1013_g X 0.00793154f $X=9.275 $Y=2.505 $X2=0 $Y2=0
cc_562 N_A_1348_111#_M1001_g N_VGND_c_1265_n 0.0125264f $X=9.225 $Y=0.87 $X2=0
+ $Y2=0
cc_563 N_A_1348_111#_c_759_n N_VGND_c_1265_n 0.00158737f $X=9.275 $Y=1.575 $X2=0
+ $Y2=0
cc_564 N_A_1348_111#_c_762_n N_VGND_c_1265_n 0.00386627f $X=9.585 $Y=0.55 $X2=0
+ $Y2=0
cc_565 N_A_1348_111#_c_765_n N_VGND_c_1265_n 6.46283e-19 $X=9.02 $Y=0.385 $X2=0
+ $Y2=0
cc_566 N_A_1348_111#_M1001_g N_VGND_c_1210_n 0.00405014f $X=9.225 $Y=0.87 $X2=0
+ $Y2=0
cc_567 N_A_1348_111#_c_761_n N_VGND_c_1210_n 0.0145327f $X=9.51 $Y=0.475 $X2=0
+ $Y2=0
cc_568 N_A_1348_111#_c_762_n N_VGND_c_1210_n 0.00555249f $X=9.585 $Y=0.55 $X2=0
+ $Y2=0
cc_569 N_A_1348_111#_c_765_n N_VGND_c_1210_n 0.0206124f $X=9.02 $Y=0.385 $X2=0
+ $Y2=0
cc_570 N_A_1348_111#_c_767_n N_VGND_c_1210_n 0.00542684f $X=9.3 $Y=0.385 $X2=0
+ $Y2=0
cc_571 N_A_1348_111#_M1001_g N_VGND_c_1213_n 0.00654256f $X=9.225 $Y=0.87 $X2=0
+ $Y2=0
cc_572 N_A_1348_111#_c_762_n N_VGND_c_1213_n 6.42933e-19 $X=9.585 $Y=0.55 $X2=0
+ $Y2=0
cc_573 N_A_1348_111#_c_765_n N_VGND_c_1213_n 0.0205545f $X=9.02 $Y=0.385 $X2=0
+ $Y2=0
cc_574 N_A_1348_111#_c_766_n N_VGND_c_1213_n 3.97099e-19 $X=8.855 $Y=0.407 $X2=0
+ $Y2=0
cc_575 N_A_1348_111#_c_767_n N_VGND_c_1213_n 0.00636571f $X=9.3 $Y=0.385 $X2=0
+ $Y2=0
cc_576 N_A_1348_111#_c_761_n N_VGND_c_1214_n 0.0015682f $X=9.51 $Y=0.475 $X2=0
+ $Y2=0
cc_577 N_A_1348_111#_c_764_n N_VGND_c_1214_n 0.0168561f $X=6.965 $Y=0.35 $X2=0
+ $Y2=0
cc_578 N_A_1348_111#_c_766_n N_VGND_c_1214_n 0.134275f $X=8.855 $Y=0.407 $X2=0
+ $Y2=0
cc_579 N_A_1348_111#_c_767_n N_VGND_c_1214_n 0.00859812f $X=9.3 $Y=0.385 $X2=0
+ $Y2=0
cc_580 N_A_1348_111#_c_761_n N_VGND_c_1217_n 0.0038983f $X=9.51 $Y=0.475 $X2=0
+ $Y2=0
cc_581 N_A_1348_111#_c_761_n N_VGND_c_1218_n 0.00633754f $X=9.51 $Y=0.475 $X2=0
+ $Y2=0
cc_582 N_A_1348_111#_c_764_n N_VGND_c_1218_n 0.00967329f $X=6.965 $Y=0.35 $X2=0
+ $Y2=0
cc_583 N_A_1348_111#_c_766_n N_VGND_c_1218_n 0.0815909f $X=8.855 $Y=0.407 $X2=0
+ $Y2=0
cc_584 N_A_1348_111#_c_767_n N_VGND_c_1218_n 0.0117385f $X=9.3 $Y=0.385 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_841_n N_A_265_409#_c_908_n 0.0428289f $X=0.935 $Y=2.19 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_846_n N_A_265_409#_c_908_n 0.0219574f $X=2.6 $Y=3.33 $X2=0 $Y2=0
cc_587 N_VPWR_c_840_n N_A_265_409#_c_908_n 0.0125652f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_588 N_VPWR_M1003_s N_A_265_409#_c_910_n 0.00991155f $X=2.62 $Y=1.835 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_842_n N_A_265_409#_c_910_n 0.0255507f $X=2.765 $Y=2.76 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_841_n N_A_265_409#_c_912_n 0.02688f $X=0.935 $Y=2.19 $X2=0 $Y2=0
cc_591 N_VPWR_c_847_n N_A_763_347#_c_975_n 0.0478559f $X=8.845 $Y=3.33 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_840_n N_A_763_347#_c_975_n 0.0263693f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_593 N_VPWR_c_847_n N_A_763_347#_c_977_n 0.0741759f $X=8.845 $Y=3.33 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_840_n N_A_763_347#_c_977_n 0.0411363f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_847_n N_A_763_347#_c_979_n 0.0825594f $X=8.845 $Y=3.33 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_840_n N_A_763_347#_c_979_n 0.0466377f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_847_n N_A_763_347#_c_983_n 0.0215054f $X=8.845 $Y=3.33 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_840_n N_A_763_347#_c_983_n 0.0112592f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_VPWR_c_847_n N_A_763_347#_c_984_n 0.0112749f $X=8.845 $Y=3.33 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_840_n N_A_763_347#_c_984_n 0.0058379f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_847_n N_A_763_347#_c_985_n 0.0218455f $X=8.845 $Y=3.33 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_840_n N_A_763_347#_c_985_n 0.0125874f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_843_n X 0.0420241f $X=9.01 $Y=2.15 $X2=0 $Y2=0
cc_604 N_VPWR_c_843_n X 0.0293627f $X=9.01 $Y=2.15 $X2=0 $Y2=0
cc_605 N_VPWR_c_848_n X 0.0263342f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_606 N_VPWR_c_840_n X 0.0214424f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_607 N_A_265_409#_c_910_n N_A_763_347#_M1011_s 0.0102945f $X=4.405 $Y=2.33
+ $X2=0 $Y2=0
cc_608 N_A_265_409#_c_910_n N_A_763_347#_c_975_n 0.0304643f $X=4.405 $Y=2.33
+ $X2=0 $Y2=0
cc_609 N_A_265_409#_M1011_d N_A_763_347#_c_976_n 0.00751289f $X=4.43 $Y=1.735
+ $X2=0 $Y2=0
cc_610 N_A_265_409#_c_910_n N_A_763_347#_c_976_n 0.0353261f $X=4.405 $Y=2.33
+ $X2=0 $Y2=0
cc_611 N_A_265_409#_c_911_n N_A_763_347#_c_976_n 0.0204345f $X=4.57 $Y=1.88
+ $X2=0 $Y2=0
cc_612 N_A_265_409#_c_906_n N_A_763_347#_c_987_n 8.37456e-19 $X=4.57 $Y=1.415
+ $X2=0 $Y2=0
cc_613 N_A_265_409#_M1011_d N_A_763_347#_c_1006_n 0.00281591f $X=4.43 $Y=1.735
+ $X2=0 $Y2=0
cc_614 N_A_265_409#_c_906_n N_A_763_347#_c_1006_n 0.0069487f $X=4.57 $Y=1.415
+ $X2=0 $Y2=0
cc_615 N_A_265_409#_c_911_n N_A_763_347#_c_1006_n 0.0139033f $X=4.57 $Y=1.88
+ $X2=0 $Y2=0
cc_616 N_A_265_409#_c_906_n N_A_763_347#_c_972_n 0.0258114f $X=4.57 $Y=1.415
+ $X2=0 $Y2=0
cc_617 N_A_265_409#_c_911_n N_A_763_347#_c_972_n 0.0115926f $X=4.57 $Y=1.88
+ $X2=0 $Y2=0
cc_618 N_A_265_409#_c_910_n N_A_763_347#_c_983_n 0.0247986f $X=4.405 $Y=2.33
+ $X2=0 $Y2=0
cc_619 N_A_763_347#_c_987_n N_A_803_81#_M1014_d 0.00188202f $X=5.285 $Y=1.88
+ $X2=0 $Y2=0
cc_620 N_A_763_347#_c_981_n N_A_803_81#_M1022_d 0.012912f $X=7.895 $Y=2.06 $X2=0
+ $Y2=0
cc_621 N_A_763_347#_c_976_n N_A_803_81#_c_1127_n 0.0265673f $X=5 $Y=2.895 $X2=0
+ $Y2=0
cc_622 N_A_763_347#_c_977_n N_A_803_81#_c_1127_n 0.0196464f $X=6.325 $Y=2.98
+ $X2=0 $Y2=0
cc_623 N_A_763_347#_c_987_n N_A_803_81#_c_1119_n 0.00132326f $X=5.285 $Y=1.88
+ $X2=0 $Y2=0
cc_624 N_A_763_347#_c_977_n N_A_803_81#_c_1119_n 0.0185263f $X=6.325 $Y=2.98
+ $X2=0 $Y2=0
cc_625 N_A_763_347#_c_976_n N_A_803_81#_c_1129_n 0.0130518f $X=5 $Y=2.895 $X2=0
+ $Y2=0
cc_626 N_A_763_347#_c_987_n N_A_803_81#_c_1129_n 0.0179065f $X=5.285 $Y=1.88
+ $X2=0 $Y2=0
cc_627 N_A_763_347#_M1016_d N_A_803_81#_c_1107_n 0.00522312f $X=6.35 $Y=1.735
+ $X2=0 $Y2=0
cc_628 N_A_763_347#_M1016_d N_A_803_81#_c_1144_n 0.00730313f $X=6.35 $Y=1.735
+ $X2=0 $Y2=0
cc_629 N_A_763_347#_c_978_n N_A_803_81#_c_1144_n 0.0136235f $X=6.49 $Y=2.59
+ $X2=0 $Y2=0
cc_630 N_A_763_347#_c_979_n N_A_803_81#_c_1144_n 0.00398181f $X=7.895 $Y=2.98
+ $X2=0 $Y2=0
cc_631 N_A_763_347#_c_979_n N_A_803_81#_c_1146_n 0.0146388f $X=7.895 $Y=2.98
+ $X2=0 $Y2=0
cc_632 N_A_763_347#_c_1034_n N_A_803_81#_c_1146_n 0.00723403f $X=7.535 $Y=2.06
+ $X2=0 $Y2=0
cc_633 N_A_763_347#_M1016_d N_A_803_81#_c_1140_n 7.59612e-19 $X=6.35 $Y=1.735
+ $X2=0 $Y2=0
cc_634 N_A_763_347#_c_977_n N_A_803_81#_c_1140_n 5.32803e-19 $X=6.325 $Y=2.98
+ $X2=0 $Y2=0
cc_635 N_A_763_347#_c_978_n N_A_803_81#_c_1140_n 0.00761838f $X=6.49 $Y=2.59
+ $X2=0 $Y2=0
cc_636 N_A_763_347#_c_979_n N_A_803_81#_c_1141_n 0.00472935f $X=7.895 $Y=2.98
+ $X2=0 $Y2=0
cc_637 N_A_763_347#_c_979_n N_A_803_81#_c_1109_n 0.0156564f $X=7.895 $Y=2.98
+ $X2=0 $Y2=0
cc_638 N_A_763_347#_c_981_n N_A_803_81#_c_1109_n 0.0123718f $X=7.895 $Y=2.06
+ $X2=0 $Y2=0
cc_639 N_A_763_347#_c_1034_n N_A_803_81#_c_1109_n 0.00181339f $X=7.535 $Y=2.06
+ $X2=0 $Y2=0
cc_640 N_A_763_347#_c_982_n N_A_803_81#_c_1109_n 0.0263226f $X=7.98 $Y=2.895
+ $X2=0 $Y2=0
cc_641 N_A_803_81#_c_1105_n N_VGND_c_1214_n 0.131782f $X=6.305 $Y=0.35 $X2=0
+ $Y2=0
cc_642 N_A_803_81#_c_1106_n N_VGND_c_1214_n 0.0105618f $X=4.245 $Y=0.35 $X2=0
+ $Y2=0
cc_643 N_A_803_81#_c_1105_n N_VGND_c_1218_n 0.0763154f $X=6.305 $Y=0.35 $X2=0
+ $Y2=0
cc_644 N_A_803_81#_c_1106_n N_VGND_c_1218_n 0.00572509f $X=4.245 $Y=0.35 $X2=0
+ $Y2=0
cc_645 X N_VGND_c_1265_n 0.0082067f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_646 N_X_c_1186_n N_VGND_c_1210_n 0.00360907f $X=9.8 $Y=0.87 $X2=0 $Y2=0
cc_647 N_X_c_1186_n N_VGND_c_1213_n 0.00327227f $X=9.8 $Y=0.87 $X2=0 $Y2=0
cc_648 N_X_c_1186_n N_VGND_c_1217_n 0.00497092f $X=9.8 $Y=0.87 $X2=0 $Y2=0
cc_649 N_X_c_1186_n N_VGND_c_1218_n 0.00749824f $X=9.8 $Y=0.87 $X2=0 $Y2=0
cc_650 N_VGND_c_1265_n A_1860_132# 0.00146512f $X=9.365 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_651 N_VGND_c_1210_n A_1860_132# 7.6006e-19 $X=9.45 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
