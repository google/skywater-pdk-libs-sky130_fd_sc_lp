* File: sky130_fd_sc_lp__dlrbn_lp.pex.spice
* Created: Fri Aug 28 10:25:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%D 3 7 11 15 17 18 19 23 24
c45 24 0 1.43466e-19 $X=0.605 $Y=1.255
c46 7 0 9.04602e-20 $X=0.605 $Y=2.48
r47 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.255 $X2=0.605 $Y2=1.255
r48 18 19 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.637 $Y=1.295
+ $X2=0.637 $Y2=1.665
r49 18 24 1.16703 $w=3.93e-07 $l=4e-08 $layer=LI1_cond $X=0.637 $Y=1.295
+ $X2=0.637 $Y2=1.255
r50 16 23 54.4068 $w=3.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.595 $Y=1.585
+ $X2=0.595 $Y2=1.255
r51 16 17 31.5166 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.585
+ $X2=0.595 $Y2=1.76
r52 15 23 2.47304 $w=3.5e-07 $l=1.5e-08 $layer=POLY_cond $X=0.595 $Y=1.24
+ $X2=0.595 $Y2=1.255
r53 7 17 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.605 $Y=2.48
+ $X2=0.605 $Y2=1.76
r54 1 15 26.0701 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=1.09
+ $X2=0.675 $Y2=1.24
r55 1 11 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.855 $Y=1.09
+ $X2=0.855 $Y2=0.55
r56 1 3 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.495 $Y=1.09
+ $X2=0.495 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%GATE_N 3 7 11 15 20 22 23 27 28
c54 28 0 1.90141e-20 $X=1.335 $Y=1.125
c55 20 0 1.43466e-19 $X=1.645 $Y=1.035
r56 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.335
+ $Y=1.125 $X2=1.335 $Y2=1.125
r57 22 23 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.292 $Y=1.295
+ $X2=1.292 $Y2=1.665
r58 22 28 4.72085 $w=4.13e-07 $l=1.7e-07 $layer=LI1_cond $X=1.292 $Y=1.295
+ $X2=1.292 $Y2=1.125
r59 19 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.335 $Y=1.11
+ $X2=1.335 $Y2=1.125
r60 19 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.335 $Y=1.035
+ $X2=1.645 $Y2=1.035
r61 16 19 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=1.285 $Y=1.035
+ $X2=1.335 $Y2=1.035
r62 14 27 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.335 $Y=1.48
+ $X2=1.335 $Y2=1.125
r63 14 15 29.7575 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.255 $Y=1.48
+ $X2=1.255 $Y2=1.63
r64 9 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.645 $Y=0.96
+ $X2=1.645 $Y2=1.035
r65 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.645 $Y=0.96
+ $X2=1.645 $Y2=0.55
r66 5 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.285 $Y=0.96
+ $X2=1.285 $Y2=1.035
r67 5 7 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.285 $Y=0.96
+ $X2=1.285 $Y2=0.55
r68 3 15 211.186 $w=2.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.135 $Y=2.48
+ $X2=1.135 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%A_252_396# 1 2 7 8 9 11 14 17 20 24 27 28
+ 30 38 41 42 45 47 48 54 60 63 64 66 67 68 72
c152 68 0 1.52433e-20 $X=4.195 $Y=0.94
c153 38 0 1.53546e-19 $X=2.995 $Y=0.93
c154 17 0 1.65112e-19 $X=2.715 $Y=1.87
r155 72 79 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=4.195 $Y=1.02
+ $X2=4.315 $Y2=1.02
r156 72 77 13.7714 $w=3.15e-07 $l=9e-08 $layer=POLY_cond $X=4.195 $Y=1.02
+ $X2=4.105 $Y2=1.02
r157 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.195
+ $Y=1.02 $X2=4.195 $Y2=1.02
r158 68 71 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.195 $Y=0.94
+ $X2=4.195 $Y2=1.02
r159 66 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.595
+ $Y=1.02 $X2=2.595 $Y2=1.02
r160 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.865
+ $Y=2.125 $X2=1.865 $Y2=2.125
r161 61 66 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.695 $Y=0.94
+ $X2=2.595 $Y2=0.94
r162 60 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=0.94
+ $X2=4.195 $Y2=0.94
r163 60 61 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=4.03 $Y=0.94
+ $X2=2.695 $Y2=0.94
r164 52 63 4.84325 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=1.96
+ $X2=1.83 $Y2=2.085
r165 52 54 60.1831 $w=2.68e-07 $l=1.41e-06 $layer=LI1_cond $X=1.83 $Y=1.96
+ $X2=1.83 $Y2=0.55
r166 48 63 1.62111 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=1.695 $Y=2.085
+ $X2=1.83 $Y2=2.085
r167 48 50 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.695 $Y=2.085
+ $X2=1.4 $Y2=2.085
r168 43 45 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=4.315 $Y=1.6
+ $X2=4.445 $Y2=1.6
r169 40 67 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=2.61 $Y=1.345
+ $X2=2.61 $Y2=1.02
r170 40 41 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=2.61 $Y=1.345
+ $X2=2.61 $Y2=1.525
r171 37 38 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.635 $Y=0.93
+ $X2=2.995 $Y2=0.93
r172 35 67 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=2.61 $Y=1.005
+ $X2=2.61 $Y2=1.02
r173 35 37 12.8191 $w=1.5e-07 $l=2.5e-08 $layer=POLY_cond $X=2.61 $Y=0.93
+ $X2=2.635 $Y2=0.93
r174 33 64 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.865 $Y=2.02
+ $X2=1.865 $Y2=2.125
r175 31 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.445 $Y=1.675
+ $X2=4.445 $Y2=1.6
r176 31 47 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.445 $Y=1.675
+ $X2=4.445 $Y2=1.885
r177 28 47 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.395 $Y=2.01
+ $X2=4.395 $Y2=1.885
r178 28 30 112.788 $w=2.5e-07 $l=5.85e-07 $layer=POLY_cond $X=4.395 $Y=2.01
+ $X2=4.395 $Y2=2.595
r179 27 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.315 $Y=1.525
+ $X2=4.315 $Y2=1.6
r180 26 79 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.185
+ $X2=4.315 $Y2=1.02
r181 26 27 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.315 $Y=1.185
+ $X2=4.315 $Y2=1.525
r182 22 77 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=0.855
+ $X2=4.105 $Y2=1.02
r183 22 24 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.105 $Y=0.855
+ $X2=4.105 $Y2=0.445
r184 18 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.995 $Y=0.855
+ $X2=2.995 $Y2=0.93
r185 18 20 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.995 $Y=0.855
+ $X2=2.995 $Y2=0.445
r186 17 42 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=2.715 $Y=1.87
+ $X2=2.665 $Y2=1.945
r187 17 41 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.715 $Y=1.87
+ $X2=2.715 $Y2=1.525
r188 12 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.635 $Y=0.855
+ $X2=2.635 $Y2=0.93
r189 12 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.635 $Y=0.855
+ $X2=2.635 $Y2=0.445
r190 9 42 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=2.665 $Y=2.02
+ $X2=2.665 $Y2=1.945
r191 9 11 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.665 $Y=2.02
+ $X2=2.665 $Y2=2.595
r192 8 33 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.03 $Y=1.945
+ $X2=1.865 $Y2=2.02
r193 7 42 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.54 $Y=1.945
+ $X2=2.665 $Y2=1.945
r194 7 8 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.54 $Y=1.945
+ $X2=2.03 $Y2=1.945
r195 2 50 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=1.98 $X2=1.4 $Y2=2.125
r196 1 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.34 $X2=1.86 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%A_27_68# 1 2 9 13 14 15 17 21 24 26 29 30
+ 31 33 34 35 38 39 42 46 47 48 50
c124 39 0 5.71049e-20 $X=3.325 $Y=1.77
c125 38 0 3.46692e-19 $X=3.325 $Y=1.77
c126 31 0 7.14461e-20 $X=1.385 $Y=2.98
c127 13 0 1.52433e-20 $X=3.64 $Y=0.805
c128 9 0 1.85755e-19 $X=3.365 $Y=2.595
r129 46 47 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.297 $Y=2.125
+ $X2=0.297 $Y2=1.96
r130 44 47 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=0.175 $Y=0.78
+ $X2=0.175 $Y2=1.96
r131 42 44 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=0.267 $Y=0.55
+ $X2=0.267 $Y2=0.78
r132 39 51 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.325 $Y=1.77
+ $X2=3.325 $Y2=1.935
r133 39 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.325 $Y=1.77
+ $X2=3.325 $Y2=1.605
r134 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.325
+ $Y=1.77 $X2=3.325 $Y2=1.77
r135 36 38 12.3942 $w=2.63e-07 $l=2.85e-07 $layer=LI1_cond $X=3.357 $Y=2.055
+ $X2=3.357 $Y2=1.77
r136 34 36 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.225 $Y=2.14
+ $X2=3.357 $Y2=2.055
r137 34 35 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.225 $Y=2.14
+ $X2=2.835 $Y2=2.14
r138 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.75 $Y=2.225
+ $X2=2.835 $Y2=2.14
r139 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.75 $Y=2.225
+ $X2=2.75 $Y2=2.895
r140 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.665 $Y=2.98
+ $X2=2.75 $Y2=2.895
r141 30 31 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=2.665 $Y=2.98
+ $X2=1.385 $Y2=2.98
r142 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.3 $Y=2.895
+ $X2=1.385 $Y2=2.98
r143 28 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.3 $Y=2.56
+ $X2=1.3 $Y2=2.895
r144 27 48 4.68428 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.505 $Y=2.475
+ $X2=0.297 $Y2=2.475
r145 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.215 $Y=2.475
+ $X2=1.3 $Y2=2.56
r146 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.215 $Y=2.475
+ $X2=0.505 $Y2=2.475
r147 22 48 2.337 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=2.56
+ $X2=0.297 $Y2=2.475
r148 22 24 7.63667 $w=4.13e-07 $l=2.75e-07 $layer=LI1_cond $X=0.297 $Y=2.56
+ $X2=0.297 $Y2=2.835
r149 21 48 2.337 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=2.39
+ $X2=0.297 $Y2=2.475
r150 20 46 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=0.297 $Y=2.167
+ $X2=0.297 $Y2=2.125
r151 20 21 6.19265 $w=4.13e-07 $l=2.23e-07 $layer=LI1_cond $X=0.297 $Y=2.167
+ $X2=0.297 $Y2=2.39
r152 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.715 $Y=0.73
+ $X2=3.715 $Y2=0.445
r153 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.64 $Y=0.805
+ $X2=3.715 $Y2=0.73
r154 13 14 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.64 $Y=0.805
+ $X2=3.46 $Y2=0.805
r155 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.385 $Y=0.88
+ $X2=3.46 $Y2=0.805
r156 11 50 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=3.385 $Y=0.88
+ $X2=3.385 $Y2=1.605
r157 9 51 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.365 $Y=2.595
+ $X2=3.365 $Y2=1.935
r158 2 46 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.98 $X2=0.34 $Y2=2.125
r159 2 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.98 $X2=0.34 $Y2=2.835
r160 1 42 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.34 $X2=0.28 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%A_451_419# 1 2 9 13 16 19 21 24 25 26 27 30
+ 34 36 38 41 43 44
c136 41 0 1.8158e-19 $X=3.865 $Y=1.59
c137 25 0 1.53546e-19 $X=3.68 $Y=1.34
r138 44 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.765 $Y=1.12
+ $X2=4.765 $Y2=0.955
r139 43 46 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=1.12
+ $X2=4.765 $Y2=1.285
r140 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.765
+ $Y=1.12 $X2=4.765 $Y2=1.12
r141 41 49 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.865 $Y=1.59
+ $X2=3.865 $Y2=1.755
r142 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.865
+ $Y=1.59 $X2=3.865 $Y2=1.59
r143 38 40 3.38889 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=3.855 $Y=1.51
+ $X2=3.855 $Y2=1.59
r144 31 34 5.34059 $w=4.08e-07 $l=1.9e-07 $layer=LI1_cond $X=2.23 $Y=0.47
+ $X2=2.42 $Y2=0.47
r145 30 46 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.685 $Y=1.425
+ $X2=4.685 $Y2=1.285
r146 28 38 3.82142 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.03 $Y=1.51
+ $X2=3.855 $Y2=1.51
r147 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.6 $Y=1.51
+ $X2=4.685 $Y2=1.425
r148 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.6 $Y=1.51
+ $X2=4.03 $Y2=1.51
r149 25 38 7.20139 $w=2.88e-07 $l=2.45713e-07 $layer=LI1_cond $X=3.68 $Y=1.34
+ $X2=3.855 $Y2=1.51
r150 25 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.68 $Y=1.34
+ $X2=3.045 $Y2=1.34
r151 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.96 $Y=1.425
+ $X2=3.045 $Y2=1.34
r152 23 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.96 $Y=1.425
+ $X2=2.96 $Y2=1.705
r153 22 36 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.485 $Y=1.79
+ $X2=2.315 $Y2=1.79
r154 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.875 $Y=1.79
+ $X2=2.96 $Y2=1.705
r155 21 22 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.875 $Y=1.79
+ $X2=2.485 $Y2=1.79
r156 17 36 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=1.875
+ $X2=2.315 $Y2=1.79
r157 17 19 17.6256 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=2.315 $Y=1.875
+ $X2=2.315 $Y2=2.395
r158 16 36 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.23 $Y=1.705
+ $X2=2.315 $Y2=1.79
r159 15 31 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.23 $Y=0.675
+ $X2=2.23 $Y2=0.47
r160 15 16 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.23 $Y=0.675
+ $X2=2.23 $Y2=1.705
r161 13 51 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.675 $Y=0.445
+ $X2=4.675 $Y2=0.955
r162 9 49 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.855 $Y=2.595
+ $X2=3.855 $Y2=1.755
r163 2 19 600 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=1 $X=2.255
+ $Y=2.095 $X2=2.4 $Y2=2.395
r164 1 34 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.42 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%A_952_305# 1 2 9 13 15 17 18 20 23 25 29 33
+ 37 41 46 49 51 52 56 58 60 63 68 70 76 83
c163 83 0 1.61435e-20 $X=7.75 $Y=1.46
c164 63 0 3.08053e-20 $X=6.095 $Y=1.04
r165 82 83 39.217 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.625 $Y=1.46
+ $X2=7.75 $Y2=1.46
r166 81 82 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.46
+ $X2=7.625 $Y2=1.46
r167 71 81 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=7.165 $Y=1.46
+ $X2=7.46 $Y2=1.46
r168 71 78 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.165 $Y=1.46
+ $X2=7.1 $Y2=1.46
r169 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.165
+ $Y=1.46 $X2=7.165 $Y2=1.46
r170 67 70 7.31957 $w=3.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.93 $Y=1.44
+ $X2=7.165 $Y2=1.44
r171 67 68 6.04704 $w=3.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=1.44
+ $X2=6.845 $Y2=1.44
r172 63 65 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.175 $Y=1.04
+ $X2=6.175 $Y2=1.34
r173 59 76 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.13 $Y=1.69
+ $X2=5.215 $Y2=1.69
r174 59 73 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=5.13 $Y=1.69
+ $X2=4.885 $Y2=1.69
r175 58 60 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=1.69
+ $X2=5.13 $Y2=1.525
r176 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.69 $X2=5.13 $Y2=1.69
r177 55 67 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.93 $Y=1.625
+ $X2=6.93 $Y2=1.44
r178 55 56 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=6.93 $Y=1.625
+ $X2=6.93 $Y2=2.7
r179 54 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=1.34
+ $X2=6.175 $Y2=1.34
r180 54 68 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.26 $Y=1.34
+ $X2=6.845 $Y2=1.34
r181 51 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.845 $Y=2.785
+ $X2=6.93 $Y2=2.7
r182 51 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.845 $Y=2.785
+ $X2=6.155 $Y2=2.785
r183 47 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.99 $Y=2.7
+ $X2=6.155 $Y2=2.785
r184 47 49 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5.99 $Y=2.7
+ $X2=5.99 $Y2=2.24
r185 46 63 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=5.295 $Y=1.08
+ $X2=6.09 $Y2=1.08
r186 43 46 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.21 $Y=1.205
+ $X2=5.295 $Y2=1.08
r187 43 60 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.21 $Y=1.205
+ $X2=5.21 $Y2=1.525
r188 35 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.8 $Y=1.295
+ $X2=8.8 $Y2=1.37
r189 35 37 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=8.8 $Y=1.295 $X2=8.8
+ $Y2=0.59
r190 31 41 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=8.75 $Y=1.37 $X2=8.8
+ $Y2=1.37
r191 31 39 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=8.75 $Y=1.37
+ $X2=8.44 $Y2=1.37
r192 31 33 229.82 $w=2.5e-07 $l=9.25e-07 $layer=POLY_cond $X=8.75 $Y=1.445
+ $X2=8.75 $Y2=2.37
r193 27 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.44 $Y=1.295
+ $X2=8.44 $Y2=1.37
r194 27 29 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=8.44 $Y=1.295
+ $X2=8.44 $Y2=0.59
r195 25 39 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.365 $Y=1.37
+ $X2=8.44 $Y2=1.37
r196 25 83 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=8.365 $Y=1.37
+ $X2=7.75 $Y2=1.37
r197 21 82 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.625 $Y=1.625
+ $X2=7.625 $Y2=1.46
r198 21 23 241 $w=2.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.625 $Y=1.625
+ $X2=7.625 $Y2=2.595
r199 18 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.295
+ $X2=7.46 $Y2=1.46
r200 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.46 $Y=1.295
+ $X2=7.46 $Y2=0.975
r201 15 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.1 $Y=1.295
+ $X2=7.1 $Y2=1.46
r202 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.1 $Y=1.295
+ $X2=7.1 $Y2=0.975
r203 11 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.215 $Y=1.525
+ $X2=5.215 $Y2=1.69
r204 11 13 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=5.215 $Y=1.525
+ $X2=5.215 $Y2=0.445
r205 7 73 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.885 $Y=1.855
+ $X2=4.885 $Y2=1.69
r206 7 9 183.856 $w=2.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.885 $Y=1.855
+ $X2=4.885 $Y2=2.595
r207 2 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.85
+ $Y=2.095 $X2=5.99 $Y2=2.24
r208 1 63 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.955
+ $Y=0.765 $X2=6.095 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%A_796_419# 1 2 9 13 15 18 20 21 22 25 27 32
+ 33 36 37 42
c110 36 0 4.84139e-20 $X=6.02 $Y=0.49
c111 21 0 1.85755e-19 $X=4.295 $Y=2.12
c112 13 0 8.17573e-20 $X=6.31 $Y=0.655
r113 37 43 37.6836 $w=2.75e-07 $l=2.15e-07 $layer=POLY_cond $X=6.02 $Y=0.49
+ $X2=5.805 $Y2=0.49
r114 36 39 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6.02 $Y=0.49 $X2=6.02
+ $Y2=0.69
r115 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.02
+ $Y=0.49 $X2=6.02 $Y2=0.49
r116 33 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=1.73
+ $X2=5.725 $Y2=1.565
r117 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=1.73 $X2=5.725 $Y2=1.73
r118 29 32 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=1.73
+ $X2=5.725 $Y2=1.73
r119 24 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=1.895
+ $X2=5.56 $Y2=1.73
r120 24 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.56 $Y=1.895
+ $X2=5.56 $Y2=2.035
r121 23 27 7.33333 $w=3.66e-07 $l=3.06855e-07 $layer=LI1_cond $X=4.71 $Y=0.69
+ $X2=4.502 $Y2=0.47
r122 22 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.855 $Y=0.69
+ $X2=6.02 $Y2=0.69
r123 22 23 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=5.855 $Y=0.69
+ $X2=4.71 $Y2=0.69
r124 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.475 $Y=2.12
+ $X2=5.56 $Y2=2.035
r125 20 21 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=5.475 $Y=2.12
+ $X2=4.295 $Y2=2.12
r126 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.13 $Y=2.205
+ $X2=4.295 $Y2=2.12
r127 16 18 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=4.13 $Y=2.205
+ $X2=4.13 $Y2=2.24
r128 13 37 50.8291 $w=2.75e-07 $l=3.63249e-07 $layer=POLY_cond $X=6.31 $Y=0.655
+ $X2=6.02 $Y2=0.49
r129 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.31 $Y=0.655
+ $X2=6.31 $Y2=0.975
r130 11 43 16.9318 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.805 $Y=0.655
+ $X2=5.805 $Y2=0.49
r131 11 42 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=5.805 $Y=0.655
+ $X2=5.805 $Y2=1.565
r132 7 33 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=1.895
+ $X2=5.725 $Y2=1.73
r133 7 9 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=5.725 $Y=1.895
+ $X2=5.725 $Y2=2.595
r134 2 18 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.98
+ $Y=2.095 $X2=4.13 $Y2=2.24
r135 1 27 182 $w=1.7e-07 $l=3.79737e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.235 $X2=4.46 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%RESET_B 3 7 9 10 17 18
c41 17 0 6.70955e-20 $X=6.5 $Y=1.77
c42 7 0 4.84139e-20 $X=6.67 $Y=0.975
r43 16 18 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=6.5 $Y=1.77 $X2=6.67
+ $Y2=1.77
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.5
+ $Y=1.77 $X2=6.5 $Y2=1.77
r45 13 16 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=6.255 $Y=1.77
+ $X2=6.5 $Y2=1.77
r46 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.5 $Y=2.035 $X2=6.5
+ $Y2=2.405
r47 9 17 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.5 $Y=2.035 $X2=6.5
+ $Y2=1.77
r48 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.67 $Y=1.605
+ $X2=6.67 $Y2=1.77
r49 5 7 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=6.67 $Y=1.605 $X2=6.67
+ $Y2=0.975
r50 1 13 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.935
+ $X2=6.255 $Y2=1.77
r51 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.255 $Y=1.935
+ $X2=6.255 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%A_1617_76# 1 2 9 13 17 23 26 28 31 35 40 43
+ 45 46
r66 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.32
+ $Y=1.165 $X2=9.32 $Y2=1.165
r67 40 42 10.6507 $w=3.43e-07 $l=2.3e-07 $layer=LI1_cond $X=8.232 $Y=0.59
+ $X2=8.232 $Y2=0.82
r68 36 43 3.35233 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=8.65 $Y=1.085
+ $X2=8.442 $Y2=1.085
r69 35 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.155 $Y=1.085
+ $X2=9.32 $Y2=1.085
r70 35 36 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=9.155 $Y=1.085
+ $X2=8.65 $Y2=1.085
r71 31 33 19.7165 $w=4.13e-07 $l=7.1e-07 $layer=LI1_cond $X=8.442 $Y=2.015
+ $X2=8.442 $Y2=2.725
r72 29 43 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=8.442 $Y=1.17
+ $X2=8.442 $Y2=1.085
r73 29 31 23.4654 $w=4.13e-07 $l=8.45e-07 $layer=LI1_cond $X=8.442 $Y=1.17
+ $X2=8.442 $Y2=2.015
r74 28 43 3.22182 $w=2.92e-07 $l=1.58915e-07 $layer=LI1_cond $X=8.32 $Y=1
+ $X2=8.442 $Y2=1.085
r75 28 42 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.32 $Y=1 $X2=8.32
+ $Y2=0.82
r76 25 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.32 $Y=1.505
+ $X2=9.32 $Y2=1.165
r77 25 26 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.32 $Y=1.505
+ $X2=9.32 $Y2=1.67
r78 22 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.32 $Y=1.15
+ $X2=9.32 $Y2=1.165
r79 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.32 $Y=1.075
+ $X2=9.59 $Y2=1.075
r80 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.23 $Y=1.075 $X2=9.32
+ $Y2=1.075
r81 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.59 $Y=1 $X2=9.59
+ $Y2=1.075
r82 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.59 $Y=1 $X2=9.59
+ $Y2=0.59
r83 13 26 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=9.28 $Y=2.37 $X2=9.28
+ $Y2=1.67
r84 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.23 $Y=1 $X2=9.23
+ $Y2=1.075
r85 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.23 $Y=1 $X2=9.23
+ $Y2=0.59
r86 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.34
+ $Y=1.87 $X2=8.485 $Y2=2.725
r87 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.34
+ $Y=1.87 $X2=8.485 $Y2=2.015
r88 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.085
+ $Y=0.38 $X2=8.225 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%VPWR 1 2 3 4 5 20 24 28 32 38 42 44 52 57
+ 65 72 73 76 79 82 85 88
c99 24 0 5.71049e-20 $X=3.1 $Y=2.57
r100 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r101 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r102 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 73 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r105 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r106 70 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.18 $Y=3.33
+ $X2=9.015 $Y2=3.33
r107 70 72 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=9.18 $Y=3.33
+ $X2=9.84 $Y2=3.33
r108 69 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r109 69 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 66 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.525 $Y=3.33
+ $X2=7.36 $Y2=3.33
r112 66 68 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.525 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 65 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.85 $Y=3.33
+ $X2=9.015 $Y2=3.33
r114 65 68 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=8.85 $Y=3.33
+ $X2=7.92 $Y2=3.33
r115 64 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 61 64 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 60 63 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r120 58 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.15 $Y2=3.33
r121 58 60 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.52 $Y2=3.33
r122 57 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.195 $Y=3.33
+ $X2=7.36 $Y2=3.33
r123 57 63 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.195 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 56 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r126 53 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.14 $Y2=3.33
r127 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.6 $Y2=3.33
r128 52 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=5.15 $Y2=3.33
r129 52 55 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r130 51 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r132 48 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 48 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 47 50 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 45 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.87 $Y2=3.33
r137 45 47 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 44 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.015 $Y=3.33
+ $X2=3.14 $Y2=3.33
r139 44 50 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.015 $Y=3.33
+ $X2=2.64 $Y2=3.33
r140 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r141 42 56 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r142 42 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r143 38 41 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.015 $Y=2.015
+ $X2=9.015 $Y2=2.725
r144 36 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.015 $Y=3.245
+ $X2=9.015 $Y2=3.33
r145 36 41 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=9.015 $Y=3.245
+ $X2=9.015 $Y2=2.725
r146 32 35 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.36 $Y=2.24
+ $X2=7.36 $Y2=2.95
r147 30 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=3.245
+ $X2=7.36 $Y2=3.33
r148 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.36 $Y=3.245
+ $X2=7.36 $Y2=2.95
r149 26 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=3.33
r150 26 28 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=2.55
r151 22 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=3.33
r152 22 24 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=2.57
r153 18 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=3.33
r154 18 20 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=2.83
r155 5 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.875
+ $Y=1.87 $X2=9.015 $Y2=2.725
r156 5 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.875
+ $Y=1.87 $X2=9.015 $Y2=2.015
r157 4 35 400 $w=1.7e-07 $l=1.34101e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.095 $X2=7.36 $Y2=2.95
r158 4 32 400 $w=1.7e-07 $l=1.05e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.095 $X2=7.36 $Y2=2.24
r159 3 28 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=5.01
+ $Y=2.095 $X2=5.15 $Y2=2.55
r160 2 24 300 $w=1.7e-07 $l=6.10635e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=2.095 $X2=3.1 $Y2=2.57
r161 1 20 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=1.98 $X2=0.87 $Y2=2.83
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%Q 1 2 9 13 14 15 16 17 18
r28 17 18 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.88 $Y=2.405
+ $X2=7.88 $Y2=2.775
r29 17 31 5.43295 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.88 $Y=2.405
+ $X2=7.88 $Y2=2.24
r30 16 31 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=7.88 $Y=2.035
+ $X2=7.88 $Y2=2.24
r31 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.88 $Y=1.665
+ $X2=7.88 $Y2=2.035
r32 14 15 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.88 $Y=1.295
+ $X2=7.88 $Y2=1.665
r33 13 14 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=7.88 $Y=1.205 $X2=7.88
+ $Y2=1.295
r34 12 13 0.789345 $w=3.63e-07 $l=2.5e-08 $layer=LI1_cond $X=7.782 $Y=1.18
+ $X2=7.782 $Y2=1.205
r35 9 12 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=7.692 $Y=0.975
+ $X2=7.692 $Y2=1.18
r36 2 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.75
+ $Y=2.095 $X2=7.89 $Y2=2.24
r37 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.535
+ $Y=0.765 $X2=7.675 $Y2=0.975
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%Q_N 1 2 10 13 14 15 28 29
r23 28 29 10.0909 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=9.675 $Y=2.015
+ $X2=9.675 $Y2=1.85
r24 15 23 1.01363 $w=5.88e-07 $l=5e-08 $layer=LI1_cond $X=9.675 $Y=2.775
+ $X2=9.675 $Y2=2.725
r25 14 23 6.48721 $w=5.88e-07 $l=3.2e-07 $layer=LI1_cond $X=9.675 $Y=2.405
+ $X2=9.675 $Y2=2.725
r26 14 19 5.27085 $w=5.88e-07 $l=2.6e-07 $layer=LI1_cond $X=9.675 $Y=2.405
+ $X2=9.675 $Y2=2.145
r27 13 19 2.22998 $w=5.88e-07 $l=1.1e-07 $layer=LI1_cond $X=9.675 $Y=2.035
+ $X2=9.675 $Y2=2.145
r28 13 28 0.40545 $w=5.88e-07 $l=2e-08 $layer=LI1_cond $X=9.675 $Y=2.035
+ $X2=9.675 $Y2=2.015
r29 12 29 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=9.885 $Y=0.82
+ $X2=9.885 $Y2=1.85
r30 10 12 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=9.805 $Y=0.59
+ $X2=9.805 $Y2=0.82
r31 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.405
+ $Y=1.87 $X2=9.545 $Y2=2.015
r32 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.405
+ $Y=1.87 $X2=9.545 $Y2=2.725
r33 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.665
+ $Y=0.38 $X2=9.805 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_LP%VGND 1 2 3 4 5 18 20 24 28 32 36 38 40 45
+ 53 58 65 66 69 72 75 78 81
r119 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r120 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r121 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r122 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r123 70 73 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r124 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r125 66 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=8.88
+ $Y2=0
r126 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r127 63 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.18 $Y=0 $X2=9.015
+ $Y2=0
r128 63 65 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=9.18 $Y=0 $X2=9.84
+ $Y2=0
r129 62 82 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.88 $Y2=0
r130 62 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r131 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r132 59 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.05 $Y=0 $X2=6.885
+ $Y2=0
r133 59 61 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.05 $Y=0 $X2=7.44
+ $Y2=0
r134 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.85 $Y=0 $X2=9.015
+ $Y2=0
r135 58 61 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=8.85 $Y=0 $X2=7.44
+ $Y2=0
r136 57 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r137 57 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=5.52
+ $Y2=0
r138 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r139 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=0 $X2=5.51
+ $Y2=0
r140 54 56 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=5.675 $Y=0
+ $X2=6.48 $Y2=0
r141 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.72 $Y=0 $X2=6.885
+ $Y2=0
r142 53 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.72 $Y=0 $X2=6.48
+ $Y2=0
r143 49 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r144 48 51 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r145 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 46 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.21
+ $Y2=0
r147 46 48 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.6
+ $Y2=0
r148 45 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.345 $Y=0 $X2=5.51
+ $Y2=0
r149 45 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.04 $Y2=0
r150 43 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r151 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r152 40 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r153 40 42 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r154 38 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r155 38 49 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r156 38 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r157 34 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.015 $Y=0.085
+ $X2=9.015 $Y2=0
r158 34 36 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=9.015 $Y=0.085
+ $X2=9.015 $Y2=0.59
r159 30 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.885 $Y=0.085
+ $X2=6.885 $Y2=0
r160 30 32 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=6.885 $Y=0.085
+ $X2=6.885 $Y2=0.91
r161 26 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=0.085
+ $X2=5.51 $Y2=0
r162 26 28 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.51 $Y=0.085
+ $X2=5.51 $Y2=0.34
r163 22 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r164 22 24 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.445
r165 21 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r166 20 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.21
+ $Y2=0
r167 20 21 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=3.045 $Y=0
+ $X2=1.235 $Y2=0
r168 16 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r169 16 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.55
r170 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.875
+ $Y=0.38 $X2=9.015 $Y2=0.59
r171 4 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.745
+ $Y=0.765 $X2=6.885 $Y2=0.91
r172 3 28 182 $w=1.7e-07 $l=2.67395e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.235 $X2=5.51 $Y2=0.34
r173 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.235 $X2=3.21 $Y2=0.445
r174 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.34 $X2=1.07 $Y2=0.55
.ends

