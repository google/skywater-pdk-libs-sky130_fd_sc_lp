* File: sky130_fd_sc_lp__dlrbp_lp.spice
* Created: Fri Aug 28 10:26:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dlrbp_lp  VNB VPB D GATE RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1014 A_114_112# N_D_M1014_g N_A_27_112#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_D_M1006_g A_114_112# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1008 A_272_112# N_GATE_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_272_419#_M1000_d N_GATE_M1000_g A_272_112# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 A_542_49# N_A_272_419#_M1016_g N_A_455_49#_M1016_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_272_419#_M1010_g A_542_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1018 A_700_49# N_A_27_112#_M1018_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1026 N_A_778_49#_M1026_d N_A_455_49#_M1026_g A_700_49# VNB NSHORT L=0.15
+ W=0.42 AD=0.1428 AS=0.0504 PD=1.1 PS=0.66 NRD=101.424 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1019 A_944_49# N_A_272_419#_M1019_g N_A_778_49#_M1026_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.1428 PD=0.84 PS=1.1 NRD=44.28 NRS=12.852 M=1 R=2.8
+ SA=75002.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_1028_23#_M1028_g A_944_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.1554 AS=0.0882 PD=1.58 PS=0.84 NRD=24.276 NRS=44.28 M=1 R=2.8 SA=75002.8
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1020 A_1273_49# N_A_778_49#_M1020_g N_A_1028_23#_M1020_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_RESET_B_M1023_g A_1273_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_1431_49# N_A_1028_23#_M1005_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_Q_M1024_d N_A_1028_23#_M1024_g A_1431_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 A_1701_74# N_A_1028_23#_M1029_g N_A_1614_74#_M1029_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1028_23#_M1001_g A_1701_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1017 A_1859_74# N_A_1614_74#_M1017_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_Q_N_M1012_d N_A_1614_74#_M1012_g A_1859_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_D_M1027_g N_A_27_112#_M1027_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1013 N_A_272_419#_M1013_d N_GATE_M1013_g N_VPWR_M1027_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1011 N_VPWR_M1011_d N_A_272_419#_M1011_g N_A_455_49#_M1011_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.194 AS=0.285 PD=1.52 PS=2.57 NRD=16.7253 NRS=0 M=1 R=4
+ SA=125000 SB=125004 A=0.25 P=2.5 MULT=1
MM1025 A_692_367# N_A_27_112#_M1025_g N_VPWR_M1011_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.194 PD=1.24 PS=1.52 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1007 N_A_778_49#_M1007_d N_A_272_419#_M1007_g A_692_367# VPB PHIGHVT L=0.25
+ W=1 AD=0.2875 AS=0.12 PD=1.575 PS=1.24 NRD=50.2153 NRS=12.7853 M=1 R=4
+ SA=125001 SB=125003 A=0.25 P=2.5 MULT=1
MM1009 A_955_367# N_A_455_49#_M1009_g N_A_778_49#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1825 AS=0.2875 PD=1.365 PS=1.575 NRD=25.0978 NRS=7.8603 M=1 R=4 SA=125002
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_A_1028_23#_M1002_g A_955_367# VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.1825 PD=1.32 PS=1.365 NRD=0 NRS=25.0978 M=1 R=4 SA=125003
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1021 N_A_1028_23#_M1021_d N_A_778_49#_M1021_g N_VPWR_M1002_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.2345 AS=0.16 PD=1.54 PS=1.32 NRD=16.0752 NRS=7.8603 M=1 R=4
+ SA=125003 SB=125001 A=0.25 P=2.5 MULT=1
MM1015 N_VPWR_M1015_d N_RESET_B_M1015_g N_A_1028_23#_M1021_d VPB PHIGHVT L=0.25
+ W=1 AD=0.1425 AS=0.2345 PD=1.285 PS=1.54 NRD=0 NRS=16.0752 M=1 R=4 SA=125004
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1003 N_Q_M1003_d N_A_1028_23#_M1003_g N_VPWR_M1015_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1425 PD=2.57 PS=1.285 NRD=0 NRS=0.9653 M=1 R=4 SA=125004
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_1028_23#_M1004_g N_A_1614_74#_M1004_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1022 N_Q_N_M1022_d N_A_1614_74#_M1022_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX30_noxref VNB VPB NWDIODE A=20.3903 P=24.97
*
.include "sky130_fd_sc_lp__dlrbp_lp.pxi.spice"
*
.ends
*
*
