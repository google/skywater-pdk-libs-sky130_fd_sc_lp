# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ha_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__ha_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.075000 1.345000 4.715000 1.675000 ;
        RECT 4.545000 1.675000 4.715000 1.695000 ;
        RECT 4.545000 1.695000 7.375000 1.750000 ;
        RECT 4.545000 1.750000 6.120000 1.875000 ;
        RECT 5.440000 1.425000 5.770000 1.580000 ;
        RECT 5.440000 1.580000 7.375000 1.695000 ;
        RECT 6.875000 1.425000 7.375000 1.580000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.895000 1.345000 5.260000 1.515000 ;
        RECT 5.090000 1.085000 7.725000 1.255000 ;
        RECT 5.090000 1.255000 5.260000 1.345000 ;
        RECT 5.980000 1.255000 6.310000 1.345000 ;
        RECT 7.555000 1.255000 7.725000 1.345000 ;
        RECT 7.555000 1.345000 8.425000 1.515000 ;
        RECT 7.835000 1.515000 8.425000 1.750000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 1.045000 3.550000 1.215000 ;
        RECT 2.425000 1.215000 2.595000 1.755000 ;
        RECT 2.425000 1.755000 3.515000 1.925000 ;
        RECT 2.425000 1.925000 2.725000 3.075000 ;
        RECT 2.500000 0.255000 2.690000 1.045000 ;
        RECT 3.280000 1.925000 3.515000 3.075000 ;
        RECT 3.360000 0.255000 3.550000 1.045000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.045000 1.830000 1.215000 ;
        RECT 0.090000 1.215000 0.405000 1.755000 ;
        RECT 0.090000 1.755000 1.830000 1.925000 ;
        RECT 0.745000 1.925000 0.935000 3.075000 ;
        RECT 0.780000 0.255000 0.970000 1.045000 ;
        RECT 1.605000 1.925000 1.830000 3.075000 ;
        RECT 1.640000 0.255000 1.830000 1.045000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.245000  2.095000  0.575000 3.245000 ;
      RECT 0.280000  0.085000  0.610000 0.875000 ;
      RECT 0.675000  1.395000  2.245000 1.565000 ;
      RECT 1.105000  2.095000  1.435000 3.245000 ;
      RECT 1.140000  0.085000  1.470000 0.865000 ;
      RECT 2.000000  0.085000  2.330000 0.670000 ;
      RECT 2.000000  1.810000  2.255000 3.245000 ;
      RECT 2.075000  0.840000  2.245000 1.395000 ;
      RECT 2.775000  1.395000  3.890000 1.565000 ;
      RECT 2.860000  0.085000  3.190000 0.865000 ;
      RECT 2.895000  2.095000  3.110000 3.245000 ;
      RECT 3.685000  2.195000  4.015000 3.245000 ;
      RECT 3.720000  0.085000  4.060000 0.805000 ;
      RECT 3.720000  0.995000  4.920000 1.165000 ;
      RECT 3.720000  1.165000  3.890000 1.395000 ;
      RECT 3.720000  1.565000  3.890000 1.855000 ;
      RECT 3.720000  1.855000  4.365000 2.025000 ;
      RECT 4.195000  2.025000  4.365000 2.045000 ;
      RECT 4.195000  2.045000  8.775000 2.100000 ;
      RECT 4.195000  2.100000  6.470000 2.215000 ;
      RECT 4.195000  2.215000  4.510000 3.055000 ;
      RECT 4.230000  0.265000  5.435000 0.435000 ;
      RECT 4.230000  0.435000  4.560000 0.815000 ;
      RECT 4.680000  2.385000  5.010000 3.245000 ;
      RECT 4.730000  0.605000  4.920000 0.995000 ;
      RECT 5.105000  0.435000  5.435000 0.825000 ;
      RECT 5.180000  2.215000  5.390000 3.075000 ;
      RECT 5.560000  2.385000  5.890000 3.245000 ;
      RECT 5.605000  0.085000  5.890000 0.915000 ;
      RECT 6.300000  1.930000  8.775000 2.045000 ;
      RECT 6.380000  0.365000  6.710000 0.725000 ;
      RECT 6.380000  0.725000  7.660000 0.735000 ;
      RECT 6.380000  0.735000  8.075000 0.915000 ;
      RECT 6.380000  2.395000  9.125000 2.440000 ;
      RECT 6.380000  2.440000  6.820000 2.565000 ;
      RECT 6.380000  2.565000  6.640000 3.075000 ;
      RECT 6.650000  2.270000  9.125000 2.395000 ;
      RECT 6.810000  2.745000  8.270000 2.780000 ;
      RECT 6.810000  2.780000  7.170000 2.955000 ;
      RECT 6.890000  0.085000  7.220000 0.535000 ;
      RECT 7.000000  2.610000  8.270000 2.745000 ;
      RECT 7.340000  2.950000  7.685000 3.245000 ;
      RECT 7.400000  0.285000  7.660000 0.725000 ;
      RECT 7.830000  0.085000  8.445000 0.565000 ;
      RECT 7.905000  0.915000  8.075000 0.925000 ;
      RECT 7.905000  0.925000  8.855000 1.095000 ;
      RECT 7.940000  2.780000  8.270000 2.960000 ;
      RECT 8.245000  0.565000  8.445000 0.755000 ;
      RECT 8.450000  2.440000  9.125000 2.450000 ;
      RECT 8.450000  2.450000  8.780000 3.075000 ;
      RECT 8.605000  1.405000  9.170000 1.575000 ;
      RECT 8.605000  1.575000  8.775000 1.930000 ;
      RECT 8.665000  0.265000  9.930000 0.435000 ;
      RECT 8.665000  0.435000  8.855000 0.925000 ;
      RECT 8.950000  2.630000  9.520000 3.245000 ;
      RECT 8.955000  1.755000  9.985000 1.925000 ;
      RECT 8.955000  1.925000  9.125000 2.270000 ;
      RECT 9.035000  0.615000  9.510000 1.145000 ;
      RECT 9.295000  2.105000  9.520000 2.630000 ;
      RECT 9.340000  1.145000  9.510000 1.755000 ;
      RECT 9.680000  0.435000  9.930000 1.185000 ;
      RECT 9.690000  1.925000  9.985000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  0.840000 9.445000 1.010000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 0.810000 2.305000 0.855000 ;
      RECT 2.015000 0.855000 9.505000 0.995000 ;
      RECT 2.015000 0.995000 2.305000 1.040000 ;
      RECT 9.215000 0.810000 9.505000 0.855000 ;
      RECT 9.215000 0.995000 9.505000 1.040000 ;
  END
END sky130_fd_sc_lp__ha_4
END LIBRARY
