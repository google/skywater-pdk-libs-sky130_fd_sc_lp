* File: sky130_fd_sc_lp__a21oi_lp.pxi.spice
* Created: Wed Sep  2 09:20:51 2020
* 
x_PM_SKY130_FD_SC_LP__A21OI_LP%A2 N_A2_c_48_n N_A2_c_54_n N_A2_M1005_g
+ N_A2_M1002_g N_A2_c_50_n N_A2_c_51_n A2 N_A2_c_52_n N_A2_c_53_n
+ PM_SKY130_FD_SC_LP__A21OI_LP%A2
x_PM_SKY130_FD_SC_LP__A21OI_LP%A1 N_A1_M1006_g N_A1_M1001_g N_A1_c_87_n
+ N_A1_c_88_n A1 N_A1_c_90_n PM_SKY130_FD_SC_LP__A21OI_LP%A1
x_PM_SKY130_FD_SC_LP__A21OI_LP%B1 N_B1_M1003_g N_B1_M1000_g N_B1_M1004_g B1
+ N_B1_c_130_n PM_SKY130_FD_SC_LP__A21OI_LP%B1
x_PM_SKY130_FD_SC_LP__A21OI_LP%A_31_409# N_A_31_409#_M1005_s N_A_31_409#_M1001_d
+ N_A_31_409#_c_167_n N_A_31_409#_c_168_n N_A_31_409#_c_169_n
+ N_A_31_409#_c_170_n PM_SKY130_FD_SC_LP__A21OI_LP%A_31_409#
x_PM_SKY130_FD_SC_LP__A21OI_LP%VPWR N_VPWR_M1005_d N_VPWR_c_200_n VPWR
+ N_VPWR_c_201_n N_VPWR_c_199_n N_VPWR_c_203_n PM_SKY130_FD_SC_LP__A21OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A21OI_LP%Y N_Y_M1006_d N_Y_M1000_d N_Y_c_223_n N_Y_c_224_n
+ Y Y Y Y Y Y N_Y_c_226_n Y Y PM_SKY130_FD_SC_LP__A21OI_LP%Y
x_PM_SKY130_FD_SC_LP__A21OI_LP%VGND N_VGND_M1002_s N_VGND_M1004_d N_VGND_c_266_n
+ N_VGND_c_267_n N_VGND_c_268_n N_VGND_c_269_n VGND N_VGND_c_270_n
+ N_VGND_c_271_n PM_SKY130_FD_SC_LP__A21OI_LP%VGND
cc_1 VNB N_A2_c_48_n 0.0212633f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.305
cc_2 VNB N_A2_M1002_g 0.0279149f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_3 VNB N_A2_c_50_n 0.0283125f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.525
cc_4 VNB N_A2_c_51_n 0.0107227f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.765
cc_5 VNB N_A2_c_52_n 0.028108f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.02
cc_6 VNB N_A2_c_53_n 0.0290358f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.02
cc_7 VNB N_A1_M1006_g 0.0351259f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.525
cc_8 VNB N_A1_c_87_n 0.0198243f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_9 VNB N_A1_c_88_n 0.00458524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A1 0.00954574f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.525
cc_11 VNB N_A1_c_90_n 0.0176475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_M1003_g 0.0315368f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.525
cc_13 VNB N_B1_M1004_g 0.0360067f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_14 VNB B1 2.87194e-19 $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.525
cc_15 VNB N_B1_c_130_n 0.0568203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_199_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.02
cc_17 VNB N_Y_c_223_n 0.0010022f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.855
cc_18 VNB N_Y_c_224_n 0.0100728f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_19 VNB Y 0.00905392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_226_n 0.0094116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB Y 0.0371346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_266_n 0.0138745f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.545
cc_23 VNB N_VGND_c_267_n 0.0213411f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.855
cc_24 VNB N_VGND_c_268_n 0.0109752f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_25 VNB N_VGND_c_269_n 0.0148317f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.525
cc_26 VNB N_VGND_c_270_n 0.0382869f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.02
cc_27 VNB N_VGND_c_271_n 0.150585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A2_c_54_n 0.0147112f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.89
cc_29 VPB N_A2_M1005_g 0.0294926f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.545
cc_30 VPB N_A2_c_51_n 0.00909031f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.765
cc_31 VPB N_A1_M1001_g 0.0335111f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.545
cc_32 VPB N_A1_c_88_n 0.00758005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB A1 0.00242956f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.525
cc_34 VPB N_B1_M1000_g 0.0392486f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.545
cc_35 VPB B1 8.39373e-19 $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.525
cc_36 VPB N_B1_c_130_n 0.015854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_31_409#_c_167_n 0.0391242f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.855
cc_38 VPB N_A_31_409#_c_168_n 0.0151311f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.525
cc_39 VPB N_A_31_409#_c_169_n 0.0107391f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.765
cc_40 VPB N_A_31_409#_c_170_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.02
cc_41 VPB N_VPWR_c_200_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_201_n 0.0380539f $X=-0.19 $Y=1.655 $X2=0.44 $Y2=1.02
cc_43 VPB N_VPWR_c_199_n 0.0550536f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.02
cc_44 VPB N_VPWR_c_203_n 0.0245402f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.19
cc_45 VPB Y 0.0410226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB Y 0.0192317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB Y 0.0197913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 N_A2_M1002_g N_A1_M1006_g 0.0255934f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_49 N_A2_c_53_n N_A1_M1006_g 0.00103847f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_50 N_A2_c_54_n N_A1_M1001_g 0.0323667f $X=0.565 $Y=1.89 $X2=0 $Y2=0
cc_51 N_A2_c_51_n N_A1_M1001_g 7.61622e-19 $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_52 N_A2_c_48_n N_A1_c_87_n 0.0255934f $X=0.44 $Y=1.305 $X2=0 $Y2=0
cc_53 N_A2_c_51_n N_A1_c_87_n 0.00804429f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_54 N_A2_c_48_n A1 0.0018594f $X=0.44 $Y=1.305 $X2=0 $Y2=0
cc_55 N_A2_c_51_n A1 0.00133377f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A2_c_53_n A1 0.0196065f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_57 N_A2_c_52_n N_A1_c_90_n 0.0255934f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_58 N_A2_c_53_n N_A1_c_90_n 4.84182e-19 $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_59 N_A2_M1005_g N_A_31_409#_c_167_n 0.0174312f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_60 N_A2_M1005_g N_A_31_409#_c_168_n 0.0205163f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_61 N_A2_c_50_n N_A_31_409#_c_168_n 3.8461e-19 $X=0.44 $Y=1.525 $X2=0 $Y2=0
cc_62 N_A2_c_53_n N_A_31_409#_c_168_n 0.00321236f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_63 N_A2_M1005_g N_A_31_409#_c_169_n 0.00338134f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_64 N_A2_c_50_n N_A_31_409#_c_169_n 0.00505179f $X=0.44 $Y=1.525 $X2=0 $Y2=0
cc_65 N_A2_c_53_n N_A_31_409#_c_169_n 0.0157182f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_66 N_A2_M1005_g N_A_31_409#_c_170_n 9.43535e-19 $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_67 N_A2_M1005_g N_VPWR_c_200_n 0.0199441f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_68 N_A2_M1005_g N_VPWR_c_199_n 0.014097f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_69 N_A2_M1005_g N_VPWR_c_203_n 0.00769046f $X=0.565 $Y=2.545 $X2=0 $Y2=0
cc_70 N_A2_c_53_n N_Y_c_224_n 0.0012559f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_71 N_A2_M1002_g N_VGND_c_267_n 0.0154869f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A2_c_52_n N_VGND_c_267_n 0.00776823f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_73 N_A2_c_53_n N_VGND_c_267_n 0.0270777f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_74 N_A2_M1002_g N_VGND_c_270_n 0.00486043f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A2_M1002_g N_VGND_c_271_n 0.00780343f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A2_c_53_n N_VGND_c_271_n 0.00472631f $X=0.385 $Y=1.02 $X2=0 $Y2=0
cc_77 N_A1_M1006_g N_B1_M1003_g 0.0207188f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_78 N_A1_M1001_g N_B1_M1000_g 0.0217656f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_79 A1 B1 0.0518188f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A1_c_90_n B1 6.91441e-19 $X=1.065 $Y=1.24 $X2=0 $Y2=0
cc_81 A1 N_B1_c_130_n 0.00459954f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A1_c_90_n N_B1_c_130_n 0.0363231f $X=1.065 $Y=1.24 $X2=0 $Y2=0
cc_83 N_A1_M1001_g N_A_31_409#_c_167_n 9.43535e-19 $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A1_M1001_g N_A_31_409#_c_168_n 0.0200288f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_85 N_A1_c_88_n N_A_31_409#_c_168_n 0.00209912f $X=1.065 $Y=1.745 $X2=0 $Y2=0
cc_86 A1 N_A_31_409#_c_168_n 0.0320267f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A1_M1001_g N_A_31_409#_c_170_n 0.0172711f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_88 N_A1_M1001_g N_VPWR_c_200_n 0.0188592f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_89 N_A1_M1001_g N_VPWR_c_201_n 0.00769046f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_90 N_A1_M1001_g N_VPWR_c_199_n 0.0134474f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_91 N_A1_M1006_g N_Y_c_223_n 0.00707393f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A1_M1006_g N_Y_c_224_n 0.00466564f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_93 A1 N_Y_c_224_n 0.0130477f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A1_c_90_n N_Y_c_224_n 0.00175043f $X=1.065 $Y=1.24 $X2=0 $Y2=0
cc_95 N_A1_M1001_g Y 2.75256e-19 $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_96 N_A1_M1006_g N_VGND_c_267_n 0.00247402f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A1_M1006_g N_VGND_c_270_n 0.00585385f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A1_M1006_g N_VGND_c_271_n 0.0112502f $X=0.975 $Y=0.445 $X2=0 $Y2=0
cc_99 N_B1_M1000_g N_A_31_409#_c_168_n 0.00525764f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_100 B1 N_A_31_409#_c_168_n 0.00235924f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B1_c_130_n N_A_31_409#_c_168_n 0.00124451f $X=1.66 $Y=1.24 $X2=0 $Y2=0
cc_102 N_B1_M1000_g N_A_31_409#_c_170_n 0.0173747f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_103 N_B1_M1000_g N_VPWR_c_200_n 8.7471e-19 $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_104 N_B1_M1000_g N_VPWR_c_201_n 0.00826654f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_105 N_B1_M1000_g N_VPWR_c_199_n 0.0156484f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_106 N_B1_M1003_g N_Y_c_223_n 0.00881509f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_107 N_B1_M1004_g N_Y_c_223_n 0.00166179f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B1_M1003_g N_Y_c_224_n 0.00390232f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_109 N_B1_M1003_g Y 0.00834974f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_110 N_B1_M1004_g Y 0.017381f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_111 B1 Y 0.0246023f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B1_c_130_n Y 2.06137e-19 $X=1.66 $Y=1.24 $X2=0 $Y2=0
cc_113 N_B1_M1000_g Y 0.0136661f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_114 N_B1_M1000_g Y 0.00771081f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_115 N_B1_M1004_g Y 0.0255355f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_116 B1 Y 0.0382076f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_M1000_g Y 0.00558148f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_118 B1 Y 0.00588764f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B1_c_130_n Y 0.00725566f $X=1.66 $Y=1.24 $X2=0 $Y2=0
cc_120 N_B1_M1003_g N_VGND_c_269_n 0.0020441f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_121 N_B1_M1004_g N_VGND_c_269_n 0.0112017f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_122 N_B1_M1003_g N_VGND_c_270_n 0.00426341f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B1_M1004_g N_VGND_c_270_n 0.00364083f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_124 N_B1_M1003_g N_VGND_c_271_n 0.00623968f $X=1.545 $Y=0.445 $X2=0 $Y2=0
cc_125 N_B1_M1004_g N_VGND_c_271_n 0.00416707f $X=1.905 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_31_409#_c_168_n N_VPWR_M1005_d 0.00180746f $X=1.195 $Y=2.01 $X2=-0.19
+ $Y2=1.655
cc_127 N_A_31_409#_c_167_n N_VPWR_c_200_n 0.0520536f $X=0.3 $Y=2.19 $X2=0 $Y2=0
cc_128 N_A_31_409#_c_168_n N_VPWR_c_200_n 0.0163515f $X=1.195 $Y=2.01 $X2=0
+ $Y2=0
cc_129 N_A_31_409#_c_170_n N_VPWR_c_200_n 0.0520536f $X=1.36 $Y=2.19 $X2=0 $Y2=0
cc_130 N_A_31_409#_c_170_n N_VPWR_c_201_n 0.021949f $X=1.36 $Y=2.19 $X2=0 $Y2=0
cc_131 N_A_31_409#_c_167_n N_VPWR_c_199_n 0.0125808f $X=0.3 $Y=2.19 $X2=0 $Y2=0
cc_132 N_A_31_409#_c_170_n N_VPWR_c_199_n 0.0124703f $X=1.36 $Y=2.19 $X2=0 $Y2=0
cc_133 N_A_31_409#_c_167_n N_VPWR_c_203_n 0.0220321f $X=0.3 $Y=2.19 $X2=0 $Y2=0
cc_134 N_A_31_409#_c_168_n Y 0.00328883f $X=1.195 $Y=2.01 $X2=0 $Y2=0
cc_135 N_A_31_409#_c_168_n Y 0.00509062f $X=1.195 $Y=2.01 $X2=0 $Y2=0
cc_136 N_A_31_409#_c_170_n Y 0.0664415f $X=1.36 $Y=2.19 $X2=0 $Y2=0
cc_137 N_VPWR_c_201_n Y 0.0368655f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_138 N_VPWR_c_199_n Y 0.0210933f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_139 N_Y_c_223_n N_VGND_c_267_n 0.0113057f $X=1.33 $Y=0.47 $X2=0 $Y2=0
cc_140 N_Y_c_223_n N_VGND_c_269_n 0.00936806f $X=1.33 $Y=0.47 $X2=0 $Y2=0
cc_141 Y N_VGND_c_269_n 0.00636087f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_142 N_Y_c_226_n N_VGND_c_269_n 0.0167824f $X=2.175 $Y=0.895 $X2=0 $Y2=0
cc_143 N_Y_c_223_n N_VGND_c_270_n 0.0196636f $X=1.33 $Y=0.47 $X2=0 $Y2=0
cc_144 Y N_VGND_c_270_n 0.00652017f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_145 N_Y_M1006_d N_VGND_c_271_n 0.00743588f $X=1.05 $Y=0.235 $X2=0 $Y2=0
cc_146 N_Y_c_223_n N_VGND_c_271_n 0.0125545f $X=1.33 $Y=0.47 $X2=0 $Y2=0
cc_147 Y N_VGND_c_271_n 0.0114914f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_148 N_Y_c_226_n N_VGND_c_271_n 8.95026e-19 $X=2.175 $Y=0.895 $X2=0 $Y2=0
cc_149 N_VGND_c_271_n A_132_47# 0.010279f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_150 N_VGND_c_271_n A_324_47# 0.00271994f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
