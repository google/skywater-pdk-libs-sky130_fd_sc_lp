# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a221o_0
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a221o_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.540000 0.840000 1.845000 1.605000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.900000 1.065000 1.360000 1.615000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 0.840000 2.270000 1.510000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 1.050000 2.840000 1.585000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 0.995000 3.755000 1.665000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.280000 0.535000 0.555000 ;
        RECT 0.090000 0.555000 0.335000 1.390000 ;
        RECT 0.090000 1.390000 0.270000 2.400000 ;
        RECT 0.090000 2.400000 0.475000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.440000  1.560000 0.675000 2.230000 ;
      RECT 0.505000  0.725000 1.370000 0.895000 ;
      RECT 0.505000  0.895000 0.675000 1.560000 ;
      RECT 0.645000  2.400000 0.925000 3.245000 ;
      RECT 0.715000  0.085000 1.030000 0.555000 ;
      RECT 1.095000  1.785000 2.785000 1.955000 ;
      RECT 1.095000  1.955000 1.350000 3.075000 ;
      RECT 1.200000  0.280000 2.610000 0.610000 ;
      RECT 1.200000  0.610000 1.370000 0.725000 ;
      RECT 1.520000  2.400000 1.815000 3.245000 ;
      RECT 2.005000  2.135000 2.285000 2.905000 ;
      RECT 2.005000  2.905000 3.285000 3.075000 ;
      RECT 2.440000  0.610000 2.610000 0.645000 ;
      RECT 2.440000  0.645000 3.575000 0.815000 ;
      RECT 2.455000  1.955000 2.785000 2.735000 ;
      RECT 2.780000  0.085000 3.110000 0.475000 ;
      RECT 2.955000  2.185000 3.285000 2.905000 ;
      RECT 3.010000  0.815000 3.190000 1.845000 ;
      RECT 3.010000  1.845000 3.715000 2.015000 ;
      RECT 3.280000  0.280000 3.575000 0.645000 ;
      RECT 3.455000  2.015000 3.715000 2.795000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__a221o_0
