* NGSPICE file created from sky130_fd_sc_lp__xnor2_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__xnor2_lp A B VGND VNB VPB VPWR Y
M1000 Y a_82_66# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=8.4e+11p ps=7.68e+06u
M1001 a_112_92# B VGND VNB nshort w=420000u l=150000u
+  ad=3.003e+11p pd=3.11e+06u as=2.331e+11p ps=2.79e+06u
M1002 VPWR A a_280_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1003 VPWR B a_82_66# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1004 VGND A a_112_92# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_510_125# A VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1006 a_280_419# B Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_82_66# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_82_66# B a_510_125# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1009 a_112_92# a_82_66# Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
.ends

