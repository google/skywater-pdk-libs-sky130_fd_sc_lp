# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a211o_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a211o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 1.195000 2.470000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.195000 1.845000 1.525000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 1.195000 3.215000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.195000 3.755000 1.515000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.255000 0.825000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.095000  0.085000 0.385000 1.095000 ;
      RECT 0.095000  1.815000 0.385000 3.245000 ;
      RECT 0.995000  0.085000 1.805000 0.685000 ;
      RECT 1.000000  1.345000 1.415000 1.675000 ;
      RECT 1.000000  2.045000 1.285000 3.245000 ;
      RECT 1.245000  0.855000 3.675000 1.025000 ;
      RECT 1.245000  1.025000 1.415000 1.345000 ;
      RECT 1.245000  1.675000 1.415000 1.695000 ;
      RECT 1.245000  1.695000 3.675000 1.875000 ;
      RECT 1.475000  2.045000 2.790000 2.225000 ;
      RECT 1.475000  2.225000 1.790000 3.075000 ;
      RECT 1.960000  2.395000 2.290000 3.245000 ;
      RECT 2.365000  0.255000 2.695000 0.855000 ;
      RECT 2.460000  2.225000 2.790000 3.065000 ;
      RECT 2.915000  0.085000 3.245000 0.685000 ;
      RECT 3.345000  1.875000 3.675000 3.075000 ;
      RECT 3.415000  0.255000 3.675000 0.855000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__a211o_2
END LIBRARY
