* File: sky130_fd_sc_lp__a41oi_2.pxi.spice
* Created: Wed Sep  2 09:29:41 2020
* 
x_PM_SKY130_FD_SC_LP__A41OI_2%B1 N_B1_c_94_n N_B1_M1011_g N_B1_M1001_g
+ N_B1_c_96_n N_B1_M1012_g N_B1_M1007_g B1 B1 N_B1_c_99_n
+ PM_SKY130_FD_SC_LP__A41OI_2%B1
x_PM_SKY130_FD_SC_LP__A41OI_2%A1 N_A1_M1000_g N_A1_c_140_n N_A1_M1004_g
+ N_A1_M1015_g N_A1_c_142_n N_A1_M1016_g A1 A1 N_A1_c_143_n N_A1_c_144_n
+ PM_SKY130_FD_SC_LP__A41OI_2%A1
x_PM_SKY130_FD_SC_LP__A41OI_2%A2 N_A2_M1010_g N_A2_M1002_g N_A2_M1014_g
+ N_A2_M1018_g N_A2_c_201_n N_A2_c_202_n A2 A2 PM_SKY130_FD_SC_LP__A41OI_2%A2
x_PM_SKY130_FD_SC_LP__A41OI_2%A3 N_A3_M1006_g N_A3_c_253_n N_A3_M1005_g
+ N_A3_c_254_n N_A3_M1017_g N_A3_M1008_g N_A3_c_256_n A3 N_A3_c_258_n
+ PM_SKY130_FD_SC_LP__A41OI_2%A3
x_PM_SKY130_FD_SC_LP__A41OI_2%A4 N_A4_M1009_g N_A4_M1003_g N_A4_M1019_g
+ N_A4_M1013_g A4 A4 N_A4_c_318_n PM_SKY130_FD_SC_LP__A41OI_2%A4
x_PM_SKY130_FD_SC_LP__A41OI_2%A_103_367# N_A_103_367#_M1001_d
+ N_A_103_367#_M1007_d N_A_103_367#_M1015_d N_A_103_367#_M1018_s
+ N_A_103_367#_M1008_s N_A_103_367#_M1013_s N_A_103_367#_c_356_n
+ N_A_103_367#_c_357_n N_A_103_367#_c_365_n N_A_103_367#_c_368_n
+ N_A_103_367#_c_367_n N_A_103_367#_c_371_n N_A_103_367#_c_374_n
+ N_A_103_367#_c_378_n N_A_103_367#_c_385_n N_A_103_367#_c_387_n
+ N_A_103_367#_c_358_n N_A_103_367#_c_359_n N_A_103_367#_c_360_n
+ N_A_103_367#_c_397_n N_A_103_367#_c_401_n N_A_103_367#_c_361_n
+ N_A_103_367#_c_362_n N_A_103_367#_c_376_n N_A_103_367#_c_398_n
+ PM_SKY130_FD_SC_LP__A41OI_2%A_103_367#
x_PM_SKY130_FD_SC_LP__A41OI_2%Y N_Y_M1011_d N_Y_M1004_s N_Y_M1001_s N_Y_c_505_p
+ N_Y_c_453_n N_Y_c_461_n N_Y_c_463_n N_Y_c_456_n N_Y_c_454_n N_Y_c_478_n Y Y
+ N_Y_c_458_n PM_SKY130_FD_SC_LP__A41OI_2%Y
x_PM_SKY130_FD_SC_LP__A41OI_2%VPWR N_VPWR_M1000_s N_VPWR_M1010_d N_VPWR_M1006_d
+ N_VPWR_M1003_d N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_520_n
+ N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n VPWR N_VPWR_c_524_n
+ N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_516_n N_VPWR_c_528_n N_VPWR_c_529_n
+ PM_SKY130_FD_SC_LP__A41OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A41OI_2%VGND N_VGND_M1011_s N_VGND_M1012_s N_VGND_M1009_d
+ N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n N_VGND_c_600_n N_VGND_c_601_n
+ N_VGND_c_602_n VGND N_VGND_c_603_n N_VGND_c_604_n N_VGND_c_605_n
+ N_VGND_c_606_n PM_SKY130_FD_SC_LP__A41OI_2%VGND
x_PM_SKY130_FD_SC_LP__A41OI_2%A_318_69# N_A_318_69#_M1004_d N_A_318_69#_M1016_d
+ N_A_318_69#_M1014_d N_A_318_69#_c_661_n N_A_318_69#_c_662_n
+ N_A_318_69#_c_663_n N_A_318_69#_c_664_n N_A_318_69#_c_665_n
+ PM_SKY130_FD_SC_LP__A41OI_2%A_318_69#
x_PM_SKY130_FD_SC_LP__A41OI_2%A_577_69# N_A_577_69#_M1002_s N_A_577_69#_M1005_s
+ N_A_577_69#_c_703_n N_A_577_69#_c_700_n N_A_577_69#_c_701_n
+ N_A_577_69#_c_702_n PM_SKY130_FD_SC_LP__A41OI_2%A_577_69#
x_PM_SKY130_FD_SC_LP__A41OI_2%A_788_69# N_A_788_69#_M1005_d N_A_788_69#_M1017_d
+ N_A_788_69#_M1019_s N_A_788_69#_c_737_n N_A_788_69#_c_731_n
+ N_A_788_69#_c_732_n N_A_788_69#_c_733_n N_A_788_69#_c_734_n
+ N_A_788_69#_c_735_n PM_SKY130_FD_SC_LP__A41OI_2%A_788_69#
cc_1 VNB N_B1_c_94_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.185
cc_2 VNB N_B1_M1001_g 0.00860042f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_3 VNB N_B1_c_96_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.185
cc_4 VNB N_B1_M1007_g 0.00603408f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_5 VNB B1 0.0279053f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_B1_c_99_n 0.067308f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.35
cc_7 VNB N_A1_M1000_g 0.00168888f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.655
cc_8 VNB N_A1_c_140_n 0.0187791f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_9 VNB N_A1_M1015_g 0.00139613f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.655
cc_10 VNB N_A1_c_142_n 0.0159543f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_11 VNB N_A1_c_143_n 0.00835596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_c_144_n 0.0604064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_M1002_g 0.0188471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_M1014_g 0.0241444f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.515
cc_15 VNB N_A2_c_201_n 0.0298279f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_A2_c_202_n 0.0392252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_M1006_g 0.00170456f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.655
cc_18 VNB N_A3_c_253_n 0.0200101f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_19 VNB N_A3_c_254_n 0.0165868f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.185
cc_20 VNB N_A3_M1008_g 0.00170419f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_21 VNB N_A3_c_256_n 0.00168242f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB A3 0.00259769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A3_c_258_n 0.0539493f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.35
cc_24 VNB N_A4_M1009_g 0.0186546f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.655
cc_25 VNB N_A4_M1019_g 0.0250995f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.515
cc_26 VNB A4 0.0193793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A4_c_318_n 0.0384835f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.35
cc_28 VNB N_Y_c_453_n 0.011216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_454_n 7.26827e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.35
cc_30 VNB Y 0.0036898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_516_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_597_n 0.012758f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.655
cc_33 VNB N_VGND_c_598_n 0.0340406f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_34 VNB N_VGND_c_599_n 0.00733726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_600_n 0.00332106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_601_n 0.0930956f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_37 VNB N_VGND_c_602_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_603_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.35
cc_39 VNB N_VGND_c_604_n 0.0203883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_605_n 0.35179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_606_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_318_69#_c_661_n 0.0049363f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.655
cc_43 VNB N_A_318_69#_c_662_n 0.00920641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_318_69#_c_663_n 0.00220982f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_45 VNB N_A_318_69#_c_664_n 0.00497646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_318_69#_c_665_n 0.00681636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_577_69#_c_700_n 0.0176559f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.515
cc_48 VNB N_A_577_69#_c_701_n 0.00203727f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_49 VNB N_A_577_69#_c_702_n 0.00202358f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_50 VNB N_A_788_69#_c_731_n 0.00189245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_788_69#_c_732_n 0.013217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_788_69#_c_733_n 0.0309544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_788_69#_c_734_n 0.0101648f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_54 VNB N_A_788_69#_c_735_n 0.00313214f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.35
cc_55 VPB N_B1_M1001_g 0.0260435f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.465
cc_56 VPB N_B1_M1007_g 0.0195822f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_57 VPB B1 0.024905f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_58 VPB N_A1_M1000_g 0.0213402f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.655
cc_59 VPB N_A1_M1015_g 0.0200914f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=0.655
cc_60 VPB N_A2_M1010_g 0.0216543f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.655
cc_61 VPB N_A2_M1018_g 0.0226972f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_62 VPB N_A2_c_201_n 0.0135674f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_63 VPB N_A2_c_202_n 0.00916969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB A2 0.00900425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A3_M1006_g 0.0207694f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.655
cc_66 VPB N_A3_M1008_g 0.0207686f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_67 VPB N_A4_M1003_g 0.0185257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A4_M1013_g 0.0242504f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_69 VPB A4 0.0152373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A4_c_318_n 0.00505959f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.35
cc_71 VPB N_A_103_367#_c_356_n 0.00788844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_103_367#_c_357_n 0.036931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_103_367#_c_358_n 0.00359109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_103_367#_c_359_n 0.00592706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_103_367#_c_360_n 0.00454365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_103_367#_c_361_n 0.00755451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_103_367#_c_362_n 0.0371313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_Y_c_456_n 0.00445338f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.35
cc_79 VPB Y 0.00155091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_Y_c_458_n 0.00499367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_517_n 0.00563065f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_82 VPB N_VPWR_c_518_n 0.00445303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_519_n 4.13242e-19 $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.35
cc_84 VPB N_VPWR_c_520_n 0.0492775f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.35
cc_85 VPB N_VPWR_c_521_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.35
cc_86 VPB N_VPWR_c_522_n 0.0159054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_523_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.48
cc_88 VPB N_VPWR_c_524_n 0.0184545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_525_n 0.0159314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_526_n 0.0193536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_516_n 0.0660573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_528_n 0.0205011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_529_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 N_B1_M1007_g N_A1_M1000_g 0.0284415f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_95 N_B1_c_99_n N_A1_c_140_n 0.00239306f $X=1.285 $Y=1.35 $X2=0 $Y2=0
cc_96 N_B1_M1001_g N_A1_c_143_n 7.80594e-19 $X=0.855 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B1_M1007_g N_A1_c_143_n 0.00483077f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_98 B1 N_A1_c_143_n 0.0212471f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B1_c_99_n N_A1_c_143_n 0.0181281f $X=1.285 $Y=1.35 $X2=0 $Y2=0
cc_100 N_B1_c_99_n N_A1_c_144_n 0.0216536f $X=1.285 $Y=1.35 $X2=0 $Y2=0
cc_101 B1 N_A_103_367#_c_357_n 0.0227746f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B1_c_99_n N_A_103_367#_c_357_n 0.00117246f $X=1.285 $Y=1.35 $X2=0 $Y2=0
cc_103 N_B1_M1001_g N_A_103_367#_c_365_n 0.0118004f $X=0.855 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_B1_M1007_g N_A_103_367#_c_365_n 0.010053f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_105 N_B1_M1007_g N_A_103_367#_c_367_n 0.00187497f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_106 N_B1_c_96_n N_Y_c_453_n 0.0188026f $X=0.98 $Y=1.185 $X2=0 $Y2=0
cc_107 N_B1_c_99_n N_Y_c_453_n 0.00792852f $X=1.285 $Y=1.35 $X2=0 $Y2=0
cc_108 B1 N_Y_c_461_n 0.0110079f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B1_c_99_n N_Y_c_461_n 0.00275918f $X=1.285 $Y=1.35 $X2=0 $Y2=0
cc_110 N_B1_M1001_g N_Y_c_463_n 0.00857378f $X=0.855 $Y=2.465 $X2=0 $Y2=0
cc_111 N_B1_M1007_g N_Y_c_463_n 0.00952563f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B1_M1001_g N_Y_c_456_n 0.00471333f $X=0.855 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B1_M1007_g N_Y_c_456_n 0.00125224f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B1_c_99_n N_Y_c_456_n 0.00396901f $X=1.285 $Y=1.35 $X2=0 $Y2=0
cc_115 N_B1_M1007_g N_Y_c_458_n 0.0111034f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B1_M1001_g N_VPWR_c_520_n 0.00357877f $X=0.855 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B1_M1007_g N_VPWR_c_520_n 0.00357842f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B1_M1001_g N_VPWR_c_516_n 0.00665089f $X=0.855 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B1_M1007_g N_VPWR_c_516_n 0.00537652f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_c_94_n N_VGND_c_598_n 0.0165374f $X=0.55 $Y=1.185 $X2=0 $Y2=0
cc_121 N_B1_c_96_n N_VGND_c_598_n 6.73275e-19 $X=0.98 $Y=1.185 $X2=0 $Y2=0
cc_122 B1 N_VGND_c_598_n 0.026791f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B1_c_94_n N_VGND_c_599_n 5.75816e-19 $X=0.55 $Y=1.185 $X2=0 $Y2=0
cc_124 N_B1_c_96_n N_VGND_c_599_n 0.0128375f $X=0.98 $Y=1.185 $X2=0 $Y2=0
cc_125 N_B1_c_94_n N_VGND_c_603_n 0.00486043f $X=0.55 $Y=1.185 $X2=0 $Y2=0
cc_126 N_B1_c_96_n N_VGND_c_603_n 0.00486043f $X=0.98 $Y=1.185 $X2=0 $Y2=0
cc_127 N_B1_c_94_n N_VGND_c_605_n 0.00824727f $X=0.55 $Y=1.185 $X2=0 $Y2=0
cc_128 N_B1_c_96_n N_VGND_c_605_n 0.00824727f $X=0.98 $Y=1.185 $X2=0 $Y2=0
cc_129 N_B1_c_96_n N_A_318_69#_c_665_n 9.59572e-19 $X=0.98 $Y=1.185 $X2=0 $Y2=0
cc_130 N_A1_M1015_g N_A2_M1010_g 0.0162174f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A1_c_142_n N_A2_M1002_g 0.0183956f $X=2.38 $Y=1.295 $X2=0 $Y2=0
cc_132 N_A1_c_144_n N_A2_c_201_n 0.0237589f $X=2.31 $Y=1.46 $X2=0 $Y2=0
cc_133 N_A1_M1000_g N_A_103_367#_c_368_n 7.32094e-19 $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A1_M1000_g N_A_103_367#_c_367_n 0.0101308f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A1_M1015_g N_A_103_367#_c_367_n 8.49982e-19 $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A1_M1000_g N_A_103_367#_c_371_n 0.0119714f $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A1_M1015_g N_A_103_367#_c_371_n 0.0119714f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A1_c_144_n N_A_103_367#_c_371_n 2.60653e-19 $X=2.31 $Y=1.46 $X2=0 $Y2=0
cc_139 N_A1_M1000_g N_A_103_367#_c_374_n 7.30796e-19 $X=1.715 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A1_M1015_g N_A_103_367#_c_374_n 0.00955916f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A1_M1015_g N_A_103_367#_c_376_n 0.00151803f $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A1_c_140_n N_Y_c_453_n 0.0144824f $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_143 N_A1_c_143_n N_Y_c_453_n 0.059245f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_144 N_A1_c_144_n N_Y_c_453_n 0.00159907f $X=2.31 $Y=1.46 $X2=0 $Y2=0
cc_145 N_A1_M1000_g N_Y_c_463_n 7.61432e-19 $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A1_c_143_n N_Y_c_456_n 0.0105448f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_147 N_A1_c_140_n N_Y_c_454_n 0.00127782f $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_148 N_A1_c_142_n N_Y_c_454_n 0.00384706f $X=2.38 $Y=1.295 $X2=0 $Y2=0
cc_149 N_A1_c_143_n N_Y_c_454_n 0.0170828f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_150 N_A1_c_144_n N_Y_c_454_n 0.0101181f $X=2.31 $Y=1.46 $X2=0 $Y2=0
cc_151 N_A1_c_140_n N_Y_c_478_n 0.0108323f $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_152 N_A1_c_142_n N_Y_c_478_n 0.00482495f $X=2.38 $Y=1.295 $X2=0 $Y2=0
cc_153 N_A1_M1000_g Y 0.00396119f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A1_M1015_g Y 0.0150323f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A1_c_143_n Y 0.0154911f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_156 N_A1_c_144_n Y 0.0220568f $X=2.31 $Y=1.46 $X2=0 $Y2=0
cc_157 N_A1_M1000_g N_Y_c_458_n 0.0112664f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A1_c_143_n N_Y_c_458_n 0.0505521f $X=1.735 $Y=1.46 $X2=0 $Y2=0
cc_159 N_A1_c_144_n N_Y_c_458_n 0.00928761f $X=2.31 $Y=1.46 $X2=0 $Y2=0
cc_160 N_A1_M1000_g N_VPWR_c_517_n 0.00709273f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A1_M1015_g N_VPWR_c_517_n 0.00947696f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A1_M1000_g N_VPWR_c_520_n 0.00547432f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A1_M1015_g N_VPWR_c_524_n 0.0054895f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A1_M1000_g N_VPWR_c_516_n 0.0102865f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A1_M1015_g N_VPWR_c_516_n 0.0103372f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A1_c_140_n N_VGND_c_599_n 7.33568e-19 $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_167 N_A1_c_140_n N_VGND_c_601_n 0.0029147f $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_168 N_A1_c_142_n N_VGND_c_601_n 0.0029147f $X=2.38 $Y=1.295 $X2=0 $Y2=0
cc_169 N_A1_c_140_n N_VGND_c_605_n 0.00428625f $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_170 N_A1_c_142_n N_VGND_c_605_n 0.00399217f $X=2.38 $Y=1.295 $X2=0 $Y2=0
cc_171 N_A1_c_140_n N_A_318_69#_c_661_n 0.00970681f $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_172 N_A1_c_142_n N_A_318_69#_c_661_n 0.0118596f $X=2.38 $Y=1.295 $X2=0 $Y2=0
cc_173 N_A1_c_142_n N_A_318_69#_c_663_n 5.73473e-19 $X=2.38 $Y=1.295 $X2=0 $Y2=0
cc_174 N_A1_c_140_n N_A_318_69#_c_665_n 8.76155e-19 $X=1.95 $Y=1.295 $X2=0 $Y2=0
cc_175 N_A2_M1018_g N_A3_M1006_g 0.0182808f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A2_c_202_n N_A3_c_256_n 9.33813e-19 $X=3.675 $Y=1.51 $X2=0 $Y2=0
cc_177 A2 N_A3_c_256_n 0.00480345f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A2_c_202_n N_A3_c_258_n 0.0182808f $X=3.675 $Y=1.51 $X2=0 $Y2=0
cc_179 A2 N_A3_c_258_n 9.93491e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A2_M1010_g N_A_103_367#_c_374_n 0.0140269f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A2_M1010_g N_A_103_367#_c_378_n 0.0150475f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A2_M1018_g N_A_103_367#_c_378_n 0.0210774f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A2_c_201_n N_A_103_367#_c_378_n 0.00496877f $X=3.315 $Y=1.51 $X2=0
+ $Y2=0
cc_184 A2 N_A_103_367#_c_378_n 0.0377216f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A2_M1018_g N_A_103_367#_c_359_n 0.0011358f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_186 A2 N_A_103_367#_c_359_n 0.010199f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A2_M1010_g N_A_103_367#_c_376_n 8.11192e-19 $X=2.74 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A2_M1002_g N_Y_c_454_n 5.16772e-19 $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_189 N_A2_c_201_n N_Y_c_454_n 4.67438e-19 $X=3.315 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A2_M1010_g Y 0.0145707f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A2_c_201_n Y 0.0111316f $X=3.315 $Y=1.51 $X2=0 $Y2=0
cc_192 A2 Y 0.0349007f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_M1010_g N_VPWR_c_524_n 0.0054895f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A2_M1018_g N_VPWR_c_525_n 0.00487821f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A2_M1010_g N_VPWR_c_516_n 0.0112981f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A2_M1018_g N_VPWR_c_516_n 0.00827265f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A2_M1010_g N_VPWR_c_528_n 0.0163163f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A2_M1018_g N_VPWR_c_528_n 0.0118433f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A2_M1002_g N_VGND_c_601_n 0.00450424f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_200 N_A2_M1014_g N_VGND_c_601_n 0.00291444f $X=3.24 $Y=0.765 $X2=0 $Y2=0
cc_201 N_A2_M1002_g N_VGND_c_605_n 0.00862457f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_202 N_A2_M1014_g N_VGND_c_605_n 0.00428623f $X=3.24 $Y=0.765 $X2=0 $Y2=0
cc_203 N_A2_M1002_g N_A_318_69#_c_661_n 7.3655e-19 $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_204 N_A2_M1002_g N_A_318_69#_c_662_n 0.0155059f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_205 N_A2_M1014_g N_A_318_69#_c_662_n 0.0138552f $X=3.24 $Y=0.765 $X2=0 $Y2=0
cc_206 N_A2_c_201_n N_A_318_69#_c_662_n 0.00376468f $X=3.315 $Y=1.51 $X2=0 $Y2=0
cc_207 N_A2_c_202_n N_A_318_69#_c_662_n 0.010072f $X=3.675 $Y=1.51 $X2=0 $Y2=0
cc_208 A2 N_A_318_69#_c_662_n 0.0568281f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A2_c_201_n N_A_318_69#_c_663_n 7.49468e-19 $X=3.315 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A2_M1002_g N_A_577_69#_c_703_n 0.00527422f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_211 N_A2_M1014_g N_A_577_69#_c_703_n 0.0110663f $X=3.24 $Y=0.765 $X2=0 $Y2=0
cc_212 N_A2_M1014_g N_A_577_69#_c_700_n 0.0102755f $X=3.24 $Y=0.765 $X2=0 $Y2=0
cc_213 N_A2_M1002_g N_A_577_69#_c_701_n 0.00291412f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_214 N_A2_M1014_g N_A_577_69#_c_701_n 0.00159238f $X=3.24 $Y=0.765 $X2=0 $Y2=0
cc_215 N_A2_M1014_g N_A_788_69#_c_734_n 0.00114518f $X=3.24 $Y=0.765 $X2=0 $Y2=0
cc_216 N_A3_c_254_n N_A4_M1009_g 0.0183223f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_217 A3 N_A4_M1009_g 6.40299e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A3_M1008_g N_A4_M1003_g 0.0183223f $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_219 A3 A4 0.00442422f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A3_c_258_n A4 0.00136683f $X=4.78 $Y=1.46 $X2=0 $Y2=0
cc_221 A3 N_A4_c_318_n 8.00014e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_222 N_A3_c_258_n N_A4_c_318_n 0.0183223f $X=4.78 $Y=1.46 $X2=0 $Y2=0
cc_223 N_A3_M1006_g N_A_103_367#_c_385_n 0.00413617f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_224 N_A3_M1008_g N_A_103_367#_c_385_n 7.7589e-19 $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A3_M1006_g N_A_103_367#_c_387_n 0.00892035f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_226 N_A3_M1006_g N_A_103_367#_c_358_n 0.0119774f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A3_M1008_g N_A_103_367#_c_358_n 0.0126609f $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A3_c_256_n N_A_103_367#_c_358_n 0.0187768f $X=4.4 $Y=1.46 $X2=0 $Y2=0
cc_229 A3 N_A_103_367#_c_358_n 0.0286078f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_230 N_A3_c_258_n N_A_103_367#_c_358_n 0.00738242f $X=4.78 $Y=1.46 $X2=0 $Y2=0
cc_231 N_A3_M1006_g N_A_103_367#_c_359_n 0.00189415f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_A3_c_256_n N_A_103_367#_c_359_n 0.00190438f $X=4.4 $Y=1.46 $X2=0 $Y2=0
cc_233 N_A3_M1006_g N_A_103_367#_c_360_n 7.67971e-19 $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A3_M1008_g N_A_103_367#_c_360_n 0.00642042f $X=4.78 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A3_M1008_g N_A_103_367#_c_397_n 0.0120846f $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A3_M1006_g N_A_103_367#_c_398_n 0.0030869f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A3_M1006_g N_VPWR_c_518_n 0.0118485f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A3_M1008_g N_VPWR_c_518_n 0.0118513f $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A3_M1008_g N_VPWR_c_519_n 7.47121e-19 $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A3_M1008_g N_VPWR_c_522_n 0.0054895f $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A3_M1006_g N_VPWR_c_525_n 0.0054895f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_242 N_A3_M1006_g N_VPWR_c_516_n 0.0103474f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A3_M1008_g N_VPWR_c_516_n 0.0103474f $X=4.78 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A3_M1006_g N_VPWR_c_528_n 6.97376e-19 $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A3_c_254_n N_VGND_c_600_n 6.40654e-19 $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_246 N_A3_c_253_n N_VGND_c_601_n 0.00292717f $X=4.35 $Y=1.295 $X2=0 $Y2=0
cc_247 N_A3_c_254_n N_VGND_c_601_n 0.00451696f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_248 N_A3_c_253_n N_VGND_c_605_n 0.00427714f $X=4.35 $Y=1.295 $X2=0 $Y2=0
cc_249 N_A3_c_254_n N_VGND_c_605_n 0.00866163f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_250 N_A3_c_253_n N_A_318_69#_c_662_n 0.00154513f $X=4.35 $Y=1.295 $X2=0 $Y2=0
cc_251 N_A3_c_253_n N_A_577_69#_c_700_n 0.0106221f $X=4.35 $Y=1.295 $X2=0 $Y2=0
cc_252 N_A3_c_253_n N_A_577_69#_c_702_n 0.0113942f $X=4.35 $Y=1.295 $X2=0 $Y2=0
cc_253 N_A3_c_254_n N_A_577_69#_c_702_n 0.00696754f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_254 N_A3_c_253_n N_A_788_69#_c_737_n 0.0128846f $X=4.35 $Y=1.295 $X2=0 $Y2=0
cc_255 N_A3_c_254_n N_A_788_69#_c_737_n 0.0134234f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_256 N_A3_c_256_n N_A_788_69#_c_737_n 0.00578606f $X=4.4 $Y=1.46 $X2=0 $Y2=0
cc_257 A3 N_A_788_69#_c_737_n 0.0235645f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_258 N_A3_c_258_n N_A_788_69#_c_737_n 5.6365e-19 $X=4.78 $Y=1.46 $X2=0 $Y2=0
cc_259 N_A3_c_254_n N_A_788_69#_c_731_n 8.28776e-19 $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_260 N_A3_c_253_n N_A_788_69#_c_734_n 0.00365483f $X=4.35 $Y=1.295 $X2=0 $Y2=0
cc_261 N_A3_c_256_n N_A_788_69#_c_734_n 0.00990997f $X=4.4 $Y=1.46 $X2=0 $Y2=0
cc_262 N_A3_c_258_n N_A_788_69#_c_734_n 0.00370085f $X=4.78 $Y=1.46 $X2=0 $Y2=0
cc_263 N_A3_c_254_n N_A_788_69#_c_735_n 0.00113557f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_264 A3 N_A_788_69#_c_735_n 0.00365123f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_265 N_A4_M1003_g N_A_103_367#_c_360_n 0.00296783f $X=5.21 $Y=2.465 $X2=0
+ $Y2=0
cc_266 A4 N_A_103_367#_c_360_n 0.00303083f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_267 N_A4_M1003_g N_A_103_367#_c_401_n 0.0139984f $X=5.21 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A4_M1013_g N_A_103_367#_c_401_n 0.01229f $X=5.64 $Y=2.465 $X2=0 $Y2=0
cc_269 A4 N_A_103_367#_c_401_n 0.0319853f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_270 N_A4_c_318_n N_A_103_367#_c_401_n 5.76518e-19 $X=5.64 $Y=1.51 $X2=0 $Y2=0
cc_271 A4 N_A_103_367#_c_361_n 0.0215874f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_272 N_A4_M1003_g N_VPWR_c_519_n 0.0147983f $X=5.21 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A4_M1013_g N_VPWR_c_519_n 0.0164949f $X=5.64 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A4_M1003_g N_VPWR_c_522_n 0.00486043f $X=5.21 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A4_M1013_g N_VPWR_c_526_n 0.00486043f $X=5.64 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A4_M1003_g N_VPWR_c_516_n 0.0082726f $X=5.21 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A4_M1013_g N_VPWR_c_516_n 0.00927852f $X=5.64 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A4_M1009_g N_VGND_c_600_n 0.0103699f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_279 N_A4_M1019_g N_VGND_c_600_n 0.0127653f $X=5.64 $Y=0.765 $X2=0 $Y2=0
cc_280 N_A4_M1009_g N_VGND_c_601_n 0.00400407f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_281 N_A4_M1019_g N_VGND_c_604_n 0.00400407f $X=5.64 $Y=0.765 $X2=0 $Y2=0
cc_282 N_A4_M1009_g N_VGND_c_605_n 0.00775088f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_283 N_A4_M1019_g N_VGND_c_605_n 0.00798302f $X=5.64 $Y=0.765 $X2=0 $Y2=0
cc_284 N_A4_M1009_g N_A_577_69#_c_702_n 3.12158e-19 $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_285 N_A4_M1009_g N_A_788_69#_c_731_n 8.28776e-19 $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_286 N_A4_M1009_g N_A_788_69#_c_732_n 0.0146436f $X=5.21 $Y=0.765 $X2=0 $Y2=0
cc_287 N_A4_M1019_g N_A_788_69#_c_732_n 0.0136069f $X=5.64 $Y=0.765 $X2=0 $Y2=0
cc_288 A4 N_A_788_69#_c_732_n 0.0607174f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_289 N_A4_c_318_n N_A_788_69#_c_732_n 0.00246472f $X=5.64 $Y=1.51 $X2=0 $Y2=0
cc_290 N_A4_M1019_g N_A_788_69#_c_733_n 0.00354556f $X=5.64 $Y=0.765 $X2=0 $Y2=0
cc_291 N_A_103_367#_c_365_n N_Y_M1001_s 0.00332931f $X=1.335 $Y=2.985 $X2=0
+ $Y2=0
cc_292 N_A_103_367#_c_365_n N_Y_c_463_n 0.0160814f $X=1.335 $Y=2.985 $X2=0 $Y2=0
cc_293 N_A_103_367#_M1015_d Y 0.00182683f $X=2.385 $Y=1.835 $X2=0 $Y2=0
cc_294 N_A_103_367#_c_378_n Y 0.00823312f $X=3.855 $Y=2.222 $X2=0 $Y2=0
cc_295 N_A_103_367#_c_376_n Y 0.018662f $X=2.525 $Y=2.205 $X2=0 $Y2=0
cc_296 N_A_103_367#_M1007_d N_Y_c_458_n 0.00176461f $X=1.36 $Y=1.835 $X2=0 $Y2=0
cc_297 N_A_103_367#_c_368_n N_Y_c_458_n 0.0153678f $X=1.535 $Y=2.29 $X2=0 $Y2=0
cc_298 N_A_103_367#_c_371_n N_Y_c_458_n 0.0424013f $X=2.36 $Y=2.205 $X2=0 $Y2=0
cc_299 N_A_103_367#_c_371_n N_VPWR_M1000_s 0.00747546f $X=2.36 $Y=2.205
+ $X2=-0.19 $Y2=1.655
cc_300 N_A_103_367#_c_378_n N_VPWR_M1010_d 0.0236999f $X=3.855 $Y=2.222 $X2=0
+ $Y2=0
cc_301 N_A_103_367#_c_358_n N_VPWR_M1006_d 0.0037308f $X=4.83 $Y=1.8 $X2=0 $Y2=0
cc_302 N_A_103_367#_c_401_n N_VPWR_M1003_d 0.0033481f $X=5.76 $Y=2.01 $X2=0
+ $Y2=0
cc_303 N_A_103_367#_c_371_n N_VPWR_c_517_n 0.0266042f $X=2.36 $Y=2.205 $X2=0
+ $Y2=0
cc_304 N_A_103_367#_c_374_n N_VPWR_c_517_n 0.0447249f $X=2.525 $Y=2.94 $X2=0
+ $Y2=0
cc_305 N_A_103_367#_c_385_n N_VPWR_c_518_n 0.00463015f $X=3.965 $Y=1.98 $X2=0
+ $Y2=0
cc_306 N_A_103_367#_c_387_n N_VPWR_c_518_n 0.0535654f $X=3.965 $Y=2.445 $X2=0
+ $Y2=0
cc_307 N_A_103_367#_c_358_n N_VPWR_c_518_n 0.0266856f $X=4.83 $Y=1.8 $X2=0 $Y2=0
cc_308 N_A_103_367#_c_360_n N_VPWR_c_518_n 0.00308638f $X=4.96 $Y=2.095 $X2=0
+ $Y2=0
cc_309 N_A_103_367#_c_397_n N_VPWR_c_518_n 0.0700025f $X=4.995 $Y=2.445 $X2=0
+ $Y2=0
cc_310 N_A_103_367#_c_398_n N_VPWR_c_518_n 0.0158177f $X=3.992 $Y=2.222 $X2=0
+ $Y2=0
cc_311 N_A_103_367#_c_401_n N_VPWR_c_519_n 0.0170777f $X=5.76 $Y=2.01 $X2=0
+ $Y2=0
cc_312 N_A_103_367#_c_356_n N_VPWR_c_520_n 0.0179183f $X=0.605 $Y=2.895 $X2=0
+ $Y2=0
cc_313 N_A_103_367#_c_365_n N_VPWR_c_520_n 0.0330957f $X=1.335 $Y=2.985 $X2=0
+ $Y2=0
cc_314 N_A_103_367#_c_367_n N_VPWR_c_520_n 0.0189216f $X=1.535 $Y=2.885 $X2=0
+ $Y2=0
cc_315 N_A_103_367#_c_397_n N_VPWR_c_522_n 0.015688f $X=4.995 $Y=2.445 $X2=0
+ $Y2=0
cc_316 N_A_103_367#_c_374_n N_VPWR_c_524_n 0.0189236f $X=2.525 $Y=2.94 $X2=0
+ $Y2=0
cc_317 N_A_103_367#_c_387_n N_VPWR_c_525_n 0.015688f $X=3.965 $Y=2.445 $X2=0
+ $Y2=0
cc_318 N_A_103_367#_c_362_n N_VPWR_c_526_n 0.0178111f $X=5.855 $Y=2.91 $X2=0
+ $Y2=0
cc_319 N_A_103_367#_M1001_d N_VPWR_c_516_n 0.00215161f $X=0.515 $Y=1.835 $X2=0
+ $Y2=0
cc_320 N_A_103_367#_M1007_d N_VPWR_c_516_n 0.00223559f $X=1.36 $Y=1.835 $X2=0
+ $Y2=0
cc_321 N_A_103_367#_M1015_d N_VPWR_c_516_n 0.00223559f $X=2.385 $Y=1.835 $X2=0
+ $Y2=0
cc_322 N_A_103_367#_M1018_s N_VPWR_c_516_n 0.00380103f $X=3.825 $Y=1.835 $X2=0
+ $Y2=0
cc_323 N_A_103_367#_M1008_s N_VPWR_c_516_n 0.00380103f $X=4.855 $Y=1.835 $X2=0
+ $Y2=0
cc_324 N_A_103_367#_M1013_s N_VPWR_c_516_n 0.00371702f $X=5.715 $Y=1.835 $X2=0
+ $Y2=0
cc_325 N_A_103_367#_c_356_n N_VPWR_c_516_n 0.0101082f $X=0.605 $Y=2.895 $X2=0
+ $Y2=0
cc_326 N_A_103_367#_c_365_n N_VPWR_c_516_n 0.0212559f $X=1.335 $Y=2.985 $X2=0
+ $Y2=0
cc_327 N_A_103_367#_c_367_n N_VPWR_c_516_n 0.0123762f $X=1.535 $Y=2.885 $X2=0
+ $Y2=0
cc_328 N_A_103_367#_c_374_n N_VPWR_c_516_n 0.0123859f $X=2.525 $Y=2.94 $X2=0
+ $Y2=0
cc_329 N_A_103_367#_c_387_n N_VPWR_c_516_n 0.00984745f $X=3.965 $Y=2.445 $X2=0
+ $Y2=0
cc_330 N_A_103_367#_c_397_n N_VPWR_c_516_n 0.0098316f $X=4.995 $Y=2.445 $X2=0
+ $Y2=0
cc_331 N_A_103_367#_c_362_n N_VPWR_c_516_n 0.0100304f $X=5.855 $Y=2.91 $X2=0
+ $Y2=0
cc_332 N_A_103_367#_c_378_n N_VPWR_c_528_n 0.0606239f $X=3.855 $Y=2.222 $X2=0
+ $Y2=0
cc_333 N_A_103_367#_c_358_n N_A_788_69#_c_737_n 9.51656e-19 $X=4.83 $Y=1.8 $X2=0
+ $Y2=0
cc_334 N_A_103_367#_c_360_n N_A_788_69#_c_737_n 0.00138667f $X=4.96 $Y=2.095
+ $X2=0 $Y2=0
cc_335 N_A_103_367#_c_401_n N_A_788_69#_c_732_n 0.00310167f $X=5.76 $Y=2.01
+ $X2=0 $Y2=0
cc_336 N_A_103_367#_c_359_n N_A_788_69#_c_734_n 0.00881426f $X=4.13 $Y=1.8 $X2=0
+ $Y2=0
cc_337 N_A_103_367#_c_360_n N_A_788_69#_c_735_n 0.00796346f $X=4.96 $Y=2.095
+ $X2=0 $Y2=0
cc_338 Y N_VPWR_M1000_s 0.00114732f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_339 N_Y_c_458_n N_VPWR_M1000_s 0.002902f $X=2.07 $Y=1.687 $X2=-0.19
+ $Y2=-0.245
cc_340 N_Y_M1001_s N_VPWR_c_516_n 0.00225186f $X=0.93 $Y=1.835 $X2=0 $Y2=0
cc_341 N_Y_c_453_n N_VGND_M1012_s 0.00466584f $X=2 $Y=0.955 $X2=0 $Y2=0
cc_342 N_Y_c_453_n N_VGND_c_599_n 0.0220026f $X=2 $Y=0.955 $X2=0 $Y2=0
cc_343 N_Y_c_505_p N_VGND_c_603_n 0.0124525f $X=0.765 $Y=0.42 $X2=0 $Y2=0
cc_344 N_Y_M1011_d N_VGND_c_605_n 0.00536646f $X=0.625 $Y=0.235 $X2=0 $Y2=0
cc_345 N_Y_c_505_p N_VGND_c_605_n 0.00730901f $X=0.765 $Y=0.42 $X2=0 $Y2=0
cc_346 N_Y_c_453_n N_A_318_69#_M1004_d 0.00536966f $X=2 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_347 N_Y_M1004_s N_A_318_69#_c_661_n 0.00176461f $X=2.025 $Y=0.345 $X2=0 $Y2=0
cc_348 N_Y_c_453_n N_A_318_69#_c_661_n 0.00387154f $X=2 $Y=0.955 $X2=0 $Y2=0
cc_349 N_Y_c_478_n N_A_318_69#_c_661_n 0.015927f $X=2.165 $Y=0.68 $X2=0 $Y2=0
cc_350 Y N_A_318_69#_c_662_n 0.00828959f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_351 N_Y_c_454_n N_A_318_69#_c_663_n 0.00939595f $X=2.165 $Y=1.06 $X2=0 $Y2=0
cc_352 Y N_A_318_69#_c_663_n 0.0172749f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_353 N_Y_c_453_n N_A_318_69#_c_665_n 0.0211076f $X=2 $Y=0.955 $X2=0 $Y2=0
cc_354 N_VGND_c_601_n N_A_318_69#_c_661_n 0.0558783f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_605_n N_A_318_69#_c_661_n 0.0312081f $X=6 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_599_n N_A_318_69#_c_665_n 0.0338453f $X=1.195 $Y=0.575 $X2=0
+ $Y2=0
cc_357 N_VGND_c_601_n N_A_318_69#_c_665_n 0.0193073f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_605_n N_A_318_69#_c_665_n 0.0106918f $X=6 $Y=0 $X2=0 $Y2=0
cc_359 N_VGND_c_601_n N_A_577_69#_c_700_n 0.0771922f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_605_n N_A_577_69#_c_700_n 0.0443523f $X=6 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_601_n N_A_577_69#_c_701_n 0.0234284f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_605_n N_A_577_69#_c_701_n 0.0125908f $X=6 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_600_n N_A_577_69#_c_702_n 0.00206987f $X=5.425 $Y=0.47 $X2=0
+ $Y2=0
cc_364 N_VGND_c_601_n N_A_577_69#_c_702_n 0.0226204f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_605_n N_A_577_69#_c_702_n 0.0123953f $X=6 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_600_n N_A_788_69#_c_731_n 0.0211767f $X=5.425 $Y=0.47 $X2=0
+ $Y2=0
cc_367 N_VGND_c_601_n N_A_788_69#_c_731_n 0.00932315f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_605_n N_A_788_69#_c_731_n 0.00704664f $X=6 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_M1009_d N_A_788_69#_c_732_n 0.00176461f $X=5.285 $Y=0.345 $X2=0
+ $Y2=0
cc_370 N_VGND_c_600_n N_A_788_69#_c_732_n 0.0170777f $X=5.425 $Y=0.47 $X2=0
+ $Y2=0
cc_371 N_VGND_c_600_n N_A_788_69#_c_733_n 0.0229007f $X=5.425 $Y=0.47 $X2=0
+ $Y2=0
cc_372 N_VGND_c_604_n N_A_788_69#_c_733_n 0.0127923f $X=6 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_c_605_n N_A_788_69#_c_733_n 0.00966963f $X=6 $Y=0 $X2=0 $Y2=0
cc_374 N_A_318_69#_c_662_n N_A_577_69#_M1002_s 0.00176461f $X=3.36 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_375 N_A_318_69#_c_662_n N_A_577_69#_c_703_n 0.017036f $X=3.36 $Y=1.17 $X2=0
+ $Y2=0
cc_376 N_A_318_69#_M1014_d N_A_577_69#_c_700_n 0.00363296f $X=3.315 $Y=0.345
+ $X2=0 $Y2=0
cc_377 N_A_318_69#_c_662_n N_A_577_69#_c_700_n 0.00272017f $X=3.36 $Y=1.17 $X2=0
+ $Y2=0
cc_378 N_A_318_69#_c_664_n N_A_577_69#_c_700_n 0.0241848f $X=3.525 $Y=0.68 $X2=0
+ $Y2=0
cc_379 N_A_318_69#_c_661_n N_A_577_69#_c_701_n 0.011362f $X=2.5 $Y=0.34 $X2=0
+ $Y2=0
cc_380 N_A_318_69#_c_662_n N_A_788_69#_c_734_n 0.00914659f $X=3.36 $Y=1.17 $X2=0
+ $Y2=0
cc_381 N_A_318_69#_c_664_n N_A_788_69#_c_734_n 0.0351506f $X=3.525 $Y=0.68 $X2=0
+ $Y2=0
cc_382 N_A_577_69#_c_700_n N_A_788_69#_M1005_d 0.00363296f $X=4.4 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_383 N_A_577_69#_M1005_s N_A_788_69#_c_737_n 0.00332815f $X=4.425 $Y=0.345
+ $X2=0 $Y2=0
cc_384 N_A_577_69#_c_700_n N_A_788_69#_c_737_n 0.00388708f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_385 N_A_577_69#_c_702_n N_A_788_69#_c_737_n 0.0165025f $X=4.565 $Y=0.34 $X2=0
+ $Y2=0
cc_386 N_A_577_69#_c_702_n N_A_788_69#_c_731_n 0.0147979f $X=4.565 $Y=0.34 $X2=0
+ $Y2=0
cc_387 N_A_577_69#_c_700_n N_A_788_69#_c_734_n 0.0240386f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
