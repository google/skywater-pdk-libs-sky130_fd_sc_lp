* File: sky130_fd_sc_lp__xnor3_1.pxi.spice
* Created: Wed Sep  2 10:40:41 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR3_1%A_81_259# N_A_81_259#_M1010_d N_A_81_259#_M1011_d
+ N_A_81_259#_M1020_g N_A_81_259#_M1019_g N_A_81_259#_c_160_n
+ N_A_81_259#_c_161_n N_A_81_259#_c_237_p N_A_81_259#_c_168_n
+ N_A_81_259#_c_169_n N_A_81_259#_c_170_n N_A_81_259#_c_162_n
+ N_A_81_259#_c_163_n N_A_81_259#_c_164_n N_A_81_259#_c_179_p
+ N_A_81_259#_c_165_n PM_SKY130_FD_SC_LP__XNOR3_1%A_81_259#
x_PM_SKY130_FD_SC_LP__XNOR3_1%C N_C_M1006_g N_C_M1014_g N_C_c_249_n N_C_M1010_g
+ N_C_M1011_g N_C_c_252_n C N_C_c_253_n N_C_c_254_n
+ PM_SKY130_FD_SC_LP__XNOR3_1%C
x_PM_SKY130_FD_SC_LP__XNOR3_1%A_244_137# N_A_244_137#_M1006_d
+ N_A_244_137#_M1014_d N_A_244_137#_M1009_g N_A_244_137#_M1016_g
+ N_A_244_137#_c_319_n N_A_244_137#_c_320_n N_A_244_137#_c_321_n
+ N_A_244_137#_c_322_n N_A_244_137#_c_323_n
+ PM_SKY130_FD_SC_LP__XNOR3_1%A_244_137#
x_PM_SKY130_FD_SC_LP__XNOR3_1%A_754_367# N_A_754_367#_M1002_d
+ N_A_754_367#_M1021_d N_A_754_367#_M1012_g N_A_754_367#_M1000_g
+ N_A_754_367#_c_385_n N_A_754_367#_c_386_n N_A_754_367#_M1008_g
+ N_A_754_367#_M1001_g N_A_754_367#_c_389_n N_A_754_367#_c_390_n
+ N_A_754_367#_c_397_n N_A_754_367#_c_398_n N_A_754_367#_c_399_n
+ N_A_754_367#_c_391_n N_A_754_367#_c_392_n N_A_754_367#_c_393_n
+ PM_SKY130_FD_SC_LP__XNOR3_1%A_754_367#
x_PM_SKY130_FD_SC_LP__XNOR3_1%B N_B_M1021_g N_B_M1002_g N_B_c_500_n N_B_c_509_n
+ N_B_c_510_n N_B_c_511_n N_B_M1017_g N_B_M1004_g N_B_c_513_n N_B_M1013_g
+ N_B_M1007_g N_B_c_503_n N_B_c_516_n N_B_c_504_n B N_B_c_505_n N_B_c_506_n
+ PM_SKY130_FD_SC_LP__XNOR3_1%B
x_PM_SKY130_FD_SC_LP__XNOR3_1%A N_A_M1003_g N_A_M1018_g A N_A_c_632_n
+ PM_SKY130_FD_SC_LP__XNOR3_1%A
x_PM_SKY130_FD_SC_LP__XNOR3_1%A_871_373# N_A_871_373#_M1000_s
+ N_A_871_373#_M1007_d N_A_871_373#_M1012_s N_A_871_373#_M1013_d
+ N_A_871_373#_M1015_g N_A_871_373#_M1005_g N_A_871_373#_c_688_n
+ N_A_871_373#_c_681_n N_A_871_373#_c_720_n N_A_871_373#_c_689_n
+ N_A_871_373#_c_690_n N_A_871_373#_c_724_n N_A_871_373#_c_727_n
+ N_A_871_373#_c_691_n N_A_871_373#_c_682_n N_A_871_373#_c_693_n
+ N_A_871_373#_c_683_n N_A_871_373#_c_684_n N_A_871_373#_c_685_n
+ N_A_871_373#_c_686_n PM_SKY130_FD_SC_LP__XNOR3_1%A_871_373#
x_PM_SKY130_FD_SC_LP__XNOR3_1%X N_X_M1019_s N_X_M1020_s N_X_c_804_n N_X_c_805_n
+ N_X_c_801_n X X N_X_c_803_n X PM_SKY130_FD_SC_LP__XNOR3_1%X
x_PM_SKY130_FD_SC_LP__XNOR3_1%VPWR N_VPWR_M1020_d N_VPWR_M1021_s N_VPWR_M1018_d
+ N_VPWR_c_824_n N_VPWR_c_825_n N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n
+ VPWR N_VPWR_c_829_n N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_823_n
+ N_VPWR_c_833_n N_VPWR_c_834_n PM_SKY130_FD_SC_LP__XNOR3_1%VPWR
x_PM_SKY130_FD_SC_LP__XNOR3_1%A_355_451# N_A_355_451#_M1009_d
+ N_A_355_451#_M1001_d N_A_355_451#_M1011_s N_A_355_451#_M1012_d
+ N_A_355_451#_c_906_n N_A_355_451#_c_907_n N_A_355_451#_c_915_n
+ N_A_355_451#_c_901_n N_A_355_451#_c_902_n N_A_355_451#_c_909_n
+ N_A_355_451#_c_910_n N_A_355_451#_c_943_n N_A_355_451#_c_903_n
+ N_A_355_451#_c_911_n N_A_355_451#_c_904_n N_A_355_451#_c_905_n
+ N_A_355_451#_c_953_n PM_SKY130_FD_SC_LP__XNOR3_1%A_355_451#
x_PM_SKY130_FD_SC_LP__XNOR3_1%A_354_109# N_A_354_109#_M1010_s
+ N_A_354_109#_M1000_d N_A_354_109#_M1016_d N_A_354_109#_M1008_d
+ N_A_354_109#_c_1049_n N_A_354_109#_c_1037_n N_A_354_109#_c_1038_n
+ N_A_354_109#_c_1039_n N_A_354_109#_c_1040_n N_A_354_109#_c_1041_n
+ N_A_354_109#_c_1042_n N_A_354_109#_c_1081_n N_A_354_109#_c_1043_n
+ N_A_354_109#_c_1044_n N_A_354_109#_c_1088_n N_A_354_109#_c_1045_n
+ PM_SKY130_FD_SC_LP__XNOR3_1%A_354_109#
x_PM_SKY130_FD_SC_LP__XNOR3_1%A_1090_373# N_A_1090_373#_M1004_d
+ N_A_1090_373#_M1015_d N_A_1090_373#_M1017_d N_A_1090_373#_M1005_d
+ N_A_1090_373#_c_1148_n N_A_1090_373#_c_1149_n N_A_1090_373#_c_1141_n
+ N_A_1090_373#_c_1142_n N_A_1090_373#_c_1150_n N_A_1090_373#_c_1143_n
+ N_A_1090_373#_c_1144_n N_A_1090_373#_c_1145_n N_A_1090_373#_c_1146_n
+ N_A_1090_373#_c_1151_n N_A_1090_373#_c_1147_n N_A_1090_373#_c_1164_n
+ N_A_1090_373#_c_1178_n N_A_1090_373#_c_1218_n N_A_1090_373#_c_1153_n
+ N_A_1090_373#_c_1154_n PM_SKY130_FD_SC_LP__XNOR3_1%A_1090_373#
x_PM_SKY130_FD_SC_LP__XNOR3_1%VGND N_VGND_M1019_d N_VGND_M1002_s N_VGND_M1003_d
+ N_VGND_c_1249_n N_VGND_c_1250_n N_VGND_c_1251_n N_VGND_c_1252_n VGND
+ N_VGND_c_1253_n N_VGND_c_1254_n N_VGND_c_1255_n N_VGND_c_1256_n
+ N_VGND_c_1257_n PM_SKY130_FD_SC_LP__XNOR3_1%VGND
cc_1 VNB N_A_81_259#_M1020_g 0.00181071f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_2 VNB N_A_81_259#_M1019_g 0.0278454f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.685
cc_3 VNB N_A_81_259#_c_160_n 4.15939e-19 $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.95
cc_4 VNB N_A_81_259#_c_161_n 0.0177864f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=0.62
cc_5 VNB N_A_81_259#_c_162_n 0.00517772f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_6 VNB N_A_81_259#_c_163_n 0.034243f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_7 VNB N_A_81_259#_c_164_n 0.00336775f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.295
cc_8 VNB N_A_81_259#_c_165_n 0.00355747f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.62
cc_9 VNB N_C_M1006_g 0.0281378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_C_c_249_n 0.0449953f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_11 VNB N_C_M1010_g 0.0246813f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.685
cc_12 VNB N_C_M1011_g 0.00892937f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.625
cc_13 VNB N_C_c_252_n 0.00550773f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=0.62
cc_14 VNB N_C_c_253_n 0.0241114f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.865
cc_15 VNB N_C_c_254_n 7.37582e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_244_137#_M1009_g 0.0364918f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_17 VNB N_A_244_137#_c_319_n 0.0073928f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.705
cc_18 VNB N_A_244_137#_c_320_n 0.00502554f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.62
cc_19 VNB N_A_244_137#_c_321_n 6.04008e-19 $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.12
cc_20 VNB N_A_244_137#_c_322_n 0.00505475f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.95
cc_21 VNB N_A_244_137#_c_323_n 0.011456f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.95
cc_22 VNB N_A_754_367#_M1000_g 0.0373199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_754_367#_c_385_n 0.071246f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.705
cc_24 VNB N_A_754_367#_c_386_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.295
cc_25 VNB N_A_754_367#_M1008_g 0.00832643f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=0.62
cc_26 VNB N_A_754_367#_M1001_g 0.0417898f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.95
cc_27 VNB N_A_754_367#_c_389_n 0.0184075f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_28 VNB N_A_754_367#_c_390_n 0.00779566f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.295
cc_29 VNB N_A_754_367#_c_391_n 0.00307974f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_30 VNB N_A_754_367#_c_392_n 0.00330803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_754_367#_c_393_n 0.0378451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_M1002_g 0.0269235f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.625
cc_33 VNB N_B_c_500_n 0.0199589f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_34 VNB N_B_M1004_g 0.0276903f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.12
cc_35 VNB N_B_M1007_g 0.0419532f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.625
cc_36 VNB N_B_c_503_n 0.00363501f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.035
cc_37 VNB N_B_c_504_n 0.00956473f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.765
cc_38 VNB N_B_c_505_n 0.0310399f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.625
cc_39 VNB N_B_c_506_n 0.0017732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_M1003_g 0.0233906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_M1018_g 0.00890692f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.625
cc_42 VNB A 0.00468049f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_43 VNB N_A_c_632_n 0.0286655f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.685
cc_44 VNB N_A_871_373#_M1015_g 0.0291693f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.705
cc_45 VNB N_A_871_373#_M1005_g 0.00802354f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=0.62
cc_46 VNB N_A_871_373#_c_681_n 0.0235101f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.95
cc_47 VNB N_A_871_373#_c_682_n 0.00223267f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.295
cc_48 VNB N_A_871_373#_c_683_n 0.00390434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_871_373#_c_684_n 0.00540028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_871_373#_c_685_n 0.0354638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_871_373#_c_686_n 0.00340132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_X_c_801_n 0.0245825f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.705
cc_53 VNB X 0.0122585f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.625
cc_54 VNB N_X_c_803_n 0.029348f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.95
cc_55 VNB N_VPWR_c_823_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.625
cc_56 VNB N_A_355_451#_c_901_n 0.0119806f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.62
cc_57 VNB N_A_355_451#_c_902_n 0.0141472f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.865
cc_58 VNB N_A_355_451#_c_903_n 0.00228752f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_59 VNB N_A_355_451#_c_904_n 0.00973476f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.765
cc_60 VNB N_A_355_451#_c_905_n 7.89398e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_354_109#_c_1037_n 0.00529317f $X=-0.19 $Y=-0.245 $X2=2.245
+ $Y2=0.62
cc_62 VNB N_A_354_109#_c_1038_n 0.0105359f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.12
cc_63 VNB N_A_354_109#_c_1039_n 0.00638811f $X=-0.19 $Y=-0.245 $X2=1.035
+ $Y2=2.865
cc_64 VNB N_A_354_109#_c_1040_n 4.46741e-19 $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.95
cc_65 VNB N_A_354_109#_c_1041_n 0.00122885f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_66 VNB N_A_354_109#_c_1042_n 0.00737405f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_67 VNB N_A_354_109#_c_1043_n 0.034226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_354_109#_c_1044_n 0.0030999f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.62
cc_69 VNB N_A_354_109#_c_1045_n 0.0018135f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.625
cc_70 VNB N_A_1090_373#_c_1141_n 0.0139513f $X=-0.19 $Y=-0.245 $X2=0.695
+ $Y2=0.705
cc_71 VNB N_A_1090_373#_c_1142_n 0.00235852f $X=-0.19 $Y=-0.245 $X2=0.695
+ $Y2=1.95
cc_72 VNB N_A_1090_373#_c_1143_n 0.0228529f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.95
cc_73 VNB N_A_1090_373#_c_1144_n 0.004114f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.46
cc_74 VNB N_A_1090_373#_c_1145_n 8.47722e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1090_373#_c_1146_n 0.0114231f $X=-0.19 $Y=-0.245 $X2=1.035
+ $Y2=2.035
cc_76 VNB N_A_1090_373#_c_1147_n 0.0319635f $X=-0.19 $Y=-0.245 $X2=2.41
+ $Y2=0.765
cc_77 VNB N_VGND_c_1249_n 0.0138784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1250_n 0.00912322f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.95
cc_79 VNB N_VGND_c_1251_n 0.0827263f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.12
cc_80 VNB N_VGND_c_1252_n 0.00631837f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.865
cc_81 VNB N_VGND_c_1253_n 0.0623852f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.95
cc_82 VNB N_VGND_c_1254_n 0.0218847f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.765
cc_83 VNB N_VGND_c_1255_n 0.437587f $X=-0.19 $Y=-0.245 $X2=2.41 $Y2=0.765
cc_84 VNB N_VGND_c_1256_n 0.0354693f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.625
cc_85 VNB N_VGND_c_1257_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VPB N_A_81_259#_M1020_g 0.0265497f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_87 VPB N_A_81_259#_c_160_n 0.00297631f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.95
cc_88 VPB N_A_81_259#_c_168_n 0.012027f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.865
cc_89 VPB N_A_81_259#_c_169_n 0.00357423f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.95
cc_90 VPB N_A_81_259#_c_170_n 0.0232634f $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.95
cc_91 VPB N_C_M1014_g 0.0230855f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.625
cc_92 VPB N_C_M1011_g 0.0525786f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.625
cc_93 VPB N_C_c_253_n 0.0066751f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.865
cc_94 VPB N_C_c_254_n 0.00471071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_244_137#_M1016_g 0.0225781f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.685
cc_96 VPB N_A_244_137#_c_321_n 0.0168878f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.12
cc_97 VPB N_A_244_137#_c_322_n 0.014288f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.95
cc_98 VPB N_A_244_137#_c_323_n 0.0222005f $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.95
cc_99 VPB N_A_754_367#_M1012_g 0.0210757f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_100 VPB N_A_754_367#_M1008_g 0.0216325f $X=-0.19 $Y=1.655 $X2=2.245 $Y2=0.62
cc_101 VPB N_A_754_367#_c_390_n 0.00143665f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.295
cc_102 VPB N_A_754_367#_c_397_n 0.00326551f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.625
cc_103 VPB N_A_754_367#_c_398_n 0.00241234f $X=-0.19 $Y=1.655 $X2=1.035
+ $Y2=2.035
cc_104 VPB N_A_754_367#_c_399_n 8.99775e-19 $X=-0.19 $Y=1.655 $X2=2.41 $Y2=0.765
cc_105 VPB N_A_754_367#_c_392_n 0.00161385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_754_367#_c_393_n 0.0117573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_B_M1021_g 0.0224788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_B_c_500_n 0.00522803f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_109 VPB N_B_c_509_n 0.0804008f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.685
cc_110 VPB N_B_c_510_n 0.0678146f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.685
cc_111 VPB N_B_c_511_n 0.0100054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_B_M1017_g 0.0483219f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.95
cc_113 VPB N_B_c_513_n 0.0746931f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.95
cc_114 VPB N_B_M1013_g 0.0388612f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.46
cc_115 VPB N_B_c_503_n 0.00680233f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.035
cc_116 VPB N_B_c_516_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_B_c_504_n 0.00733062f $X=-0.19 $Y=1.655 $X2=2.41 $Y2=0.765
cc_118 VPB N_B_c_505_n 0.00468161f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.625
cc_119 VPB N_B_c_506_n 0.00401429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_M1018_g 0.0275196f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.625
cc_121 VPB N_A_871_373#_M1005_g 0.0316312f $X=-0.19 $Y=1.655 $X2=2.245 $Y2=0.62
cc_122 VPB N_A_871_373#_c_688_n 0.0369721f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.12
cc_123 VPB N_A_871_373#_c_689_n 0.0105015f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.46
cc_124 VPB N_A_871_373#_c_690_n 0.00188369f $X=-0.19 $Y=1.655 $X2=0.695
+ $Y2=2.035
cc_125 VPB N_A_871_373#_c_691_n 0.00808616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_871_373#_c_682_n 0.00395774f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.295
cc_127 VPB N_A_871_373#_c_693_n 0.00978916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_X_c_804_n 0.0081627f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_129 VPB N_X_c_805_n 0.042522f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.295
cc_130 VPB N_X_c_801_n 0.00759794f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=0.705
cc_131 VPB N_VPWR_c_824_n 0.00240024f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.685
cc_132 VPB N_VPWR_c_825_n 0.00814293f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.295
cc_133 VPB N_VPWR_c_826_n 0.00892355f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.62
cc_134 VPB N_VPWR_c_827_n 0.0867021f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.95
cc_135 VPB N_VPWR_c_828_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.95
cc_136 VPB N_VPWR_c_829_n 0.015629f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_137 VPB N_VPWR_c_830_n 0.0634919f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.035
cc_138 VPB N_VPWR_c_831_n 0.0207606f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.295
cc_139 VPB N_VPWR_c_823_n 0.0849448f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.625
cc_140 VPB N_VPWR_c_833_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_834_n 0.00510127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_355_451#_c_906_n 0.00297234f $X=-0.19 $Y=1.655 $X2=0.695
+ $Y2=0.705
cc_143 VPB N_A_355_451#_c_907_n 0.00625075f $X=-0.19 $Y=1.655 $X2=0.695
+ $Y2=1.625
cc_144 VPB N_A_355_451#_c_901_n 0.0105771f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.62
cc_145 VPB N_A_355_451#_c_909_n 0.00369969f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.95
cc_146 VPB N_A_355_451#_c_910_n 0.00355932f $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.95
cc_147 VPB N_A_355_451#_c_911_n 0.00616001f $X=-0.19 $Y=1.655 $X2=1.035
+ $Y2=2.035
cc_148 VPB N_A_354_109#_c_1037_n 0.00804255f $X=-0.19 $Y=1.655 $X2=2.245
+ $Y2=0.62
cc_149 VPB N_A_354_109#_c_1040_n 0.00376233f $X=-0.19 $Y=1.655 $X2=2.34 $Y2=2.95
cc_150 VPB N_A_1090_373#_c_1148_n 0.00476697f $X=-0.19 $Y=1.655 $X2=0.49
+ $Y2=0.685
cc_151 VPB N_A_1090_373#_c_1149_n 0.00223847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_1090_373#_c_1150_n 0.00128196f $X=-0.19 $Y=1.655 $X2=0.78
+ $Y2=0.62
cc_153 VPB N_A_1090_373#_c_1151_n 0.0114989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_1090_373#_c_1147_n 0.0118607f $X=-0.19 $Y=1.655 $X2=2.41
+ $Y2=0.765
cc_155 VPB N_A_1090_373#_c_1153_n 0.0377127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_1090_373#_c_1154_n 0.0027702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 N_A_81_259#_M1019_g N_C_M1006_g 0.0113372f $X=0.49 $Y=0.685 $X2=0 $Y2=0
cc_158 N_A_81_259#_c_161_n N_C_M1006_g 0.0141776f $X=2.245 $Y=0.62 $X2=0 $Y2=0
cc_159 N_A_81_259#_c_163_n N_C_M1006_g 0.00162617f $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_160 N_A_81_259#_c_164_n N_C_M1006_g 0.0098163f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_161 N_A_81_259#_M1020_g N_C_M1014_g 0.0118766f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_81_259#_c_160_n N_C_M1014_g 0.00367621f $X=0.695 $Y=1.95 $X2=0 $Y2=0
cc_163 N_A_81_259#_c_168_n N_C_M1014_g 0.01528f $X=1.035 $Y=2.865 $X2=0 $Y2=0
cc_164 N_A_81_259#_c_170_n N_C_M1014_g 0.00431838f $X=2.34 $Y=2.95 $X2=0 $Y2=0
cc_165 N_A_81_259#_c_179_p N_C_M1014_g 0.0053908f $X=1.035 $Y=2.035 $X2=0 $Y2=0
cc_166 N_A_81_259#_c_161_n N_C_c_249_n 0.00461816f $X=2.245 $Y=0.62 $X2=0 $Y2=0
cc_167 N_A_81_259#_c_161_n N_C_M1010_g 0.0129392f $X=2.245 $Y=0.62 $X2=0 $Y2=0
cc_168 N_A_81_259#_c_165_n N_C_M1010_g 7.56449e-19 $X=2.41 $Y=0.62 $X2=0 $Y2=0
cc_169 N_A_81_259#_c_170_n N_C_M1011_g 0.00999283f $X=2.34 $Y=2.95 $X2=0 $Y2=0
cc_170 N_A_81_259#_M1020_g N_C_c_253_n 8.77977e-19 $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A_81_259#_c_162_n N_C_c_253_n 0.00237623f $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_172 N_A_81_259#_c_163_n N_C_c_253_n 0.0120679f $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_173 N_A_81_259#_c_179_p N_C_c_253_n 2.15032e-19 $X=1.035 $Y=2.035 $X2=0 $Y2=0
cc_174 N_A_81_259#_c_161_n N_C_c_254_n 0.00360792f $X=2.245 $Y=0.62 $X2=0 $Y2=0
cc_175 N_A_81_259#_c_162_n N_C_c_254_n 0.0259512f $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_176 N_A_81_259#_c_163_n N_C_c_254_n 3.35357e-19 $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_177 N_A_81_259#_c_179_p N_C_c_254_n 0.00521588f $X=1.035 $Y=2.035 $X2=0 $Y2=0
cc_178 N_A_81_259#_c_161_n N_A_244_137#_M1006_d 0.0023192f $X=2.245 $Y=0.62
+ $X2=-0.19 $Y2=-0.245
cc_179 N_A_81_259#_c_165_n N_A_244_137#_M1009_g 0.0069702f $X=2.41 $Y=0.62 $X2=0
+ $Y2=0
cc_180 N_A_81_259#_c_170_n N_A_244_137#_M1016_g 0.0047198f $X=2.34 $Y=2.95 $X2=0
+ $Y2=0
cc_181 N_A_81_259#_c_161_n N_A_244_137#_c_319_n 0.0315404f $X=2.245 $Y=0.62
+ $X2=0 $Y2=0
cc_182 N_A_81_259#_c_164_n N_A_244_137#_c_319_n 0.00947787f $X=0.61 $Y=1.295
+ $X2=0 $Y2=0
cc_183 N_A_81_259#_c_168_n N_A_244_137#_c_321_n 0.0135758f $X=1.035 $Y=2.865
+ $X2=0 $Y2=0
cc_184 N_A_81_259#_c_170_n N_A_244_137#_c_321_n 0.0153442f $X=2.34 $Y=2.95 $X2=0
+ $Y2=0
cc_185 N_A_81_259#_M1020_g N_X_c_804_n 0.00334092f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_81_259#_c_160_n N_X_c_804_n 0.00109453f $X=0.695 $Y=1.95 $X2=0 $Y2=0
cc_187 N_A_81_259#_M1019_g N_X_c_801_n 0.00365947f $X=0.49 $Y=0.685 $X2=0 $Y2=0
cc_188 N_A_81_259#_c_160_n N_X_c_801_n 0.00878088f $X=0.695 $Y=1.95 $X2=0 $Y2=0
cc_189 N_A_81_259#_c_162_n N_X_c_801_n 0.0248573f $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_190 N_A_81_259#_c_163_n N_X_c_801_n 0.011854f $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_191 N_A_81_259#_c_164_n N_X_c_801_n 0.00785193f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_192 N_A_81_259#_M1019_g X 0.00340332f $X=0.49 $Y=0.685 $X2=0 $Y2=0
cc_193 N_A_81_259#_c_163_n X 4.83855e-19 $X=0.57 $Y=1.46 $X2=0 $Y2=0
cc_194 N_A_81_259#_M1019_g N_X_c_803_n 0.0164689f $X=0.49 $Y=0.685 $X2=0 $Y2=0
cc_195 N_A_81_259#_c_164_n N_X_c_803_n 0.0165087f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_196 N_A_81_259#_c_160_n N_VPWR_M1020_d 0.00304226f $X=0.695 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_81_259#_c_168_n N_VPWR_M1020_d 0.00459015f $X=1.035 $Y=2.865
+ $X2=-0.19 $Y2=-0.245
cc_198 N_A_81_259#_c_179_p N_VPWR_M1020_d 0.0210977f $X=1.035 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_81_259#_M1020_g N_VPWR_c_824_n 0.0175594f $X=0.48 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_81_259#_c_168_n N_VPWR_c_824_n 0.0434875f $X=1.035 $Y=2.865 $X2=0
+ $Y2=0
cc_201 N_A_81_259#_c_169_n N_VPWR_c_824_n 0.0145003f $X=1.12 $Y=2.95 $X2=0 $Y2=0
cc_202 N_A_81_259#_c_162_n N_VPWR_c_824_n 0.00126179f $X=0.57 $Y=1.46 $X2=0
+ $Y2=0
cc_203 N_A_81_259#_c_179_p N_VPWR_c_824_n 0.0135869f $X=1.035 $Y=2.035 $X2=0
+ $Y2=0
cc_204 N_A_81_259#_M1020_g N_VPWR_c_829_n 0.00486043f $X=0.48 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_A_81_259#_c_169_n N_VPWR_c_830_n 0.00971923f $X=1.12 $Y=2.95 $X2=0
+ $Y2=0
cc_206 N_A_81_259#_c_170_n N_VPWR_c_830_n 0.0678664f $X=2.34 $Y=2.95 $X2=0 $Y2=0
cc_207 N_A_81_259#_M1011_d N_VPWR_c_823_n 0.0023412f $X=2.2 $Y=2.255 $X2=0 $Y2=0
cc_208 N_A_81_259#_M1020_g N_VPWR_c_823_n 0.00918457f $X=0.48 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_A_81_259#_c_169_n N_VPWR_c_823_n 0.00647808f $X=1.12 $Y=2.95 $X2=0
+ $Y2=0
cc_210 N_A_81_259#_c_170_n N_VPWR_c_823_n 0.0500311f $X=2.34 $Y=2.95 $X2=0 $Y2=0
cc_211 N_A_81_259#_c_170_n N_A_355_451#_M1011_s 0.00679513f $X=2.34 $Y=2.95
+ $X2=0 $Y2=0
cc_212 N_A_81_259#_M1011_d N_A_355_451#_c_907_n 0.00888391f $X=2.2 $Y=2.255
+ $X2=0 $Y2=0
cc_213 N_A_81_259#_c_170_n N_A_355_451#_c_907_n 0.0250481f $X=2.34 $Y=2.95 $X2=0
+ $Y2=0
cc_214 N_A_81_259#_c_170_n N_A_355_451#_c_915_n 0.0142188f $X=2.34 $Y=2.95 $X2=0
+ $Y2=0
cc_215 N_A_81_259#_c_165_n N_A_355_451#_c_902_n 0.0190793f $X=2.41 $Y=0.62 $X2=0
+ $Y2=0
cc_216 N_A_81_259#_c_161_n N_A_354_109#_M1010_s 0.00349817f $X=2.245 $Y=0.62
+ $X2=-0.19 $Y2=-0.245
cc_217 N_A_81_259#_c_161_n N_A_354_109#_c_1049_n 0.0150184f $X=2.245 $Y=0.62
+ $X2=0 $Y2=0
cc_218 N_A_81_259#_M1010_d N_A_354_109#_c_1042_n 0.00252325f $X=2.2 $Y=0.545
+ $X2=0 $Y2=0
cc_219 N_A_81_259#_c_161_n N_A_354_109#_c_1042_n 0.00371431f $X=2.245 $Y=0.62
+ $X2=0 $Y2=0
cc_220 N_A_81_259#_c_165_n N_A_354_109#_c_1042_n 0.0214744f $X=2.41 $Y=0.62
+ $X2=0 $Y2=0
cc_221 N_A_81_259#_c_165_n N_A_354_109#_c_1044_n 0.00212153f $X=2.41 $Y=0.62
+ $X2=0 $Y2=0
cc_222 N_A_81_259#_c_161_n N_VGND_M1019_d 0.0116534f $X=2.245 $Y=0.62 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_81_259#_c_237_p N_VGND_M1019_d 0.00327702f $X=0.78 $Y=0.62 $X2=-0.19
+ $Y2=-0.245
cc_224 N_A_81_259#_c_164_n N_VGND_M1019_d 0.0085574f $X=0.61 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A_81_259#_c_161_n N_VGND_c_1253_n 0.0286737f $X=2.245 $Y=0.62 $X2=0
+ $Y2=0
cc_226 N_A_81_259#_c_165_n N_VGND_c_1253_n 0.00824997f $X=2.41 $Y=0.62 $X2=0
+ $Y2=0
cc_227 N_A_81_259#_M1019_g N_VGND_c_1255_n 0.0116231f $X=0.49 $Y=0.685 $X2=0
+ $Y2=0
cc_228 N_A_81_259#_c_161_n N_VGND_c_1255_n 0.0400247f $X=2.245 $Y=0.62 $X2=0
+ $Y2=0
cc_229 N_A_81_259#_c_237_p N_VGND_c_1255_n 0.00215545f $X=0.78 $Y=0.62 $X2=0
+ $Y2=0
cc_230 N_A_81_259#_c_165_n N_VGND_c_1255_n 0.0106026f $X=2.41 $Y=0.62 $X2=0
+ $Y2=0
cc_231 N_A_81_259#_M1019_g N_VGND_c_1256_n 0.0116681f $X=0.49 $Y=0.685 $X2=0
+ $Y2=0
cc_232 N_A_81_259#_c_161_n N_VGND_c_1256_n 0.0146677f $X=2.245 $Y=0.62 $X2=0
+ $Y2=0
cc_233 N_A_81_259#_c_237_p N_VGND_c_1256_n 0.0113155f $X=0.78 $Y=0.62 $X2=0
+ $Y2=0
cc_234 N_C_M1010_g N_A_244_137#_M1009_g 0.0328214f $X=2.125 $Y=0.865 $X2=0 $Y2=0
cc_235 N_C_M1011_g N_A_244_137#_M1016_g 0.0309529f $X=2.125 $Y=2.675 $X2=0 $Y2=0
cc_236 N_C_M1006_g N_A_244_137#_c_319_n 0.00513609f $X=1.145 $Y=0.895 $X2=0
+ $Y2=0
cc_237 N_C_c_253_n N_A_244_137#_c_319_n 0.00590429f $X=1.19 $Y=1.42 $X2=0 $Y2=0
cc_238 N_C_c_254_n N_A_244_137#_c_319_n 0.0076841f $X=1.19 $Y=1.51 $X2=0 $Y2=0
cc_239 N_C_M1006_g N_A_244_137#_c_320_n 0.00677201f $X=1.145 $Y=0.895 $X2=0
+ $Y2=0
cc_240 N_C_c_249_n N_A_244_137#_c_320_n 0.0173732f $X=2.05 $Y=1.42 $X2=0 $Y2=0
cc_241 N_C_M1010_g N_A_244_137#_c_320_n 7.6185e-19 $X=2.125 $Y=0.865 $X2=0 $Y2=0
cc_242 N_C_M1011_g N_A_244_137#_c_320_n 0.0010898f $X=2.125 $Y=2.675 $X2=0 $Y2=0
cc_243 N_C_c_253_n N_A_244_137#_c_320_n 6.90109e-19 $X=1.19 $Y=1.42 $X2=0 $Y2=0
cc_244 N_C_c_254_n N_A_244_137#_c_320_n 0.015029f $X=1.19 $Y=1.51 $X2=0 $Y2=0
cc_245 N_C_M1014_g N_A_244_137#_c_321_n 0.00972533f $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_246 N_C_c_249_n N_A_244_137#_c_321_n 0.00380226f $X=2.05 $Y=1.42 $X2=0 $Y2=0
cc_247 N_C_M1011_g N_A_244_137#_c_321_n 0.0107514f $X=2.125 $Y=2.675 $X2=0 $Y2=0
cc_248 N_C_c_253_n N_A_244_137#_c_321_n 0.00320802f $X=1.19 $Y=1.42 $X2=0 $Y2=0
cc_249 N_C_c_254_n N_A_244_137#_c_321_n 0.0212441f $X=1.19 $Y=1.51 $X2=0 $Y2=0
cc_250 N_C_c_249_n N_A_244_137#_c_322_n 0.0128003f $X=2.05 $Y=1.42 $X2=0 $Y2=0
cc_251 N_C_M1011_g N_A_244_137#_c_322_n 0.0209879f $X=2.125 $Y=2.675 $X2=0 $Y2=0
cc_252 N_C_M1011_g N_A_244_137#_c_323_n 0.0213346f $X=2.125 $Y=2.675 $X2=0 $Y2=0
cc_253 N_C_M1014_g N_VPWR_c_824_n 9.14078e-19 $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_254 N_C_M1011_g N_VPWR_c_830_n 0.00366111f $X=2.125 $Y=2.675 $X2=0 $Y2=0
cc_255 N_C_M1011_g N_VPWR_c_823_n 0.00806346f $X=2.125 $Y=2.675 $X2=0 $Y2=0
cc_256 N_C_M1014_g N_A_355_451#_c_906_n 9.72484e-19 $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_257 N_C_M1011_g N_A_355_451#_c_906_n 0.00678071f $X=2.125 $Y=2.675 $X2=0
+ $Y2=0
cc_258 N_C_M1011_g N_A_355_451#_c_907_n 0.00968645f $X=2.125 $Y=2.675 $X2=0
+ $Y2=0
cc_259 N_C_M1014_g N_A_355_451#_c_915_n 0.00212542f $X=1.16 $Y=2.155 $X2=0 $Y2=0
cc_260 N_C_M1011_g N_A_355_451#_c_915_n 0.00138548f $X=2.125 $Y=2.675 $X2=0
+ $Y2=0
cc_261 N_C_M1006_g N_A_354_109#_c_1049_n 3.77434e-19 $X=1.145 $Y=0.895 $X2=0
+ $Y2=0
cc_262 N_C_M1010_g N_A_354_109#_c_1049_n 0.00487813f $X=2.125 $Y=0.865 $X2=0
+ $Y2=0
cc_263 N_C_c_249_n N_A_354_109#_c_1041_n 0.0061982f $X=2.05 $Y=1.42 $X2=0 $Y2=0
cc_264 N_C_M1010_g N_A_354_109#_c_1041_n 0.00336487f $X=2.125 $Y=0.865 $X2=0
+ $Y2=0
cc_265 N_C_c_252_n N_A_354_109#_c_1041_n 4.37774e-19 $X=2.125 $Y=1.42 $X2=0
+ $Y2=0
cc_266 N_C_M1010_g N_A_354_109#_c_1042_n 0.00718423f $X=2.125 $Y=0.865 $X2=0
+ $Y2=0
cc_267 N_C_c_252_n N_A_354_109#_c_1042_n 0.00272336f $X=2.125 $Y=1.42 $X2=0
+ $Y2=0
cc_268 N_C_M1010_g N_A_354_109#_c_1044_n 4.10504e-19 $X=2.125 $Y=0.865 $X2=0
+ $Y2=0
cc_269 N_C_M1006_g N_VGND_c_1253_n 6.43532e-19 $X=1.145 $Y=0.895 $X2=0 $Y2=0
cc_270 N_C_M1010_g N_VGND_c_1253_n 0.0034654f $X=2.125 $Y=0.865 $X2=0 $Y2=0
cc_271 N_C_M1010_g N_VGND_c_1255_n 0.00492109f $X=2.125 $Y=0.865 $X2=0 $Y2=0
cc_272 N_A_244_137#_M1016_g N_VPWR_c_825_n 0.0036689f $X=2.67 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_A_244_137#_M1016_g N_VPWR_c_830_n 0.00401801f $X=2.67 $Y=2.465 $X2=0
+ $Y2=0
cc_274 N_A_244_137#_M1016_g N_VPWR_c_823_n 0.0052212f $X=2.67 $Y=2.465 $X2=0
+ $Y2=0
cc_275 N_A_244_137#_M1016_g N_A_355_451#_c_906_n 0.00134279f $X=2.67 $Y=2.465
+ $X2=0 $Y2=0
cc_276 N_A_244_137#_c_321_n N_A_355_451#_c_906_n 0.0211225f $X=1.655 $Y=1.72
+ $X2=0 $Y2=0
cc_277 N_A_244_137#_c_322_n N_A_355_451#_c_906_n 0.0126771f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_278 N_A_244_137#_M1016_g N_A_355_451#_c_907_n 0.0171856f $X=2.67 $Y=2.465
+ $X2=0 $Y2=0
cc_279 N_A_244_137#_c_322_n N_A_355_451#_c_907_n 0.0141558f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_280 N_A_244_137#_c_323_n N_A_355_451#_c_907_n 0.00281036f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_281 N_A_244_137#_M1009_g N_A_355_451#_c_901_n 0.00512668f $X=2.625 $Y=0.865
+ $X2=0 $Y2=0
cc_282 N_A_244_137#_M1016_g N_A_355_451#_c_901_n 0.00512877f $X=2.67 $Y=2.465
+ $X2=0 $Y2=0
cc_283 N_A_244_137#_M1009_g N_A_355_451#_c_902_n 0.00946614f $X=2.625 $Y=0.865
+ $X2=0 $Y2=0
cc_284 N_A_244_137#_M1016_g N_A_355_451#_c_911_n 4.44828e-19 $X=2.67 $Y=2.465
+ $X2=0 $Y2=0
cc_285 N_A_244_137#_M1009_g N_A_354_109#_c_1049_n 8.59078e-19 $X=2.625 $Y=0.865
+ $X2=0 $Y2=0
cc_286 N_A_244_137#_c_319_n N_A_354_109#_c_1049_n 0.0206636f $X=1.485 $Y=1 $X2=0
+ $Y2=0
cc_287 N_A_244_137#_c_320_n N_A_354_109#_c_1049_n 0.00411073f $X=1.57 $Y=1.555
+ $X2=0 $Y2=0
cc_288 N_A_244_137#_M1009_g N_A_354_109#_c_1037_n 0.0059287f $X=2.625 $Y=0.865
+ $X2=0 $Y2=0
cc_289 N_A_244_137#_c_322_n N_A_354_109#_c_1037_n 0.0262099f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_290 N_A_244_137#_c_323_n N_A_354_109#_c_1037_n 0.020008f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_291 N_A_244_137#_c_320_n N_A_354_109#_c_1041_n 0.0169738f $X=1.57 $Y=1.555
+ $X2=0 $Y2=0
cc_292 N_A_244_137#_c_322_n N_A_354_109#_c_1041_n 0.0203863f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_293 N_A_244_137#_M1009_g N_A_354_109#_c_1042_n 0.0147106f $X=2.625 $Y=0.865
+ $X2=0 $Y2=0
cc_294 N_A_244_137#_c_322_n N_A_354_109#_c_1042_n 0.0431772f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_295 N_A_244_137#_c_323_n N_A_354_109#_c_1042_n 0.00483958f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_296 N_A_244_137#_M1009_g N_A_354_109#_c_1044_n 0.0084367f $X=2.625 $Y=0.865
+ $X2=0 $Y2=0
cc_297 N_A_244_137#_c_322_n N_A_354_109#_c_1044_n 0.00434951f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_298 N_A_244_137#_c_323_n N_A_354_109#_c_1044_n 0.0027957f $X=2.575 $Y=1.72
+ $X2=0 $Y2=0
cc_299 N_A_244_137#_M1009_g N_VGND_c_1249_n 7.08668e-19 $X=2.625 $Y=0.865 $X2=0
+ $Y2=0
cc_300 N_A_244_137#_M1009_g N_VGND_c_1253_n 0.00441768f $X=2.625 $Y=0.865 $X2=0
+ $Y2=0
cc_301 N_A_244_137#_M1009_g N_VGND_c_1255_n 0.00492109f $X=2.625 $Y=0.865 $X2=0
+ $Y2=0
cc_302 N_A_754_367#_c_390_n N_B_M1021_g 0.00156901f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_303 N_A_754_367#_c_399_n N_B_M1021_g 0.00477187f $X=4.185 $Y=2.075 $X2=0
+ $Y2=0
cc_304 N_A_754_367#_c_390_n N_B_M1002_g 0.00605717f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_305 N_A_754_367#_c_391_n N_B_M1002_g 0.00386051f $X=4.015 $Y=1.04 $X2=0 $Y2=0
cc_306 N_A_754_367#_c_390_n N_B_c_500_n 0.00997133f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_307 N_A_754_367#_c_391_n N_B_c_500_n 0.0034492f $X=4.015 $Y=1.04 $X2=0 $Y2=0
cc_308 N_A_754_367#_c_392_n N_B_c_500_n 7.39742e-19 $X=4.655 $Y=1.54 $X2=0 $Y2=0
cc_309 N_A_754_367#_c_393_n N_B_c_500_n 0.0118049f $X=4.83 $Y=1.54 $X2=0 $Y2=0
cc_310 N_A_754_367#_M1012_g N_B_c_509_n 0.0229707f $X=4.83 $Y=2.285 $X2=0 $Y2=0
cc_311 N_A_754_367#_c_390_n N_B_c_509_n 0.0067109f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_312 N_A_754_367#_c_397_n N_B_c_509_n 0.00927453f $X=4.49 $Y=2.115 $X2=0 $Y2=0
cc_313 N_A_754_367#_c_398_n N_B_c_509_n 0.00271318f $X=4.575 $Y=2.03 $X2=0 $Y2=0
cc_314 N_A_754_367#_c_399_n N_B_c_509_n 0.00666007f $X=4.185 $Y=2.075 $X2=0
+ $Y2=0
cc_315 N_A_754_367#_M1012_g N_B_c_510_n 0.00737233f $X=4.83 $Y=2.285 $X2=0 $Y2=0
cc_316 N_A_754_367#_M1012_g N_B_M1017_g 0.0116783f $X=4.83 $Y=2.285 $X2=0 $Y2=0
cc_317 N_A_754_367#_M1008_g N_B_M1017_g 0.0109056f $X=5.805 $Y=2.185 $X2=0 $Y2=0
cc_318 N_A_754_367#_M1000_g N_B_M1004_g 0.0276f $X=4.905 $Y=0.945 $X2=0 $Y2=0
cc_319 N_A_754_367#_c_385_n N_B_M1004_g 0.00737859f $X=5.875 $Y=0.18 $X2=0 $Y2=0
cc_320 N_A_754_367#_M1001_g N_B_M1004_g 0.0201816f $X=5.95 $Y=0.79 $X2=0 $Y2=0
cc_321 N_A_754_367#_c_389_n N_B_M1004_g 0.0109506f $X=5.95 $Y=1.415 $X2=0 $Y2=0
cc_322 N_A_754_367#_c_393_n N_B_M1004_g 0.00186419f $X=4.83 $Y=1.54 $X2=0 $Y2=0
cc_323 N_A_754_367#_M1008_g N_B_c_513_n 0.00313411f $X=5.805 $Y=2.185 $X2=0
+ $Y2=0
cc_324 N_A_754_367#_c_385_n N_B_M1007_g 0.0265308f $X=5.875 $Y=0.18 $X2=0 $Y2=0
cc_325 N_A_754_367#_M1008_g N_B_M1007_g 9.12991e-19 $X=5.805 $Y=2.185 $X2=0
+ $Y2=0
cc_326 N_A_754_367#_M1008_g N_B_c_503_n 0.0109506f $X=5.805 $Y=2.185 $X2=0 $Y2=0
cc_327 N_A_754_367#_c_392_n N_B_c_503_n 3.97414e-19 $X=4.655 $Y=1.54 $X2=0 $Y2=0
cc_328 N_A_754_367#_c_393_n N_B_c_503_n 0.0116783f $X=4.83 $Y=1.54 $X2=0 $Y2=0
cc_329 N_A_754_367#_M1008_g N_B_c_504_n 0.0168967f $X=5.805 $Y=2.185 $X2=0 $Y2=0
cc_330 N_A_754_367#_c_399_n N_B_c_505_n 0.00507989f $X=4.185 $Y=2.075 $X2=0
+ $Y2=0
cc_331 N_A_754_367#_c_393_n N_B_c_505_n 0.00194619f $X=4.83 $Y=1.54 $X2=0 $Y2=0
cc_332 N_A_754_367#_c_390_n N_B_c_506_n 0.0324176f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_333 N_A_754_367#_c_399_n N_B_c_506_n 0.00565864f $X=4.185 $Y=2.075 $X2=0
+ $Y2=0
cc_334 N_A_754_367#_c_397_n N_A_871_373#_M1012_s 0.011836f $X=4.49 $Y=2.115
+ $X2=0 $Y2=0
cc_335 N_A_754_367#_c_398_n N_A_871_373#_M1012_s 0.00436247f $X=4.575 $Y=2.03
+ $X2=0 $Y2=0
cc_336 N_A_754_367#_M1012_g N_A_871_373#_c_688_n 0.00150696f $X=4.83 $Y=2.285
+ $X2=0 $Y2=0
cc_337 N_A_754_367#_M1008_g N_A_871_373#_c_688_n 4.90186e-19 $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_338 N_A_754_367#_M1000_g N_A_871_373#_c_681_n 0.0134795f $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_339 N_A_754_367#_c_385_n N_A_871_373#_c_681_n 0.0143559f $X=5.875 $Y=0.18
+ $X2=0 $Y2=0
cc_340 N_A_754_367#_M1001_g N_A_871_373#_c_681_n 0.0125001f $X=5.95 $Y=0.79
+ $X2=0 $Y2=0
cc_341 N_A_754_367#_M1012_g N_A_871_373#_c_693_n 0.00324719f $X=4.83 $Y=2.285
+ $X2=0 $Y2=0
cc_342 N_A_754_367#_M1000_g N_A_871_373#_c_683_n 7.70316e-19 $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_343 N_A_754_367#_M1021_d N_VPWR_c_823_n 0.00396876f $X=3.77 $Y=1.835 $X2=0
+ $Y2=0
cc_344 N_A_754_367#_c_390_n N_A_355_451#_c_901_n 0.0089317f $X=4.1 $Y=1.95 $X2=0
+ $Y2=0
cc_345 N_A_754_367#_c_399_n N_A_355_451#_c_901_n 0.00992574f $X=4.185 $Y=2.075
+ $X2=0 $Y2=0
cc_346 N_A_754_367#_c_391_n N_A_355_451#_c_901_n 0.00360118f $X=4.015 $Y=1.04
+ $X2=0 $Y2=0
cc_347 N_A_754_367#_c_391_n N_A_355_451#_c_902_n 0.00189861f $X=4.015 $Y=1.04
+ $X2=0 $Y2=0
cc_348 N_A_754_367#_M1021_d N_A_355_451#_c_909_n 0.00668987f $X=3.77 $Y=1.835
+ $X2=0 $Y2=0
cc_349 N_A_754_367#_M1012_g N_A_355_451#_c_909_n 0.0117915f $X=4.83 $Y=2.285
+ $X2=0 $Y2=0
cc_350 N_A_754_367#_c_397_n N_A_355_451#_c_909_n 0.0137412f $X=4.49 $Y=2.115
+ $X2=0 $Y2=0
cc_351 N_A_754_367#_c_399_n N_A_355_451#_c_909_n 0.0502087f $X=4.185 $Y=2.075
+ $X2=0 $Y2=0
cc_352 N_A_754_367#_c_392_n N_A_355_451#_c_909_n 0.0023023f $X=4.655 $Y=1.54
+ $X2=0 $Y2=0
cc_353 N_A_754_367#_c_393_n N_A_355_451#_c_909_n 7.29728e-19 $X=4.83 $Y=1.54
+ $X2=0 $Y2=0
cc_354 N_A_754_367#_M1012_g N_A_355_451#_c_910_n 0.0046037f $X=4.83 $Y=2.285
+ $X2=0 $Y2=0
cc_355 N_A_754_367#_M1012_g N_A_355_451#_c_943_n 0.00960332f $X=4.83 $Y=2.285
+ $X2=0 $Y2=0
cc_356 N_A_754_367#_c_397_n N_A_355_451#_c_943_n 0.0115078f $X=4.49 $Y=2.115
+ $X2=0 $Y2=0
cc_357 N_A_754_367#_c_398_n N_A_355_451#_c_943_n 0.00935411f $X=4.575 $Y=2.03
+ $X2=0 $Y2=0
cc_358 N_A_754_367#_M1001_g N_A_355_451#_c_903_n 0.0115021f $X=5.95 $Y=0.79
+ $X2=0 $Y2=0
cc_359 N_A_754_367#_M1002_d N_A_355_451#_c_904_n 0.00720902f $X=3.875 $Y=0.345
+ $X2=0 $Y2=0
cc_360 N_A_754_367#_M1000_g N_A_355_451#_c_904_n 0.00805876f $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_361 N_A_754_367#_c_391_n N_A_355_451#_c_904_n 0.019222f $X=4.015 $Y=1.04
+ $X2=0 $Y2=0
cc_362 N_A_754_367#_c_392_n N_A_355_451#_c_904_n 0.00353465f $X=4.655 $Y=1.54
+ $X2=0 $Y2=0
cc_363 N_A_754_367#_c_393_n N_A_355_451#_c_904_n 0.00146026f $X=4.83 $Y=1.54
+ $X2=0 $Y2=0
cc_364 N_A_754_367#_M1000_g N_A_355_451#_c_905_n 0.00657907f $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_365 N_A_754_367#_M1001_g N_A_355_451#_c_953_n 0.00518245f $X=5.95 $Y=0.79
+ $X2=0 $Y2=0
cc_366 N_A_754_367#_M1008_g N_A_354_109#_c_1038_n 0.0110561f $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_367 N_A_754_367#_c_389_n N_A_354_109#_c_1038_n 0.00809459f $X=5.95 $Y=1.415
+ $X2=0 $Y2=0
cc_368 N_A_754_367#_c_392_n N_A_354_109#_c_1039_n 0.0139107f $X=4.655 $Y=1.54
+ $X2=0 $Y2=0
cc_369 N_A_754_367#_c_393_n N_A_354_109#_c_1039_n 0.00372716f $X=4.83 $Y=1.54
+ $X2=0 $Y2=0
cc_370 N_A_754_367#_M1008_g N_A_354_109#_c_1040_n 0.00660777f $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_371 N_A_754_367#_M1000_g N_A_354_109#_c_1081_n 0.0122102f $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_372 N_A_754_367#_M1000_g N_A_354_109#_c_1043_n 0.00538948f $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_373 N_A_754_367#_c_390_n N_A_354_109#_c_1043_n 0.016028f $X=4.1 $Y=1.95 $X2=0
+ $Y2=0
cc_374 N_A_754_367#_c_399_n N_A_354_109#_c_1043_n 0.00606516f $X=4.185 $Y=2.075
+ $X2=0 $Y2=0
cc_375 N_A_754_367#_c_391_n N_A_354_109#_c_1043_n 0.00902348f $X=4.015 $Y=1.04
+ $X2=0 $Y2=0
cc_376 N_A_754_367#_c_392_n N_A_354_109#_c_1043_n 0.0114219f $X=4.655 $Y=1.54
+ $X2=0 $Y2=0
cc_377 N_A_754_367#_c_393_n N_A_354_109#_c_1043_n 0.00143542f $X=4.83 $Y=1.54
+ $X2=0 $Y2=0
cc_378 N_A_754_367#_M1000_g N_A_354_109#_c_1088_n 0.00241343f $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_379 N_A_754_367#_c_392_n N_A_354_109#_c_1088_n 9.29202e-19 $X=4.655 $Y=1.54
+ $X2=0 $Y2=0
cc_380 N_A_754_367#_c_393_n N_A_354_109#_c_1088_n 0.00100415f $X=4.83 $Y=1.54
+ $X2=0 $Y2=0
cc_381 N_A_754_367#_M1000_g N_A_354_109#_c_1045_n 0.00528553f $X=4.905 $Y=0.945
+ $X2=0 $Y2=0
cc_382 N_A_754_367#_c_392_n N_A_354_109#_c_1045_n 0.00547347f $X=4.655 $Y=1.54
+ $X2=0 $Y2=0
cc_383 N_A_754_367#_c_393_n N_A_354_109#_c_1045_n 0.00201052f $X=4.83 $Y=1.54
+ $X2=0 $Y2=0
cc_384 N_A_754_367#_M1008_g N_A_1090_373#_c_1148_n 0.00620628f $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_385 N_A_754_367#_M1008_g N_A_1090_373#_c_1149_n 0.00187682f $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_386 N_A_754_367#_M1001_g N_A_1090_373#_c_1141_n 0.0115819f $X=5.95 $Y=0.79
+ $X2=0 $Y2=0
cc_387 N_A_754_367#_c_389_n N_A_1090_373#_c_1141_n 0.00271571f $X=5.95 $Y=1.415
+ $X2=0 $Y2=0
cc_388 N_A_754_367#_M1008_g N_A_1090_373#_c_1142_n 3.24546e-19 $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_389 N_A_754_367#_M1001_g N_A_1090_373#_c_1142_n 0.00384234f $X=5.95 $Y=0.79
+ $X2=0 $Y2=0
cc_390 N_A_754_367#_M1001_g N_A_1090_373#_c_1144_n 0.00520007f $X=5.95 $Y=0.79
+ $X2=0 $Y2=0
cc_391 N_A_754_367#_c_389_n N_A_1090_373#_c_1144_n 0.00165782f $X=5.95 $Y=1.415
+ $X2=0 $Y2=0
cc_392 N_A_754_367#_M1008_g N_A_1090_373#_c_1145_n 0.00200133f $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_393 N_A_754_367#_M1008_g N_A_1090_373#_c_1164_n 0.00745199f $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_394 N_A_754_367#_M1012_g N_A_1090_373#_c_1154_n 4.19892e-19 $X=4.83 $Y=2.285
+ $X2=0 $Y2=0
cc_395 N_A_754_367#_M1008_g N_A_1090_373#_c_1154_n 0.00837795f $X=5.805 $Y=2.185
+ $X2=0 $Y2=0
cc_396 N_A_754_367#_c_386_n N_VGND_c_1251_n 0.0258037f $X=4.98 $Y=0.18 $X2=0
+ $Y2=0
cc_397 N_A_754_367#_c_385_n N_VGND_c_1255_n 0.0269927f $X=5.875 $Y=0.18 $X2=0
+ $Y2=0
cc_398 N_A_754_367#_c_386_n N_VGND_c_1255_n 0.00604517f $X=4.98 $Y=0.18 $X2=0
+ $Y2=0
cc_399 N_B_M1007_g N_A_M1003_g 0.0134071f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_400 N_B_M1013_g N_A_M1018_g 0.0227776f $X=6.45 $Y=2.285 $X2=0 $Y2=0
cc_401 N_B_M1007_g N_A_M1018_g 0.00595579f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_402 N_B_M1007_g A 0.00203113f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_403 N_B_M1007_g N_A_c_632_n 0.0166463f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_404 N_B_c_510_n N_A_871_373#_c_688_n 0.0103141f $X=5.3 $Y=3.15 $X2=0 $Y2=0
cc_405 N_B_M1017_g N_A_871_373#_c_688_n 0.01639f $X=5.375 $Y=2.185 $X2=0 $Y2=0
cc_406 N_B_c_513_n N_A_871_373#_c_688_n 0.0153957f $X=6.375 $Y=3.15 $X2=0 $Y2=0
cc_407 N_B_M1013_g N_A_871_373#_c_688_n 0.0132952f $X=6.45 $Y=2.285 $X2=0 $Y2=0
cc_408 N_B_M1004_g N_A_871_373#_c_681_n 0.00116683f $X=5.405 $Y=0.945 $X2=0
+ $Y2=0
cc_409 N_B_M1007_g N_A_871_373#_c_681_n 0.0137612f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_410 N_B_M1013_g N_A_871_373#_c_689_n 0.00333379f $X=6.45 $Y=2.285 $X2=0 $Y2=0
cc_411 N_B_M1013_g N_A_871_373#_c_690_n 0.0105755f $X=6.45 $Y=2.285 $X2=0 $Y2=0
cc_412 N_B_c_509_n N_A_871_373#_c_693_n 0.0133569f $X=4.205 $Y=3.075 $X2=0 $Y2=0
cc_413 N_B_c_510_n N_A_871_373#_c_693_n 0.007046f $X=5.3 $Y=3.15 $X2=0 $Y2=0
cc_414 N_B_M1017_g N_A_871_373#_c_693_n 0.00193355f $X=5.375 $Y=2.185 $X2=0
+ $Y2=0
cc_415 N_B_M1002_g N_A_871_373#_c_683_n 0.00522618f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_416 N_B_M1021_g N_VPWR_c_825_n 0.0108066f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_417 N_B_c_509_n N_VPWR_c_825_n 0.00205689f $X=4.205 $Y=3.075 $X2=0 $Y2=0
cc_418 N_B_M1013_g N_VPWR_c_826_n 0.0027318f $X=6.45 $Y=2.285 $X2=0 $Y2=0
cc_419 N_B_M1021_g N_VPWR_c_827_n 0.00486043f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_420 N_B_c_511_n N_VPWR_c_827_n 0.0545884f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_421 N_B_M1021_g N_VPWR_c_823_n 0.00472306f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_422 N_B_c_510_n N_VPWR_c_823_n 0.0243376f $X=5.3 $Y=3.15 $X2=0 $Y2=0
cc_423 N_B_c_511_n N_VPWR_c_823_n 0.00576054f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_424 N_B_c_513_n N_VPWR_c_823_n 0.0278168f $X=6.375 $Y=3.15 $X2=0 $Y2=0
cc_425 N_B_c_516_n N_VPWR_c_823_n 0.00371014f $X=5.375 $Y=3.15 $X2=0 $Y2=0
cc_426 N_B_M1021_g N_A_355_451#_c_901_n 0.0141185f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_427 N_B_M1002_g N_A_355_451#_c_901_n 0.00536253f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_428 N_B_c_505_n N_A_355_451#_c_901_n 0.00794046f $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_429 N_B_c_506_n N_A_355_451#_c_901_n 0.0329807f $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_430 N_B_M1002_g N_A_355_451#_c_902_n 0.00854083f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_431 N_B_M1021_g N_A_355_451#_c_909_n 0.0152242f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_432 N_B_c_509_n N_A_355_451#_c_909_n 0.0131984f $X=4.205 $Y=3.075 $X2=0 $Y2=0
cc_433 N_B_c_510_n N_A_355_451#_c_909_n 4.24983e-19 $X=5.3 $Y=3.15 $X2=0 $Y2=0
cc_434 N_B_c_505_n N_A_355_451#_c_909_n 2.98676e-19 $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_435 N_B_c_506_n N_A_355_451#_c_909_n 0.00585355f $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_436 N_B_c_509_n N_A_355_451#_c_910_n 7.57393e-19 $X=4.205 $Y=3.075 $X2=0
+ $Y2=0
cc_437 N_B_M1017_g N_A_355_451#_c_910_n 0.00405215f $X=5.375 $Y=2.185 $X2=0
+ $Y2=0
cc_438 N_B_c_509_n N_A_355_451#_c_943_n 9.04782e-19 $X=4.205 $Y=3.075 $X2=0
+ $Y2=0
cc_439 N_B_M1017_g N_A_355_451#_c_943_n 0.00445018f $X=5.375 $Y=2.185 $X2=0
+ $Y2=0
cc_440 N_B_M1004_g N_A_355_451#_c_903_n 0.0142268f $X=5.405 $Y=0.945 $X2=0 $Y2=0
cc_441 N_B_M1021_g N_A_355_451#_c_911_n 0.005392f $X=3.695 $Y=2.465 $X2=0 $Y2=0
cc_442 N_B_M1002_g N_A_355_451#_c_904_n 0.0171219f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_443 N_B_c_505_n N_A_355_451#_c_904_n 9.05893e-19 $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_444 N_B_c_506_n N_A_355_451#_c_904_n 0.00404934f $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_445 N_B_M1004_g N_A_355_451#_c_905_n 4.8835e-19 $X=5.405 $Y=0.945 $X2=0 $Y2=0
cc_446 N_B_M1004_g N_A_354_109#_c_1038_n 0.0116551f $X=5.405 $Y=0.945 $X2=0
+ $Y2=0
cc_447 N_B_M1007_g N_A_354_109#_c_1038_n 3.05157e-19 $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_448 N_B_c_503_n N_A_354_109#_c_1038_n 0.00754489f $X=5.39 $Y=1.755 $X2=0
+ $Y2=0
cc_449 N_B_c_504_n N_A_354_109#_c_1038_n 2.52658e-19 $X=6.54 $Y=1.63 $X2=0 $Y2=0
cc_450 N_B_c_504_n N_A_354_109#_c_1040_n 0.00209523f $X=6.54 $Y=1.63 $X2=0 $Y2=0
cc_451 N_B_M1002_g N_A_354_109#_c_1043_n 0.00572974f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_452 N_B_c_500_n N_A_354_109#_c_1043_n 0.00568412f $X=4.13 $Y=1.6 $X2=0 $Y2=0
cc_453 N_B_c_505_n N_A_354_109#_c_1043_n 0.00319431f $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_454 N_B_c_506_n N_A_354_109#_c_1043_n 0.0184615f $X=3.68 $Y=1.51 $X2=0 $Y2=0
cc_455 N_B_M1004_g N_A_354_109#_c_1045_n 0.00658191f $X=5.405 $Y=0.945 $X2=0
+ $Y2=0
cc_456 N_B_M1013_g N_A_1090_373#_c_1148_n 0.00671037f $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_457 N_B_M1017_g N_A_1090_373#_c_1149_n 0.00493539f $X=5.375 $Y=2.185 $X2=0
+ $Y2=0
cc_458 N_B_M1007_g N_A_1090_373#_c_1141_n 0.0112752f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_459 N_B_M1007_g N_A_1090_373#_c_1142_n 0.00729132f $X=6.54 $Y=0.68 $X2=0
+ $Y2=0
cc_460 N_B_M1013_g N_A_1090_373#_c_1150_n 0.0199861f $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_461 N_B_c_504_n N_A_1090_373#_c_1150_n 9.96368e-19 $X=6.54 $Y=1.63 $X2=0
+ $Y2=0
cc_462 N_B_M1004_g N_A_1090_373#_c_1144_n 0.0046255f $X=5.405 $Y=0.945 $X2=0
+ $Y2=0
cc_463 N_B_M1007_g N_A_1090_373#_c_1145_n 9.43675e-19 $X=6.54 $Y=0.68 $X2=0
+ $Y2=0
cc_464 N_B_c_504_n N_A_1090_373#_c_1145_n 0.0130109f $X=6.54 $Y=1.63 $X2=0 $Y2=0
cc_465 N_B_M1013_g N_A_1090_373#_c_1164_n 0.00568419f $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_466 N_B_c_504_n N_A_1090_373#_c_1164_n 0.0019161f $X=6.54 $Y=1.63 $X2=0 $Y2=0
cc_467 N_B_M1017_g N_A_1090_373#_c_1178_n 0.00472971f $X=5.375 $Y=2.185 $X2=0
+ $Y2=0
cc_468 N_B_M1017_g N_A_1090_373#_c_1154_n 0.00773019f $X=5.375 $Y=2.185 $X2=0
+ $Y2=0
cc_469 N_B_M1013_g N_A_1090_373#_c_1154_n 3.25743e-19 $X=6.45 $Y=2.285 $X2=0
+ $Y2=0
cc_470 N_B_c_503_n N_A_1090_373#_c_1154_n 9.27963e-19 $X=5.39 $Y=1.755 $X2=0
+ $Y2=0
cc_471 N_B_M1002_g N_VGND_c_1249_n 0.00907008f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_472 N_B_M1002_g N_VGND_c_1251_n 0.00340157f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_473 N_B_M1007_g N_VGND_c_1251_n 0.00283474f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_474 N_B_M1002_g N_VGND_c_1255_n 0.00512888f $X=3.8 $Y=0.765 $X2=0 $Y2=0
cc_475 N_B_M1007_g N_VGND_c_1255_n 0.0037669f $X=6.54 $Y=0.68 $X2=0 $Y2=0
cc_476 N_A_M1003_g N_A_871_373#_M1015_g 0.0154938f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_477 N_A_c_632_n N_A_871_373#_M1015_g 2.52004e-19 $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_478 N_A_M1018_g N_A_871_373#_M1005_g 0.0294008f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_479 N_A_M1018_g N_A_871_373#_c_688_n 0.00164434f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_480 N_A_M1003_g N_A_871_373#_c_681_n 0.00321881f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_481 N_A_M1003_g N_A_871_373#_c_720_n 0.00550663f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_482 A N_A_871_373#_c_689_n 0.00513609f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_483 N_A_c_632_n N_A_871_373#_c_689_n 0.00198334f $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_484 N_A_M1018_g N_A_871_373#_c_690_n 0.0101465f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_485 N_A_M1003_g N_A_871_373#_c_724_n 0.00943917f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_486 A N_A_871_373#_c_724_n 0.0118553f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_487 N_A_c_632_n N_A_871_373#_c_724_n 0.00274244f $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_488 N_A_M1003_g N_A_871_373#_c_727_n 7.98126e-19 $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_489 A N_A_871_373#_c_727_n 0.00436704f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_490 N_A_c_632_n N_A_871_373#_c_727_n 0.001256f $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_491 N_A_M1018_g N_A_871_373#_c_691_n 0.0198082f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_492 A N_A_871_373#_c_691_n 0.0108135f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_493 N_A_c_632_n N_A_871_373#_c_691_n 0.0021322f $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_494 N_A_M1018_g N_A_871_373#_c_682_n 0.00363864f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_495 N_A_c_632_n N_A_871_373#_c_684_n 0.00363864f $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_496 A N_A_871_373#_c_685_n 3.679e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_497 N_A_c_632_n N_A_871_373#_c_685_n 0.0213355f $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_498 N_A_M1003_g N_A_871_373#_c_686_n 0.00462885f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_499 A N_A_871_373#_c_686_n 0.0258091f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_500 N_A_c_632_n N_A_871_373#_c_686_n 0.0010524f $X=7.02 $Y=1.345 $X2=0 $Y2=0
cc_501 N_A_M1018_g N_VPWR_c_826_n 0.00986627f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_502 N_A_M1018_g N_VPWR_c_827_n 0.00452954f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_503 N_A_M1018_g N_VPWR_c_823_n 0.0044646f $X=7.11 $Y=2.415 $X2=0 $Y2=0
cc_504 N_A_M1003_g N_A_1090_373#_c_1141_n 3.55535e-19 $X=6.995 $Y=0.68 $X2=0
+ $Y2=0
cc_505 A N_A_1090_373#_c_1141_n 0.00603357f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_506 N_A_M1018_g N_A_1090_373#_c_1142_n 8.48787e-19 $X=7.11 $Y=2.415 $X2=0
+ $Y2=0
cc_507 A N_A_1090_373#_c_1142_n 0.0121613f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_508 N_A_c_632_n N_A_1090_373#_c_1142_n 2.6045e-19 $X=7.02 $Y=1.345 $X2=0
+ $Y2=0
cc_509 N_A_M1018_g N_A_1090_373#_c_1150_n 0.00109976f $X=7.11 $Y=2.415 $X2=0
+ $Y2=0
cc_510 N_A_M1003_g N_A_1090_373#_c_1143_n 9.09739e-19 $X=6.995 $Y=0.68 $X2=0
+ $Y2=0
cc_511 N_A_M1018_g N_A_1090_373#_c_1164_n 0.00797812f $X=7.11 $Y=2.415 $X2=0
+ $Y2=0
cc_512 N_A_M1018_g N_A_1090_373#_c_1153_n 7.62644e-19 $X=7.11 $Y=2.415 $X2=0
+ $Y2=0
cc_513 N_A_M1003_g N_VGND_c_1250_n 0.00345875f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_514 N_A_M1003_g N_VGND_c_1251_n 0.0043861f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_515 N_A_M1003_g N_VGND_c_1255_n 0.00453346f $X=6.995 $Y=0.68 $X2=0 $Y2=0
cc_516 N_A_871_373#_c_691_n N_VPWR_M1018_d 0.00493663f $X=7.355 $Y=2.01 $X2=0
+ $Y2=0
cc_517 N_A_871_373#_M1005_g N_VPWR_c_826_n 0.00807479f $X=7.645 $Y=2.415 $X2=0
+ $Y2=0
cc_518 N_A_871_373#_c_688_n N_VPWR_c_826_n 0.0120703f $X=6.615 $Y=2.98 $X2=0
+ $Y2=0
cc_519 N_A_871_373#_c_690_n N_VPWR_c_826_n 0.0340074f $X=6.78 $Y=2.43 $X2=0
+ $Y2=0
cc_520 N_A_871_373#_c_691_n N_VPWR_c_826_n 0.0199569f $X=7.355 $Y=2.01 $X2=0
+ $Y2=0
cc_521 N_A_871_373#_c_688_n N_VPWR_c_827_n 0.139571f $X=6.615 $Y=2.98 $X2=0
+ $Y2=0
cc_522 N_A_871_373#_c_693_n N_VPWR_c_827_n 0.0210718f $X=4.5 $Y=2.795 $X2=0
+ $Y2=0
cc_523 N_A_871_373#_M1005_g N_VPWR_c_831_n 0.00520606f $X=7.645 $Y=2.415 $X2=0
+ $Y2=0
cc_524 N_A_871_373#_M1005_g N_VPWR_c_823_n 0.005315f $X=7.645 $Y=2.415 $X2=0
+ $Y2=0
cc_525 N_A_871_373#_c_688_n N_VPWR_c_823_n 0.0779583f $X=6.615 $Y=2.98 $X2=0
+ $Y2=0
cc_526 N_A_871_373#_c_693_n N_VPWR_c_823_n 0.0111709f $X=4.5 $Y=2.795 $X2=0
+ $Y2=0
cc_527 N_A_871_373#_c_681_n N_A_355_451#_M1001_d 0.00318544f $X=6.615 $Y=0.34
+ $X2=0 $Y2=0
cc_528 N_A_871_373#_M1012_s N_A_355_451#_c_909_n 0.00819962f $X=4.355 $Y=1.865
+ $X2=0 $Y2=0
cc_529 N_A_871_373#_c_688_n N_A_355_451#_c_909_n 0.00709861f $X=6.615 $Y=2.98
+ $X2=0 $Y2=0
cc_530 N_A_871_373#_c_693_n N_A_355_451#_c_909_n 0.0247092f $X=4.5 $Y=2.795
+ $X2=0 $Y2=0
cc_531 N_A_871_373#_c_688_n N_A_355_451#_c_910_n 0.0260267f $X=6.615 $Y=2.98
+ $X2=0 $Y2=0
cc_532 N_A_871_373#_c_693_n N_A_355_451#_c_910_n 9.99622e-19 $X=4.5 $Y=2.795
+ $X2=0 $Y2=0
cc_533 N_A_871_373#_M1000_s N_A_355_451#_c_904_n 0.0104928f $X=4.43 $Y=0.215
+ $X2=0 $Y2=0
cc_534 N_A_871_373#_c_681_n N_A_355_451#_c_904_n 0.0103843f $X=6.615 $Y=0.34
+ $X2=0 $Y2=0
cc_535 N_A_871_373#_c_683_n N_A_355_451#_c_904_n 0.022946f $X=4.74 $Y=0.35 $X2=0
+ $Y2=0
cc_536 N_A_871_373#_c_681_n N_A_355_451#_c_905_n 0.0793336f $X=6.615 $Y=0.34
+ $X2=0 $Y2=0
cc_537 N_A_871_373#_c_681_n N_A_355_451#_c_953_n 0.0211422f $X=6.615 $Y=0.34
+ $X2=0 $Y2=0
cc_538 N_A_871_373#_M1000_s N_A_354_109#_c_1043_n 0.00468586f $X=4.43 $Y=0.215
+ $X2=0 $Y2=0
cc_539 N_A_871_373#_c_688_n N_A_1090_373#_c_1148_n 0.0363857f $X=6.615 $Y=2.98
+ $X2=0 $Y2=0
cc_540 N_A_871_373#_c_690_n N_A_1090_373#_c_1148_n 0.0140086f $X=6.78 $Y=2.43
+ $X2=0 $Y2=0
cc_541 N_A_871_373#_c_688_n N_A_1090_373#_c_1149_n 0.0200859f $X=6.615 $Y=2.98
+ $X2=0 $Y2=0
cc_542 N_A_871_373#_c_689_n N_A_1090_373#_c_1150_n 0.0260818f $X=6.78 $Y=2.175
+ $X2=0 $Y2=0
cc_543 N_A_871_373#_c_690_n N_A_1090_373#_c_1150_n 0.0241479f $X=6.78 $Y=2.43
+ $X2=0 $Y2=0
cc_544 N_A_871_373#_M1015_g N_A_1090_373#_c_1143_n 0.00817688f $X=7.645 $Y=0.68
+ $X2=0 $Y2=0
cc_545 N_A_871_373#_M1015_g N_A_1090_373#_c_1146_n 0.00361034f $X=7.645 $Y=0.68
+ $X2=0 $Y2=0
cc_546 N_A_871_373#_c_685_n N_A_1090_373#_c_1146_n 0.00154448f $X=7.56 $Y=1.355
+ $X2=0 $Y2=0
cc_547 N_A_871_373#_c_686_n N_A_1090_373#_c_1146_n 0.00359045f $X=7.5 $Y=1.19
+ $X2=0 $Y2=0
cc_548 N_A_871_373#_M1005_g N_A_1090_373#_c_1151_n 0.00359158f $X=7.645 $Y=2.415
+ $X2=0 $Y2=0
cc_549 N_A_871_373#_c_691_n N_A_1090_373#_c_1151_n 0.0116338f $X=7.355 $Y=2.01
+ $X2=0 $Y2=0
cc_550 N_A_871_373#_c_685_n N_A_1090_373#_c_1151_n 0.0012513f $X=7.56 $Y=1.355
+ $X2=0 $Y2=0
cc_551 N_A_871_373#_M1015_g N_A_1090_373#_c_1147_n 0.0026807f $X=7.645 $Y=0.68
+ $X2=0 $Y2=0
cc_552 N_A_871_373#_M1005_g N_A_1090_373#_c_1147_n 0.00729087f $X=7.645 $Y=2.415
+ $X2=0 $Y2=0
cc_553 N_A_871_373#_c_682_n N_A_1090_373#_c_1147_n 0.0164784f $X=7.44 $Y=1.845
+ $X2=0 $Y2=0
cc_554 N_A_871_373#_c_684_n N_A_1090_373#_c_1147_n 0.0232021f $X=7.56 $Y=1.355
+ $X2=0 $Y2=0
cc_555 N_A_871_373#_c_685_n N_A_1090_373#_c_1147_n 0.00855199f $X=7.56 $Y=1.355
+ $X2=0 $Y2=0
cc_556 N_A_871_373#_c_686_n N_A_1090_373#_c_1147_n 0.00607787f $X=7.5 $Y=1.19
+ $X2=0 $Y2=0
cc_557 N_A_871_373#_M1013_d N_A_1090_373#_c_1164_n 0.00677677f $X=6.525 $Y=1.865
+ $X2=0 $Y2=0
cc_558 N_A_871_373#_M1005_g N_A_1090_373#_c_1164_n 0.0115321f $X=7.645 $Y=2.415
+ $X2=0 $Y2=0
cc_559 N_A_871_373#_c_688_n N_A_1090_373#_c_1164_n 0.00793215f $X=6.615 $Y=2.98
+ $X2=0 $Y2=0
cc_560 N_A_871_373#_c_690_n N_A_1090_373#_c_1164_n 0.0419918f $X=6.78 $Y=2.43
+ $X2=0 $Y2=0
cc_561 N_A_871_373#_c_691_n N_A_1090_373#_c_1164_n 0.0199617f $X=7.355 $Y=2.01
+ $X2=0 $Y2=0
cc_562 N_A_871_373#_c_688_n N_A_1090_373#_c_1178_n 0.00282038f $X=6.615 $Y=2.98
+ $X2=0 $Y2=0
cc_563 N_A_871_373#_M1005_g N_A_1090_373#_c_1153_n 0.0110729f $X=7.645 $Y=2.415
+ $X2=0 $Y2=0
cc_564 N_A_871_373#_c_724_n N_VGND_M1003_d 0.0143465f $X=7.355 $Y=0.86 $X2=0
+ $Y2=0
cc_565 N_A_871_373#_c_686_n N_VGND_M1003_d 0.00115462f $X=7.5 $Y=1.19 $X2=0
+ $Y2=0
cc_566 N_A_871_373#_M1015_g N_VGND_c_1250_n 0.00553533f $X=7.645 $Y=0.68 $X2=0
+ $Y2=0
cc_567 N_A_871_373#_c_681_n N_VGND_c_1250_n 0.0115062f $X=6.615 $Y=0.34 $X2=0
+ $Y2=0
cc_568 N_A_871_373#_c_724_n N_VGND_c_1250_n 0.0258044f $X=7.355 $Y=0.86 $X2=0
+ $Y2=0
cc_569 N_A_871_373#_c_681_n N_VGND_c_1251_n 0.0235948f $X=6.615 $Y=0.34 $X2=0
+ $Y2=0
cc_570 N_A_871_373#_c_683_n N_VGND_c_1251_n 0.140519f $X=4.74 $Y=0.35 $X2=0
+ $Y2=0
cc_571 N_A_871_373#_M1015_g N_VGND_c_1254_n 0.00441827f $X=7.645 $Y=0.68 $X2=0
+ $Y2=0
cc_572 N_A_871_373#_M1000_s N_VGND_c_1255_n 0.00255417f $X=4.43 $Y=0.215 $X2=0
+ $Y2=0
cc_573 N_A_871_373#_M1015_g N_VGND_c_1255_n 0.00855758f $X=7.645 $Y=0.68 $X2=0
+ $Y2=0
cc_574 N_A_871_373#_c_681_n N_VGND_c_1255_n 0.0127202f $X=6.615 $Y=0.34 $X2=0
+ $Y2=0
cc_575 N_A_871_373#_c_724_n N_VGND_c_1255_n 0.00992058f $X=7.355 $Y=0.86 $X2=0
+ $Y2=0
cc_576 N_A_871_373#_c_683_n N_VGND_c_1255_n 0.0772519f $X=4.74 $Y=0.35 $X2=0
+ $Y2=0
cc_577 N_X_c_805_n N_VPWR_c_829_n 0.0174494f $X=0.265 $Y=1.98 $X2=0 $Y2=0
cc_578 N_X_M1020_s N_VPWR_c_823_n 0.00410679f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_579 N_X_c_805_n N_VPWR_c_823_n 0.00963638f $X=0.265 $Y=1.98 $X2=0 $Y2=0
cc_580 N_X_c_803_n N_VGND_c_1255_n 0.0130308f $X=0.275 $Y=0.42 $X2=0 $Y2=0
cc_581 N_X_c_803_n N_VGND_c_1256_n 0.0314354f $X=0.275 $Y=0.42 $X2=0 $Y2=0
cc_582 N_VPWR_c_823_n N_A_355_451#_M1011_s 0.00226477f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_830_n N_A_355_451#_c_907_n 0.0107404f $X=3.315 $Y=3.33 $X2=0
+ $Y2=0
cc_584 N_VPWR_c_823_n N_A_355_451#_c_907_n 0.0197795f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_585 N_VPWR_M1021_s N_A_355_451#_c_901_n 0.00727384f $X=3.335 $Y=1.835 $X2=0
+ $Y2=0
cc_586 N_VPWR_M1021_s N_A_355_451#_c_909_n 0.0117446f $X=3.335 $Y=1.835 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_825_n N_A_355_451#_c_909_n 0.0106199f $X=3.48 $Y=2.95 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_823_n N_A_355_451#_c_909_n 0.0252473f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_589 N_VPWR_M1021_s N_A_355_451#_c_911_n 0.0026413f $X=3.335 $Y=1.835 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_825_n N_A_355_451#_c_911_n 0.00241991f $X=3.48 $Y=2.95 $X2=0
+ $Y2=0
cc_591 N_VPWR_c_830_n N_A_355_451#_c_911_n 0.00280522f $X=3.315 $Y=3.33 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_823_n N_A_355_451#_c_911_n 0.00440799f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_593 N_VPWR_M1018_d N_A_1090_373#_c_1164_n 0.00744031f $X=7.185 $Y=1.915 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_826_n N_A_1090_373#_c_1164_n 0.0257612f $X=7.325 $Y=2.43 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_826_n N_A_1090_373#_c_1218_n 2.9203e-19 $X=7.325 $Y=2.43 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_826_n N_A_1090_373#_c_1153_n 0.0381441f $X=7.325 $Y=2.43 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_831_n N_A_1090_373#_c_1153_n 0.0142109f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_823_n N_A_1090_373#_c_1153_n 0.0135539f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_A_355_451#_c_903_n N_A_354_109#_M1000_d 0.00209751f $X=6.115 $Y=0.68
+ $X2=0 $Y2=0
cc_600 N_A_355_451#_c_905_n N_A_354_109#_M1000_d 7.17773e-19 $X=5.08 $Y=0.69
+ $X2=0 $Y2=0
cc_601 N_A_355_451#_c_907_n N_A_354_109#_M1016_d 0.011292f $X=3.175 $Y=2.61
+ $X2=0 $Y2=0
cc_602 N_A_355_451#_c_907_n N_A_354_109#_c_1037_n 0.0136682f $X=3.175 $Y=2.61
+ $X2=0 $Y2=0
cc_603 N_A_355_451#_c_901_n N_A_354_109#_c_1037_n 0.0724917f $X=3.26 $Y=2.37
+ $X2=0 $Y2=0
cc_604 N_A_355_451#_c_943_n N_A_354_109#_c_1039_n 0.0160727f $X=5.045 $Y=2.04
+ $X2=0 $Y2=0
cc_605 N_A_355_451#_M1009_d N_A_354_109#_c_1042_n 0.00262724f $X=2.7 $Y=0.545
+ $X2=0 $Y2=0
cc_606 N_A_355_451#_c_901_n N_A_354_109#_c_1042_n 0.0153897f $X=3.26 $Y=2.37
+ $X2=0 $Y2=0
cc_607 N_A_355_451#_c_902_n N_A_354_109#_c_1042_n 0.0194915f $X=3.345 $Y=0.7
+ $X2=0 $Y2=0
cc_608 N_A_355_451#_c_903_n N_A_354_109#_c_1081_n 0.0139792f $X=6.115 $Y=0.68
+ $X2=0 $Y2=0
cc_609 N_A_355_451#_c_905_n N_A_354_109#_c_1081_n 0.00710005f $X=5.08 $Y=0.69
+ $X2=0 $Y2=0
cc_610 N_A_355_451#_c_901_n N_A_354_109#_c_1043_n 0.0252875f $X=3.26 $Y=2.37
+ $X2=0 $Y2=0
cc_611 N_A_355_451#_c_902_n N_A_354_109#_c_1043_n 0.00978294f $X=3.345 $Y=0.7
+ $X2=0 $Y2=0
cc_612 N_A_355_451#_c_943_n N_A_354_109#_c_1043_n 4.17134e-19 $X=5.045 $Y=2.04
+ $X2=0 $Y2=0
cc_613 N_A_355_451#_c_904_n N_A_354_109#_c_1043_n 0.0340249f $X=4.91 $Y=0.69
+ $X2=0 $Y2=0
cc_614 N_A_355_451#_M1009_d N_A_354_109#_c_1044_n 2.3149e-19 $X=2.7 $Y=0.545
+ $X2=0 $Y2=0
cc_615 N_A_355_451#_c_901_n N_A_354_109#_c_1044_n 3.59929e-19 $X=3.26 $Y=2.37
+ $X2=0 $Y2=0
cc_616 N_A_355_451#_c_902_n N_A_354_109#_c_1044_n 0.00112681f $X=3.345 $Y=0.7
+ $X2=0 $Y2=0
cc_617 N_A_355_451#_c_943_n N_A_354_109#_c_1088_n 0.00303583f $X=5.045 $Y=2.04
+ $X2=0 $Y2=0
cc_618 N_A_355_451#_c_903_n N_A_354_109#_c_1088_n 4.82901e-19 $X=6.115 $Y=0.68
+ $X2=0 $Y2=0
cc_619 N_A_355_451#_c_904_n N_A_354_109#_c_1088_n 9.5383e-19 $X=4.91 $Y=0.69
+ $X2=0 $Y2=0
cc_620 N_A_355_451#_c_905_n N_A_354_109#_c_1088_n 6.90726e-19 $X=5.08 $Y=0.69
+ $X2=0 $Y2=0
cc_621 N_A_355_451#_c_903_n N_A_1090_373#_M1004_d 0.00503454f $X=6.115 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_622 N_A_355_451#_c_910_n N_A_1090_373#_c_1149_n 0.0119961f $X=5.045 $Y=2.37
+ $X2=0 $Y2=0
cc_623 N_A_355_451#_c_903_n N_A_1090_373#_c_1141_n 0.0112199f $X=6.115 $Y=0.68
+ $X2=0 $Y2=0
cc_624 N_A_355_451#_c_953_n N_A_1090_373#_c_1141_n 0.0252261f $X=6.28 $Y=0.68
+ $X2=0 $Y2=0
cc_625 N_A_355_451#_c_903_n N_A_1090_373#_c_1144_n 0.0207486f $X=6.115 $Y=0.68
+ $X2=0 $Y2=0
cc_626 N_A_355_451#_c_953_n N_A_1090_373#_c_1144_n 2.46087e-19 $X=6.28 $Y=0.68
+ $X2=0 $Y2=0
cc_627 N_A_355_451#_c_910_n N_A_1090_373#_c_1178_n 0.00448337f $X=5.045 $Y=2.37
+ $X2=0 $Y2=0
cc_628 N_A_355_451#_c_943_n N_A_1090_373#_c_1178_n 0.00224094f $X=5.045 $Y=2.04
+ $X2=0 $Y2=0
cc_629 N_A_355_451#_c_910_n N_A_1090_373#_c_1154_n 0.00765064f $X=5.045 $Y=2.37
+ $X2=0 $Y2=0
cc_630 N_A_355_451#_c_943_n N_A_1090_373#_c_1154_n 0.0308497f $X=5.045 $Y=2.04
+ $X2=0 $Y2=0
cc_631 N_A_355_451#_c_901_n N_VGND_M1002_s 0.00279669f $X=3.26 $Y=2.37 $X2=0
+ $Y2=0
cc_632 N_A_355_451#_c_902_n N_VGND_M1002_s 0.0042174f $X=3.345 $Y=0.7 $X2=0
+ $Y2=0
cc_633 N_A_355_451#_c_904_n N_VGND_M1002_s 0.0106113f $X=4.91 $Y=0.69 $X2=0
+ $Y2=0
cc_634 N_A_355_451#_c_902_n N_VGND_c_1249_n 0.00332414f $X=3.345 $Y=0.7 $X2=0
+ $Y2=0
cc_635 N_A_355_451#_c_904_n N_VGND_c_1249_n 0.0218575f $X=4.91 $Y=0.69 $X2=0
+ $Y2=0
cc_636 N_A_355_451#_c_904_n N_VGND_c_1251_n 0.0132589f $X=4.91 $Y=0.69 $X2=0
+ $Y2=0
cc_637 N_A_355_451#_c_902_n N_VGND_c_1253_n 0.0131199f $X=3.345 $Y=0.7 $X2=0
+ $Y2=0
cc_638 N_A_355_451#_c_902_n N_VGND_c_1255_n 0.0179564f $X=3.345 $Y=0.7 $X2=0
+ $Y2=0
cc_639 N_A_355_451#_c_904_n N_VGND_c_1255_n 0.0241417f $X=4.91 $Y=0.69 $X2=0
+ $Y2=0
cc_640 N_A_354_109#_M1008_d N_A_1090_373#_c_1148_n 0.00431306f $X=5.88 $Y=1.865
+ $X2=0 $Y2=0
cc_641 N_A_354_109#_c_1040_n N_A_1090_373#_c_1148_n 0.010916f $X=6.02 $Y=2.095
+ $X2=0 $Y2=0
cc_642 N_A_354_109#_c_1038_n N_A_1090_373#_c_1141_n 0.0240818f $X=5.935 $Y=1.54
+ $X2=0 $Y2=0
cc_643 N_A_354_109#_c_1038_n N_A_1090_373#_c_1142_n 0.0148582f $X=5.935 $Y=1.54
+ $X2=0 $Y2=0
cc_644 N_A_354_109#_M1008_d N_A_1090_373#_c_1150_n 0.00635265f $X=5.88 $Y=1.865
+ $X2=0 $Y2=0
cc_645 N_A_354_109#_c_1038_n N_A_1090_373#_c_1144_n 0.0258547f $X=5.935 $Y=1.54
+ $X2=0 $Y2=0
cc_646 N_A_354_109#_c_1088_n N_A_1090_373#_c_1144_n 5.86627e-19 $X=5.04 $Y=1.295
+ $X2=0 $Y2=0
cc_647 N_A_354_109#_c_1045_n N_A_1090_373#_c_1144_n 0.0125846f $X=5.04 $Y=1.295
+ $X2=0 $Y2=0
cc_648 N_A_354_109#_c_1040_n N_A_1090_373#_c_1145_n 0.0529031f $X=6.02 $Y=2.095
+ $X2=0 $Y2=0
cc_649 N_A_354_109#_M1008_d N_A_1090_373#_c_1164_n 0.0115511f $X=5.88 $Y=1.865
+ $X2=0 $Y2=0
cc_650 N_A_354_109#_c_1040_n N_A_1090_373#_c_1164_n 0.0104279f $X=6.02 $Y=2.095
+ $X2=0 $Y2=0
cc_651 N_A_354_109#_c_1040_n N_A_1090_373#_c_1178_n 2.6899e-19 $X=6.02 $Y=2.095
+ $X2=0 $Y2=0
cc_652 N_A_354_109#_c_1038_n N_A_1090_373#_c_1154_n 0.0225811f $X=5.935 $Y=1.54
+ $X2=0 $Y2=0
cc_653 N_A_354_109#_c_1040_n N_A_1090_373#_c_1154_n 0.0187216f $X=6.02 $Y=2.095
+ $X2=0 $Y2=0
cc_654 N_A_1090_373#_c_1143_n N_VGND_c_1250_n 0.0154946f $X=7.86 $Y=0.505 $X2=0
+ $Y2=0
cc_655 N_A_1090_373#_c_1143_n N_VGND_c_1254_n 0.017498f $X=7.86 $Y=0.505 $X2=0
+ $Y2=0
cc_656 N_A_1090_373#_c_1143_n N_VGND_c_1255_n 0.0139289f $X=7.86 $Y=0.505 $X2=0
+ $Y2=0
