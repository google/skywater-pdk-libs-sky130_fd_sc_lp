# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.210000 2.315000 1.390000 ;
        RECT 2.030000 1.390000 2.575000 2.155000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.573300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.090000 0.965000 10.430000 1.165000 ;
        RECT 10.170000 1.845000 10.430000 3.075000 ;
        RECT 10.225000 1.165000 10.430000 1.845000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.581700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.035000 1.820000 11.435000 3.075000 ;
        RECT 11.165000 0.255000 11.435000 1.095000 ;
        RECT 11.185000 1.095000 11.435000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.535000 1.920000 1.825000 1.965000 ;
        RECT 1.535000 1.965000 8.065000 2.105000 ;
        RECT 1.535000 2.105000 1.825000 2.150000 ;
        RECT 4.415000 1.920000 4.705000 1.965000 ;
        RECT 4.415000 2.105000 4.705000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.530000 1.580000 0.915000 2.180000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.100000  0.585000  0.430000 1.070000 ;
      RECT  0.100000  1.070000  1.035000 1.400000 ;
      RECT  0.100000  1.400000  0.360000 3.020000 ;
      RECT  0.530000  2.350000  0.860000 3.245000 ;
      RECT  0.600000  0.085000  0.810000 0.900000 ;
      RECT  0.980000  0.585000  1.375000 0.870000 ;
      RECT  0.980000  0.870000  2.255000 0.900000 ;
      RECT  1.030000  2.350000  1.350000 3.020000 ;
      RECT  1.110000  1.580000  1.395000 2.100000 ;
      RECT  1.110000  2.100000  1.350000 2.350000 ;
      RECT  1.205000  0.900000  2.255000 1.040000 ;
      RECT  1.205000  1.040000  1.395000 1.580000 ;
      RECT  1.520000  2.325000  3.345000 2.495000 ;
      RECT  1.520000  2.495000  1.730000 2.735000 ;
      RECT  1.545000  0.085000  1.875000 0.700000 ;
      RECT  1.595000  1.450000  1.860000 2.155000 ;
      RECT  1.970000  2.665000  2.320000 3.245000 ;
      RECT  2.045000  0.630000  4.755000 0.720000 ;
      RECT  2.045000  0.720000  6.450000 0.800000 ;
      RECT  2.045000  0.800000  2.255000 0.870000 ;
      RECT  2.485000  0.980000  2.925000 1.220000 ;
      RECT  2.540000  2.495000  3.345000 2.735000 ;
      RECT  2.755000  1.220000  2.925000 2.115000 ;
      RECT  2.755000  2.115000  3.150000 2.300000 ;
      RECT  2.755000  2.300000  3.345000 2.325000 ;
      RECT  3.095000  0.800000  3.265000 1.615000 ;
      RECT  3.095000  1.615000  3.500000 1.945000 ;
      RECT  3.435000  0.970000  4.215000 1.060000 ;
      RECT  3.435000  1.060000  5.600000 1.260000 ;
      RECT  3.435000  1.260000  3.860000 1.300000 ;
      RECT  3.515000  2.370000  5.095000 2.470000 ;
      RECT  3.515000  2.470000  3.965000 2.735000 ;
      RECT  3.680000  1.300000  3.860000 2.300000 ;
      RECT  3.680000  2.300000  5.095000 2.370000 ;
      RECT  4.040000  1.440000  5.240000 1.610000 ;
      RECT  4.040000  1.610000  4.295000 2.030000 ;
      RECT  4.340000  2.650000  4.670000 3.245000 ;
      RECT  4.475000  1.790000  4.900000 2.120000 ;
      RECT  4.540000  0.800000  6.450000 0.890000 ;
      RECT  4.850000  2.470000  5.095000 2.735000 ;
      RECT  5.070000  1.610000  5.240000 1.900000 ;
      RECT  5.070000  1.900000  6.145000 2.070000 ;
      RECT  5.225000  0.085000  5.555000 0.550000 ;
      RECT  5.350000  2.240000  5.680000 3.245000 ;
      RECT  5.410000  1.260000  5.600000 1.720000 ;
      RECT  5.770000  1.060000  6.100000 1.320000 ;
      RECT  5.930000  1.320000  6.100000 1.900000 ;
      RECT  5.930000  2.070000  6.145000 2.910000 ;
      RECT  6.270000  0.890000  6.450000 1.720000 ;
      RECT  6.500000  2.040000  6.820000 2.915000 ;
      RECT  6.620000  0.630000  6.820000 1.250000 ;
      RECT  6.620000  1.250000  8.430000 1.430000 ;
      RECT  6.620000  1.430000  6.820000 2.040000 ;
      RECT  7.200000  1.600000  8.790000 1.770000 ;
      RECT  7.200000  1.770000  7.530000 2.190000 ;
      RECT  7.325000  2.405000  7.995000 3.245000 ;
      RECT  7.495000  0.085000  7.685000 0.950000 ;
      RECT  7.740000  1.940000  8.070000 2.200000 ;
      RECT  7.875000  0.345000  9.130000 0.515000 ;
      RECT  7.875000  0.515000  8.045000 1.190000 ;
      RECT  7.875000  1.190000  8.430000 1.250000 ;
      RECT  8.165000  2.345000  8.420000 2.735000 ;
      RECT  8.225000  0.685000  8.790000 1.015000 ;
      RECT  8.250000  1.770000  8.790000 1.970000 ;
      RECT  8.250000  1.970000  8.420000 2.345000 ;
      RECT  8.590000  2.405000  8.825000 3.245000 ;
      RECT  8.610000  1.015000  8.790000 1.600000 ;
      RECT  8.960000  0.515000  9.130000 0.625000 ;
      RECT  8.960000  0.625000 10.995000 0.795000 ;
      RECT  8.960000  0.965000  9.290000 1.145000 ;
      RECT  8.960000  1.145000  9.165000 1.250000 ;
      RECT  8.995000  1.250000  9.165000 2.165000 ;
      RECT  8.995000  2.165000 10.000000 2.335000 ;
      RECT  8.995000  2.335000  9.325000 3.065000 ;
      RECT  9.345000  1.325000  9.640000 1.995000 ;
      RECT  9.460000  0.795000  9.640000 1.325000 ;
      RECT  9.505000  2.505000  9.835000 3.245000 ;
      RECT  9.600000  0.085000  9.930000 0.455000 ;
      RECT  9.830000  1.345000 10.055000 1.675000 ;
      RECT  9.830000  1.675000 10.000000 2.165000 ;
      RECT 10.600000  1.820000 10.865000 3.245000 ;
      RECT 10.665000  0.085000 10.995000 0.455000 ;
      RECT 10.825000  0.795000 10.995000 1.185000 ;
      RECT 10.825000  1.185000 11.015000 1.515000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  1.950000  1.765000 2.120000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  1.950000  4.645000 2.120000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
  END
END sky130_fd_sc_lp__dfrbp_1
END LIBRARY
