* File: sky130_fd_sc_lp__inv_0.pex.spice
* Created: Wed Sep  2 09:55:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_0%A 3 7 9 10 11 16 17
r18 16 19 88.6355 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=0.332 $Y=1.12
+ $X2=0.332 $Y2=1.625
r19 16 18 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.332 $Y=1.12
+ $X2=0.332 $Y2=0.955
r20 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r21 10 11 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.665
+ $X2=0.242 $Y2=2.035
r22 9 10 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.665
r23 9 17 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.12
r24 7 19 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=0.485 $Y=2.63
+ $X2=0.485 $Y2=1.625
r25 3 18 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.485 $Y=0.56
+ $X2=0.485 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__INV_0%VPWR 1 4 6 8 12 13
r13 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r14 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r15 10 16 4.4377 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.2
+ $Y2=3.33
r16 10 12 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.72
+ $Y2=3.33
r17 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.72 $Y2=3.33
r18 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 4 16 3.03982 $w=2.95e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.2 $Y2=3.33
r20 4 6 30.862 $w=2.93e-07 $l=7.9e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.252 $Y2=2.455
r21 1 6 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=2.31 $X2=0.27 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__INV_0%Y 1 2 7 8 9 10 11 12 20
r9 11 12 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=2.405
+ $X2=0.722 $Y2=2.775
r10 10 11 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=2.035
+ $X2=0.722 $Y2=2.405
r11 9 10 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=1.665
+ $X2=0.722 $Y2=2.035
r12 8 9 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=1.295
+ $X2=0.722 $Y2=1.665
r13 7 8 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=0.925
+ $X2=0.722 $Y2=1.295
r14 7 20 13.7915 $w=3.03e-07 $l=3.65e-07 $layer=LI1_cond $X=0.722 $Y=0.925
+ $X2=0.722 $Y2=0.56
r15 2 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=2.31 $X2=0.7 $Y2=2.455
r16 1 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.35 $X2=0.7 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__INV_0%VGND 1 4 6 8 12 13
r11 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r12 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r13 10 16 4.4377 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.2 $Y2=0
r14 10 12 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.72
+ $Y2=0
r15 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r16 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r17 4 16 3.03982 $w=2.95e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.252 $Y=0.085
+ $X2=0.2 $Y2=0
r18 4 6 18.5563 $w=2.93e-07 $l=4.75e-07 $layer=LI1_cond $X=0.252 $Y=0.085
+ $X2=0.252 $Y2=0.56
r19 1 6 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.35 $X2=0.27 $Y2=0.56
.ends

