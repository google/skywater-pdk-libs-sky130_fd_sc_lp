* File: sky130_fd_sc_lp__dlrtn_lp.pxi.spice
* Created: Wed Sep  2 09:47:10 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTN_LP%D N_D_c_157_n N_D_M1003_g N_D_c_158_n N_D_M1000_g
+ N_D_c_159_n N_D_c_160_n N_D_M1019_g N_D_c_161_n N_D_c_162_n D D N_D_c_163_n
+ N_D_c_164_n N_D_c_165_n PM_SKY130_FD_SC_LP__DLRTN_LP%D
x_PM_SKY130_FD_SC_LP__DLRTN_LP%GATE_N N_GATE_N_c_201_n N_GATE_N_M1012_g
+ N_GATE_N_M1004_g N_GATE_N_c_203_n N_GATE_N_M1005_g N_GATE_N_c_205_n GATE_N
+ GATE_N N_GATE_N_c_207_n PM_SKY130_FD_SC_LP__DLRTN_LP%GATE_N
x_PM_SKY130_FD_SC_LP__DLRTN_LP%A_264_415# N_A_264_415#_M1005_d
+ N_A_264_415#_M1012_d N_A_264_415#_c_254_n N_A_264_415#_M1015_g
+ N_A_264_415#_c_255_n N_A_264_415#_c_256_n N_A_264_415#_M1018_g
+ N_A_264_415#_c_258_n N_A_264_415#_M1010_g N_A_264_415#_M1020_g
+ N_A_264_415#_c_261_n N_A_264_415#_c_271_n N_A_264_415#_M1023_g
+ N_A_264_415#_c_262_n N_A_264_415#_c_274_n N_A_264_415#_c_263_n
+ N_A_264_415#_c_264_n N_A_264_415#_c_265_n N_A_264_415#_c_266_n
+ N_A_264_415#_c_267_n PM_SKY130_FD_SC_LP__DLRTN_LP%A_264_415#
x_PM_SKY130_FD_SC_LP__DLRTN_LP%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1000_s
+ N_A_27_47#_M1016_g N_A_27_47#_c_388_n N_A_27_47#_c_389_n N_A_27_47#_M1022_g
+ N_A_27_47#_c_404_n N_A_27_47#_c_398_n N_A_27_47#_c_399_n N_A_27_47#_c_391_n
+ N_A_27_47#_c_392_n N_A_27_47#_c_393_n N_A_27_47#_c_394_n N_A_27_47#_c_402_n
+ N_A_27_47#_c_395_n N_A_27_47#_c_413_n N_A_27_47#_c_396_n
+ PM_SKY130_FD_SC_LP__DLRTN_LP%A_27_47#
x_PM_SKY130_FD_SC_LP__DLRTN_LP%A_399_415# N_A_399_415#_M1018_s
+ N_A_399_415#_M1015_s N_A_399_415#_M1002_g N_A_399_415#_M1007_g
+ N_A_399_415#_c_481_n N_A_399_415#_c_482_n N_A_399_415#_c_483_n
+ N_A_399_415#_c_484_n N_A_399_415#_c_485_n N_A_399_415#_c_486_n
+ N_A_399_415#_c_487_n N_A_399_415#_c_488_n N_A_399_415#_c_489_n
+ N_A_399_415#_c_490_n N_A_399_415#_c_491_n N_A_399_415#_c_492_n
+ PM_SKY130_FD_SC_LP__DLRTN_LP%A_399_415#
x_PM_SKY130_FD_SC_LP__DLRTN_LP%A_949_335# N_A_949_335#_M1001_s
+ N_A_949_335#_M1021_d N_A_949_335#_M1009_g N_A_949_335#_M1013_g
+ N_A_949_335#_M1011_g N_A_949_335#_M1017_g N_A_949_335#_M1014_g
+ N_A_949_335#_c_598_n N_A_949_335#_c_614_n N_A_949_335#_c_599_n
+ N_A_949_335#_c_600_n N_A_949_335#_c_601_n N_A_949_335#_c_602_n
+ N_A_949_335#_c_615_n N_A_949_335#_c_632_p N_A_949_335#_c_603_n
+ N_A_949_335#_c_604_n N_A_949_335#_c_616_n N_A_949_335#_c_605_n
+ N_A_949_335#_c_606_n N_A_949_335#_c_607_n N_A_949_335#_c_608_n
+ N_A_949_335#_c_609_n N_A_949_335#_c_610_n
+ PM_SKY130_FD_SC_LP__DLRTN_LP%A_949_335#
x_PM_SKY130_FD_SC_LP__DLRTN_LP%A_744_415# N_A_744_415#_M1020_d
+ N_A_744_415#_M1002_d N_A_744_415#_M1021_g N_A_744_415#_c_729_n
+ N_A_744_415#_c_730_n N_A_744_415#_M1001_g N_A_744_415#_c_731_n
+ N_A_744_415#_c_737_n N_A_744_415#_c_744_n N_A_744_415#_c_745_n
+ N_A_744_415#_c_738_n N_A_744_415#_c_732_n N_A_744_415#_c_747_n
+ N_A_744_415#_c_733_n N_A_744_415#_c_734_n N_A_744_415#_c_735_n
+ PM_SKY130_FD_SC_LP__DLRTN_LP%A_744_415#
x_PM_SKY130_FD_SC_LP__DLRTN_LP%RESET_B N_RESET_B_M1008_g N_RESET_B_M1006_g
+ N_RESET_B_c_829_n N_RESET_B_c_834_n RESET_B N_RESET_B_c_830_n
+ N_RESET_B_c_831_n PM_SKY130_FD_SC_LP__DLRTN_LP%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTN_LP%VPWR N_VPWR_M1000_d N_VPWR_M1015_d N_VPWR_M1009_d
+ N_VPWR_M1008_d N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n
+ N_VPWR_c_883_n N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n
+ N_VPWR_c_888_n VPWR N_VPWR_c_889_n N_VPWR_c_890_n N_VPWR_c_878_n
+ N_VPWR_c_892_n PM_SKY130_FD_SC_LP__DLRTN_LP%VPWR
x_PM_SKY130_FD_SC_LP__DLRTN_LP%Q N_Q_M1014_d N_Q_M1017_d Q Q Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DLRTN_LP%Q
x_PM_SKY130_FD_SC_LP__DLRTN_LP%VGND N_VGND_M1019_d N_VGND_M1010_d N_VGND_M1013_d
+ N_VGND_M1006_d N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n
+ N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n VGND N_VGND_c_983_n
+ N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n
+ N_VGND_c_989_n PM_SKY130_FD_SC_LP__DLRTN_LP%VGND
cc_1 VNB N_D_c_157_n 0.0180432f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_D_c_158_n 0.0223277f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.595
cc_3 VNB N_D_c_159_n 0.0194214f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_4 VNB N_D_c_160_n 0.0135378f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_5 VNB N_D_c_161_n 0.00611761f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_6 VNB N_D_c_162_n 0.00449551f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.78
cc_7 VNB N_D_c_163_n 0.0163556f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.275
cc_8 VNB N_D_c_164_n 0.00669862f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.275
cc_9 VNB N_D_c_165_n 0.0108193f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.11
cc_10 VNB N_GATE_N_c_201_n 0.00208313f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_11 VNB N_GATE_N_M1004_g 0.0392434f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.595
cc_12 VNB N_GATE_N_c_203_n 0.0260776f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.575
cc_13 VNB N_GATE_N_M1005_g 0.0383543f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.805
cc_14 VNB N_GATE_N_c_205_n 0.0130941f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_15 VNB GATE_N 0.00251617f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.78
cc_16 VNB N_GATE_N_c_207_n 0.0270751f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.275
cc_17 VNB N_A_264_415#_c_254_n 0.0175077f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.595
cc_18 VNB N_A_264_415#_c_255_n 0.0528264f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.805
cc_19 VNB N_A_264_415#_c_256_n 0.0156858f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_20 VNB N_A_264_415#_M1018_g 0.0210279f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_21 VNB N_A_264_415#_c_258_n 0.0186614f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_A_264_415#_M1010_g 0.0160228f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.275
cc_23 VNB N_A_264_415#_M1020_g 0.0293444f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.275
cc_24 VNB N_A_264_415#_c_261_n 0.02366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_264_415#_c_262_n 0.0085456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_264_415#_c_263_n 0.0145844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_264_415#_c_264_n 0.0135821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_264_415#_c_265_n 0.0282399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_264_415#_c_266_n 0.00262036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_264_415#_c_267_n 0.0111433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_388_n 0.0242565f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.805
cc_32 VNB N_A_27_47#_c_389_n 0.00798099f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_33 VNB N_A_27_47#_M1022_g 0.0370024f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_34 VNB N_A_27_47#_c_391_n 3.20109e-19 $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.275
cc_35 VNB N_A_27_47#_c_392_n 0.00297314f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.295
cc_36 VNB N_A_27_47#_c_393_n 0.00967168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_c_394_n 0.021289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_395_n 0.0466843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_c_396_n 0.0216297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_399_415#_c_481_n 0.0176316f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_41 VNB N_A_399_415#_c_482_n 0.0158429f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.78
cc_42 VNB N_A_399_415#_c_483_n 0.00514715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_399_415#_c_484_n 0.0256696f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.275
cc_44 VNB N_A_399_415#_c_485_n 0.0153274f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.275
cc_45 VNB N_A_399_415#_c_486_n 0.00834f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.11
cc_46 VNB N_A_399_415#_c_487_n 0.00374908f $X=-0.19 $Y=-0.245 $X2=0.647
+ $Y2=1.665
cc_47 VNB N_A_399_415#_c_488_n 0.055775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_399_415#_c_489_n 0.00274086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_399_415#_c_490_n 0.003035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_399_415#_c_491_n 0.011644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_399_415#_c_492_n 0.0040006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_949_335#_M1013_g 0.0259927f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.805
cc_53 VNB N_A_949_335#_M1011_g 0.0175998f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_54 VNB N_A_949_335#_M1017_g 0.00831986f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.275
cc_55 VNB N_A_949_335#_M1014_g 0.021956f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.275
cc_56 VNB N_A_949_335#_c_598_n 0.0312778f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.295
cc_57 VNB N_A_949_335#_c_599_n 0.00907443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_949_335#_c_600_n 0.0274633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_949_335#_c_601_n 0.0149589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_949_335#_c_602_n 0.00831903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_949_335#_c_603_n 0.0145056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_949_335#_c_604_n 0.0148142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_949_335#_c_605_n 0.00125664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_949_335#_c_606_n 0.00279621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_949_335#_c_607_n 7.90679e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_949_335#_c_608_n 0.0442661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_949_335#_c_609_n 0.0248887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_949_335#_c_610_n 0.00111775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_744_415#_c_729_n 0.0297411f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_70 VNB N_A_744_415#_c_730_n 0.0195698f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.805
cc_71 VNB N_A_744_415#_c_731_n 0.0177771f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.78
cc_72 VNB N_A_744_415#_c_732_n 0.00477688f $X=-0.19 $Y=-0.245 $X2=0.647
+ $Y2=1.665
cc_73 VNB N_A_744_415#_c_733_n 0.00266761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_744_415#_c_734_n 0.00232024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_744_415#_c_735_n 0.0313696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_RESET_B_M1006_g 0.0347417f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.595
cc_77 VNB N_RESET_B_c_829_n 0.0162651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_RESET_B_c_830_n 0.0138487f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_79 VNB N_RESET_B_c_831_n 0.00443907f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_80 VNB N_VPWR_c_878_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB Q 0.0667137f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.595
cc_82 VNB N_VGND_c_976_n 0.00642294f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_83 VNB N_VGND_c_977_n 0.0470907f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_84 VNB N_VGND_c_978_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_979_n 0.0110755f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.275
cc_86 VNB N_VGND_c_980_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.295
cc_87 VNB N_VGND_c_981_n 0.043414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_982_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_983_n 0.0268233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_984_n 0.0286512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_985_n 0.0271986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_986_n 0.388248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_987_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_988_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_989_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VPB N_D_M1000_g 0.04017f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.575
cc_97 VPB N_D_c_162_n 0.0127696f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.78
cc_98 VPB N_D_c_164_n 0.00348152f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.275
cc_99 VPB N_GATE_N_c_201_n 0.0116021f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.73
cc_100 VPB N_GATE_N_M1012_g 0.0373453f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_101 VPB GATE_N 0.00201838f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.78
cc_102 VPB N_A_264_415#_c_254_n 0.0179089f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.595
cc_103 VPB N_A_264_415#_M1015_g 0.041369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_264_415#_c_261_n 0.00104039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_264_415#_c_271_n 0.0280946f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=1.665
cc_106 VPB N_A_264_415#_M1023_g 0.0339876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_264_415#_c_262_n 0.00344964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_264_415#_c_274_n 0.0152979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_264_415#_c_263_n 0.00249886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_264_415#_c_267_n 0.0274205f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_M1016_g 0.0269222f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.575
cc_112 VPB N_A_27_47#_c_398_n 0.013971f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.275
cc_113 VPB N_A_27_47#_c_399_n 0.00185706f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.11
cc_114 VPB N_A_27_47#_c_392_n 0.00989857f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=1.295
cc_115 VPB N_A_27_47#_c_393_n 0.0179895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_402_n 0.0524834f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_395_n 0.0195691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_399_415#_M1002_g 0.0279676f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.575
cc_119 VPB N_A_399_415#_c_482_n 0.00557345f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.78
cc_120 VPB N_A_399_415#_c_486_n 0.00670756f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.11
cc_121 VPB N_A_399_415#_c_490_n 0.0029091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_399_415#_c_491_n 0.0202319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_949_335#_M1009_g 0.0351718f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.575
cc_124 VPB N_A_949_335#_M1017_g 0.0465107f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.275
cc_125 VPB N_A_949_335#_c_598_n 0.00112658f $X=-0.19 $Y=1.655 $X2=0.647
+ $Y2=1.295
cc_126 VPB N_A_949_335#_c_614_n 0.0213554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_949_335#_c_615_n 0.00247894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_949_335#_c_616_n 0.00665803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_949_335#_c_607_n 0.00318489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_744_415#_M1021_g 0.040426f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.575
cc_131 VPB N_A_744_415#_c_737_n 0.00279184f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_132 VPB N_A_744_415#_c_738_n 0.00482835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_744_415#_c_733_n 0.00662121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_744_415#_c_734_n 2.06056e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_744_415#_c_735_n 0.0210176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_RESET_B_M1008_g 0.0292411f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_137 VPB N_RESET_B_c_829_n 0.00321417f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_RESET_B_c_834_n 0.0122621f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.805
cc_139 VPB N_RESET_B_c_831_n 0.00413963f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.805
cc_140 VPB N_VPWR_c_879_n 0.00100404f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_141 VPB N_VPWR_c_880_n 0.00292294f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_142 VPB N_VPWR_c_881_n 0.0102257f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.275
cc_143 VPB N_VPWR_c_882_n 0.0034231f $X=-0.19 $Y=1.655 $X2=0.647 $Y2=1.295
cc_144 VPB N_VPWR_c_883_n 0.0205471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_884_n 0.00460685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_885_n 0.0434575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_886_n 0.00372128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_887_n 0.065049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_888_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_889_n 0.0243168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_890_n 0.027616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_878_n 0.11886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_892_n 0.00526006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB Q 0.0229543f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.595
cc_155 VPB Q 0.0201773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB Q 0.037144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 N_D_c_162_n N_GATE_N_c_201_n 0.011958f $X=0.605 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_158 N_D_M1000_g N_GATE_N_M1012_g 0.0522092f $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_159 N_D_c_160_n N_GATE_N_M1004_g 0.0185179f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_160 N_D_c_163_n N_GATE_N_M1004_g 2.30929e-19 $X=0.625 $Y=1.275 $X2=0 $Y2=0
cc_161 N_D_c_165_n N_GATE_N_M1004_g 0.00118442f $X=0.605 $Y=1.11 $X2=0 $Y2=0
cc_162 N_D_c_163_n N_GATE_N_c_205_n 0.011958f $X=0.625 $Y=1.275 $X2=0 $Y2=0
cc_163 N_D_c_164_n N_GATE_N_c_205_n 0.00415243f $X=0.625 $Y=1.275 $X2=0 $Y2=0
cc_164 N_D_c_163_n GATE_N 7.68828e-19 $X=0.625 $Y=1.275 $X2=0 $Y2=0
cc_165 N_D_c_164_n GATE_N 0.0475486f $X=0.625 $Y=1.275 $X2=0 $Y2=0
cc_166 N_D_c_158_n N_GATE_N_c_207_n 0.011958f $X=0.605 $Y=1.595 $X2=0 $Y2=0
cc_167 N_D_M1000_g N_A_264_415#_c_274_n 0.00110366f $X=0.665 $Y=2.575 $X2=0
+ $Y2=0
cc_168 N_D_M1000_g N_A_27_47#_c_404_n 0.0210641f $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_169 N_D_c_157_n N_A_27_47#_c_394_n 0.00850964f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_170 N_D_c_160_n N_A_27_47#_c_394_n 0.00111582f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_171 N_D_M1000_g N_A_27_47#_c_402_n 0.0187074f $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_172 N_D_c_162_n N_A_27_47#_c_402_n 0.002357f $X=0.605 $Y=1.78 $X2=0 $Y2=0
cc_173 N_D_c_164_n N_A_27_47#_c_402_n 0.00627901f $X=0.625 $Y=1.275 $X2=0 $Y2=0
cc_174 N_D_c_157_n N_A_27_47#_c_395_n 0.0317162f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_175 N_D_M1000_g N_A_27_47#_c_395_n 0.00740404f $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_176 N_D_c_164_n N_A_27_47#_c_395_n 0.0486307f $X=0.625 $Y=1.275 $X2=0 $Y2=0
cc_177 N_D_M1000_g N_A_27_47#_c_413_n 6.186e-19 $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_178 N_D_M1000_g N_VPWR_c_879_n 0.00980888f $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_179 N_D_M1000_g N_VPWR_c_883_n 0.00608873f $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_180 N_D_M1000_g N_VPWR_c_878_n 0.00792977f $X=0.665 $Y=2.575 $X2=0 $Y2=0
cc_181 N_D_c_157_n N_VGND_c_976_n 0.00239794f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_182 N_D_c_160_n N_VGND_c_976_n 0.01353f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_183 N_D_c_157_n N_VGND_c_983_n 0.00549284f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_184 N_D_c_159_n N_VGND_c_983_n 4.87571e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_185 N_D_c_160_n N_VGND_c_983_n 0.00486043f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_186 N_D_c_157_n N_VGND_c_986_n 0.010905f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_187 N_D_c_159_n N_VGND_c_986_n 6.51792e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_188 N_D_c_160_n N_VGND_c_986_n 0.00814425f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_189 N_GATE_N_M1005_g N_A_264_415#_c_255_n 0.00305873f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_190 N_GATE_N_c_201_n N_A_264_415#_c_274_n 2.58585e-19 $X=1.195 $Y=1.79 $X2=0
+ $Y2=0
cc_191 N_GATE_N_M1012_g N_A_264_415#_c_274_n 0.00676661f $X=1.195 $Y=2.575 $X2=0
+ $Y2=0
cc_192 GATE_N N_A_264_415#_c_274_n 0.00367208f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_193 N_GATE_N_M1012_g N_A_264_415#_c_263_n 0.00581063f $X=1.195 $Y=2.575 $X2=0
+ $Y2=0
cc_194 N_GATE_N_M1004_g N_A_264_415#_c_263_n 0.0102409f $X=1.285 $Y=0.445 $X2=0
+ $Y2=0
cc_195 N_GATE_N_c_203_n N_A_264_415#_c_263_n 0.00910596f $X=1.6 $Y=1.195 $X2=0
+ $Y2=0
cc_196 N_GATE_N_M1005_g N_A_264_415#_c_263_n 0.0201758f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_197 GATE_N N_A_264_415#_c_263_n 0.0434507f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_198 N_GATE_N_c_207_n N_A_264_415#_c_263_n 0.0076821f $X=1.195 $Y=1.285 $X2=0
+ $Y2=0
cc_199 N_GATE_N_M1005_g N_A_264_415#_c_266_n 0.00520773f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_GATE_N_M1012_g N_A_264_415#_c_267_n 0.00689064f $X=1.195 $Y=2.575 $X2=0
+ $Y2=0
cc_201 N_GATE_N_c_203_n N_A_264_415#_c_267_n 0.00704159f $X=1.6 $Y=1.195 $X2=0
+ $Y2=0
cc_202 GATE_N N_A_264_415#_c_267_n 7.96549e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_203 N_GATE_N_c_207_n N_A_264_415#_c_267_n 0.0130346f $X=1.195 $Y=1.285 $X2=0
+ $Y2=0
cc_204 N_GATE_N_M1012_g N_A_27_47#_c_404_n 0.0193917f $X=1.195 $Y=2.575 $X2=0
+ $Y2=0
cc_205 N_GATE_N_M1012_g N_A_27_47#_c_398_n 9.86509e-19 $X=1.195 $Y=2.575 $X2=0
+ $Y2=0
cc_206 N_GATE_N_M1012_g N_A_27_47#_c_402_n 0.00249872f $X=1.195 $Y=2.575 $X2=0
+ $Y2=0
cc_207 N_GATE_N_M1012_g N_A_27_47#_c_413_n 0.0124846f $X=1.195 $Y=2.575 $X2=0
+ $Y2=0
cc_208 N_GATE_N_M1005_g N_A_399_415#_c_482_n 0.00169243f $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_GATE_N_M1005_g N_A_399_415#_c_483_n 7.00968e-19 $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_210 N_GATE_N_M1005_g N_A_399_415#_c_485_n 9.92157e-19 $X=1.675 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_GATE_N_M1012_g N_VPWR_c_879_n 0.0157608f $X=1.195 $Y=2.575 $X2=0 $Y2=0
cc_212 N_GATE_N_M1012_g N_VPWR_c_885_n 0.00612037f $X=1.195 $Y=2.575 $X2=0 $Y2=0
cc_213 N_GATE_N_M1012_g N_VPWR_c_878_n 0.00818443f $X=1.195 $Y=2.575 $X2=0 $Y2=0
cc_214 N_GATE_N_M1004_g N_VGND_c_976_n 0.0122138f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_215 N_GATE_N_M1005_g N_VGND_c_976_n 0.00177822f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_216 N_GATE_N_c_205_n N_VGND_c_976_n 0.00122441f $X=1.195 $Y=1.195 $X2=0 $Y2=0
cc_217 GATE_N N_VGND_c_976_n 0.00866099f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_218 N_GATE_N_M1004_g N_VGND_c_977_n 0.00486043f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_219 N_GATE_N_M1005_g N_VGND_c_977_n 0.00366111f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_220 N_GATE_N_M1004_g N_VGND_c_986_n 0.00823808f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_221 N_GATE_N_M1005_g N_VGND_c_986_n 0.00654681f $X=1.675 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_264_415#_M1015_g N_A_27_47#_M1016_g 0.0213982f $X=2.405 $Y=2.575
+ $X2=0 $Y2=0
cc_223 N_A_264_415#_c_264_n N_A_27_47#_c_388_n 0.018275f $X=3.965 $Y=1.18 $X2=0
+ $Y2=0
cc_224 N_A_264_415#_c_265_n N_A_27_47#_c_388_n 0.0344181f $X=3.965 $Y=1.18 $X2=0
+ $Y2=0
cc_225 N_A_264_415#_c_255_n N_A_27_47#_c_389_n 0.0060033f $X=2.455 $Y=1.345
+ $X2=0 $Y2=0
cc_226 N_A_264_415#_c_258_n N_A_27_47#_c_389_n 0.00276269f $X=2.98 $Y=0.88 $X2=0
+ $Y2=0
cc_227 N_A_264_415#_c_264_n N_A_27_47#_c_389_n 0.00872219f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_228 N_A_264_415#_c_255_n N_A_27_47#_M1022_g 0.00356628f $X=2.455 $Y=1.345
+ $X2=0 $Y2=0
cc_229 N_A_264_415#_M1010_g N_A_27_47#_M1022_g 0.0242879f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_230 N_A_264_415#_M1020_g N_A_27_47#_M1022_g 0.0344181f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_231 N_A_264_415#_c_264_n N_A_27_47#_M1022_g 0.0100442f $X=3.965 $Y=1.18 $X2=0
+ $Y2=0
cc_232 N_A_264_415#_M1012_d N_A_27_47#_c_398_n 0.00608748f $X=1.32 $Y=2.075
+ $X2=0 $Y2=0
cc_233 N_A_264_415#_M1015_g N_A_27_47#_c_398_n 0.0193692f $X=2.405 $Y=2.575
+ $X2=0 $Y2=0
cc_234 N_A_264_415#_c_274_n N_A_27_47#_c_398_n 0.0209736f $X=1.57 $Y=2.185 $X2=0
+ $Y2=0
cc_235 N_A_264_415#_M1015_g N_A_27_47#_c_399_n 0.0263229f $X=2.405 $Y=2.575
+ $X2=0 $Y2=0
cc_236 N_A_264_415#_M1015_g N_A_27_47#_c_391_n 0.00620561f $X=2.405 $Y=2.575
+ $X2=0 $Y2=0
cc_237 N_A_264_415#_c_255_n N_A_27_47#_c_391_n 0.00100947f $X=2.455 $Y=1.345
+ $X2=0 $Y2=0
cc_238 N_A_264_415#_c_262_n N_A_27_47#_c_391_n 0.00953098f $X=2.405 $Y=1.66
+ $X2=0 $Y2=0
cc_239 N_A_264_415#_c_264_n N_A_27_47#_c_391_n 0.00837986f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_240 N_A_264_415#_c_255_n N_A_27_47#_c_392_n 0.00479981f $X=2.455 $Y=1.345
+ $X2=0 $Y2=0
cc_241 N_A_264_415#_c_264_n N_A_27_47#_c_392_n 0.0399732f $X=3.965 $Y=1.18 $X2=0
+ $Y2=0
cc_242 N_A_264_415#_c_258_n N_A_27_47#_c_393_n 0.00226448f $X=2.98 $Y=0.88 $X2=0
+ $Y2=0
cc_243 N_A_264_415#_c_262_n N_A_27_47#_c_393_n 0.0103254f $X=2.405 $Y=1.66 $X2=0
+ $Y2=0
cc_244 N_A_264_415#_c_264_n N_A_27_47#_c_393_n 0.0019391f $X=3.965 $Y=1.18 $X2=0
+ $Y2=0
cc_245 N_A_264_415#_M1012_d N_A_27_47#_c_413_n 0.00875823f $X=1.32 $Y=2.075
+ $X2=0 $Y2=0
cc_246 N_A_264_415#_c_274_n N_A_27_47#_c_413_n 0.00683325f $X=1.57 $Y=2.185
+ $X2=0 $Y2=0
cc_247 N_A_264_415#_c_256_n N_A_27_47#_c_396_n 0.00651864f $X=2.455 $Y=1.585
+ $X2=0 $Y2=0
cc_248 N_A_264_415#_M1023_g N_A_399_415#_M1002_g 0.0152634f $X=4.38 $Y=2.575
+ $X2=0 $Y2=0
cc_249 N_A_264_415#_M1020_g N_A_399_415#_c_481_n 0.0222629f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_250 N_A_264_415#_c_254_n N_A_399_415#_c_482_n 0.0145746f $X=2.28 $Y=1.66
+ $X2=0 $Y2=0
cc_251 N_A_264_415#_M1015_g N_A_399_415#_c_482_n 0.00596513f $X=2.405 $Y=2.575
+ $X2=0 $Y2=0
cc_252 N_A_264_415#_c_255_n N_A_399_415#_c_482_n 0.0183918f $X=2.455 $Y=1.345
+ $X2=0 $Y2=0
cc_253 N_A_264_415#_c_274_n N_A_399_415#_c_482_n 0.0204881f $X=1.57 $Y=2.185
+ $X2=0 $Y2=0
cc_254 N_A_264_415#_c_263_n N_A_399_415#_c_482_n 0.0903607f $X=1.735 $Y=1.75
+ $X2=0 $Y2=0
cc_255 N_A_264_415#_c_264_n N_A_399_415#_c_482_n 0.0219418f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_256 N_A_264_415#_c_267_n N_A_399_415#_c_482_n 0.00139703f $X=1.735 $Y=1.66
+ $X2=0 $Y2=0
cc_257 N_A_264_415#_M1018_g N_A_399_415#_c_483_n 0.00729198f $X=2.695 $Y=0.445
+ $X2=0 $Y2=0
cc_258 N_A_264_415#_M1010_g N_A_399_415#_c_483_n 0.00150162f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_259 N_A_264_415#_c_263_n N_A_399_415#_c_483_n 0.00743872f $X=1.735 $Y=1.75
+ $X2=0 $Y2=0
cc_260 N_A_264_415#_c_266_n N_A_399_415#_c_483_n 0.0120321f $X=1.89 $Y=0.39
+ $X2=0 $Y2=0
cc_261 N_A_264_415#_c_255_n N_A_399_415#_c_484_n 0.00208665f $X=2.455 $Y=1.345
+ $X2=0 $Y2=0
cc_262 N_A_264_415#_M1018_g N_A_399_415#_c_484_n 0.00581098f $X=2.695 $Y=0.445
+ $X2=0 $Y2=0
cc_263 N_A_264_415#_c_258_n N_A_399_415#_c_484_n 0.00488849f $X=2.98 $Y=0.88
+ $X2=0 $Y2=0
cc_264 N_A_264_415#_M1010_g N_A_399_415#_c_484_n 0.0081165f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_265 N_A_264_415#_M1020_g N_A_399_415#_c_484_n 0.0122822f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_266 N_A_264_415#_c_265_n N_A_399_415#_c_484_n 0.00459442f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_267 N_A_264_415#_c_255_n N_A_399_415#_c_485_n 0.00791294f $X=2.455 $Y=1.345
+ $X2=0 $Y2=0
cc_268 N_A_264_415#_M1018_g N_A_399_415#_c_485_n 0.00364314f $X=2.695 $Y=0.445
+ $X2=0 $Y2=0
cc_269 N_A_264_415#_c_263_n N_A_399_415#_c_485_n 0.01419f $X=1.735 $Y=1.75 $X2=0
+ $Y2=0
cc_270 N_A_264_415#_c_264_n N_A_399_415#_c_485_n 0.122154f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_271 N_A_264_415#_c_261_n N_A_399_415#_c_486_n 0.00633293f $X=4.055 $Y=1.675
+ $X2=0 $Y2=0
cc_272 N_A_264_415#_c_271_n N_A_399_415#_c_486_n 0.0174302f $X=4.38 $Y=1.825
+ $X2=0 $Y2=0
cc_273 N_A_264_415#_c_264_n N_A_399_415#_c_486_n 0.0204544f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_274 N_A_264_415#_c_265_n N_A_399_415#_c_486_n 0.00439769f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_275 N_A_264_415#_M1020_g N_A_399_415#_c_487_n 0.00352815f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_276 N_A_264_415#_c_264_n N_A_399_415#_c_487_n 0.0263463f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_277 N_A_264_415#_c_265_n N_A_399_415#_c_487_n 0.00109506f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_278 N_A_264_415#_c_271_n N_A_399_415#_c_488_n 0.00918315f $X=4.38 $Y=1.825
+ $X2=0 $Y2=0
cc_279 N_A_264_415#_c_264_n N_A_399_415#_c_488_n 3.86936e-19 $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_280 N_A_264_415#_c_265_n N_A_399_415#_c_488_n 0.0267159f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_281 N_A_264_415#_c_261_n N_A_399_415#_c_489_n 0.00354908f $X=4.055 $Y=1.675
+ $X2=0 $Y2=0
cc_282 N_A_264_415#_c_271_n N_A_399_415#_c_490_n 5.29207e-19 $X=4.38 $Y=1.825
+ $X2=0 $Y2=0
cc_283 N_A_264_415#_M1023_g N_A_399_415#_c_490_n 5.17698e-19 $X=4.38 $Y=2.575
+ $X2=0 $Y2=0
cc_284 N_A_264_415#_c_264_n N_A_399_415#_c_490_n 0.0196409f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_285 N_A_264_415#_c_261_n N_A_399_415#_c_491_n 0.0158864f $X=4.055 $Y=1.675
+ $X2=0 $Y2=0
cc_286 N_A_264_415#_M1023_g N_A_399_415#_c_491_n 0.00250189f $X=4.38 $Y=2.575
+ $X2=0 $Y2=0
cc_287 N_A_264_415#_c_264_n N_A_399_415#_c_491_n 0.00159907f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_288 N_A_264_415#_c_265_n N_A_399_415#_c_492_n 0.00354908f $X=3.965 $Y=1.18
+ $X2=0 $Y2=0
cc_289 N_A_264_415#_M1023_g N_A_949_335#_M1009_g 0.0433935f $X=4.38 $Y=2.575
+ $X2=0 $Y2=0
cc_290 N_A_264_415#_c_271_n N_A_949_335#_c_614_n 0.0433935f $X=4.38 $Y=1.825
+ $X2=0 $Y2=0
cc_291 N_A_264_415#_c_271_n N_A_744_415#_c_737_n 0.00663538f $X=4.38 $Y=1.825
+ $X2=0 $Y2=0
cc_292 N_A_264_415#_M1023_g N_A_744_415#_c_737_n 0.00116699f $X=4.38 $Y=2.575
+ $X2=0 $Y2=0
cc_293 N_A_264_415#_M1023_g N_A_744_415#_c_744_n 0.0166867f $X=4.38 $Y=2.575
+ $X2=0 $Y2=0
cc_294 N_A_264_415#_M1020_g N_A_744_415#_c_745_n 0.00300383f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_295 N_A_264_415#_M1023_g N_A_744_415#_c_738_n 0.0192958f $X=4.38 $Y=2.575
+ $X2=0 $Y2=0
cc_296 N_A_264_415#_c_271_n N_A_744_415#_c_747_n 0.00174512f $X=4.38 $Y=1.825
+ $X2=0 $Y2=0
cc_297 N_A_264_415#_c_261_n N_A_744_415#_c_734_n 7.16315e-19 $X=4.055 $Y=1.675
+ $X2=0 $Y2=0
cc_298 N_A_264_415#_c_271_n N_A_744_415#_c_734_n 2.86866e-19 $X=4.38 $Y=1.825
+ $X2=0 $Y2=0
cc_299 N_A_264_415#_M1015_g N_VPWR_c_880_n 0.0102998f $X=2.405 $Y=2.575 $X2=0
+ $Y2=0
cc_300 N_A_264_415#_M1015_g N_VPWR_c_885_n 0.00645804f $X=2.405 $Y=2.575 $X2=0
+ $Y2=0
cc_301 N_A_264_415#_M1023_g N_VPWR_c_887_n 0.00906878f $X=4.38 $Y=2.575 $X2=0
+ $Y2=0
cc_302 N_A_264_415#_M1015_g N_VPWR_c_878_n 0.00974819f $X=2.405 $Y=2.575 $X2=0
+ $Y2=0
cc_303 N_A_264_415#_M1023_g N_VPWR_c_878_n 0.0164887f $X=4.38 $Y=2.575 $X2=0
+ $Y2=0
cc_304 N_A_264_415#_c_263_n N_VGND_c_976_n 0.0046278f $X=1.735 $Y=1.75 $X2=0
+ $Y2=0
cc_305 N_A_264_415#_M1018_g N_VGND_c_977_n 0.00418312f $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_306 N_A_264_415#_M1010_g N_VGND_c_977_n 0.0035715f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_307 N_A_264_415#_c_266_n N_VGND_c_977_n 0.022491f $X=1.89 $Y=0.39 $X2=0 $Y2=0
cc_308 N_A_264_415#_M1018_g N_VGND_c_978_n 0.00188079f $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_309 N_A_264_415#_M1010_g N_VGND_c_978_n 0.00914585f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_310 N_A_264_415#_M1020_g N_VGND_c_978_n 0.00195503f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_311 N_A_264_415#_M1020_g N_VGND_c_981_n 0.00429465f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_312 N_A_264_415#_M1005_d N_VGND_c_986_n 0.0023412f $X=1.75 $Y=0.235 $X2=0
+ $Y2=0
cc_313 N_A_264_415#_M1018_g N_VGND_c_986_n 0.0071786f $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_314 N_A_264_415#_M1010_g N_VGND_c_986_n 0.00404234f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_315 N_A_264_415#_M1020_g N_VGND_c_986_n 0.00630445f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_316 N_A_264_415#_c_266_n N_VGND_c_986_n 0.0170706f $X=1.89 $Y=0.39 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_398_n N_A_399_415#_M1015_s 0.00842335f $X=2.405 $Y=2.75
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_M1016_g N_A_399_415#_M1002_g 0.0767523f $X=3.105 $Y=2.575
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_398_n N_A_399_415#_c_482_n 0.0126095f $X=2.405 $Y=2.75 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_399_n N_A_399_415#_c_482_n 0.0241651f $X=2.49 $Y=2.665 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_391_n N_A_399_415#_c_482_n 0.0246417f $X=2.575 $Y=1.75 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_389_n N_A_399_415#_c_484_n 0.00132122f $X=3.23 $Y=1.27 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1022_g N_A_399_415#_c_484_n 0.0114565f $X=3.485 $Y=0.445
+ $X2=0 $Y2=0
cc_324 N_A_27_47#_c_388_n N_A_399_415#_c_490_n 5.09316e-19 $X=3.41 $Y=1.27 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_392_n N_A_399_415#_c_490_n 0.02209f $X=3.065 $Y=1.75 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_393_n N_A_399_415#_c_490_n 4.14293e-19 $X=3.065 $Y=1.75
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_388_n N_A_399_415#_c_491_n 0.00682692f $X=3.41 $Y=1.27 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_392_n N_A_399_415#_c_491_n 0.00114003f $X=3.065 $Y=1.75
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_393_n N_A_399_415#_c_491_n 0.0207808f $X=3.065 $Y=1.75 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_404_n N_VPWR_M1000_d 0.00807879f $X=1.275 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_331 N_A_27_47#_c_404_n N_VPWR_c_879_n 0.0153414f $X=1.275 $Y=2.58 $X2=0 $Y2=0
cc_332 N_A_27_47#_c_402_n N_VPWR_c_879_n 0.014861f $X=0.4 $Y=2.22 $X2=0 $Y2=0
cc_333 N_A_27_47#_M1016_g N_VPWR_c_880_n 0.0275616f $X=3.105 $Y=2.575 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_392_n N_VPWR_c_880_n 0.0176322f $X=3.065 $Y=1.75 $X2=0 $Y2=0
cc_335 N_A_27_47#_c_393_n N_VPWR_c_880_n 0.00167493f $X=3.065 $Y=1.75 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_404_n N_VPWR_c_883_n 0.00304017f $X=1.275 $Y=2.58 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_402_n N_VPWR_c_883_n 0.0281861f $X=0.4 $Y=2.22 $X2=0 $Y2=0
cc_338 N_A_27_47#_c_404_n N_VPWR_c_885_n 0.00273525f $X=1.275 $Y=2.58 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_398_n N_VPWR_c_885_n 0.02698f $X=2.405 $Y=2.75 $X2=0 $Y2=0
cc_340 N_A_27_47#_c_413_n N_VPWR_c_885_n 0.00361883f $X=1.36 $Y=2.58 $X2=0 $Y2=0
cc_341 N_A_27_47#_M1016_g N_VPWR_c_887_n 0.00845957f $X=3.105 $Y=2.575 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_M1016_g N_VPWR_c_878_n 0.0143819f $X=3.105 $Y=2.575 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_404_n N_VPWR_c_878_n 0.010179f $X=1.275 $Y=2.58 $X2=0 $Y2=0
cc_344 N_A_27_47#_c_398_n N_VPWR_c_878_n 0.0349914f $X=2.405 $Y=2.75 $X2=0 $Y2=0
cc_345 N_A_27_47#_c_402_n N_VPWR_c_878_n 0.0174072f $X=0.4 $Y=2.22 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_413_n N_VPWR_c_878_n 0.00526615f $X=1.36 $Y=2.58 $X2=0 $Y2=0
cc_347 N_A_27_47#_c_394_n N_VGND_c_976_n 0.0137333f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_348 N_A_27_47#_M1022_g N_VGND_c_978_n 0.0096431f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_M1022_g N_VGND_c_981_n 0.0035715f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_394_n N_VGND_c_983_n 0.019876f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_351 N_A_27_47#_M1003_s N_VGND_c_986_n 0.00232985f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_M1022_g N_VGND_c_986_n 0.00417192f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_394_n N_VGND_c_986_n 0.0126907f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_354 N_A_399_415#_c_481_n N_A_949_335#_M1013_g 0.0176904f $X=4.505 $Y=0.765
+ $X2=0 $Y2=0
cc_355 N_A_399_415#_c_484_n N_A_949_335#_M1013_g 4.38684e-19 $X=4.31 $Y=0.75
+ $X2=0 $Y2=0
cc_356 N_A_399_415#_c_487_n N_A_949_335#_M1013_g 3.11485e-19 $X=4.505 $Y=0.93
+ $X2=0 $Y2=0
cc_357 N_A_399_415#_c_488_n N_A_949_335#_M1013_g 0.0175551f $X=4.505 $Y=0.93
+ $X2=0 $Y2=0
cc_358 N_A_399_415#_c_486_n N_A_949_335#_c_598_n 5.56491e-19 $X=4.31 $Y=1.67
+ $X2=0 $Y2=0
cc_359 N_A_399_415#_c_489_n N_A_949_335#_c_598_n 7.76352e-19 $X=4.395 $Y=1.585
+ $X2=0 $Y2=0
cc_360 N_A_399_415#_c_486_n N_A_949_335#_c_614_n 2.93746e-19 $X=4.31 $Y=1.67
+ $X2=0 $Y2=0
cc_361 N_A_399_415#_c_488_n N_A_949_335#_c_599_n 0.0175551f $X=4.505 $Y=0.93
+ $X2=0 $Y2=0
cc_362 N_A_399_415#_c_492_n N_A_949_335#_c_599_n 3.11485e-19 $X=4.477 $Y=1.435
+ $X2=0 $Y2=0
cc_363 N_A_399_415#_M1002_g N_A_744_415#_c_737_n 0.00485005f $X=3.595 $Y=2.575
+ $X2=0 $Y2=0
cc_364 N_A_399_415#_c_486_n N_A_744_415#_c_737_n 0.0174719f $X=4.31 $Y=1.67
+ $X2=0 $Y2=0
cc_365 N_A_399_415#_M1002_g N_A_744_415#_c_744_n 0.0207918f $X=3.595 $Y=2.575
+ $X2=0 $Y2=0
cc_366 N_A_399_415#_c_481_n N_A_744_415#_c_745_n 0.00926342f $X=4.505 $Y=0.765
+ $X2=0 $Y2=0
cc_367 N_A_399_415#_c_484_n N_A_744_415#_c_745_n 0.038845f $X=4.31 $Y=0.75 $X2=0
+ $Y2=0
cc_368 N_A_399_415#_c_488_n N_A_744_415#_c_745_n 0.00165244f $X=4.505 $Y=0.93
+ $X2=0 $Y2=0
cc_369 N_A_399_415#_c_486_n N_A_744_415#_c_738_n 0.00945374f $X=4.31 $Y=1.67
+ $X2=0 $Y2=0
cc_370 N_A_399_415#_c_488_n N_A_744_415#_c_738_n 0.00145181f $X=4.505 $Y=0.93
+ $X2=0 $Y2=0
cc_371 N_A_399_415#_c_492_n N_A_744_415#_c_738_n 0.00476986f $X=4.477 $Y=1.435
+ $X2=0 $Y2=0
cc_372 N_A_399_415#_c_481_n N_A_744_415#_c_732_n 0.00348143f $X=4.505 $Y=0.765
+ $X2=0 $Y2=0
cc_373 N_A_399_415#_c_484_n N_A_744_415#_c_732_n 0.0134649f $X=4.31 $Y=0.75
+ $X2=0 $Y2=0
cc_374 N_A_399_415#_c_487_n N_A_744_415#_c_732_n 0.0423764f $X=4.505 $Y=0.93
+ $X2=0 $Y2=0
cc_375 N_A_399_415#_c_488_n N_A_744_415#_c_732_n 0.0039312f $X=4.505 $Y=0.93
+ $X2=0 $Y2=0
cc_376 N_A_399_415#_c_486_n N_A_744_415#_c_734_n 0.00899499f $X=4.31 $Y=1.67
+ $X2=0 $Y2=0
cc_377 N_A_399_415#_c_489_n N_A_744_415#_c_734_n 0.0077007f $X=4.395 $Y=1.585
+ $X2=0 $Y2=0
cc_378 N_A_399_415#_c_492_n N_A_744_415#_c_734_n 8.086e-19 $X=4.477 $Y=1.435
+ $X2=0 $Y2=0
cc_379 N_A_399_415#_M1002_g N_VPWR_c_880_n 0.0050932f $X=3.595 $Y=2.575 $X2=0
+ $Y2=0
cc_380 N_A_399_415#_M1002_g N_VPWR_c_887_n 0.00941859f $X=3.595 $Y=2.575 $X2=0
+ $Y2=0
cc_381 N_A_399_415#_M1002_g N_VPWR_c_878_n 0.0173779f $X=3.595 $Y=2.575 $X2=0
+ $Y2=0
cc_382 N_A_399_415#_c_483_n N_VGND_c_977_n 0.0191205f $X=2.48 $Y=0.47 $X2=0
+ $Y2=0
cc_383 N_A_399_415#_c_485_n N_VGND_c_977_n 0.0118783f $X=2.645 $Y=0.75 $X2=0
+ $Y2=0
cc_384 N_A_399_415#_c_483_n N_VGND_c_978_n 0.00736062f $X=2.48 $Y=0.47 $X2=0
+ $Y2=0
cc_385 N_A_399_415#_c_484_n N_VGND_c_978_n 0.019245f $X=4.31 $Y=0.75 $X2=0 $Y2=0
cc_386 N_A_399_415#_c_481_n N_VGND_c_981_n 0.00366111f $X=4.505 $Y=0.765 $X2=0
+ $Y2=0
cc_387 N_A_399_415#_c_484_n N_VGND_c_981_n 0.00974987f $X=4.31 $Y=0.75 $X2=0
+ $Y2=0
cc_388 N_A_399_415#_M1018_s N_VGND_c_986_n 0.00232985f $X=2.335 $Y=0.235 $X2=0
+ $Y2=0
cc_389 N_A_399_415#_c_481_n N_VGND_c_986_n 0.0059822f $X=4.505 $Y=0.765 $X2=0
+ $Y2=0
cc_390 N_A_399_415#_c_483_n N_VGND_c_986_n 0.0124057f $X=2.48 $Y=0.47 $X2=0
+ $Y2=0
cc_391 N_A_399_415#_c_484_n N_VGND_c_986_n 0.0173529f $X=4.31 $Y=0.75 $X2=0
+ $Y2=0
cc_392 N_A_399_415#_c_485_n N_VGND_c_986_n 0.018931f $X=2.645 $Y=0.75 $X2=0
+ $Y2=0
cc_393 N_A_949_335#_M1009_g N_A_744_415#_M1021_g 0.0176611f $X=4.87 $Y=2.575
+ $X2=0 $Y2=0
cc_394 N_A_949_335#_c_614_n N_A_744_415#_M1021_g 0.00163556f $X=4.902 $Y=1.825
+ $X2=0 $Y2=0
cc_395 N_A_949_335#_c_615_n N_A_744_415#_M1021_g 0.00436783f $X=6.03 $Y=2.225
+ $X2=0 $Y2=0
cc_396 N_A_949_335#_c_632_p N_A_744_415#_M1021_g 0.0150723f $X=6.03 $Y=2.9 $X2=0
+ $Y2=0
cc_397 N_A_949_335#_c_604_n N_A_744_415#_c_729_n 0.00840989f $X=5.985 $Y=0.94
+ $X2=0 $Y2=0
cc_398 N_A_949_335#_c_602_n N_A_744_415#_c_730_n 0.0123432f $X=5.82 $Y=0.495
+ $X2=0 $Y2=0
cc_399 N_A_949_335#_c_602_n N_A_744_415#_c_731_n 0.00534835f $X=5.82 $Y=0.495
+ $X2=0 $Y2=0
cc_400 N_A_949_335#_c_603_n N_A_744_415#_c_731_n 0.00717156f $X=6.68 $Y=0.94
+ $X2=0 $Y2=0
cc_401 N_A_949_335#_c_604_n N_A_744_415#_c_731_n 0.00358703f $X=5.985 $Y=0.94
+ $X2=0 $Y2=0
cc_402 N_A_949_335#_c_608_n N_A_744_415#_c_731_n 0.0129126f $X=5.34 $Y=1.02
+ $X2=0 $Y2=0
cc_403 N_A_949_335#_M1009_g N_A_744_415#_c_744_n 0.00362885f $X=4.87 $Y=2.575
+ $X2=0 $Y2=0
cc_404 N_A_949_335#_M1013_g N_A_744_415#_c_745_n 0.00674168f $X=4.985 $Y=0.445
+ $X2=0 $Y2=0
cc_405 N_A_949_335#_M1009_g N_A_744_415#_c_738_n 0.0211488f $X=4.87 $Y=2.575
+ $X2=0 $Y2=0
cc_406 N_A_949_335#_M1013_g N_A_744_415#_c_732_n 0.0103405f $X=4.985 $Y=0.445
+ $X2=0 $Y2=0
cc_407 N_A_949_335#_c_598_n N_A_744_415#_c_732_n 0.0118777f $X=4.902 $Y=1.675
+ $X2=0 $Y2=0
cc_408 N_A_949_335#_c_599_n N_A_744_415#_c_732_n 0.00878822f $X=4.985 $Y=1.02
+ $X2=0 $Y2=0
cc_409 N_A_949_335#_c_602_n N_A_744_415#_c_732_n 0.00484282f $X=5.82 $Y=0.495
+ $X2=0 $Y2=0
cc_410 N_A_949_335#_c_604_n N_A_744_415#_c_732_n 0.0233345f $X=5.985 $Y=0.94
+ $X2=0 $Y2=0
cc_411 N_A_949_335#_M1009_g N_A_744_415#_c_747_n 0.010683f $X=4.87 $Y=2.575
+ $X2=0 $Y2=0
cc_412 N_A_949_335#_c_614_n N_A_744_415#_c_747_n 0.00326272f $X=4.902 $Y=1.825
+ $X2=0 $Y2=0
cc_413 N_A_949_335#_c_598_n N_A_744_415#_c_733_n 0.00773684f $X=4.902 $Y=1.675
+ $X2=0 $Y2=0
cc_414 N_A_949_335#_c_614_n N_A_744_415#_c_733_n 0.0040907f $X=4.902 $Y=1.825
+ $X2=0 $Y2=0
cc_415 N_A_949_335#_c_604_n N_A_744_415#_c_733_n 0.027914f $X=5.985 $Y=0.94
+ $X2=0 $Y2=0
cc_416 N_A_949_335#_c_608_n N_A_744_415#_c_733_n 0.005857f $X=5.34 $Y=1.02 $X2=0
+ $Y2=0
cc_417 N_A_949_335#_c_598_n N_A_744_415#_c_734_n 0.00583722f $X=4.902 $Y=1.675
+ $X2=0 $Y2=0
cc_418 N_A_949_335#_c_614_n N_A_744_415#_c_734_n 0.00425033f $X=4.902 $Y=1.825
+ $X2=0 $Y2=0
cc_419 N_A_949_335#_c_598_n N_A_744_415#_c_735_n 0.0128703f $X=4.902 $Y=1.675
+ $X2=0 $Y2=0
cc_420 N_A_949_335#_c_615_n N_A_744_415#_c_735_n 4.08477e-19 $X=6.03 $Y=2.225
+ $X2=0 $Y2=0
cc_421 N_A_949_335#_c_604_n N_A_744_415#_c_735_n 0.00851725f $X=5.985 $Y=0.94
+ $X2=0 $Y2=0
cc_422 N_A_949_335#_c_608_n N_A_744_415#_c_735_n 0.00693868f $X=5.34 $Y=1.02
+ $X2=0 $Y2=0
cc_423 N_A_949_335#_M1017_g N_RESET_B_M1008_g 0.0272672f $X=6.93 $Y=2.575 $X2=0
+ $Y2=0
cc_424 N_A_949_335#_c_615_n N_RESET_B_M1008_g 9.82838e-19 $X=6.03 $Y=2.225 $X2=0
+ $Y2=0
cc_425 N_A_949_335#_c_632_p N_RESET_B_M1008_g 0.0153275f $X=6.03 $Y=2.9 $X2=0
+ $Y2=0
cc_426 N_A_949_335#_c_616_n N_RESET_B_M1008_g 0.0184094f $X=6.68 $Y=2.14 $X2=0
+ $Y2=0
cc_427 N_A_949_335#_c_607_n N_RESET_B_M1008_g 0.00356794f $X=6.765 $Y=2.055
+ $X2=0 $Y2=0
cc_428 N_A_949_335#_M1011_g N_RESET_B_M1006_g 0.0154215f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_429 N_A_949_335#_c_600_n N_RESET_B_M1006_g 0.0183319f $X=7.185 $Y=0.93 $X2=0
+ $Y2=0
cc_430 N_A_949_335#_c_602_n N_RESET_B_M1006_g 0.00201249f $X=5.82 $Y=0.495 $X2=0
+ $Y2=0
cc_431 N_A_949_335#_c_603_n N_RESET_B_M1006_g 0.0114183f $X=6.68 $Y=0.94 $X2=0
+ $Y2=0
cc_432 N_A_949_335#_c_606_n N_RESET_B_M1006_g 0.00401419f $X=6.86 $Y=1.345 $X2=0
+ $Y2=0
cc_433 N_A_949_335#_M1017_g N_RESET_B_c_829_n 0.0141794f $X=6.93 $Y=2.575 $X2=0
+ $Y2=0
cc_434 N_A_949_335#_c_601_n N_RESET_B_c_829_n 0.0103532f $X=6.882 $Y=1.525 $X2=0
+ $Y2=0
cc_435 N_A_949_335#_c_610_n N_RESET_B_c_829_n 7.36481e-19 $X=6.86 $Y=1.525 $X2=0
+ $Y2=0
cc_436 N_A_949_335#_c_616_n N_RESET_B_c_834_n 0.00208225f $X=6.68 $Y=2.14 $X2=0
+ $Y2=0
cc_437 N_A_949_335#_c_607_n N_RESET_B_c_834_n 7.36481e-19 $X=6.765 $Y=2.055
+ $X2=0 $Y2=0
cc_438 N_A_949_335#_c_603_n N_RESET_B_c_830_n 0.00469967f $X=6.68 $Y=0.94 $X2=0
+ $Y2=0
cc_439 N_A_949_335#_c_606_n N_RESET_B_c_830_n 7.36481e-19 $X=6.86 $Y=1.345 $X2=0
+ $Y2=0
cc_440 N_A_949_335#_c_609_n N_RESET_B_c_830_n 0.0103532f $X=6.875 $Y=1.02 $X2=0
+ $Y2=0
cc_441 N_A_949_335#_M1017_g N_RESET_B_c_831_n 3.61355e-19 $X=6.93 $Y=2.575 $X2=0
+ $Y2=0
cc_442 N_A_949_335#_c_615_n N_RESET_B_c_831_n 0.0274639f $X=6.03 $Y=2.225 $X2=0
+ $Y2=0
cc_443 N_A_949_335#_c_603_n N_RESET_B_c_831_n 0.0394278f $X=6.68 $Y=0.94 $X2=0
+ $Y2=0
cc_444 N_A_949_335#_c_604_n N_RESET_B_c_831_n 0.00826237f $X=5.985 $Y=0.94 $X2=0
+ $Y2=0
cc_445 N_A_949_335#_c_616_n N_RESET_B_c_831_n 0.0223243f $X=6.68 $Y=2.14 $X2=0
+ $Y2=0
cc_446 N_A_949_335#_c_606_n N_RESET_B_c_831_n 0.0519429f $X=6.86 $Y=1.345 $X2=0
+ $Y2=0
cc_447 N_A_949_335#_c_609_n N_RESET_B_c_831_n 3.75692e-19 $X=6.875 $Y=1.02 $X2=0
+ $Y2=0
cc_448 N_A_949_335#_c_616_n N_VPWR_M1008_d 0.00398712f $X=6.68 $Y=2.14 $X2=0
+ $Y2=0
cc_449 N_A_949_335#_M1009_g N_VPWR_c_881_n 0.0267415f $X=4.87 $Y=2.575 $X2=0
+ $Y2=0
cc_450 N_A_949_335#_c_615_n N_VPWR_c_881_n 0.00787512f $X=6.03 $Y=2.225 $X2=0
+ $Y2=0
cc_451 N_A_949_335#_c_632_p N_VPWR_c_881_n 0.0366224f $X=6.03 $Y=2.9 $X2=0 $Y2=0
cc_452 N_A_949_335#_M1017_g N_VPWR_c_882_n 0.0105403f $X=6.93 $Y=2.575 $X2=0
+ $Y2=0
cc_453 N_A_949_335#_c_632_p N_VPWR_c_882_n 0.0434878f $X=6.03 $Y=2.9 $X2=0 $Y2=0
cc_454 N_A_949_335#_c_616_n N_VPWR_c_882_n 0.0212953f $X=6.68 $Y=2.14 $X2=0
+ $Y2=0
cc_455 N_A_949_335#_M1009_g N_VPWR_c_887_n 0.00941859f $X=4.87 $Y=2.575 $X2=0
+ $Y2=0
cc_456 N_A_949_335#_c_632_p N_VPWR_c_889_n 0.0177952f $X=6.03 $Y=2.9 $X2=0 $Y2=0
cc_457 N_A_949_335#_M1017_g N_VPWR_c_890_n 0.00906878f $X=6.93 $Y=2.575 $X2=0
+ $Y2=0
cc_458 N_A_949_335#_M1009_g N_VPWR_c_878_n 0.0175196f $X=4.87 $Y=2.575 $X2=0
+ $Y2=0
cc_459 N_A_949_335#_M1017_g N_VPWR_c_878_n 0.0172612f $X=6.93 $Y=2.575 $X2=0
+ $Y2=0
cc_460 N_A_949_335#_c_632_p N_VPWR_c_878_n 0.0124497f $X=6.03 $Y=2.9 $X2=0 $Y2=0
cc_461 N_A_949_335#_M1011_g Q 0.00201375f $X=6.825 $Y=0.495 $X2=0 $Y2=0
cc_462 N_A_949_335#_M1014_g Q 0.013846f $X=7.185 $Y=0.495 $X2=0 $Y2=0
cc_463 N_A_949_335#_c_600_n Q 0.00623432f $X=7.185 $Y=0.93 $X2=0 $Y2=0
cc_464 N_A_949_335#_c_605_n Q 0.0121963f $X=6.86 $Y=1.025 $X2=0 $Y2=0
cc_465 N_A_949_335#_c_606_n Q 0.0358261f $X=6.86 $Y=1.345 $X2=0 $Y2=0
cc_466 N_A_949_335#_c_607_n Q 0.0217473f $X=6.765 $Y=2.055 $X2=0 $Y2=0
cc_467 N_A_949_335#_c_609_n Q 0.0246345f $X=6.875 $Y=1.02 $X2=0 $Y2=0
cc_468 N_A_949_335#_M1017_g Q 0.00648543f $X=6.93 $Y=2.575 $X2=0 $Y2=0
cc_469 N_A_949_335#_c_616_n Q 0.013428f $X=6.68 $Y=2.14 $X2=0 $Y2=0
cc_470 N_A_949_335#_c_610_n Q 2.65009e-19 $X=6.86 $Y=1.525 $X2=0 $Y2=0
cc_471 N_A_949_335#_M1017_g Q 0.012507f $X=6.93 $Y=2.575 $X2=0 $Y2=0
cc_472 N_A_949_335#_M1013_g N_VGND_c_979_n 0.0140723f $X=4.985 $Y=0.445 $X2=0
+ $Y2=0
cc_473 N_A_949_335#_c_602_n N_VGND_c_979_n 0.0270728f $X=5.82 $Y=0.495 $X2=0
+ $Y2=0
cc_474 N_A_949_335#_c_604_n N_VGND_c_979_n 0.0196411f $X=5.985 $Y=0.94 $X2=0
+ $Y2=0
cc_475 N_A_949_335#_c_608_n N_VGND_c_979_n 0.00194826f $X=5.34 $Y=1.02 $X2=0
+ $Y2=0
cc_476 N_A_949_335#_M1011_g N_VGND_c_980_n 0.0112546f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_477 N_A_949_335#_M1014_g N_VGND_c_980_n 0.00197591f $X=7.185 $Y=0.495 $X2=0
+ $Y2=0
cc_478 N_A_949_335#_c_602_n N_VGND_c_980_n 0.0137175f $X=5.82 $Y=0.495 $X2=0
+ $Y2=0
cc_479 N_A_949_335#_c_603_n N_VGND_c_980_n 0.0154557f $X=6.68 $Y=0.94 $X2=0
+ $Y2=0
cc_480 N_A_949_335#_c_605_n N_VGND_c_980_n 0.00525394f $X=6.86 $Y=1.025 $X2=0
+ $Y2=0
cc_481 N_A_949_335#_M1013_g N_VGND_c_981_n 0.00461015f $X=4.985 $Y=0.445 $X2=0
+ $Y2=0
cc_482 N_A_949_335#_c_602_n N_VGND_c_984_n 0.0220321f $X=5.82 $Y=0.495 $X2=0
+ $Y2=0
cc_483 N_A_949_335#_M1011_g N_VGND_c_985_n 0.00445056f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_484 N_A_949_335#_M1014_g N_VGND_c_985_n 0.00502664f $X=7.185 $Y=0.495 $X2=0
+ $Y2=0
cc_485 N_A_949_335#_M1013_g N_VGND_c_986_n 0.00958812f $X=4.985 $Y=0.445 $X2=0
+ $Y2=0
cc_486 N_A_949_335#_M1011_g N_VGND_c_986_n 0.00425628f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_487 N_A_949_335#_M1014_g N_VGND_c_986_n 0.0100616f $X=7.185 $Y=0.495 $X2=0
+ $Y2=0
cc_488 N_A_949_335#_c_602_n N_VGND_c_986_n 0.0125808f $X=5.82 $Y=0.495 $X2=0
+ $Y2=0
cc_489 N_A_949_335#_c_603_n N_VGND_c_986_n 0.0146623f $X=6.68 $Y=0.94 $X2=0
+ $Y2=0
cc_490 N_A_949_335#_c_604_n N_VGND_c_986_n 0.00853275f $X=5.985 $Y=0.94 $X2=0
+ $Y2=0
cc_491 N_A_949_335#_c_605_n N_VGND_c_986_n 0.0091484f $X=6.86 $Y=1.025 $X2=0
+ $Y2=0
cc_492 N_A_949_335#_c_608_n N_VGND_c_986_n 0.00258753f $X=5.34 $Y=1.02 $X2=0
+ $Y2=0
cc_493 N_A_744_415#_c_729_n N_RESET_B_M1006_g 0.00918799f $X=5.885 $Y=1.425
+ $X2=0 $Y2=0
cc_494 N_A_744_415#_c_730_n N_RESET_B_M1006_g 0.0489213f $X=6.035 $Y=0.815 $X2=0
+ $Y2=0
cc_495 N_A_744_415#_c_735_n N_RESET_B_c_829_n 0.0178008f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_496 N_A_744_415#_M1021_g N_RESET_B_c_834_n 0.022787f $X=5.765 $Y=2.575 $X2=0
+ $Y2=0
cc_497 N_A_744_415#_c_729_n N_RESET_B_c_830_n 0.0178008f $X=5.885 $Y=1.425 $X2=0
+ $Y2=0
cc_498 N_A_744_415#_M1021_g N_RESET_B_c_831_n 0.00692274f $X=5.765 $Y=2.575
+ $X2=0 $Y2=0
cc_499 N_A_744_415#_c_729_n N_RESET_B_c_831_n 0.0141128f $X=5.885 $Y=1.425 $X2=0
+ $Y2=0
cc_500 N_A_744_415#_c_731_n N_RESET_B_c_831_n 0.00101235f $X=6.035 $Y=0.89 $X2=0
+ $Y2=0
cc_501 N_A_744_415#_c_733_n N_RESET_B_c_831_n 0.0263058f $X=5.54 $Y=1.59 $X2=0
+ $Y2=0
cc_502 N_A_744_415#_c_735_n N_RESET_B_c_831_n 0.0113798f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_503 N_A_744_415#_M1021_g N_VPWR_c_881_n 0.016764f $X=5.765 $Y=2.575 $X2=0
+ $Y2=0
cc_504 N_A_744_415#_c_738_n N_VPWR_c_881_n 0.0134301f $X=4.825 $Y=2.14 $X2=0
+ $Y2=0
cc_505 N_A_744_415#_c_733_n N_VPWR_c_881_n 0.0189814f $X=5.54 $Y=1.59 $X2=0
+ $Y2=0
cc_506 N_A_744_415#_c_735_n N_VPWR_c_881_n 0.00278824f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_507 N_A_744_415#_M1021_g N_VPWR_c_882_n 8.39432e-19 $X=5.765 $Y=2.575 $X2=0
+ $Y2=0
cc_508 N_A_744_415#_c_744_n N_VPWR_c_887_n 0.0197322f $X=4.115 $Y=2.9 $X2=0
+ $Y2=0
cc_509 N_A_744_415#_M1021_g N_VPWR_c_889_n 0.00906878f $X=5.765 $Y=2.575 $X2=0
+ $Y2=0
cc_510 N_A_744_415#_M1021_g N_VPWR_c_878_n 0.016724f $X=5.765 $Y=2.575 $X2=0
+ $Y2=0
cc_511 N_A_744_415#_c_744_n N_VPWR_c_878_n 0.0125705f $X=4.115 $Y=2.9 $X2=0
+ $Y2=0
cc_512 N_A_744_415#_c_738_n A_901_415# 0.0048076f $X=4.825 $Y=2.14 $X2=-0.19
+ $Y2=-0.245
cc_513 N_A_744_415#_c_745_n N_VGND_c_978_n 0.00573659f $X=4.825 $Y=0.39 $X2=0
+ $Y2=0
cc_514 N_A_744_415#_c_730_n N_VGND_c_979_n 0.00254767f $X=6.035 $Y=0.815 $X2=0
+ $Y2=0
cc_515 N_A_744_415#_c_745_n N_VGND_c_979_n 0.0146778f $X=4.825 $Y=0.39 $X2=0
+ $Y2=0
cc_516 N_A_744_415#_c_732_n N_VGND_c_979_n 0.013153f $X=4.91 $Y=1.425 $X2=0
+ $Y2=0
cc_517 N_A_744_415#_c_730_n N_VGND_c_980_n 0.00197591f $X=6.035 $Y=0.815 $X2=0
+ $Y2=0
cc_518 N_A_744_415#_c_745_n N_VGND_c_981_n 0.0451579f $X=4.825 $Y=0.39 $X2=0
+ $Y2=0
cc_519 N_A_744_415#_c_730_n N_VGND_c_984_n 0.00502664f $X=6.035 $Y=0.815 $X2=0
+ $Y2=0
cc_520 N_A_744_415#_M1020_d N_VGND_c_986_n 0.00350385f $X=3.95 $Y=0.235 $X2=0
+ $Y2=0
cc_521 N_A_744_415#_c_730_n N_VGND_c_986_n 0.0066094f $X=6.035 $Y=0.815 $X2=0
+ $Y2=0
cc_522 N_A_744_415#_c_745_n N_VGND_c_986_n 0.0343632f $X=4.825 $Y=0.39 $X2=0
+ $Y2=0
cc_523 N_A_744_415#_c_745_n A_898_47# 0.0109154f $X=4.825 $Y=0.39 $X2=-0.19
+ $Y2=-0.245
cc_524 N_A_744_415#_c_732_n A_898_47# 0.0022425f $X=4.91 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_525 N_RESET_B_M1008_g N_VPWR_c_882_n 0.0166465f $X=6.295 $Y=2.575 $X2=0 $Y2=0
cc_526 N_RESET_B_M1008_g N_VPWR_c_889_n 0.00810976f $X=6.295 $Y=2.575 $X2=0
+ $Y2=0
cc_527 N_RESET_B_M1008_g N_VPWR_c_878_n 0.0135863f $X=6.295 $Y=2.575 $X2=0 $Y2=0
cc_528 N_RESET_B_M1008_g Q 7.7349e-19 $X=6.295 $Y=2.575 $X2=0 $Y2=0
cc_529 N_RESET_B_M1006_g N_VGND_c_980_n 0.0112556f $X=6.395 $Y=0.495 $X2=0 $Y2=0
cc_530 N_RESET_B_M1006_g N_VGND_c_984_n 0.00445056f $X=6.395 $Y=0.495 $X2=0
+ $Y2=0
cc_531 N_RESET_B_M1006_g N_VGND_c_986_n 0.00428592f $X=6.395 $Y=0.495 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_882_n Q 0.0339178f $X=6.56 $Y=2.57 $X2=0 $Y2=0
cc_533 N_VPWR_c_890_n Q 0.03358f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_534 N_VPWR_c_878_n Q 0.0205026f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_535 Q N_VGND_c_980_n 0.0137175f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_536 Q N_VGND_c_985_n 0.0220321f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_537 Q N_VGND_c_986_n 0.0125808f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_538 A_114_47# N_VGND_c_986_n 0.00829524f $X=0.57 $Y=0.235 $X2=7.44 $Y2=0
cc_539 N_VGND_c_986_n A_272_47# 0.00922959f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
cc_540 N_VGND_c_986_n A_554_47# 0.00253354f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
cc_541 N_VGND_c_986_n A_712_47# 0.00289547f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
cc_542 N_VGND_c_986_n A_898_47# 0.00343004f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
