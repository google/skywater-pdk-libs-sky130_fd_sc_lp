* NGSPICE file created from sky130_fd_sc_lp__buf_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__buf_4 A VGND VNB VPB VPWR X
M1000 a_122_23# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=1.0647e+12p ps=9.25e+06u
M1001 a_122_23# A VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=6.93e+11p ps=6.69e+06u
M1002 VGND a_122_23# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1003 X a_122_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_122_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1005 VPWR a_122_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_122_23# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_122_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_122_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_122_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

