* File: sky130_fd_sc_lp__o221ai_lp.pxi.spice
* Created: Wed Sep  2 10:19:26 2020
* 
x_PM_SKY130_FD_SC_LP__O221AI_LP%C1 N_C1_c_77_n N_C1_M1003_g N_C1_M1004_g C1
+ PM_SKY130_FD_SC_LP__O221AI_LP%C1
x_PM_SKY130_FD_SC_LP__O221AI_LP%B1 N_B1_M1006_g N_B1_c_113_n N_B1_M1007_g
+ N_B1_c_118_n B1 B1 N_B1_c_115_n PM_SKY130_FD_SC_LP__O221AI_LP%B1
x_PM_SKY130_FD_SC_LP__O221AI_LP%B2 N_B2_M1001_g N_B2_M1002_g N_B2_c_165_n
+ N_B2_c_160_n N_B2_c_161_n B2 B2 N_B2_c_162_n N_B2_c_163_n
+ PM_SKY130_FD_SC_LP__O221AI_LP%B2
x_PM_SKY130_FD_SC_LP__O221AI_LP%A2 N_A2_M1000_g N_A2_c_221_n N_A2_c_222_n
+ N_A2_c_228_n N_A2_M1005_g N_A2_c_223_n N_A2_c_224_n N_A2_c_225_n A2 A2
+ N_A2_c_227_n PM_SKY130_FD_SC_LP__O221AI_LP%A2
x_PM_SKY130_FD_SC_LP__O221AI_LP%A1 N_A1_c_289_n N_A1_M1008_g N_A1_M1009_g
+ N_A1_c_284_n N_A1_c_285_n N_A1_c_286_n A1 N_A1_c_287_n N_A1_c_288_n
+ PM_SKY130_FD_SC_LP__O221AI_LP%A1
x_PM_SKY130_FD_SC_LP__O221AI_LP%Y N_Y_M1004_s N_Y_M1003_s N_Y_M1001_d
+ N_Y_c_331_n N_Y_c_332_n N_Y_c_339_n N_Y_c_348_n Y Y N_Y_c_333_n
+ PM_SKY130_FD_SC_LP__O221AI_LP%Y
x_PM_SKY130_FD_SC_LP__O221AI_LP%VPWR N_VPWR_M1003_d N_VPWR_M1008_d
+ N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n VPWR
+ N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_375_n N_VPWR_c_383_n
+ PM_SKY130_FD_SC_LP__O221AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O221AI_LP%A_216_55# N_A_216_55#_M1004_d
+ N_A_216_55#_M1002_d N_A_216_55#_c_422_n N_A_216_55#_c_423_n
+ N_A_216_55#_c_428_n N_A_216_55#_c_435_n N_A_216_55#_c_424_n
+ N_A_216_55#_c_425_n N_A_216_55#_c_426_n
+ PM_SKY130_FD_SC_LP__O221AI_LP%A_216_55#
x_PM_SKY130_FD_SC_LP__O221AI_LP%A_302_55# N_A_302_55#_M1006_d
+ N_A_302_55#_M1009_d N_A_302_55#_c_480_n N_A_302_55#_c_481_n
+ N_A_302_55#_c_482_n N_A_302_55#_c_483_n N_A_302_55#_c_484_n
+ N_A_302_55#_c_485_n PM_SKY130_FD_SC_LP__O221AI_LP%A_302_55#
x_PM_SKY130_FD_SC_LP__O221AI_LP%VGND N_VGND_M1000_d N_VGND_c_529_n VGND
+ N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n
+ PM_SKY130_FD_SC_LP__O221AI_LP%VGND
cc_1 VNB N_C1_c_77_n 0.0717242f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.72
cc_2 VNB N_C1_M1004_g 0.034644f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.485
cc_3 VNB C1 0.00403307f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_B1_M1006_g 0.0387699f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.595
cc_5 VNB N_B1_c_113_n 0.0242722f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.485
cc_6 VNB B1 0.0144939f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.215
cc_7 VNB N_B1_c_115_n 0.01999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B2_M1002_g 0.025415f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.485
cc_9 VNB N_B2_c_160_n 0.00256479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B2_c_161_n 0.00785218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_c_162_n 0.0619855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B2_c_163_n 0.0100346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_221_n 0.0225036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_222_n 0.0118532f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.05
cc_15 VNB N_A2_c_223_n 0.019116f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.215
cc_16 VNB N_A2_c_224_n 0.0330781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_225_n 0.0210016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A2 0.0153631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_227_n 0.0222551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_M1009_g 0.0276414f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_21 VNB N_A1_c_284_n 0.025285f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.215
cc_22 VNB N_A1_c_285_n 0.0154921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_286_n 0.00425307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_287_n 0.0186157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_288_n 0.0032218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_331_n 0.0224164f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.215
cc_27 VNB N_Y_c_332_n 0.0228906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_333_n 0.0471932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_375_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_216_55#_c_422_n 0.00207321f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_31 VNB N_A_216_55#_c_423_n 0.00552788f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.215
cc_32 VNB N_A_216_55#_c_424_n 0.0455692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_216_55#_c_425_n 0.00544733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_216_55#_c_426_n 0.0324748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_302_55#_c_480_n 0.00234627f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_36 VNB N_A_302_55#_c_481_n 0.00227415f $X=-0.19 $Y=-0.245 $X2=0.822 $Y2=1.215
cc_37 VNB N_A_302_55#_c_482_n 0.00685853f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.215
cc_38 VNB N_A_302_55#_c_483_n 0.00725966f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.215
cc_39 VNB N_A_302_55#_c_484_n 0.00420729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_302_55#_c_485_n 0.0110917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_529_n 0.00711907f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.485
cc_42 VNB N_VGND_c_530_n 0.0544804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_531_n 0.0516634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_532_n 0.260757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_533_n 0.00631679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_C1_c_77_n 0.0150605f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.72
cc_47 VPB N_C1_M1003_g 0.0452217f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.595
cc_48 VPB C1 0.00301611f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_49 VPB N_B1_c_113_n 4.90082e-19 $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.485
cc_50 VPB N_B1_M1007_g 0.0322116f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_51 VPB N_B1_c_118_n 0.0166279f $X=-0.19 $Y=1.655 $X2=0.822 $Y2=1.215
cc_52 VPB B1 0.00274635f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.215
cc_53 VPB N_B2_M1001_g 0.0259225f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.595
cc_54 VPB N_B2_c_165_n 0.0313584f $X=-0.19 $Y=1.655 $X2=0.822 $Y2=1.215
cc_55 VPB N_B2_c_160_n 7.47102e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_B2_c_161_n 0.0210125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_B2_c_163_n 0.00254836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A2_c_228_n 0.0093012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A2_M1005_g 0.0249422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A2_c_225_n 0.00858189f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A1_c_289_n 0.00982817f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.595
cc_62 VPB N_A1_M1008_g 0.0322697f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.05
cc_63 VPB N_A1_c_286_n 0.00910519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB Y 0.0813675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_Y_c_333_n 0.013851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_376_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_67 VPB N_VPWR_c_377_n 0.0267058f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.215
cc_68 VPB N_VPWR_c_378_n 0.0517503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_379_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_380_n 0.027607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_381_n 0.0253733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_375_n 0.0753475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_383_n 0.0051042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_216_55#_c_423_n 0.00369645f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.215
cc_75 VPB N_A_216_55#_c_428_n 0.0404892f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.215
cc_76 VPB N_A_216_55#_c_424_n 0.027389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 N_C1_M1004_g N_B1_M1006_g 0.0226088f $X=1.005 $Y=0.485 $X2=0 $Y2=0
cc_78 N_C1_c_77_n N_B1_c_113_n 0.0066511f $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_79 N_C1_M1003_g N_B1_M1007_g 0.0362644f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_80 N_C1_M1003_g N_B1_c_118_n 0.0066511f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_81 N_C1_c_77_n B1 6.24965e-19 $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_82 N_C1_c_77_n N_B1_c_115_n 0.0226088f $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_83 N_C1_c_77_n N_Y_c_332_n 0.00222488f $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_84 N_C1_M1004_g N_Y_c_332_n 0.00121798f $X=1.005 $Y=0.485 $X2=0 $Y2=0
cc_85 C1 N_Y_c_332_n 0.0169485f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_86 N_C1_M1003_g N_Y_c_339_n 0.0204364f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_87 N_C1_c_77_n Y 0.0023335f $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_88 N_C1_M1003_g Y 0.031324f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_89 C1 Y 0.0257173f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_C1_c_77_n N_Y_c_333_n 0.0157026f $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_91 N_C1_M1003_g N_Y_c_333_n 0.00483835f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_92 N_C1_M1004_g N_Y_c_333_n 0.00706922f $X=1.005 $Y=0.485 $X2=0 $Y2=0
cc_93 C1 N_Y_c_333_n 0.0377432f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_94 N_C1_M1003_g N_VPWR_c_376_n 0.0109035f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_95 N_C1_M1003_g N_VPWR_c_380_n 0.00638986f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_96 N_C1_M1003_g N_VPWR_c_375_n 0.00840643f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_97 N_C1_M1004_g N_A_216_55#_c_422_n 0.00659327f $X=1.005 $Y=0.485 $X2=0 $Y2=0
cc_98 N_C1_c_77_n N_A_216_55#_c_423_n 0.0164688f $X=0.975 $Y=1.72 $X2=0 $Y2=0
cc_99 N_C1_M1003_g N_A_216_55#_c_423_n 0.0153102f $X=0.975 $Y=2.595 $X2=0 $Y2=0
cc_100 N_C1_M1004_g N_A_216_55#_c_423_n 0.00728832f $X=1.005 $Y=0.485 $X2=0
+ $Y2=0
cc_101 C1 N_A_216_55#_c_423_n 0.0457028f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_102 N_C1_M1003_g N_A_216_55#_c_435_n 0.00647071f $X=0.975 $Y=2.595 $X2=0
+ $Y2=0
cc_103 N_C1_M1004_g N_A_216_55#_c_425_n 0.00909172f $X=1.005 $Y=0.485 $X2=0
+ $Y2=0
cc_104 N_C1_M1004_g N_VGND_c_530_n 0.00511657f $X=1.005 $Y=0.485 $X2=0 $Y2=0
cc_105 N_C1_M1004_g N_VGND_c_532_n 0.0106692f $X=1.005 $Y=0.485 $X2=0 $Y2=0
cc_106 N_B1_c_118_n N_B2_M1001_g 0.0466345f $X=1.547 $Y=1.85 $X2=0 $Y2=0
cc_107 N_B1_c_113_n N_B2_c_160_n 2.76303e-19 $X=1.547 $Y=1.663 $X2=0 $Y2=0
cc_108 N_B1_M1007_g N_B2_c_160_n 5.7458e-19 $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_109 B1 N_B2_c_160_n 0.0188249f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_B1_c_113_n N_B2_c_161_n 0.0466345f $X=1.547 $Y=1.663 $X2=0 $Y2=0
cc_111 B1 N_B2_c_161_n 0.00150812f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B1_M1006_g N_A2_c_223_n 0.0181547f $X=1.435 $Y=0.485 $X2=0 $Y2=0
cc_113 N_B1_M1006_g A2 7.57481e-19 $X=1.435 $Y=0.485 $X2=0 $Y2=0
cc_114 B1 A2 0.015932f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B1_c_115_n A2 5.02821e-19 $X=1.57 $Y=1.345 $X2=0 $Y2=0
cc_116 N_B1_M1006_g N_A2_c_227_n 0.00564752f $X=1.435 $Y=0.485 $X2=0 $Y2=0
cc_117 B1 N_A2_c_227_n 7.1075e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B1_c_115_n N_A2_c_227_n 0.00821742f $X=1.57 $Y=1.345 $X2=0 $Y2=0
cc_119 N_B1_M1007_g N_Y_c_339_n 0.017863f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_120 N_B1_M1007_g N_Y_c_348_n 0.00185644f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_121 N_B1_M1007_g Y 0.00174529f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_122 N_B1_M1007_g N_VPWR_c_376_n 0.0107066f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_123 N_B1_M1007_g N_VPWR_c_378_n 0.00722861f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_124 N_B1_M1007_g N_VPWR_c_375_n 0.00929854f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_125 N_B1_M1006_g N_A_216_55#_c_422_n 0.00590914f $X=1.435 $Y=0.485 $X2=0
+ $Y2=0
cc_126 N_B1_M1006_g N_A_216_55#_c_423_n 0.0106602f $X=1.435 $Y=0.485 $X2=0 $Y2=0
cc_127 N_B1_M1007_g N_A_216_55#_c_423_n 0.00526221f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_128 B1 N_A_216_55#_c_423_n 0.0487772f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B1_M1007_g N_A_216_55#_c_428_n 0.0160611f $X=1.61 $Y=2.595 $X2=0 $Y2=0
cc_130 N_B1_c_118_n N_A_216_55#_c_428_n 0.00207057f $X=1.547 $Y=1.85 $X2=0 $Y2=0
cc_131 B1 N_A_216_55#_c_428_n 0.0182867f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_M1006_g N_A_216_55#_c_425_n 0.00525934f $X=1.435 $Y=0.485 $X2=0
+ $Y2=0
cc_133 N_B1_M1006_g N_A_302_55#_c_480_n 0.00222789f $X=1.435 $Y=0.485 $X2=0
+ $Y2=0
cc_134 N_B1_M1006_g N_A_302_55#_c_482_n 0.00153797f $X=1.435 $Y=0.485 $X2=0
+ $Y2=0
cc_135 B1 N_A_302_55#_c_482_n 0.012682f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B1_c_115_n N_A_302_55#_c_482_n 0.00119949f $X=1.57 $Y=1.345 $X2=0 $Y2=0
cc_137 N_B1_M1006_g N_VGND_c_530_n 0.00511657f $X=1.435 $Y=0.485 $X2=0 $Y2=0
cc_138 N_B1_M1006_g N_VGND_c_532_n 0.00982809f $X=1.435 $Y=0.485 $X2=0 $Y2=0
cc_139 N_B2_c_165_n N_A2_c_222_n 0.00132975f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_140 N_B2_c_160_n N_A2_c_222_n 3.30281e-19 $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_141 N_B2_c_161_n N_A2_c_222_n 0.0157718f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_142 N_B2_M1001_g N_A2_c_228_n 0.038348f $X=2.1 $Y=2.595 $X2=0 $Y2=0
cc_143 N_B2_c_165_n N_A2_c_228_n 0.00985244f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_144 N_B2_c_160_n N_A2_c_224_n 2.66635e-19 $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_145 N_B2_c_161_n N_A2_c_224_n 6.48064e-19 $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_146 N_B2_c_165_n N_A2_c_225_n 0.00527006f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_147 N_B2_c_160_n N_A2_c_225_n 0.00115151f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_148 N_B2_c_161_n N_A2_c_225_n 0.0182524f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_149 N_B2_c_165_n A2 0.0204335f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_150 N_B2_c_160_n A2 0.0205769f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_151 N_B2_c_161_n A2 0.0010147f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_152 N_B2_c_165_n N_A1_c_289_n 0.0076706f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_153 N_B2_c_165_n N_A1_M1008_g 0.00359488f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_154 N_B2_M1002_g N_A1_M1009_g 0.0186797f $X=3.58 $Y=0.485 $X2=0 $Y2=0
cc_155 N_B2_c_163_n N_A1_M1009_g 4.25215e-19 $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_156 N_B2_c_162_n N_A1_c_284_n 0.0172421f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_157 N_B2_c_165_n N_A1_c_285_n 9.16733e-19 $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_158 N_B2_c_165_n N_A1_c_286_n 0.00405814f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_159 N_B2_c_163_n N_A1_c_286_n 0.00582181f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_160 N_B2_c_162_n N_A1_c_287_n 0.0172421f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_161 N_B2_c_163_n N_A1_c_287_n 0.00442226f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_162 N_B2_c_165_n N_A1_c_288_n 0.0245014f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_163 N_B2_c_162_n N_A1_c_288_n 7.99251e-19 $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_164 N_B2_c_163_n N_A1_c_288_n 0.0438819f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_165 N_B2_M1001_g N_Y_c_339_n 0.0158545f $X=2.1 $Y=2.595 $X2=0 $Y2=0
cc_166 N_B2_M1001_g N_Y_c_348_n 0.00985205f $X=2.1 $Y=2.595 $X2=0 $Y2=0
cc_167 N_B2_M1001_g N_VPWR_c_378_n 0.00712039f $X=2.1 $Y=2.595 $X2=0 $Y2=0
cc_168 N_B2_M1001_g N_VPWR_c_375_n 0.00906658f $X=2.1 $Y=2.595 $X2=0 $Y2=0
cc_169 N_B2_M1001_g N_A_216_55#_c_428_n 0.0149049f $X=2.1 $Y=2.595 $X2=0 $Y2=0
cc_170 N_B2_c_165_n N_A_216_55#_c_428_n 0.100841f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_171 N_B2_c_160_n N_A_216_55#_c_428_n 0.020685f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_172 N_B2_c_161_n N_A_216_55#_c_428_n 4.21457e-19 $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_173 N_B2_c_162_n N_A_216_55#_c_428_n 0.00105409f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_174 N_B2_M1002_g N_A_216_55#_c_424_n 0.00502213f $X=3.58 $Y=0.485 $X2=0 $Y2=0
cc_175 N_B2_c_165_n N_A_216_55#_c_424_n 0.0137879f $X=3.485 $Y=1.85 $X2=0 $Y2=0
cc_176 N_B2_c_162_n N_A_216_55#_c_424_n 0.0149053f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_177 N_B2_c_163_n N_A_216_55#_c_424_n 0.0636755f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_178 N_B2_M1002_g N_A_216_55#_c_426_n 0.0086871f $X=3.58 $Y=0.485 $X2=0 $Y2=0
cc_179 N_B2_c_162_n N_A_216_55#_c_426_n 9.23196e-19 $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_180 N_B2_c_163_n N_A_216_55#_c_426_n 0.0102029f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_181 N_B2_M1002_g N_A_302_55#_c_485_n 0.00612002f $X=3.58 $Y=0.485 $X2=0 $Y2=0
cc_182 N_B2_c_163_n N_A_302_55#_c_485_n 0.00353815f $X=3.67 $Y=1.06 $X2=0 $Y2=0
cc_183 N_B2_M1002_g N_VGND_c_531_n 0.00511657f $X=3.58 $Y=0.485 $X2=0 $Y2=0
cc_184 N_B2_M1002_g N_VGND_c_532_n 0.0105196f $X=3.58 $Y=0.485 $X2=0 $Y2=0
cc_185 N_A2_c_228_n N_A1_c_289_n 0.0402984f $X=2.67 $Y=1.95 $X2=0 $Y2=0
cc_186 N_A2_M1005_g N_A1_M1008_g 0.0402984f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_187 N_A2_c_221_n N_A1_c_284_n 0.0100162f $X=2.545 $Y=1.29 $X2=0 $Y2=0
cc_188 N_A2_c_227_n N_A1_c_284_n 0.00264104f $X=2.185 $Y=1.2 $X2=0 $Y2=0
cc_189 N_A2_c_225_n N_A1_c_285_n 0.0100162f $X=2.67 $Y=1.825 $X2=0 $Y2=0
cc_190 N_A2_c_225_n N_A1_c_286_n 0.00972034f $X=2.67 $Y=1.825 $X2=0 $Y2=0
cc_191 N_A2_c_224_n N_A1_c_287_n 0.00264104f $X=2.11 $Y=0.94 $X2=0 $Y2=0
cc_192 A2 N_A1_c_287_n 0.00314382f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_193 N_A2_c_221_n N_A1_c_288_n 2.17403e-19 $X=2.545 $Y=1.29 $X2=0 $Y2=0
cc_194 N_A2_c_224_n N_A1_c_288_n 6.87341e-19 $X=2.11 $Y=0.94 $X2=0 $Y2=0
cc_195 N_A2_c_225_n N_A1_c_288_n 0.00113647f $X=2.67 $Y=1.825 $X2=0 $Y2=0
cc_196 A2 N_A1_c_288_n 0.0300951f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A2_M1005_g N_VPWR_c_377_n 0.00362925f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_198 N_A2_M1005_g N_VPWR_c_378_n 0.00975641f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_199 N_A2_M1005_g N_VPWR_c_375_n 0.0172159f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_200 N_A2_M1005_g N_A_216_55#_c_428_n 0.0224632f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_201 N_A2_c_224_n N_A_216_55#_c_425_n 3.33984e-19 $X=2.11 $Y=0.94 $X2=0 $Y2=0
cc_202 N_A2_c_223_n N_A_302_55#_c_480_n 0.0109397f $X=2.11 $Y=0.79 $X2=0 $Y2=0
cc_203 N_A2_c_221_n N_A_302_55#_c_481_n 0.0010806f $X=2.545 $Y=1.29 $X2=0 $Y2=0
cc_204 N_A2_c_223_n N_A_302_55#_c_481_n 0.00654871f $X=2.11 $Y=0.79 $X2=0 $Y2=0
cc_205 N_A2_c_224_n N_A_302_55#_c_481_n 0.0186593f $X=2.11 $Y=0.94 $X2=0 $Y2=0
cc_206 A2 N_A_302_55#_c_481_n 0.040823f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_207 N_A2_c_223_n N_A_302_55#_c_482_n 0.00151577f $X=2.11 $Y=0.79 $X2=0 $Y2=0
cc_208 N_A2_c_224_n N_A_302_55#_c_482_n 0.00199177f $X=2.11 $Y=0.94 $X2=0 $Y2=0
cc_209 N_A2_c_221_n N_A_302_55#_c_484_n 5.19793e-19 $X=2.545 $Y=1.29 $X2=0 $Y2=0
cc_210 N_A2_c_223_n N_A_302_55#_c_484_n 0.00341398f $X=2.11 $Y=0.79 $X2=0 $Y2=0
cc_211 N_A2_c_224_n N_A_302_55#_c_484_n 2.54031e-19 $X=2.11 $Y=0.94 $X2=0 $Y2=0
cc_212 A2 N_A_302_55#_c_484_n 0.013564f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_213 N_A2_c_223_n N_VGND_c_529_n 0.00893094f $X=2.11 $Y=0.79 $X2=0 $Y2=0
cc_214 N_A2_c_224_n N_VGND_c_529_n 0.00162313f $X=2.11 $Y=0.94 $X2=0 $Y2=0
cc_215 N_A2_c_223_n N_VGND_c_530_n 0.00389854f $X=2.11 $Y=0.79 $X2=0 $Y2=0
cc_216 N_A2_c_223_n N_VGND_c_532_n 0.00661355f $X=2.11 $Y=0.79 $X2=0 $Y2=0
cc_217 N_A1_M1008_g N_VPWR_c_377_n 0.023694f $X=3.16 $Y=2.595 $X2=0 $Y2=0
cc_218 N_A1_M1008_g N_VPWR_c_378_n 0.008763f $X=3.16 $Y=2.595 $X2=0 $Y2=0
cc_219 N_A1_M1008_g N_VPWR_c_375_n 0.0144563f $X=3.16 $Y=2.595 $X2=0 $Y2=0
cc_220 N_A1_M1008_g N_A_216_55#_c_428_n 0.0235917f $X=3.16 $Y=2.595 $X2=0 $Y2=0
cc_221 N_A1_M1009_g N_A_302_55#_c_483_n 0.0102146f $X=3.15 $Y=0.485 $X2=0 $Y2=0
cc_222 N_A1_c_287_n N_A_302_55#_c_483_n 9.35231e-19 $X=3.1 $Y=1.08 $X2=0 $Y2=0
cc_223 N_A1_c_288_n N_A_302_55#_c_483_n 0.0181527f $X=3.1 $Y=1.08 $X2=0 $Y2=0
cc_224 N_A1_M1009_g N_A_302_55#_c_484_n 0.00465998f $X=3.15 $Y=0.485 $X2=0 $Y2=0
cc_225 N_A1_M1009_g N_A_302_55#_c_485_n 0.0142807f $X=3.15 $Y=0.485 $X2=0 $Y2=0
cc_226 N_A1_c_287_n N_A_302_55#_c_485_n 2.8619e-19 $X=3.1 $Y=1.08 $X2=0 $Y2=0
cc_227 N_A1_c_288_n N_A_302_55#_c_485_n 0.00469802f $X=3.1 $Y=1.08 $X2=0 $Y2=0
cc_228 N_A1_M1009_g N_VGND_c_529_n 0.00693297f $X=3.15 $Y=0.485 $X2=0 $Y2=0
cc_229 N_A1_M1009_g N_VGND_c_531_n 0.00373861f $X=3.15 $Y=0.485 $X2=0 $Y2=0
cc_230 N_A1_M1009_g N_VGND_c_532_n 0.00631877f $X=3.15 $Y=0.485 $X2=0 $Y2=0
cc_231 N_Y_c_339_n N_VPWR_M1003_d 0.0061526f $X=2.2 $Y=2.55 $X2=-0.19 $Y2=-0.245
cc_232 N_Y_c_339_n N_VPWR_c_376_n 0.0198473f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_233 Y N_VPWR_c_376_n 0.0174391f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_234 N_Y_c_339_n N_VPWR_c_378_n 0.0104803f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_235 N_Y_c_348_n N_VPWR_c_378_n 0.0182904f $X=2.365 $Y=2.765 $X2=0 $Y2=0
cc_236 N_Y_c_339_n N_VPWR_c_380_n 0.00284377f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_237 Y N_VPWR_c_380_n 0.0480763f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_238 N_Y_M1003_s N_VPWR_c_375_n 0.0023218f $X=0.565 $Y=2.095 $X2=0 $Y2=0
cc_239 N_Y_M1001_d N_VPWR_c_375_n 0.00313279f $X=2.225 $Y=2.095 $X2=0 $Y2=0
cc_240 N_Y_c_339_n N_VPWR_c_375_n 0.0251718f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_241 N_Y_c_348_n N_VPWR_c_375_n 0.0125379f $X=2.365 $Y=2.765 $X2=0 $Y2=0
cc_242 Y N_VPWR_c_375_n 0.0287592f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_243 N_Y_c_339_n A_347_419# 0.00369683f $X=2.2 $Y=2.55 $X2=-0.19 $Y2=-0.245
cc_244 N_Y_c_332_n N_A_216_55#_c_422_n 0.0172926f $X=0.79 $Y=0.49 $X2=0 $Y2=0
cc_245 Y N_A_216_55#_c_423_n 0.0140893f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_246 N_Y_M1001_d N_A_216_55#_c_428_n 0.00442863f $X=2.225 $Y=2.095 $X2=0 $Y2=0
cc_247 N_Y_c_339_n N_A_216_55#_c_428_n 0.0712841f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_248 N_Y_c_339_n N_A_216_55#_c_435_n 0.00849102f $X=2.2 $Y=2.55 $X2=0 $Y2=0
cc_249 Y N_A_216_55#_c_435_n 0.0136768f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_250 N_Y_c_331_n N_VGND_c_530_n 0.0114622f $X=0.295 $Y=0.49 $X2=0 $Y2=0
cc_251 N_Y_c_332_n N_VGND_c_530_n 0.037654f $X=0.79 $Y=0.49 $X2=0 $Y2=0
cc_252 N_Y_c_331_n N_VGND_c_532_n 0.00657784f $X=0.295 $Y=0.49 $X2=0 $Y2=0
cc_253 N_Y_c_332_n N_VGND_c_532_n 0.022179f $X=0.79 $Y=0.49 $X2=0 $Y2=0
cc_254 N_VPWR_c_375_n A_347_419# 0.00300148f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_255 N_VPWR_c_375_n A_559_419# 0.010279f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_256 N_VPWR_M1003_d N_A_216_55#_c_423_n 2.36033e-19 $X=1.1 $Y=2.095 $X2=0
+ $Y2=0
cc_257 N_VPWR_M1003_d N_A_216_55#_c_428_n 0.0083518f $X=1.1 $Y=2.095 $X2=0 $Y2=0
cc_258 N_VPWR_M1008_d N_A_216_55#_c_428_n 0.00587508f $X=3.285 $Y=2.095 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_377_n N_A_216_55#_c_428_n 0.0210602f $X=3.425 $Y=2.79 $X2=0
+ $Y2=0
cc_260 N_VPWR_M1003_d N_A_216_55#_c_435_n 7.61421e-19 $X=1.1 $Y=2.095 $X2=0
+ $Y2=0
cc_261 A_347_419# N_A_216_55#_c_428_n 0.00610645f $X=1.735 $Y=2.095 $X2=0.79
+ $Y2=0.49
cc_262 A_559_419# N_A_216_55#_c_428_n 0.00613492f $X=2.795 $Y=2.095 $X2=3.425
+ $Y2=2.79
cc_263 N_A_216_55#_c_422_n N_A_302_55#_c_480_n 0.015413f $X=1.22 $Y=0.49 $X2=0
+ $Y2=0
cc_264 N_A_216_55#_c_422_n N_A_302_55#_c_482_n 0.0132018f $X=1.22 $Y=0.49 $X2=0
+ $Y2=0
cc_265 N_A_216_55#_c_426_n N_A_302_55#_c_485_n 0.0172315f $X=4.1 $Y=0.49 $X2=0
+ $Y2=0
cc_266 N_A_216_55#_c_422_n N_VGND_c_530_n 0.0218883f $X=1.22 $Y=0.49 $X2=0 $Y2=0
cc_267 N_A_216_55#_c_426_n N_VGND_c_531_n 0.0308633f $X=4.1 $Y=0.49 $X2=0 $Y2=0
cc_268 N_A_216_55#_c_422_n N_VGND_c_532_n 0.0124575f $X=1.22 $Y=0.49 $X2=0 $Y2=0
cc_269 N_A_216_55#_c_426_n N_VGND_c_532_n 0.018168f $X=4.1 $Y=0.49 $X2=0 $Y2=0
cc_270 N_A_302_55#_c_481_n N_VGND_M1000_d 0.00681332f $X=2.585 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_271 N_A_302_55#_c_483_n N_VGND_M1000_d 0.00568386f $X=3.2 $Y=0.63 $X2=-0.19
+ $Y2=-0.245
cc_272 N_A_302_55#_c_484_n N_VGND_M1000_d 0.00675779f $X=2.67 $Y=0.63 $X2=-0.19
+ $Y2=-0.245
cc_273 N_A_302_55#_c_480_n N_VGND_c_529_n 0.00896155f $X=1.73 $Y=0.49 $X2=0
+ $Y2=0
cc_274 N_A_302_55#_c_481_n N_VGND_c_529_n 0.0240681f $X=2.585 $Y=0.77 $X2=0
+ $Y2=0
cc_275 N_A_302_55#_c_480_n N_VGND_c_530_n 0.0217987f $X=1.73 $Y=0.49 $X2=0 $Y2=0
cc_276 N_A_302_55#_c_481_n N_VGND_c_530_n 0.00228033f $X=2.585 $Y=0.77 $X2=0
+ $Y2=0
cc_277 N_A_302_55#_c_481_n N_VGND_c_531_n 0.00281466f $X=2.585 $Y=0.77 $X2=0
+ $Y2=0
cc_278 N_A_302_55#_c_483_n N_VGND_c_531_n 0.0089265f $X=3.2 $Y=0.63 $X2=0 $Y2=0
cc_279 N_A_302_55#_c_484_n N_VGND_c_531_n 0.0037773f $X=2.67 $Y=0.63 $X2=0 $Y2=0
cc_280 N_A_302_55#_c_485_n N_VGND_c_531_n 0.0212883f $X=3.365 $Y=0.49 $X2=0
+ $Y2=0
cc_281 N_A_302_55#_c_480_n N_VGND_c_532_n 0.0125322f $X=1.73 $Y=0.49 $X2=0 $Y2=0
cc_282 N_A_302_55#_c_481_n N_VGND_c_532_n 0.0107211f $X=2.585 $Y=0.77 $X2=0
+ $Y2=0
cc_283 N_A_302_55#_c_483_n N_VGND_c_532_n 0.0130074f $X=3.2 $Y=0.63 $X2=0 $Y2=0
cc_284 N_A_302_55#_c_484_n N_VGND_c_532_n 0.00526871f $X=2.67 $Y=0.63 $X2=0
+ $Y2=0
cc_285 N_A_302_55#_c_485_n N_VGND_c_532_n 0.0123326f $X=3.365 $Y=0.49 $X2=0
+ $Y2=0
