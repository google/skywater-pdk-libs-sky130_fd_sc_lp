* File: sky130_fd_sc_lp__dfxbp_2.pxi.spice
* Created: Fri Aug 28 10:23:49 2020
* 
x_PM_SKY130_FD_SC_LP__DFXBP_2%CLK N_CLK_M1008_g N_CLK_M1002_g N_CLK_c_193_n
+ N_CLK_c_194_n N_CLK_c_195_n CLK CLK CLK N_CLK_c_197_n
+ PM_SKY130_FD_SC_LP__DFXBP_2%CLK
x_PM_SKY130_FD_SC_LP__DFXBP_2%D N_D_M1024_g N_D_M1027_g N_D_c_221_n N_D_c_222_n
+ N_D_c_223_n D D D N_D_c_225_n PM_SKY130_FD_SC_LP__DFXBP_2%D
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_236_463# N_A_236_463#_M1028_s
+ N_A_236_463#_M1015_s N_A_236_463#_M1016_g N_A_236_463#_c_267_n
+ N_A_236_463#_M1000_g N_A_236_463#_M1025_g N_A_236_463#_c_261_n
+ N_A_236_463#_c_262_n N_A_236_463#_M1019_g N_A_236_463#_c_263_n
+ N_A_236_463#_c_272_n N_A_236_463#_c_273_n N_A_236_463#_c_274_n
+ N_A_236_463#_c_275_n N_A_236_463#_c_276_n N_A_236_463#_c_298_p
+ N_A_236_463#_c_277_n N_A_236_463#_c_264_n N_A_236_463#_c_279_n
+ N_A_236_463#_c_280_n N_A_236_463#_c_281_n N_A_236_463#_c_265_n
+ PM_SKY130_FD_SC_LP__DFXBP_2%A_236_463#
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_670_93# N_A_670_93#_M1022_d N_A_670_93#_M1009_d
+ N_A_670_93#_c_426_n N_A_670_93#_M1006_g N_A_670_93#_M1007_g
+ N_A_670_93#_c_427_n N_A_670_93#_c_436_n N_A_670_93#_c_428_n
+ N_A_670_93#_c_429_n N_A_670_93#_c_430_n N_A_670_93#_c_431_n
+ N_A_670_93#_c_432_n N_A_670_93#_c_433_n PM_SKY130_FD_SC_LP__DFXBP_2%A_670_93#
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_537_119# N_A_537_119#_M1001_d
+ N_A_537_119#_M1016_d N_A_537_119#_c_499_n N_A_537_119#_M1022_g
+ N_A_537_119#_M1009_g N_A_537_119#_c_500_n N_A_537_119#_c_506_n
+ N_A_537_119#_c_501_n N_A_537_119#_c_502_n N_A_537_119#_c_509_n
+ N_A_537_119#_c_503_n N_A_537_119#_c_504_n
+ PM_SKY130_FD_SC_LP__DFXBP_2%A_537_119#
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_110_70# N_A_110_70#_M1008_d N_A_110_70#_M1002_d
+ N_A_110_70#_c_575_n N_A_110_70#_c_576_n N_A_110_70#_M1015_g
+ N_A_110_70#_M1028_g N_A_110_70#_c_590_n N_A_110_70#_c_591_n
+ N_A_110_70#_c_579_n N_A_110_70#_c_580_n N_A_110_70#_M1001_g
+ N_A_110_70#_c_582_n N_A_110_70#_M1017_g N_A_110_70#_c_593_n
+ N_A_110_70#_M1023_g N_A_110_70#_M1026_g N_A_110_70#_c_584_n
+ N_A_110_70#_c_585_n N_A_110_70#_c_595_n N_A_110_70#_c_596_n
+ N_A_110_70#_c_597_n N_A_110_70#_c_586_n N_A_110_70#_c_587_n
+ N_A_110_70#_c_588_n PM_SKY130_FD_SC_LP__DFXBP_2%A_110_70#
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_1169_93# N_A_1169_93#_M1005_d
+ N_A_1169_93#_M1030_d N_A_1169_93#_c_708_n N_A_1169_93#_M1004_g
+ N_A_1169_93#_M1010_g N_A_1169_93#_c_709_n N_A_1169_93#_M1018_g
+ N_A_1169_93#_M1021_g N_A_1169_93#_M1003_g N_A_1169_93#_M1013_g
+ N_A_1169_93#_M1012_g N_A_1169_93#_M1014_g N_A_1169_93#_c_714_n
+ N_A_1169_93#_c_715_n N_A_1169_93#_c_716_n N_A_1169_93#_c_733_n
+ N_A_1169_93#_c_717_n N_A_1169_93#_c_743_n N_A_1169_93#_c_718_n
+ N_A_1169_93#_c_734_n N_A_1169_93#_c_735_n N_A_1169_93#_c_736_n
+ N_A_1169_93#_c_719_n N_A_1169_93#_c_720_n N_A_1169_93#_c_721_n
+ N_A_1169_93#_c_722_n N_A_1169_93#_c_738_n N_A_1169_93#_c_723_n
+ N_A_1169_93#_c_724_n N_A_1169_93#_c_725_n N_A_1169_93#_c_726_n
+ N_A_1169_93#_c_727_n PM_SKY130_FD_SC_LP__DFXBP_2%A_1169_93#
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_982_369# N_A_982_369#_M1025_d
+ N_A_982_369#_M1023_d N_A_982_369#_M1005_g N_A_982_369#_M1030_g
+ N_A_982_369#_c_873_n N_A_982_369#_c_874_n N_A_982_369#_c_875_n
+ N_A_982_369#_c_876_n N_A_982_369#_c_877_n N_A_982_369#_c_895_n
+ N_A_982_369#_c_878_n N_A_982_369#_c_879_n N_A_982_369#_c_880_n
+ PM_SKY130_FD_SC_LP__DFXBP_2%A_982_369#
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_1513_137# N_A_1513_137#_M1018_s
+ N_A_1513_137#_M1021_s N_A_1513_137#_c_962_n N_A_1513_137#_M1020_g
+ N_A_1513_137#_M1011_g N_A_1513_137#_c_964_n N_A_1513_137#_M1029_g
+ N_A_1513_137#_M1031_g N_A_1513_137#_c_966_n N_A_1513_137#_c_967_n
+ N_A_1513_137#_c_972_n N_A_1513_137#_c_968_n
+ PM_SKY130_FD_SC_LP__DFXBP_2%A_1513_137#
x_PM_SKY130_FD_SC_LP__DFXBP_2%VPWR N_VPWR_M1002_s N_VPWR_M1015_d N_VPWR_M1007_d
+ N_VPWR_M1010_d N_VPWR_M1021_d N_VPWR_M1031_d N_VPWR_M1012_s N_VPWR_c_1027_n
+ N_VPWR_c_1028_n N_VPWR_c_1029_n N_VPWR_c_1030_n N_VPWR_c_1031_n
+ N_VPWR_c_1032_n N_VPWR_c_1033_n N_VPWR_c_1034_n N_VPWR_c_1035_n
+ N_VPWR_c_1036_n N_VPWR_c_1037_n VPWR N_VPWR_c_1038_n N_VPWR_c_1039_n
+ N_VPWR_c_1040_n N_VPWR_c_1041_n N_VPWR_c_1042_n N_VPWR_c_1043_n
+ N_VPWR_c_1044_n N_VPWR_c_1045_n N_VPWR_c_1046_n N_VPWR_c_1026_n
+ PM_SKY130_FD_SC_LP__DFXBP_2%VPWR
x_PM_SKY130_FD_SC_LP__DFXBP_2%A_429_119# N_A_429_119#_M1024_d
+ N_A_429_119#_M1027_d N_A_429_119#_c_1140_n N_A_429_119#_c_1138_n
+ N_A_429_119#_c_1137_n PM_SKY130_FD_SC_LP__DFXBP_2%A_429_119#
x_PM_SKY130_FD_SC_LP__DFXBP_2%Q_N N_Q_N_M1020_d N_Q_N_M1011_s Q_N Q_N Q_N Q_N
+ Q_N N_Q_N_c_1165_n PM_SKY130_FD_SC_LP__DFXBP_2%Q_N
x_PM_SKY130_FD_SC_LP__DFXBP_2%Q N_Q_M1013_d N_Q_M1003_d N_Q_c_1183_n Q Q Q Q Q Q
+ Q N_Q_c_1185_n PM_SKY130_FD_SC_LP__DFXBP_2%Q
x_PM_SKY130_FD_SC_LP__DFXBP_2%VGND N_VGND_M1008_s N_VGND_M1028_d N_VGND_M1006_d
+ N_VGND_M1004_d N_VGND_M1018_d N_VGND_M1029_s N_VGND_M1014_s N_VGND_c_1205_n
+ N_VGND_c_1206_n N_VGND_c_1207_n N_VGND_c_1208_n N_VGND_c_1209_n
+ N_VGND_c_1210_n N_VGND_c_1211_n N_VGND_c_1212_n VGND N_VGND_c_1213_n
+ N_VGND_c_1214_n N_VGND_c_1215_n N_VGND_c_1216_n N_VGND_c_1217_n
+ N_VGND_c_1218_n N_VGND_c_1219_n N_VGND_c_1220_n N_VGND_c_1221_n
+ N_VGND_c_1222_n PM_SKY130_FD_SC_LP__DFXBP_2%VGND
cc_1 VNB N_CLK_M1002_g 0.00644914f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.61
cc_2 VNB N_CLK_c_193_n 0.0246852f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.88
cc_3 VNB N_CLK_c_194_n 0.0300413f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.385
cc_4 VNB N_CLK_c_195_n 0.0189125f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.55
cc_5 VNB CLK 0.0337136f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_CLK_c_197_n 0.019803f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_7 VNB N_D_c_221_n 0.0167562f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.88
cc_8 VNB N_D_c_222_n 0.0291574f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.385
cc_9 VNB N_D_c_223_n 0.00221227f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.55
cc_10 VNB D 0.00212036f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_11 VNB N_D_c_225_n 0.0188734f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_12 VNB N_A_236_463#_M1000_g 0.0452396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_236_463#_M1025_g 0.0208801f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_14 VNB N_A_236_463#_c_261_n 0.0210174f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.925
cc_15 VNB N_A_236_463#_c_262_n 0.0233173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_236_463#_c_263_n 0.0135758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_236_463#_c_264_n 0.00558902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_236_463#_c_265_n 0.0431095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_670_93#_c_426_n 0.0168672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_670_93#_c_427_n 0.0105403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_670_93#_c_428_n 0.00238816f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_22 VNB N_A_670_93#_c_429_n 0.00468056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_670_93#_c_430_n 0.00237791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_670_93#_c_431_n 2.53684e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_670_93#_c_432_n 0.00162017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_670_93#_c_433_n 0.0458833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_537_119#_c_499_n 0.0181199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_537_119#_c_500_n 0.004404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_537_119#_c_501_n 0.0127306f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_30 VNB N_A_537_119#_c_502_n 8.76593e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_537_119#_c_503_n 0.00244472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_537_119#_c_504_n 0.0341774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_110_70#_c_575_n 0.0211279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_110_70#_c_576_n 0.0195214f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_35 VNB N_A_110_70#_M1015_g 0.00401081f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_36 VNB N_A_110_70#_M1028_g 0.0481567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_110_70#_c_579_n 0.0593361f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_38 VNB N_A_110_70#_c_580_n 0.0126405f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_39 VNB N_A_110_70#_M1001_g 0.0404198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_110_70#_c_582_n 0.218613f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_41 VNB N_A_110_70#_M1026_g 0.0346662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_110_70#_c_584_n 0.0143406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_110_70#_c_585_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_110_70#_c_586_n 0.0158631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_110_70#_c_587_n 0.00531277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_110_70#_c_588_n 0.0119702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1169_93#_c_708_n 0.0180111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1169_93#_c_709_n 0.0319732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1169_93#_M1018_g 0.0260387f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.045
cc_50 VNB N_A_1169_93#_M1021_g 0.00871546f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.045
cc_51 VNB N_A_1169_93#_M1013_g 0.022661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1169_93#_M1014_g 0.0297671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1169_93#_c_714_n 0.0191009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1169_93#_c_715_n 0.00918414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1169_93#_c_716_n 0.00437251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1169_93#_c_717_n 0.00391059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1169_93#_c_718_n 0.016343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1169_93#_c_719_n 0.00581751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1169_93#_c_720_n 0.00276457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1169_93#_c_721_n 0.0193037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1169_93#_c_722_n 0.0248069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1169_93#_c_723_n 0.00308383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1169_93#_c_724_n 0.0441073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1169_93#_c_725_n 0.00308927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1169_93#_c_726_n 0.00183541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1169_93#_c_727_n 0.0711847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_982_369#_M1005_g 0.0242764f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.88
cc_68 VNB N_A_982_369#_c_873_n 0.0249015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_982_369#_c_874_n 3.74969e-19 $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.045
cc_70 VNB N_A_982_369#_c_875_n 0.00127379f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.045
cc_71 VNB N_A_982_369#_c_876_n 0.00210888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_982_369#_c_877_n 0.0268808f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_73 VNB N_A_982_369#_c_878_n 0.0011396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_982_369#_c_879_n 0.00102128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_982_369#_c_880_n 0.0167318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1513_137#_c_962_n 0.019115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1513_137#_M1011_g 0.00602303f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_78 VNB N_A_1513_137#_c_964_n 0.017407f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_79 VNB N_A_1513_137#_M1031_g 0.00499822f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.045
cc_80 VNB N_A_1513_137#_c_966_n 6.63573e-19 $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=1.045
cc_81 VNB N_A_1513_137#_c_967_n 0.0146077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1513_137#_c_968_n 0.0650667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VPWR_c_1026_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_429_119#_c_1137_n 0.00966395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_Q_c_1183_n 0.00132092f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.88
cc_86 VNB Q 0.00284409f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_87 VNB N_Q_c_1185_n 0.00189031f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_88 VNB N_VGND_c_1205_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1206_n 0.0216486f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.045
cc_90 VNB N_VGND_c_1207_n 0.00556671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1208_n 0.013088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1209_n 0.012341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1210_n 0.0513872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1211_n 0.0167433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1212_n 0.042272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1213_n 0.0326727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1214_n 0.0426277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1215_n 0.0468841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1216_n 0.0192204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1217_n 0.0179821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1218_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1219_n 0.0321229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1220_n 0.0100021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1221_n 0.0111602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1222_n 0.541316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VPB N_CLK_M1002_g 0.0638844f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.61
cc_107 VPB CLK 0.0102843f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_108 VPB N_D_M1027_g 0.0421262f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.61
cc_109 VPB N_D_c_223_n 0.0181729f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.55
cc_110 VPB D 0.00475698f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_111 VPB N_A_236_463#_M1016_g 0.0183981f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.88
cc_112 VPB N_A_236_463#_c_267_n 0.012166f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_113 VPB N_A_236_463#_M1000_g 0.0113352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_236_463#_c_262_n 0.00662927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_236_463#_M1019_g 0.0483364f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.295
cc_116 VPB N_A_236_463#_c_263_n 0.00549713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_236_463#_c_272_n 0.0150589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_236_463#_c_273_n 0.00249239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_236_463#_c_274_n 0.0202236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_236_463#_c_275_n 0.00136338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_236_463#_c_276_n 0.00949722f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_236_463#_c_277_n 0.00473113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_236_463#_c_264_n 0.00358934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_236_463#_c_279_n 0.0126606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_236_463#_c_280_n 0.0433659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_236_463#_c_281_n 0.0202603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_670_93#_M1007_g 0.0254434f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_128 VPB N_A_670_93#_c_427_n 0.0165484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_670_93#_c_436_n 0.0114584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_670_93#_c_429_n 5.57542e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_537_119#_M1009_g 0.0199458f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_132 VPB N_A_537_119#_c_506_n 0.0072139f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.045
cc_133 VPB N_A_537_119#_c_501_n 0.0081012f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.045
cc_134 VPB N_A_537_119#_c_502_n 0.00117194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_537_119#_c_509_n 0.00110606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_537_119#_c_503_n 0.00414724f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_537_119#_c_504_n 0.0114435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_110_70#_M1015_g 0.051364f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_139 VPB N_A_110_70#_c_590_n 0.110297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_110_70#_c_591_n 0.0126953f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.045
cc_141 VPB N_A_110_70#_M1017_g 0.0211864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_110_70#_c_593_n 0.114934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_110_70#_M1023_g 0.0459163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_110_70#_c_595_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_110_70#_c_596_n 0.0142436f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_110_70#_c_597_n 0.00987469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_110_70#_c_587_n 0.0473067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_1169_93#_M1010_g 0.0209859f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_149 VPB N_A_1169_93#_M1021_g 0.0262932f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.045
cc_150 VPB N_A_1169_93#_M1003_g 0.0217499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_1169_93#_M1012_g 0.0272177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_1169_93#_c_716_n 0.0195167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_1169_93#_c_733_n 0.0161488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_1169_93#_c_734_n 0.0107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_1169_93#_c_735_n 0.00789126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_1169_93#_c_736_n 0.0250353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_1169_93#_c_720_n 0.00752175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_1169_93#_c_738_n 0.00539079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_982_369#_M1030_g 0.0419815f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_160 VPB N_A_982_369#_c_874_n 0.0171076f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.045
cc_161 VPB N_A_982_369#_c_876_n 0.0109223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_982_369#_c_879_n 0.00168047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_1513_137#_M1011_g 0.0233713f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_164 VPB N_A_1513_137#_M1031_g 0.0210447f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.045
cc_165 VPB N_A_1513_137#_c_966_n 0.0039199f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.045
cc_166 VPB N_A_1513_137#_c_972_n 0.0152568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1027_n 0.0110658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1028_n 0.0416867f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.045
cc_169 VPB N_VPWR_c_1029_n 0.00159565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1030_n 0.0101028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1031_n 0.0151034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1032_n 0.0335075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1033_n 0.0129973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1034_n 0.0123785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1035_n 0.0654309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1036_n 0.0382142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1037_n 0.00814555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1038_n 0.0321999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1039_n 0.0511365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1040_n 0.0612483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1041_n 0.0182639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1042_n 0.0184107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1043_n 0.00330333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1044_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1045_n 0.00766811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1046_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1026_n 0.134266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_429_119#_c_1138_n 0.0028671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_429_119#_c_1137_n 0.00779519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB Q 0.00327718f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_191 N_CLK_M1002_g N_A_236_463#_c_263_n 3.91236e-19 $X=0.475 $Y=2.61 $X2=0
+ $Y2=0
cc_192 N_CLK_M1002_g N_A_236_463#_c_279_n 0.00123398f $X=0.475 $Y=2.61 $X2=0
+ $Y2=0
cc_193 N_CLK_c_195_n N_A_110_70#_c_576_n 0.0174403f $X=0.385 $Y=1.55 $X2=0 $Y2=0
cc_194 CLK N_A_110_70#_c_576_n 0.00126181f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_195 N_CLK_M1002_g N_A_110_70#_c_596_n 0.00835349f $X=0.475 $Y=2.61 $X2=0
+ $Y2=0
cc_196 N_CLK_M1002_g N_A_110_70#_c_597_n 0.00496861f $X=0.475 $Y=2.61 $X2=0
+ $Y2=0
cc_197 N_CLK_c_193_n N_A_110_70#_c_586_n 0.0166013f $X=0.385 $Y=0.88 $X2=0 $Y2=0
cc_198 N_CLK_c_195_n N_A_110_70#_c_586_n 0.00216729f $X=0.385 $Y=1.55 $X2=0
+ $Y2=0
cc_199 CLK N_A_110_70#_c_586_n 0.0450417f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_200 N_CLK_M1002_g N_A_110_70#_c_587_n 0.0174403f $X=0.475 $Y=2.61 $X2=0 $Y2=0
cc_201 N_CLK_c_193_n N_A_110_70#_c_588_n 6.25862e-19 $X=0.385 $Y=0.88 $X2=0
+ $Y2=0
cc_202 N_CLK_M1002_g N_VPWR_c_1028_n 0.0135641f $X=0.475 $Y=2.61 $X2=0 $Y2=0
cc_203 CLK N_VPWR_c_1028_n 0.0138645f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_204 N_CLK_M1002_g N_VPWR_c_1038_n 0.00536147f $X=0.475 $Y=2.61 $X2=0 $Y2=0
cc_205 N_CLK_M1002_g N_VPWR_c_1026_n 0.00521957f $X=0.475 $Y=2.61 $X2=0 $Y2=0
cc_206 N_CLK_c_193_n N_VGND_c_1206_n 0.0115229f $X=0.385 $Y=0.88 $X2=0 $Y2=0
cc_207 CLK N_VGND_c_1206_n 0.0266998f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_208 N_CLK_c_197_n N_VGND_c_1206_n 0.00110489f $X=0.385 $Y=1.045 $X2=0 $Y2=0
cc_209 N_CLK_c_193_n N_VGND_c_1213_n 0.00396895f $X=0.385 $Y=0.88 $X2=0 $Y2=0
cc_210 N_CLK_c_193_n N_VGND_c_1222_n 0.00662739f $X=0.385 $Y=0.88 $X2=0 $Y2=0
cc_211 CLK N_VGND_c_1222_n 0.00281011f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_212 N_D_M1027_g N_A_236_463#_c_267_n 0.02154f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_213 N_D_M1027_g N_A_236_463#_M1000_g 0.00186986f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_214 N_D_c_225_n N_A_236_463#_M1000_g 0.0067306f $X=2.16 $Y=1.29 $X2=0 $Y2=0
cc_215 N_D_M1027_g N_A_236_463#_c_263_n 0.0010281f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_216 N_D_c_222_n N_A_236_463#_c_263_n 0.00120439f $X=2.16 $Y=1.63 $X2=0 $Y2=0
cc_217 D N_A_236_463#_c_263_n 0.0312606f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_218 N_D_M1027_g N_A_236_463#_c_272_n 0.00528965f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_219 N_D_c_223_n N_A_236_463#_c_272_n 5.7175e-19 $X=2.16 $Y=1.795 $X2=0 $Y2=0
cc_220 D N_A_236_463#_c_272_n 0.0150634f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_221 N_D_M1027_g N_A_236_463#_c_273_n 0.0108324f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_222 N_D_M1027_g N_A_236_463#_c_274_n 0.00307819f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_223 N_D_M1027_g N_A_110_70#_M1015_g 0.016175f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_224 N_D_c_222_n N_A_110_70#_M1015_g 0.00582195f $X=2.16 $Y=1.63 $X2=0 $Y2=0
cc_225 D N_A_110_70#_M1015_g 0.00347857f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_226 N_D_c_221_n N_A_110_70#_M1028_g 0.0132366f $X=2.16 $Y=1.125 $X2=0 $Y2=0
cc_227 D N_A_110_70#_M1028_g 0.00191771f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_228 N_D_M1027_g N_A_110_70#_c_590_n 0.00897756f $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_229 N_D_c_221_n N_A_110_70#_c_579_n 0.0104164f $X=2.16 $Y=1.125 $X2=0 $Y2=0
cc_230 N_D_c_221_n N_A_110_70#_M1001_g 0.0123561f $X=2.16 $Y=1.125 $X2=0 $Y2=0
cc_231 N_D_c_225_n N_A_110_70#_M1001_g 0.00123393f $X=2.16 $Y=1.29 $X2=0 $Y2=0
cc_232 N_D_c_225_n N_A_110_70#_c_584_n 0.0132366f $X=2.16 $Y=1.29 $X2=0 $Y2=0
cc_233 N_D_M1027_g N_VPWR_c_1029_n 6.45389e-19 $X=2.22 $Y=2.525 $X2=0 $Y2=0
cc_234 D N_A_429_119#_c_1140_n 0.00521176f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_235 N_D_c_225_n N_A_429_119#_c_1140_n 0.00362353f $X=2.16 $Y=1.29 $X2=0 $Y2=0
cc_236 N_D_M1027_g N_A_429_119#_c_1137_n 0.00668021f $X=2.22 $Y=2.525 $X2=0
+ $Y2=0
cc_237 N_D_c_221_n N_A_429_119#_c_1137_n 0.00323441f $X=2.16 $Y=1.125 $X2=0
+ $Y2=0
cc_238 D N_A_429_119#_c_1137_n 0.0733272f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_239 N_D_c_225_n N_A_429_119#_c_1137_n 0.00784094f $X=2.16 $Y=1.29 $X2=0 $Y2=0
cc_240 N_D_c_221_n N_VGND_c_1207_n 0.0038173f $X=2.16 $Y=1.125 $X2=0 $Y2=0
cc_241 N_D_c_221_n N_VGND_c_1222_n 9.39239e-19 $X=2.16 $Y=1.125 $X2=0 $Y2=0
cc_242 N_A_236_463#_c_277_n N_A_670_93#_M1009_d 0.00537986f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_243 N_A_236_463#_M1000_g N_A_670_93#_c_426_n 0.0597399f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_244 N_A_236_463#_c_276_n N_A_670_93#_M1007_g 0.00432585f $X=3.39 $Y=2.405
+ $X2=0 $Y2=0
cc_245 N_A_236_463#_c_298_p N_A_670_93#_M1007_g 0.00585183f $X=3.39 $Y=2.905
+ $X2=0 $Y2=0
cc_246 N_A_236_463#_c_277_n N_A_670_93#_M1007_g 0.0151719f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_247 N_A_236_463#_c_280_n N_A_670_93#_M1007_g 0.00381934f $X=3.29 $Y=1.99
+ $X2=0 $Y2=0
cc_248 N_A_236_463#_M1000_g N_A_670_93#_c_427_n 0.0082442f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_249 N_A_236_463#_c_276_n N_A_670_93#_c_427_n 0.00407928f $X=3.39 $Y=2.405
+ $X2=0 $Y2=0
cc_250 N_A_236_463#_c_280_n N_A_670_93#_c_427_n 0.0158717f $X=3.29 $Y=1.99 $X2=0
+ $Y2=0
cc_251 N_A_236_463#_c_277_n N_A_670_93#_c_436_n 0.00121144f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_252 N_A_236_463#_c_277_n N_A_670_93#_c_429_n 0.0170777f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_253 N_A_236_463#_c_264_n N_A_670_93#_c_429_n 0.0599192f $X=5.05 $Y=1.34 $X2=0
+ $Y2=0
cc_254 N_A_236_463#_c_265_n N_A_670_93#_c_429_n 0.00331343f $X=5.215 $Y=1.34
+ $X2=0 $Y2=0
cc_255 N_A_236_463#_M1025_g N_A_670_93#_c_430_n 0.00524217f $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_256 N_A_236_463#_M1000_g N_A_670_93#_c_431_n 0.00101718f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_257 N_A_236_463#_M1025_g N_A_670_93#_c_432_n 0.00258989f $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_258 N_A_236_463#_c_280_n N_A_670_93#_c_433_n 0.00294089f $X=3.29 $Y=1.99
+ $X2=0 $Y2=0
cc_259 N_A_236_463#_c_274_n N_A_537_119#_M1016_d 0.00367596f $X=3.305 $Y=2.99
+ $X2=0 $Y2=0
cc_260 N_A_236_463#_M1025_g N_A_537_119#_c_499_n 0.00973929f $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_261 N_A_236_463#_c_264_n N_A_537_119#_c_499_n 2.09706e-19 $X=5.05 $Y=1.34
+ $X2=0 $Y2=0
cc_262 N_A_236_463#_c_277_n N_A_537_119#_M1009_g 0.0161016f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_263 N_A_236_463#_M1000_g N_A_537_119#_c_500_n 0.0234094f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_264 N_A_236_463#_M1016_g N_A_537_119#_c_506_n 0.00480121f $X=2.65 $Y=2.525
+ $X2=0 $Y2=0
cc_265 N_A_236_463#_M1000_g N_A_537_119#_c_506_n 0.00669536f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_266 N_A_236_463#_c_276_n N_A_537_119#_c_506_n 0.030248f $X=3.39 $Y=2.405
+ $X2=0 $Y2=0
cc_267 N_A_236_463#_c_281_n N_A_537_119#_c_506_n 0.0143033f $X=2.99 $Y=1.99
+ $X2=0 $Y2=0
cc_268 N_A_236_463#_M1000_g N_A_537_119#_c_501_n 0.0151764f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_269 N_A_236_463#_c_276_n N_A_537_119#_c_501_n 0.0269712f $X=3.39 $Y=2.405
+ $X2=0 $Y2=0
cc_270 N_A_236_463#_c_277_n N_A_537_119#_c_501_n 0.0181082f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_271 N_A_236_463#_c_280_n N_A_537_119#_c_501_n 0.00599042f $X=3.29 $Y=1.99
+ $X2=0 $Y2=0
cc_272 N_A_236_463#_M1000_g N_A_537_119#_c_502_n 0.00420066f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_273 N_A_236_463#_c_281_n N_A_537_119#_c_502_n 0.00162933f $X=2.99 $Y=1.99
+ $X2=0 $Y2=0
cc_274 N_A_236_463#_c_274_n N_A_537_119#_c_509_n 0.0253006f $X=3.305 $Y=2.99
+ $X2=0 $Y2=0
cc_275 N_A_236_463#_c_298_p N_A_537_119#_c_509_n 0.0236381f $X=3.39 $Y=2.905
+ $X2=0 $Y2=0
cc_276 N_A_236_463#_c_281_n N_A_537_119#_c_509_n 0.007746f $X=2.99 $Y=1.99 $X2=0
+ $Y2=0
cc_277 N_A_236_463#_c_277_n N_A_537_119#_c_503_n 0.00909937f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_278 N_A_236_463#_c_277_n N_A_537_119#_c_504_n 0.00127167f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_279 N_A_236_463#_c_264_n N_A_537_119#_c_504_n 8.13416e-19 $X=5.05 $Y=1.34
+ $X2=0 $Y2=0
cc_280 N_A_236_463#_c_265_n N_A_537_119#_c_504_n 0.00973929f $X=5.215 $Y=1.34
+ $X2=0 $Y2=0
cc_281 N_A_236_463#_c_263_n N_A_110_70#_c_575_n 0.014223f $X=1.38 $Y=0.805 $X2=0
+ $Y2=0
cc_282 N_A_236_463#_c_263_n N_A_110_70#_M1015_g 0.0228027f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_283 N_A_236_463#_c_272_n N_A_110_70#_M1015_g 0.0130125f $X=2 $Y=2.385 $X2=0
+ $Y2=0
cc_284 N_A_236_463#_c_273_n N_A_110_70#_M1015_g 0.00126741f $X=2.085 $Y=2.905
+ $X2=0 $Y2=0
cc_285 N_A_236_463#_c_275_n N_A_110_70#_M1015_g 6.62719e-19 $X=2.17 $Y=2.99
+ $X2=0 $Y2=0
cc_286 N_A_236_463#_c_279_n N_A_110_70#_M1015_g 0.00199203f $X=1.305 $Y=2.46
+ $X2=0 $Y2=0
cc_287 N_A_236_463#_c_263_n N_A_110_70#_M1028_g 0.0131946f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_288 N_A_236_463#_M1016_g N_A_110_70#_c_590_n 0.00882199f $X=2.65 $Y=2.525
+ $X2=0 $Y2=0
cc_289 N_A_236_463#_c_272_n N_A_110_70#_c_590_n 0.00414112f $X=2 $Y=2.385 $X2=0
+ $Y2=0
cc_290 N_A_236_463#_c_274_n N_A_110_70#_c_590_n 0.017362f $X=3.305 $Y=2.99 $X2=0
+ $Y2=0
cc_291 N_A_236_463#_c_275_n N_A_110_70#_c_590_n 0.00378523f $X=2.17 $Y=2.99
+ $X2=0 $Y2=0
cc_292 N_A_236_463#_M1000_g N_A_110_70#_M1001_g 0.0119936f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_293 N_A_236_463#_M1000_g N_A_110_70#_c_582_n 0.0103162f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_294 N_A_236_463#_M1025_g N_A_110_70#_c_582_n 0.0104164f $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_295 N_A_236_463#_M1016_g N_A_110_70#_M1017_g 0.00939635f $X=2.65 $Y=2.525
+ $X2=0 $Y2=0
cc_296 N_A_236_463#_c_274_n N_A_110_70#_M1017_g 0.014792f $X=3.305 $Y=2.99 $X2=0
+ $Y2=0
cc_297 N_A_236_463#_c_276_n N_A_110_70#_M1017_g 0.00242663f $X=3.39 $Y=2.405
+ $X2=0 $Y2=0
cc_298 N_A_236_463#_c_298_p N_A_110_70#_M1017_g 0.0128121f $X=3.39 $Y=2.905
+ $X2=0 $Y2=0
cc_299 N_A_236_463#_c_280_n N_A_110_70#_M1017_g 0.00994476f $X=3.29 $Y=1.99
+ $X2=0 $Y2=0
cc_300 N_A_236_463#_c_274_n N_A_110_70#_c_593_n 0.00206861f $X=3.305 $Y=2.99
+ $X2=0 $Y2=0
cc_301 N_A_236_463#_c_277_n N_A_110_70#_c_593_n 0.0104204f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_302 N_A_236_463#_c_277_n N_A_110_70#_M1023_g 0.0197751f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_303 N_A_236_463#_c_264_n N_A_110_70#_M1023_g 0.0104466f $X=5.05 $Y=1.34 $X2=0
+ $Y2=0
cc_304 N_A_236_463#_c_265_n N_A_110_70#_M1023_g 0.00459855f $X=5.215 $Y=1.34
+ $X2=0 $Y2=0
cc_305 N_A_236_463#_M1025_g N_A_110_70#_M1026_g 0.0149483f $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_306 N_A_236_463#_c_261_n N_A_110_70#_M1026_g 0.00953991f $X=5.485 $Y=1.43
+ $X2=0 $Y2=0
cc_307 N_A_236_463#_c_263_n N_A_110_70#_c_584_n 0.00369941f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_308 N_A_236_463#_c_274_n N_A_110_70#_c_595_n 3.42637e-19 $X=3.305 $Y=2.99
+ $X2=0 $Y2=0
cc_309 N_A_236_463#_c_263_n N_A_110_70#_c_596_n 0.00935191f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_310 N_A_236_463#_c_279_n N_A_110_70#_c_596_n 0.0377874f $X=1.305 $Y=2.46
+ $X2=0 $Y2=0
cc_311 N_A_236_463#_c_263_n N_A_110_70#_c_597_n 0.0131572f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_312 N_A_236_463#_c_263_n N_A_110_70#_c_586_n 0.0922999f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_313 N_A_236_463#_c_263_n N_A_110_70#_c_587_n 0.00428335f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_314 N_A_236_463#_c_263_n N_A_110_70#_c_588_n 0.00650832f $X=1.38 $Y=0.805
+ $X2=0 $Y2=0
cc_315 N_A_236_463#_M1019_g N_A_1169_93#_M1010_g 0.0230476f $X=5.71 $Y=2.475
+ $X2=0 $Y2=0
cc_316 N_A_236_463#_c_265_n N_A_1169_93#_c_714_n 0.0011781f $X=5.215 $Y=1.34
+ $X2=0 $Y2=0
cc_317 N_A_236_463#_c_262_n N_A_1169_93#_c_715_n 0.00647014f $X=5.71 $Y=1.665
+ $X2=0 $Y2=0
cc_318 N_A_236_463#_M1019_g N_A_1169_93#_c_716_n 0.0175495f $X=5.71 $Y=2.475
+ $X2=0 $Y2=0
cc_319 N_A_236_463#_c_262_n N_A_1169_93#_c_743_n 0.00177191f $X=5.71 $Y=1.665
+ $X2=0 $Y2=0
cc_320 N_A_236_463#_c_262_n N_A_1169_93#_c_718_n 0.0175495f $X=5.71 $Y=1.665
+ $X2=0 $Y2=0
cc_321 N_A_236_463#_M1019_g N_A_1169_93#_c_735_n 0.00111397f $X=5.71 $Y=2.475
+ $X2=0 $Y2=0
cc_322 N_A_236_463#_c_277_n N_A_982_369#_M1023_d 0.0101725f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_323 N_A_236_463#_c_264_n N_A_982_369#_M1023_d 0.00628409f $X=5.05 $Y=1.34
+ $X2=0 $Y2=0
cc_324 N_A_236_463#_M1025_g N_A_982_369#_c_875_n 0.00153486f $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_325 N_A_236_463#_c_261_n N_A_982_369#_c_876_n 0.011967f $X=5.485 $Y=1.43
+ $X2=0 $Y2=0
cc_326 N_A_236_463#_c_262_n N_A_982_369#_c_876_n 0.0126038f $X=5.71 $Y=1.665
+ $X2=0 $Y2=0
cc_327 N_A_236_463#_M1019_g N_A_982_369#_c_876_n 0.0343008f $X=5.71 $Y=2.475
+ $X2=0 $Y2=0
cc_328 N_A_236_463#_c_277_n N_A_982_369#_c_876_n 0.0141997f $X=4.955 $Y=2.32
+ $X2=0 $Y2=0
cc_329 N_A_236_463#_c_264_n N_A_982_369#_c_876_n 0.0694623f $X=5.05 $Y=1.34
+ $X2=0 $Y2=0
cc_330 N_A_236_463#_c_265_n N_A_982_369#_c_876_n 9.98304e-19 $X=5.215 $Y=1.34
+ $X2=0 $Y2=0
cc_331 N_A_236_463#_c_262_n N_A_982_369#_c_877_n 0.00787426f $X=5.71 $Y=1.665
+ $X2=0 $Y2=0
cc_332 N_A_236_463#_M1025_g N_A_982_369#_c_895_n 0.00395845f $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_333 N_A_236_463#_c_261_n N_A_982_369#_c_895_n 0.00348696f $X=5.485 $Y=1.43
+ $X2=0 $Y2=0
cc_334 N_A_236_463#_c_264_n N_A_982_369#_c_895_n 0.0050179f $X=5.05 $Y=1.34
+ $X2=0 $Y2=0
cc_335 N_A_236_463#_c_265_n N_A_982_369#_c_895_n 0.0032813f $X=5.215 $Y=1.34
+ $X2=0 $Y2=0
cc_336 N_A_236_463#_M1025_g N_A_982_369#_c_878_n 6.14431e-19 $X=4.93 $Y=0.805
+ $X2=0 $Y2=0
cc_337 N_A_236_463#_c_264_n N_A_982_369#_c_878_n 0.0113769f $X=5.05 $Y=1.34
+ $X2=0 $Y2=0
cc_338 N_A_236_463#_c_265_n N_A_982_369#_c_878_n 0.00230333f $X=5.215 $Y=1.34
+ $X2=0 $Y2=0
cc_339 N_A_236_463#_c_272_n N_VPWR_M1015_d 0.0048841f $X=2 $Y=2.385 $X2=0 $Y2=0
cc_340 N_A_236_463#_c_273_n N_VPWR_M1015_d 0.00336363f $X=2.085 $Y=2.905 $X2=0
+ $Y2=0
cc_341 N_A_236_463#_c_277_n N_VPWR_M1007_d 0.00986464f $X=4.955 $Y=2.32 $X2=0
+ $Y2=0
cc_342 N_A_236_463#_c_272_n N_VPWR_c_1029_n 0.015111f $X=2 $Y=2.385 $X2=0 $Y2=0
cc_343 N_A_236_463#_c_273_n N_VPWR_c_1029_n 0.0200088f $X=2.085 $Y=2.905 $X2=0
+ $Y2=0
cc_344 N_A_236_463#_c_275_n N_VPWR_c_1029_n 0.0146734f $X=2.17 $Y=2.99 $X2=0
+ $Y2=0
cc_345 N_A_236_463#_c_279_n N_VPWR_c_1029_n 0.0120501f $X=1.305 $Y=2.46 $X2=0
+ $Y2=0
cc_346 N_A_236_463#_c_274_n N_VPWR_c_1030_n 0.00740565f $X=3.305 $Y=2.99 $X2=0
+ $Y2=0
cc_347 N_A_236_463#_c_298_p N_VPWR_c_1030_n 0.0121244f $X=3.39 $Y=2.905 $X2=0
+ $Y2=0
cc_348 N_A_236_463#_c_277_n N_VPWR_c_1030_n 0.0266042f $X=4.955 $Y=2.32 $X2=0
+ $Y2=0
cc_349 N_A_236_463#_M1019_g N_VPWR_c_1031_n 0.00247929f $X=5.71 $Y=2.475 $X2=0
+ $Y2=0
cc_350 N_A_236_463#_c_279_n N_VPWR_c_1038_n 0.0112754f $X=1.305 $Y=2.46 $X2=0
+ $Y2=0
cc_351 N_A_236_463#_c_274_n N_VPWR_c_1039_n 0.0842755f $X=3.305 $Y=2.99 $X2=0
+ $Y2=0
cc_352 N_A_236_463#_c_275_n N_VPWR_c_1039_n 0.0115893f $X=2.17 $Y=2.99 $X2=0
+ $Y2=0
cc_353 N_A_236_463#_M1019_g N_VPWR_c_1040_n 0.00404937f $X=5.71 $Y=2.475 $X2=0
+ $Y2=0
cc_354 N_A_236_463#_M1019_g N_VPWR_c_1026_n 0.0046394f $X=5.71 $Y=2.475 $X2=0
+ $Y2=0
cc_355 N_A_236_463#_c_272_n N_VPWR_c_1026_n 0.00874693f $X=2 $Y=2.385 $X2=0
+ $Y2=0
cc_356 N_A_236_463#_c_274_n N_VPWR_c_1026_n 0.0438485f $X=3.305 $Y=2.99 $X2=0
+ $Y2=0
cc_357 N_A_236_463#_c_275_n N_VPWR_c_1026_n 0.00583135f $X=2.17 $Y=2.99 $X2=0
+ $Y2=0
cc_358 N_A_236_463#_c_279_n N_VPWR_c_1026_n 0.0120432f $X=1.305 $Y=2.46 $X2=0
+ $Y2=0
cc_359 N_A_236_463#_M1016_g N_A_429_119#_c_1138_n 0.00366715f $X=2.65 $Y=2.525
+ $X2=0 $Y2=0
cc_360 N_A_236_463#_c_272_n N_A_429_119#_c_1138_n 0.00737527f $X=2 $Y=2.385
+ $X2=0 $Y2=0
cc_361 N_A_236_463#_c_274_n N_A_429_119#_c_1138_n 0.0108977f $X=3.305 $Y=2.99
+ $X2=0 $Y2=0
cc_362 N_A_236_463#_M1016_g N_A_429_119#_c_1137_n 0.00254542f $X=2.65 $Y=2.525
+ $X2=0 $Y2=0
cc_363 N_A_236_463#_c_267_n N_A_429_119#_c_1137_n 0.00390877f $X=2.725 $Y=2.08
+ $X2=0 $Y2=0
cc_364 N_A_236_463#_M1000_g N_A_429_119#_c_1137_n 0.00153455f $X=3.065 $Y=0.805
+ $X2=0 $Y2=0
cc_365 N_A_236_463#_c_298_p A_669_499# 0.00653665f $X=3.39 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_366 N_A_236_463#_c_277_n A_669_499# 0.00304701f $X=4.955 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_367 N_A_236_463#_c_263_n N_VGND_c_1213_n 0.00485468f $X=1.38 $Y=0.805 $X2=0
+ $Y2=0
cc_368 N_A_236_463#_M1000_g N_VGND_c_1219_n 0.00139459f $X=3.065 $Y=0.805 $X2=0
+ $Y2=0
cc_369 N_A_236_463#_M1025_g N_VGND_c_1219_n 6.09261e-19 $X=4.93 $Y=0.805 $X2=0
+ $Y2=0
cc_370 N_A_236_463#_M1000_g N_VGND_c_1222_n 9.39239e-19 $X=3.065 $Y=0.805 $X2=0
+ $Y2=0
cc_371 N_A_236_463#_M1025_g N_VGND_c_1222_n 9.39239e-19 $X=4.93 $Y=0.805 $X2=0
+ $Y2=0
cc_372 N_A_236_463#_c_263_n N_VGND_c_1222_n 0.00780059f $X=1.38 $Y=0.805 $X2=0
+ $Y2=0
cc_373 N_A_670_93#_c_428_n N_A_537_119#_c_499_n 0.0155503f $X=4.455 $Y=1.09
+ $X2=0 $Y2=0
cc_374 N_A_670_93#_c_429_n N_A_537_119#_c_499_n 0.00510561f $X=4.62 $Y=1.97
+ $X2=0 $Y2=0
cc_375 N_A_670_93#_c_431_n N_A_537_119#_c_499_n 9.81335e-19 $X=3.65 $Y=1.09
+ $X2=0 $Y2=0
cc_376 N_A_670_93#_c_432_n N_A_537_119#_c_499_n 0.00156298f $X=4.62 $Y=1.09
+ $X2=0 $Y2=0
cc_377 N_A_670_93#_c_433_n N_A_537_119#_c_499_n 0.00465836f $X=3.74 $Y=1.29
+ $X2=0 $Y2=0
cc_378 N_A_670_93#_c_427_n N_A_537_119#_M1009_g 0.00550493f $X=3.76 $Y=1.925
+ $X2=0 $Y2=0
cc_379 N_A_670_93#_c_436_n N_A_537_119#_M1009_g 0.0217958f $X=3.76 $Y=2.075
+ $X2=0 $Y2=0
cc_380 N_A_670_93#_c_429_n N_A_537_119#_M1009_g 0.0101619f $X=4.62 $Y=1.97 $X2=0
+ $Y2=0
cc_381 N_A_670_93#_c_426_n N_A_537_119#_c_500_n 0.00296414f $X=3.425 $Y=1.125
+ $X2=0 $Y2=0
cc_382 N_A_670_93#_c_427_n N_A_537_119#_c_500_n 4.27344e-19 $X=3.76 $Y=1.925
+ $X2=0 $Y2=0
cc_383 N_A_670_93#_c_431_n N_A_537_119#_c_500_n 0.0122044f $X=3.65 $Y=1.09 $X2=0
+ $Y2=0
cc_384 N_A_670_93#_c_427_n N_A_537_119#_c_501_n 0.0127034f $X=3.76 $Y=1.925
+ $X2=0 $Y2=0
cc_385 N_A_670_93#_c_436_n N_A_537_119#_c_501_n 0.00115332f $X=3.76 $Y=2.075
+ $X2=0 $Y2=0
cc_386 N_A_670_93#_c_428_n N_A_537_119#_c_501_n 0.00901096f $X=4.455 $Y=1.09
+ $X2=0 $Y2=0
cc_387 N_A_670_93#_c_431_n N_A_537_119#_c_501_n 0.0244829f $X=3.65 $Y=1.09 $X2=0
+ $Y2=0
cc_388 N_A_670_93#_c_433_n N_A_537_119#_c_501_n 0.00850401f $X=3.74 $Y=1.29
+ $X2=0 $Y2=0
cc_389 N_A_670_93#_c_428_n N_A_537_119#_c_503_n 0.0180925f $X=4.455 $Y=1.09
+ $X2=0 $Y2=0
cc_390 N_A_670_93#_c_429_n N_A_537_119#_c_503_n 0.0273892f $X=4.62 $Y=1.97 $X2=0
+ $Y2=0
cc_391 N_A_670_93#_c_431_n N_A_537_119#_c_503_n 0.00186711f $X=3.65 $Y=1.09
+ $X2=0 $Y2=0
cc_392 N_A_670_93#_c_433_n N_A_537_119#_c_503_n 0.00130265f $X=3.74 $Y=1.29
+ $X2=0 $Y2=0
cc_393 N_A_670_93#_c_428_n N_A_537_119#_c_504_n 0.00177146f $X=4.455 $Y=1.09
+ $X2=0 $Y2=0
cc_394 N_A_670_93#_c_429_n N_A_537_119#_c_504_n 0.0107738f $X=4.62 $Y=1.97 $X2=0
+ $Y2=0
cc_395 N_A_670_93#_c_433_n N_A_537_119#_c_504_n 0.0218931f $X=3.74 $Y=1.29 $X2=0
+ $Y2=0
cc_396 N_A_670_93#_c_426_n N_A_110_70#_c_582_n 0.0103107f $X=3.425 $Y=1.125
+ $X2=0 $Y2=0
cc_397 N_A_670_93#_c_430_n N_A_110_70#_c_582_n 0.00520087f $X=4.62 $Y=0.75 $X2=0
+ $Y2=0
cc_398 N_A_670_93#_M1007_g N_A_110_70#_M1017_g 0.0146656f $X=3.78 $Y=2.525 $X2=0
+ $Y2=0
cc_399 N_A_670_93#_M1007_g N_A_110_70#_c_593_n 0.0101316f $X=3.78 $Y=2.525 $X2=0
+ $Y2=0
cc_400 N_A_670_93#_c_429_n N_A_110_70#_M1023_g 0.0061824f $X=4.62 $Y=1.97 $X2=0
+ $Y2=0
cc_401 N_A_670_93#_c_430_n N_A_982_369#_c_875_n 9.75027e-19 $X=4.62 $Y=0.75
+ $X2=0 $Y2=0
cc_402 N_A_670_93#_c_432_n N_A_982_369#_c_875_n 0.00541131f $X=4.62 $Y=1.09
+ $X2=0 $Y2=0
cc_403 N_A_670_93#_c_430_n N_A_982_369#_c_895_n 0.0183071f $X=4.62 $Y=0.75 $X2=0
+ $Y2=0
cc_404 N_A_670_93#_c_432_n N_A_982_369#_c_878_n 0.00126132f $X=4.62 $Y=1.09
+ $X2=0 $Y2=0
cc_405 N_A_670_93#_M1007_g N_VPWR_c_1030_n 0.00451394f $X=3.78 $Y=2.525 $X2=0
+ $Y2=0
cc_406 N_A_670_93#_M1007_g N_VPWR_c_1026_n 9.39239e-19 $X=3.78 $Y=2.525 $X2=0
+ $Y2=0
cc_407 N_A_670_93#_c_428_n N_VGND_M1006_d 0.00908184f $X=4.455 $Y=1.09 $X2=0
+ $Y2=0
cc_408 N_A_670_93#_c_431_n N_VGND_M1006_d 0.00281835f $X=3.65 $Y=1.09 $X2=0
+ $Y2=0
cc_409 N_A_670_93#_c_430_n N_VGND_c_1215_n 0.00580769f $X=4.62 $Y=0.75 $X2=0
+ $Y2=0
cc_410 N_A_670_93#_c_426_n N_VGND_c_1219_n 0.0103896f $X=3.425 $Y=1.125 $X2=0
+ $Y2=0
cc_411 N_A_670_93#_c_428_n N_VGND_c_1219_n 0.0390483f $X=4.455 $Y=1.09 $X2=0
+ $Y2=0
cc_412 N_A_670_93#_c_430_n N_VGND_c_1219_n 0.0108424f $X=4.62 $Y=0.75 $X2=0
+ $Y2=0
cc_413 N_A_670_93#_c_431_n N_VGND_c_1219_n 0.023306f $X=3.65 $Y=1.09 $X2=0 $Y2=0
cc_414 N_A_670_93#_c_433_n N_VGND_c_1219_n 0.00170059f $X=3.74 $Y=1.29 $X2=0
+ $Y2=0
cc_415 N_A_670_93#_c_426_n N_VGND_c_1222_n 7.88961e-19 $X=3.425 $Y=1.125 $X2=0
+ $Y2=0
cc_416 N_A_670_93#_c_430_n N_VGND_c_1222_n 0.00710006f $X=4.62 $Y=0.75 $X2=0
+ $Y2=0
cc_417 N_A_537_119#_c_500_n N_A_110_70#_M1001_g 0.00209302f $X=2.85 $Y=0.805
+ $X2=0 $Y2=0
cc_418 N_A_537_119#_c_499_n N_A_110_70#_c_582_n 0.0103107f $X=4.405 $Y=1.355
+ $X2=0 $Y2=0
cc_419 N_A_537_119#_c_500_n N_A_110_70#_c_582_n 0.00387959f $X=2.85 $Y=0.805
+ $X2=0 $Y2=0
cc_420 N_A_537_119#_c_506_n N_A_110_70#_M1017_g 3.29355e-19 $X=2.855 $Y=2.405
+ $X2=0 $Y2=0
cc_421 N_A_537_119#_c_509_n N_A_110_70#_M1017_g 0.00318518f $X=2.96 $Y=2.57
+ $X2=0 $Y2=0
cc_422 N_A_537_119#_M1009_g N_A_110_70#_c_593_n 0.00794568f $X=4.405 $Y=2.265
+ $X2=0 $Y2=0
cc_423 N_A_537_119#_M1009_g N_A_110_70#_M1023_g 0.0365182f $X=4.405 $Y=2.265
+ $X2=0 $Y2=0
cc_424 N_A_537_119#_M1009_g N_VPWR_c_1030_n 0.00453309f $X=4.405 $Y=2.265 $X2=0
+ $Y2=0
cc_425 N_A_537_119#_M1009_g N_VPWR_c_1026_n 9.55878e-19 $X=4.405 $Y=2.265 $X2=0
+ $Y2=0
cc_426 N_A_537_119#_c_500_n N_A_429_119#_c_1140_n 0.0244033f $X=2.85 $Y=0.805
+ $X2=0 $Y2=0
cc_427 N_A_537_119#_c_500_n N_A_429_119#_c_1137_n 0.0456969f $X=2.85 $Y=0.805
+ $X2=0 $Y2=0
cc_428 N_A_537_119#_c_506_n N_A_429_119#_c_1137_n 0.0459942f $X=2.855 $Y=2.405
+ $X2=0 $Y2=0
cc_429 N_A_537_119#_c_502_n N_A_429_119#_c_1137_n 0.0143577f $X=2.89 $Y=1.64
+ $X2=0 $Y2=0
cc_430 N_A_537_119#_c_500_n N_VGND_c_1214_n 0.00415173f $X=2.85 $Y=0.805 $X2=0
+ $Y2=0
cc_431 N_A_537_119#_c_499_n N_VGND_c_1219_n 0.00878485f $X=4.405 $Y=1.355 $X2=0
+ $Y2=0
cc_432 N_A_537_119#_c_500_n N_VGND_c_1219_n 0.00677107f $X=2.85 $Y=0.805 $X2=0
+ $Y2=0
cc_433 N_A_537_119#_c_499_n N_VGND_c_1222_n 7.88961e-19 $X=4.405 $Y=1.355 $X2=0
+ $Y2=0
cc_434 N_A_537_119#_c_500_n N_VGND_c_1222_n 0.00648087f $X=2.85 $Y=0.805 $X2=0
+ $Y2=0
cc_435 N_A_110_70#_M1026_g N_A_1169_93#_c_708_n 0.0378272f $X=5.55 $Y=0.805
+ $X2=0 $Y2=0
cc_436 N_A_110_70#_M1026_g N_A_982_369#_c_875_n 0.00591586f $X=5.55 $Y=0.805
+ $X2=0 $Y2=0
cc_437 N_A_110_70#_M1023_g N_A_982_369#_c_876_n 0.00993905f $X=4.835 $Y=2.265
+ $X2=0 $Y2=0
cc_438 N_A_110_70#_M1026_g N_A_982_369#_c_877_n 0.00154629f $X=5.55 $Y=0.805
+ $X2=0 $Y2=0
cc_439 N_A_110_70#_c_582_n N_A_982_369#_c_895_n 0.00568984f $X=5.475 $Y=0.18
+ $X2=0 $Y2=0
cc_440 N_A_110_70#_M1026_g N_A_982_369#_c_895_n 0.0139659f $X=5.55 $Y=0.805
+ $X2=0 $Y2=0
cc_441 N_A_110_70#_M1026_g N_A_982_369#_c_878_n 8.26078e-19 $X=5.55 $Y=0.805
+ $X2=0 $Y2=0
cc_442 N_A_110_70#_c_596_n N_VPWR_c_1028_n 0.0260368f $X=0.69 $Y=2.445 $X2=0
+ $Y2=0
cc_443 N_A_110_70#_M1015_g N_VPWR_c_1029_n 0.0101741f $X=1.52 $Y=2.635 $X2=0
+ $Y2=0
cc_444 N_A_110_70#_c_590_n N_VPWR_c_1029_n 0.0145012f $X=3.195 $Y=3.15 $X2=0
+ $Y2=0
cc_445 N_A_110_70#_c_591_n N_VPWR_c_1029_n 0.0035753f $X=1.595 $Y=3.15 $X2=0
+ $Y2=0
cc_446 N_A_110_70#_M1017_g N_VPWR_c_1030_n 0.00114631f $X=3.27 $Y=2.705 $X2=0
+ $Y2=0
cc_447 N_A_110_70#_c_593_n N_VPWR_c_1030_n 0.025556f $X=4.76 $Y=3.15 $X2=0 $Y2=0
cc_448 N_A_110_70#_M1023_g N_VPWR_c_1030_n 0.00736786f $X=4.835 $Y=2.265 $X2=0
+ $Y2=0
cc_449 N_A_110_70#_c_591_n N_VPWR_c_1038_n 0.00525069f $X=1.595 $Y=3.15 $X2=0
+ $Y2=0
cc_450 N_A_110_70#_c_596_n N_VPWR_c_1038_n 0.0110688f $X=0.69 $Y=2.445 $X2=0
+ $Y2=0
cc_451 N_A_110_70#_c_590_n N_VPWR_c_1039_n 0.0534324f $X=3.195 $Y=3.15 $X2=0
+ $Y2=0
cc_452 N_A_110_70#_c_593_n N_VPWR_c_1040_n 0.0232701f $X=4.76 $Y=3.15 $X2=0
+ $Y2=0
cc_453 N_A_110_70#_c_590_n N_VPWR_c_1026_n 0.0327646f $X=3.195 $Y=3.15 $X2=0
+ $Y2=0
cc_454 N_A_110_70#_c_591_n N_VPWR_c_1026_n 0.00646524f $X=1.595 $Y=3.15 $X2=0
+ $Y2=0
cc_455 N_A_110_70#_c_593_n N_VPWR_c_1026_n 0.0604531f $X=4.76 $Y=3.15 $X2=0
+ $Y2=0
cc_456 N_A_110_70#_c_595_n N_VPWR_c_1026_n 0.00370843f $X=3.27 $Y=3.15 $X2=0
+ $Y2=0
cc_457 N_A_110_70#_c_596_n N_VPWR_c_1026_n 0.0100797f $X=0.69 $Y=2.445 $X2=0
+ $Y2=0
cc_458 N_A_110_70#_c_579_n N_A_429_119#_c_1140_n 0.00481166f $X=2.535 $Y=0.18
+ $X2=0 $Y2=0
cc_459 N_A_110_70#_M1001_g N_A_429_119#_c_1140_n 0.00576121f $X=2.61 $Y=0.805
+ $X2=0 $Y2=0
cc_460 N_A_110_70#_M1001_g N_A_429_119#_c_1137_n 0.00523045f $X=2.61 $Y=0.805
+ $X2=0 $Y2=0
cc_461 N_A_110_70#_c_588_n N_VGND_c_1206_n 0.0135678f $X=0.915 $Y=0.525 $X2=0
+ $Y2=0
cc_462 N_A_110_70#_M1028_g N_VGND_c_1207_n 0.020159f $X=1.595 $Y=0.805 $X2=0
+ $Y2=0
cc_463 N_A_110_70#_c_579_n N_VGND_c_1207_n 0.0187123f $X=2.535 $Y=0.18 $X2=0
+ $Y2=0
cc_464 N_A_110_70#_c_580_n N_VGND_c_1207_n 0.00388727f $X=1.67 $Y=0.18 $X2=0
+ $Y2=0
cc_465 N_A_110_70#_M1001_g N_VGND_c_1207_n 0.00550178f $X=2.61 $Y=0.805 $X2=0
+ $Y2=0
cc_466 N_A_110_70#_c_588_n N_VGND_c_1207_n 0.00962588f $X=0.915 $Y=0.525 $X2=0
+ $Y2=0
cc_467 N_A_110_70#_c_582_n N_VGND_c_1208_n 0.010516f $X=5.475 $Y=0.18 $X2=0
+ $Y2=0
cc_468 N_A_110_70#_M1026_g N_VGND_c_1208_n 0.00176088f $X=5.55 $Y=0.805 $X2=0
+ $Y2=0
cc_469 N_A_110_70#_c_580_n N_VGND_c_1213_n 0.00486043f $X=1.67 $Y=0.18 $X2=0
+ $Y2=0
cc_470 N_A_110_70#_c_588_n N_VGND_c_1213_n 0.0206407f $X=0.915 $Y=0.525 $X2=0
+ $Y2=0
cc_471 N_A_110_70#_c_579_n N_VGND_c_1214_n 0.0470016f $X=2.535 $Y=0.18 $X2=0
+ $Y2=0
cc_472 N_A_110_70#_c_582_n N_VGND_c_1215_n 0.0376009f $X=5.475 $Y=0.18 $X2=0
+ $Y2=0
cc_473 N_A_110_70#_c_582_n N_VGND_c_1219_n 0.0557164f $X=5.475 $Y=0.18 $X2=0
+ $Y2=0
cc_474 N_A_110_70#_c_579_n N_VGND_c_1222_n 0.0172617f $X=2.535 $Y=0.18 $X2=0
+ $Y2=0
cc_475 N_A_110_70#_c_580_n N_VGND_c_1222_n 0.00983503f $X=1.67 $Y=0.18 $X2=0
+ $Y2=0
cc_476 N_A_110_70#_c_582_n N_VGND_c_1222_n 0.0761814f $X=5.475 $Y=0.18 $X2=0
+ $Y2=0
cc_477 N_A_110_70#_c_585_n N_VGND_c_1222_n 0.00727527f $X=2.61 $Y=0.18 $X2=0
+ $Y2=0
cc_478 N_A_110_70#_c_588_n N_VGND_c_1222_n 0.0163302f $X=0.915 $Y=0.525 $X2=0
+ $Y2=0
cc_479 N_A_1169_93#_c_708_n N_A_982_369#_M1005_g 0.00691713f $X=5.92 $Y=1.125
+ $X2=0 $Y2=0
cc_480 N_A_1169_93#_c_714_n N_A_982_369#_M1005_g 0.00469429f $X=6.07 $Y=1.2
+ $X2=0 $Y2=0
cc_481 N_A_1169_93#_c_719_n N_A_982_369#_M1005_g 0.00454254f $X=7.05 $Y=1.255
+ $X2=0 $Y2=0
cc_482 N_A_1169_93#_c_722_n N_A_982_369#_M1005_g 0.00748575f $X=6.825 $Y=0.52
+ $X2=0 $Y2=0
cc_483 N_A_1169_93#_M1010_g N_A_982_369#_M1030_g 0.013388f $X=6.22 $Y=2.465
+ $X2=0 $Y2=0
cc_484 N_A_1169_93#_c_716_n N_A_982_369#_M1030_g 0.00809514f $X=6.16 $Y=1.93
+ $X2=0 $Y2=0
cc_485 N_A_1169_93#_c_743_n N_A_982_369#_M1030_g 6.64418e-19 $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_486 N_A_1169_93#_c_734_n N_A_982_369#_M1030_g 0.0193288f $X=6.9 $Y=2.075
+ $X2=0 $Y2=0
cc_487 N_A_1169_93#_c_736_n N_A_982_369#_M1030_g 0.00607936f $X=7.005 $Y=2.4
+ $X2=0 $Y2=0
cc_488 N_A_1169_93#_c_743_n N_A_982_369#_c_873_n 0.00107622f $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_489 N_A_1169_93#_c_718_n N_A_982_369#_c_873_n 0.0121203f $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_490 N_A_1169_93#_c_720_n N_A_982_369#_c_873_n 0.0117806f $X=7.067 $Y=1.985
+ $X2=0 $Y2=0
cc_491 N_A_1169_93#_c_716_n N_A_982_369#_c_874_n 0.0121203f $X=6.16 $Y=1.93
+ $X2=0 $Y2=0
cc_492 N_A_1169_93#_c_734_n N_A_982_369#_c_874_n 0.00125045f $X=6.9 $Y=2.075
+ $X2=0 $Y2=0
cc_493 N_A_1169_93#_c_708_n N_A_982_369#_c_875_n 9.80256e-19 $X=5.92 $Y=1.125
+ $X2=0 $Y2=0
cc_494 N_A_1169_93#_c_715_n N_A_982_369#_c_876_n 0.00230655f $X=6.16 $Y=1.425
+ $X2=0 $Y2=0
cc_495 N_A_1169_93#_c_743_n N_A_982_369#_c_876_n 0.0178487f $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_496 N_A_1169_93#_c_735_n N_A_982_369#_c_876_n 0.00765521f $X=6.325 $Y=2.075
+ $X2=0 $Y2=0
cc_497 N_A_1169_93#_c_714_n N_A_982_369#_c_877_n 0.0170757f $X=6.07 $Y=1.2 $X2=0
+ $Y2=0
cc_498 N_A_1169_93#_c_715_n N_A_982_369#_c_877_n 0.00416367f $X=6.16 $Y=1.425
+ $X2=0 $Y2=0
cc_499 N_A_1169_93#_c_743_n N_A_982_369#_c_877_n 0.0234645f $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_500 N_A_1169_93#_c_718_n N_A_982_369#_c_877_n 0.00513735f $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_501 N_A_1169_93#_c_734_n N_A_982_369#_c_877_n 0.0060642f $X=6.9 $Y=2.075
+ $X2=0 $Y2=0
cc_502 N_A_1169_93#_c_708_n N_A_982_369#_c_895_n 0.00101961f $X=5.92 $Y=1.125
+ $X2=0 $Y2=0
cc_503 N_A_1169_93#_c_715_n N_A_982_369#_c_879_n 6.32206e-19 $X=6.16 $Y=1.425
+ $X2=0 $Y2=0
cc_504 N_A_1169_93#_c_743_n N_A_982_369#_c_879_n 0.0192312f $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_505 N_A_1169_93#_c_718_n N_A_982_369#_c_879_n 0.00165031f $X=6.16 $Y=1.59
+ $X2=0 $Y2=0
cc_506 N_A_1169_93#_c_734_n N_A_982_369#_c_879_n 0.0203812f $X=6.9 $Y=2.075
+ $X2=0 $Y2=0
cc_507 N_A_1169_93#_c_719_n N_A_982_369#_c_879_n 0.00879f $X=7.05 $Y=1.255 $X2=0
+ $Y2=0
cc_508 N_A_1169_93#_c_720_n N_A_982_369#_c_879_n 0.0224308f $X=7.067 $Y=1.985
+ $X2=0 $Y2=0
cc_509 N_A_1169_93#_c_722_n N_A_982_369#_c_879_n 0.00897551f $X=6.825 $Y=0.52
+ $X2=0 $Y2=0
cc_510 N_A_1169_93#_c_723_n N_A_982_369#_c_879_n 0.021042f $X=7.27 $Y=1.35 $X2=0
+ $Y2=0
cc_511 N_A_1169_93#_c_715_n N_A_982_369#_c_880_n 0.00469429f $X=6.16 $Y=1.425
+ $X2=0 $Y2=0
cc_512 N_A_1169_93#_c_719_n N_A_982_369#_c_880_n 0.00142989f $X=7.05 $Y=1.255
+ $X2=0 $Y2=0
cc_513 N_A_1169_93#_c_722_n N_A_982_369#_c_880_n 0.00401256f $X=6.825 $Y=0.52
+ $X2=0 $Y2=0
cc_514 N_A_1169_93#_c_723_n N_A_982_369#_c_880_n 0.00185208f $X=7.27 $Y=1.35
+ $X2=0 $Y2=0
cc_515 N_A_1169_93#_c_724_n N_A_982_369#_c_880_n 0.0172518f $X=7.27 $Y=1.35
+ $X2=0 $Y2=0
cc_516 N_A_1169_93#_c_721_n N_A_1513_137#_M1018_s 0.00246333f $X=9.37 $Y=0.63
+ $X2=-0.19 $Y2=-0.245
cc_517 N_A_1169_93#_M1018_g N_A_1513_137#_c_962_n 0.0132154f $X=7.925 $Y=0.895
+ $X2=0 $Y2=0
cc_518 N_A_1169_93#_c_721_n N_A_1513_137#_c_962_n 0.0162938f $X=9.37 $Y=0.63
+ $X2=0 $Y2=0
cc_519 N_A_1169_93#_M1021_g N_A_1513_137#_M1011_g 0.0117051f $X=7.925 $Y=2.155
+ $X2=0 $Y2=0
cc_520 N_A_1169_93#_M1013_g N_A_1513_137#_c_964_n 0.0279828f $X=9.61 $Y=0.685
+ $X2=0 $Y2=0
cc_521 N_A_1169_93#_c_721_n N_A_1513_137#_c_964_n 0.015972f $X=9.37 $Y=0.63
+ $X2=0 $Y2=0
cc_522 N_A_1169_93#_c_726_n N_A_1513_137#_c_964_n 0.00693582f $X=9.462 $Y=1.32
+ $X2=0 $Y2=0
cc_523 N_A_1169_93#_M1003_g N_A_1513_137#_M1031_g 0.0311107f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_524 N_A_1169_93#_M1021_g N_A_1513_137#_c_966_n 0.00768702f $X=7.925 $Y=2.155
+ $X2=0 $Y2=0
cc_525 N_A_1169_93#_c_720_n N_A_1513_137#_c_966_n 0.00766485f $X=7.067 $Y=1.985
+ $X2=0 $Y2=0
cc_526 N_A_1169_93#_c_709_n N_A_1513_137#_c_967_n 0.0185008f $X=7.85 $Y=1.44
+ $X2=0 $Y2=0
cc_527 N_A_1169_93#_M1018_g N_A_1513_137#_c_967_n 0.0192788f $X=7.925 $Y=0.895
+ $X2=0 $Y2=0
cc_528 N_A_1169_93#_M1021_g N_A_1513_137#_c_967_n 0.012068f $X=7.925 $Y=2.155
+ $X2=0 $Y2=0
cc_529 N_A_1169_93#_c_717_n N_A_1513_137#_c_967_n 0.00349549f $X=7.925 $Y=1.44
+ $X2=0 $Y2=0
cc_530 N_A_1169_93#_c_719_n N_A_1513_137#_c_967_n 0.00677497f $X=7.05 $Y=1.255
+ $X2=0 $Y2=0
cc_531 N_A_1169_93#_c_720_n N_A_1513_137#_c_967_n 0.00490455f $X=7.067 $Y=1.985
+ $X2=0 $Y2=0
cc_532 N_A_1169_93#_c_721_n N_A_1513_137#_c_967_n 0.0610733f $X=9.37 $Y=0.63
+ $X2=0 $Y2=0
cc_533 N_A_1169_93#_c_722_n N_A_1513_137#_c_967_n 0.00897033f $X=6.825 $Y=0.52
+ $X2=0 $Y2=0
cc_534 N_A_1169_93#_c_723_n N_A_1513_137#_c_967_n 0.021734f $X=7.27 $Y=1.35
+ $X2=0 $Y2=0
cc_535 N_A_1169_93#_c_724_n N_A_1513_137#_c_967_n 0.00142824f $X=7.27 $Y=1.35
+ $X2=0 $Y2=0
cc_536 N_A_1169_93#_c_709_n N_A_1513_137#_c_972_n 0.00233385f $X=7.85 $Y=1.44
+ $X2=0 $Y2=0
cc_537 N_A_1169_93#_M1021_g N_A_1513_137#_c_972_n 0.00826205f $X=7.925 $Y=2.155
+ $X2=0 $Y2=0
cc_538 N_A_1169_93#_c_736_n N_A_1513_137#_c_972_n 0.0151699f $X=7.005 $Y=2.4
+ $X2=0 $Y2=0
cc_539 N_A_1169_93#_c_720_n N_A_1513_137#_c_972_n 0.00789392f $X=7.067 $Y=1.985
+ $X2=0 $Y2=0
cc_540 N_A_1169_93#_c_738_n N_A_1513_137#_c_972_n 0.00917249f $X=7.035 $Y=2.075
+ $X2=0 $Y2=0
cc_541 N_A_1169_93#_M1018_g N_A_1513_137#_c_968_n 0.0214264f $X=7.925 $Y=0.895
+ $X2=0 $Y2=0
cc_542 N_A_1169_93#_c_721_n N_A_1513_137#_c_968_n 0.0012495f $X=9.37 $Y=0.63
+ $X2=0 $Y2=0
cc_543 N_A_1169_93#_c_725_n N_A_1513_137#_c_968_n 0.00119517f $X=9.47 $Y=1.485
+ $X2=0 $Y2=0
cc_544 N_A_1169_93#_c_727_n N_A_1513_137#_c_968_n 0.0226188f $X=10.04 $Y=1.485
+ $X2=0 $Y2=0
cc_545 N_A_1169_93#_M1010_g N_VPWR_c_1031_n 0.0128203f $X=6.22 $Y=2.465 $X2=0
+ $Y2=0
cc_546 N_A_1169_93#_c_734_n N_VPWR_c_1031_n 0.0296402f $X=6.9 $Y=2.075 $X2=0
+ $Y2=0
cc_547 N_A_1169_93#_c_735_n N_VPWR_c_1031_n 0.00338407f $X=6.325 $Y=2.075 $X2=0
+ $Y2=0
cc_548 N_A_1169_93#_M1021_g N_VPWR_c_1032_n 0.00627954f $X=7.925 $Y=2.155 $X2=0
+ $Y2=0
cc_549 N_A_1169_93#_M1003_g N_VPWR_c_1033_n 0.00972049f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_550 N_A_1169_93#_c_725_n N_VPWR_c_1033_n 0.00962869f $X=9.47 $Y=1.485 $X2=0
+ $Y2=0
cc_551 N_A_1169_93#_c_727_n N_VPWR_c_1033_n 0.00378792f $X=10.04 $Y=1.485 $X2=0
+ $Y2=0
cc_552 N_A_1169_93#_M1012_g N_VPWR_c_1035_n 0.00772993f $X=10.035 $Y=2.465 $X2=0
+ $Y2=0
cc_553 N_A_1169_93#_M1021_g N_VPWR_c_1036_n 0.00312414f $X=7.925 $Y=2.155 $X2=0
+ $Y2=0
cc_554 N_A_1169_93#_c_736_n N_VPWR_c_1036_n 0.0181659f $X=7.005 $Y=2.4 $X2=0
+ $Y2=0
cc_555 N_A_1169_93#_M1010_g N_VPWR_c_1040_n 0.00332367f $X=6.22 $Y=2.465 $X2=0
+ $Y2=0
cc_556 N_A_1169_93#_M1003_g N_VPWR_c_1042_n 0.00585385f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_557 N_A_1169_93#_M1012_g N_VPWR_c_1042_n 0.00585385f $X=10.035 $Y=2.465 $X2=0
+ $Y2=0
cc_558 N_A_1169_93#_M1030_d N_VPWR_c_1026_n 0.00336915f $X=6.865 $Y=2.255 $X2=0
+ $Y2=0
cc_559 N_A_1169_93#_M1010_g N_VPWR_c_1026_n 0.00387424f $X=6.22 $Y=2.465 $X2=0
+ $Y2=0
cc_560 N_A_1169_93#_M1021_g N_VPWR_c_1026_n 0.00410284f $X=7.925 $Y=2.155 $X2=0
+ $Y2=0
cc_561 N_A_1169_93#_M1003_g N_VPWR_c_1026_n 0.0111197f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_562 N_A_1169_93#_M1012_g N_VPWR_c_1026_n 0.0115127f $X=10.035 $Y=2.465 $X2=0
+ $Y2=0
cc_563 N_A_1169_93#_c_736_n N_VPWR_c_1026_n 0.0104192f $X=7.005 $Y=2.4 $X2=0
+ $Y2=0
cc_564 N_A_1169_93#_c_721_n N_Q_N_M1020_d 0.00422717f $X=9.37 $Y=0.63 $X2=-0.19
+ $Y2=-0.245
cc_565 N_A_1169_93#_M1018_g N_Q_N_c_1165_n 4.01888e-19 $X=7.925 $Y=0.895 $X2=0
+ $Y2=0
cc_566 N_A_1169_93#_M1021_g N_Q_N_c_1165_n 9.49157e-19 $X=7.925 $Y=2.155 $X2=0
+ $Y2=0
cc_567 N_A_1169_93#_M1003_g N_Q_N_c_1165_n 0.00102144f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_568 N_A_1169_93#_M1013_g N_Q_N_c_1165_n 3.80281e-19 $X=9.61 $Y=0.685 $X2=0
+ $Y2=0
cc_569 N_A_1169_93#_c_721_n N_Q_N_c_1165_n 0.0170777f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_570 N_A_1169_93#_c_726_n N_Q_N_c_1165_n 0.0287566f $X=9.462 $Y=1.32 $X2=0
+ $Y2=0
cc_571 N_A_1169_93#_c_727_n N_Q_N_c_1165_n 0.00113285f $X=10.04 $Y=1.485 $X2=0
+ $Y2=0
cc_572 N_A_1169_93#_c_726_n N_Q_c_1183_n 0.0150162f $X=9.462 $Y=1.32 $X2=0 $Y2=0
cc_573 N_A_1169_93#_M1003_g Q 0.00509559f $X=9.605 $Y=2.465 $X2=0 $Y2=0
cc_574 N_A_1169_93#_M1013_g Q 0.00136561f $X=9.61 $Y=0.685 $X2=0 $Y2=0
cc_575 N_A_1169_93#_M1012_g Q 0.0053545f $X=10.035 $Y=2.465 $X2=0 $Y2=0
cc_576 N_A_1169_93#_c_725_n Q 0.0219374f $X=9.47 $Y=1.485 $X2=0 $Y2=0
cc_577 N_A_1169_93#_c_726_n Q 0.0117936f $X=9.462 $Y=1.32 $X2=0 $Y2=0
cc_578 N_A_1169_93#_c_727_n Q 0.0293723f $X=10.04 $Y=1.485 $X2=0 $Y2=0
cc_579 N_A_1169_93#_M1013_g N_Q_c_1185_n 0.00107166f $X=9.61 $Y=0.685 $X2=0
+ $Y2=0
cc_580 N_A_1169_93#_M1014_g N_Q_c_1185_n 0.00614953f $X=10.04 $Y=0.685 $X2=0
+ $Y2=0
cc_581 N_A_1169_93#_c_721_n N_VGND_M1018_d 0.00911084f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_582 N_A_1169_93#_c_721_n N_VGND_M1029_s 0.0109575f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_583 N_A_1169_93#_c_726_n N_VGND_M1029_s 0.00487338f $X=9.462 $Y=1.32 $X2=0
+ $Y2=0
cc_584 N_A_1169_93#_c_708_n N_VGND_c_1208_n 0.012591f $X=5.92 $Y=1.125 $X2=0
+ $Y2=0
cc_585 N_A_1169_93#_c_714_n N_VGND_c_1208_n 0.00400331f $X=6.07 $Y=1.2 $X2=0
+ $Y2=0
cc_586 N_A_1169_93#_c_722_n N_VGND_c_1208_n 0.0254434f $X=6.825 $Y=0.52 $X2=0
+ $Y2=0
cc_587 N_A_1169_93#_M1014_g N_VGND_c_1210_n 0.00715682f $X=10.04 $Y=0.685 $X2=0
+ $Y2=0
cc_588 N_A_1169_93#_c_721_n N_VGND_c_1211_n 0.0242865f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_589 N_A_1169_93#_M1018_g N_VGND_c_1212_n 6.49089e-19 $X=7.925 $Y=0.895 $X2=0
+ $Y2=0
cc_590 N_A_1169_93#_c_721_n N_VGND_c_1212_n 0.021458f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_591 N_A_1169_93#_c_722_n N_VGND_c_1212_n 0.0205312f $X=6.825 $Y=0.52 $X2=0
+ $Y2=0
cc_592 N_A_1169_93#_c_708_n N_VGND_c_1215_n 0.0035863f $X=5.92 $Y=1.125 $X2=0
+ $Y2=0
cc_593 N_A_1169_93#_c_721_n N_VGND_c_1216_n 0.0132159f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_594 N_A_1169_93#_M1013_g N_VGND_c_1217_n 0.00549656f $X=9.61 $Y=0.685 $X2=0
+ $Y2=0
cc_595 N_A_1169_93#_M1014_g N_VGND_c_1217_n 0.00555245f $X=10.04 $Y=0.685 $X2=0
+ $Y2=0
cc_596 N_A_1169_93#_c_721_n N_VGND_c_1217_n 7.9879e-19 $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_597 N_A_1169_93#_M1013_g N_VGND_c_1221_n 0.00239955f $X=9.61 $Y=0.685 $X2=0
+ $Y2=0
cc_598 N_A_1169_93#_c_721_n N_VGND_c_1221_n 0.0248835f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_599 N_A_1169_93#_c_708_n N_VGND_c_1222_n 0.00401353f $X=5.92 $Y=1.125 $X2=0
+ $Y2=0
cc_600 N_A_1169_93#_M1013_g N_VGND_c_1222_n 0.0106644f $X=9.61 $Y=0.685 $X2=0
+ $Y2=0
cc_601 N_A_1169_93#_M1014_g N_VGND_c_1222_n 0.0112297f $X=10.04 $Y=0.685 $X2=0
+ $Y2=0
cc_602 N_A_1169_93#_c_721_n N_VGND_c_1222_n 0.0558038f $X=9.37 $Y=0.63 $X2=0
+ $Y2=0
cc_603 N_A_1169_93#_c_722_n N_VGND_c_1222_n 0.0172655f $X=6.825 $Y=0.52 $X2=0
+ $Y2=0
cc_604 N_A_982_369#_M1030_g N_A_1513_137#_c_972_n 0.00176197f $X=6.79 $Y=2.675
+ $X2=0 $Y2=0
cc_605 N_A_982_369#_M1030_g N_VPWR_c_1031_n 0.0206935f $X=6.79 $Y=2.675 $X2=0
+ $Y2=0
cc_606 N_A_982_369#_M1030_g N_VPWR_c_1036_n 0.00525069f $X=6.79 $Y=2.675 $X2=0
+ $Y2=0
cc_607 N_A_982_369#_c_876_n N_VPWR_c_1040_n 0.00512837f $X=5.4 $Y=1.99 $X2=0
+ $Y2=0
cc_608 N_A_982_369#_M1030_g N_VPWR_c_1026_n 0.0101648f $X=6.79 $Y=2.675 $X2=0
+ $Y2=0
cc_609 N_A_982_369#_c_876_n N_VPWR_c_1026_n 0.0075815f $X=5.4 $Y=1.99 $X2=0
+ $Y2=0
cc_610 N_A_982_369#_M1005_g N_VGND_c_1208_n 0.00734531f $X=6.61 $Y=0.695 $X2=0
+ $Y2=0
cc_611 N_A_982_369#_c_877_n N_VGND_c_1208_n 0.0390191f $X=6.535 $Y=1.23 $X2=0
+ $Y2=0
cc_612 N_A_982_369#_c_895_n N_VGND_c_1208_n 0.0132749f $X=5.44 $Y=0.807 $X2=0
+ $Y2=0
cc_613 N_A_982_369#_M1005_g N_VGND_c_1212_n 0.00430542f $X=6.61 $Y=0.695 $X2=0
+ $Y2=0
cc_614 N_A_982_369#_c_895_n N_VGND_c_1215_n 0.00826777f $X=5.44 $Y=0.807 $X2=0
+ $Y2=0
cc_615 N_A_982_369#_M1005_g N_VGND_c_1222_n 0.00544287f $X=6.61 $Y=0.695 $X2=0
+ $Y2=0
cc_616 N_A_982_369#_c_895_n N_VGND_c_1222_n 0.0122895f $X=5.44 $Y=0.807 $X2=0
+ $Y2=0
cc_617 N_A_1513_137#_M1011_g N_VPWR_c_1032_n 0.0109648f $X=8.59 $Y=2.465 $X2=0
+ $Y2=0
cc_618 N_A_1513_137#_c_967_n N_VPWR_c_1032_n 0.036614f $X=7.71 $Y=0.98 $X2=0
+ $Y2=0
cc_619 N_A_1513_137#_c_972_n N_VPWR_c_1032_n 0.0261555f $X=7.71 $Y=1.98 $X2=0
+ $Y2=0
cc_620 N_A_1513_137#_c_968_n N_VPWR_c_1032_n 0.00166391f $X=9.02 $Y=1.38 $X2=0
+ $Y2=0
cc_621 N_A_1513_137#_M1031_g N_VPWR_c_1033_n 0.0109758f $X=9.02 $Y=2.465 $X2=0
+ $Y2=0
cc_622 N_A_1513_137#_M1011_g N_VPWR_c_1041_n 0.0054895f $X=8.59 $Y=2.465 $X2=0
+ $Y2=0
cc_623 N_A_1513_137#_M1031_g N_VPWR_c_1041_n 0.0054895f $X=9.02 $Y=2.465 $X2=0
+ $Y2=0
cc_624 N_A_1513_137#_M1011_g N_VPWR_c_1026_n 0.0110654f $X=8.59 $Y=2.465 $X2=0
+ $Y2=0
cc_625 N_A_1513_137#_M1031_g N_VPWR_c_1026_n 0.010281f $X=9.02 $Y=2.465 $X2=0
+ $Y2=0
cc_626 N_A_1513_137#_c_972_n N_VPWR_c_1026_n 0.012771f $X=7.71 $Y=1.98 $X2=0
+ $Y2=0
cc_627 N_A_1513_137#_c_962_n N_Q_N_c_1165_n 0.00516625f $X=8.59 $Y=1.215 $X2=0
+ $Y2=0
cc_628 N_A_1513_137#_M1011_g N_Q_N_c_1165_n 0.0239069f $X=8.59 $Y=2.465 $X2=0
+ $Y2=0
cc_629 N_A_1513_137#_c_964_n N_Q_N_c_1165_n 0.00677698f $X=9.02 $Y=1.215 $X2=0
+ $Y2=0
cc_630 N_A_1513_137#_M1031_g N_Q_N_c_1165_n 0.0240204f $X=9.02 $Y=2.465 $X2=0
+ $Y2=0
cc_631 N_A_1513_137#_c_967_n N_Q_N_c_1165_n 0.0501581f $X=7.71 $Y=0.98 $X2=0
+ $Y2=0
cc_632 N_A_1513_137#_c_968_n N_Q_N_c_1165_n 0.023481f $X=9.02 $Y=1.38 $X2=0
+ $Y2=0
cc_633 N_A_1513_137#_c_967_n N_VGND_M1018_d 0.00671139f $X=7.71 $Y=0.98 $X2=0
+ $Y2=0
cc_634 N_A_1513_137#_c_962_n N_VGND_c_1211_n 0.00884127f $X=8.59 $Y=1.215 $X2=0
+ $Y2=0
cc_635 N_A_1513_137#_c_962_n N_VGND_c_1216_n 0.00387708f $X=8.59 $Y=1.215 $X2=0
+ $Y2=0
cc_636 N_A_1513_137#_c_964_n N_VGND_c_1216_n 0.00387708f $X=9.02 $Y=1.215 $X2=0
+ $Y2=0
cc_637 N_A_1513_137#_c_964_n N_VGND_c_1221_n 0.00381978f $X=9.02 $Y=1.215 $X2=0
+ $Y2=0
cc_638 N_A_1513_137#_c_962_n N_VGND_c_1222_n 0.00656008f $X=8.59 $Y=1.215 $X2=0
+ $Y2=0
cc_639 N_A_1513_137#_c_964_n N_VGND_c_1222_n 0.00567145f $X=9.02 $Y=1.215 $X2=0
+ $Y2=0
cc_640 N_VPWR_c_1026_n N_Q_N_M1011_s 0.00223559f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_641 N_VPWR_c_1032_n N_Q_N_c_1165_n 0.0480995f $X=8.14 $Y=1.98 $X2=0 $Y2=0
cc_642 N_VPWR_c_1033_n N_Q_N_c_1165_n 0.0455403f $X=9.315 $Y=1.985 $X2=0 $Y2=0
cc_643 N_VPWR_c_1041_n N_Q_N_c_1165_n 0.0189236f $X=9.15 $Y=3.33 $X2=0 $Y2=0
cc_644 N_VPWR_c_1026_n N_Q_N_c_1165_n 0.0123859f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_645 N_VPWR_c_1026_n N_Q_M1003_d 0.00432284f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_646 N_VPWR_c_1033_n Q 8.51311e-19 $X=9.315 $Y=1.985 $X2=0 $Y2=0
cc_647 N_VPWR_c_1035_n Q 0.00151856f $X=10.25 $Y=1.98 $X2=0 $Y2=0
cc_648 N_VPWR_c_1042_n Q 0.0135169f $X=10.125 $Y=3.33 $X2=0 $Y2=0
cc_649 N_VPWR_c_1026_n Q 0.00847005f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_650 N_A_429_119#_c_1140_n N_VGND_c_1214_n 0.00698304f $X=2.51 $Y=0.79 $X2=0
+ $Y2=0
cc_651 N_A_429_119#_c_1140_n N_VGND_c_1222_n 0.0105404f $X=2.51 $Y=0.79 $X2=0
+ $Y2=0
cc_652 N_Q_c_1185_n N_VGND_c_1210_n 0.00225185f $X=9.825 $Y=0.42 $X2=0 $Y2=0
cc_653 N_Q_c_1185_n N_VGND_c_1217_n 0.016703f $X=9.825 $Y=0.42 $X2=0 $Y2=0
cc_654 N_Q_c_1185_n N_VGND_c_1221_n 5.73528e-19 $X=9.825 $Y=0.42 $X2=0 $Y2=0
cc_655 N_Q_c_1185_n N_VGND_c_1222_n 0.0090585f $X=9.825 $Y=0.42 $X2=0 $Y2=0
