* File: sky130_fd_sc_lp__nor4b_m.pex.spice
* Created: Wed Sep  2 10:11:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4B_M%D_N 3 9 11 12 13 14 15 16 17 24
r46 24 26 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.627 $Y=1.615
+ $X2=0.627 $Y2=1.45
r47 16 17 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.69 $Y=1.615
+ $X2=0.69 $Y2=2.035
r48 16 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.66
+ $Y=1.615 $X2=0.66 $Y2=1.615
r49 15 16 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.69 $Y=1.295
+ $X2=0.69 $Y2=1.615
r50 14 15 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=0.925
+ $X2=0.69 $Y2=1.295
r51 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=0.555
+ $X2=0.69 $Y2=0.925
r52 11 12 43.452 $w=3.95e-07 $l=1.5e-07 $layer=POLY_cond $X=0.725 $Y=1.97
+ $X2=0.725 $Y2=2.12
r53 9 12 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.945 $Y=2.69
+ $X2=0.945 $Y2=2.12
r54 5 24 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.627 $Y=1.647
+ $X2=0.627 $Y2=1.615
r55 5 11 45.4779 $w=3.95e-07 $l=3.23e-07 $layer=POLY_cond $X=0.627 $Y=1.647
+ $X2=0.627 $Y2=1.97
r56 3 26 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.505 $Y=0.55 $X2=0.505
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_M%A 2 5 8 11 13 16 18 19 20 21 27
r55 27 29 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.207 $Y=1.225
+ $X2=1.207 $Y2=1.06
r56 20 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.2
+ $Y2=2.035
r57 19 20 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.2 $Y=1.225 $X2=1.2
+ $Y2=1.665
r58 19 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2
+ $Y=1.225 $X2=1.2 $Y2=1.225
r59 18 19 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=1.225
r60 14 16 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.305 $Y=2.195
+ $X2=1.485 $Y2=2.195
r61 9 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.485 $Y=2.27
+ $X2=1.485 $Y2=2.195
r62 9 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.485 $Y=2.27
+ $X2=1.485 $Y2=2.69
r63 8 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.305 $Y=2.12
+ $X2=1.305 $Y2=2.195
r64 8 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.305 $Y=2.12
+ $X2=1.305 $Y2=1.73
r65 5 29 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.305 $Y=0.55
+ $X2=1.305 $Y2=1.06
r66 2 13 47.5363 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=1.207 $Y=1.558
+ $X2=1.207 $Y2=1.73
r67 1 27 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=1.207 $Y=1.232
+ $X2=1.207 $Y2=1.225
r68 1 2 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=1.207 $Y=1.232
+ $X2=1.207 $Y2=1.558
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_M%B 3 7 11 12 13 14 15 20
c44 13 0 4.85574e-20 $X=1.68 $Y=1.295
r45 14 15 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.665
+ $X2=1.717 $Y2=2.035
r46 13 14 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.295
+ $X2=1.717 $Y2=1.665
r47 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.755
+ $Y=1.375 $X2=1.755 $Y2=1.375
r48 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.755 $Y=1.715
+ $X2=1.755 $Y2=1.375
r49 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.715
+ $X2=1.755 $Y2=1.88
r50 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.21
+ $X2=1.755 $Y2=1.375
r51 7 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.845 $Y=2.69
+ $X2=1.845 $Y2=1.88
r52 3 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.735 $Y=0.55
+ $X2=1.735 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_M%C 3 7 11 12 13 14 15 20
c45 7 0 1.25011e-19 $X=2.245 $Y=0.55
r46 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.295
+ $Y=1.425 $X2=2.295 $Y2=1.425
r47 14 15 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.227 $Y=1.665
+ $X2=2.227 $Y2=2.035
r48 14 21 9.0684 $w=3.03e-07 $l=2.4e-07 $layer=LI1_cond $X=2.227 $Y=1.665
+ $X2=2.227 $Y2=1.425
r49 13 21 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=2.227 $Y=1.295
+ $X2=2.227 $Y2=1.425
r50 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=1.425
r51 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=1.93
r52 10 20 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.26
+ $X2=2.295 $Y2=1.425
r53 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.245 $Y=0.55
+ $X2=2.245 $Y2=1.26
r54 3 12 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.205 $Y=2.69
+ $X2=2.205 $Y2=1.93
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_M%A_33_68# 1 2 9 11 13 19 23 26 29 31 32 35 37
+ 41 42 44
r75 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.835
+ $Y=1.815 $X2=2.835 $Y2=1.815
r76 39 41 15.526 $w=3.58e-07 $l=4.85e-07 $layer=LI1_cond $X=2.74 $Y=2.3 $X2=2.74
+ $Y2=1.815
r77 38 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.835 $Y=2.385
+ $X2=0.73 $Y2=2.385
r78 37 39 31.798 $w=6.6e-08 $l=2.18403e-07 $layer=LI1_cond $X=2.56 $Y=2.385
+ $X2=2.74 $Y2=2.3
r79 37 38 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=2.56 $Y=2.385
+ $X2=0.835 $Y2=2.385
r80 33 44 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.47
+ $X2=0.73 $Y2=2.385
r81 33 35 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.73 $Y=2.47
+ $X2=0.73 $Y2=2.625
r82 31 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.625 $Y=2.385
+ $X2=0.73 $Y2=2.385
r83 31 32 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.625 $Y=2.385
+ $X2=0.395 $Y2=2.385
r84 27 32 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.29 $Y=2.3
+ $X2=0.395 $Y2=2.385
r85 27 29 88.9913 $w=2.08e-07 $l=1.685e-06 $layer=LI1_cond $X=0.29 $Y=2.3
+ $X2=0.29 $Y2=0.615
r86 26 42 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.65
+ $X2=2.835 $Y2=1.815
r87 21 23 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.675 $Y=0.945
+ $X2=2.775 $Y2=0.945
r88 19 42 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.835 $Y=2.17
+ $X2=2.835 $Y2=1.815
r89 16 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.565 $Y=2.245
+ $X2=2.835 $Y2=2.245
r90 14 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.775 $Y=1.02
+ $X2=2.775 $Y2=0.945
r91 14 26 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.775 $Y=1.02
+ $X2=2.775 $Y2=1.65
r92 11 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.675 $Y=0.87
+ $X2=2.675 $Y2=0.945
r93 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.675 $Y=0.87
+ $X2=2.675 $Y2=0.55
r94 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.565 $Y=2.32
+ $X2=2.565 $Y2=2.245
r95 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.565 $Y=2.32
+ $X2=2.565 $Y2=2.69
r96 2 35 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=2.48 $X2=0.73 $Y2=2.625
r97 1 29 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.34 $X2=0.29 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_M%VPWR 1 6 8 10 20 21 24
r26 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r27 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r28 17 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r29 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r30 15 17 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r31 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r34 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 8 21 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33 $X2=1.2
+ $Y2=3.33
r37 8 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245 $X2=1.18
+ $Y2=3.33
r39 4 6 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.18 $Y=3.245 $X2=1.18
+ $Y2=2.755
r40 1 6 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=2.48 $X2=1.18 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_M%Y 1 2 3 12 17 21 22 26 27 29 30 31 32 45
c51 17 0 7.64536e-20 $X=1.6 $Y=0.555
r52 32 45 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.925
+ $X2=3.1 $Y2=0.925
r53 32 45 2.15294 $w=1.68e-07 $l=3.3e-08 $layer=LI1_cond $X=3.067 $Y=0.925
+ $X2=3.1 $Y2=0.925
r54 31 32 27.8578 $w=1.68e-07 $l=4.27e-07 $layer=LI1_cond $X=2.64 $Y=0.925
+ $X2=3.067 $Y2=0.925
r55 29 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=0.925
+ $X2=1.685 $Y2=0.925
r56 29 30 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.725 $Y=0.925
+ $X2=2.16 $Y2=0.925
r57 29 41 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.725 $Y=0.925
+ $X2=1.685 $Y2=0.925
r58 27 32 63.6674 $w=2.73e-07 $l=1.49e-06 $layer=LI1_cond $X=3.185 $Y=2.5
+ $X2=3.185 $Y2=1.01
r59 26 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=2.665
+ $X2=3.185 $Y2=2.5
r60 24 26 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.995 $Y=2.665
+ $X2=3.185 $Y2=2.665
r61 21 30 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.355 $Y=0.925
+ $X2=2.16 $Y2=0.925
r62 21 22 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.355 $Y=0.925
+ $X2=2.45 $Y2=0.925
r63 20 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.545 $Y=0.925
+ $X2=2.64 $Y2=0.925
r64 20 22 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.545 $Y=0.925
+ $X2=2.45 $Y2=0.925
r65 18 29 9.22049 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.6 $Y=0.66 $X2=1.6
+ $Y2=0.84
r66 17 18 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.6 $Y=0.555 $X2=1.6
+ $Y2=0.66
r67 15 17 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.52 $Y=0.555 $X2=1.6
+ $Y2=0.555
r68 10 22 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.84
+ $X2=2.45 $Y2=0.925
r69 10 12 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=2.45 $Y=0.84
+ $X2=2.45 $Y2=0.615
r70 3 24 600 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=2.48 $X2=2.995 $Y2=2.665
r71 2 12 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.34 $X2=2.46 $Y2=0.615
r72 1 15 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.38
+ $Y=0.34 $X2=1.52 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_M%VGND 1 2 3 12 16 20 23 24 26 27 28 29 30 31
+ 45
r46 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r48 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 31 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r51 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r52 31 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 29 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.64
+ $Y2=0
r54 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.89
+ $Y2=0
r55 28 44 4.66471 $w=1.7e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.12
+ $Y2=0
r56 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.89
+ $Y2=0
r57 26 38 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.68
+ $Y2=0
r58 26 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.97
+ $Y2=0
r59 25 41 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.64
+ $Y2=0
r60 25 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=1.97
+ $Y2=0
r61 23 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r62 23 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.08
+ $Y2=0
r63 22 38 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.68
+ $Y2=0
r64 22 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.08
+ $Y2=0
r65 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0
r66 18 20 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.89 $Y=0.085 $X2=2.89
+ $Y2=0.485
r67 14 27 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=0.085
+ $X2=1.97 $Y2=0
r68 14 16 21.1255 $w=2.08e-07 $l=4e-07 $layer=LI1_cond $X=1.97 $Y=0.085 $X2=1.97
+ $Y2=0.485
r69 10 24 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=0.085
+ $X2=1.08 $Y2=0
r70 10 12 23.3493 $w=1.88e-07 $l=4e-07 $layer=LI1_cond $X=1.08 $Y=0.085 $X2=1.08
+ $Y2=0.485
r71 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.75
+ $Y=0.34 $X2=2.89 $Y2=0.485
r72 2 16 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=0.34 $X2=1.97 $Y2=0.485
r73 1 12 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.34 $X2=1.07 $Y2=0.485
.ends

