* File: sky130_fd_sc_lp__a311oi_2.pxi.spice
* Created: Fri Aug 28 09:58:26 2020
* 
x_PM_SKY130_FD_SC_LP__A311OI_2%A3 N_A3_M1014_g N_A3_M1013_g N_A3_M1015_g
+ N_A3_M1018_g N_A3_c_102_n A3 N_A3_c_103_n N_A3_c_104_n
+ PM_SKY130_FD_SC_LP__A311OI_2%A3
x_PM_SKY130_FD_SC_LP__A311OI_2%A2 N_A2_M1005_g N_A2_M1002_g N_A2_M1012_g
+ N_A2_M1010_g A2 A2 N_A2_c_148_n N_A2_c_154_n N_A2_c_149_n
+ PM_SKY130_FD_SC_LP__A311OI_2%A2
x_PM_SKY130_FD_SC_LP__A311OI_2%A1 N_A1_M1000_g N_A1_c_207_n N_A1_c_208_n
+ N_A1_M1011_g N_A1_M1007_g N_A1_M1008_g A1 N_A1_c_211_n N_A1_c_212_n
+ PM_SKY130_FD_SC_LP__A311OI_2%A1
x_PM_SKY130_FD_SC_LP__A311OI_2%B1 N_B1_M1006_g N_B1_M1003_g N_B1_M1017_g
+ N_B1_M1019_g B1 N_B1_c_279_n N_B1_c_276_n PM_SKY130_FD_SC_LP__A311OI_2%B1
x_PM_SKY130_FD_SC_LP__A311OI_2%C1 N_C1_M1004_g N_C1_M1001_g N_C1_M1016_g
+ N_C1_M1009_g C1 C1 C1 N_C1_c_320_n PM_SKY130_FD_SC_LP__A311OI_2%C1
x_PM_SKY130_FD_SC_LP__A311OI_2%VPWR N_VPWR_M1013_s N_VPWR_M1018_s N_VPWR_M1010_d
+ N_VPWR_M1011_s N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_362_n
+ N_VPWR_c_363_n VPWR N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n
+ N_VPWR_c_367_n N_VPWR_c_358_n N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n
+ PM_SKY130_FD_SC_LP__A311OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A311OI_2%A_135_367# N_A_135_367#_M1013_d
+ N_A_135_367#_M1002_s N_A_135_367#_M1000_d N_A_135_367#_M1003_d
+ N_A_135_367#_c_465_n N_A_135_367#_c_438_n N_A_135_367#_c_439_n
+ N_A_135_367#_c_450_n N_A_135_367#_c_453_n N_A_135_367#_c_440_n
+ N_A_135_367#_c_454_n N_A_135_367#_c_459_n
+ PM_SKY130_FD_SC_LP__A311OI_2%A_135_367#
x_PM_SKY130_FD_SC_LP__A311OI_2%A_727_367# N_A_727_367#_M1003_s
+ N_A_727_367#_M1019_s N_A_727_367#_M1009_d N_A_727_367#_c_491_n
+ N_A_727_367#_c_518_p N_A_727_367#_c_497_n N_A_727_367#_c_492_n
+ N_A_727_367#_c_493_n N_A_727_367#_c_510_n
+ PM_SKY130_FD_SC_LP__A311OI_2%A_727_367#
x_PM_SKY130_FD_SC_LP__A311OI_2%Y N_Y_M1007_s N_Y_M1008_s N_Y_M1017_d N_Y_M1016_d
+ N_Y_M1001_s N_Y_c_520_n N_Y_c_521_n N_Y_c_522_n N_Y_c_523_n N_Y_c_524_n
+ N_Y_c_525_n N_Y_c_526_n N_Y_c_527_n N_Y_c_528_n N_Y_c_529_n N_Y_c_530_n
+ N_Y_c_532_n N_Y_c_580_n Y Y Y Y Y N_Y_c_538_n Y PM_SKY130_FD_SC_LP__A311OI_2%Y
x_PM_SKY130_FD_SC_LP__A311OI_2%A_48_69# N_A_48_69#_M1014_s N_A_48_69#_M1015_s
+ N_A_48_69#_M1012_s N_A_48_69#_c_621_n N_A_48_69#_c_622_n N_A_48_69#_c_623_n
+ N_A_48_69#_c_624_n N_A_48_69#_c_625_n N_A_48_69#_c_626_n N_A_48_69#_c_627_n
+ PM_SKY130_FD_SC_LP__A311OI_2%A_48_69#
x_PM_SKY130_FD_SC_LP__A311OI_2%VGND N_VGND_M1014_d N_VGND_M1006_s N_VGND_M1004_s
+ N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n VGND N_VGND_c_666_n
+ N_VGND_c_667_n N_VGND_c_668_n N_VGND_c_669_n N_VGND_c_670_n N_VGND_c_671_n
+ N_VGND_c_672_n PM_SKY130_FD_SC_LP__A311OI_2%VGND
x_PM_SKY130_FD_SC_LP__A311OI_2%A_307_69# N_A_307_69#_M1005_d N_A_307_69#_M1007_d
+ N_A_307_69#_c_734_n N_A_307_69#_c_731_n N_A_307_69#_c_732_n
+ N_A_307_69#_c_741_n PM_SKY130_FD_SC_LP__A311OI_2%A_307_69#
cc_1 VNB N_A3_M1014_g 0.0245211f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.765
cc_2 VNB N_A3_M1015_g 0.0182362f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.765
cc_3 VNB N_A3_c_102_n 0.00129035f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.5
cc_4 VNB N_A3_c_103_n 0.0557607f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.505
cc_5 VNB N_A3_c_104_n 0.0119784f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.582
cc_6 VNB N_A2_M1005_g 0.0184468f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.765
cc_7 VNB N_A2_M1012_g 0.0235659f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.765
cc_8 VNB A2 0.0135347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_c_148_n 0.0520168f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.505
cc_10 VNB N_A2_c_149_n 0.00129035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_207_n 0.011234f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.675
cc_12 VNB N_A1_c_208_n 0.00767002f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_13 VNB N_A1_M1007_g 0.0237181f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.675
cc_14 VNB N_A1_M1008_g 0.0195969f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.5
cc_15 VNB N_A1_c_211_n 0.0367082f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.505
cc_16 VNB N_A1_c_212_n 0.00213611f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_17 VNB N_B1_M1006_g 0.019408f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.765
cc_18 VNB N_B1_M1017_g 0.0194073f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.765
cc_19 VNB N_B1_c_276_n 0.032197f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.505
cc_20 VNB N_C1_M1004_g 0.0194073f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.765
cc_21 VNB N_C1_M1016_g 0.0259905f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.765
cc_22 VNB C1 0.0166233f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.5
cc_23 VNB N_C1_c_320_n 0.0369905f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.505
cc_24 VNB N_VPWR_c_358_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_520_n 0.00522425f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.5
cc_26 VNB N_Y_c_521_n 0.00490807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_522_n 0.00320383f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_Y_c_523_n 0.00183929f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_29 VNB N_Y_c_524_n 0.00387041f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.505
cc_30 VNB N_Y_c_525_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_526_n 0.0132586f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.582
cc_32 VNB N_Y_c_527_n 0.0326282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_528_n 0.00476715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_529_n 0.00276309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_530_n 0.00178419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_48_69#_c_621_n 0.0300387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_48_69#_c_622_n 0.0031384f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=2.465
cc_38 VNB N_A_48_69#_c_623_n 0.00878964f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=2.465
cc_39 VNB N_A_48_69#_c_624_n 0.00189149f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.5
cc_40 VNB N_A_48_69#_c_625_n 0.00767986f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.5
cc_41 VNB N_A_48_69#_c_626_n 0.00591013f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.505
cc_42 VNB N_A_48_69#_c_627_n 0.00286334f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_43 VNB N_VGND_c_663_n 0.00332106f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=2.465
cc_44 VNB N_VGND_c_664_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.5
cc_45 VNB N_VGND_c_665_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_VGND_c_666_n 0.0737279f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_47 VNB N_VGND_c_667_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_668_n 0.0166602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_669_n 0.328188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_670_n 0.0261255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_671_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_672_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_307_69#_c_731_n 0.0241728f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.765
cc_54 VNB N_A_307_69#_c_732_n 0.00203674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_A3_M1013_g 0.0238666f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_56 VPB N_A3_M1018_g 0.0179917f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=2.465
cc_57 VPB N_A3_c_103_n 0.0138688f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.505
cc_58 VPB N_A3_c_104_n 0.00886774f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.582
cc_59 VPB N_A2_M1002_g 0.0179917f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_60 VPB N_A2_M1010_g 0.0207915f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=2.465
cc_61 VPB A2 0.00332745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A2_c_148_n 0.0135296f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.505
cc_63 VPB N_A2_c_154_n 0.00294131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A1_M1000_g 0.0204986f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=0.765
cc_65 VPB N_A1_c_207_n 0.00300811f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.675
cc_66 VPB N_A1_c_208_n 5.21411e-19 $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_67 VPB N_A1_M1011_g 0.0215831f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.335
cc_68 VPB N_A1_c_211_n 0.0174746f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.505
cc_69 VPB N_A1_c_212_n 0.00478185f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_70 VPB N_B1_M1003_g 0.0239943f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_71 VPB N_B1_M1019_g 0.0186259f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=2.465
cc_72 VPB N_B1_c_279_n 0.00209697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_B1_c_276_n 0.00471452f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.505
cc_74 VPB N_C1_M1001_g 0.0183424f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_75 VPB N_C1_M1009_g 0.0244533f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=2.465
cc_76 VPB C1 0.0142626f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.5
cc_77 VPB N_C1_c_320_n 0.00492723f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.505
cc_78 VPB N_VPWR_c_359_n 0.0143271f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.675
cc_79 VPB N_VPWR_c_360_n 0.048246f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=2.465
cc_80 VPB N_VPWR_c_361_n 3.28374e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_362_n 0.00452823f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.505
cc_82 VPB N_VPWR_c_363_n 0.00877349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_364_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_365_n 0.0170192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_366_n 0.0168601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_367_n 0.0585533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_358_n 0.0603153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_369_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_370_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_371_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_135_367#_c_438_n 0.00740227f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.5
cc_92 VPB N_A_135_367#_c_439_n 0.00231254f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.5
cc_93 VPB N_A_135_367#_c_440_n 0.0130663f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.582
cc_94 VPB N_A_727_367#_c_491_n 0.00342647f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=0.765
cc_95 VPB N_A_727_367#_c_492_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.5
cc_96 VPB N_A_727_367#_c_493_n 0.0377269f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_97 VPB N_Y_c_521_n 0.00498917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_Y_c_532_n 0.00710593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 N_A3_M1015_g N_A2_M1005_g 0.0192544f $X=1.03 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A3_M1018_g N_A2_M1002_g 0.0192544f $X=1.03 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A3_c_102_n N_A2_c_148_n 2.12097e-19 $X=0.94 $Y=1.5 $X2=0 $Y2=0
cc_102 N_A3_c_103_n N_A2_c_148_n 0.0192544f $X=1.03 $Y=1.505 $X2=0 $Y2=0
cc_103 N_A3_c_102_n N_A2_c_149_n 0.00950855f $X=0.94 $Y=1.5 $X2=0 $Y2=0
cc_104 N_A3_c_103_n N_A2_c_149_n 2.12097e-19 $X=1.03 $Y=1.505 $X2=0 $Y2=0
cc_105 N_A3_M1013_g N_VPWR_c_360_n 0.0203576f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A3_M1018_g N_VPWR_c_360_n 7.75547e-19 $X=1.03 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A3_c_103_n N_VPWR_c_360_n 0.00183513f $X=1.03 $Y=1.505 $X2=0 $Y2=0
cc_108 N_A3_c_104_n N_VPWR_c_360_n 0.0257689f $X=0.55 $Y=1.582 $X2=0 $Y2=0
cc_109 N_A3_M1013_g N_VPWR_c_361_n 7.42371e-19 $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A3_M1018_g N_VPWR_c_361_n 0.0145847f $X=1.03 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A3_M1013_g N_VPWR_c_364_n 0.00486043f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A3_M1018_g N_VPWR_c_364_n 0.00486043f $X=1.03 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A3_M1013_g N_VPWR_c_358_n 0.00824727f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A3_M1018_g N_VPWR_c_358_n 0.00824727f $X=1.03 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A3_M1018_g N_A_135_367#_c_438_n 0.0129569f $X=1.03 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A3_c_102_n N_A_135_367#_c_438_n 0.0140641f $X=0.94 $Y=1.5 $X2=0 $Y2=0
cc_117 N_A3_M1013_g N_A_135_367#_c_439_n 0.00253514f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A3_c_102_n N_A_135_367#_c_439_n 0.0145237f $X=0.94 $Y=1.5 $X2=0 $Y2=0
cc_119 N_A3_c_103_n N_A_135_367#_c_439_n 0.00261475f $X=1.03 $Y=1.505 $X2=0
+ $Y2=0
cc_120 N_A3_M1014_g N_A_48_69#_c_621_n 0.00354556f $X=0.6 $Y=0.765 $X2=0 $Y2=0
cc_121 N_A3_M1014_g N_A_48_69#_c_622_n 0.0134505f $X=0.6 $Y=0.765 $X2=0 $Y2=0
cc_122 N_A3_M1015_g N_A_48_69#_c_622_n 0.0129554f $X=1.03 $Y=0.765 $X2=0 $Y2=0
cc_123 N_A3_c_103_n N_A_48_69#_c_622_n 0.00357321f $X=1.03 $Y=1.505 $X2=0 $Y2=0
cc_124 N_A3_c_104_n N_A_48_69#_c_622_n 0.0437702f $X=0.55 $Y=1.582 $X2=0 $Y2=0
cc_125 N_A3_c_103_n N_A_48_69#_c_623_n 0.0065941f $X=1.03 $Y=1.505 $X2=0 $Y2=0
cc_126 N_A3_c_104_n N_A_48_69#_c_623_n 0.0219471f $X=0.55 $Y=1.582 $X2=0 $Y2=0
cc_127 N_A3_M1015_g N_A_48_69#_c_624_n 8.28776e-19 $X=1.03 $Y=0.765 $X2=0 $Y2=0
cc_128 N_A3_M1014_g N_VGND_c_663_n 0.0126588f $X=0.6 $Y=0.765 $X2=0 $Y2=0
cc_129 N_A3_M1015_g N_VGND_c_663_n 0.0102767f $X=1.03 $Y=0.765 $X2=0 $Y2=0
cc_130 N_A3_M1015_g N_VGND_c_666_n 0.00400407f $X=1.03 $Y=0.765 $X2=0 $Y2=0
cc_131 N_A3_M1014_g N_VGND_c_669_n 0.00798302f $X=0.6 $Y=0.765 $X2=0 $Y2=0
cc_132 N_A3_M1015_g N_VGND_c_669_n 0.00775088f $X=1.03 $Y=0.765 $X2=0 $Y2=0
cc_133 N_A3_M1014_g N_VGND_c_670_n 0.00400407f $X=0.6 $Y=0.765 $X2=0 $Y2=0
cc_134 N_A3_M1015_g N_A_307_69#_c_732_n 2.32983e-19 $X=1.03 $Y=0.765 $X2=0 $Y2=0
cc_135 N_A2_M1010_g N_A1_M1000_g 0.0306047f $X=1.89 $Y=2.465 $X2=0 $Y2=0
cc_136 A2 N_A1_M1000_g 0.00490542f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_137 A2 N_A1_c_207_n 0.0055887f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_138 A2 N_A1_c_208_n 0.00596328f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A2_c_148_n N_A1_c_208_n 0.00981137f $X=1.89 $Y=1.505 $X2=0 $Y2=0
cc_140 A2 N_A1_M1011_g 2.93669e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_141 A2 N_A1_c_211_n 6.17233e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A2_M1002_g N_VPWR_c_361_n 0.0146036f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A2_M1010_g N_VPWR_c_361_n 7.53251e-19 $X=1.89 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A2_M1010_g N_VPWR_c_362_n 0.00648836f $X=1.89 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A2_M1002_g N_VPWR_c_365_n 0.00486043f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A2_M1010_g N_VPWR_c_365_n 0.0054895f $X=1.89 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A2_M1002_g N_VPWR_c_358_n 0.00824727f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A2_M1010_g N_VPWR_c_358_n 0.0105372f $X=1.89 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A2_M1002_g N_A_135_367#_c_438_n 0.0129569f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A2_M1010_g N_A_135_367#_c_438_n 0.00253514f $X=1.89 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A2_c_148_n N_A_135_367#_c_438_n 0.00261475f $X=1.89 $Y=1.505 $X2=0
+ $Y2=0
cc_152 N_A2_c_149_n N_A_135_367#_c_438_n 0.0286794f $X=1.94 $Y=1.582 $X2=0 $Y2=0
cc_153 N_A2_M1010_g N_A_135_367#_c_450_n 0.0154709f $X=1.89 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A2_c_148_n N_A_135_367#_c_450_n 2.62763e-19 $X=1.89 $Y=1.505 $X2=0
+ $Y2=0
cc_155 N_A2_c_154_n N_A_135_367#_c_450_n 8.80305e-19 $X=2.275 $Y=1.582 $X2=0
+ $Y2=0
cc_156 N_A2_M1010_g N_A_135_367#_c_453_n 8.25449e-19 $X=1.89 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A2_M1010_g N_A_135_367#_c_454_n 0.0113002f $X=1.89 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A2_M1012_g N_Y_c_520_n 8.87163e-19 $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_159 A2 N_Y_c_521_n 0.0268798f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A2_c_148_n N_Y_c_521_n 0.00217335f $X=1.89 $Y=1.505 $X2=0 $Y2=0
cc_161 N_A2_M1012_g N_Y_c_528_n 6.03765e-19 $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_162 A2 N_Y_c_528_n 0.00705895f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_163 N_A2_c_148_n N_Y_c_538_n 0.0016349f $X=1.89 $Y=1.505 $X2=0 $Y2=0
cc_164 N_A2_c_154_n N_Y_c_538_n 0.0529752f $X=2.275 $Y=1.582 $X2=0 $Y2=0
cc_165 N_A2_M1005_g N_A_48_69#_c_624_n 8.28478e-19 $X=1.46 $Y=0.765 $X2=0 $Y2=0
cc_166 N_A2_M1005_g N_A_48_69#_c_625_n 0.0129554f $X=1.46 $Y=0.765 $X2=0 $Y2=0
cc_167 N_A2_M1012_g N_A_48_69#_c_625_n 0.0138953f $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_168 N_A2_c_148_n N_A_48_69#_c_625_n 0.0101463f $X=1.89 $Y=1.505 $X2=0 $Y2=0
cc_169 N_A2_c_154_n N_A_48_69#_c_625_n 0.0288831f $X=2.275 $Y=1.582 $X2=0 $Y2=0
cc_170 N_A2_c_149_n N_A_48_69#_c_625_n 0.0437702f $X=1.94 $Y=1.582 $X2=0 $Y2=0
cc_171 N_A2_M1005_g N_VGND_c_663_n 6.50188e-19 $X=1.46 $Y=0.765 $X2=0 $Y2=0
cc_172 N_A2_M1005_g N_VGND_c_666_n 0.00450424f $X=1.46 $Y=0.765 $X2=0 $Y2=0
cc_173 N_A2_M1012_g N_VGND_c_666_n 0.00291444f $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_174 N_A2_M1005_g N_VGND_c_669_n 0.00862457f $X=1.46 $Y=0.765 $X2=0 $Y2=0
cc_175 N_A2_M1012_g N_VGND_c_669_n 0.00428623f $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_176 N_A2_M1005_g N_A_307_69#_c_734_n 0.00517295f $X=1.46 $Y=0.765 $X2=0 $Y2=0
cc_177 N_A2_M1012_g N_A_307_69#_c_734_n 0.0109596f $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_178 N_A2_M1012_g N_A_307_69#_c_731_n 0.0102482f $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_179 N_A2_M1005_g N_A_307_69#_c_732_n 0.00344817f $X=1.46 $Y=0.765 $X2=0 $Y2=0
cc_180 N_A2_M1012_g N_A_307_69#_c_732_n 0.00159238f $X=1.89 $Y=0.765 $X2=0 $Y2=0
cc_181 N_A1_M1008_g N_B1_M1006_g 0.0181033f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_182 N_A1_c_211_n N_B1_c_279_n 2.84704e-19 $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A1_c_212_n N_B1_c_279_n 0.0218651f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A1_c_211_n N_B1_c_276_n 0.0181033f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A1_c_212_n N_B1_c_276_n 0.00321615f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A1_M1000_g N_VPWR_c_362_n 0.0065171f $X=2.555 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A1_M1000_g N_VPWR_c_363_n 6.59962e-19 $X=2.555 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A1_M1011_g N_VPWR_c_363_n 0.0129895f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A1_M1000_g N_VPWR_c_366_n 0.0054895f $X=2.555 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A1_M1011_g N_VPWR_c_366_n 0.00486043f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A1_M1000_g N_VPWR_c_358_n 0.0105235f $X=2.555 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A1_M1011_g N_VPWR_c_358_n 0.00824727f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A1_M1000_g N_A_135_367#_c_450_n 0.0121441f $X=2.555 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A1_M1000_g N_A_135_367#_c_453_n 0.0102695f $X=2.555 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A1_M1011_g N_A_135_367#_c_440_n 0.0142939f $X=2.985 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A1_M1000_g N_A_135_367#_c_454_n 8.27389e-19 $X=2.555 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A1_M1000_g N_A_135_367#_c_459_n 7.32094e-19 $X=2.555 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A1_M1011_g N_A_727_367#_c_491_n 8.26507e-19 $X=2.985 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A1_M1000_g N_Y_c_521_n 0.00196482f $X=2.555 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A1_c_207_n N_Y_c_521_n 0.00203121f $X=2.91 $Y=1.6 $X2=0 $Y2=0
cc_201 N_A1_M1011_g N_Y_c_521_n 0.00757533f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A1_M1007_g N_Y_c_521_n 0.0030745f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_203 N_A1_M1008_g N_Y_c_521_n 4.43558e-19 $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_204 N_A1_c_211_n N_Y_c_521_n 0.0166271f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_205 N_A1_c_212_n N_Y_c_521_n 0.0201297f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_206 N_A1_M1007_g N_Y_c_522_n 0.00955927f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_207 N_A1_M1008_g N_Y_c_522_n 0.0133191f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_208 N_A1_c_211_n N_Y_c_522_n 0.00252537f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_209 N_A1_c_212_n N_Y_c_522_n 0.0278016f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A1_M1008_g N_Y_c_523_n 8.28478e-19 $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_211 N_A1_c_207_n N_Y_c_528_n 0.00494297f $X=2.91 $Y=1.6 $X2=0 $Y2=0
cc_212 N_A1_M1007_g N_Y_c_528_n 0.0052097f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_213 N_A1_c_212_n N_Y_c_529_n 0.00168673f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_214 N_A1_c_211_n N_Y_c_532_n 0.0077983f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_215 N_A1_c_212_n N_Y_c_532_n 0.0315212f $X=3.455 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A1_M1011_g Y 0.0122062f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A1_M1000_g N_Y_c_538_n 0.0127097f $X=2.555 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A1_c_207_n N_Y_c_538_n 0.00196563f $X=2.91 $Y=1.6 $X2=0 $Y2=0
cc_219 N_A1_M1007_g N_A_48_69#_c_625_n 6.07562e-19 $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_220 N_A1_M1008_g N_VGND_c_664_n 7.54061e-19 $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_221 N_A1_M1007_g N_VGND_c_666_n 0.00302473f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_222 N_A1_M1008_g N_VGND_c_666_n 0.00466675f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_223 N_A1_M1007_g N_VGND_c_669_n 0.00484658f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_224 N_A1_M1008_g N_VGND_c_669_n 0.00898886f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_225 N_A1_M1007_g N_A_307_69#_c_731_n 0.0117119f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_226 N_A1_M1008_g N_A_307_69#_c_731_n 0.00307433f $X=3.545 $Y=0.745 $X2=0
+ $Y2=0
cc_227 N_A1_M1007_g N_A_307_69#_c_741_n 0.0108727f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_228 N_A1_M1008_g N_A_307_69#_c_741_n 0.00509157f $X=3.545 $Y=0.745 $X2=0
+ $Y2=0
cc_229 N_B1_M1017_g N_C1_M1004_g 0.0241477f $X=4.405 $Y=0.745 $X2=0 $Y2=0
cc_230 N_B1_M1019_g N_C1_M1001_g 0.0241477f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_231 N_B1_M1019_g C1 0.0029952f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_232 N_B1_c_279_n C1 0.0260434f $X=4.065 $Y=1.51 $X2=0 $Y2=0
cc_233 N_B1_c_276_n C1 0.00957912f $X=4.405 $Y=1.51 $X2=0 $Y2=0
cc_234 N_B1_c_276_n N_C1_c_320_n 0.0241477f $X=4.405 $Y=1.51 $X2=0 $Y2=0
cc_235 N_B1_M1003_g N_VPWR_c_363_n 0.00555871f $X=3.975 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B1_M1003_g N_VPWR_c_367_n 0.00357877f $X=3.975 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1019_g N_VPWR_c_367_n 0.00357877f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_M1003_g N_VPWR_c_358_n 0.00665089f $X=3.975 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1019_g N_VPWR_c_358_n 0.00537654f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_M1003_g N_A_135_367#_c_440_n 0.0200342f $X=3.975 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_B1_M1003_g N_A_727_367#_c_491_n 0.0112106f $X=3.975 $Y=2.465 $X2=0
+ $Y2=0
cc_242 N_B1_M1019_g N_A_727_367#_c_491_n 0.0153414f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_B1_M1006_g N_Y_c_523_n 8.28776e-19 $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_244 N_B1_M1006_g N_Y_c_524_n 0.0132884f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_245 N_B1_M1017_g N_Y_c_524_n 0.0143319f $X=4.405 $Y=0.745 $X2=0 $Y2=0
cc_246 N_B1_c_279_n N_Y_c_524_n 0.0241876f $X=4.065 $Y=1.51 $X2=0 $Y2=0
cc_247 N_B1_c_276_n N_Y_c_524_n 0.00252537f $X=4.405 $Y=1.51 $X2=0 $Y2=0
cc_248 N_B1_M1017_g N_Y_c_525_n 8.28776e-19 $X=4.405 $Y=0.745 $X2=0 $Y2=0
cc_249 N_B1_M1003_g N_Y_c_532_n 0.0140186f $X=3.975 $Y=2.465 $X2=0 $Y2=0
cc_250 N_B1_M1019_g N_Y_c_532_n 0.0173168f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B1_c_279_n N_Y_c_532_n 0.0228449f $X=4.065 $Y=1.51 $X2=0 $Y2=0
cc_252 N_B1_c_276_n N_Y_c_532_n 7.9609e-19 $X=4.405 $Y=1.51 $X2=0 $Y2=0
cc_253 N_B1_M1006_g N_VGND_c_664_n 0.0106526f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_254 N_B1_M1017_g N_VGND_c_664_n 0.0102222f $X=4.405 $Y=0.745 $X2=0 $Y2=0
cc_255 N_B1_M1017_g N_VGND_c_665_n 5.123e-19 $X=4.405 $Y=0.745 $X2=0 $Y2=0
cc_256 N_B1_M1006_g N_VGND_c_666_n 0.00414769f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_257 N_B1_M1017_g N_VGND_c_667_n 0.00414769f $X=4.405 $Y=0.745 $X2=0 $Y2=0
cc_258 N_B1_M1006_g N_VGND_c_669_n 0.0078848f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_259 N_B1_M1017_g N_VGND_c_669_n 0.0078848f $X=4.405 $Y=0.745 $X2=0 $Y2=0
cc_260 N_C1_M1001_g N_VPWR_c_367_n 0.00357877f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_261 N_C1_M1009_g N_VPWR_c_367_n 0.00357877f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_262 N_C1_M1001_g N_VPWR_c_358_n 0.00537654f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_263 N_C1_M1009_g N_VPWR_c_358_n 0.00626584f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_264 N_C1_M1001_g N_A_727_367#_c_497_n 0.012237f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_265 N_C1_M1009_g N_A_727_367#_c_497_n 0.0120601f $X=5.265 $Y=2.465 $X2=0
+ $Y2=0
cc_266 C1 N_A_727_367#_c_493_n 0.022751f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_267 C1 N_Y_c_524_n 0.00923187f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_268 N_C1_M1004_g N_Y_c_525_n 8.28776e-19 $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_269 N_C1_M1004_g N_Y_c_526_n 0.0133082f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_270 N_C1_M1016_g N_Y_c_526_n 0.0140857f $X=5.265 $Y=0.745 $X2=0 $Y2=0
cc_271 C1 N_Y_c_526_n 0.0742129f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_272 N_C1_c_320_n N_Y_c_526_n 0.00246472f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_273 N_C1_M1016_g N_Y_c_527_n 0.00354659f $X=5.265 $Y=0.745 $X2=0 $Y2=0
cc_274 C1 N_Y_c_530_n 0.0167894f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_275 N_C1_M1001_g N_Y_c_532_n 0.0138576f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_276 C1 N_Y_c_532_n 0.0347909f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_277 N_C1_M1009_g N_Y_c_580_n 0.00820169f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_278 C1 N_Y_c_580_n 0.0190692f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_279 N_C1_c_320_n N_Y_c_580_n 6.52992e-19 $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_280 N_C1_M1004_g N_VGND_c_664_n 5.123e-19 $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_281 N_C1_M1004_g N_VGND_c_665_n 0.0102222f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_282 N_C1_M1016_g N_VGND_c_665_n 0.012533f $X=5.265 $Y=0.745 $X2=0 $Y2=0
cc_283 N_C1_M1004_g N_VGND_c_667_n 0.00414769f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_284 N_C1_M1016_g N_VGND_c_668_n 0.00414769f $X=5.265 $Y=0.745 $X2=0 $Y2=0
cc_285 N_C1_M1004_g N_VGND_c_669_n 0.0078848f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_286 N_C1_M1016_g N_VGND_c_669_n 0.00824082f $X=5.265 $Y=0.745 $X2=0 $Y2=0
cc_287 N_VPWR_c_358_n N_A_135_367#_M1013_d 0.00571434f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_288 N_VPWR_c_358_n N_A_135_367#_M1002_s 0.00380103f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_358_n N_A_135_367#_M1000_d 0.00380103f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_358_n N_A_135_367#_M1003_d 0.00225186f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_364_n N_A_135_367#_c_465_n 0.0120977f $X=1.08 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_358_n N_A_135_367#_c_465_n 0.00691495f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_M1018_s N_A_135_367#_c_438_n 0.00176461f $X=1.105 $Y=1.835 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_361_n N_A_135_367#_c_438_n 0.0170777f $X=1.245 $Y=2.18 $X2=0
+ $Y2=0
cc_295 N_VPWR_M1010_d N_A_135_367#_c_450_n 0.0117692f $X=1.965 $Y=1.835 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_362_n N_A_135_367#_c_450_n 0.0266856f $X=2.225 $Y=2.76 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_362_n N_A_135_367#_c_453_n 0.028341f $X=2.225 $Y=2.76 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_366_n N_A_135_367#_c_453_n 0.015688f $X=3.035 $Y=3.33 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_358_n N_A_135_367#_c_453_n 0.00984745f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_M1011_s N_A_135_367#_c_440_n 0.00503575f $X=3.06 $Y=1.835 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_363_n N_A_135_367#_c_440_n 0.0220026f $X=3.2 $Y=2.76 $X2=0 $Y2=0
cc_302 N_VPWR_c_362_n N_A_135_367#_c_454_n 0.0278473f $X=2.225 $Y=2.76 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_365_n N_A_135_367#_c_454_n 0.015688f $X=2.06 $Y=3.33 $X2=0 $Y2=0
cc_304 N_VPWR_c_358_n N_A_135_367#_c_454_n 0.00984217f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_358_n N_A_727_367#_M1003_s 0.00215176f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_306 N_VPWR_c_358_n N_A_727_367#_M1019_s 0.0022356f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_358_n N_A_727_367#_M1009_d 0.0021516f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_363_n N_A_727_367#_c_491_n 0.0195302f $X=3.2 $Y=2.76 $X2=0 $Y2=0
cc_309 N_VPWR_c_367_n N_A_727_367#_c_491_n 0.0525397f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_358_n N_A_727_367#_c_491_n 0.0324915f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_367_n N_A_727_367#_c_497_n 0.0341772f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_358_n N_A_727_367#_c_497_n 0.0216081f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_367_n N_A_727_367#_c_492_n 0.0186279f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_358_n N_A_727_367#_c_492_n 0.0108858f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_367_n N_A_727_367#_c_510_n 0.0150071f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_358_n N_A_727_367#_c_510_n 0.0101082f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_358_n N_Y_M1001_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_318 N_VPWR_M1011_s N_Y_c_532_n 0.00596908f $X=3.06 $Y=1.835 $X2=0 $Y2=0
cc_319 N_VPWR_M1010_d N_Y_c_538_n 0.0110156f $X=1.965 $Y=1.835 $X2=0 $Y2=0
cc_320 N_A_135_367#_c_440_n N_A_727_367#_M1003_s 0.00607338f $X=4.025 $Y=2.375
+ $X2=-0.19 $Y2=1.655
cc_321 N_A_135_367#_M1003_d N_A_727_367#_c_491_n 0.00337304f $X=4.05 $Y=1.835
+ $X2=0 $Y2=0
cc_322 N_A_135_367#_c_440_n N_A_727_367#_c_491_n 0.0307161f $X=4.025 $Y=2.375
+ $X2=0 $Y2=0
cc_323 N_A_135_367#_M1003_d N_Y_c_532_n 0.00371129f $X=4.05 $Y=1.835 $X2=0 $Y2=0
cc_324 N_A_135_367#_c_440_n N_Y_c_532_n 0.0773713f $X=4.025 $Y=2.375 $X2=0 $Y2=0
cc_325 N_A_135_367#_c_440_n Y 0.0113922f $X=4.025 $Y=2.375 $X2=0 $Y2=0
cc_326 N_A_135_367#_M1000_d N_Y_c_538_n 0.00415747f $X=2.63 $Y=1.835 $X2=0 $Y2=0
cc_327 N_A_135_367#_c_450_n N_Y_c_538_n 0.0380311f $X=2.605 $Y=2.375 $X2=0 $Y2=0
cc_328 N_A_135_367#_c_459_n N_Y_c_538_n 0.0155387f $X=2.77 $Y=2.375 $X2=0 $Y2=0
cc_329 N_A_135_367#_c_438_n N_A_48_69#_c_622_n 0.00156656f $X=1.58 $Y=1.84 $X2=0
+ $Y2=0
cc_330 N_A_135_367#_c_438_n N_A_48_69#_c_625_n 0.00156656f $X=1.58 $Y=1.84 $X2=0
+ $Y2=0
cc_331 N_A_135_367#_c_438_n N_A_48_69#_c_627_n 0.00748144f $X=1.58 $Y=1.84 $X2=0
+ $Y2=0
cc_332 N_A_727_367#_c_497_n N_Y_M1001_s 0.00332344f $X=5.365 $Y=2.99 $X2=0 $Y2=0
cc_333 N_A_727_367#_M1003_s N_Y_c_532_n 0.00685112f $X=3.635 $Y=1.835 $X2=0
+ $Y2=0
cc_334 N_A_727_367#_M1019_s N_Y_c_532_n 0.00355129f $X=4.48 $Y=1.835 $X2=0 $Y2=0
cc_335 N_A_727_367#_c_518_p N_Y_c_532_n 0.0136549f $X=4.62 $Y=2.455 $X2=0 $Y2=0
cc_336 N_A_727_367#_c_497_n N_Y_c_580_n 0.0128826f $X=5.365 $Y=2.99 $X2=0 $Y2=0
cc_337 N_Y_c_520_n N_A_48_69#_c_625_n 5.62116e-19 $X=2.83 $Y=0.68 $X2=0 $Y2=0
cc_338 N_Y_c_528_n N_A_48_69#_c_625_n 0.00995927f $X=2.655 $Y=1.085 $X2=0 $Y2=0
cc_339 N_Y_c_520_n N_A_48_69#_c_626_n 0.0267481f $X=2.83 $Y=0.68 $X2=0 $Y2=0
cc_340 N_Y_c_524_n N_VGND_M1006_s 0.00176461f $X=4.525 $Y=1.17 $X2=0 $Y2=0
cc_341 N_Y_c_526_n N_VGND_M1004_s 0.00176461f $X=5.385 $Y=1.17 $X2=0 $Y2=0
cc_342 N_Y_c_523_n N_VGND_c_664_n 0.0236157f $X=3.76 $Y=0.47 $X2=0 $Y2=0
cc_343 N_Y_c_524_n N_VGND_c_664_n 0.0170777f $X=4.525 $Y=1.17 $X2=0 $Y2=0
cc_344 N_Y_c_525_n N_VGND_c_664_n 0.0236157f $X=4.62 $Y=0.47 $X2=0 $Y2=0
cc_345 N_Y_c_525_n N_VGND_c_665_n 0.0236157f $X=4.62 $Y=0.47 $X2=0 $Y2=0
cc_346 N_Y_c_526_n N_VGND_c_665_n 0.0170777f $X=5.385 $Y=1.17 $X2=0 $Y2=0
cc_347 N_Y_c_527_n N_VGND_c_665_n 0.0236597f $X=5.48 $Y=0.47 $X2=0 $Y2=0
cc_348 N_Y_c_523_n N_VGND_c_666_n 0.0102275f $X=3.76 $Y=0.47 $X2=0 $Y2=0
cc_349 N_Y_c_525_n N_VGND_c_667_n 0.0102275f $X=4.62 $Y=0.47 $X2=0 $Y2=0
cc_350 N_Y_c_527_n N_VGND_c_668_n 0.0151237f $X=5.48 $Y=0.47 $X2=0 $Y2=0
cc_351 N_Y_c_523_n N_VGND_c_669_n 0.00712543f $X=3.76 $Y=0.47 $X2=0 $Y2=0
cc_352 N_Y_c_525_n N_VGND_c_669_n 0.00712543f $X=4.62 $Y=0.47 $X2=0 $Y2=0
cc_353 N_Y_c_527_n N_VGND_c_669_n 0.0105365f $X=5.48 $Y=0.47 $X2=0 $Y2=0
cc_354 N_Y_c_522_n N_A_307_69#_M1007_d 0.00184993f $X=3.665 $Y=1.17 $X2=0 $Y2=0
cc_355 N_Y_M1007_s N_A_307_69#_c_731_n 0.00428784f $X=2.675 $Y=0.325 $X2=0 $Y2=0
cc_356 N_Y_c_520_n N_A_307_69#_c_731_n 0.0248779f $X=2.83 $Y=0.68 $X2=0 $Y2=0
cc_357 N_Y_c_522_n N_A_307_69#_c_731_n 0.00194454f $X=3.665 $Y=1.17 $X2=0 $Y2=0
cc_358 N_Y_c_523_n N_A_307_69#_c_731_n 0.00578498f $X=3.76 $Y=0.47 $X2=0 $Y2=0
cc_359 N_Y_c_528_n N_A_307_69#_c_731_n 8.56591e-19 $X=2.655 $Y=1.085 $X2=0 $Y2=0
cc_360 N_Y_c_522_n N_A_307_69#_c_741_n 0.0156176f $X=3.665 $Y=1.17 $X2=0 $Y2=0
cc_361 N_A_48_69#_c_622_n N_VGND_M1014_d 0.00176461f $X=1.15 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_362 N_A_48_69#_c_621_n N_VGND_c_663_n 0.0225255f $X=0.385 $Y=0.49 $X2=0 $Y2=0
cc_363 N_A_48_69#_c_622_n N_VGND_c_663_n 0.0170777f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_364 N_A_48_69#_c_624_n N_VGND_c_663_n 0.02249f $X=1.245 $Y=0.49 $X2=0 $Y2=0
cc_365 N_A_48_69#_c_624_n N_VGND_c_666_n 0.00932149f $X=1.245 $Y=0.49 $X2=0
+ $Y2=0
cc_366 N_A_48_69#_c_621_n N_VGND_c_669_n 0.00966963f $X=0.385 $Y=0.49 $X2=0
+ $Y2=0
cc_367 N_A_48_69#_c_624_n N_VGND_c_669_n 0.00704609f $X=1.245 $Y=0.49 $X2=0
+ $Y2=0
cc_368 N_A_48_69#_c_621_n N_VGND_c_670_n 0.0127923f $X=0.385 $Y=0.49 $X2=0 $Y2=0
cc_369 N_A_48_69#_c_625_n N_A_307_69#_M1005_d 0.00176461f $X=2.01 $Y=1.16
+ $X2=-0.19 $Y2=-0.245
cc_370 N_A_48_69#_c_625_n N_A_307_69#_c_734_n 0.0170147f $X=2.01 $Y=1.16 $X2=0
+ $Y2=0
cc_371 N_A_48_69#_M1012_s N_A_307_69#_c_731_n 0.00363296f $X=1.965 $Y=0.345
+ $X2=0 $Y2=0
cc_372 N_A_48_69#_c_625_n N_A_307_69#_c_731_n 0.00275981f $X=2.01 $Y=1.16 $X2=0
+ $Y2=0
cc_373 N_A_48_69#_c_626_n N_A_307_69#_c_731_n 0.0249437f $X=2.175 $Y=0.68 $X2=0
+ $Y2=0
cc_374 N_A_48_69#_c_624_n N_A_307_69#_c_732_n 0.0049425f $X=1.245 $Y=0.49 $X2=0
+ $Y2=0
cc_375 N_VGND_c_664_n N_A_307_69#_c_731_n 0.00156784f $X=4.19 $Y=0.45 $X2=0
+ $Y2=0
cc_376 N_VGND_c_666_n N_A_307_69#_c_731_n 0.107949f $X=4.025 $Y=0 $X2=0 $Y2=0
cc_377 N_VGND_c_669_n N_A_307_69#_c_731_n 0.0612531f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_663_n N_A_307_69#_c_732_n 0.00219498f $X=0.815 $Y=0.47 $X2=0
+ $Y2=0
cc_379 N_VGND_c_666_n N_A_307_69#_c_732_n 0.0234016f $X=4.025 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_669_n N_A_307_69#_c_732_n 0.0125857f $X=5.52 $Y=0 $X2=0 $Y2=0
