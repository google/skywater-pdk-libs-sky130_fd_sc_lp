* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sleep_sergate_plv_14 VIRTPWR VPWR SLEEP VPB
X0 VIRTPWR SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=7e+06u l=150000u
X1 VPWR SLEEP VIRTPWR VPB sky130_fd_pr__pfet_01v8_hvt w=7e+06u l=150000u
.ends
