* File: sky130_fd_sc_lp__ebufn_lp2.pex.spice
* Created: Wed Sep  2 09:51:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EBUFN_LP2%A 1 3 6 10 13 15 16 17 18 23
c40 13 0 1.57086e-19 $X=0.69 $Y=0.915
r41 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=0.925
+ $X2=0.71 $Y2=1.295
r42 17 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=0.93 $X2=0.71 $Y2=0.93
r43 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=0.555
+ $X2=0.71 $Y2=0.925
r44 14 23 33.9804 $w=4.55e-07 $l=2.78e-07 $layer=POLY_cond $X=0.647 $Y=1.208
+ $X2=0.647 $Y2=0.93
r45 14 15 38.953 $w=4.55e-07 $l=2.27e-07 $layer=POLY_cond $X=0.647 $Y=1.208
+ $X2=0.647 $Y2=1.435
r46 13 23 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=0.647 $Y=0.915
+ $X2=0.647 $Y2=0.93
r47 6 15 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.545 $Y=2.545
+ $X2=0.545 $Y2=1.435
r48 1 13 24.7927 $w=4.55e-07 $l=1.5e-07 $layer=POLY_cond $X=0.69 $Y=0.765
+ $X2=0.69 $Y2=0.915
r49 1 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.885 $Y=0.765
+ $X2=0.885 $Y2=0.445
r50 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.495 $Y=0.765
+ $X2=0.495 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP2%A_27_47# 1 2 7 8 11 15 18 21 25 29 33 34
+ 36
c68 11 0 1.07755e-19 $X=2.05 $Y=1.175
r69 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.325
+ $Y=1.89 $X2=1.325 $Y2=1.89
r70 31 33 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.325 $Y=1.845
+ $X2=1.325 $Y2=1.89
r71 30 36 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.76
+ $X2=0.28 $Y2=1.76
r72 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.16 $Y=1.76
+ $X2=1.325 $Y2=1.845
r73 29 30 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.16 $Y=1.76
+ $X2=0.445 $Y2=1.76
r74 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.19 $X2=0.28
+ $Y2=2.9
r75 23 36 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=1.845
+ $X2=0.28 $Y2=1.76
r76 23 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.28 $Y=1.845
+ $X2=0.28 $Y2=2.19
r77 19 36 3.24686 $w=2.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.24 $Y=1.675
+ $X2=0.28 $Y2=1.76
r78 19 21 55.5478 $w=2.48e-07 $l=1.205e-06 $layer=LI1_cond $X=0.24 $Y=1.675
+ $X2=0.24 $Y2=0.47
r79 17 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.325 $Y=1.875
+ $X2=1.325 $Y2=1.89
r80 13 18 15.9654 $w=2e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.25 $Y=1.875
+ $X2=2.175 $Y2=1.8
r81 13 15 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.25 $Y=1.875
+ $X2=2.25 $Y2=2.595
r82 9 18 15.9654 $w=2e-07 $l=1.58114e-07 $layer=POLY_cond $X=2.05 $Y=1.725
+ $X2=2.175 $Y2=1.8
r83 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.05 $Y=1.725
+ $X2=2.05 $Y2=1.175
r84 8 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.49 $Y=1.8
+ $X2=1.325 $Y2=1.875
r85 7 18 9.46703 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.975 $Y=1.8 $X2=2.175
+ $Y2=1.8
r86 7 8 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.975 $Y=1.8 $X2=1.49
+ $Y2=1.8
r87 2 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r88 2 25 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r89 1 21 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP2%A_232_231# 1 2 8 9 10 13 17 20 21 23 24 25
+ 30 35 36 37 40
c87 13 0 9.30966e-20 $X=2.525 $Y=0.975
r88 35 36 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.547 $Y=2.495
+ $X2=3.547 $Y2=2.33
r89 32 37 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.64 $Y=1.425
+ $X2=3.56 $Y2=1.34
r90 32 36 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=3.64 $Y=1.425
+ $X2=3.64 $Y2=2.33
r91 28 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=1.255
+ $X2=3.56 $Y2=1.34
r92 28 30 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.56 $Y=1.255
+ $X2=3.56 $Y2=0.975
r93 24 37 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=1.34
+ $X2=3.56 $Y2=1.34
r94 24 25 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=3.395 $Y=1.34
+ $X2=2.35 $Y2=1.34
r95 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=1.255
+ $X2=2.35 $Y2=1.34
r96 22 23 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.265 $Y=0.895
+ $X2=2.265 $Y2=1.255
r97 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.18 $Y=0.81
+ $X2=2.265 $Y2=0.895
r98 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.18 $Y=0.81 $X2=1.49
+ $Y2=0.81
r99 18 40 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.325 $Y=1.32
+ $X2=1.515 $Y2=1.32
r100 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.32 $X2=1.325 $Y2=1.32
r101 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.325 $Y=0.895
+ $X2=1.49 $Y2=0.81
r102 15 17 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.325 $Y=0.895
+ $X2=1.325 $Y2=1.32
r103 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.525 $Y=0.595
+ $X2=2.525 $Y2=0.975
r104 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.45 $Y=0.52
+ $X2=2.525 $Y2=0.595
r105 9 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.45 $Y=0.52
+ $X2=1.59 $Y2=0.52
r106 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.155
+ $X2=1.515 $Y2=1.32
r107 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.515 $Y=0.595
+ $X2=1.59 $Y2=0.52
r108 7 8 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.515 $Y=0.595
+ $X2=1.515 $Y2=1.155
r109 2 35 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=3.395
+ $Y=2.095 $X2=3.535 $Y2=2.495
r110 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.765 $X2=3.56 $Y2=0.975
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP2%TE_B 3 7 11 15 17 18 26
c47 26 0 1.76476e-19 $X=3.27 $Y=1.77
r48 26 27 11.1574 $w=3.24e-07 $l=7.5e-08 $layer=POLY_cond $X=3.27 $Y=1.77
+ $X2=3.345 $Y2=1.77
r49 25 26 46.8611 $w=3.24e-07 $l=3.15e-07 $layer=POLY_cond $X=2.955 $Y=1.77
+ $X2=3.27 $Y2=1.77
r50 23 25 26.034 $w=3.24e-07 $l=1.75e-07 $layer=POLY_cond $X=2.78 $Y=1.77
+ $X2=2.955 $Y2=1.77
r51 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.77 $X2=2.78 $Y2=1.77
r52 21 23 5.95062 $w=3.24e-07 $l=4e-08 $layer=POLY_cond $X=2.74 $Y=1.77 $X2=2.78
+ $Y2=1.77
r53 18 24 7.46177 $w=5.43e-07 $l=3.4e-07 $layer=LI1_cond $X=3.12 $Y=1.877
+ $X2=2.78 $Y2=1.877
r54 17 24 3.07249 $w=5.43e-07 $l=1.4e-07 $layer=LI1_cond $X=2.64 $Y=1.877
+ $X2=2.78 $Y2=1.877
r55 13 27 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.605
+ $X2=3.345 $Y2=1.77
r56 13 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.345 $Y=1.605
+ $X2=3.345 $Y2=0.975
r57 9 26 8.92133 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.935
+ $X2=3.27 $Y2=1.77
r58 9 11 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.27 $Y=1.935
+ $X2=3.27 $Y2=2.595
r59 5 25 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.605
+ $X2=2.955 $Y2=1.77
r60 5 7 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.955 $Y=1.605
+ $X2=2.955 $Y2=0.975
r61 1 21 8.92133 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.935
+ $X2=2.74 $Y2=1.77
r62 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.74 $Y=1.935 $X2=2.74
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP2%VPWR 1 2 11 17 20 21 22 32 33 36
r38 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r40 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r41 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r46 24 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 22 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 22 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 20 29 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.84 $Y=3.33 $X2=2.64
+ $Y2=3.33
r50 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=3.33
+ $X2=3.005 $Y2=3.33
r51 19 32 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.17 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=3.33
+ $X2=3.005 $Y2=3.33
r53 15 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=3.245
+ $X2=3.005 $Y2=3.33
r54 15 17 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.005 $Y=3.245
+ $X2=3.005 $Y2=2.495
r55 11 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19 $X2=0.81
+ $Y2=2.9
r56 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245 $X2=0.81
+ $Y2=3.33
r57 9 14 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r58 2 17 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=2.865
+ $Y=2.095 $X2=3.005 $Y2=2.495
r59 1 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r60 1 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP2%Z 1 2 9 14 16 17 18 26
c31 16 0 1.76476e-19 $X=2.075 $Y=1.95
c32 9 0 9.30966e-20 $X=1.835 $Y=1.24
r33 27 36 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=2.047 $Y=2.302
+ $X2=2.047 $Y2=2.24
r34 26 34 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=2.16 $Y=2.035 $X2=2.16
+ $Y2=2.075
r35 17 18 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.047 $Y=2.405
+ $X2=2.047 $Y2=2.775
r36 17 27 2.70761 $w=4.53e-07 $l=1.03e-07 $layer=LI1_cond $X=2.047 $Y=2.405
+ $X2=2.047 $Y2=2.302
r37 16 36 3.7591 $w=4.53e-07 $l=1.43e-07 $layer=LI1_cond $X=2.047 $Y=2.097
+ $X2=2.047 $Y2=2.24
r38 16 34 3.49812 $w=4.53e-07 $l=2.2e-08 $layer=LI1_cond $X=2.047 $Y=2.097
+ $X2=2.047 $Y2=2.075
r39 16 26 1.15244 $w=2.28e-07 $l=2.3e-08 $layer=LI1_cond $X=2.16 $Y=2.012
+ $X2=2.16 $Y2=2.035
r40 14 16 11.8752 $w=2.28e-07 $l=2.37e-07 $layer=LI1_cond $X=2.16 $Y=1.775
+ $X2=2.16 $Y2=2.012
r41 7 14 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.835 $Y=1.69
+ $X2=2.16 $Y2=1.69
r42 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.835 $Y=1.605
+ $X2=1.835 $Y2=1.24
r43 2 36 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.095 $X2=1.985 $Y2=2.24
r44 1 9 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=1.69
+ $Y=0.965 $X2=1.835 $Y2=1.24
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP2%VGND 1 2 9 13 15 17 22 29 30 33 36
c41 17 0 1.57086e-19 $X=1.055 $Y=0
c42 13 0 1.07755e-19 $X=2.74 $Y=0.91
r43 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r46 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.74
+ $Y2=0
r48 27 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.6
+ $Y2=0
r49 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r50 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r52 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r53 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.74
+ $Y2=0
r54 22 25 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=1.68
+ $Y2=0
r55 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r56 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r58 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.72
+ $Y2=0
r59 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r61 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0
r62 11 13 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0.91
r63 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085 $X2=1.22
+ $Y2=0
r64 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.38
r65 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.765 $X2=2.74 $Y2=0.91
r66 1 9 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.235 $X2=1.22 $Y2=0.38
.ends

