* File: sky130_fd_sc_lp__a22o_2.pex.spice
* Created: Wed Sep  2 09:22:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22O_2%A_94_249# 1 2 3 4 15 19 23 27 29 30 33 36 37
+ 38 39 40 45 47 49 54
c116 54 0 1.99348e-19 $X=0.995 $Y=1.41
c117 38 0 7.77818e-20 $X=2.62 $Y=1.08
r118 54 63 11.2331 $w=2.36e-07 $l=5.5e-08 $layer=POLY_cond $X=0.995 $Y=1.485
+ $X2=1.05 $Y2=1.485
r119 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.41 $X2=0.995 $Y2=1.41
r120 47 58 3.09071 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=3.615 $Y=2.14
+ $X2=3.615 $Y2=2.035
r121 47 49 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=3.615 $Y=2.14
+ $X2=3.615 $Y2=2.475
r122 43 45 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=3.55 $Y=0.995
+ $X2=3.55 $Y2=0.42
r123 40 42 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.72 $Y2=2.035
r124 39 58 3.8266 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.615 $Y2=2.035
r125 39 42 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=2.72 $Y2=2.035
r126 38 56 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.08
+ $X2=2.535 $Y2=1.08
r127 37 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.385 $Y=1.08
+ $X2=3.55 $Y2=0.995
r128 37 38 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.385 $Y=1.08
+ $X2=2.62 $Y2=1.08
r129 36 40 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.535 $Y=1.93
+ $X2=2.62 $Y2=2.035
r130 35 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=1.165
+ $X2=2.535 $Y2=1.08
r131 35 36 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.535 $Y=1.165
+ $X2=2.535 $Y2=1.93
r132 31 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.2 $Y=1.08
+ $X2=2.535 $Y2=1.08
r133 31 33 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=2.2 $Y=0.995
+ $X2=2.2 $Y2=0.42
r134 30 53 14.1263 $w=2.85e-07 $l=4.1225e-07 $layer=LI1_cond $X=1.28 $Y=1.08
+ $X2=1.095 $Y2=1.41
r135 29 31 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=1.08
+ $X2=2.2 $Y2=1.08
r136 29 30 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.035 $Y=1.08
+ $X2=1.28 $Y2=1.08
r137 25 63 13.389 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.05 $Y=1.245
+ $X2=1.05 $Y2=1.485
r138 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.05 $Y=1.245
+ $X2=1.05 $Y2=0.665
r139 21 54 4.08475 $w=2.36e-07 $l=2e-08 $layer=POLY_cond $X=0.975 $Y=1.485
+ $X2=0.995 $Y2=1.485
r140 21 23 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.975 $Y=1.575
+ $X2=0.975 $Y2=2.465
r141 17 21 72.5042 $w=2.36e-07 $l=4.59592e-07 $layer=POLY_cond $X=0.62 $Y=1.245
+ $X2=0.975 $Y2=1.485
r142 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.62 $Y=1.245
+ $X2=0.62 $Y2=0.665
r143 13 17 15.3178 $w=2.36e-07 $l=1.83712e-07 $layer=POLY_cond $X=0.545 $Y=1.395
+ $X2=0.62 $Y2=1.245
r144 13 15 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.545 $Y=1.395
+ $X2=0.545 $Y2=2.465
r145 4 58 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=2.015
r146 4 49 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=2.475
r147 3 42 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=1.835 $X2=2.72 $Y2=2.035
r148 2 45 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.245 $X2=3.55 $Y2=0.42
r149 1 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.245 $X2=2.2 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%A2 3 7 9 12 13
c40 13 0 1.99348e-19 $X=1.535 $Y=1.51
r41 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.51
+ $X2=1.535 $Y2=1.675
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.51
+ $X2=1.535 $Y2=1.345
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.535
+ $Y=1.51 $X2=1.535 $Y2=1.51
r44 9 13 4.10641 $w=4.33e-07 $l=1.55e-07 $layer=LI1_cond $X=1.667 $Y=1.665
+ $X2=1.667 $Y2=1.51
r45 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.625 $Y=0.665
+ $X2=1.625 $Y2=1.345
r46 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.555 $Y=2.465
+ $X2=1.555 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%A1 3 7 9 10 16 17
r35 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.51 $X2=2.16 $Y2=1.51
r36 13 16 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.985 $Y=1.51
+ $X2=2.16 $Y2=1.51
r37 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.15 $Y=1.665
+ $X2=2.15 $Y2=2.035
r38 9 17 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.15 $Y=1.665
+ $X2=2.15 $Y2=1.51
r39 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.675
+ $X2=1.985 $Y2=1.51
r40 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.985 $Y=1.675
+ $X2=1.985 $Y2=2.465
r41 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.345
+ $X2=1.985 $Y2=1.51
r42 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.985 $Y=1.345
+ $X2=1.985 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%B2 3 7 9 12
c33 3 0 5.97839e-20 $X=2.935 $Y=2.465
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.51
+ $X2=2.885 $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.51
+ $X2=2.885 $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.885
+ $Y=1.51 $X2=2.885 $Y2=1.51
r37 9 13 6.68702 $w=4.03e-07 $l=2.35e-07 $layer=LI1_cond $X=3.12 $Y=1.547
+ $X2=2.885 $Y2=1.547
r38 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.975 $Y=0.665
+ $X2=2.975 $Y2=1.345
r39 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.935 $Y=2.465
+ $X2=2.935 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%B1 3 7 9 12 15
c27 15 0 5.97839e-20 $X=3.55 $Y=1.46
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.46 $X2=3.55 $Y2=1.46
r29 12 14 28.0409 $w=3.18e-07 $l=1.85e-07 $layer=POLY_cond $X=3.365 $Y=1.46
+ $X2=3.55 $Y2=1.46
r30 11 12 4.54717 $w=3.18e-07 $l=3e-08 $layer=POLY_cond $X=3.335 $Y=1.46
+ $X2=3.365 $Y2=1.46
r31 9 15 6.56252 $w=3.58e-07 $l=2.05e-07 $layer=LI1_cond $X=3.565 $Y=1.665
+ $X2=3.565 $Y2=1.46
r32 5 12 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.625
+ $X2=3.365 $Y2=1.46
r33 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.365 $Y=1.625
+ $X2=3.365 $Y2=2.465
r34 1 11 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=1.295
+ $X2=3.335 $Y2=1.46
r35 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.335 $Y=1.295
+ $X2=3.335 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%VPWR 1 2 3 10 12 18 24 26 28 33 43 44 50 53
r51 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 41 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 38 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.2 $Y2=3.33
r60 38 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.43 $Y=3.33
+ $X2=1.265 $Y2=3.33
r64 34 36 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.43 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 33 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.2 $Y2=3.33
r66 33 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 29 47 3.95154 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.207 $Y2=3.33
r71 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 28 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=1.265 $Y2=3.33
r73 28 31 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r74 26 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 26 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 22 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=3.245 $X2=2.2
+ $Y2=3.33
r77 22 24 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.2 $Y=3.245 $X2=2.2
+ $Y2=2.765
r78 18 21 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=1.265 $Y=2.005
+ $X2=1.265 $Y2=2.95
r79 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.245
+ $X2=1.265 $Y2=3.33
r80 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.265 $Y=3.245
+ $X2=1.265 $Y2=2.95
r81 12 15 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=0.29 $Y=2.165
+ $X2=0.29 $Y2=2.95
r82 10 47 3.19163 $w=2.5e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.207 $Y2=3.33
r83 10 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.95
r84 3 24 600 $w=1.7e-07 $l=9.97547e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=1.835 $X2=2.2 $Y2=2.765
r85 2 21 400 $w=1.7e-07 $l=1.21776e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.265 $Y2=2.95
r86 2 18 400 $w=1.7e-07 $l=2.87706e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.265 $Y2=2.005
r87 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.95
r88 1 12 400 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%X 1 2 11 15 16 17 18 24 30
r27 22 30 1.40162 $w=3.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.755 $Y=0.88
+ $X2=0.755 $Y2=0.925
r28 18 32 7.13719 $w=3.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.755 $Y=0.945
+ $X2=0.755 $Y2=1.065
r29 18 30 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=0.755 $Y=0.945
+ $X2=0.755 $Y2=0.925
r30 18 22 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=0.755 $Y=0.86
+ $X2=0.755 $Y2=0.88
r31 17 18 9.49987 $w=3.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.755 $Y=0.555
+ $X2=0.755 $Y2=0.86
r32 17 24 4.20486 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.755 $Y=0.555
+ $X2=0.755 $Y2=0.42
r33 15 16 8.63747 $w=3.23e-07 $l=1.7e-07 $layer=LI1_cond $X=0.75 $Y=1.755
+ $X2=0.75 $Y2=1.925
r34 15 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.655 $Y=1.755
+ $X2=0.655 $Y2=1.065
r35 11 13 32.9776 $w=3.23e-07 $l=9.3e-07 $layer=LI1_cond $X=0.767 $Y=1.98
+ $X2=0.767 $Y2=2.91
r36 11 16 1.95029 $w=3.23e-07 $l=5.5e-08 $layer=LI1_cond $X=0.767 $Y=1.98
+ $X2=0.767 $Y2=1.925
r37 2 13 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.91
r38 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=1.98
r39 1 24 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.695
+ $Y=0.245 $X2=0.835 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%A_326_367# 1 2 9 13 15 19 21
r28 17 19 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.15 $Y=2.48 $X2=3.15
+ $Y2=2.485
r29 16 21 3.05049 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.885 $Y=2.395
+ $X2=1.745 $Y2=2.395
r30 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.985 $Y=2.395
+ $X2=3.15 $Y2=2.48
r31 15 16 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.985 $Y=2.395
+ $X2=1.885 $Y2=2.395
r32 11 21 3.46198 $w=2.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.735 $Y=2.48
+ $X2=1.745 $Y2=2.395
r33 11 13 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=1.735 $Y=2.48
+ $X2=1.735 $Y2=2.5
r34 7 21 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=2.31
+ $X2=1.745 $Y2=2.395
r35 7 9 9.2607 $w=2.78e-07 $l=2.25e-07 $layer=LI1_cond $X=1.745 $Y=2.31
+ $X2=1.745 $Y2=2.085
r36 2 19 300 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=2 $X=3.01
+ $Y=1.835 $X2=3.15 $Y2=2.485
r37 1 13 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=1.63
+ $Y=1.835 $X2=1.77 $Y2=2.5
r38 1 9 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.835 $X2=1.77 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_2%VGND 1 2 3 10 12 14 18 22 24 26 33 34 40 43
c48 3 0 7.77818e-20 $X=2.615 $Y=0.245
r49 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r52 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 34 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r54 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 31 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.76
+ $Y2=0
r56 31 33 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.6
+ $Y2=0
r57 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r58 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 27 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.345
+ $Y2=0
r60 27 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.68
+ $Y2=0
r61 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.76
+ $Y2=0
r62 26 29 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=1.68
+ $Y2=0
r63 24 44 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r64 24 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r65 20 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0
r66 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0.37
r67 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.345 $Y=0.085
+ $X2=1.345 $Y2=0
r68 16 18 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.345 $Y=0.085
+ $X2=1.345 $Y2=0.37
r69 15 37 4.16268 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.2 $Y2=0
r70 14 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.345
+ $Y2=0
r71 14 15 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=0.4
+ $Y2=0
r72 10 37 3.12201 $w=2.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.2 $Y2=0
r73 10 12 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.39
r74 3 22 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.615
+ $Y=0.245 $X2=2.76 $Y2=0.37
r75 2 18 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.245 $X2=1.345 $Y2=0.37
r76 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.245 $X2=0.295 $Y2=0.39
.ends

