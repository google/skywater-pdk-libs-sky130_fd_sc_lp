* File: sky130_fd_sc_lp__dlxbn_2.pxi.spice
* Created: Wed Sep  2 09:47:57 2020
* 
x_PM_SKY130_FD_SC_LP__DLXBN_2%D N_D_M1014_g N_D_M1011_g N_D_c_163_n N_D_c_164_n
+ N_D_c_169_n D D N_D_c_166_n PM_SKY130_FD_SC_LP__DLXBN_2%D
x_PM_SKY130_FD_SC_LP__DLXBN_2%GATE_N N_GATE_N_c_196_n N_GATE_N_M1013_g
+ N_GATE_N_M1019_g N_GATE_N_c_198_n N_GATE_N_c_199_n N_GATE_N_c_200_n GATE_N
+ N_GATE_N_c_201_n N_GATE_N_c_202_n PM_SKY130_FD_SC_LP__DLXBN_2%GATE_N
x_PM_SKY130_FD_SC_LP__DLXBN_2%A_214_136# N_A_214_136#_M1013_d
+ N_A_214_136#_M1019_d N_A_214_136#_c_237_n N_A_214_136#_M1010_g
+ N_A_214_136#_M1000_g N_A_214_136#_M1022_g N_A_214_136#_c_239_n
+ N_A_214_136#_M1006_g N_A_214_136#_c_240_n N_A_214_136#_c_241_n
+ N_A_214_136#_c_250_n N_A_214_136#_c_251_n N_A_214_136#_c_242_n
+ N_A_214_136#_c_243_n N_A_214_136#_c_244_n N_A_214_136#_c_245_n
+ PM_SKY130_FD_SC_LP__DLXBN_2%A_214_136#
x_PM_SKY130_FD_SC_LP__DLXBN_2%A_45_136# N_A_45_136#_M1014_s N_A_45_136#_M1011_s
+ N_A_45_136#_c_349_n N_A_45_136#_c_350_n N_A_45_136#_M1001_g
+ N_A_45_136#_c_355_n N_A_45_136#_M1023_g N_A_45_136#_c_351_n
+ N_A_45_136#_c_352_n N_A_45_136#_c_358_n N_A_45_136#_c_359_n
+ N_A_45_136#_c_353_n N_A_45_136#_c_360_n PM_SKY130_FD_SC_LP__DLXBN_2%A_45_136#
x_PM_SKY130_FD_SC_LP__DLXBN_2%A_354_47# N_A_354_47#_M1010_s N_A_354_47#_M1000_s
+ N_A_354_47#_M1020_g N_A_354_47#_M1002_g N_A_354_47#_c_445_n
+ N_A_354_47#_c_434_n N_A_354_47#_c_435_n N_A_354_47#_c_462_n
+ N_A_354_47#_c_439_n N_A_354_47#_c_440_n N_A_354_47#_c_441_n
+ N_A_354_47#_c_442_n N_A_354_47#_c_436_n N_A_354_47#_c_437_n
+ N_A_354_47#_c_444_n PM_SKY130_FD_SC_LP__DLXBN_2%A_354_47#
x_PM_SKY130_FD_SC_LP__DLXBN_2%A_805_21# N_A_805_21#_M1012_d N_A_805_21#_M1016_d
+ N_A_805_21#_M1017_g N_A_805_21#_M1005_g N_A_805_21#_M1018_g
+ N_A_805_21#_M1009_g N_A_805_21#_M1004_g N_A_805_21#_c_550_n
+ N_A_805_21#_M1008_g N_A_805_21#_M1021_g N_A_805_21#_c_552_n
+ N_A_805_21#_M1025_g N_A_805_21#_c_553_n N_A_805_21#_c_554_n
+ N_A_805_21#_c_555_n N_A_805_21#_c_556_n N_A_805_21#_c_577_n
+ N_A_805_21#_c_557_n N_A_805_21#_c_558_n N_A_805_21#_c_578_n
+ N_A_805_21#_c_559_n N_A_805_21#_c_579_n N_A_805_21#_c_560_n
+ N_A_805_21#_c_561_n N_A_805_21#_c_562_n N_A_805_21#_c_706_p
+ N_A_805_21#_c_563_n N_A_805_21#_c_564_n N_A_805_21#_c_565_n
+ N_A_805_21#_c_566_n N_A_805_21#_c_582_n N_A_805_21#_c_652_p
+ N_A_805_21#_c_567_n N_A_805_21#_c_568_n N_A_805_21#_c_569_n
+ N_A_805_21#_c_570_n N_A_805_21#_c_585_n N_A_805_21#_c_586_n
+ N_A_805_21#_c_571_n N_A_805_21#_c_572_n PM_SKY130_FD_SC_LP__DLXBN_2%A_805_21#
x_PM_SKY130_FD_SC_LP__DLXBN_2%A_619_47# N_A_619_47#_M1022_d N_A_619_47#_M1020_d
+ N_A_619_47#_M1012_g N_A_619_47#_M1016_g N_A_619_47#_c_755_n
+ N_A_619_47#_c_741_n N_A_619_47#_c_742_n N_A_619_47#_c_743_n
+ N_A_619_47#_c_734_n N_A_619_47#_c_735_n N_A_619_47#_c_736_n
+ N_A_619_47#_c_737_n N_A_619_47#_c_738_n N_A_619_47#_c_739_n
+ PM_SKY130_FD_SC_LP__DLXBN_2%A_619_47#
x_PM_SKY130_FD_SC_LP__DLXBN_2%A_1138_153# N_A_1138_153#_M1018_s
+ N_A_1138_153#_M1009_s N_A_1138_153#_c_827_n N_A_1138_153#_M1007_g
+ N_A_1138_153#_M1003_g N_A_1138_153#_c_829_n N_A_1138_153#_c_830_n
+ N_A_1138_153#_M1024_g N_A_1138_153#_M1015_g N_A_1138_153#_c_832_n
+ N_A_1138_153#_c_833_n N_A_1138_153#_c_834_n N_A_1138_153#_c_835_n
+ N_A_1138_153#_c_836_n PM_SKY130_FD_SC_LP__DLXBN_2%A_1138_153#
x_PM_SKY130_FD_SC_LP__DLXBN_2%VPWR N_VPWR_M1011_d N_VPWR_M1000_d N_VPWR_M1005_d
+ N_VPWR_M1009_d N_VPWR_M1015_d N_VPWR_M1021_s N_VPWR_c_892_n N_VPWR_c_893_n
+ N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n N_VPWR_c_897_n N_VPWR_c_898_n
+ VPWR N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_901_n N_VPWR_c_902_n
+ N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_905_n N_VPWR_c_906_n N_VPWR_c_907_n
+ N_VPWR_c_908_n N_VPWR_c_891_n PM_SKY130_FD_SC_LP__DLXBN_2%VPWR
x_PM_SKY130_FD_SC_LP__DLXBN_2%Q_N N_Q_N_M1007_s N_Q_N_M1003_s Q_N Q_N Q_N Q_N
+ Q_N N_Q_N_c_1002_n PM_SKY130_FD_SC_LP__DLXBN_2%Q_N
x_PM_SKY130_FD_SC_LP__DLXBN_2%Q N_Q_M1008_d N_Q_M1004_d N_Q_c_1021_n Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DLXBN_2%Q
x_PM_SKY130_FD_SC_LP__DLXBN_2%VGND N_VGND_M1014_d N_VGND_M1010_d N_VGND_M1017_d
+ N_VGND_M1018_d N_VGND_M1024_d N_VGND_M1025_s N_VGND_c_1044_n N_VGND_c_1045_n
+ N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n N_VGND_c_1049_n
+ N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n N_VGND_c_1053_n
+ N_VGND_c_1054_n VGND N_VGND_c_1055_n N_VGND_c_1056_n N_VGND_c_1057_n
+ N_VGND_c_1058_n N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n
+ PM_SKY130_FD_SC_LP__DLXBN_2%VGND
cc_1 VNB N_D_c_163_n 0.0217977f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.21
cc_2 VNB N_D_c_164_n 0.020011f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.715
cc_3 VNB D 0.00759673f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_D_c_166_n 0.0163166f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_5 VNB N_GATE_N_c_196_n 0.0181198f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.21
cc_6 VNB N_GATE_N_M1019_g 0.0143014f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.395
cc_7 VNB N_GATE_N_c_198_n 0.0291649f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_8 VNB N_GATE_N_c_199_n 0.033696f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.88
cc_9 VNB N_GATE_N_c_200_n 0.00990067f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_GATE_N_c_201_n 0.042988f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_11 VNB N_GATE_N_c_202_n 0.00966433f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_12 VNB N_A_214_136#_c_237_n 0.0478158f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.21
cc_13 VNB N_A_214_136#_M1022_g 0.0321797f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_14 VNB N_A_214_136#_c_239_n 0.0325664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_214_136#_c_240_n 0.0213705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_214_136#_c_241_n 0.00975313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_214_136#_c_242_n 0.0165016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_214_136#_c_243_n 0.01793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_214_136#_c_244_n 0.00475675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_214_136#_c_245_n 0.042672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_45_136#_c_349_n 0.0351576f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_22 VNB N_A_45_136#_c_350_n 0.0141248f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.21
cc_23 VNB N_A_45_136#_c_351_n 0.0169061f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_24 VNB N_A_45_136#_c_352_n 0.0286807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_45_136#_c_353_n 0.0161893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_354_47#_M1002_g 0.0227841f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB N_A_354_47#_c_434_n 0.0071735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_354_47#_c_435_n 0.00319793f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.375
cc_29 VNB N_A_354_47#_c_436_n 0.00379772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_354_47#_c_437_n 0.0343064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_805_21#_M1018_g 0.0438901f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_32 VNB N_A_805_21#_M1004_g 0.0106154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_805_21#_c_550_n 0.0179856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_805_21#_M1021_g 0.00146541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_805_21#_c_552_n 0.0215764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_805_21#_c_553_n 0.0202134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_805_21#_c_554_n 0.0116541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_805_21#_c_555_n 0.0283848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_805_21#_c_556_n 0.0114734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_805_21#_c_557_n 0.00121107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_805_21#_c_558_n 0.0164489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_805_21#_c_559_n 0.0107436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_805_21#_c_560_n 0.0119813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_805_21#_c_561_n 0.0198483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_805_21#_c_562_n 0.00563806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_805_21#_c_563_n 0.00115717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_805_21#_c_564_n 0.00136131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_805_21#_c_565_n 0.00182267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_805_21#_c_566_n 0.00890428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_805_21#_c_567_n 0.0155352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_805_21#_c_568_n 0.0452747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_805_21#_c_569_n 0.00299682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_805_21#_c_570_n 0.00517036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_805_21#_c_571_n 0.0550612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_805_21#_c_572_n 0.00886383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_619_47#_c_734_n 0.00729557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_619_47#_c_735_n 0.00411008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_619_47#_c_736_n 0.0161014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_619_47#_c_737_n 0.00156342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_619_47#_c_738_n 0.0292988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_619_47#_c_739_n 0.0207668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1138_153#_c_827_n 0.0186261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1138_153#_M1003_g 0.00162504f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_64 VNB N_A_1138_153#_c_829_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1138_153#_c_830_n 0.018048f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.375
cc_66 VNB N_A_1138_153#_M1015_g 0.0105993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1138_153#_c_832_n 0.00576598f $X=-0.19 $Y=-0.245 $X2=0.68
+ $Y2=1.665
cc_68 VNB N_A_1138_153#_c_833_n 7.9666e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1138_153#_c_834_n 0.00534319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1138_153#_c_835_n 0.0116189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1138_153#_c_836_n 0.0398654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VPWR_c_891_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB Q 0.00204696f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.715
cc_74 VNB Q 0.00107534f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.88
cc_75 VNB N_VGND_c_1044_n 0.0244686f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.665
cc_76 VNB N_VGND_c_1045_n 0.00529921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1046_n 0.0084905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1047_n 0.0086011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1048_n 0.00711089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1049_n 0.0111997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1050_n 0.03987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1051_n 0.0354642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1052_n 0.00631381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1053_n 0.0393725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1054_n 0.00631381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1055_n 0.044037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1056_n 0.0197306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1057_n 0.0165399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1058_n 0.0257546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1059_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1060_n 0.00631381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1061_n 0.450405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_D_M1011_g 0.0254744f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.395
cc_94 VPB N_D_c_164_n 0.00423171f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.715
cc_95 VPB N_D_c_169_n 0.0167996f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.88
cc_96 VPB D 0.00570572f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_97 VPB N_GATE_N_M1019_g 0.0426274f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.395
cc_98 VPB N_A_214_136#_M1000_g 0.0283415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_214_136#_c_239_n 0.0231193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_214_136#_M1006_g 0.0425531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_214_136#_c_241_n 0.00726959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_214_136#_c_250_n 0.032401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_214_136#_c_251_n 0.0149567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_214_136#_c_243_n 0.0157623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_214_136#_c_244_n 0.00254424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_214_136#_c_245_n 0.0126246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_45_136#_c_349_n 0.00107597f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.375
cc_108 VPB N_A_45_136#_c_355_n 0.0783172f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_109 VPB N_A_45_136#_M1023_g 0.0201424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_45_136#_c_352_n 0.019461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_45_136#_c_358_n 0.0270075f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.375
cc_112 VPB N_A_45_136#_c_359_n 0.00607342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_45_136#_c_360_n 0.0401955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_354_47#_M1020_g 0.0213375f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.21
cc_115 VPB N_A_354_47#_c_439_n 0.00190513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_354_47#_c_440_n 0.00508577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_354_47#_c_441_n 0.00225981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_354_47#_c_442_n 0.0295605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_354_47#_c_436_n 0.00393111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_354_47#_c_444_n 0.0157374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_805_21#_M1005_g 0.035411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_805_21#_M1018_g 0.0281743f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.375
cc_123 VPB N_A_805_21#_M1004_g 0.0200373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_805_21#_M1021_g 0.0215219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_805_21#_c_577_n 0.00249134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_805_21#_c_578_n 0.00372484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_805_21#_c_579_n 0.0306223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_805_21#_c_560_n 0.00496188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_805_21#_c_566_n 0.00339569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_805_21#_c_582_n 0.00819791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_805_21#_c_567_n 0.0260177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_805_21#_c_569_n 0.0216135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_805_21#_c_585_n 0.00402953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_805_21#_c_586_n 0.0165144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_619_47#_M1016_g 0.0246695f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_136 VPB N_A_619_47#_c_741_n 0.00297301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_619_47#_c_742_n 0.00160268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_619_47#_c_743_n 0.00209131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_619_47#_c_735_n 0.00531637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_619_47#_c_736_n 0.00296304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_619_47#_c_738_n 0.00759571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_1138_153#_M1003_g 0.0233363f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_143 VPB N_A_1138_153#_M1015_g 0.0202119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_1138_153#_c_833_n 0.0206591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_892_n 0.0246391f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.665
cc_146 VPB N_VPWR_c_893_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_894_n 0.0165524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_895_n 0.0352153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_896_n 0.00275572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_897_n 0.0128916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_898_n 0.0202992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_899_n 0.0378742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_900_n 0.0450458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_901_n 0.0381602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_902_n 0.0182639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_903_n 0.0150267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_904_n 0.0283221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_905_n 0.00631622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_906_n 0.0104886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_907_n 0.00862975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_908_n 0.00516427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_891_n 0.126684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 N_D_c_163_n N_GATE_N_c_196_n 0.0106198f $X=0.545 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_164 D N_GATE_N_M1019_g 0.00509751f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_165 N_D_c_166_n N_GATE_N_M1019_g 0.0506925f $X=0.545 $Y=1.375 $X2=0 $Y2=0
cc_166 D N_GATE_N_c_200_n 0.00176788f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_167 N_D_c_166_n N_GATE_N_c_200_n 0.00976199f $X=0.545 $Y=1.375 $X2=0 $Y2=0
cc_168 N_D_c_163_n N_A_214_136#_c_243_n 2.38257e-19 $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_169 D N_A_214_136#_c_243_n 0.0382872f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_170 N_D_M1011_g N_A_45_136#_c_352_n 0.00544769f $X=0.635 $Y=2.395 $X2=0 $Y2=0
cc_171 N_D_c_163_n N_A_45_136#_c_352_n 0.00507313f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_172 D N_A_45_136#_c_352_n 0.0515816f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_173 N_D_c_166_n N_A_45_136#_c_352_n 0.0162737f $X=0.545 $Y=1.375 $X2=0 $Y2=0
cc_174 N_D_M1011_g N_A_45_136#_c_358_n 0.0125212f $X=0.635 $Y=2.395 $X2=0 $Y2=0
cc_175 D N_A_45_136#_c_358_n 0.0188405f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_176 N_D_c_166_n N_A_45_136#_c_353_n 0.00276578f $X=0.545 $Y=1.375 $X2=0 $Y2=0
cc_177 N_D_M1011_g N_A_45_136#_c_360_n 9.83956e-19 $X=0.635 $Y=2.395 $X2=0 $Y2=0
cc_178 N_D_c_169_n N_A_45_136#_c_360_n 0.003944f $X=0.545 $Y=1.88 $X2=0 $Y2=0
cc_179 D N_A_45_136#_c_360_n 0.00664099f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_180 N_D_M1011_g N_VPWR_c_892_n 0.00988584f $X=0.635 $Y=2.395 $X2=0 $Y2=0
cc_181 N_D_M1011_g N_VPWR_c_904_n 0.00349617f $X=0.635 $Y=2.395 $X2=0 $Y2=0
cc_182 N_D_M1011_g N_VPWR_c_891_n 0.00396651f $X=0.635 $Y=2.395 $X2=0 $Y2=0
cc_183 N_D_c_163_n N_VGND_c_1044_n 0.00340737f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_184 D N_VGND_c_1044_n 0.0174299f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_185 N_D_c_166_n N_VGND_c_1044_n 2.98046e-19 $X=0.545 $Y=1.375 $X2=0 $Y2=0
cc_186 N_D_c_163_n N_VGND_c_1058_n 0.0038748f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_187 N_D_c_163_n N_VGND_c_1061_n 0.00454494f $X=0.545 $Y=1.21 $X2=0 $Y2=0
cc_188 N_GATE_N_c_199_n N_A_214_136#_c_237_n 0.0202107f $X=1.535 $Y=1.21 $X2=0
+ $Y2=0
cc_189 N_GATE_N_c_201_n N_A_214_136#_c_237_n 0.00725133f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_190 N_GATE_N_M1019_g N_A_214_136#_c_240_n 0.00260108f $X=1.065 $Y=2.395 $X2=0
+ $Y2=0
cc_191 N_GATE_N_c_198_n N_A_214_136#_c_240_n 0.0127692f $X=1.46 $Y=1.285 $X2=0
+ $Y2=0
cc_192 N_GATE_N_c_196_n N_A_214_136#_c_243_n 0.00830403f $X=0.995 $Y=1.21 $X2=0
+ $Y2=0
cc_193 N_GATE_N_M1019_g N_A_214_136#_c_243_n 0.0146191f $X=1.065 $Y=2.395 $X2=0
+ $Y2=0
cc_194 N_GATE_N_c_198_n N_A_214_136#_c_243_n 0.0231904f $X=1.46 $Y=1.285 $X2=0
+ $Y2=0
cc_195 N_GATE_N_c_199_n N_A_214_136#_c_243_n 0.0161455f $X=1.535 $Y=1.21 $X2=0
+ $Y2=0
cc_196 N_GATE_N_c_201_n N_A_214_136#_c_243_n 9.34848e-19 $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_197 N_GATE_N_c_202_n N_A_214_136#_c_243_n 0.0338156f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_198 N_GATE_N_M1019_g N_A_45_136#_c_358_n 0.0206238f $X=1.065 $Y=2.395 $X2=0
+ $Y2=0
cc_199 N_GATE_N_c_201_n N_A_354_47#_c_445_n 0.00218246f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_200 N_GATE_N_c_202_n N_A_354_47#_c_445_n 0.0240062f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_201 N_GATE_N_c_199_n N_A_354_47#_c_435_n 0.00431916f $X=1.535 $Y=1.21 $X2=0
+ $Y2=0
cc_202 N_GATE_N_c_202_n N_A_354_47#_c_435_n 0.00204979f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_203 N_GATE_N_M1019_g N_A_354_47#_c_444_n 0.00847689f $X=1.065 $Y=2.395 $X2=0
+ $Y2=0
cc_204 N_GATE_N_M1019_g N_VPWR_c_892_n 0.0175735f $X=1.065 $Y=2.395 $X2=0 $Y2=0
cc_205 N_GATE_N_M1019_g N_VPWR_c_899_n 0.00349617f $X=1.065 $Y=2.395 $X2=0 $Y2=0
cc_206 N_GATE_N_M1019_g N_VPWR_c_891_n 0.00396651f $X=1.065 $Y=2.395 $X2=0 $Y2=0
cc_207 N_GATE_N_c_196_n N_VGND_c_1044_n 0.00159683f $X=0.995 $Y=1.21 $X2=0 $Y2=0
cc_208 N_GATE_N_c_201_n N_VGND_c_1044_n 0.00348299f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_209 N_GATE_N_c_202_n N_VGND_c_1044_n 0.0215698f $X=1.445 $Y=0.405 $X2=0 $Y2=0
cc_210 N_GATE_N_c_196_n N_VGND_c_1051_n 0.0038748f $X=0.995 $Y=1.21 $X2=0 $Y2=0
cc_211 N_GATE_N_c_201_n N_VGND_c_1051_n 0.00604998f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_212 N_GATE_N_c_202_n N_VGND_c_1051_n 0.0227751f $X=1.445 $Y=0.405 $X2=0 $Y2=0
cc_213 N_GATE_N_c_196_n N_VGND_c_1061_n 0.00454494f $X=0.995 $Y=1.21 $X2=0 $Y2=0
cc_214 N_GATE_N_c_201_n N_VGND_c_1061_n 0.00762569f $X=1.445 $Y=0.405 $X2=0
+ $Y2=0
cc_215 N_GATE_N_c_202_n N_VGND_c_1061_n 0.0166253f $X=1.445 $Y=0.405 $X2=0 $Y2=0
cc_216 N_A_214_136#_c_237_n N_A_45_136#_c_349_n 0.031722f $X=2.11 $Y=0.73 $X2=0
+ $Y2=0
cc_217 N_A_214_136#_M1022_g N_A_45_136#_c_349_n 0.00739727f $X=3.02 $Y=0.445
+ $X2=0 $Y2=0
cc_218 N_A_214_136#_c_242_n N_A_45_136#_c_349_n 0.0200311f $X=2.935 $Y=1.17
+ $X2=0 $Y2=0
cc_219 N_A_214_136#_c_243_n N_A_45_136#_c_349_n 0.00625171f $X=1.615 $Y=1.17
+ $X2=0 $Y2=0
cc_220 N_A_214_136#_c_244_n N_A_45_136#_c_349_n 0.00145765f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_221 N_A_214_136#_c_245_n N_A_45_136#_c_349_n 0.026688f $X=2.995 $Y=1.25 $X2=0
+ $Y2=0
cc_222 N_A_214_136#_c_237_n N_A_45_136#_c_350_n 0.0172601f $X=2.11 $Y=0.73 $X2=0
+ $Y2=0
cc_223 N_A_214_136#_M1022_g N_A_45_136#_c_350_n 0.049778f $X=3.02 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_214_136#_c_241_n N_A_45_136#_c_355_n 0.0205259f $X=1.985 $Y=1.635
+ $X2=0 $Y2=0
cc_225 N_A_214_136#_c_250_n N_A_45_136#_c_355_n 0.00885584f $X=2.112 $Y=2.145
+ $X2=0 $Y2=0
cc_226 N_A_214_136#_c_251_n N_A_45_136#_c_355_n 0.00977373f $X=2.112 $Y=2.295
+ $X2=0 $Y2=0
cc_227 N_A_214_136#_c_242_n N_A_45_136#_c_355_n 0.00401735f $X=2.935 $Y=1.17
+ $X2=0 $Y2=0
cc_228 N_A_214_136#_c_243_n N_A_45_136#_c_355_n 0.00242567f $X=1.615 $Y=1.17
+ $X2=0 $Y2=0
cc_229 N_A_214_136#_c_245_n N_A_45_136#_c_355_n 0.00737532f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_230 N_A_214_136#_M1000_g N_A_45_136#_M1023_g 0.0170704f $X=2.15 $Y=2.775
+ $X2=0 $Y2=0
cc_231 N_A_214_136#_c_237_n N_A_45_136#_c_351_n 0.0083414f $X=2.11 $Y=0.73 $X2=0
+ $Y2=0
cc_232 N_A_214_136#_c_242_n N_A_45_136#_c_351_n 0.00430684f $X=2.935 $Y=1.17
+ $X2=0 $Y2=0
cc_233 N_A_214_136#_M1019_d N_A_45_136#_c_358_n 0.0196876f $X=1.14 $Y=2.075
+ $X2=0 $Y2=0
cc_234 N_A_214_136#_M1000_g N_A_45_136#_c_358_n 0.00363223f $X=2.15 $Y=2.775
+ $X2=0 $Y2=0
cc_235 N_A_214_136#_c_241_n N_A_45_136#_c_358_n 6.29725e-19 $X=1.985 $Y=1.635
+ $X2=0 $Y2=0
cc_236 N_A_214_136#_c_251_n N_A_45_136#_c_358_n 0.0125673f $X=2.112 $Y=2.295
+ $X2=0 $Y2=0
cc_237 N_A_214_136#_c_243_n N_A_45_136#_c_358_n 0.0726051f $X=1.615 $Y=1.17
+ $X2=0 $Y2=0
cc_238 N_A_214_136#_c_241_n N_A_45_136#_c_359_n 3.51413e-19 $X=1.985 $Y=1.635
+ $X2=0 $Y2=0
cc_239 N_A_214_136#_c_250_n N_A_45_136#_c_359_n 0.00118364f $X=2.112 $Y=2.145
+ $X2=0 $Y2=0
cc_240 N_A_214_136#_c_242_n N_A_45_136#_c_359_n 0.0203452f $X=2.935 $Y=1.17
+ $X2=0 $Y2=0
cc_241 N_A_214_136#_c_243_n N_A_45_136#_c_359_n 0.0208455f $X=1.615 $Y=1.17
+ $X2=0 $Y2=0
cc_242 N_A_214_136#_c_244_n N_A_45_136#_c_359_n 0.00992286f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_243 N_A_214_136#_c_245_n N_A_45_136#_c_359_n 8.81898e-19 $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_244 N_A_214_136#_M1006_g N_A_354_47#_M1020_g 0.0107719f $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_245 N_A_214_136#_M1022_g N_A_354_47#_M1002_g 0.0190576f $X=3.02 $Y=0.445
+ $X2=0 $Y2=0
cc_246 N_A_214_136#_c_237_n N_A_354_47#_c_445_n 0.00500058f $X=2.11 $Y=0.73
+ $X2=0 $Y2=0
cc_247 N_A_214_136#_c_237_n N_A_354_47#_c_434_n 0.00900697f $X=2.11 $Y=0.73
+ $X2=0 $Y2=0
cc_248 N_A_214_136#_M1022_g N_A_354_47#_c_434_n 0.0120444f $X=3.02 $Y=0.445
+ $X2=0 $Y2=0
cc_249 N_A_214_136#_c_239_n N_A_354_47#_c_434_n 0.003898f $X=3.695 $Y=1.59 $X2=0
+ $Y2=0
cc_250 N_A_214_136#_c_242_n N_A_354_47#_c_434_n 0.0586706f $X=2.935 $Y=1.17
+ $X2=0 $Y2=0
cc_251 N_A_214_136#_c_243_n N_A_354_47#_c_434_n 0.0104071f $X=1.615 $Y=1.17
+ $X2=0 $Y2=0
cc_252 N_A_214_136#_c_244_n N_A_354_47#_c_434_n 0.0219834f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_253 N_A_214_136#_c_245_n N_A_354_47#_c_434_n 9.47341e-19 $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_254 N_A_214_136#_c_237_n N_A_354_47#_c_435_n 0.00514392f $X=2.11 $Y=0.73
+ $X2=0 $Y2=0
cc_255 N_A_214_136#_c_243_n N_A_354_47#_c_435_n 0.0235226f $X=1.615 $Y=1.17
+ $X2=0 $Y2=0
cc_256 N_A_214_136#_M1000_g N_A_354_47#_c_462_n 0.00976509f $X=2.15 $Y=2.775
+ $X2=0 $Y2=0
cc_257 N_A_214_136#_c_239_n N_A_354_47#_c_440_n 0.00122064f $X=3.695 $Y=1.59
+ $X2=0 $Y2=0
cc_258 N_A_214_136#_M1006_g N_A_354_47#_c_440_n 0.00173152f $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_259 N_A_214_136#_c_244_n N_A_354_47#_c_440_n 0.00735921f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_260 N_A_214_136#_c_245_n N_A_354_47#_c_440_n 4.44763e-19 $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_261 N_A_214_136#_c_244_n N_A_354_47#_c_441_n 0.0124907f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_262 N_A_214_136#_c_245_n N_A_354_47#_c_441_n 0.00131017f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_263 N_A_214_136#_M1006_g N_A_354_47#_c_442_n 0.0195821f $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_264 N_A_214_136#_c_244_n N_A_354_47#_c_442_n 2.17072e-19 $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_265 N_A_214_136#_c_245_n N_A_354_47#_c_442_n 0.022397f $X=2.995 $Y=1.25 $X2=0
+ $Y2=0
cc_266 N_A_214_136#_M1022_g N_A_354_47#_c_436_n 0.00202319f $X=3.02 $Y=0.445
+ $X2=0 $Y2=0
cc_267 N_A_214_136#_c_239_n N_A_354_47#_c_436_n 0.0226266f $X=3.695 $Y=1.59
+ $X2=0 $Y2=0
cc_268 N_A_214_136#_M1006_g N_A_354_47#_c_436_n 0.00451918f $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_269 N_A_214_136#_c_244_n N_A_354_47#_c_436_n 0.0623909f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_270 N_A_214_136#_c_245_n N_A_354_47#_c_436_n 0.00164068f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_271 N_A_214_136#_M1022_g N_A_354_47#_c_437_n 0.0105835f $X=3.02 $Y=0.445
+ $X2=0 $Y2=0
cc_272 N_A_214_136#_c_239_n N_A_354_47#_c_437_n 0.0193933f $X=3.695 $Y=1.59
+ $X2=0 $Y2=0
cc_273 N_A_214_136#_c_244_n N_A_354_47#_c_437_n 0.001481f $X=2.995 $Y=1.25 $X2=0
+ $Y2=0
cc_274 N_A_214_136#_c_245_n N_A_354_47#_c_437_n 0.00624125f $X=2.995 $Y=1.25
+ $X2=0 $Y2=0
cc_275 N_A_214_136#_M1000_g N_A_354_47#_c_444_n 0.00766049f $X=2.15 $Y=2.775
+ $X2=0 $Y2=0
cc_276 N_A_214_136#_c_251_n N_A_354_47#_c_444_n 3.75142e-19 $X=2.112 $Y=2.295
+ $X2=0 $Y2=0
cc_277 N_A_214_136#_M1006_g N_A_805_21#_c_577_n 2.39957e-19 $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_278 N_A_214_136#_c_239_n N_A_805_21#_c_557_n 3.26215e-19 $X=3.695 $Y=1.59
+ $X2=0 $Y2=0
cc_279 N_A_214_136#_c_239_n N_A_805_21#_c_558_n 0.047185f $X=3.695 $Y=1.59 $X2=0
+ $Y2=0
cc_280 N_A_214_136#_M1006_g N_A_805_21#_c_586_n 0.047185f $X=3.77 $Y=2.665 $X2=0
+ $Y2=0
cc_281 N_A_214_136#_M1006_g N_A_619_47#_c_741_n 0.00648594f $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_282 N_A_214_136#_c_239_n N_A_619_47#_c_742_n 0.00176671f $X=3.695 $Y=1.59
+ $X2=0 $Y2=0
cc_283 N_A_214_136#_M1006_g N_A_619_47#_c_742_n 0.0131841f $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_284 N_A_214_136#_c_239_n N_A_619_47#_c_743_n 4.11197e-19 $X=3.695 $Y=1.59
+ $X2=0 $Y2=0
cc_285 N_A_214_136#_c_239_n N_A_619_47#_c_735_n 0.00911424f $X=3.695 $Y=1.59
+ $X2=0 $Y2=0
cc_286 N_A_214_136#_M1006_g N_A_619_47#_c_735_n 0.0121086f $X=3.77 $Y=2.665
+ $X2=0 $Y2=0
cc_287 N_A_214_136#_M1000_g N_VPWR_c_893_n 0.00591224f $X=2.15 $Y=2.775 $X2=0
+ $Y2=0
cc_288 N_A_214_136#_M1000_g N_VPWR_c_899_n 0.00419017f $X=2.15 $Y=2.775 $X2=0
+ $Y2=0
cc_289 N_A_214_136#_M1006_g N_VPWR_c_900_n 0.00517164f $X=3.77 $Y=2.665 $X2=0
+ $Y2=0
cc_290 N_A_214_136#_M1000_g N_VPWR_c_891_n 0.00782163f $X=2.15 $Y=2.775 $X2=0
+ $Y2=0
cc_291 N_A_214_136#_M1006_g N_VPWR_c_891_n 0.00519032f $X=3.77 $Y=2.665 $X2=0
+ $Y2=0
cc_292 N_A_214_136#_c_237_n N_VGND_c_1045_n 0.00450413f $X=2.11 $Y=0.73 $X2=0
+ $Y2=0
cc_293 N_A_214_136#_c_237_n N_VGND_c_1051_n 0.00427248f $X=2.11 $Y=0.73 $X2=0
+ $Y2=0
cc_294 N_A_214_136#_M1022_g N_VGND_c_1055_n 0.0042361f $X=3.02 $Y=0.445 $X2=0
+ $Y2=0
cc_295 N_A_214_136#_c_237_n N_VGND_c_1061_n 0.00743109f $X=2.11 $Y=0.73 $X2=0
+ $Y2=0
cc_296 N_A_214_136#_M1022_g N_VGND_c_1061_n 0.0062231f $X=3.02 $Y=0.445 $X2=0
+ $Y2=0
cc_297 N_A_214_136#_c_243_n N_VGND_c_1061_n 0.00295661f $X=1.615 $Y=1.17 $X2=0
+ $Y2=0
cc_298 N_A_45_136#_M1023_g N_A_354_47#_M1020_g 0.0328299f $X=2.87 $Y=2.775 $X2=0
+ $Y2=0
cc_299 N_A_45_136#_c_350_n N_A_354_47#_c_445_n 8.06329e-19 $X=2.66 $Y=0.73 $X2=0
+ $Y2=0
cc_300 N_A_45_136#_c_350_n N_A_354_47#_c_434_n 0.00733797f $X=2.66 $Y=0.73 $X2=0
+ $Y2=0
cc_301 N_A_45_136#_c_351_n N_A_354_47#_c_434_n 0.00853354f $X=2.66 $Y=0.805
+ $X2=0 $Y2=0
cc_302 N_A_45_136#_c_355_n N_A_354_47#_c_462_n 0.00203795f $X=2.87 $Y=2.295
+ $X2=0 $Y2=0
cc_303 N_A_45_136#_M1023_g N_A_354_47#_c_462_n 0.0154473f $X=2.87 $Y=2.775 $X2=0
+ $Y2=0
cc_304 N_A_45_136#_c_358_n N_A_354_47#_c_462_n 0.0481441f $X=2.435 $Y=2.24 $X2=0
+ $Y2=0
cc_305 N_A_45_136#_c_355_n N_A_354_47#_c_439_n 0.00153319f $X=2.87 $Y=2.295
+ $X2=0 $Y2=0
cc_306 N_A_45_136#_M1023_g N_A_354_47#_c_439_n 0.00811312f $X=2.87 $Y=2.775
+ $X2=0 $Y2=0
cc_307 N_A_45_136#_c_358_n N_A_354_47#_c_439_n 0.00806515f $X=2.435 $Y=2.24
+ $X2=0 $Y2=0
cc_308 N_A_45_136#_c_355_n N_A_354_47#_c_441_n 0.00358092f $X=2.87 $Y=2.295
+ $X2=0 $Y2=0
cc_309 N_A_45_136#_c_358_n N_A_354_47#_c_441_n 0.00550842f $X=2.435 $Y=2.24
+ $X2=0 $Y2=0
cc_310 N_A_45_136#_c_359_n N_A_354_47#_c_441_n 0.0159432f $X=2.525 $Y=1.79 $X2=0
+ $Y2=0
cc_311 N_A_45_136#_c_355_n N_A_354_47#_c_442_n 0.0376891f $X=2.87 $Y=2.295 $X2=0
+ $Y2=0
cc_312 N_A_45_136#_c_355_n N_A_354_47#_c_436_n 9.88848e-19 $X=2.87 $Y=2.295
+ $X2=0 $Y2=0
cc_313 N_A_45_136#_c_359_n N_A_354_47#_c_436_n 0.00691128f $X=2.525 $Y=1.79
+ $X2=0 $Y2=0
cc_314 N_A_45_136#_M1023_g N_A_354_47#_c_444_n 7.57809e-19 $X=2.87 $Y=2.775
+ $X2=0 $Y2=0
cc_315 N_A_45_136#_c_358_n N_A_354_47#_c_444_n 0.0243113f $X=2.435 $Y=2.24 $X2=0
+ $Y2=0
cc_316 N_A_45_136#_M1023_g N_A_619_47#_c_741_n 0.00164123f $X=2.87 $Y=2.775
+ $X2=0 $Y2=0
cc_317 N_A_45_136#_c_358_n N_VPWR_M1011_d 0.0045589f $X=2.435 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_318 N_A_45_136#_c_358_n N_VPWR_c_892_n 0.0170777f $X=2.435 $Y=2.24 $X2=0
+ $Y2=0
cc_319 N_A_45_136#_c_360_n N_VPWR_c_892_n 0.00946338f $X=0.32 $Y=2.24 $X2=0
+ $Y2=0
cc_320 N_A_45_136#_M1023_g N_VPWR_c_893_n 0.00689433f $X=2.87 $Y=2.775 $X2=0
+ $Y2=0
cc_321 N_A_45_136#_M1023_g N_VPWR_c_900_n 0.00429451f $X=2.87 $Y=2.775 $X2=0
+ $Y2=0
cc_322 N_A_45_136#_c_360_n N_VPWR_c_904_n 0.00881807f $X=0.32 $Y=2.24 $X2=0
+ $Y2=0
cc_323 N_A_45_136#_M1023_g N_VPWR_c_891_n 0.0065462f $X=2.87 $Y=2.775 $X2=0
+ $Y2=0
cc_324 N_A_45_136#_c_360_n N_VPWR_c_891_n 0.0125978f $X=0.32 $Y=2.24 $X2=0 $Y2=0
cc_325 N_A_45_136#_c_350_n N_VGND_c_1045_n 0.00450413f $X=2.66 $Y=0.73 $X2=0
+ $Y2=0
cc_326 N_A_45_136#_c_351_n N_VGND_c_1045_n 5.90728e-19 $X=2.66 $Y=0.805 $X2=0
+ $Y2=0
cc_327 N_A_45_136#_c_350_n N_VGND_c_1055_n 0.0042361f $X=2.66 $Y=0.73 $X2=0
+ $Y2=0
cc_328 N_A_45_136#_c_353_n N_VGND_c_1058_n 0.00568364f $X=0.35 $Y=0.875 $X2=0
+ $Y2=0
cc_329 N_A_45_136#_c_350_n N_VGND_c_1061_n 0.005967f $X=2.66 $Y=0.73 $X2=0 $Y2=0
cc_330 N_A_45_136#_c_353_n N_VGND_c_1061_n 0.0104907f $X=0.35 $Y=0.875 $X2=0
+ $Y2=0
cc_331 N_A_354_47#_M1002_g N_A_805_21#_c_553_n 0.0227787f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_332 N_A_354_47#_c_437_n N_A_805_21#_c_554_n 0.00182696f $X=3.535 $Y=1.02
+ $X2=0 $Y2=0
cc_333 N_A_354_47#_c_436_n N_A_805_21#_c_555_n 6.02025e-19 $X=3.535 $Y=1.02
+ $X2=0 $Y2=0
cc_334 N_A_354_47#_c_437_n N_A_805_21#_c_555_n 0.00764169f $X=3.535 $Y=1.02
+ $X2=0 $Y2=0
cc_335 N_A_354_47#_c_434_n N_A_619_47#_M1022_d 0.00349126f $X=3.38 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_336 N_A_354_47#_M1002_g N_A_619_47#_c_755_n 0.0133598f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_337 N_A_354_47#_c_434_n N_A_619_47#_c_755_n 0.0296077f $X=3.38 $Y=0.71 $X2=0
+ $Y2=0
cc_338 N_A_354_47#_c_437_n N_A_619_47#_c_755_n 5.96694e-19 $X=3.535 $Y=1.02
+ $X2=0 $Y2=0
cc_339 N_A_354_47#_M1020_g N_A_619_47#_c_741_n 0.00858091f $X=3.23 $Y=2.775
+ $X2=0 $Y2=0
cc_340 N_A_354_47#_c_440_n N_A_619_47#_c_742_n 8.06796e-19 $X=3.38 $Y=2.092
+ $X2=0 $Y2=0
cc_341 N_A_354_47#_M1020_g N_A_619_47#_c_743_n 0.00304709f $X=3.23 $Y=2.775
+ $X2=0 $Y2=0
cc_342 N_A_354_47#_c_439_n N_A_619_47#_c_743_n 0.00654547f $X=3.015 $Y=2.495
+ $X2=0 $Y2=0
cc_343 N_A_354_47#_c_440_n N_A_619_47#_c_743_n 0.0292269f $X=3.38 $Y=2.092 $X2=0
+ $Y2=0
cc_344 N_A_354_47#_c_442_n N_A_619_47#_c_743_n 0.00458407f $X=3.32 $Y=2.13 $X2=0
+ $Y2=0
cc_345 N_A_354_47#_M1002_g N_A_619_47#_c_734_n 0.0055153f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_346 N_A_354_47#_c_434_n N_A_619_47#_c_734_n 0.0135453f $X=3.38 $Y=0.71 $X2=0
+ $Y2=0
cc_347 N_A_354_47#_c_436_n N_A_619_47#_c_734_n 0.018965f $X=3.535 $Y=1.02 $X2=0
+ $Y2=0
cc_348 N_A_354_47#_c_437_n N_A_619_47#_c_734_n 0.00164161f $X=3.535 $Y=1.02
+ $X2=0 $Y2=0
cc_349 N_A_354_47#_M1020_g N_A_619_47#_c_735_n 4.62241e-19 $X=3.23 $Y=2.775
+ $X2=0 $Y2=0
cc_350 N_A_354_47#_c_440_n N_A_619_47#_c_735_n 0.0205977f $X=3.38 $Y=2.092 $X2=0
+ $Y2=0
cc_351 N_A_354_47#_c_442_n N_A_619_47#_c_735_n 6.47686e-19 $X=3.32 $Y=2.13 $X2=0
+ $Y2=0
cc_352 N_A_354_47#_c_436_n N_A_619_47#_c_735_n 0.0537729f $X=3.535 $Y=1.02 $X2=0
+ $Y2=0
cc_353 N_A_354_47#_c_436_n N_A_619_47#_c_737_n 0.0141883f $X=3.535 $Y=1.02 $X2=0
+ $Y2=0
cc_354 N_A_354_47#_c_437_n N_A_619_47#_c_737_n 0.00121729f $X=3.535 $Y=1.02
+ $X2=0 $Y2=0
cc_355 N_A_354_47#_c_462_n N_VPWR_M1000_d 0.011699f $X=2.93 $Y=2.58 $X2=0 $Y2=0
cc_356 N_A_354_47#_c_462_n N_VPWR_c_893_n 0.0252358f $X=2.93 $Y=2.58 $X2=0 $Y2=0
cc_357 N_A_354_47#_c_444_n N_VPWR_c_893_n 0.0142983f $X=1.935 $Y=2.61 $X2=0
+ $Y2=0
cc_358 N_A_354_47#_c_462_n N_VPWR_c_899_n 0.00335527f $X=2.93 $Y=2.58 $X2=0
+ $Y2=0
cc_359 N_A_354_47#_c_444_n N_VPWR_c_899_n 0.0208264f $X=1.935 $Y=2.61 $X2=0
+ $Y2=0
cc_360 N_A_354_47#_M1020_g N_VPWR_c_900_n 0.0054895f $X=3.23 $Y=2.775 $X2=0
+ $Y2=0
cc_361 N_A_354_47#_c_462_n N_VPWR_c_900_n 0.00619062f $X=2.93 $Y=2.58 $X2=0
+ $Y2=0
cc_362 N_A_354_47#_M1000_s N_VPWR_c_891_n 0.00215158f $X=1.81 $Y=2.455 $X2=0
+ $Y2=0
cc_363 N_A_354_47#_M1020_g N_VPWR_c_891_n 0.0111524f $X=3.23 $Y=2.775 $X2=0
+ $Y2=0
cc_364 N_A_354_47#_c_462_n N_VPWR_c_891_n 0.0190748f $X=2.93 $Y=2.58 $X2=0 $Y2=0
cc_365 N_A_354_47#_c_444_n N_VPWR_c_891_n 0.0125165f $X=1.935 $Y=2.61 $X2=0
+ $Y2=0
cc_366 N_A_354_47#_c_462_n A_589_491# 0.0018152f $X=2.93 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_367 N_A_354_47#_c_434_n N_VGND_M1010_d 0.00291642f $X=3.38 $Y=0.71 $X2=0
+ $Y2=0
cc_368 N_A_354_47#_c_434_n N_VGND_c_1045_n 0.0217336f $X=3.38 $Y=0.71 $X2=0
+ $Y2=0
cc_369 N_A_354_47#_c_445_n N_VGND_c_1051_n 0.014234f $X=1.895 $Y=0.445 $X2=0
+ $Y2=0
cc_370 N_A_354_47#_c_434_n N_VGND_c_1051_n 0.00259169f $X=3.38 $Y=0.71 $X2=0
+ $Y2=0
cc_371 N_A_354_47#_M1002_g N_VGND_c_1055_n 0.00357877f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_372 N_A_354_47#_c_434_n N_VGND_c_1055_n 0.00876875f $X=3.38 $Y=0.71 $X2=0
+ $Y2=0
cc_373 N_A_354_47#_M1010_s N_VGND_c_1061_n 0.00254447f $X=1.77 $Y=0.235 $X2=0
+ $Y2=0
cc_374 N_A_354_47#_M1002_g N_VGND_c_1061_n 0.00598834f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_375 N_A_354_47#_c_445_n N_VGND_c_1061_n 0.0101374f $X=1.895 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_A_354_47#_c_434_n N_VGND_c_1061_n 0.0219364f $X=3.38 $Y=0.71 $X2=0
+ $Y2=0
cc_377 N_A_354_47#_c_434_n A_547_47# 0.00165214f $X=3.38 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_378 N_A_805_21#_M1005_g N_A_619_47#_M1016_g 0.00660083f $X=4.13 $Y=2.665
+ $X2=0 $Y2=0
cc_379 N_A_805_21#_c_557_n N_A_619_47#_M1016_g 8.77977e-19 $X=4.22 $Y=1.56 $X2=0
+ $Y2=0
cc_380 N_A_805_21#_c_578_n N_A_619_47#_M1016_g 0.0167962f $X=5.005 $Y=1.93 $X2=0
+ $Y2=0
cc_381 N_A_805_21#_c_579_n N_A_619_47#_M1016_g 0.00435155f $X=5.1 $Y=2.425 $X2=0
+ $Y2=0
cc_382 N_A_805_21#_c_569_n N_A_619_47#_M1016_g 0.0121701f $X=4.22 $Y=1.9 $X2=0
+ $Y2=0
cc_383 N_A_805_21#_c_553_n N_A_619_47#_c_755_n 0.00225576f $X=4.115 $Y=0.765
+ $X2=0 $Y2=0
cc_384 N_A_805_21#_M1005_g N_A_619_47#_c_742_n 0.00145989f $X=4.13 $Y=2.665
+ $X2=0 $Y2=0
cc_385 N_A_805_21#_c_553_n N_A_619_47#_c_734_n 0.00481104f $X=4.115 $Y=0.765
+ $X2=0 $Y2=0
cc_386 N_A_805_21#_c_555_n N_A_619_47#_c_734_n 0.00327784f $X=4.22 $Y=1.395
+ $X2=0 $Y2=0
cc_387 N_A_805_21#_c_555_n N_A_619_47#_c_735_n 0.0137235f $X=4.22 $Y=1.395 $X2=0
+ $Y2=0
cc_388 N_A_805_21#_c_577_n N_A_619_47#_c_735_n 0.0215332f $X=4.232 $Y=1.795
+ $X2=0 $Y2=0
cc_389 N_A_805_21#_c_557_n N_A_619_47#_c_735_n 0.0289332f $X=4.22 $Y=1.56 $X2=0
+ $Y2=0
cc_390 N_A_805_21#_c_554_n N_A_619_47#_c_736_n 0.00128631f $X=4.115 $Y=0.915
+ $X2=0 $Y2=0
cc_391 N_A_805_21#_c_555_n N_A_619_47#_c_736_n 0.0198097f $X=4.22 $Y=1.395 $X2=0
+ $Y2=0
cc_392 N_A_805_21#_c_557_n N_A_619_47#_c_736_n 0.033891f $X=4.22 $Y=1.56 $X2=0
+ $Y2=0
cc_393 N_A_805_21#_c_558_n N_A_619_47#_c_736_n 0.00390517f $X=4.22 $Y=1.56 $X2=0
+ $Y2=0
cc_394 N_A_805_21#_c_578_n N_A_619_47#_c_736_n 0.0355086f $X=5.005 $Y=1.93 $X2=0
+ $Y2=0
cc_395 N_A_805_21#_c_560_n N_A_619_47#_c_736_n 0.0312645f $X=5.175 $Y=1.795
+ $X2=0 $Y2=0
cc_396 N_A_805_21#_c_570_n N_A_619_47#_c_736_n 0.003653f $X=5.055 $Y=1.125 $X2=0
+ $Y2=0
cc_397 N_A_805_21#_c_555_n N_A_619_47#_c_738_n 0.00263468f $X=4.22 $Y=1.395
+ $X2=0 $Y2=0
cc_398 N_A_805_21#_c_557_n N_A_619_47#_c_738_n 2.21651e-19 $X=4.22 $Y=1.56 $X2=0
+ $Y2=0
cc_399 N_A_805_21#_c_558_n N_A_619_47#_c_738_n 0.0142581f $X=4.22 $Y=1.56 $X2=0
+ $Y2=0
cc_400 N_A_805_21#_c_578_n N_A_619_47#_c_738_n 0.00141825f $X=5.005 $Y=1.93
+ $X2=0 $Y2=0
cc_401 N_A_805_21#_c_560_n N_A_619_47#_c_738_n 0.0139094f $X=5.175 $Y=1.795
+ $X2=0 $Y2=0
cc_402 N_A_805_21#_c_570_n N_A_619_47#_c_738_n 0.00193562f $X=5.055 $Y=1.125
+ $X2=0 $Y2=0
cc_403 N_A_805_21#_c_553_n N_A_619_47#_c_739_n 0.00801971f $X=4.115 $Y=0.765
+ $X2=0 $Y2=0
cc_404 N_A_805_21#_c_554_n N_A_619_47#_c_739_n 0.010567f $X=4.115 $Y=0.915 $X2=0
+ $Y2=0
cc_405 N_A_805_21#_c_560_n N_A_619_47#_c_739_n 0.00286135f $X=5.175 $Y=1.795
+ $X2=0 $Y2=0
cc_406 N_A_805_21#_c_562_n N_A_619_47#_c_739_n 0.00234955f $X=5.265 $Y=0.355
+ $X2=0 $Y2=0
cc_407 N_A_805_21#_c_565_n N_A_1138_153#_M1018_s 0.00288932f $X=6.04 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_408 N_A_805_21#_c_563_n N_A_1138_153#_c_827_n 7.78143e-19 $X=5.875 $Y=0.625
+ $X2=0 $Y2=0
cc_409 N_A_805_21#_c_564_n N_A_1138_153#_c_827_n 0.0164573f $X=7.275 $Y=0.71
+ $X2=0 $Y2=0
cc_410 N_A_805_21#_c_571_n N_A_1138_153#_c_827_n 0.0227081f $X=6.05 $Y=0.36
+ $X2=0 $Y2=0
cc_411 N_A_805_21#_M1018_g N_A_1138_153#_M1003_g 0.00890174f $X=6.05 $Y=0.975
+ $X2=0 $Y2=0
cc_412 N_A_805_21#_c_564_n N_A_1138_153#_c_829_n 3.51054e-19 $X=7.275 $Y=0.71
+ $X2=0 $Y2=0
cc_413 N_A_805_21#_c_550_n N_A_1138_153#_c_830_n 0.0222175f $X=7.735 $Y=1.295
+ $X2=0 $Y2=0
cc_414 N_A_805_21#_c_564_n N_A_1138_153#_c_830_n 0.0155624f $X=7.275 $Y=0.71
+ $X2=0 $Y2=0
cc_415 N_A_805_21#_c_566_n N_A_1138_153#_c_830_n 0.010599f $X=7.36 $Y=2.305
+ $X2=0 $Y2=0
cc_416 N_A_805_21#_M1004_g N_A_1138_153#_M1015_g 0.0237416f $X=7.655 $Y=2.465
+ $X2=0 $Y2=0
cc_417 N_A_805_21#_c_556_n N_A_1138_153#_c_832_n 0.0237416f $X=7.695 $Y=1.37
+ $X2=0 $Y2=0
cc_418 N_A_805_21#_M1018_g N_A_1138_153#_c_833_n 0.00855912f $X=6.05 $Y=0.975
+ $X2=0 $Y2=0
cc_419 N_A_805_21#_c_579_n N_A_1138_153#_c_833_n 0.0186768f $X=5.1 $Y=2.425
+ $X2=0 $Y2=0
cc_420 N_A_805_21#_c_560_n N_A_1138_153#_c_833_n 0.0183029f $X=5.175 $Y=1.795
+ $X2=0 $Y2=0
cc_421 N_A_805_21#_c_585_n N_A_1138_153#_c_833_n 0.0129766f $X=5.1 $Y=1.93 $X2=0
+ $Y2=0
cc_422 N_A_805_21#_M1018_g N_A_1138_153#_c_834_n 0.0169663f $X=6.05 $Y=0.975
+ $X2=0 $Y2=0
cc_423 N_A_805_21#_c_564_n N_A_1138_153#_c_834_n 0.0170912f $X=7.275 $Y=0.71
+ $X2=0 $Y2=0
cc_424 N_A_805_21#_c_565_n N_A_1138_153#_c_834_n 0.00128009f $X=6.04 $Y=0.71
+ $X2=0 $Y2=0
cc_425 N_A_805_21#_M1018_g N_A_1138_153#_c_835_n 0.0193619f $X=6.05 $Y=0.975
+ $X2=0 $Y2=0
cc_426 N_A_805_21#_c_561_n N_A_1138_153#_c_835_n 0.00149626f $X=5.71 $Y=0.355
+ $X2=0 $Y2=0
cc_427 N_A_805_21#_c_565_n N_A_1138_153#_c_835_n 0.0203883f $X=6.04 $Y=0.71
+ $X2=0 $Y2=0
cc_428 N_A_805_21#_c_570_n N_A_1138_153#_c_835_n 0.0183029f $X=5.055 $Y=1.125
+ $X2=0 $Y2=0
cc_429 N_A_805_21#_c_571_n N_A_1138_153#_c_835_n 0.00105015f $X=6.05 $Y=0.36
+ $X2=0 $Y2=0
cc_430 N_A_805_21#_M1018_g N_A_1138_153#_c_836_n 0.0213976f $X=6.05 $Y=0.975
+ $X2=0 $Y2=0
cc_431 N_A_805_21#_c_564_n N_A_1138_153#_c_836_n 0.00514989f $X=7.275 $Y=0.71
+ $X2=0 $Y2=0
cc_432 N_A_805_21#_c_578_n N_VPWR_M1005_d 0.00505212f $X=5.005 $Y=1.93 $X2=0
+ $Y2=0
cc_433 N_A_805_21#_c_566_n N_VPWR_M1015_d 0.00876168f $X=7.36 $Y=2.305 $X2=0
+ $Y2=0
cc_434 N_A_805_21#_c_582_n N_VPWR_M1015_d 0.00374628f $X=8.225 $Y=2.39 $X2=0
+ $Y2=0
cc_435 N_A_805_21#_c_652_p N_VPWR_M1015_d 0.00298231f $X=7.445 $Y=2.39 $X2=0
+ $Y2=0
cc_436 N_A_805_21#_c_582_n N_VPWR_M1021_s 0.00317287f $X=8.225 $Y=2.39 $X2=0
+ $Y2=0
cc_437 N_A_805_21#_c_567_n N_VPWR_M1021_s 0.00853892f $X=8.32 $Y=1.46 $X2=0
+ $Y2=0
cc_438 N_A_805_21#_M1005_g N_VPWR_c_894_n 0.00650631f $X=4.13 $Y=2.665 $X2=0
+ $Y2=0
cc_439 N_A_805_21#_c_577_n N_VPWR_c_894_n 0.00792636f $X=4.232 $Y=1.795 $X2=0
+ $Y2=0
cc_440 N_A_805_21#_c_578_n N_VPWR_c_894_n 0.0373898f $X=5.005 $Y=1.93 $X2=0
+ $Y2=0
cc_441 N_A_805_21#_c_579_n N_VPWR_c_894_n 0.0356104f $X=5.1 $Y=2.425 $X2=0 $Y2=0
cc_442 N_A_805_21#_c_586_n N_VPWR_c_894_n 0.00203907f $X=4.22 $Y=2.065 $X2=0
+ $Y2=0
cc_443 N_A_805_21#_M1018_g N_VPWR_c_895_n 0.00458918f $X=6.05 $Y=0.975 $X2=0
+ $Y2=0
cc_444 N_A_805_21#_M1004_g N_VPWR_c_896_n 0.0128734f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_445 N_A_805_21#_M1021_g N_VPWR_c_896_n 0.00172455f $X=8.085 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_A_805_21#_c_582_n N_VPWR_c_896_n 0.00718224f $X=8.225 $Y=2.39 $X2=0
+ $Y2=0
cc_447 N_A_805_21#_c_652_p N_VPWR_c_896_n 0.0147597f $X=7.445 $Y=2.39 $X2=0
+ $Y2=0
cc_448 N_A_805_21#_M1004_g N_VPWR_c_898_n 0.00176135f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A_805_21#_M1021_g N_VPWR_c_898_n 0.015633f $X=8.085 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_805_21#_c_582_n N_VPWR_c_898_n 0.0235013f $X=8.225 $Y=2.39 $X2=0
+ $Y2=0
cc_451 N_A_805_21#_M1005_g N_VPWR_c_900_n 0.00517164f $X=4.13 $Y=2.665 $X2=0
+ $Y2=0
cc_452 N_A_805_21#_M1018_g N_VPWR_c_901_n 0.00312414f $X=6.05 $Y=0.975 $X2=0
+ $Y2=0
cc_453 N_A_805_21#_c_579_n N_VPWR_c_901_n 0.0184952f $X=5.1 $Y=2.425 $X2=0 $Y2=0
cc_454 N_A_805_21#_M1004_g N_VPWR_c_903_n 0.00525069f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_455 N_A_805_21#_M1021_g N_VPWR_c_903_n 0.00486043f $X=8.085 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A_805_21#_M1005_g N_VPWR_c_891_n 0.00519032f $X=4.13 $Y=2.665 $X2=0
+ $Y2=0
cc_457 N_A_805_21#_M1018_g N_VPWR_c_891_n 0.00410284f $X=6.05 $Y=0.975 $X2=0
+ $Y2=0
cc_458 N_A_805_21#_M1004_g N_VPWR_c_891_n 0.0049745f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_459 N_A_805_21#_M1021_g N_VPWR_c_891_n 0.00465068f $X=8.085 $Y=2.465 $X2=0
+ $Y2=0
cc_460 N_A_805_21#_c_579_n N_VPWR_c_891_n 0.0100304f $X=5.1 $Y=2.425 $X2=0 $Y2=0
cc_461 N_A_805_21#_c_582_n N_VPWR_c_891_n 0.0191888f $X=8.225 $Y=2.39 $X2=0
+ $Y2=0
cc_462 N_A_805_21#_c_652_p N_VPWR_c_891_n 5.99846e-19 $X=7.445 $Y=2.39 $X2=0
+ $Y2=0
cc_463 N_A_805_21#_c_564_n N_Q_N_M1007_s 0.0045033f $X=7.275 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_464 N_A_805_21#_M1018_g N_Q_N_c_1002_n 0.00242382f $X=6.05 $Y=0.975 $X2=0
+ $Y2=0
cc_465 N_A_805_21#_M1004_g N_Q_N_c_1002_n 0.00115274f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_466 N_A_805_21#_c_564_n N_Q_N_c_1002_n 0.0170777f $X=7.275 $Y=0.71 $X2=0
+ $Y2=0
cc_467 N_A_805_21#_c_566_n N_Q_N_c_1002_n 0.0713712f $X=7.36 $Y=2.305 $X2=0
+ $Y2=0
cc_468 N_A_805_21#_c_582_n N_Q_M1004_d 0.00514444f $X=8.225 $Y=2.39 $X2=0 $Y2=0
cc_469 N_A_805_21#_c_550_n N_Q_c_1021_n 0.00581818f $X=7.735 $Y=1.295 $X2=0
+ $Y2=0
cc_470 N_A_805_21#_c_564_n N_Q_c_1021_n 0.00835692f $X=7.275 $Y=0.71 $X2=0 $Y2=0
cc_471 N_A_805_21#_c_566_n N_Q_c_1021_n 0.0723693f $X=7.36 $Y=2.305 $X2=0 $Y2=0
cc_472 N_A_805_21#_c_550_n Q 0.0058123f $X=7.735 $Y=1.295 $X2=0 $Y2=0
cc_473 N_A_805_21#_c_552_n Q 0.00386983f $X=8.165 $Y=1.295 $X2=0 $Y2=0
cc_474 N_A_805_21#_c_564_n Q 0.00144661f $X=7.275 $Y=0.71 $X2=0 $Y2=0
cc_475 N_A_805_21#_M1004_g Q 0.0135109f $X=7.655 $Y=2.465 $X2=0 $Y2=0
cc_476 N_A_805_21#_c_550_n Q 0.00969072f $X=7.735 $Y=1.295 $X2=0 $Y2=0
cc_477 N_A_805_21#_M1021_g Q 0.00888381f $X=8.085 $Y=2.465 $X2=0 $Y2=0
cc_478 N_A_805_21#_c_556_n Q 0.00299603f $X=7.695 $Y=1.37 $X2=0 $Y2=0
cc_479 N_A_805_21#_c_582_n Q 0.0178394f $X=8.225 $Y=2.39 $X2=0 $Y2=0
cc_480 N_A_805_21#_c_567_n Q 0.0609212f $X=8.32 $Y=1.46 $X2=0 $Y2=0
cc_481 N_A_805_21#_c_568_n Q 0.00800124f $X=8.32 $Y=1.46 $X2=0 $Y2=0
cc_482 N_A_805_21#_c_572_n Q 0.00766458f $X=8.01 $Y=1.46 $X2=0 $Y2=0
cc_483 N_A_805_21#_c_564_n N_VGND_M1018_d 0.0117022f $X=7.275 $Y=0.71 $X2=0
+ $Y2=0
cc_484 N_A_805_21#_c_564_n N_VGND_M1024_d 0.00402952f $X=7.275 $Y=0.71 $X2=0
+ $Y2=0
cc_485 N_A_805_21#_c_566_n N_VGND_M1024_d 0.00630766f $X=7.36 $Y=2.305 $X2=0
+ $Y2=0
cc_486 N_A_805_21#_c_553_n N_VGND_c_1046_n 0.0104384f $X=4.115 $Y=0.765 $X2=0
+ $Y2=0
cc_487 N_A_805_21#_c_554_n N_VGND_c_1046_n 0.00146965f $X=4.115 $Y=0.915 $X2=0
+ $Y2=0
cc_488 N_A_805_21#_c_562_n N_VGND_c_1046_n 0.00936016f $X=5.265 $Y=0.355 $X2=0
+ $Y2=0
cc_489 N_A_805_21#_c_706_p N_VGND_c_1047_n 0.0160692f $X=5.875 $Y=0.455 $X2=0
+ $Y2=0
cc_490 N_A_805_21#_c_564_n N_VGND_c_1047_n 0.02498f $X=7.275 $Y=0.71 $X2=0 $Y2=0
cc_491 N_A_805_21#_c_571_n N_VGND_c_1047_n 0.00394083f $X=6.05 $Y=0.36 $X2=0
+ $Y2=0
cc_492 N_A_805_21#_c_550_n N_VGND_c_1048_n 0.00254608f $X=7.735 $Y=1.295 $X2=0
+ $Y2=0
cc_493 N_A_805_21#_c_564_n N_VGND_c_1048_n 0.0140995f $X=7.275 $Y=0.71 $X2=0
+ $Y2=0
cc_494 N_A_805_21#_c_550_n N_VGND_c_1050_n 6.75831e-19 $X=7.735 $Y=1.295 $X2=0
+ $Y2=0
cc_495 N_A_805_21#_c_552_n N_VGND_c_1050_n 0.0170688f $X=8.165 $Y=1.295 $X2=0
+ $Y2=0
cc_496 N_A_805_21#_c_567_n N_VGND_c_1050_n 0.0203551f $X=8.32 $Y=1.46 $X2=0
+ $Y2=0
cc_497 N_A_805_21#_c_568_n N_VGND_c_1050_n 0.00176637f $X=8.32 $Y=1.46 $X2=0
+ $Y2=0
cc_498 N_A_805_21#_c_561_n N_VGND_c_1053_n 0.0289308f $X=5.71 $Y=0.355 $X2=0
+ $Y2=0
cc_499 N_A_805_21#_c_562_n N_VGND_c_1053_n 0.0301084f $X=5.265 $Y=0.355 $X2=0
+ $Y2=0
cc_500 N_A_805_21#_c_706_p N_VGND_c_1053_n 0.022125f $X=5.875 $Y=0.455 $X2=0
+ $Y2=0
cc_501 N_A_805_21#_c_564_n N_VGND_c_1053_n 0.00317388f $X=7.275 $Y=0.71 $X2=0
+ $Y2=0
cc_502 N_A_805_21#_c_571_n N_VGND_c_1053_n 0.008223f $X=6.05 $Y=0.36 $X2=0 $Y2=0
cc_503 N_A_805_21#_c_553_n N_VGND_c_1055_n 0.00585385f $X=4.115 $Y=0.765 $X2=0
+ $Y2=0
cc_504 N_A_805_21#_c_554_n N_VGND_c_1055_n 5.95547e-19 $X=4.115 $Y=0.915 $X2=0
+ $Y2=0
cc_505 N_A_805_21#_c_564_n N_VGND_c_1056_n 0.010819f $X=7.275 $Y=0.71 $X2=0
+ $Y2=0
cc_506 N_A_805_21#_c_550_n N_VGND_c_1057_n 0.00378237f $X=7.735 $Y=1.295 $X2=0
+ $Y2=0
cc_507 N_A_805_21#_c_552_n N_VGND_c_1057_n 0.00400407f $X=8.165 $Y=1.295 $X2=0
+ $Y2=0
cc_508 N_A_805_21#_c_550_n N_VGND_c_1061_n 0.00601326f $X=7.735 $Y=1.295 $X2=0
+ $Y2=0
cc_509 N_A_805_21#_c_552_n N_VGND_c_1061_n 0.00774504f $X=8.165 $Y=1.295 $X2=0
+ $Y2=0
cc_510 N_A_805_21#_c_553_n N_VGND_c_1061_n 0.0123431f $X=4.115 $Y=0.765 $X2=0
+ $Y2=0
cc_511 N_A_805_21#_c_554_n N_VGND_c_1061_n 8.01698e-19 $X=4.115 $Y=0.915 $X2=0
+ $Y2=0
cc_512 N_A_805_21#_c_561_n N_VGND_c_1061_n 0.016781f $X=5.71 $Y=0.355 $X2=0
+ $Y2=0
cc_513 N_A_805_21#_c_562_n N_VGND_c_1061_n 0.0163286f $X=5.265 $Y=0.355 $X2=0
+ $Y2=0
cc_514 N_A_805_21#_c_706_p N_VGND_c_1061_n 0.011244f $X=5.875 $Y=0.455 $X2=0
+ $Y2=0
cc_515 N_A_805_21#_c_564_n N_VGND_c_1061_n 0.0265757f $X=7.275 $Y=0.71 $X2=0
+ $Y2=0
cc_516 N_A_805_21#_c_571_n N_VGND_c_1061_n 0.0117988f $X=6.05 $Y=0.36 $X2=0
+ $Y2=0
cc_517 N_A_619_47#_c_741_n N_VPWR_c_893_n 0.00679097f $X=3.445 $Y=2.6 $X2=0
+ $Y2=0
cc_518 N_A_619_47#_M1016_g N_VPWR_c_894_n 0.0190971f $X=4.885 $Y=2.415 $X2=0
+ $Y2=0
cc_519 N_A_619_47#_c_741_n N_VPWR_c_894_n 0.0114891f $X=3.445 $Y=2.6 $X2=0 $Y2=0
cc_520 N_A_619_47#_c_742_n N_VPWR_c_894_n 0.00735747f $X=3.79 $Y=2.475 $X2=0
+ $Y2=0
cc_521 N_A_619_47#_c_735_n N_VPWR_c_894_n 0.00895169f $X=3.875 $Y=2.39 $X2=0
+ $Y2=0
cc_522 N_A_619_47#_c_741_n N_VPWR_c_900_n 0.0210569f $X=3.445 $Y=2.6 $X2=0 $Y2=0
cc_523 N_A_619_47#_M1016_g N_VPWR_c_901_n 0.00445056f $X=4.885 $Y=2.415 $X2=0
+ $Y2=0
cc_524 N_A_619_47#_M1020_d N_VPWR_c_891_n 0.00215158f $X=3.305 $Y=2.455 $X2=0
+ $Y2=0
cc_525 N_A_619_47#_M1016_g N_VPWR_c_891_n 0.00899805f $X=4.885 $Y=2.415 $X2=0
+ $Y2=0
cc_526 N_A_619_47#_c_741_n N_VPWR_c_891_n 0.0125713f $X=3.445 $Y=2.6 $X2=0 $Y2=0
cc_527 N_A_619_47#_c_742_n N_VPWR_c_891_n 0.0131576f $X=3.79 $Y=2.475 $X2=0
+ $Y2=0
cc_528 N_A_619_47#_c_742_n A_769_491# 0.00239886f $X=3.79 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_529 N_A_619_47#_c_736_n N_VGND_M1017_d 0.00572264f $X=4.505 $Y=1.14 $X2=0
+ $Y2=0
cc_530 N_A_619_47#_c_755_n N_VGND_c_1046_n 0.0110535f $X=3.79 $Y=0.355 $X2=0
+ $Y2=0
cc_531 N_A_619_47#_c_734_n N_VGND_c_1046_n 0.0220426f $X=3.875 $Y=1.055 $X2=0
+ $Y2=0
cc_532 N_A_619_47#_c_736_n N_VGND_c_1046_n 0.0273879f $X=4.505 $Y=1.14 $X2=0
+ $Y2=0
cc_533 N_A_619_47#_c_739_n N_VGND_c_1046_n 0.00770369f $X=4.777 $Y=1.295 $X2=0
+ $Y2=0
cc_534 N_A_619_47#_c_739_n N_VGND_c_1053_n 0.00482246f $X=4.777 $Y=1.295 $X2=0
+ $Y2=0
cc_535 N_A_619_47#_c_755_n N_VGND_c_1055_n 0.0493072f $X=3.79 $Y=0.355 $X2=0
+ $Y2=0
cc_536 N_A_619_47#_M1022_d N_VGND_c_1061_n 0.00378179f $X=3.095 $Y=0.235 $X2=0
+ $Y2=0
cc_537 N_A_619_47#_c_755_n N_VGND_c_1061_n 0.0300599f $X=3.79 $Y=0.355 $X2=0
+ $Y2=0
cc_538 N_A_619_47#_c_739_n N_VGND_c_1061_n 0.00994426f $X=4.777 $Y=1.295 $X2=0
+ $Y2=0
cc_539 N_A_619_47#_c_755_n A_737_47# 0.00714088f $X=3.79 $Y=0.355 $X2=-0.19
+ $Y2=-0.245
cc_540 N_A_619_47#_c_734_n A_737_47# 0.00529158f $X=3.875 $Y=1.055 $X2=-0.19
+ $Y2=-0.245
cc_541 N_A_1138_153#_M1003_g N_VPWR_c_895_n 0.00931197f $X=6.715 $Y=2.465 $X2=0
+ $Y2=0
cc_542 N_A_1138_153#_c_833_n N_VPWR_c_895_n 0.00405624f $X=5.835 $Y=1.98 $X2=0
+ $Y2=0
cc_543 N_A_1138_153#_c_834_n N_VPWR_c_895_n 0.0386028f $X=6.5 $Y=1.46 $X2=0
+ $Y2=0
cc_544 N_A_1138_153#_c_836_n N_VPWR_c_895_n 0.00580062f $X=6.79 $Y=1.46 $X2=0
+ $Y2=0
cc_545 N_A_1138_153#_M1015_g N_VPWR_c_896_n 0.00547999f $X=7.145 $Y=2.465 $X2=0
+ $Y2=0
cc_546 N_A_1138_153#_M1003_g N_VPWR_c_902_n 0.0054895f $X=6.715 $Y=2.465 $X2=0
+ $Y2=0
cc_547 N_A_1138_153#_M1015_g N_VPWR_c_902_n 0.0054895f $X=7.145 $Y=2.465 $X2=0
+ $Y2=0
cc_548 N_A_1138_153#_M1003_g N_VPWR_c_891_n 0.0110927f $X=6.715 $Y=2.465 $X2=0
+ $Y2=0
cc_549 N_A_1138_153#_M1015_g N_VPWR_c_891_n 0.0100951f $X=7.145 $Y=2.465 $X2=0
+ $Y2=0
cc_550 N_A_1138_153#_c_833_n N_VPWR_c_891_n 0.0115026f $X=5.835 $Y=1.98 $X2=0
+ $Y2=0
cc_551 N_A_1138_153#_c_827_n N_Q_N_c_1002_n 0.00880335f $X=6.715 $Y=1.295 $X2=0
+ $Y2=0
cc_552 N_A_1138_153#_M1003_g N_Q_N_c_1002_n 0.0215912f $X=6.715 $Y=2.465 $X2=0
+ $Y2=0
cc_553 N_A_1138_153#_c_829_n N_Q_N_c_1002_n 0.00839308f $X=7.07 $Y=1.37 $X2=0
+ $Y2=0
cc_554 N_A_1138_153#_c_830_n N_Q_N_c_1002_n 0.00511386f $X=7.145 $Y=1.295 $X2=0
+ $Y2=0
cc_555 N_A_1138_153#_M1015_g N_Q_N_c_1002_n 0.024771f $X=7.145 $Y=2.465 $X2=0
+ $Y2=0
cc_556 N_A_1138_153#_c_832_n N_Q_N_c_1002_n 0.00158441f $X=7.145 $Y=1.37 $X2=0
+ $Y2=0
cc_557 N_A_1138_153#_c_834_n N_Q_N_c_1002_n 0.0247039f $X=6.5 $Y=1.46 $X2=0
+ $Y2=0
cc_558 N_A_1138_153#_c_836_n N_Q_N_c_1002_n 0.00750545f $X=6.79 $Y=1.46 $X2=0
+ $Y2=0
cc_559 N_A_1138_153#_c_830_n N_Q_c_1021_n 5.83282e-19 $X=7.145 $Y=1.295 $X2=0
+ $Y2=0
cc_560 N_A_1138_153#_c_830_n Q 8.33023e-19 $X=7.145 $Y=1.295 $X2=0 $Y2=0
cc_561 N_A_1138_153#_c_827_n N_VGND_c_1047_n 0.00668067f $X=6.715 $Y=1.295 $X2=0
+ $Y2=0
cc_562 N_A_1138_153#_c_830_n N_VGND_c_1048_n 0.00426942f $X=7.145 $Y=1.295 $X2=0
+ $Y2=0
cc_563 N_A_1138_153#_c_827_n N_VGND_c_1056_n 0.00341315f $X=6.715 $Y=1.295 $X2=0
+ $Y2=0
cc_564 N_A_1138_153#_c_830_n N_VGND_c_1056_n 0.00341315f $X=7.145 $Y=1.295 $X2=0
+ $Y2=0
cc_565 N_A_1138_153#_c_827_n N_VGND_c_1061_n 0.00466594f $X=6.715 $Y=1.295 $X2=0
+ $Y2=0
cc_566 N_A_1138_153#_c_830_n N_VGND_c_1061_n 0.00458952f $X=7.145 $Y=1.295 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_891_n A_589_491# 0.00422333f $X=8.4 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_568 N_VPWR_c_891_n N_Q_N_M1003_s 0.00223559f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_569 N_VPWR_c_895_n N_Q_N_c_1002_n 0.0475101f $X=6.265 $Y=1.96 $X2=0 $Y2=0
cc_570 N_VPWR_c_902_n N_Q_N_c_1002_n 0.0189236f $X=7.265 $Y=3.33 $X2=0 $Y2=0
cc_571 N_VPWR_c_891_n N_Q_N_c_1002_n 0.0123859f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_572 N_VPWR_c_891_n N_Q_M1004_d 0.00417163f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_573 Q N_VGND_c_1048_n 0.00513078f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_574 Q N_VGND_c_1050_n 0.0303953f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_575 N_Q_c_1021_n N_VGND_c_1057_n 0.00118198f $X=7.875 $Y=0.825 $X2=0 $Y2=0
cc_576 Q N_VGND_c_1057_n 0.0128944f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_577 N_Q_c_1021_n N_VGND_c_1061_n 0.00170782f $X=7.875 $Y=0.825 $X2=0 $Y2=0
cc_578 Q N_VGND_c_1061_n 0.00985309f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_579 N_VGND_c_1061_n A_547_47# 0.00241193f $X=8.4 $Y=0 $X2=-0.19 $Y2=-0.245
cc_580 N_VGND_c_1061_n A_737_47# 0.00499543f $X=8.4 $Y=0 $X2=-0.19 $Y2=-0.245
