* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_58_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.1214e+12p ps=9.34e+06u
M1001 a_326_69# A1 Y VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=3.36e+11p ps=2.48e+06u
M1002 a_58_367# B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A3 a_58_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1151e+12p pd=6.81e+06u as=0p ps=0u
M1004 Y B1 a_141_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.89e+11p ps=2.13e+06u
M1005 VPWR A1 a_58_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_141_69# B2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.452e+11p ps=4.42e+06u
M1007 a_58_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_434_69# A2 a_326_69# VNB nshort w=840000u l=150000u
+  ad=3.696e+11p pd=2.56e+06u as=0p ps=0u
M1009 VGND A3 a_434_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
