* File: sky130_fd_sc_lp__a2111oi_4.spice
* Created: Fri Aug 28 09:46:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111oi_4.pex.spice"
.subckt sky130_fd_sc_lp__a2111oi_4  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1014 N_Y_M1014_d N_D1_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75005
+ A=0.126 P=1.98 MULT=1
MM1022 N_Y_M1014_d N_D1_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.6 A=0.126 P=1.98 MULT=1
MM1023 N_Y_M1023_d N_D1_M1023_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.2 A=0.126 P=1.98 MULT=1
MM1039 N_Y_M1023_d N_D1_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1039_s N_C1_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_C1_M1018_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1018_d N_C1_M1031_g N_Y_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1034 N_VGND_M1034_d N_C1_M1034_g N_Y_M1031_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1176 PD=1.23 PS=1.12 NRD=8.568 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VGND_M1034_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=7.14 M=1 R=5.6 SA=75003.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1001_d N_B1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1019 N_Y_M1019_d N_B1_M1019_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1025 N_Y_M1019_d N_B1_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75005 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1002_d N_A1_M1002_g N_A_1201_47#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1013 N_Y_M1002_d N_A1_M1013_g N_A_1201_47#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1015 N_Y_M1015_d N_A1_M1015_g N_A_1201_47#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1029 N_Y_M1015_d N_A1_M1029_g N_A_1201_47#_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1575 PD=1.12 PS=1.215 NRD=0 NRS=12.852 M=1 R=5.6 SA=75001.5
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1004 N_A_1201_47#_M1029_s N_A2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1575 AS=0.1176 PD=1.215 PS=1.12 NRD=0.708 NRS=0 M=1 R=5.6 SA=75002
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_A_1201_47#_M1005_d N_A2_M1005_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1021 N_A_1201_47#_M1005_d N_A2_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1026 N_A_1201_47#_M1026_d N_A2_M1026_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_D1_M1000_g N_A_27_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1000_d N_D1_M1016_g N_A_27_367#_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1027 N_Y_M1027_d N_D1_M1027_g N_A_27_367#_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1038 N_Y_M1027_d N_D1_M1038_g N_A_27_367#_M1038_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 N_A_454_367#_M1006_d N_C1_M1006_g N_A_27_367#_M1038_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_A_454_367#_M1006_d N_C1_M1010_g N_A_27_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1030 N_A_454_367#_M1030_d N_C1_M1030_g N_A_27_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1032 N_A_454_367#_M1030_d N_C1_M1032_g N_A_27_367#_M1032_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_A_454_367#_M1007_d N_B1_M1007_g N_A_819_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1011 N_A_454_367#_M1007_d N_B1_M1011_g N_A_819_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1033 N_A_454_367#_M1033_d N_B1_M1033_g N_A_819_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1035 N_A_454_367#_M1033_d N_B1_M1035_g N_A_819_367#_M1035_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1008 N_A_819_367#_M1035_s N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1020 N_A_819_367#_M1020_d N_A1_M1020_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1024 N_A_819_367#_M1020_d N_A1_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.189 PD=1.54 PS=1.56 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1028 N_A_819_367#_M1028_d N_A1_M1028_g N_VPWR_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.252 AS=0.189 PD=1.66 PS=1.56 NRD=5.2008 NRS=3.1126 M=1 R=8.4
+ SA=75003.2 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A2_M1012_g N_A_819_367#_M1028_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.252 PD=1.54 PS=1.66 NRD=0 NRS=13.5339 M=1 R=8.4
+ SA=75003.8 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1012_d N_A2_M1017_g N_A_819_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2331 PD=1.54 PS=1.63 NRD=0 NRS=9.3772 M=1 R=8.4
+ SA=75004.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1036 N_VPWR_M1036_d N_A2_M1036_g N_A_819_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2331 PD=1.54 PS=1.63 NRD=0 NRS=4.6886 M=1 R=8.4
+ SA=75004.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1036_d N_A2_M1037_g N_A_819_367#_M1037_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.5079 P=24.65
c_92 VNB 0 1.34154e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a2111oi_4.pxi.spice"
*
.ends
*
*
