* File: sky130_fd_sc_lp__fah_1.spice
* Created: Wed Sep  2 09:53:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fah_1.pex.spice"
.subckt sky130_fd_sc_lp__fah_1  VNB VPB CI B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* CI	CI
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_84_21#_M1006_g N_SUM_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.241812 AS=0.2394 PD=1.6573 PS=2.25 NRD=17.136 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_A_239_135#_M1008_d N_CI_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.184238 PD=1.85 PS=1.2627 NRD=0 NRS=43.656 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A_413_34#_M1004_g N_COUT_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.317497 AS=0.2394 PD=1.84459 PS=2.25 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1027 N_A_630_100#_M1027_d N_A_239_135#_M1027_g N_VGND_M1004_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.29515 AS=0.241903 PD=2.35 PS=1.40541 NRD=22.488 NRS=95.616
+ M=1 R=4.26667 SA=75001.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1024 N_A_413_34#_M1024_d N_A_814_384#_M1024_g N_A_878_41#_M1024_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.37535 PD=0.92 PS=2.93 NRD=0 NRS=99.648 M=1
+ R=4.26667 SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 N_A_239_135#_M1002_d N_A_1022_362#_M1002_g N_A_413_34#_M1024_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1023 N_A_84_21#_M1023_d N_A_814_384#_M1023_g N_A_239_135#_M1002_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.13795 AS=0.0896 PD=1.2 PS=0.92 NRD=22.5 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_630_100#_M1017_d N_A_1022_362#_M1017_g N_A_84_21#_M1023_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.13795 PD=1.85 PS=1.2 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1028 N_VGND_M1028_d N_B_M1028_g N_A_878_41#_M1028_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.2394 PD=2.25 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_1022_362#_M1005_d N_A_878_41#_M1005_g N_A_1741_367#_M1005_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1025 N_A_1930_367#_M1025_d N_B_M1025_g N_A_1022_362#_M1005_d VNB NSHORT L=0.15
+ W=0.64 AD=0.16755 AS=0.0896 PD=1.18 PS=0.92 NRD=21.552 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75002 A=0.096 P=1.58 MULT=1
MM1014 N_A_814_384#_M1014_d N_A_878_41#_M1014_g N_A_1930_367#_M1025_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.16755 PD=0.92 PS=1.18 NRD=0 NRS=21.552 M=1
+ R=4.26667 SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1009 N_A_1741_367#_M1009_d N_B_M1009_g N_A_814_384#_M1014_d VNB NSHORT L=0.15
+ W=0.64 AD=0.133968 AS=0.0896 PD=1.06811 PS=0.92 NRD=21.552 NRS=0 M=1 R=4.26667
+ SA=75001.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1019 N_VGND_M1019_d N_A_2229_269#_M1019_g N_A_1741_367#_M1009_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.481775 AS=0.175832 PD=2.86 PS=1.40189 NRD=38.568 NRS=0 M=1
+ R=5.6 SA=75001.7 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1026 N_VGND_M1026_d N_A_M1026_g N_A_1930_367#_M1026_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_2229_269#_M1010_d N_A_M1010_g N_VGND_M1026_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1018_d N_A_84_21#_M1018_g N_SUM_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.342876 AS=0.3591 PD=2.01823 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1011 N_A_239_135#_M1011_d N_CI_M1011_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.272124 PD=2.57 PS=1.60177 NRD=0 NRS=53.1703 M=1 R=6.66667
+ SA=75000.9 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_413_34#_M1007_g N_COUT_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.414741 AS=0.3591 PD=2.20779 PS=3.09 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.6 A=0.189 P=2.82 MULT=1
MM1012 N_A_630_100#_M1012_d N_A_239_135#_M1012_g N_VPWR_M1007_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.293614 AS=0.329159 PD=1.82065 PS=1.75221 NRD=22.6353
+ NRS=53.9977 M=1 R=6.66667 SA=75001 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1013 N_A_84_21#_M1013_d N_A_814_384#_M1013_g N_A_630_100#_M1012_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.35235 AS=0.246636 PD=1.84 PS=1.52935 NRD=0 NRS=55.948 M=1
+ R=5.6 SA=75001.4 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1001 N_A_239_135#_M1001_d N_A_1022_362#_M1001_g N_A_84_21#_M1013_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.239575 AS=0.35235 PD=1.525 PS=1.84 NRD=26.9693 NRS=143.042
+ M=1 R=5.6 SA=75002.3 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1020 N_A_413_34#_M1020_d N_A_814_384#_M1020_g N_A_239_135#_M1001_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2163 AS=0.239575 PD=1.355 PS=1.525 NRD=0 NRS=53.978 M=1
+ R=5.6 SA=75002.4 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1015 N_A_878_41#_M1015_d N_A_1022_362#_M1015_g N_A_413_34#_M1020_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1806 AS=0.2163 PD=1.324 PS=1.355 NRD=26.9693 NRS=55.1009
+ M=1 R=5.6 SA=75003 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1022 N_VPWR_M1022_d N_B_M1022_g N_A_878_41#_M1015_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.2709 PD=3.09 PS=1.986 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_A_814_384#_M1003_d N_A_878_41#_M1003_g N_A_1741_367#_M1003_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1176 AS=0.3066 PD=1.12 PS=2.41 NRD=0 NRS=18.7544
+ M=1 R=5.6 SA=75000.3 SB=75002.6 A=0.126 P=1.98 MULT=1
MM1021 N_A_1930_367#_M1021_d N_B_M1021_g N_A_814_384#_M1003_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.233575 AS=0.1176 PD=1.55 PS=1.12 NRD=52.3035 NRS=0 M=1 R=5.6
+ SA=75000.7 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1029 N_A_1022_362#_M1029_d N_A_878_41#_M1029_g N_A_1930_367#_M1021_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1512 AS=0.233575 PD=1.2 PS=1.55 NRD=0 NRS=52.3035
+ M=1 R=5.6 SA=75001.3 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1031 N_A_1741_367#_M1031_d N_B_M1031_g N_A_1022_362#_M1029_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.16296 AS=0.1512 PD=1.296 PS=1.2 NRD=0 NRS=18.7544 M=1 R=5.6
+ SA=75001.9 SB=75001 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_2229_269#_M1000_g N_A_1741_367#_M1031_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.732675 AS=0.24444 PD=3.78 PS=1.944 NRD=42.9854 NRS=12.4898
+ M=1 R=8.4 SA=75001.6 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_1930_367#_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1016 N_A_2229_269#_M1016_d N_A_M1016_g N_VPWR_M1030_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=25.7743 P=31.37
c_141 VNB 0 1.67676e-19 $X=0 $Y=0
c_264 VPB 0 2.56143e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__fah_1.pxi.spice"
*
.ends
*
*
