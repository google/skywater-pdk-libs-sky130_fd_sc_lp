* File: sky130_fd_sc_lp__o21a_lp.pxi.spice
* Created: Wed Sep  2 10:15:35 2020
* 
x_PM_SKY130_FD_SC_LP__O21A_LP%A1 N_A1_c_61_n N_A1_M1004_g N_A1_c_66_n
+ N_A1_M1000_g A1 A1 N_A1_c_64_n PM_SKY130_FD_SC_LP__O21A_LP%A1
x_PM_SKY130_FD_SC_LP__O21A_LP%A2 N_A2_M1003_g N_A2_c_99_n N_A2_M1002_g
+ N_A2_c_96_n A2 A2 A2 A2 A2 N_A2_c_98_n PM_SKY130_FD_SC_LP__O21A_LP%A2
x_PM_SKY130_FD_SC_LP__O21A_LP%B1 N_B1_M1005_g N_B1_M1001_g B1 N_B1_c_147_n
+ PM_SKY130_FD_SC_LP__O21A_LP%B1
x_PM_SKY130_FD_SC_LP__O21A_LP%A_244_409# N_A_244_409#_M1005_d
+ N_A_244_409#_M1002_d N_A_244_409#_M1006_g N_A_244_409#_M1007_g
+ N_A_244_409#_M1008_g N_A_244_409#_c_185_n N_A_244_409#_c_186_n
+ N_A_244_409#_c_194_n N_A_244_409#_c_187_n N_A_244_409#_c_195_n
+ N_A_244_409#_c_196_n N_A_244_409#_c_188_n N_A_244_409#_c_189_n
+ N_A_244_409#_c_190_n N_A_244_409#_c_191_n N_A_244_409#_c_192_n
+ PM_SKY130_FD_SC_LP__O21A_LP%A_244_409#
x_PM_SKY130_FD_SC_LP__O21A_LP%VPWR N_VPWR_M1000_s N_VPWR_M1001_d N_VPWR_c_256_n
+ N_VPWR_c_257_n N_VPWR_c_258_n VPWR N_VPWR_c_259_n N_VPWR_c_260_n
+ N_VPWR_c_255_n N_VPWR_c_262_n PM_SKY130_FD_SC_LP__O21A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O21A_LP%X N_X_M1008_d N_X_M1006_d N_X_c_291_n N_X_c_292_n
+ X X X X N_X_c_290_n PM_SKY130_FD_SC_LP__O21A_LP%X
x_PM_SKY130_FD_SC_LP__O21A_LP%A_27_57# N_A_27_57#_M1004_s N_A_27_57#_M1003_d
+ N_A_27_57#_c_314_n N_A_27_57#_c_315_n N_A_27_57#_c_316_n N_A_27_57#_c_317_n
+ PM_SKY130_FD_SC_LP__O21A_LP%A_27_57#
x_PM_SKY130_FD_SC_LP__O21A_LP%VGND N_VGND_M1004_d N_VGND_M1007_s N_VGND_c_343_n
+ N_VGND_c_344_n VGND N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n
+ N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n PM_SKY130_FD_SC_LP__O21A_LP%VGND
cc_1 VNB N_A1_c_61_n 0.0251214f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.64
cc_2 VNB N_A1_M1004_g 0.0475617f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_3 VNB A1 0.0212606f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_64_n 0.0257603f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.34
cc_5 VNB N_A2_M1003_g 0.0373652f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.175
cc_6 VNB N_A2_c_96_n 0.00793161f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB A2 0.00808691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_98_n 0.0301908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_M1005_g 0.0443373f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.175
cc_10 VNB N_B1_M1001_g 0.0104437f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.97
cc_11 VNB B1 0.00508234f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.545
cc_12 VNB N_B1_c_147_n 0.0562627f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.34
cc_13 VNB N_A_244_409#_M1006_g 0.011453f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.545
cc_14 VNB N_A_244_409#_M1007_g 0.0220446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_244_409#_M1008_g 0.0228408f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.175
cc_16 VNB N_A_244_409#_c_185_n 0.0353439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_244_409#_c_186_n 0.0175393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_244_409#_c_187_n 0.00950696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_244_409#_c_188_n 0.00633173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_244_409#_c_189_n 0.00665366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_244_409#_c_190_n 0.0112087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_244_409#_c_191_n 0.0028678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_244_409#_c_192_n 0.0291425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_255_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_290_n 0.0649419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_57#_c_314_n 0.0240181f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.545
cc_27 VNB N_A_27_57#_c_315_n 0.0198721f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_A_27_57#_c_316_n 0.010309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_57#_c_317_n 0.00370575f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.34
cc_30 VNB N_VGND_c_343_n 0.00651576f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.545
cc_31 VNB N_VGND_c_344_n 0.00682676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_345_n 0.019006f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.175
cc_33 VNB N_VGND_c_346_n 0.0336618f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_34 VNB N_VGND_c_347_n 0.0270417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_348_n 0.20311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_349_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_350_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A1_c_61_n 0.0424902f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.64
cc_39 VPB N_A1_c_66_n 0.0237725f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.97
cc_40 VPB A1 0.012241f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_41 VPB N_A2_c_99_n 0.00937461f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.97
cc_42 VPB N_A2_M1002_g 0.0273479f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.545
cc_43 VPB N_A2_c_96_n 0.00490217f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_44 VPB A2 0.00663286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B1_M1001_g 0.0420358f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.97
cc_46 VPB N_A_244_409#_M1006_g 0.0461481f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.545
cc_47 VPB N_A_244_409#_c_194_n 0.00467056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_244_409#_c_195_n 0.00309935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_244_409#_c_196_n 0.00383443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_244_409#_c_188_n 2.7562e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_256_n 0.0132707f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.97
cc_52 VPB N_VPWR_c_257_n 0.0461962f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.545
cc_53 VPB N_VPWR_c_258_n 0.00927422f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.34
cc_54 VPB N_VPWR_c_259_n 0.0409445f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.34
cc_55 VPB N_VPWR_c_260_n 0.0303808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_255_n 0.0820293f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_262_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_X_c_291_n 0.0323816f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.545
cc_59 VPB N_X_c_292_n 0.0243257f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.34
cc_60 VPB N_X_c_290_n 0.0284283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 N_A1_M1004_g N_A2_M1003_g 0.0268164f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_62 N_A1_c_64_n N_A2_M1003_g 2.11782e-19 $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_63 N_A1_c_61_n N_A2_c_99_n 0.0352525f $X=0.425 $Y=1.64 $X2=0 $Y2=0
cc_64 N_A1_c_66_n N_A2_M1002_g 0.0352525f $X=0.605 $Y=1.97 $X2=0 $Y2=0
cc_65 N_A1_c_61_n N_A2_c_96_n 0.0113231f $X=0.425 $Y=1.64 $X2=0 $Y2=0
cc_66 A1 N_A2_c_96_n 3.33801e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A1_c_61_n A2 0.0154892f $X=0.425 $Y=1.64 $X2=0 $Y2=0
cc_68 A1 A2 0.0327997f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A1_c_64_n A2 0.00132278f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_70 A1 N_A2_c_98_n 0.00107341f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A1_c_64_n N_A2_c_98_n 0.0176376f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_72 N_A1_c_61_n N_VPWR_c_257_n 0.00202045f $X=0.425 $Y=1.64 $X2=0 $Y2=0
cc_73 N_A1_c_66_n N_VPWR_c_257_n 0.0241304f $X=0.605 $Y=1.97 $X2=0 $Y2=0
cc_74 A1 N_VPWR_c_257_n 0.0280615f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A1_c_66_n N_VPWR_c_259_n 0.00802402f $X=0.605 $Y=1.97 $X2=0 $Y2=0
cc_76 N_A1_c_66_n N_VPWR_c_255_n 0.0142664f $X=0.605 $Y=1.97 $X2=0 $Y2=0
cc_77 N_A1_M1004_g N_A_27_57#_c_314_n 0.0110202f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_78 N_A1_M1004_g N_A_27_57#_c_315_n 0.00958284f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_79 A1 N_A_27_57#_c_315_n 0.00752329f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A1_c_64_n N_A_27_57#_c_315_n 0.00246363f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_81 N_A1_M1004_g N_A_27_57#_c_316_n 0.004207f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_82 A1 N_A_27_57#_c_316_n 0.0275186f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A1_c_64_n N_A_27_57#_c_316_n 0.00155458f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_84 N_A1_M1004_g N_A_27_57#_c_317_n 6.34679e-19 $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_85 N_A1_M1004_g N_VGND_c_343_n 0.00268233f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_86 N_A1_M1004_g N_VGND_c_345_n 0.00502664f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_87 N_A1_M1004_g N_VGND_c_348_n 0.00643613f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_88 N_A2_M1003_g N_B1_M1005_g 0.0258632f $X=1.005 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A2_c_99_n N_B1_M1001_g 0.0142969f $X=1.095 $Y=1.87 $X2=0 $Y2=0
cc_90 N_A2_c_96_n N_B1_M1001_g 0.00259293f $X=1.095 $Y=1.745 $X2=0 $Y2=0
cc_91 A2 N_B1_M1001_g 0.00581352f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_92 A2 B1 0.0252378f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A2_c_98_n B1 3.06363e-19 $X=1.035 $Y=1.345 $X2=0 $Y2=0
cc_94 A2 N_B1_c_147_n 0.00244926f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_A2_c_98_n N_B1_c_147_n 0.0177911f $X=1.035 $Y=1.345 $X2=0 $Y2=0
cc_96 A2 N_A_244_409#_M1002_d 0.0089034f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A2_c_99_n N_A_244_409#_c_194_n 0.00354297f $X=1.095 $Y=1.87 $X2=0 $Y2=0
cc_98 N_A2_M1002_g N_A_244_409#_c_194_n 0.00416482f $X=1.095 $Y=2.545 $X2=0
+ $Y2=0
cc_99 A2 N_A_244_409#_c_194_n 0.081944f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A2_M1003_g N_A_244_409#_c_187_n 2.16745e-19 $X=1.005 $Y=0.495 $X2=0
+ $Y2=0
cc_101 N_A2_c_99_n N_A_244_409#_c_196_n 4.20151e-19 $X=1.095 $Y=1.87 $X2=0 $Y2=0
cc_102 A2 N_A_244_409#_c_196_n 0.0147551f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A2_M1002_g N_VPWR_c_257_n 0.00216219f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_104 A2 N_VPWR_c_257_n 0.0382647f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A2_M1002_g N_VPWR_c_259_n 0.00595064f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_106 A2 N_VPWR_c_259_n 0.0119421f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A2_M1002_g N_VPWR_c_255_n 0.00804775f $X=1.095 $Y=2.545 $X2=0 $Y2=0
cc_108 A2 N_VPWR_c_255_n 0.0142002f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 A2 A_146_409# 0.0104886f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_110 N_A2_M1003_g N_A_27_57#_c_314_n 6.46493e-19 $X=1.005 $Y=0.495 $X2=0 $Y2=0
cc_111 N_A2_M1003_g N_A_27_57#_c_315_n 0.0118052f $X=1.005 $Y=0.495 $X2=0 $Y2=0
cc_112 A2 N_A_27_57#_c_315_n 0.03535f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_113 N_A2_c_98_n N_A_27_57#_c_315_n 0.0013442f $X=1.035 $Y=1.345 $X2=0 $Y2=0
cc_114 N_A2_M1003_g N_A_27_57#_c_317_n 0.009671f $X=1.005 $Y=0.495 $X2=0 $Y2=0
cc_115 N_A2_M1003_g N_VGND_c_343_n 0.00456564f $X=1.005 $Y=0.495 $X2=0 $Y2=0
cc_116 N_A2_M1003_g N_VGND_c_346_n 0.00502664f $X=1.005 $Y=0.495 $X2=0 $Y2=0
cc_117 N_A2_M1003_g N_VGND_c_348_n 0.00592049f $X=1.005 $Y=0.495 $X2=0 $Y2=0
cc_118 N_B1_M1001_g N_A_244_409#_c_186_n 0.0221591f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_119 N_B1_M1001_g N_A_244_409#_c_194_n 0.0243264f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_120 N_B1_M1005_g N_A_244_409#_c_187_n 0.00957422f $X=1.515 $Y=0.495 $X2=0
+ $Y2=0
cc_121 N_B1_M1001_g N_A_244_409#_c_195_n 0.0214069f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_122 N_B1_M1001_g N_A_244_409#_c_196_n 0.0034891f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_123 B1 N_A_244_409#_c_196_n 0.026509f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B1_c_147_n N_A_244_409#_c_196_n 0.0023796f $X=1.925 $Y=1.34 $X2=0 $Y2=0
cc_125 N_B1_M1005_g N_A_244_409#_c_188_n 0.00474335f $X=1.515 $Y=0.495 $X2=0
+ $Y2=0
cc_126 N_B1_M1001_g N_A_244_409#_c_188_n 0.00889074f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_127 B1 N_A_244_409#_c_188_n 0.0225103f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B1_c_147_n N_A_244_409#_c_188_n 0.00904119f $X=1.925 $Y=1.34 $X2=0
+ $Y2=0
cc_129 N_B1_M1005_g N_A_244_409#_c_190_n 0.00631629f $X=1.515 $Y=0.495 $X2=0
+ $Y2=0
cc_130 B1 N_A_244_409#_c_190_n 0.0186377f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B1_c_147_n N_A_244_409#_c_190_n 0.00930368f $X=1.925 $Y=1.34 $X2=0
+ $Y2=0
cc_132 N_B1_c_147_n N_A_244_409#_c_191_n 3.13953e-19 $X=1.925 $Y=1.34 $X2=0
+ $Y2=0
cc_133 N_B1_c_147_n N_A_244_409#_c_192_n 0.0221591f $X=1.925 $Y=1.34 $X2=0 $Y2=0
cc_134 N_B1_M1001_g N_VPWR_c_258_n 0.0234358f $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_135 N_B1_M1001_g N_VPWR_c_259_n 0.00769046f $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_136 N_B1_M1001_g N_VPWR_c_255_n 0.013839f $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_137 N_B1_M1001_g N_X_c_291_n 2.08302e-19 $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_138 N_B1_M1005_g N_A_27_57#_c_315_n 0.00162595f $X=1.515 $Y=0.495 $X2=0 $Y2=0
cc_139 N_B1_M1005_g N_A_27_57#_c_317_n 0.00339679f $X=1.515 $Y=0.495 $X2=0 $Y2=0
cc_140 N_B1_M1005_g N_VGND_c_344_n 0.00258029f $X=1.515 $Y=0.495 $X2=0 $Y2=0
cc_141 N_B1_M1005_g N_VGND_c_346_n 0.00502664f $X=1.515 $Y=0.495 $X2=0 $Y2=0
cc_142 N_B1_M1005_g N_VGND_c_348_n 0.0105351f $X=1.515 $Y=0.495 $X2=0 $Y2=0
cc_143 N_A_244_409#_M1006_g N_VPWR_c_258_n 0.0246202f $X=2.455 $Y=2.545 $X2=0
+ $Y2=0
cc_144 N_A_244_409#_c_194_n N_VPWR_c_258_n 0.0678674f $X=1.66 $Y=2.19 $X2=0
+ $Y2=0
cc_145 N_A_244_409#_c_195_n N_VPWR_c_258_n 0.0131386f $X=2.005 $Y=1.77 $X2=0
+ $Y2=0
cc_146 N_A_244_409#_c_194_n N_VPWR_c_259_n 0.0220321f $X=1.66 $Y=2.19 $X2=0
+ $Y2=0
cc_147 N_A_244_409#_M1006_g N_VPWR_c_260_n 0.00769046f $X=2.455 $Y=2.545 $X2=0
+ $Y2=0
cc_148 N_A_244_409#_M1006_g N_VPWR_c_255_n 0.0143431f $X=2.455 $Y=2.545 $X2=0
+ $Y2=0
cc_149 N_A_244_409#_c_194_n N_VPWR_c_255_n 0.0125808f $X=1.66 $Y=2.19 $X2=0
+ $Y2=0
cc_150 N_A_244_409#_M1006_g N_X_c_291_n 0.013875f $X=2.455 $Y=2.545 $X2=0 $Y2=0
cc_151 N_A_244_409#_M1006_g N_X_c_292_n 0.00363507f $X=2.455 $Y=2.545 $X2=0
+ $Y2=0
cc_152 N_A_244_409#_c_186_n N_X_c_292_n 3.40936e-19 $X=2.507 $Y=1.495 $X2=0
+ $Y2=0
cc_153 N_A_244_409#_c_191_n N_X_c_292_n 0.00281512f $X=2.52 $Y=0.99 $X2=0 $Y2=0
cc_154 N_A_244_409#_M1006_g N_X_c_290_n 0.0182681f $X=2.455 $Y=2.545 $X2=0 $Y2=0
cc_155 N_A_244_409#_M1007_g N_X_c_290_n 0.00185044f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_156 N_A_244_409#_M1008_g N_X_c_290_n 0.0126368f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A_244_409#_c_185_n N_X_c_290_n 0.00644564f $X=2.865 $Y=0.9 $X2=0 $Y2=0
cc_158 N_A_244_409#_c_191_n N_X_c_290_n 0.0422161f $X=2.52 $Y=0.99 $X2=0 $Y2=0
cc_159 N_A_244_409#_c_192_n N_X_c_290_n 0.0112572f $X=2.52 $Y=0.99 $X2=0 $Y2=0
cc_160 N_A_244_409#_c_190_n N_A_27_57#_c_315_n 0.0143385f $X=2.175 $Y=0.91 $X2=0
+ $Y2=0
cc_161 N_A_244_409#_c_187_n N_A_27_57#_c_317_n 0.0255455f $X=1.73 $Y=0.495 $X2=0
+ $Y2=0
cc_162 N_A_244_409#_M1007_g N_VGND_c_344_n 0.0132554f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_163 N_A_244_409#_M1008_g N_VGND_c_344_n 0.0023851f $X=2.865 $Y=0.445 $X2=0
+ $Y2=0
cc_164 N_A_244_409#_c_185_n N_VGND_c_344_n 0.00108079f $X=2.865 $Y=0.9 $X2=0
+ $Y2=0
cc_165 N_A_244_409#_c_187_n N_VGND_c_344_n 0.025619f $X=1.73 $Y=0.495 $X2=0
+ $Y2=0
cc_166 N_A_244_409#_c_190_n N_VGND_c_344_n 0.0175357f $X=2.175 $Y=0.91 $X2=0
+ $Y2=0
cc_167 N_A_244_409#_c_191_n N_VGND_c_344_n 0.00549803f $X=2.52 $Y=0.99 $X2=0
+ $Y2=0
cc_168 N_A_244_409#_c_187_n N_VGND_c_346_n 0.0217141f $X=1.73 $Y=0.495 $X2=0
+ $Y2=0
cc_169 N_A_244_409#_M1007_g N_VGND_c_347_n 0.00486043f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_170 N_A_244_409#_M1008_g N_VGND_c_347_n 0.00550269f $X=2.865 $Y=0.445 $X2=0
+ $Y2=0
cc_171 N_A_244_409#_M1007_g N_VGND_c_348_n 0.00437501f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_172 N_A_244_409#_M1008_g N_VGND_c_348_n 0.0109068f $X=2.865 $Y=0.445 $X2=0
+ $Y2=0
cc_173 N_A_244_409#_c_185_n N_VGND_c_348_n 3.08405e-19 $X=2.865 $Y=0.9 $X2=0
+ $Y2=0
cc_174 N_A_244_409#_c_187_n N_VGND_c_348_n 0.0125146f $X=1.73 $Y=0.495 $X2=0
+ $Y2=0
cc_175 N_A_244_409#_c_190_n N_VGND_c_348_n 0.00891189f $X=2.175 $Y=0.91 $X2=0
+ $Y2=0
cc_176 N_A_244_409#_c_191_n N_VGND_c_348_n 0.00817171f $X=2.52 $Y=0.99 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_258_n N_X_c_291_n 0.0520536f $X=2.19 $Y=2.2 $X2=0 $Y2=0
cc_178 N_VPWR_c_260_n N_X_c_291_n 0.0220321f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_255_n N_X_c_291_n 0.0125808f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_180 N_VPWR_c_258_n N_X_c_292_n 0.0117799f $X=2.19 $Y=2.2 $X2=0 $Y2=0
cc_181 N_VPWR_c_258_n N_X_c_290_n 0.00225454f $X=2.19 $Y=2.2 $X2=0 $Y2=0
cc_182 N_X_c_290_n N_VGND_c_344_n 0.0117101f $X=3.08 $Y=0.445 $X2=0 $Y2=0
cc_183 N_X_c_290_n N_VGND_c_347_n 0.0167325f $X=3.08 $Y=0.445 $X2=0 $Y2=0
cc_184 N_X_M1008_d N_VGND_c_348_n 0.00234843f $X=2.94 $Y=0.235 $X2=0 $Y2=0
cc_185 N_X_c_290_n N_VGND_c_348_n 0.0123752f $X=3.08 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A_27_57#_c_314_n N_VGND_c_343_n 0.0143477f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_187 N_A_27_57#_c_315_n N_VGND_c_343_n 0.019034f $X=1.055 $Y=0.91 $X2=0 $Y2=0
cc_188 N_A_27_57#_c_317_n N_VGND_c_343_n 0.0143477f $X=1.22 $Y=0.495 $X2=0 $Y2=0
cc_189 N_A_27_57#_c_314_n N_VGND_c_345_n 0.0220321f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_190 N_A_27_57#_c_317_n N_VGND_c_346_n 0.0220321f $X=1.22 $Y=0.495 $X2=0 $Y2=0
cc_191 N_A_27_57#_c_314_n N_VGND_c_348_n 0.0125808f $X=0.28 $Y=0.495 $X2=0 $Y2=0
cc_192 N_A_27_57#_c_315_n N_VGND_c_348_n 0.011685f $X=1.055 $Y=0.91 $X2=0 $Y2=0
cc_193 N_A_27_57#_c_317_n N_VGND_c_348_n 0.0125808f $X=1.22 $Y=0.495 $X2=0 $Y2=0
cc_194 N_VGND_c_348_n A_516_47# 0.00567374f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
