* File: sky130_fd_sc_lp__dlymetal6s6s_1.pxi.spice
* Created: Fri Aug 28 10:31:23 2020
* 
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A N_A_M1008_g N_A_M1010_g A N_A_c_95_n
+ N_A_c_96_n PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_27_131# N_A_27_131#_M1008_s
+ N_A_27_131#_M1010_s N_A_27_131#_M1006_g N_A_27_131#_M1001_g
+ N_A_27_131#_c_123_n N_A_27_131#_c_136_n N_A_27_131#_c_124_n
+ N_A_27_131#_c_125_n N_A_27_131#_c_126_n N_A_27_131#_c_130_n
+ N_A_27_131#_c_127_n PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_27_131#
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_208_47# N_A_208_47#_M1006_d
+ N_A_208_47#_M1001_d N_A_208_47#_M1011_g N_A_208_47#_M1005_g
+ N_A_208_47#_c_183_n N_A_208_47#_c_184_n N_A_208_47#_c_185_n
+ N_A_208_47#_c_186_n N_A_208_47#_c_191_n N_A_208_47#_c_187_n
+ N_A_208_47#_c_188_n N_A_208_47#_c_189_n N_A_208_47#_c_193_n
+ PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_208_47#
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_315_131# N_A_315_131#_M1011_s
+ N_A_315_131#_M1005_s N_A_315_131#_M1002_g N_A_315_131#_M1000_g
+ N_A_315_131#_c_247_n N_A_315_131#_c_260_n N_A_315_131#_c_248_n
+ N_A_315_131#_c_249_n N_A_315_131#_c_250_n N_A_315_131#_c_254_n
+ N_A_315_131#_c_251_n PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_315_131#
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_496_47# N_A_496_47#_M1002_d
+ N_A_496_47#_M1000_d N_A_496_47#_M1004_g N_A_496_47#_M1003_g
+ N_A_496_47#_c_311_n N_A_496_47#_c_312_n N_A_496_47#_c_313_n
+ N_A_496_47#_c_314_n N_A_496_47#_c_319_n N_A_496_47#_c_315_n
+ N_A_496_47#_c_316_n N_A_496_47#_c_317_n N_A_496_47#_c_321_n
+ PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_496_47#
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_603_131# N_A_603_131#_M1004_s
+ N_A_603_131#_M1003_s N_A_603_131#_M1009_g N_A_603_131#_M1007_g
+ N_A_603_131#_c_376_n N_A_603_131#_c_389_n N_A_603_131#_c_377_n
+ N_A_603_131#_c_378_n N_A_603_131#_c_379_n N_A_603_131#_c_383_n
+ N_A_603_131#_c_380_n PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%A_603_131#
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%VPWR N_VPWR_M1010_d N_VPWR_M1005_d
+ N_VPWR_M1003_d N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n VPWR
+ N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_438_n
+ N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_449_n VPWR
+ PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%VPWR
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%X N_X_M1009_d N_X_M1007_d N_X_c_489_n
+ N_X_c_492_n N_X_c_490_n N_X_c_491_n X N_X_c_494_n N_X_c_503_n N_X_c_495_n X
+ PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%X
x_PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%VGND N_VGND_M1008_d N_VGND_M1011_d
+ N_VGND_M1004_d N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n VGND
+ N_VGND_c_539_n N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n
+ N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n VGND
+ PM_SKY130_FD_SC_LP__DLYMETAL6S6S_1%VGND
cc_1 VNB N_A_M1008_g 0.0305881f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.865
cc_2 VNB N_A_M1010_g 0.00321153f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.045
cc_3 VNB N_A_c_95_n 0.0367407f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_4 VNB N_A_c_96_n 0.0142689f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_5 VNB N_A_27_131#_M1006_g 0.0249043f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_131#_M1001_g 0.00287706f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_7 VNB N_A_27_131#_c_123_n 0.0060589f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.605
cc_8 VNB N_A_27_131#_c_124_n 0.00344094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_131#_c_125_n 6.31025e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_131#_c_126_n 0.0201662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_131#_c_127_n 0.0365531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_208_47#_M1011_g 0.0256351f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_A_208_47#_M1005_g 0.00318199f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_14 VNB N_A_208_47#_c_183_n 0.00995534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_208_47#_c_184_n 0.00560895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_208_47#_c_185_n 0.0192779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_208_47#_c_186_n 0.0314719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_208_47#_c_187_n 0.00125812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_208_47#_c_188_n 0.00456899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_208_47#_c_189_n 0.00344243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_315_131#_M1002_g 0.0249043f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_315_131#_M1000_g 0.00287706f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_23 VNB N_A_315_131#_c_247_n 0.006059f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.605
cc_24 VNB N_A_315_131#_c_248_n 0.00343604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_315_131#_c_249_n 8.06932e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_315_131#_c_250_n 0.00696695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_315_131#_c_251_n 0.0365429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_496_47#_M1004_g 0.0256351f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_A_496_47#_M1003_g 0.00318199f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_30 VNB N_A_496_47#_c_311_n 0.00995534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_496_47#_c_312_n 0.00560895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_496_47#_c_313_n 0.0192779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_496_47#_c_314_n 0.0314884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_496_47#_c_315_n 0.00125812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_496_47#_c_316_n 0.00456899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_496_47#_c_317_n 0.00343052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_603_131#_M1009_g 0.0249043f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_A_603_131#_M1007_g 0.00287706f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_39 VNB N_A_603_131#_c_376_n 0.006059f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.605
cc_40 VNB N_A_603_131#_c_377_n 0.00343604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_603_131#_c_378_n 8.06932e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_603_131#_c_379_n 0.00696695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_603_131#_c_380_n 0.0350929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_438_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_489_n 0.0264688f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_X_c_490_n 0.0271579f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_47 VNB N_X_c_491_n 0.00853408f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.605
cc_48 VNB N_VGND_c_536_n 0.0152805f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.44
cc_49 VNB N_VGND_c_537_n 0.00982248f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.44
cc_50 VNB N_VGND_c_538_n 0.00982248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_539_n 0.0196132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_540_n 0.0305918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_541_n 0.0305918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_542_n 0.0152818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_543_n 0.268562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_544_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_545_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_546_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_A_M1010_g 0.0323158f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.045
cc_60 VPB N_A_c_96_n 0.00704613f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_61 VPB N_A_27_131#_M1001_g 0.0265052f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_62 VPB N_A_27_131#_c_125_n 0.00285445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_27_131#_c_130_n 0.013938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_208_47#_M1005_g 0.0253109f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_65 VPB N_A_208_47#_c_191_n 0.00506407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_208_47#_c_187_n 0.00461232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_208_47#_c_193_n 0.0168145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_315_131#_M1000_g 0.0265052f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_69 VPB N_A_315_131#_c_249_n 0.00324934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_315_131#_c_254_n 0.00354173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_496_47#_M1003_g 0.0253109f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_72 VPB N_A_496_47#_c_319_n 0.00506407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_496_47#_c_315_n 0.00461232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_496_47#_c_321_n 0.0168145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_603_131#_M1007_g 0.0265052f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_76 VPB N_A_603_131#_c_378_n 0.00324934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_603_131#_c_383_n 0.00354173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_439_n 0.0332367f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_79 VPB N_VPWR_c_440_n 0.0186008f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.44
cc_80 VPB N_VPWR_c_441_n 0.0186008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_442_n 0.0207592f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_443_n 0.0336503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_444_n 0.0336503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_445_n 0.0171944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_438_n 0.121279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_447_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_448_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_449_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_X_c_492_n 0.00905053f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.44
cc_90 VPB N_X_c_490_n 0.00854167f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_91 VPB N_X_c_494_n 0.0424779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_X_c_495_n 0.0692555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 N_A_M1008_g N_A_27_131#_M1006_g 0.0169752f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_94 N_A_M1010_g N_A_27_131#_M1001_g 0.0228128f $X=0.475 $Y=2.045 $X2=0 $Y2=0
cc_95 N_A_M1008_g N_A_27_131#_c_123_n 0.0140155f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_96 N_A_c_95_n N_A_27_131#_c_123_n 2.34881e-19 $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_97 N_A_c_96_n N_A_27_131#_c_123_n 0.0117414f $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_98 N_A_M1010_g N_A_27_131#_c_136_n 0.0123302f $X=0.475 $Y=2.045 $X2=0 $Y2=0
cc_99 N_A_M1008_g N_A_27_131#_c_124_n 0.00527832f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_100 N_A_c_96_n N_A_27_131#_c_124_n 0.0233614f $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_101 N_A_M1010_g N_A_27_131#_c_125_n 0.00458359f $X=0.475 $Y=2.045 $X2=0 $Y2=0
cc_102 N_A_c_96_n N_A_27_131#_c_125_n 0.0122398f $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_103 N_A_M1008_g N_A_27_131#_c_126_n 0.00158998f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_104 N_A_c_95_n N_A_27_131#_c_126_n 0.00407112f $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_105 N_A_c_96_n N_A_27_131#_c_126_n 0.0246121f $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_106 N_A_M1010_g N_A_27_131#_c_130_n 0.00307109f $X=0.475 $Y=2.045 $X2=0 $Y2=0
cc_107 N_A_c_95_n N_A_27_131#_c_130_n 7.93987e-19 $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_108 N_A_c_96_n N_A_27_131#_c_130_n 0.0338762f $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_109 N_A_M1008_g N_A_27_131#_c_127_n 0.0214866f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_110 N_A_c_96_n N_A_27_131#_c_127_n 3.32537e-19 $X=0.385 $Y=1.44 $X2=0 $Y2=0
cc_111 N_A_M1010_g N_VPWR_c_439_n 0.00154026f $X=0.475 $Y=2.045 $X2=0 $Y2=0
cc_112 N_A_M1008_g N_VGND_c_536_n 0.00447327f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_113 N_A_M1008_g N_VGND_c_539_n 0.00399858f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_114 N_A_M1008_g N_VGND_c_543_n 0.0046122f $X=0.475 $Y=0.865 $X2=0 $Y2=0
cc_115 N_A_27_131#_M1006_g N_A_208_47#_c_184_n 0.00390403f $X=0.965 $Y=0.655
+ $X2=0 $Y2=0
cc_116 N_A_27_131#_c_124_n N_A_208_47#_c_184_n 0.0128275f $X=0.805 $Y=1.605
+ $X2=0 $Y2=0
cc_117 N_A_27_131#_c_127_n N_A_208_47#_c_184_n 8.33413e-19 $X=0.925 $Y=1.44
+ $X2=0 $Y2=0
cc_118 N_A_27_131#_c_127_n N_A_208_47#_c_186_n 0.00467288f $X=0.925 $Y=1.44
+ $X2=0 $Y2=0
cc_119 N_A_27_131#_M1001_g N_A_208_47#_c_191_n 0.00323486f $X=0.965 $Y=2.465
+ $X2=0 $Y2=0
cc_120 N_A_27_131#_c_136_n N_A_208_47#_c_191_n 0.0113721f $X=0.72 $Y=2.047 $X2=0
+ $Y2=0
cc_121 N_A_27_131#_M1001_g N_A_208_47#_c_187_n 0.00485767f $X=0.965 $Y=2.465
+ $X2=0 $Y2=0
cc_122 N_A_27_131#_c_125_n N_A_208_47#_c_187_n 0.0118249f $X=0.805 $Y=1.935
+ $X2=0 $Y2=0
cc_123 N_A_27_131#_c_124_n N_A_208_47#_c_189_n 0.0243592f $X=0.805 $Y=1.605
+ $X2=0 $Y2=0
cc_124 N_A_27_131#_c_127_n N_A_208_47#_c_189_n 0.00350342f $X=0.925 $Y=1.44
+ $X2=0 $Y2=0
cc_125 N_A_27_131#_M1001_g N_A_208_47#_c_193_n 0.00431951f $X=0.965 $Y=2.465
+ $X2=0 $Y2=0
cc_126 N_A_27_131#_c_136_n N_A_208_47#_c_193_n 0.00643722f $X=0.72 $Y=2.047
+ $X2=0 $Y2=0
cc_127 N_A_27_131#_c_124_n N_A_208_47#_c_193_n 0.00182968f $X=0.805 $Y=1.605
+ $X2=0 $Y2=0
cc_128 N_A_27_131#_c_125_n N_A_208_47#_c_193_n 4.37025e-19 $X=0.805 $Y=1.935
+ $X2=0 $Y2=0
cc_129 N_A_27_131#_c_127_n N_A_208_47#_c_193_n 4.68851e-19 $X=0.925 $Y=1.44
+ $X2=0 $Y2=0
cc_130 N_A_27_131#_c_136_n N_VPWR_M1010_d 0.00814393f $X=0.72 $Y=2.047 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_27_131#_c_125_n N_VPWR_M1010_d 0.00171264f $X=0.805 $Y=1.935
+ $X2=-0.19 $Y2=-0.245
cc_132 N_A_27_131#_M1001_g N_VPWR_c_439_n 0.00623246f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_27_131#_c_136_n N_VPWR_c_439_n 0.0204871f $X=0.72 $Y=2.047 $X2=0
+ $Y2=0
cc_134 N_A_27_131#_M1001_g N_VPWR_c_443_n 0.00585385f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_27_131#_M1001_g N_VPWR_c_438_n 0.0131218f $X=0.965 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_27_131#_M1001_g N_X_c_495_n 0.00551213f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_27_131#_c_123_n N_VGND_M1008_d 0.00119058f $X=0.72 $Y=1.06 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_27_131#_c_124_n N_VGND_M1008_d 0.00176358f $X=0.805 $Y=1.605
+ $X2=-0.19 $Y2=-0.245
cc_139 N_A_27_131#_M1006_g N_VGND_c_536_n 0.0129337f $X=0.965 $Y=0.655 $X2=0
+ $Y2=0
cc_140 N_A_27_131#_c_123_n N_VGND_c_536_n 0.00915704f $X=0.72 $Y=1.06 $X2=0
+ $Y2=0
cc_141 N_A_27_131#_c_124_n N_VGND_c_536_n 0.0110081f $X=0.805 $Y=1.605 $X2=0
+ $Y2=0
cc_142 N_A_27_131#_c_127_n N_VGND_c_536_n 4.51333e-19 $X=0.925 $Y=1.44 $X2=0
+ $Y2=0
cc_143 N_A_27_131#_c_126_n N_VGND_c_539_n 0.00444585f $X=0.26 $Y=0.865 $X2=0
+ $Y2=0
cc_144 N_A_27_131#_M1006_g N_VGND_c_540_n 0.00486043f $X=0.965 $Y=0.655 $X2=0
+ $Y2=0
cc_145 N_A_27_131#_M1006_g N_VGND_c_543_n 0.00954696f $X=0.965 $Y=0.655 $X2=0
+ $Y2=0
cc_146 N_A_27_131#_c_126_n N_VGND_c_543_n 0.00830526f $X=0.26 $Y=0.865 $X2=0
+ $Y2=0
cc_147 N_A_208_47#_M1011_g N_A_315_131#_M1002_g 0.0169752f $X=1.915 $Y=0.865
+ $X2=0 $Y2=0
cc_148 N_A_208_47#_M1005_g N_A_315_131#_M1000_g 0.0235709f $X=1.915 $Y=2.045
+ $X2=0 $Y2=0
cc_149 N_A_208_47#_M1011_g N_A_315_131#_c_247_n 0.0140353f $X=1.915 $Y=0.865
+ $X2=0 $Y2=0
cc_150 N_A_208_47#_c_185_n N_A_315_131#_c_247_n 0.0113458f $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_151 N_A_208_47#_c_186_n N_A_315_131#_c_247_n 2.3501e-19 $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_152 N_A_208_47#_M1005_g N_A_315_131#_c_260_n 0.0107574f $X=1.915 $Y=2.045
+ $X2=0 $Y2=0
cc_153 N_A_208_47#_M1011_g N_A_315_131#_c_248_n 0.00368817f $X=1.915 $Y=0.865
+ $X2=0 $Y2=0
cc_154 N_A_208_47#_c_185_n N_A_315_131#_c_248_n 0.0240545f $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_155 N_A_208_47#_c_186_n N_A_315_131#_c_248_n 9.23612e-19 $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_156 N_A_208_47#_M1005_g N_A_315_131#_c_249_n 0.00613959f $X=1.915 $Y=2.045
+ $X2=0 $Y2=0
cc_157 N_A_208_47#_M1011_g N_A_315_131#_c_250_n 0.00158998f $X=1.915 $Y=0.865
+ $X2=0 $Y2=0
cc_158 N_A_208_47#_c_183_n N_A_315_131#_c_250_n 0.0338024f $X=1.18 $Y=0.42 $X2=0
+ $Y2=0
cc_159 N_A_208_47#_c_185_n N_A_315_131#_c_250_n 0.0241515f $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_160 N_A_208_47#_c_186_n N_A_315_131#_c_250_n 0.00407385f $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_161 N_A_208_47#_M1005_g N_A_315_131#_c_254_n 0.00262595f $X=1.915 $Y=2.045
+ $X2=0 $Y2=0
cc_162 N_A_208_47#_c_185_n N_A_315_131#_c_254_n 0.0217491f $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_163 N_A_208_47#_c_186_n N_A_315_131#_c_254_n 0.00360834f $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_164 N_A_208_47#_c_191_n N_A_315_131#_c_254_n 0.0247421f $X=1.205 $Y=1.98
+ $X2=0 $Y2=0
cc_165 N_A_208_47#_c_193_n N_A_315_131#_c_254_n 0.00180002f $X=1.18 $Y=2 $X2=0
+ $Y2=0
cc_166 N_A_208_47#_M1011_g N_A_315_131#_c_251_n 0.0221797f $X=1.915 $Y=0.865
+ $X2=0 $Y2=0
cc_167 N_A_208_47#_c_185_n N_A_315_131#_c_251_n 3.28937e-19 $X=1.825 $Y=1.44
+ $X2=0 $Y2=0
cc_168 N_A_208_47#_M1005_g N_VPWR_c_440_n 7.16233e-19 $X=1.915 $Y=2.045 $X2=0
+ $Y2=0
cc_169 N_A_208_47#_c_193_n N_VPWR_c_440_n 0.0205592f $X=1.18 $Y=2 $X2=0 $Y2=0
cc_170 N_A_208_47#_c_193_n N_VPWR_c_443_n 0.0190565f $X=1.18 $Y=2 $X2=0 $Y2=0
cc_171 N_A_208_47#_M1001_d N_VPWR_c_438_n 0.00284733f $X=1.04 $Y=1.835 $X2=0
+ $Y2=0
cc_172 N_A_208_47#_c_193_n N_VPWR_c_438_n 0.0111968f $X=1.18 $Y=2 $X2=0 $Y2=0
cc_173 N_A_208_47#_M1001_d N_X_c_495_n 8.51489e-19 $X=1.04 $Y=1.835 $X2=0 $Y2=0
cc_174 N_A_208_47#_M1005_g N_X_c_495_n 0.00459273f $X=1.915 $Y=2.045 $X2=0 $Y2=0
cc_175 N_A_208_47#_c_193_n N_X_c_495_n 0.0627285f $X=1.18 $Y=2 $X2=0 $Y2=0
cc_176 N_A_208_47#_M1011_g N_VGND_c_537_n 0.00283805f $X=1.915 $Y=0.865 $X2=0
+ $Y2=0
cc_177 N_A_208_47#_c_183_n N_VGND_c_537_n 0.0131216f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_178 N_A_208_47#_M1011_g N_VGND_c_540_n 0.00399858f $X=1.915 $Y=0.865 $X2=0
+ $Y2=0
cc_179 N_A_208_47#_c_183_n N_VGND_c_540_n 0.0181695f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_180 N_A_208_47#_M1006_d N_VGND_c_543_n 0.00371702f $X=1.04 $Y=0.235 $X2=0
+ $Y2=0
cc_181 N_A_208_47#_M1011_g N_VGND_c_543_n 0.0046122f $X=1.915 $Y=0.865 $X2=0
+ $Y2=0
cc_182 N_A_208_47#_c_183_n N_VGND_c_543_n 0.0102248f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_183 N_A_315_131#_M1002_g N_A_496_47#_c_312_n 0.00390403f $X=2.405 $Y=0.655
+ $X2=0 $Y2=0
cc_184 N_A_315_131#_c_248_n N_A_496_47#_c_312_n 0.0128275f $X=2.245 $Y=1.605
+ $X2=0 $Y2=0
cc_185 N_A_315_131#_c_251_n N_A_496_47#_c_312_n 8.33413e-19 $X=2.365 $Y=1.44
+ $X2=0 $Y2=0
cc_186 N_A_315_131#_c_251_n N_A_496_47#_c_314_n 0.00467288f $X=2.365 $Y=1.44
+ $X2=0 $Y2=0
cc_187 N_A_315_131#_M1000_g N_A_496_47#_c_319_n 0.00323475f $X=2.405 $Y=2.465
+ $X2=0 $Y2=0
cc_188 N_A_315_131#_c_260_n N_A_496_47#_c_319_n 0.0131905f $X=2.16 $Y=2.027
+ $X2=0 $Y2=0
cc_189 N_A_315_131#_M1000_g N_A_496_47#_c_315_n 0.00485767f $X=2.405 $Y=2.465
+ $X2=0 $Y2=0
cc_190 N_A_315_131#_c_249_n N_A_496_47#_c_315_n 0.0118249f $X=2.245 $Y=1.895
+ $X2=0 $Y2=0
cc_191 N_A_315_131#_c_248_n N_A_496_47#_c_317_n 0.0243592f $X=2.245 $Y=1.605
+ $X2=0 $Y2=0
cc_192 N_A_315_131#_c_251_n N_A_496_47#_c_317_n 0.00350342f $X=2.365 $Y=1.44
+ $X2=0 $Y2=0
cc_193 N_A_315_131#_M1000_g N_A_496_47#_c_321_n 0.00431945f $X=2.405 $Y=2.465
+ $X2=0 $Y2=0
cc_194 N_A_315_131#_c_260_n N_A_496_47#_c_321_n 0.00688633f $X=2.16 $Y=2.027
+ $X2=0 $Y2=0
cc_195 N_A_315_131#_c_248_n N_A_496_47#_c_321_n 0.00182968f $X=2.245 $Y=1.605
+ $X2=0 $Y2=0
cc_196 N_A_315_131#_c_251_n N_A_496_47#_c_321_n 4.68851e-19 $X=2.365 $Y=1.44
+ $X2=0 $Y2=0
cc_197 N_A_315_131#_c_260_n N_VPWR_M1005_d 0.00823473f $X=2.16 $Y=2.027 $X2=0
+ $Y2=0
cc_198 N_A_315_131#_c_249_n N_VPWR_M1005_d 0.00102067f $X=2.245 $Y=1.895 $X2=0
+ $Y2=0
cc_199 N_A_315_131#_M1000_g N_VPWR_c_440_n 0.00647425f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_315_131#_c_260_n N_VPWR_c_440_n 0.0173442f $X=2.16 $Y=2.027 $X2=0
+ $Y2=0
cc_201 N_A_315_131#_M1000_g N_VPWR_c_444_n 0.00585385f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_A_315_131#_M1000_g N_VPWR_c_438_n 0.0131218f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_A_315_131#_M1000_g N_X_c_495_n 0.00982165f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_315_131#_c_260_n N_X_c_495_n 0.0153371f $X=2.16 $Y=2.027 $X2=0 $Y2=0
cc_205 N_A_315_131#_c_254_n N_X_c_495_n 0.0173796f $X=1.865 $Y=2.06 $X2=0 $Y2=0
cc_206 N_A_315_131#_c_247_n N_VGND_M1011_d 0.00119058f $X=2.16 $Y=1.06 $X2=0
+ $Y2=0
cc_207 N_A_315_131#_c_248_n N_VGND_M1011_d 0.00176358f $X=2.245 $Y=1.605 $X2=0
+ $Y2=0
cc_208 N_A_315_131#_M1002_g N_VGND_c_537_n 0.0129337f $X=2.405 $Y=0.655 $X2=0
+ $Y2=0
cc_209 N_A_315_131#_c_247_n N_VGND_c_537_n 0.00915704f $X=2.16 $Y=1.06 $X2=0
+ $Y2=0
cc_210 N_A_315_131#_c_248_n N_VGND_c_537_n 0.0110081f $X=2.245 $Y=1.605 $X2=0
+ $Y2=0
cc_211 N_A_315_131#_c_251_n N_VGND_c_537_n 4.51333e-19 $X=2.365 $Y=1.44 $X2=0
+ $Y2=0
cc_212 N_A_315_131#_c_250_n N_VGND_c_540_n 0.00444585f $X=1.7 $Y=0.865 $X2=0
+ $Y2=0
cc_213 N_A_315_131#_M1002_g N_VGND_c_541_n 0.00486043f $X=2.405 $Y=0.655 $X2=0
+ $Y2=0
cc_214 N_A_315_131#_M1002_g N_VGND_c_543_n 0.00954696f $X=2.405 $Y=0.655 $X2=0
+ $Y2=0
cc_215 N_A_315_131#_c_250_n N_VGND_c_543_n 0.00830526f $X=1.7 $Y=0.865 $X2=0
+ $Y2=0
cc_216 N_A_496_47#_M1004_g N_A_603_131#_M1009_g 0.0169752f $X=3.355 $Y=0.865
+ $X2=0 $Y2=0
cc_217 N_A_496_47#_M1003_g N_A_603_131#_M1007_g 0.0235709f $X=3.355 $Y=2.045
+ $X2=0 $Y2=0
cc_218 N_A_496_47#_M1004_g N_A_603_131#_c_376_n 0.0140353f $X=3.355 $Y=0.865
+ $X2=0 $Y2=0
cc_219 N_A_496_47#_c_313_n N_A_603_131#_c_376_n 0.0113458f $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_220 N_A_496_47#_c_314_n N_A_603_131#_c_376_n 2.3501e-19 $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_221 N_A_496_47#_M1003_g N_A_603_131#_c_389_n 0.0107574f $X=3.355 $Y=2.045
+ $X2=0 $Y2=0
cc_222 N_A_496_47#_M1004_g N_A_603_131#_c_377_n 0.00368817f $X=3.355 $Y=0.865
+ $X2=0 $Y2=0
cc_223 N_A_496_47#_c_313_n N_A_603_131#_c_377_n 0.0240545f $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_224 N_A_496_47#_c_314_n N_A_603_131#_c_377_n 9.23612e-19 $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_225 N_A_496_47#_M1003_g N_A_603_131#_c_378_n 0.00613959f $X=3.355 $Y=2.045
+ $X2=0 $Y2=0
cc_226 N_A_496_47#_M1004_g N_A_603_131#_c_379_n 0.00158998f $X=3.355 $Y=0.865
+ $X2=0 $Y2=0
cc_227 N_A_496_47#_c_311_n N_A_603_131#_c_379_n 0.0338024f $X=2.62 $Y=0.42 $X2=0
+ $Y2=0
cc_228 N_A_496_47#_c_313_n N_A_603_131#_c_379_n 0.0241515f $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_229 N_A_496_47#_c_314_n N_A_603_131#_c_379_n 0.00407385f $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_230 N_A_496_47#_M1003_g N_A_603_131#_c_383_n 0.00259526f $X=3.355 $Y=2.045
+ $X2=0 $Y2=0
cc_231 N_A_496_47#_c_313_n N_A_603_131#_c_383_n 0.0217491f $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_232 N_A_496_47#_c_314_n N_A_603_131#_c_383_n 0.00360834f $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_233 N_A_496_47#_c_319_n N_A_603_131#_c_383_n 0.0247421f $X=2.645 $Y=1.98
+ $X2=0 $Y2=0
cc_234 N_A_496_47#_c_321_n N_A_603_131#_c_383_n 0.00180002f $X=2.62 $Y=2 $X2=0
+ $Y2=0
cc_235 N_A_496_47#_M1004_g N_A_603_131#_c_380_n 0.0221773f $X=3.355 $Y=0.865
+ $X2=0 $Y2=0
cc_236 N_A_496_47#_c_313_n N_A_603_131#_c_380_n 3.28937e-19 $X=3.265 $Y=1.44
+ $X2=0 $Y2=0
cc_237 N_A_496_47#_c_321_n N_VPWR_c_440_n 0.00542266f $X=2.62 $Y=2 $X2=0 $Y2=0
cc_238 N_A_496_47#_M1003_g N_VPWR_c_441_n 7.16233e-19 $X=3.355 $Y=2.045 $X2=0
+ $Y2=0
cc_239 N_A_496_47#_c_321_n N_VPWR_c_441_n 0.0205592f $X=2.62 $Y=2 $X2=0 $Y2=0
cc_240 N_A_496_47#_c_321_n N_VPWR_c_444_n 0.0190565f $X=2.62 $Y=2 $X2=0 $Y2=0
cc_241 N_A_496_47#_M1000_d N_VPWR_c_438_n 0.00284733f $X=2.48 $Y=1.835 $X2=0
+ $Y2=0
cc_242 N_A_496_47#_c_321_n N_VPWR_c_438_n 0.0111968f $X=2.62 $Y=2 $X2=0 $Y2=0
cc_243 N_A_496_47#_M1003_g N_X_c_503_n 7.74848e-19 $X=3.355 $Y=2.045 $X2=0 $Y2=0
cc_244 N_A_496_47#_M1000_d N_X_c_495_n 8.51489e-19 $X=2.48 $Y=1.835 $X2=0 $Y2=0
cc_245 N_A_496_47#_M1003_g N_X_c_495_n 0.00459273f $X=3.355 $Y=2.045 $X2=0 $Y2=0
cc_246 N_A_496_47#_c_321_n N_X_c_495_n 0.0636761f $X=2.62 $Y=2 $X2=0 $Y2=0
cc_247 N_A_496_47#_M1004_g N_VGND_c_538_n 0.00283805f $X=3.355 $Y=0.865 $X2=0
+ $Y2=0
cc_248 N_A_496_47#_c_311_n N_VGND_c_538_n 0.0131216f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_249 N_A_496_47#_M1004_g N_VGND_c_541_n 0.00399858f $X=3.355 $Y=0.865 $X2=0
+ $Y2=0
cc_250 N_A_496_47#_c_311_n N_VGND_c_541_n 0.0181695f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_251 N_A_496_47#_M1002_d N_VGND_c_543_n 0.00371702f $X=2.48 $Y=0.235 $X2=0
+ $Y2=0
cc_252 N_A_496_47#_M1004_g N_VGND_c_543_n 0.0046122f $X=3.355 $Y=0.865 $X2=0
+ $Y2=0
cc_253 N_A_496_47#_c_311_n N_VGND_c_543_n 0.0102248f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_254 N_A_603_131#_c_389_n N_VPWR_M1003_d 0.00823473f $X=3.6 $Y=2.027 $X2=0
+ $Y2=0
cc_255 N_A_603_131#_c_378_n N_VPWR_M1003_d 0.00102067f $X=3.685 $Y=1.895 $X2=0
+ $Y2=0
cc_256 N_A_603_131#_M1007_g N_VPWR_c_441_n 0.00647425f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A_603_131#_c_389_n N_VPWR_c_441_n 0.0173442f $X=3.6 $Y=2.027 $X2=0
+ $Y2=0
cc_258 N_A_603_131#_M1007_g N_VPWR_c_445_n 0.00585385f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_259 N_A_603_131#_M1007_g N_VPWR_c_438_n 0.0127547f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_260 N_A_603_131#_M1007_g N_X_c_492_n 0.00424527f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_261 N_A_603_131#_c_389_n N_X_c_492_n 0.0132817f $X=3.6 $Y=2.027 $X2=0 $Y2=0
cc_262 N_A_603_131#_M1009_g N_X_c_490_n 0.00390868f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_263 N_A_603_131#_M1007_g N_X_c_490_n 0.00486724f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_603_131#_c_377_n N_X_c_490_n 0.0346309f $X=3.685 $Y=1.605 $X2=0 $Y2=0
cc_265 N_A_603_131#_c_378_n N_X_c_490_n 0.0118771f $X=3.685 $Y=1.895 $X2=0 $Y2=0
cc_266 N_A_603_131#_c_380_n N_X_c_490_n 0.00852845f $X=3.805 $Y=1.44 $X2=0 $Y2=0
cc_267 N_A_603_131#_M1007_g X 0.00369728f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A_603_131#_c_383_n N_X_c_494_n 6.80645e-19 $X=3.305 $Y=2.06 $X2=0 $Y2=0
cc_269 N_A_603_131#_M1007_g N_X_c_503_n 0.00723617f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_603_131#_c_389_n N_X_c_503_n 0.00718573f $X=3.6 $Y=2.027 $X2=0 $Y2=0
cc_271 N_A_603_131#_c_377_n N_X_c_503_n 0.00202145f $X=3.685 $Y=1.605 $X2=0
+ $Y2=0
cc_272 N_A_603_131#_c_383_n N_X_c_503_n 0.00127315f $X=3.305 $Y=2.06 $X2=0 $Y2=0
cc_273 N_A_603_131#_c_380_n N_X_c_503_n 5.34161e-19 $X=3.805 $Y=1.44 $X2=0 $Y2=0
cc_274 N_A_603_131#_M1007_g N_X_c_495_n 0.00568947f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_275 N_A_603_131#_c_389_n N_X_c_495_n 0.0153371f $X=3.6 $Y=2.027 $X2=0 $Y2=0
cc_276 N_A_603_131#_c_383_n N_X_c_495_n 0.0173796f $X=3.305 $Y=2.06 $X2=0 $Y2=0
cc_277 N_A_603_131#_c_376_n N_VGND_M1004_d 0.00119058f $X=3.6 $Y=1.06 $X2=0
+ $Y2=0
cc_278 N_A_603_131#_c_377_n N_VGND_M1004_d 0.00176358f $X=3.685 $Y=1.605 $X2=0
+ $Y2=0
cc_279 N_A_603_131#_M1009_g N_VGND_c_538_n 0.0129337f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_280 N_A_603_131#_c_376_n N_VGND_c_538_n 0.00915704f $X=3.6 $Y=1.06 $X2=0
+ $Y2=0
cc_281 N_A_603_131#_c_377_n N_VGND_c_538_n 0.0110081f $X=3.685 $Y=1.605 $X2=0
+ $Y2=0
cc_282 N_A_603_131#_c_380_n N_VGND_c_538_n 4.51333e-19 $X=3.805 $Y=1.44 $X2=0
+ $Y2=0
cc_283 N_A_603_131#_c_379_n N_VGND_c_541_n 0.00444585f $X=3.14 $Y=0.865 $X2=0
+ $Y2=0
cc_284 N_A_603_131#_M1009_g N_VGND_c_542_n 0.00486043f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_285 N_A_603_131#_M1009_g N_VGND_c_543_n 0.00917987f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_286 N_A_603_131#_c_379_n N_VGND_c_543_n 0.00830526f $X=3.14 $Y=0.865 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_438_n N_X_M1007_d 0.00284733f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_288 N_VPWR_c_441_n N_X_c_494_n 0.00542411f $X=3.63 $Y=2.495 $X2=0 $Y2=0
cc_289 N_VPWR_c_445_n N_X_c_494_n 0.019415f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_290 N_VPWR_c_438_n N_X_c_494_n 0.0113912f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_291 N_VPWR_M1005_d N_X_c_495_n 0.00241001f $X=1.99 $Y=1.835 $X2=0 $Y2=0
cc_292 N_VPWR_M1003_d N_X_c_495_n 0.00241001f $X=3.43 $Y=1.835 $X2=0 $Y2=0
cc_293 N_VPWR_c_439_n N_X_c_495_n 0.00532756f $X=0.75 $Y=2.495 $X2=0 $Y2=0
cc_294 N_VPWR_c_440_n N_X_c_495_n 0.0274543f $X=2.19 $Y=2.495 $X2=0 $Y2=0
cc_295 N_VPWR_c_441_n N_X_c_495_n 0.0274543f $X=3.63 $Y=2.495 $X2=0 $Y2=0
cc_296 N_X_c_489_n N_VGND_c_542_n 0.018528f $X=4.06 $Y=0.42 $X2=0 $Y2=0
cc_297 N_X_M1009_d N_VGND_c_543_n 0.00371702f $X=3.92 $Y=0.235 $X2=0 $Y2=0
cc_298 N_X_c_489_n N_VGND_c_543_n 0.0104192f $X=4.06 $Y=0.42 $X2=0 $Y2=0
