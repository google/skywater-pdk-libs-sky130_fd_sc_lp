* File: sky130_fd_sc_lp__o32ai_0.pex.spice
* Created: Fri Aug 28 11:18:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32AI_0%B1 1 3 4 6 8 9 10 11
c29 4 0 9.18442e-20 $X=0.59 $Y=1.61
c30 1 0 3.55387e-20 $X=0.505 $Y=0.94
r31 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.37
+ $Y=1.105 $X2=0.37 $Y2=1.105
r32 10 11 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=2.035
r33 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r34 9 18 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.105
r35 8 18 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.27 $Y=0.925
+ $X2=0.27 $Y2=1.105
r36 4 17 77.6914 $w=4.4e-07 $l=5.77321e-07 $layer=POLY_cond $X=0.59 $Y=1.61
+ $X2=0.435 $Y2=1.105
r37 4 6 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=0.59 $Y=1.61
+ $X2=0.59 $Y2=2.775
r38 1 17 40.446 $w=4.4e-07 $l=1.96914e-07 $layer=POLY_cond $X=0.505 $Y=0.94
+ $X2=0.435 $Y2=1.105
r39 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=0.94
+ $X2=0.505 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%B2 3 7 11 12 13 14 18
c44 7 0 1.83833e-19 $X=1.005 $Y=0.62
r45 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.07
+ $Y=1.725 $X2=1.07 $Y2=1.725
r46 14 19 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.17 $Y=2.035
+ $X2=1.17 $Y2=1.725
r47 13 19 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=1.17 $Y=1.665 $X2=1.17
+ $Y2=1.725
r48 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.07 $Y=2.065
+ $X2=1.07 $Y2=1.725
r49 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=2.065
+ $X2=1.07 $Y2=2.23
r50 10 18 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.56
+ $X2=1.07 $Y2=1.725
r51 7 10 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.005 $Y=0.62 $X2=1.005
+ $Y2=1.56
r52 3 12 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.98 $Y=2.775
+ $X2=0.98 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%A3 3 6 9 11 12 13 14 15 16 23
r45 23 26 5.70477 $w=4.45e-07 $l=1.5e-08 $layer=POLY_cond $X=1.582 $Y=1.375
+ $X2=1.582 $Y2=1.39
r46 23 25 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.582 $Y=1.375
+ $X2=1.582 $Y2=1.21
r47 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=2.405
+ $X2=1.695 $Y2=2.775
r48 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=2.035
+ $X2=1.695 $Y2=2.405
r49 13 14 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.035
r50 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=1.295
+ $X2=1.695 $Y2=1.665
r51 12 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.64
+ $Y=1.375 $X2=1.64 $Y2=1.375
r52 9 11 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=1.55 $Y=2.775
+ $X2=1.55 $Y2=1.88
r53 6 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.64 $Y=1.715
+ $X2=1.64 $Y2=1.88
r54 6 26 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=1.64 $Y=1.715
+ $X2=1.64 $Y2=1.39
r55 3 25 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.435 $Y=0.62
+ $X2=1.435 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%A2 3 7 11 12 13 14 15 16 17 24
r42 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=2.405
+ $X2=2.17 $Y2=2.775
r43 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=2.035
+ $X2=2.17 $Y2=2.405
r44 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=2.035
r45 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=1.295
+ $X2=2.17 $Y2=1.665
r46 13 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.21
+ $Y=1.375 $X2=2.21 $Y2=1.375
r47 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.21 $Y=1.715
+ $X2=2.21 $Y2=1.375
r48 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.715
+ $X2=2.21 $Y2=1.88
r49 10 24 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.21
+ $X2=2.21 $Y2=1.375
r50 7 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.26 $Y=0.62 $X2=2.26
+ $Y2=1.21
r51 3 12 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=2.12 $Y=2.775
+ $X2=2.12 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%A1 3 7 10 13 17 18 19 20 21 26
r37 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.78
+ $Y=1.375 $X2=2.78 $Y2=1.375
r38 20 21 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.73 $Y=1.665
+ $X2=2.73 $Y2=2.035
r39 20 27 7.70806 $w=4.48e-07 $l=2.9e-07 $layer=LI1_cond $X=2.73 $Y=1.665
+ $X2=2.73 $Y2=1.375
r40 19 27 2.12636 $w=4.48e-07 $l=8e-08 $layer=LI1_cond $X=2.73 $Y=1.295 $X2=2.73
+ $Y2=1.375
r41 17 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.78 $Y=1.715
+ $X2=2.78 $Y2=1.375
r42 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=1.715
+ $X2=2.78 $Y2=1.88
r43 16 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=1.21
+ $X2=2.78 $Y2=1.375
r44 11 13 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.51 $Y=2.195
+ $X2=2.69 $Y2=2.195
r45 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.69 $Y=2.12
+ $X2=2.69 $Y2=2.195
r46 10 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.69 $Y=2.12
+ $X2=2.69 $Y2=1.88
r47 7 16 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.69 $Y=0.62 $X2=2.69
+ $Y2=1.21
r48 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.51 $Y=2.27 $X2=2.51
+ $Y2=2.195
r49 1 3 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.51 $Y=2.27 $X2=2.51
+ $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%VPWR 1 2 7 9 13 15 17 24 25 31
r36 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 25 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 22 31 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.725 $Y2=3.33
r41 22 24 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 18 28 3.915 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r45 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 17 31 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.62 $Y=3.33
+ $X2=2.725 $Y2=3.33
r47 17 20 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=2.62 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 15 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 11 31 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=3.33
r51 11 13 33.5368 $w=2.08e-07 $l=6.35e-07 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=2.61
r52 7 28 3.22816 $w=2.5e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.227 $Y2=3.33
r53 7 9 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.33 $Y=3.245 $X2=0.33
+ $Y2=2.6
r54 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.585
+ $Y=2.455 $X2=2.725 $Y2=2.61
r55 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=2.455 $X2=0.37 $Y2=2.6
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%Y 1 2 7 8 9 10 11 12 23 36 38
r35 29 36 1.7512 $w=1.88e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=2.435 $X2=0.72
+ $Y2=2.405
r36 21 38 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=0.79 $Y=1.225 $X2=0.79
+ $Y2=1.295
r37 12 44 10.6457 $w=5.73e-07 $l=5e-07 $layer=LI1_cond $X=0.72 $Y=2.755 $X2=1.22
+ $Y2=2.755
r38 12 29 7.31424 $w=1.9e-07 $l=3.2e-07 $layer=LI1_cond $X=0.72 $Y=2.755
+ $X2=0.72 $Y2=2.435
r39 11 12 8.02089 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=0.72 $Y=2.462
+ $X2=0.72 $Y2=2.755
r40 11 36 1.63445 $w=1.88e-07 $l=2.8e-08 $layer=LI1_cond $X=0.72 $Y=2.377
+ $X2=0.72 $Y2=2.405
r41 10 11 19.9636 $w=1.88e-07 $l=3.42e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.377
r42 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=2.035
r43 9 40 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=1.39
r44 8 40 5.12995 $w=3.28e-07 $l=8.8e-08 $layer=LI1_cond $X=0.79 $Y=1.302
+ $X2=0.79 $Y2=1.39
r45 8 38 0.244458 $w=3.28e-07 $l=7e-09 $layer=LI1_cond $X=0.79 $Y=1.302 $X2=0.79
+ $Y2=1.295
r46 8 21 0.27938 $w=3.28e-07 $l=8e-09 $layer=LI1_cond $X=0.79 $Y=1.217 $X2=0.79
+ $Y2=1.225
r47 7 8 10.1974 $w=3.28e-07 $l=2.92e-07 $layer=LI1_cond $X=0.79 $Y=0.925
+ $X2=0.79 $Y2=1.217
r48 7 23 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.79 $Y=0.925
+ $X2=0.79 $Y2=0.705
r49 2 44 300 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=2.455 $X2=1.22 $Y2=2.6
r50 1 23 182 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.41 $X2=0.79 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%A_33_82# 1 2 3 10 15 16 17 20 22
c40 10 0 9.18442e-20 $X=1.125 $Y=0.34
r41 22 25 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.29 $Y=0.34
+ $X2=0.29 $Y2=0.565
r42 18 20 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=2.48 $Y=0.87
+ $X2=2.48 $Y2=0.62
r43 16 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.38 $Y=0.955
+ $X2=2.48 $Y2=0.87
r44 16 17 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=2.38 $Y=0.955
+ $X2=1.315 $Y2=0.955
r45 13 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.22 $Y=0.87
+ $X2=1.315 $Y2=0.955
r46 13 15 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.22 $Y=0.87
+ $X2=1.22 $Y2=0.62
r47 12 15 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.22 $Y2=0.62
r48 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=0.34
+ $X2=0.29 $Y2=0.34
r49 10 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.125 $Y=0.34
+ $X2=1.22 $Y2=0.425
r50 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.125 $Y=0.34
+ $X2=0.455 $Y2=0.34
r51 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.41 $X2=2.475 $Y2=0.62
r52 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.41 $X2=1.22 $Y2=0.62
r53 1 25 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.41 $X2=0.29 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LP__O32AI_0%VGND 1 2 9 11 12 13 14 16 30
c27 30 0 3.55387e-20 $X=3.12 $Y=0
c28 16 0 1.83833e-19 $X=1.485 $Y=0
r29 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r30 27 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r31 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r32 24 26 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.64
+ $Y2=0
r33 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r34 19 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r35 18 22 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r36 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 16 36 9.48614 $w=7.23e-07 $l=5.75e-07 $layer=LI1_cond $X=1.847 $Y=0
+ $X2=1.847 $Y2=0.575
r38 16 24 9.55322 $w=1.7e-07 $l=3.63e-07 $layer=LI1_cond $X=1.847 $Y=0 $X2=2.21
+ $Y2=0
r39 16 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.2
+ $Y2=0
r40 14 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r41 14 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r42 14 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r43 12 26 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r44 12 13 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.935
+ $Y2=0
r45 11 29 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.12
+ $Y2=0
r46 11 13 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=2.935
+ $Y2=0
r47 7 13 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=0.085
+ $X2=2.935 $Y2=0
r48 7 9 22.8354 $w=2.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.935 $Y=0.085
+ $X2=2.935 $Y2=0.62
r49 2 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.765
+ $Y=0.41 $X2=2.905 $Y2=0.62
r50 1 36 91 $w=1.7e-07 $l=6.11964e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.41 $X2=2.045 $Y2=0.575
.ends

