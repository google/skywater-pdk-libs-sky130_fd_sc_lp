* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21o_0 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_319_473# B1 a_80_275# VPB phighvt w=640000u l=150000u
+  ad=3.488e+11p pd=3.65e+06u as=1.696e+11p ps=1.81e+06u
M1001 a_319_473# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.488e+11p ps=3.65e+06u
M1002 a_80_275# B1 VGND VNB nshort w=420000u l=150000u
+  ad=1.449e+11p pd=1.53e+06u as=2.625e+11p ps=2.93e+06u
M1003 VPWR a_80_275# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1004 a_405_47# A1 a_80_275# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1005 VGND A2 a_405_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_319_473# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_80_275# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends
