* File: sky130_fd_sc_lp__invlp_1.pex.spice
* Created: Wed Sep  2 09:57:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVLP_1%A 1 3 6 8 10 12 15 17 18 19 20
r33 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.35 $X2=0.29 $Y2=1.35
r34 17 23 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.47 $Y=1.35 $X2=0.29
+ $Y2=1.35
r35 17 18 6.91837 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.47 $Y=1.35 $X2=0.56
+ $Y2=1.35
r36 13 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.935 $Y=1.335
+ $X2=0.935 $Y2=1.26
r37 13 15 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=0.935 $Y=1.335
+ $X2=0.935 $Y2=2.465
r38 10 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.935 $Y=1.185
+ $X2=0.935 $Y2=1.26
r39 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=1.185
+ $X2=0.935 $Y2=0.655
r40 9 18 6.91837 $w=1.5e-07 $l=1.27279e-07 $layer=POLY_cond $X=0.65 $Y=1.26
+ $X2=0.56 $Y2=1.35
r41 8 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.86 $Y=1.26
+ $X2=0.935 $Y2=1.26
r42 8 9 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.86 $Y=1.26 $X2=0.65
+ $Y2=1.26
r43 4 18 18.1359 $w=1.5e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.575 $Y=1.515
+ $X2=0.56 $Y2=1.35
r44 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.575 $Y=1.515
+ $X2=0.575 $Y2=2.465
r45 1 18 18.1359 $w=1.5e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.545 $Y=1.185
+ $X2=0.56 $Y2=1.35
r46 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.545 $Y=1.185
+ $X2=0.545 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_1%VPWR 1 4 6 10 14 15
r18 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r20 12 18 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.262 $Y2=3.33
r21 12 14 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=1.2 $Y2=3.33
r22 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r23 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 6 9 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=0.36 $Y=1.98 $X2=0.36
+ $Y2=2.95
r25 4 18 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.262 $Y2=3.33
r26 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.36 $Y2=2.95
r27 1 9 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.36 $Y2=2.95
r28 1 6 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.36 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_1%Y 1 2 7 8 9 10 11 12 13 22
r16 13 40 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.15 $Y=2.775
+ $X2=1.15 $Y2=2.91
r17 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=2.405
+ $X2=1.15 $Y2=2.775
r18 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.15 $Y=1.98
+ $X2=1.15 $Y2=2.405
r19 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.98
r20 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.665
r21 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.925 $X2=1.15
+ $Y2=1.295
r22 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.555 $X2=1.15
+ $Y2=0.925
r23 7 22 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.15 $Y=0.555
+ $X2=1.15 $Y2=0.42
r24 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=2.91
r25 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=1.98
r26 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_1%VGND 1 4 6 8 12 13
r17 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r18 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r19 10 16 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=0.247
+ $Y2=0
r20 10 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=1.2
+ $Y2=0
r21 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r22 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r23 4 16 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.247 $Y2=0
r24 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.33 $Y2=0.38
r25 1 6 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.185
+ $Y=0.235 $X2=0.33 $Y2=0.38
.ends

