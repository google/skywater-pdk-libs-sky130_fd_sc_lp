* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__clkbuflp_16 A VGND VNB VPB VPWR X
X0 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_1536_47# a_130_417# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X2 a_2010_47# a_130_417# X VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X3 a_130_417# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VGND a_130_417# a_1694_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X5 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_110_47# A a_130_417# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X8 VGND a_130_417# a_1062_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X9 VPWR A a_130_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X12 VPWR A a_130_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_426_47# A a_130_417# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X14 VGND a_130_417# a_1378_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X15 a_130_417# A a_584_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X16 X a_130_417# a_2168_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X17 X a_130_417# a_1220_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X18 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 VPWR A a_130_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_130_417# A a_268_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X23 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X24 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 VGND A a_426_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X27 a_904_47# a_130_417# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X28 a_130_417# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X29 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X30 a_1378_47# a_130_417# X VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X31 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 a_1694_47# a_130_417# X VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X33 a_2168_47# a_130_417# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X34 X a_130_417# a_1852_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X35 VGND a_130_417# a_746_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X36 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X37 a_1062_47# a_130_417# X VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X38 VPWR a_130_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X39 a_268_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X40 a_1852_47# a_130_417# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X41 a_746_47# a_130_417# X VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X42 VGND a_130_417# a_2010_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X43 a_130_417# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X44 a_584_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X45 X a_130_417# a_904_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X46 X a_130_417# a_1536_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X47 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X48 X a_130_417# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X49 a_1220_47# a_130_417# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
.ends
