* File: sky130_fd_sc_lp__dlxbp_lp.pxi.spice
* Created: Fri Aug 28 10:28:23 2020
* 
x_PM_SKY130_FD_SC_LP__DLXBP_LP%D N_D_c_187_n N_D_M1032_g N_D_M1021_g N_D_M1028_g
+ N_D_M1010_g N_D_c_185_n D D D N_D_c_186_n PM_SKY130_FD_SC_LP__DLXBP_LP%D
x_PM_SKY130_FD_SC_LP__DLXBP_LP%GATE N_GATE_M1011_g N_GATE_M1025_g N_GATE_M1033_g
+ N_GATE_M1023_g GATE GATE N_GATE_c_227_n PM_SKY130_FD_SC_LP__DLXBP_LP%GATE
x_PM_SKY130_FD_SC_LP__DLXBP_LP%A_350_111# N_A_350_111#_M1033_d
+ N_A_350_111#_M1023_d N_A_350_111#_M1007_g N_A_350_111#_M1012_g
+ N_A_350_111#_M1008_g N_A_350_111#_M1015_g N_A_350_111#_M1017_g
+ N_A_350_111#_M1020_g N_A_350_111#_c_297_n N_A_350_111#_c_298_n
+ N_A_350_111#_c_283_n N_A_350_111#_c_284_n N_A_350_111#_c_285_n
+ N_A_350_111#_c_286_n N_A_350_111#_c_302_n N_A_350_111#_c_287_n
+ N_A_350_111#_c_288_n N_A_350_111#_c_289_n N_A_350_111#_c_290_n
+ N_A_350_111#_c_291_n N_A_350_111#_c_292_n N_A_350_111#_c_293_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP%A_350_111#
x_PM_SKY130_FD_SC_LP__DLXBP_LP%A_27_111# N_A_27_111#_M1021_s N_A_27_111#_M1032_s
+ N_A_27_111#_M1009_g N_A_27_111#_M1013_g N_A_27_111#_c_434_n
+ N_A_27_111#_c_435_n N_A_27_111#_c_440_n N_A_27_111#_c_441_n
+ N_A_27_111#_c_442_n N_A_27_111#_c_443_n N_A_27_111#_c_444_n
+ N_A_27_111#_c_445_n N_A_27_111#_c_436_n N_A_27_111#_c_446_n
+ N_A_27_111#_c_447_n N_A_27_111#_c_448_n N_A_27_111#_c_437_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP%A_27_111#
x_PM_SKY130_FD_SC_LP__DLXBP_LP%A_469_47# N_A_469_47#_M1007_s N_A_469_47#_M1012_s
+ N_A_469_47#_M1019_g N_A_469_47#_c_540_n N_A_469_47#_c_541_n
+ N_A_469_47#_M1029_g N_A_469_47#_c_543_n N_A_469_47#_c_544_n
+ N_A_469_47#_c_545_n N_A_469_47#_c_546_n N_A_469_47#_c_547_n
+ N_A_469_47#_c_556_n N_A_469_47#_c_557_n N_A_469_47#_c_548_n
+ N_A_469_47#_c_558_n N_A_469_47#_c_549_n N_A_469_47#_c_550_n
+ N_A_469_47#_c_551_n N_A_469_47#_c_552_n N_A_469_47#_c_553_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP%A_469_47#
x_PM_SKY130_FD_SC_LP__DLXBP_LP%A_969_407# N_A_969_407#_M1022_d
+ N_A_969_407#_M1014_d N_A_969_407#_M1005_g N_A_969_407#_M1001_g
+ N_A_969_407#_M1034_g N_A_969_407#_M1018_g N_A_969_407#_M1002_g
+ N_A_969_407#_M1016_g N_A_969_407#_M1035_g N_A_969_407#_M1000_g
+ N_A_969_407#_c_679_n N_A_969_407#_c_680_n N_A_969_407#_M1024_g
+ N_A_969_407#_M1003_g N_A_969_407#_c_683_n N_A_969_407#_c_696_n
+ N_A_969_407#_c_697_n N_A_969_407#_c_684_n N_A_969_407#_c_698_n
+ N_A_969_407#_c_685_n N_A_969_407#_c_686_n N_A_969_407#_c_687_n
+ N_A_969_407#_c_699_n N_A_969_407#_c_688_n N_A_969_407#_c_689_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP%A_969_407#
x_PM_SKY130_FD_SC_LP__DLXBP_LP%A_798_47# N_A_798_47#_M1019_d N_A_798_47#_M1017_d
+ N_A_798_47#_M1031_g N_A_798_47#_M1026_g N_A_798_47#_M1022_g
+ N_A_798_47#_M1014_g N_A_798_47#_c_842_n N_A_798_47#_c_837_n
+ N_A_798_47#_c_838_n N_A_798_47#_c_839_n N_A_798_47#_c_831_n
+ N_A_798_47#_c_832_n N_A_798_47#_c_833_n N_A_798_47#_c_841_n
+ N_A_798_47#_c_834_n PM_SKY130_FD_SC_LP__DLXBP_LP%A_798_47#
x_PM_SKY130_FD_SC_LP__DLXBP_LP%A_1662_131# N_A_1662_131#_M1024_d
+ N_A_1662_131#_M1003_d N_A_1662_131#_M1027_g N_A_1662_131#_M1004_g
+ N_A_1662_131#_M1030_g N_A_1662_131#_M1006_g N_A_1662_131#_c_937_n
+ N_A_1662_131#_c_943_n N_A_1662_131#_c_938_n N_A_1662_131#_c_939_n
+ N_A_1662_131#_c_940_n PM_SKY130_FD_SC_LP__DLXBP_LP%A_1662_131#
x_PM_SKY130_FD_SC_LP__DLXBP_LP%VPWR N_VPWR_M1028_d N_VPWR_M1015_d N_VPWR_M1005_d
+ N_VPWR_M1016_d N_VPWR_M1004_s N_VPWR_c_987_n N_VPWR_c_988_n N_VPWR_c_989_n
+ N_VPWR_c_990_n N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_993_n VPWR
+ N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_996_n N_VPWR_c_997_n N_VPWR_c_998_n
+ N_VPWR_c_986_n N_VPWR_c_1000_n N_VPWR_c_1001_n N_VPWR_c_1002_n N_VPWR_c_1003_n
+ PM_SKY130_FD_SC_LP__DLXBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DLXBP_LP%Q N_Q_M1034_s N_Q_M1018_s N_Q_c_1096_n
+ N_Q_c_1100_n N_Q_c_1101_n N_Q_c_1097_n N_Q_c_1098_n N_Q_c_1102_n Q Q
+ PM_SKY130_FD_SC_LP__DLXBP_LP%Q
x_PM_SKY130_FD_SC_LP__DLXBP_LP%Q_N N_Q_N_M1030_d N_Q_N_M1006_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1164_n PM_SKY130_FD_SC_LP__DLXBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__DLXBP_LP%VGND N_VGND_M1010_d N_VGND_M1008_d N_VGND_M1001_d
+ N_VGND_M1002_d N_VGND_M1027_s N_VGND_c_1179_n N_VGND_c_1180_n N_VGND_c_1181_n
+ N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n N_VGND_c_1185_n
+ N_VGND_c_1186_n N_VGND_c_1187_n VGND N_VGND_c_1188_n N_VGND_c_1189_n
+ N_VGND_c_1190_n N_VGND_c_1191_n N_VGND_c_1192_n N_VGND_c_1193_n
+ N_VGND_c_1194_n N_VGND_c_1195_n PM_SKY130_FD_SC_LP__DLXBP_LP%VGND
cc_1 VNB N_D_M1021_g 0.0237545f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.765
cc_2 VNB N_D_M1010_g 0.0177614f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.765
cc_3 VNB N_D_c_185_n 0.0170167f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.285
cc_4 VNB N_D_c_186_n 0.0357503f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.345
cc_5 VNB N_GATE_M1011_g 0.0387582f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.725
cc_6 VNB N_GATE_M1033_g 0.0324124f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.725
cc_7 VNB GATE 0.00412791f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.7
cc_8 VNB N_GATE_c_227_n 0.00922234f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.285
cc_9 VNB N_A_350_111#_M1007_g 0.0436884f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.85
cc_10 VNB N_A_350_111#_M1008_g 0.0349027f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.85
cc_11 VNB N_A_350_111#_M1020_g 0.0219496f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.345
cc_12 VNB N_A_350_111#_c_283_n 0.00906246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_350_111#_c_284_n 0.00241836f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=2.035
cc_14 VNB N_A_350_111#_c_285_n 0.012606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_350_111#_c_286_n 0.00175436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_350_111#_c_287_n 0.00360728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_350_111#_c_288_n 0.0108757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_350_111#_c_289_n 5.74387e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_350_111#_c_290_n 0.0509677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_350_111#_c_291_n 0.00809093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_350_111#_c_292_n 0.0033547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_350_111#_c_293_n 0.0321452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_111#_M1009_g 0.0474966f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.725
cc_24 VNB N_A_27_111#_c_434_n 0.00896356f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.7
cc_25 VNB N_A_27_111#_c_435_n 0.031488f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.285
cc_26 VNB N_A_27_111#_c_436_n 0.0270979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_111#_c_437_n 0.00170034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_469_47#_M1019_g 0.0203318f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.85
cc_29 VNB N_A_469_47#_c_540_n 0.0316409f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.725
cc_30 VNB N_A_469_47#_c_541_n 0.0171819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_469_47#_M1029_g 0.0044862f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.765
cc_32 VNB N_A_469_47#_c_543_n 0.0292652f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.85
cc_33 VNB N_A_469_47#_c_544_n 0.00607939f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.135
cc_34 VNB N_A_469_47#_c_545_n 0.0214559f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.285
cc_35 VNB N_A_469_47#_c_546_n 0.00325508f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_36 VNB N_A_469_47#_c_547_n 2.85047e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_37 VNB N_A_469_47#_c_548_n 0.00533739f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.345
cc_38 VNB N_A_469_47#_c_549_n 0.0180449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_469_47#_c_550_n 0.00691027f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.035
cc_40 VNB N_A_469_47#_c_551_n 0.00904847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_469_47#_c_552_n 0.00239131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_469_47#_c_553_n 0.0152664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_969_407#_M1001_g 0.0665153f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.135
cc_44 VNB N_A_969_407#_M1034_g 0.0245555f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.7
cc_45 VNB N_A_969_407#_M1018_g 0.00111882f $X=-0.19 $Y=-0.245 $X2=0.675
+ $Y2=1.135
cc_46 VNB N_A_969_407#_M1002_g 0.0221698f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_47 VNB N_A_969_407#_M1016_g 9.81478e-19 $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.345
cc_48 VNB N_A_969_407#_M1035_g 0.0213167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_969_407#_M1000_g 8.18727e-19 $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=2.035
cc_50 VNB N_A_969_407#_c_679_n 0.00708691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_969_407#_c_680_n 0.08164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_969_407#_M1024_g 0.0263374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_969_407#_M1003_g 0.00994614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_969_407#_c_683_n 0.00822478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_969_407#_c_684_n 0.00598271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_969_407#_c_685_n 0.00402752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_969_407#_c_686_n 0.0125578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_969_407#_c_687_n 0.00308103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_969_407#_c_688_n 5.29676e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_969_407#_c_689_n 0.00496069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_798_47#_M1031_g 0.0218546f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.85
cc_62 VNB N_A_798_47#_M1026_g 0.00111192f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.135
cc_63 VNB N_A_798_47#_M1022_g 0.0234011f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.7
cc_64 VNB N_A_798_47#_M1014_g 9.79778e-19 $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.135
cc_65 VNB N_A_798_47#_c_831_n 0.00536675f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.295
cc_66 VNB N_A_798_47#_c_832_n 0.00344911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_798_47#_c_833_n 0.0179062f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.665
cc_68 VNB N_A_798_47#_c_834_n 0.0587162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1662_131#_M1027_g 0.0238669f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.85
cc_70 VNB N_A_1662_131#_M1004_g 0.00111761f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=1.135
cc_71 VNB N_A_1662_131#_M1030_g 0.0249073f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.7
cc_72 VNB N_A_1662_131#_M1006_g 0.00112085f $X=-0.19 $Y=-0.245 $X2=0.675
+ $Y2=1.135
cc_73 VNB N_A_1662_131#_c_937_n 0.011791f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_74 VNB N_A_1662_131#_c_938_n 0.0181925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1662_131#_c_939_n 0.00290493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1662_131#_c_940_n 0.043279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VPWR_c_986_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_Q_c_1096_n 0.00597105f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.85
cc_79 VNB N_Q_c_1097_n 0.00747991f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.765
cc_80 VNB N_Q_c_1098_n 0.00369896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB Q 0.00279274f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_82 VNB N_Q_N_c_1164_n 0.0576172f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.285
cc_83 VNB N_VGND_c_1179_n 0.0231364f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.7
cc_84 VNB N_VGND_c_1180_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.285
cc_85 VNB N_VGND_c_1181_n 0.00886409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1182_n 0.0149886f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.295
cc_87 VNB N_VGND_c_1183_n 0.0230144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1184_n 0.0291076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1185_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1186_n 0.0504205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1187_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1188_n 0.0455449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1189_n 0.0493886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1190_n 0.0355488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1191_n 0.0269285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1192_n 0.551196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1193_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1194_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1195_n 0.00536178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VPB N_D_c_187_n 0.0157651f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.85
cc_101 VPB N_D_M1032_g 0.0433399f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.725
cc_102 VPB N_D_M1028_g 0.0356151f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.725
cc_103 VPB D 0.00428882f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_104 VPB N_D_c_186_n 0.00416726f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.345
cc_105 VPB N_GATE_M1025_g 0.0212902f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.765
cc_106 VPB N_GATE_M1033_g 0.00790719f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.725
cc_107 VPB N_GATE_M1023_g 0.0257911f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.765
cc_108 VPB GATE 0.00504023f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.7
cc_109 VPB N_GATE_c_227_n 0.0723457f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.285
cc_110 VPB N_A_350_111#_M1012_g 0.0210934f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.765
cc_111 VPB N_A_350_111#_M1015_g 0.034792f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_112 VPB N_A_350_111#_M1017_g 0.0234023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_350_111#_c_297_n 0.0179059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_350_111#_c_298_n 0.0127397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_350_111#_c_283_n 0.00758424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_350_111#_c_284_n 0.0156273f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.035
cc_117 VPB N_A_350_111#_c_286_n 0.00654862f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_350_111#_c_302_n 0.0322916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_350_111#_c_289_n 0.00174513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_350_111#_c_290_n 0.0257515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_27_111#_M1013_g 0.0209805f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.765
cc_122 VPB N_A_27_111#_c_435_n 0.0348535f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.285
cc_123 VPB N_A_27_111#_c_440_n 0.0157024f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_124 VPB N_A_27_111#_c_441_n 0.0190339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_27_111#_c_442_n 0.00135432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_27_111#_c_443_n 0.00107343f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.345
cc_127 VPB N_A_27_111#_c_444_n 0.00646684f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.345
cc_128 VPB N_A_27_111#_c_445_n 0.0027073f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.295
cc_129 VPB N_A_27_111#_c_446_n 0.0345117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_27_111#_c_447_n 0.00459228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_27_111#_c_448_n 0.0311368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_27_111#_c_437_n 0.0139161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_469_47#_M1029_g 0.0594831f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.765
cc_134 VPB N_A_469_47#_c_547_n 0.00161798f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_135 VPB N_A_469_47#_c_556_n 0.0223985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_469_47#_c_557_n 0.00113268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_469_47#_c_558_n 0.00896572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_969_407#_M1005_g 0.0266605f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.85
cc_139 VPB N_A_969_407#_M1001_g 0.0241762f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.135
cc_140 VPB N_A_969_407#_M1018_g 0.023664f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.135
cc_141 VPB N_A_969_407#_M1016_g 0.0211901f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.345
cc_142 VPB N_A_969_407#_M1000_g 0.0198965f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.035
cc_143 VPB N_A_969_407#_M1003_g 0.0236929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_969_407#_c_696_n 0.00956945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_969_407#_c_697_n 0.0352588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_969_407#_c_698_n 0.0080435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_969_407#_c_699_n 0.0057577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_969_407#_c_688_n 0.00443255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_798_47#_M1026_g 0.0221262f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.135
cc_150 VPB N_A_798_47#_M1014_g 0.0225996f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.135
cc_151 VPB N_A_798_47#_c_837_n 0.00650625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_798_47#_c_838_n 0.0143279f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.345
cc_153 VPB N_A_798_47#_c_839_n 0.00171732f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.345
cc_154 VPB N_A_798_47#_c_832_n 0.0011066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_798_47#_c_841_n 0.0055191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_1662_131#_M1004_g 0.0225948f $X=-0.19 $Y=1.655 $X2=0.855
+ $Y2=1.135
cc_157 VPB N_A_1662_131#_M1006_g 0.023487f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.135
cc_158 VPB N_A_1662_131#_c_943_n 0.0155409f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.345
cc_159 VPB N_A_1662_131#_c_938_n 0.00560262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_987_n 0.00414835f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.7
cc_161 VPB N_VPWR_c_988_n 0.0068952f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.285
cc_162 VPB N_VPWR_c_989_n 0.00524698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_990_n 0.0244399f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.345
cc_164 VPB N_VPWR_c_991_n 0.0328362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_992_n 0.0490247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_993_n 0.005715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_994_n 0.0268803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_995_n 0.0503192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_996_n 0.0491471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_997_n 0.0350997f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_998_n 0.0262537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_986_n 0.157883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1000_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1001_n 0.00533588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1002_n 0.00533588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1003_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_Q_c_1100_n 0.00351621f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.725
cc_178 VPB N_Q_c_1101_n 0.011688f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.135
cc_179 VPB N_Q_c_1102_n 0.00657061f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.7
cc_180 VPB Q 0.00293393f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_181 VPB N_Q_N_c_1164_n 0.0554597f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.285
cc_182 N_D_M1010_g N_GATE_M1011_g 0.0205062f $X=0.855 $Y=0.765 $X2=0 $Y2=0
cc_183 D N_GATE_M1011_g 0.0012782f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_184 N_D_c_186_n N_GATE_M1011_g 0.0104124f $X=0.735 $Y=1.345 $X2=0 $Y2=0
cc_185 N_D_M1028_g N_GATE_M1025_g 0.0259566f $X=0.845 $Y=2.725 $X2=0 $Y2=0
cc_186 D GATE 0.0460589f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_187 N_D_c_186_n GATE 0.00461396f $X=0.735 $Y=1.345 $X2=0 $Y2=0
cc_188 D N_GATE_c_227_n 6.87204e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_189 N_D_c_186_n N_GATE_c_227_n 0.0414187f $X=0.735 $Y=1.345 $X2=0 $Y2=0
cc_190 N_D_c_187_n N_A_27_111#_c_435_n 0.0170475f $X=0.485 $Y=1.85 $X2=0 $Y2=0
cc_191 N_D_M1021_g N_A_27_111#_c_435_n 0.0188016f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_192 D N_A_27_111#_c_435_n 0.0494982f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_193 N_D_M1032_g N_A_27_111#_c_440_n 0.0116926f $X=0.485 $Y=2.725 $X2=0 $Y2=0
cc_194 N_D_M1028_g N_A_27_111#_c_440_n 0.0121358f $X=0.845 $Y=2.725 $X2=0 $Y2=0
cc_195 D N_A_27_111#_c_440_n 0.0209676f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_196 N_D_M1021_g N_A_27_111#_c_436_n 0.0102874f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_197 N_D_M1010_g N_A_27_111#_c_436_n 0.00125175f $X=0.855 $Y=0.765 $X2=0 $Y2=0
cc_198 N_D_M1032_g N_A_27_111#_c_446_n 0.0109377f $X=0.485 $Y=2.725 $X2=0 $Y2=0
cc_199 N_D_M1028_g N_A_27_111#_c_446_n 0.00179788f $X=0.845 $Y=2.725 $X2=0 $Y2=0
cc_200 D N_A_469_47#_c_547_n 0.00470264f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_201 D N_A_469_47#_c_551_n 0.00604029f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_202 N_D_M1032_g N_VPWR_c_987_n 0.00175817f $X=0.485 $Y=2.725 $X2=0 $Y2=0
cc_203 N_D_M1028_g N_VPWR_c_987_n 0.00976681f $X=0.845 $Y=2.725 $X2=0 $Y2=0
cc_204 N_D_M1032_g N_VPWR_c_994_n 0.00502664f $X=0.485 $Y=2.725 $X2=0 $Y2=0
cc_205 N_D_M1028_g N_VPWR_c_994_n 0.00445056f $X=0.845 $Y=2.725 $X2=0 $Y2=0
cc_206 N_D_M1032_g N_VPWR_c_986_n 0.0061677f $X=0.485 $Y=2.725 $X2=0 $Y2=0
cc_207 N_D_M1028_g N_VPWR_c_986_n 0.00409056f $X=0.845 $Y=2.725 $X2=0 $Y2=0
cc_208 N_D_M1021_g N_VGND_c_1179_n 0.00180891f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_209 N_D_M1010_g N_VGND_c_1179_n 0.0125561f $X=0.855 $Y=0.765 $X2=0 $Y2=0
cc_210 N_D_M1021_g N_VGND_c_1184_n 0.00436277f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_211 N_D_M1010_g N_VGND_c_1184_n 0.00377474f $X=0.855 $Y=0.765 $X2=0 $Y2=0
cc_212 N_D_M1021_g N_VGND_c_1192_n 0.00489211f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_213 N_D_M1010_g N_VGND_c_1192_n 0.00410937f $X=0.855 $Y=0.765 $X2=0 $Y2=0
cc_214 N_GATE_M1033_g N_A_350_111#_c_283_n 0.0105701f $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_215 N_GATE_c_227_n N_A_350_111#_c_283_n 0.00876599f $X=1.295 $Y=1.69 $X2=0
+ $Y2=0
cc_216 N_GATE_M1033_g N_A_350_111#_c_288_n 0.00563149f $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_217 N_GATE_M1025_g N_A_27_111#_c_440_n 0.0110825f $X=1.315 $Y=2.725 $X2=0
+ $Y2=0
cc_218 N_GATE_M1023_g N_A_27_111#_c_440_n 0.00112908f $X=1.675 $Y=2.725 $X2=0
+ $Y2=0
cc_219 GATE N_A_27_111#_c_440_n 0.0218641f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_220 N_GATE_c_227_n N_A_27_111#_c_440_n 0.0021478f $X=1.295 $Y=1.69 $X2=0
+ $Y2=0
cc_221 N_GATE_M1023_g N_A_27_111#_c_441_n 0.01536f $X=1.675 $Y=2.725 $X2=0 $Y2=0
cc_222 N_GATE_M1025_g N_A_27_111#_c_442_n 6.87459e-19 $X=1.315 $Y=2.725 $X2=0
+ $Y2=0
cc_223 N_GATE_M1011_g N_A_469_47#_c_544_n 0.00717607f $X=1.285 $Y=0.765 $X2=0
+ $Y2=0
cc_224 N_GATE_M1033_g N_A_469_47#_c_544_n 0.00609524f $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_225 N_GATE_M1033_g N_A_469_47#_c_545_n 0.00896008f $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_226 N_GATE_M1011_g N_A_469_47#_c_547_n 0.00167311f $X=1.285 $Y=0.765 $X2=0
+ $Y2=0
cc_227 N_GATE_M1033_g N_A_469_47#_c_547_n 0.00425908f $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_228 GATE N_A_469_47#_c_547_n 0.0345371f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_229 N_GATE_c_227_n N_A_469_47#_c_547_n 0.0233379f $X=1.295 $Y=1.69 $X2=0
+ $Y2=0
cc_230 N_GATE_M1023_g N_A_469_47#_c_556_n 5.90786e-19 $X=1.675 $Y=2.725 $X2=0
+ $Y2=0
cc_231 N_GATE_c_227_n N_A_469_47#_c_556_n 0.00451351f $X=1.295 $Y=1.69 $X2=0
+ $Y2=0
cc_232 N_GATE_M1025_g N_A_469_47#_c_557_n 2.62073e-19 $X=1.315 $Y=2.725 $X2=0
+ $Y2=0
cc_233 N_GATE_M1023_g N_A_469_47#_c_557_n 0.00740612f $X=1.675 $Y=2.725 $X2=0
+ $Y2=0
cc_234 GATE N_A_469_47#_c_557_n 0.0121273f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_235 N_GATE_c_227_n N_A_469_47#_c_557_n 0.00488426f $X=1.295 $Y=1.69 $X2=0
+ $Y2=0
cc_236 N_GATE_M1033_g N_A_469_47#_c_548_n 0.00386865f $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_237 N_GATE_M1023_g N_A_469_47#_c_558_n 0.0117409f $X=1.675 $Y=2.725 $X2=0
+ $Y2=0
cc_238 N_GATE_M1033_g N_A_469_47#_c_550_n 4.07955e-19 $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_239 N_GATE_M1011_g N_A_469_47#_c_551_n 0.00220797f $X=1.285 $Y=0.765 $X2=0
+ $Y2=0
cc_240 N_GATE_M1033_g N_A_469_47#_c_551_n 0.0106728f $X=1.675 $Y=0.765 $X2=0
+ $Y2=0
cc_241 GATE N_A_469_47#_c_551_n 0.00107018f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_242 N_GATE_c_227_n N_A_469_47#_c_551_n 0.00245195f $X=1.295 $Y=1.69 $X2=0
+ $Y2=0
cc_243 N_GATE_M1025_g N_VPWR_c_987_n 0.00291478f $X=1.315 $Y=2.725 $X2=0 $Y2=0
cc_244 N_GATE_M1025_g N_VPWR_c_992_n 0.0053602f $X=1.315 $Y=2.725 $X2=0 $Y2=0
cc_245 N_GATE_M1023_g N_VPWR_c_992_n 0.00327726f $X=1.675 $Y=2.725 $X2=0 $Y2=0
cc_246 N_GATE_M1025_g N_VPWR_c_986_n 0.00553542f $X=1.315 $Y=2.725 $X2=0 $Y2=0
cc_247 N_GATE_M1023_g N_VPWR_c_986_n 0.00563495f $X=1.675 $Y=2.725 $X2=0 $Y2=0
cc_248 N_GATE_M1011_g N_VGND_c_1179_n 0.00132515f $X=1.285 $Y=0.765 $X2=0 $Y2=0
cc_249 GATE N_VGND_c_1179_n 0.00276806f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_250 N_GATE_M1011_g N_VGND_c_1186_n 0.00454183f $X=1.285 $Y=0.765 $X2=0 $Y2=0
cc_251 N_GATE_M1033_g N_VGND_c_1186_n 6.31558e-19 $X=1.675 $Y=0.765 $X2=0 $Y2=0
cc_252 N_GATE_M1011_g N_VGND_c_1192_n 0.00489211f $X=1.285 $Y=0.765 $X2=0 $Y2=0
cc_253 N_A_350_111#_M1008_g N_A_27_111#_M1009_g 0.0321666f $X=3.095 $Y=0.445
+ $X2=0 $Y2=0
cc_254 N_A_350_111#_c_285_n N_A_27_111#_M1009_g 0.00665079f $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_255 N_A_350_111#_c_289_n N_A_27_111#_M1009_g 6.85288e-19 $X=2.795 $Y=1.34
+ $X2=0 $Y2=0
cc_256 N_A_350_111#_c_290_n N_A_27_111#_M1009_g 0.01477f $X=2.795 $Y=1.34 $X2=0
+ $Y2=0
cc_257 N_A_350_111#_M1015_g N_A_27_111#_M1013_g 0.0221576f $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_258 N_A_350_111#_M1017_g N_A_27_111#_M1013_g 0.0497071f $X=4.02 $Y=2.695
+ $X2=0 $Y2=0
cc_259 N_A_350_111#_c_285_n N_A_27_111#_c_434_n 0.00601428f $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_260 N_A_350_111#_c_286_n N_A_27_111#_c_434_n 0.00176915f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_261 N_A_350_111#_c_289_n N_A_27_111#_c_434_n 0.00140525f $X=2.795 $Y=1.34
+ $X2=0 $Y2=0
cc_262 N_A_350_111#_c_290_n N_A_27_111#_c_434_n 0.0134571f $X=2.795 $Y=1.34
+ $X2=0 $Y2=0
cc_263 N_A_350_111#_M1023_d N_A_27_111#_c_441_n 0.0144377f $X=1.75 $Y=2.405
+ $X2=0 $Y2=0
cc_264 N_A_350_111#_M1012_g N_A_27_111#_c_441_n 0.0149289f $X=2.76 $Y=2.695
+ $X2=0 $Y2=0
cc_265 N_A_350_111#_M1015_g N_A_27_111#_c_441_n 0.00353004f $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_266 N_A_350_111#_M1015_g N_A_27_111#_c_443_n 0.0125956f $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_267 N_A_350_111#_c_298_n N_A_27_111#_c_443_n 0.00727823f $X=2.732 $Y=2.235
+ $X2=0 $Y2=0
cc_268 N_A_350_111#_M1015_g N_A_27_111#_c_444_n 0.0120876f $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_269 N_A_350_111#_c_285_n N_A_27_111#_c_444_n 0.0106748f $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_270 N_A_350_111#_M1015_g N_A_27_111#_c_445_n 0.00209871f $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_271 N_A_350_111#_c_297_n N_A_27_111#_c_445_n 6.16478e-19 $X=2.732 $Y=2.085
+ $X2=0 $Y2=0
cc_272 N_A_350_111#_c_298_n N_A_27_111#_c_445_n 7.99861e-19 $X=2.732 $Y=2.235
+ $X2=0 $Y2=0
cc_273 N_A_350_111#_c_285_n N_A_27_111#_c_445_n 0.00374137f $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_274 N_A_350_111#_c_289_n N_A_27_111#_c_445_n 0.00503112f $X=2.795 $Y=1.34
+ $X2=0 $Y2=0
cc_275 N_A_350_111#_c_290_n N_A_27_111#_c_445_n 4.273e-19 $X=2.795 $Y=1.34 $X2=0
+ $Y2=0
cc_276 N_A_350_111#_M1015_g N_A_27_111#_c_447_n 0.00118187f $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_277 N_A_350_111#_c_285_n N_A_27_111#_c_447_n 0.013429f $X=3.945 $Y=1.42 $X2=0
+ $Y2=0
cc_278 N_A_350_111#_c_286_n N_A_27_111#_c_447_n 0.019012f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_279 N_A_350_111#_c_302_n N_A_27_111#_c_447_n 0.0012425f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_280 N_A_350_111#_M1015_g N_A_27_111#_c_448_n 0.021263f $X=3.12 $Y=2.695 $X2=0
+ $Y2=0
cc_281 N_A_350_111#_c_285_n N_A_27_111#_c_448_n 9.14242e-19 $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_282 N_A_350_111#_c_286_n N_A_27_111#_c_448_n 0.00104487f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_283 N_A_350_111#_c_302_n N_A_27_111#_c_448_n 0.0201811f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_284 N_A_350_111#_M1015_g N_A_27_111#_c_437_n 0.0134571f $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_285 N_A_350_111#_c_286_n N_A_27_111#_c_437_n 0.00732121f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_286 N_A_350_111#_c_302_n N_A_27_111#_c_437_n 0.00104487f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_287 N_A_350_111#_M1020_g N_A_469_47#_M1019_g 0.0179416f $X=4.425 $Y=0.445
+ $X2=0 $Y2=0
cc_288 N_A_350_111#_c_286_n N_A_469_47#_c_540_n 0.00336357f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_289 N_A_350_111#_c_287_n N_A_469_47#_c_540_n 2.76972e-19 $X=4.435 $Y=1.335
+ $X2=0 $Y2=0
cc_290 N_A_350_111#_c_291_n N_A_469_47#_c_540_n 0.0167209f $X=4.435 $Y=1.42
+ $X2=0 $Y2=0
cc_291 N_A_350_111#_c_292_n N_A_469_47#_c_540_n 5.6519e-19 $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_292 N_A_350_111#_c_293_n N_A_469_47#_c_540_n 0.0158543f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_293 N_A_350_111#_c_285_n N_A_469_47#_c_541_n 0.00733301f $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_294 N_A_350_111#_c_286_n N_A_469_47#_c_541_n 0.00434066f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_295 N_A_350_111#_c_302_n N_A_469_47#_c_541_n 0.0143658f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_296 N_A_350_111#_c_291_n N_A_469_47#_c_541_n 0.00257938f $X=4.435 $Y=1.42
+ $X2=0 $Y2=0
cc_297 N_A_350_111#_M1017_g N_A_469_47#_M1029_g 0.0214972f $X=4.02 $Y=2.695
+ $X2=0 $Y2=0
cc_298 N_A_350_111#_c_286_n N_A_469_47#_M1029_g 0.0046447f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_299 N_A_350_111#_c_302_n N_A_469_47#_M1029_g 0.0205692f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_300 N_A_350_111#_c_285_n N_A_469_47#_c_543_n 0.00312728f $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_301 N_A_350_111#_c_287_n N_A_469_47#_c_543_n 0.00646024f $X=4.435 $Y=1.335
+ $X2=0 $Y2=0
cc_302 N_A_350_111#_c_291_n N_A_469_47#_c_543_n 0.00502426f $X=4.435 $Y=1.42
+ $X2=0 $Y2=0
cc_303 N_A_350_111#_c_283_n N_A_469_47#_c_544_n 0.00779174f $X=2.005 $Y=1.525
+ $X2=0 $Y2=0
cc_304 N_A_350_111#_c_288_n N_A_469_47#_c_544_n 0.014518f $X=1.89 $Y=0.765 $X2=0
+ $Y2=0
cc_305 N_A_350_111#_M1007_g N_A_469_47#_c_545_n 0.0032944f $X=2.705 $Y=0.445
+ $X2=0 $Y2=0
cc_306 N_A_350_111#_M1008_g N_A_469_47#_c_545_n 4.79243e-19 $X=3.095 $Y=0.445
+ $X2=0 $Y2=0
cc_307 N_A_350_111#_c_288_n N_A_469_47#_c_545_n 0.0241877f $X=1.89 $Y=0.765
+ $X2=0 $Y2=0
cc_308 N_A_350_111#_c_283_n N_A_469_47#_c_547_n 0.03725f $X=2.005 $Y=1.525 $X2=0
+ $Y2=0
cc_309 N_A_350_111#_M1023_d N_A_469_47#_c_556_n 0.0173211f $X=1.75 $Y=2.405
+ $X2=0 $Y2=0
cc_310 N_A_350_111#_c_297_n N_A_469_47#_c_556_n 0.00307805f $X=2.732 $Y=2.085
+ $X2=0 $Y2=0
cc_311 N_A_350_111#_c_298_n N_A_469_47#_c_556_n 0.004794f $X=2.732 $Y=2.235
+ $X2=0 $Y2=0
cc_312 N_A_350_111#_c_283_n N_A_469_47#_c_556_n 0.0192258f $X=2.005 $Y=1.525
+ $X2=0 $Y2=0
cc_313 N_A_350_111#_c_284_n N_A_469_47#_c_556_n 0.0356832f $X=2.63 $Y=1.685
+ $X2=0 $Y2=0
cc_314 N_A_350_111#_c_289_n N_A_469_47#_c_556_n 0.00610407f $X=2.795 $Y=1.34
+ $X2=0 $Y2=0
cc_315 N_A_350_111#_M1007_g N_A_469_47#_c_548_n 0.010041f $X=2.705 $Y=0.445
+ $X2=0 $Y2=0
cc_316 N_A_350_111#_M1008_g N_A_469_47#_c_548_n 0.0014829f $X=3.095 $Y=0.445
+ $X2=0 $Y2=0
cc_317 N_A_350_111#_c_288_n N_A_469_47#_c_548_n 0.014023f $X=1.89 $Y=0.765 $X2=0
+ $Y2=0
cc_318 N_A_350_111#_M1012_g N_A_469_47#_c_558_n 0.00813087f $X=2.76 $Y=2.695
+ $X2=0 $Y2=0
cc_319 N_A_350_111#_M1015_g N_A_469_47#_c_558_n 4.10552e-19 $X=3.12 $Y=2.695
+ $X2=0 $Y2=0
cc_320 N_A_350_111#_c_298_n N_A_469_47#_c_558_n 0.00224321f $X=2.732 $Y=2.235
+ $X2=0 $Y2=0
cc_321 N_A_350_111#_M1007_g N_A_469_47#_c_549_n 0.00839695f $X=2.705 $Y=0.445
+ $X2=0 $Y2=0
cc_322 N_A_350_111#_M1008_g N_A_469_47#_c_549_n 0.0123692f $X=3.095 $Y=0.445
+ $X2=0 $Y2=0
cc_323 N_A_350_111#_c_285_n N_A_469_47#_c_549_n 0.036977f $X=3.945 $Y=1.42 $X2=0
+ $Y2=0
cc_324 N_A_350_111#_c_289_n N_A_469_47#_c_549_n 0.022731f $X=2.795 $Y=1.34 $X2=0
+ $Y2=0
cc_325 N_A_350_111#_c_290_n N_A_469_47#_c_549_n 0.00111073f $X=2.795 $Y=1.34
+ $X2=0 $Y2=0
cc_326 N_A_350_111#_M1007_g N_A_469_47#_c_550_n 0.00419211f $X=2.705 $Y=0.445
+ $X2=0 $Y2=0
cc_327 N_A_350_111#_c_284_n N_A_469_47#_c_550_n 0.0122129f $X=2.63 $Y=1.685
+ $X2=0 $Y2=0
cc_328 N_A_350_111#_c_288_n N_A_469_47#_c_550_n 0.0120685f $X=1.89 $Y=0.765
+ $X2=0 $Y2=0
cc_329 N_A_350_111#_c_289_n N_A_469_47#_c_550_n 0.00193735f $X=2.795 $Y=1.34
+ $X2=0 $Y2=0
cc_330 N_A_350_111#_c_283_n N_A_469_47#_c_551_n 0.0122439f $X=2.005 $Y=1.525
+ $X2=0 $Y2=0
cc_331 N_A_350_111#_c_288_n N_A_469_47#_c_551_n 9.7067e-19 $X=1.89 $Y=0.765
+ $X2=0 $Y2=0
cc_332 N_A_350_111#_c_285_n N_A_469_47#_c_552_n 0.0224524f $X=3.945 $Y=1.42
+ $X2=0 $Y2=0
cc_333 N_A_350_111#_c_292_n N_A_469_47#_c_552_n 0.0208816f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_334 N_A_350_111#_c_293_n N_A_469_47#_c_552_n 0.00114872f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_335 N_A_350_111#_c_292_n N_A_469_47#_c_553_n 0.00114651f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_336 N_A_350_111#_c_293_n N_A_469_47#_c_553_n 0.0200799f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_337 N_A_350_111#_M1020_g N_A_969_407#_M1001_g 0.0215946f $X=4.425 $Y=0.445
+ $X2=0 $Y2=0
cc_338 N_A_350_111#_c_287_n N_A_969_407#_M1001_g 0.00105111f $X=4.435 $Y=1.335
+ $X2=0 $Y2=0
cc_339 N_A_350_111#_c_291_n N_A_969_407#_M1001_g 5.20629e-19 $X=4.435 $Y=1.42
+ $X2=0 $Y2=0
cc_340 N_A_350_111#_c_292_n N_A_969_407#_M1001_g 3.94195e-19 $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_341 N_A_350_111#_c_293_n N_A_969_407#_M1001_g 0.0205745f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_342 N_A_350_111#_M1020_g N_A_798_47#_c_842_n 0.0140618f $X=4.425 $Y=0.445
+ $X2=0 $Y2=0
cc_343 N_A_350_111#_c_292_n N_A_798_47#_c_842_n 0.0216526f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_344 N_A_350_111#_c_293_n N_A_798_47#_c_842_n 0.00116741f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_345 N_A_350_111#_M1017_g N_A_798_47#_c_837_n 0.00708262f $X=4.02 $Y=2.695
+ $X2=0 $Y2=0
cc_346 N_A_350_111#_c_286_n N_A_798_47#_c_837_n 0.0222802f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_347 N_A_350_111#_c_302_n N_A_798_47#_c_837_n 0.00163647f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_348 N_A_350_111#_c_292_n N_A_798_47#_c_838_n 0.00167494f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_349 N_A_350_111#_c_293_n N_A_798_47#_c_838_n 2.42473e-19 $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_350 N_A_350_111#_c_286_n N_A_798_47#_c_839_n 0.0137914f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_351 N_A_350_111#_c_291_n N_A_798_47#_c_839_n 0.00483218f $X=4.435 $Y=1.42
+ $X2=0 $Y2=0
cc_352 N_A_350_111#_c_292_n N_A_798_47#_c_839_n 0.00329828f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_353 N_A_350_111#_M1020_g N_A_798_47#_c_831_n 0.00295803f $X=4.425 $Y=0.445
+ $X2=0 $Y2=0
cc_354 N_A_350_111#_c_287_n N_A_798_47#_c_831_n 0.00834199f $X=4.435 $Y=1.335
+ $X2=0 $Y2=0
cc_355 N_A_350_111#_c_292_n N_A_798_47#_c_831_n 0.0237561f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_356 N_A_350_111#_c_293_n N_A_798_47#_c_831_n 0.00174446f $X=4.515 $Y=0.99
+ $X2=0 $Y2=0
cc_357 N_A_350_111#_c_286_n N_A_798_47#_c_832_n 0.00586457f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_358 N_A_350_111#_c_291_n N_A_798_47#_c_832_n 0.00824643f $X=4.435 $Y=1.42
+ $X2=0 $Y2=0
cc_359 N_A_350_111#_M1017_g N_A_798_47#_c_841_n 0.00942285f $X=4.02 $Y=2.695
+ $X2=0 $Y2=0
cc_360 N_A_350_111#_c_286_n N_A_798_47#_c_841_n 0.00738996f $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_361 N_A_350_111#_c_302_n N_A_798_47#_c_841_n 9.57793e-19 $X=4.11 $Y=2 $X2=0
+ $Y2=0
cc_362 N_A_350_111#_M1015_g N_VPWR_c_988_n 0.00569704f $X=3.12 $Y=2.695 $X2=0
+ $Y2=0
cc_363 N_A_350_111#_M1017_g N_VPWR_c_988_n 0.00302807f $X=4.02 $Y=2.695 $X2=0
+ $Y2=0
cc_364 N_A_350_111#_M1012_g N_VPWR_c_992_n 0.00309864f $X=2.76 $Y=2.695 $X2=0
+ $Y2=0
cc_365 N_A_350_111#_M1015_g N_VPWR_c_992_n 0.00475301f $X=3.12 $Y=2.695 $X2=0
+ $Y2=0
cc_366 N_A_350_111#_M1017_g N_VPWR_c_995_n 0.00476129f $X=4.02 $Y=2.695 $X2=0
+ $Y2=0
cc_367 N_A_350_111#_M1012_g N_VPWR_c_986_n 0.00503767f $X=2.76 $Y=2.695 $X2=0
+ $Y2=0
cc_368 N_A_350_111#_M1015_g N_VPWR_c_986_n 0.00904566f $X=3.12 $Y=2.695 $X2=0
+ $Y2=0
cc_369 N_A_350_111#_M1017_g N_VPWR_c_986_n 0.00924961f $X=4.02 $Y=2.695 $X2=0
+ $Y2=0
cc_370 N_A_350_111#_M1007_g N_VGND_c_1180_n 0.00231186f $X=2.705 $Y=0.445 $X2=0
+ $Y2=0
cc_371 N_A_350_111#_M1008_g N_VGND_c_1180_n 0.0122017f $X=3.095 $Y=0.445 $X2=0
+ $Y2=0
cc_372 N_A_350_111#_M1007_g N_VGND_c_1186_n 0.0054778f $X=2.705 $Y=0.445 $X2=0
+ $Y2=0
cc_373 N_A_350_111#_M1008_g N_VGND_c_1186_n 0.00486043f $X=3.095 $Y=0.445 $X2=0
+ $Y2=0
cc_374 N_A_350_111#_M1020_g N_VGND_c_1188_n 0.00366111f $X=4.425 $Y=0.445 $X2=0
+ $Y2=0
cc_375 N_A_350_111#_M1007_g N_VGND_c_1192_n 0.00760003f $X=2.705 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_A_350_111#_M1008_g N_VGND_c_1192_n 0.00447093f $X=3.095 $Y=0.445 $X2=0
+ $Y2=0
cc_377 N_A_350_111#_M1020_g N_VGND_c_1192_n 0.00585835f $X=4.425 $Y=0.445 $X2=0
+ $Y2=0
cc_378 N_A_27_111#_c_441_n N_A_469_47#_M1012_s 0.00299939f $X=2.9 $Y=2.98 $X2=0
+ $Y2=0
cc_379 N_A_27_111#_M1009_g N_A_469_47#_M1019_g 0.0387448f $X=3.525 $Y=0.445
+ $X2=0 $Y2=0
cc_380 N_A_27_111#_c_434_n N_A_469_47#_c_543_n 0.0238323f $X=3.51 $Y=1.595 $X2=0
+ $Y2=0
cc_381 N_A_27_111#_c_443_n N_A_469_47#_c_556_n 6.99375e-19 $X=2.985 $Y=2.895
+ $X2=0 $Y2=0
cc_382 N_A_27_111#_c_445_n N_A_469_47#_c_556_n 0.0127683f $X=3.07 $Y=2.11 $X2=0
+ $Y2=0
cc_383 N_A_27_111#_c_440_n N_A_469_47#_c_557_n 4.04787e-19 $X=1.405 $Y=2.47
+ $X2=0 $Y2=0
cc_384 N_A_27_111#_c_441_n N_A_469_47#_c_558_n 0.0196147f $X=2.9 $Y=2.98 $X2=0
+ $Y2=0
cc_385 N_A_27_111#_c_443_n N_A_469_47#_c_558_n 0.0347181f $X=2.985 $Y=2.895
+ $X2=0 $Y2=0
cc_386 N_A_27_111#_M1009_g N_A_469_47#_c_549_n 0.0121639f $X=3.525 $Y=0.445
+ $X2=0 $Y2=0
cc_387 N_A_27_111#_M1009_g N_A_469_47#_c_552_n 0.00118187f $X=3.525 $Y=0.445
+ $X2=0 $Y2=0
cc_388 N_A_27_111#_M1009_g N_A_469_47#_c_553_n 0.0238323f $X=3.525 $Y=0.445
+ $X2=0 $Y2=0
cc_389 N_A_27_111#_M1013_g N_A_798_47#_c_841_n 0.00130225f $X=3.63 $Y=2.695
+ $X2=0 $Y2=0
cc_390 N_A_27_111#_c_440_n A_112_481# 0.00182165f $X=1.405 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_391 N_A_27_111#_c_440_n N_VPWR_M1028_d 0.0021985f $X=1.405 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_392 N_A_27_111#_c_440_n N_VPWR_c_987_n 0.0171834f $X=1.405 $Y=2.47 $X2=0
+ $Y2=0
cc_393 N_A_27_111#_c_442_n N_VPWR_c_987_n 0.00161266f $X=1.575 $Y=2.98 $X2=0
+ $Y2=0
cc_394 N_A_27_111#_c_446_n N_VPWR_c_987_n 0.0110409f $X=0.27 $Y=2.55 $X2=0 $Y2=0
cc_395 N_A_27_111#_M1013_g N_VPWR_c_988_n 0.0188332f $X=3.63 $Y=2.695 $X2=0
+ $Y2=0
cc_396 N_A_27_111#_c_441_n N_VPWR_c_988_n 0.00880411f $X=2.9 $Y=2.98 $X2=0 $Y2=0
cc_397 N_A_27_111#_c_444_n N_VPWR_c_988_n 0.0121706f $X=3.405 $Y=2.11 $X2=0
+ $Y2=0
cc_398 N_A_27_111#_c_447_n N_VPWR_c_988_n 0.0112045f $X=3.57 $Y=2.03 $X2=0 $Y2=0
cc_399 N_A_27_111#_c_448_n N_VPWR_c_988_n 9.79582e-19 $X=3.57 $Y=2.03 $X2=0
+ $Y2=0
cc_400 N_A_27_111#_c_441_n N_VPWR_c_992_n 0.0908025f $X=2.9 $Y=2.98 $X2=0 $Y2=0
cc_401 N_A_27_111#_c_442_n N_VPWR_c_992_n 0.0114622f $X=1.575 $Y=2.98 $X2=0
+ $Y2=0
cc_402 N_A_27_111#_c_446_n N_VPWR_c_994_n 0.0220321f $X=0.27 $Y=2.55 $X2=0 $Y2=0
cc_403 N_A_27_111#_M1013_g N_VPWR_c_995_n 0.00422142f $X=3.63 $Y=2.695 $X2=0
+ $Y2=0
cc_404 N_A_27_111#_M1013_g N_VPWR_c_986_n 0.00790489f $X=3.63 $Y=2.695 $X2=0
+ $Y2=0
cc_405 N_A_27_111#_c_440_n N_VPWR_c_986_n 0.0217306f $X=1.405 $Y=2.47 $X2=0
+ $Y2=0
cc_406 N_A_27_111#_c_441_n N_VPWR_c_986_n 0.0546003f $X=2.9 $Y=2.98 $X2=0 $Y2=0
cc_407 N_A_27_111#_c_442_n N_VPWR_c_986_n 0.00657784f $X=1.575 $Y=2.98 $X2=0
+ $Y2=0
cc_408 N_A_27_111#_c_446_n N_VPWR_c_986_n 0.0125808f $X=0.27 $Y=2.55 $X2=0 $Y2=0
cc_409 N_A_27_111#_c_441_n A_567_475# 2.67089e-19 $X=2.9 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_410 N_A_27_111#_c_443_n A_567_475# 0.00486127f $X=2.985 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_411 N_A_27_111#_c_436_n N_VGND_c_1179_n 0.0151051f $X=0.28 $Y=0.765 $X2=0
+ $Y2=0
cc_412 N_A_27_111#_M1009_g N_VGND_c_1180_n 0.0126682f $X=3.525 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_27_111#_c_436_n N_VGND_c_1184_n 0.00838453f $X=0.28 $Y=0.765 $X2=0
+ $Y2=0
cc_414 N_A_27_111#_M1009_g N_VGND_c_1188_n 0.00486043f $X=3.525 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_A_27_111#_M1009_g N_VGND_c_1192_n 0.00450668f $X=3.525 $Y=0.445 $X2=0
+ $Y2=0
cc_416 N_A_27_111#_c_436_n N_VGND_c_1192_n 0.0109142f $X=0.28 $Y=0.765 $X2=0
+ $Y2=0
cc_417 N_A_469_47#_M1029_g N_A_969_407#_M1005_g 0.040843f $X=4.56 $Y=2.805 $X2=0
+ $Y2=0
cc_418 N_A_469_47#_c_540_n N_A_969_407#_M1001_g 0.0316795f $X=4.485 $Y=1.47
+ $X2=0 $Y2=0
cc_419 N_A_469_47#_M1029_g N_A_969_407#_c_696_n 9.94903e-19 $X=4.56 $Y=2.805
+ $X2=0 $Y2=0
cc_420 N_A_469_47#_M1029_g N_A_969_407#_c_697_n 0.0196496f $X=4.56 $Y=2.805
+ $X2=0 $Y2=0
cc_421 N_A_469_47#_c_552_n N_A_798_47#_c_842_n 0.00676209f $X=3.975 $Y=0.91
+ $X2=0 $Y2=0
cc_422 N_A_469_47#_c_553_n N_A_798_47#_c_842_n 6.78885e-19 $X=3.975 $Y=0.99
+ $X2=0 $Y2=0
cc_423 N_A_469_47#_M1029_g N_A_798_47#_c_837_n 0.0192988f $X=4.56 $Y=2.805 $X2=0
+ $Y2=0
cc_424 N_A_469_47#_M1029_g N_A_798_47#_c_838_n 0.00213287f $X=4.56 $Y=2.805
+ $X2=0 $Y2=0
cc_425 N_A_469_47#_c_540_n N_A_798_47#_c_839_n 6.09117e-19 $X=4.485 $Y=1.47
+ $X2=0 $Y2=0
cc_426 N_A_469_47#_M1029_g N_A_798_47#_c_839_n 0.0069242f $X=4.56 $Y=2.805 $X2=0
+ $Y2=0
cc_427 N_A_469_47#_c_540_n N_A_798_47#_c_832_n 0.00244464f $X=4.485 $Y=1.47
+ $X2=0 $Y2=0
cc_428 N_A_469_47#_M1029_g N_A_798_47#_c_841_n 0.0180753f $X=4.56 $Y=2.805 $X2=0
+ $Y2=0
cc_429 N_A_469_47#_M1029_g N_VPWR_c_995_n 0.00366854f $X=4.56 $Y=2.805 $X2=0
+ $Y2=0
cc_430 N_A_469_47#_M1029_g N_VPWR_c_986_n 0.00543558f $X=4.56 $Y=2.805 $X2=0
+ $Y2=0
cc_431 N_A_469_47#_c_544_n N_VGND_c_1179_n 0.00889519f $X=1.46 $Y=1.175 $X2=0
+ $Y2=0
cc_432 N_A_469_47#_c_546_n N_VGND_c_1179_n 0.012299f $X=1.545 $Y=0.35 $X2=0
+ $Y2=0
cc_433 N_A_469_47#_M1019_g N_VGND_c_1180_n 0.00241777f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_434 N_A_469_47#_c_545_n N_VGND_c_1180_n 0.00571183f $X=2.325 $Y=0.35 $X2=0
+ $Y2=0
cc_435 N_A_469_47#_c_548_n N_VGND_c_1180_n 0.0066371f $X=2.49 $Y=0.47 $X2=0
+ $Y2=0
cc_436 N_A_469_47#_c_549_n N_VGND_c_1180_n 0.0200812f $X=3.81 $Y=0.91 $X2=0
+ $Y2=0
cc_437 N_A_469_47#_c_545_n N_VGND_c_1186_n 0.0671602f $X=2.325 $Y=0.35 $X2=0
+ $Y2=0
cc_438 N_A_469_47#_c_546_n N_VGND_c_1186_n 0.0114622f $X=1.545 $Y=0.35 $X2=0
+ $Y2=0
cc_439 N_A_469_47#_M1019_g N_VGND_c_1188_n 0.00585385f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_440 N_A_469_47#_M1007_s N_VGND_c_1192_n 0.00232985f $X=2.345 $Y=0.235 $X2=0
+ $Y2=0
cc_441 N_A_469_47#_M1019_g N_VGND_c_1192_n 0.00663445f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_442 N_A_469_47#_c_545_n N_VGND_c_1192_n 0.0417963f $X=2.325 $Y=0.35 $X2=0
+ $Y2=0
cc_443 N_A_469_47#_c_546_n N_VGND_c_1192_n 0.00657784f $X=1.545 $Y=0.35 $X2=0
+ $Y2=0
cc_444 N_A_469_47#_c_549_n N_VGND_c_1192_n 0.0273182f $X=3.81 $Y=0.91 $X2=0
+ $Y2=0
cc_445 N_A_469_47#_c_552_n N_VGND_c_1192_n 0.0074215f $X=3.975 $Y=0.91 $X2=0
+ $Y2=0
cc_446 N_A_469_47#_c_544_n A_272_111# 0.00252746f $X=1.46 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_447 N_A_969_407#_M1001_g N_A_798_47#_M1031_g 0.0198932f $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_448 N_A_969_407#_c_684_n N_A_798_47#_M1031_g 0.00225828f $X=6.165 $Y=0.43
+ $X2=0 $Y2=0
cc_449 N_A_969_407#_M1005_g N_A_798_47#_M1026_g 0.010107f $X=4.95 $Y=2.805 $X2=0
+ $Y2=0
cc_450 N_A_969_407#_c_696_n N_A_798_47#_M1026_g 0.0228124f $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_451 N_A_969_407#_c_697_n N_A_798_47#_M1026_g 0.00807149f $X=5.01 $Y=2.2 $X2=0
+ $Y2=0
cc_452 N_A_969_407#_c_699_n N_A_798_47#_M1026_g 0.00371875f $X=6.26 $Y=1.95
+ $X2=0 $Y2=0
cc_453 N_A_969_407#_c_684_n N_A_798_47#_M1022_g 0.0130089f $X=6.165 $Y=0.43
+ $X2=0 $Y2=0
cc_454 N_A_969_407#_c_685_n N_A_798_47#_M1022_g 0.00634725f $X=6.245 $Y=1.275
+ $X2=0 $Y2=0
cc_455 N_A_969_407#_c_687_n N_A_798_47#_M1022_g 0.00425809f $X=6.165 $Y=1.095
+ $X2=0 $Y2=0
cc_456 N_A_969_407#_c_696_n N_A_798_47#_M1014_g 0.0198244f $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_457 N_A_969_407#_c_698_n N_A_798_47#_M1014_g 0.0132884f $X=6.26 $Y=2.9 $X2=0
+ $Y2=0
cc_458 N_A_969_407#_c_699_n N_A_798_47#_M1014_g 0.00931304f $X=6.26 $Y=1.95
+ $X2=0 $Y2=0
cc_459 N_A_969_407#_c_688_n N_A_798_47#_M1014_g 0.00742602f $X=6.26 $Y=1.785
+ $X2=0 $Y2=0
cc_460 N_A_969_407#_M1001_g N_A_798_47#_c_842_n 0.0130911f $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_461 N_A_969_407#_M1005_g N_A_798_47#_c_837_n 0.00133625f $X=4.95 $Y=2.805
+ $X2=0 $Y2=0
cc_462 N_A_969_407#_M1001_g N_A_798_47#_c_837_n 0.00113028f $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_463 N_A_969_407#_c_696_n N_A_798_47#_c_837_n 0.0203086f $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_464 N_A_969_407#_c_697_n N_A_798_47#_c_837_n 4.11234e-19 $X=5.01 $Y=2.2 $X2=0
+ $Y2=0
cc_465 N_A_969_407#_M1001_g N_A_798_47#_c_838_n 4.22378e-19 $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_466 N_A_969_407#_c_696_n N_A_798_47#_c_838_n 0.00107983f $X=6.095 $Y=2.2
+ $X2=0 $Y2=0
cc_467 N_A_969_407#_c_697_n N_A_798_47#_c_838_n 3.34149e-19 $X=5.01 $Y=2.2 $X2=0
+ $Y2=0
cc_468 N_A_969_407#_M1001_g N_A_798_47#_c_831_n 0.0167806f $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_469 N_A_969_407#_M1001_g N_A_798_47#_c_832_n 0.0180679f $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_470 N_A_969_407#_c_696_n N_A_798_47#_c_832_n 0.0129383f $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_471 N_A_969_407#_c_697_n N_A_798_47#_c_832_n 7.30771e-19 $X=5.01 $Y=2.2 $X2=0
+ $Y2=0
cc_472 N_A_969_407#_M1001_g N_A_798_47#_c_833_n 0.00793664f $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_473 N_A_969_407#_c_696_n N_A_798_47#_c_833_n 0.0341464f $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_474 N_A_969_407#_c_697_n N_A_798_47#_c_833_n 0.00256698f $X=5.01 $Y=2.2 $X2=0
+ $Y2=0
cc_475 N_A_969_407#_c_689_n N_A_798_47#_c_833_n 0.0261895f $X=6.292 $Y=1.44
+ $X2=0 $Y2=0
cc_476 N_A_969_407#_M1005_g N_A_798_47#_c_841_n 0.00106984f $X=4.95 $Y=2.805
+ $X2=0 $Y2=0
cc_477 N_A_969_407#_M1001_g N_A_798_47#_c_834_n 0.0128202f $X=4.965 $Y=0.445
+ $X2=0 $Y2=0
cc_478 N_A_969_407#_c_680_n N_A_798_47#_c_834_n 0.0117001f $X=7.985 $Y=1.38
+ $X2=0 $Y2=0
cc_479 N_A_969_407#_c_696_n N_A_798_47#_c_834_n 9.3988e-19 $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_480 N_A_969_407#_c_687_n N_A_798_47#_c_834_n 0.00617392f $X=6.165 $Y=1.095
+ $X2=0 $Y2=0
cc_481 N_A_969_407#_c_699_n N_A_798_47#_c_834_n 0.00134366f $X=6.26 $Y=1.95
+ $X2=0 $Y2=0
cc_482 N_A_969_407#_c_689_n N_A_798_47#_c_834_n 0.0193011f $X=6.292 $Y=1.44
+ $X2=0 $Y2=0
cc_483 N_A_969_407#_M1035_g N_A_1662_131#_c_937_n 0.00155932f $X=7.845 $Y=0.865
+ $X2=0 $Y2=0
cc_484 N_A_969_407#_M1024_g N_A_1662_131#_c_937_n 0.0157188f $X=8.235 $Y=0.865
+ $X2=0 $Y2=0
cc_485 N_A_969_407#_M1000_g N_A_1662_131#_c_943_n 0.00230429f $X=7.91 $Y=2.125
+ $X2=0 $Y2=0
cc_486 N_A_969_407#_M1003_g N_A_1662_131#_c_943_n 0.0197942f $X=8.27 $Y=2.125
+ $X2=0 $Y2=0
cc_487 N_A_969_407#_M1003_g N_A_1662_131#_c_939_n 0.00686573f $X=8.27 $Y=2.125
+ $X2=0 $Y2=0
cc_488 N_A_969_407#_c_683_n N_A_1662_131#_c_939_n 0.00812177f $X=8.252 $Y=1.38
+ $X2=0 $Y2=0
cc_489 N_A_969_407#_c_696_n N_VPWR_M1005_d 0.00742587f $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_490 N_A_969_407#_M1005_g N_VPWR_c_989_n 0.0134114f $X=4.95 $Y=2.805 $X2=0
+ $Y2=0
cc_491 N_A_969_407#_c_696_n N_VPWR_c_989_n 0.0220816f $X=6.095 $Y=2.2 $X2=0
+ $Y2=0
cc_492 N_A_969_407#_c_698_n N_VPWR_c_989_n 0.0173978f $X=6.26 $Y=2.9 $X2=0 $Y2=0
cc_493 N_A_969_407#_M1018_g N_VPWR_c_990_n 0.00356008f $X=7.015 $Y=2.435 $X2=0
+ $Y2=0
cc_494 N_A_969_407#_M1016_g N_VPWR_c_990_n 0.0249855f $X=7.375 $Y=2.435 $X2=0
+ $Y2=0
cc_495 N_A_969_407#_M1000_g N_VPWR_c_990_n 0.00747194f $X=7.91 $Y=2.125 $X2=0
+ $Y2=0
cc_496 N_A_969_407#_M1003_g N_VPWR_c_991_n 0.00396126f $X=8.27 $Y=2.125 $X2=0
+ $Y2=0
cc_497 N_A_969_407#_M1005_g N_VPWR_c_995_n 0.00508422f $X=4.95 $Y=2.805 $X2=0
+ $Y2=0
cc_498 N_A_969_407#_M1018_g N_VPWR_c_996_n 0.00520813f $X=7.015 $Y=2.435 $X2=0
+ $Y2=0
cc_499 N_A_969_407#_M1016_g N_VPWR_c_996_n 0.00461019f $X=7.375 $Y=2.435 $X2=0
+ $Y2=0
cc_500 N_A_969_407#_c_698_n N_VPWR_c_996_n 0.0197716f $X=6.26 $Y=2.9 $X2=0 $Y2=0
cc_501 N_A_969_407#_M1000_g N_VPWR_c_997_n 0.00301355f $X=7.91 $Y=2.125 $X2=0
+ $Y2=0
cc_502 N_A_969_407#_M1003_g N_VPWR_c_997_n 0.00301355f $X=8.27 $Y=2.125 $X2=0
+ $Y2=0
cc_503 N_A_969_407#_M1005_g N_VPWR_c_986_n 0.0103247f $X=4.95 $Y=2.805 $X2=0
+ $Y2=0
cc_504 N_A_969_407#_M1018_g N_VPWR_c_986_n 0.010695f $X=7.015 $Y=2.435 $X2=0
+ $Y2=0
cc_505 N_A_969_407#_M1016_g N_VPWR_c_986_n 0.00803623f $X=7.375 $Y=2.435 $X2=0
+ $Y2=0
cc_506 N_A_969_407#_M1000_g N_VPWR_c_986_n 0.00403185f $X=7.91 $Y=2.125 $X2=0
+ $Y2=0
cc_507 N_A_969_407#_M1003_g N_VPWR_c_986_n 0.00403185f $X=8.27 $Y=2.125 $X2=0
+ $Y2=0
cc_508 N_A_969_407#_c_698_n N_VPWR_c_986_n 0.0125705f $X=6.26 $Y=2.9 $X2=0 $Y2=0
cc_509 N_A_969_407#_c_696_n A_1152_361# 0.00551744f $X=6.095 $Y=2.2 $X2=-0.19
+ $Y2=-0.245
cc_510 N_A_969_407#_M1034_g N_Q_c_1096_n 0.0131746f $X=6.94 $Y=0.655 $X2=0 $Y2=0
cc_511 N_A_969_407#_M1002_g N_Q_c_1096_n 0.00220615f $X=7.3 $Y=0.655 $X2=0 $Y2=0
cc_512 N_A_969_407#_c_684_n N_Q_c_1096_n 0.0444625f $X=6.165 $Y=0.43 $X2=0 $Y2=0
cc_513 N_A_969_407#_M1018_g N_Q_c_1100_n 0.00114325f $X=7.015 $Y=2.435 $X2=0
+ $Y2=0
cc_514 N_A_969_407#_c_680_n N_Q_c_1100_n 0.00736279f $X=7.985 $Y=1.38 $X2=0
+ $Y2=0
cc_515 N_A_969_407#_c_686_n N_Q_c_1100_n 0.0265437f $X=7.46 $Y=1.44 $X2=0 $Y2=0
cc_516 N_A_969_407#_c_699_n N_Q_c_1100_n 0.0129575f $X=6.26 $Y=1.95 $X2=0 $Y2=0
cc_517 N_A_969_407#_M1018_g N_Q_c_1101_n 0.0215393f $X=7.015 $Y=2.435 $X2=0
+ $Y2=0
cc_518 N_A_969_407#_M1016_g N_Q_c_1101_n 0.00343098f $X=7.375 $Y=2.435 $X2=0
+ $Y2=0
cc_519 N_A_969_407#_c_699_n N_Q_c_1101_n 0.0796352f $X=6.26 $Y=1.95 $X2=0 $Y2=0
cc_520 N_A_969_407#_M1034_g N_Q_c_1097_n 0.0107261f $X=6.94 $Y=0.655 $X2=0 $Y2=0
cc_521 N_A_969_407#_M1002_g N_Q_c_1097_n 0.0144513f $X=7.3 $Y=0.655 $X2=0 $Y2=0
cc_522 N_A_969_407#_M1035_g N_Q_c_1097_n 0.014349f $X=7.845 $Y=0.865 $X2=0 $Y2=0
cc_523 N_A_969_407#_c_680_n N_Q_c_1097_n 0.00668576f $X=7.985 $Y=1.38 $X2=0
+ $Y2=0
cc_524 N_A_969_407#_M1024_g N_Q_c_1097_n 0.0013479f $X=8.235 $Y=0.865 $X2=0
+ $Y2=0
cc_525 N_A_969_407#_c_686_n N_Q_c_1097_n 0.0518455f $X=7.46 $Y=1.44 $X2=0 $Y2=0
cc_526 N_A_969_407#_M1034_g N_Q_c_1098_n 0.00114325f $X=6.94 $Y=0.655 $X2=0
+ $Y2=0
cc_527 N_A_969_407#_c_680_n N_Q_c_1098_n 0.00579521f $X=7.985 $Y=1.38 $X2=0
+ $Y2=0
cc_528 N_A_969_407#_c_684_n N_Q_c_1098_n 0.0121278f $X=6.165 $Y=0.43 $X2=0 $Y2=0
cc_529 N_A_969_407#_c_686_n N_Q_c_1098_n 0.0267729f $X=7.46 $Y=1.44 $X2=0 $Y2=0
cc_530 N_A_969_407#_M1018_g N_Q_c_1102_n 0.0107261f $X=7.015 $Y=2.435 $X2=0
+ $Y2=0
cc_531 N_A_969_407#_M1016_g N_Q_c_1102_n 0.0144069f $X=7.375 $Y=2.435 $X2=0
+ $Y2=0
cc_532 N_A_969_407#_M1000_g N_Q_c_1102_n 0.0129329f $X=7.91 $Y=2.125 $X2=0 $Y2=0
cc_533 N_A_969_407#_c_680_n N_Q_c_1102_n 0.00739163f $X=7.985 $Y=1.38 $X2=0
+ $Y2=0
cc_534 N_A_969_407#_M1003_g N_Q_c_1102_n 5.31026e-19 $X=8.27 $Y=2.125 $X2=0
+ $Y2=0
cc_535 N_A_969_407#_c_686_n N_Q_c_1102_n 0.0464463f $X=7.46 $Y=1.44 $X2=0 $Y2=0
cc_536 N_A_969_407#_M1002_g Q 9.69292e-19 $X=7.3 $Y=0.655 $X2=0 $Y2=0
cc_537 N_A_969_407#_M1016_g Q 0.00329557f $X=7.375 $Y=2.435 $X2=0 $Y2=0
cc_538 N_A_969_407#_M1035_g Q 0.00561715f $X=7.845 $Y=0.865 $X2=0 $Y2=0
cc_539 N_A_969_407#_M1000_g Q 0.00409172f $X=7.91 $Y=2.125 $X2=0 $Y2=0
cc_540 N_A_969_407#_c_679_n Q 0.00373879f $X=8.16 $Y=1.38 $X2=0 $Y2=0
cc_541 N_A_969_407#_c_680_n Q 0.0106345f $X=7.985 $Y=1.38 $X2=0 $Y2=0
cc_542 N_A_969_407#_M1024_g Q 0.00142824f $X=8.235 $Y=0.865 $X2=0 $Y2=0
cc_543 N_A_969_407#_M1003_g Q 0.0019826f $X=8.27 $Y=2.125 $X2=0 $Y2=0
cc_544 N_A_969_407#_c_686_n Q 0.0243669f $X=7.46 $Y=1.44 $X2=0 $Y2=0
cc_545 N_A_969_407#_M1001_g N_VGND_c_1181_n 0.0102986f $X=4.965 $Y=0.445 $X2=0
+ $Y2=0
cc_546 N_A_969_407#_c_684_n N_VGND_c_1181_n 0.0277529f $X=6.165 $Y=0.43 $X2=0
+ $Y2=0
cc_547 N_A_969_407#_M1034_g N_VGND_c_1182_n 0.00258847f $X=6.94 $Y=0.655 $X2=0
+ $Y2=0
cc_548 N_A_969_407#_M1002_g N_VGND_c_1182_n 0.0163437f $X=7.3 $Y=0.655 $X2=0
+ $Y2=0
cc_549 N_A_969_407#_M1035_g N_VGND_c_1182_n 0.00456379f $X=7.845 $Y=0.865 $X2=0
+ $Y2=0
cc_550 N_A_969_407#_M1024_g N_VGND_c_1183_n 0.00385603f $X=8.235 $Y=0.865 $X2=0
+ $Y2=0
cc_551 N_A_969_407#_M1001_g N_VGND_c_1188_n 0.00380541f $X=4.965 $Y=0.445 $X2=0
+ $Y2=0
cc_552 N_A_969_407#_M1034_g N_VGND_c_1189_n 0.00549284f $X=6.94 $Y=0.655 $X2=0
+ $Y2=0
cc_553 N_A_969_407#_M1002_g N_VGND_c_1189_n 0.00486043f $X=7.3 $Y=0.655 $X2=0
+ $Y2=0
cc_554 N_A_969_407#_c_684_n N_VGND_c_1189_n 0.019758f $X=6.165 $Y=0.43 $X2=0
+ $Y2=0
cc_555 N_A_969_407#_M1035_g N_VGND_c_1190_n 0.00399858f $X=7.845 $Y=0.865 $X2=0
+ $Y2=0
cc_556 N_A_969_407#_M1024_g N_VGND_c_1190_n 0.00385415f $X=8.235 $Y=0.865 $X2=0
+ $Y2=0
cc_557 N_A_969_407#_M1022_d N_VGND_c_1192_n 0.0023218f $X=6.025 $Y=0.235 $X2=0
+ $Y2=0
cc_558 N_A_969_407#_M1001_g N_VGND_c_1192_n 0.00654897f $X=4.965 $Y=0.445 $X2=0
+ $Y2=0
cc_559 N_A_969_407#_M1034_g N_VGND_c_1192_n 0.0111098f $X=6.94 $Y=0.655 $X2=0
+ $Y2=0
cc_560 N_A_969_407#_M1002_g N_VGND_c_1192_n 0.00814425f $X=7.3 $Y=0.655 $X2=0
+ $Y2=0
cc_561 N_A_969_407#_M1035_g N_VGND_c_1192_n 0.0046122f $X=7.845 $Y=0.865 $X2=0
+ $Y2=0
cc_562 N_A_969_407#_M1024_g N_VGND_c_1192_n 0.0046122f $X=8.235 $Y=0.865 $X2=0
+ $Y2=0
cc_563 N_A_969_407#_c_684_n N_VGND_c_1192_n 0.012508f $X=6.165 $Y=0.43 $X2=0
+ $Y2=0
cc_564 N_A_798_47#_c_841_n N_VPWR_c_988_n 0.0148281f $X=4.235 $Y=2.805 $X2=0
+ $Y2=0
cc_565 N_A_798_47#_M1026_g N_VPWR_c_989_n 0.0161279f $X=5.685 $Y=2.435 $X2=0
+ $Y2=0
cc_566 N_A_798_47#_M1014_g N_VPWR_c_989_n 0.00244413f $X=6.045 $Y=2.435 $X2=0
+ $Y2=0
cc_567 N_A_798_47#_c_841_n N_VPWR_c_995_n 0.0222658f $X=4.235 $Y=2.805 $X2=0
+ $Y2=0
cc_568 N_A_798_47#_M1026_g N_VPWR_c_996_n 0.00461019f $X=5.685 $Y=2.435 $X2=0
+ $Y2=0
cc_569 N_A_798_47#_M1014_g N_VPWR_c_996_n 0.00520813f $X=6.045 $Y=2.435 $X2=0
+ $Y2=0
cc_570 N_A_798_47#_M1026_g N_VPWR_c_986_n 0.00803623f $X=5.685 $Y=2.435 $X2=0
+ $Y2=0
cc_571 N_A_798_47#_M1014_g N_VPWR_c_986_n 0.010695f $X=6.045 $Y=2.435 $X2=0
+ $Y2=0
cc_572 N_A_798_47#_c_841_n N_VPWR_c_986_n 0.0185853f $X=4.235 $Y=2.805 $X2=0
+ $Y2=0
cc_573 N_A_798_47#_M1022_g N_Q_c_1096_n 0.00138464f $X=5.95 $Y=0.655 $X2=0 $Y2=0
cc_574 N_A_798_47#_M1014_g N_Q_c_1100_n 3.80064e-19 $X=6.045 $Y=2.435 $X2=0
+ $Y2=0
cc_575 N_A_798_47#_M1014_g N_Q_c_1101_n 0.00221488f $X=6.045 $Y=2.435 $X2=0
+ $Y2=0
cc_576 N_A_798_47#_M1022_g N_Q_c_1098_n 3.9607e-19 $X=5.95 $Y=0.655 $X2=0 $Y2=0
cc_577 N_A_798_47#_M1031_g N_VGND_c_1181_n 0.0217652f $X=5.59 $Y=0.655 $X2=0
+ $Y2=0
cc_578 N_A_798_47#_M1022_g N_VGND_c_1181_n 0.00354111f $X=5.95 $Y=0.655 $X2=0
+ $Y2=0
cc_579 N_A_798_47#_c_842_n N_VGND_c_1181_n 0.027587f $X=4.86 $Y=0.47 $X2=0 $Y2=0
cc_580 N_A_798_47#_c_831_n N_VGND_c_1181_n 0.0325067f $X=4.945 $Y=1.275 $X2=0
+ $Y2=0
cc_581 N_A_798_47#_c_833_n N_VGND_c_1181_n 0.0276535f $X=5.805 $Y=1.44 $X2=0
+ $Y2=0
cc_582 N_A_798_47#_c_842_n N_VGND_c_1188_n 0.0478409f $X=4.86 $Y=0.47 $X2=0
+ $Y2=0
cc_583 N_A_798_47#_M1031_g N_VGND_c_1189_n 0.00486043f $X=5.59 $Y=0.655 $X2=0
+ $Y2=0
cc_584 N_A_798_47#_M1022_g N_VGND_c_1189_n 0.00549284f $X=5.95 $Y=0.655 $X2=0
+ $Y2=0
cc_585 N_A_798_47#_M1019_d N_VGND_c_1192_n 0.0032541f $X=3.99 $Y=0.235 $X2=0
+ $Y2=0
cc_586 N_A_798_47#_M1031_g N_VGND_c_1192_n 0.00814425f $X=5.59 $Y=0.655 $X2=0
+ $Y2=0
cc_587 N_A_798_47#_M1022_g N_VGND_c_1192_n 0.0111098f $X=5.95 $Y=0.655 $X2=0
+ $Y2=0
cc_588 N_A_798_47#_c_842_n N_VGND_c_1192_n 0.0354862f $X=4.86 $Y=0.47 $X2=0
+ $Y2=0
cc_589 N_A_798_47#_c_842_n A_900_47# 0.0109435f $X=4.86 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_590 N_A_1662_131#_c_943_n N_VPWR_c_990_n 0.0106412f $X=8.485 $Y=1.95 $X2=0
+ $Y2=0
cc_591 N_A_1662_131#_M1004_g N_VPWR_c_991_n 0.0305685f $X=9.24 $Y=2.465 $X2=0
+ $Y2=0
cc_592 N_A_1662_131#_M1006_g N_VPWR_c_991_n 0.004655f $X=9.6 $Y=2.465 $X2=0
+ $Y2=0
cc_593 N_A_1662_131#_c_943_n N_VPWR_c_991_n 0.0470338f $X=8.485 $Y=1.95 $X2=0
+ $Y2=0
cc_594 N_A_1662_131#_c_938_n N_VPWR_c_991_n 0.0274868f $X=9.29 $Y=1.47 $X2=0
+ $Y2=0
cc_595 N_A_1662_131#_c_940_n N_VPWR_c_991_n 9.85761e-19 $X=9.6 $Y=1.47 $X2=0
+ $Y2=0
cc_596 N_A_1662_131#_M1004_g N_VPWR_c_998_n 0.00486043f $X=9.24 $Y=2.465 $X2=0
+ $Y2=0
cc_597 N_A_1662_131#_M1006_g N_VPWR_c_998_n 0.00526721f $X=9.6 $Y=2.465 $X2=0
+ $Y2=0
cc_598 N_A_1662_131#_M1004_g N_VPWR_c_986_n 0.00814425f $X=9.24 $Y=2.465 $X2=0
+ $Y2=0
cc_599 N_A_1662_131#_M1006_g N_VPWR_c_986_n 0.0101917f $X=9.6 $Y=2.465 $X2=0
+ $Y2=0
cc_600 N_A_1662_131#_c_943_n N_VPWR_c_986_n 0.013775f $X=8.485 $Y=1.95 $X2=0
+ $Y2=0
cc_601 N_A_1662_131#_c_937_n N_Q_c_1097_n 0.0104715f $X=8.45 $Y=0.865 $X2=0
+ $Y2=0
cc_602 N_A_1662_131#_c_943_n N_Q_c_1102_n 0.00545125f $X=8.485 $Y=1.95 $X2=0
+ $Y2=0
cc_603 N_A_1662_131#_c_937_n Q 0.0120515f $X=8.45 $Y=0.865 $X2=0 $Y2=0
cc_604 N_A_1662_131#_c_943_n Q 0.0086565f $X=8.485 $Y=1.95 $X2=0 $Y2=0
cc_605 N_A_1662_131#_c_939_n Q 0.0195264f $X=8.467 $Y=1.47 $X2=0 $Y2=0
cc_606 N_A_1662_131#_M1027_g N_Q_N_c_1164_n 0.00323713f $X=9.225 $Y=0.685 $X2=0
+ $Y2=0
cc_607 N_A_1662_131#_M1004_g N_Q_N_c_1164_n 0.00440897f $X=9.24 $Y=2.465 $X2=0
+ $Y2=0
cc_608 N_A_1662_131#_M1030_g N_Q_N_c_1164_n 0.0239229f $X=9.585 $Y=0.685 $X2=0
+ $Y2=0
cc_609 N_A_1662_131#_M1006_g N_Q_N_c_1164_n 0.0313505f $X=9.6 $Y=2.465 $X2=0
+ $Y2=0
cc_610 N_A_1662_131#_c_938_n N_Q_N_c_1164_n 0.0250833f $X=9.29 $Y=1.47 $X2=0
+ $Y2=0
cc_611 N_A_1662_131#_c_940_n N_Q_N_c_1164_n 0.013006f $X=9.6 $Y=1.47 $X2=0 $Y2=0
cc_612 N_A_1662_131#_c_937_n N_VGND_c_1182_n 0.00316551f $X=8.45 $Y=0.865 $X2=0
+ $Y2=0
cc_613 N_A_1662_131#_M1027_g N_VGND_c_1183_n 0.0234518f $X=9.225 $Y=0.685 $X2=0
+ $Y2=0
cc_614 N_A_1662_131#_M1030_g N_VGND_c_1183_n 0.00336955f $X=9.585 $Y=0.685 $X2=0
+ $Y2=0
cc_615 N_A_1662_131#_c_937_n N_VGND_c_1183_n 0.033035f $X=8.45 $Y=0.865 $X2=0
+ $Y2=0
cc_616 N_A_1662_131#_c_938_n N_VGND_c_1183_n 0.0275493f $X=9.29 $Y=1.47 $X2=0
+ $Y2=0
cc_617 N_A_1662_131#_c_940_n N_VGND_c_1183_n 5.79521e-19 $X=9.6 $Y=1.47 $X2=0
+ $Y2=0
cc_618 N_A_1662_131#_c_937_n N_VGND_c_1190_n 0.00658678f $X=8.45 $Y=0.865 $X2=0
+ $Y2=0
cc_619 N_A_1662_131#_M1027_g N_VGND_c_1191_n 0.00461019f $X=9.225 $Y=0.685 $X2=0
+ $Y2=0
cc_620 N_A_1662_131#_M1030_g N_VGND_c_1191_n 0.00520813f $X=9.585 $Y=0.685 $X2=0
+ $Y2=0
cc_621 N_A_1662_131#_M1027_g N_VGND_c_1192_n 0.00803623f $X=9.225 $Y=0.685 $X2=0
+ $Y2=0
cc_622 N_A_1662_131#_M1030_g N_VGND_c_1192_n 0.0104f $X=9.585 $Y=0.685 $X2=0
+ $Y2=0
cc_623 N_A_1662_131#_c_937_n N_VGND_c_1192_n 0.00992454f $X=8.45 $Y=0.865 $X2=0
+ $Y2=0
cc_624 N_VPWR_c_990_n N_Q_c_1101_n 0.0311153f $X=7.59 $Y=2.3 $X2=0 $Y2=0
cc_625 N_VPWR_c_996_n N_Q_c_1101_n 0.0197716f $X=7.425 $Y=3.33 $X2=0 $Y2=0
cc_626 N_VPWR_c_986_n N_Q_c_1101_n 0.0125705f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_627 N_VPWR_M1016_d N_Q_c_1102_n 0.00381132f $X=7.45 $Y=1.805 $X2=0 $Y2=0
cc_628 N_VPWR_c_990_n N_Q_c_1102_n 0.0209601f $X=7.59 $Y=2.3 $X2=0 $Y2=0
cc_629 N_VPWR_c_986_n A_1863_367# 0.00899413f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_630 N_VPWR_c_986_n N_Q_N_M1006_d 0.00219599f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_631 N_VPWR_c_991_n N_Q_N_c_1164_n 0.0431709f $X=9.025 $Y=1.98 $X2=0 $Y2=0
cc_632 N_VPWR_c_998_n N_Q_N_c_1164_n 0.0207378f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_633 N_VPWR_c_986_n N_Q_N_c_1164_n 0.0130193f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_634 N_Q_c_1102_n A_1418_361# 0.00366293f $X=7.805 $Y=1.87 $X2=-0.19
+ $Y2=-0.245
cc_635 N_Q_c_1097_n N_VGND_M1002_d 0.00427535f $X=7.805 $Y=1.01 $X2=0 $Y2=0
cc_636 N_Q_c_1096_n N_VGND_c_1182_n 0.0160595f $X=6.725 $Y=0.43 $X2=0 $Y2=0
cc_637 N_Q_c_1097_n N_VGND_c_1182_n 0.0210003f $X=7.805 $Y=1.01 $X2=0 $Y2=0
cc_638 N_Q_c_1096_n N_VGND_c_1189_n 0.019758f $X=6.725 $Y=0.43 $X2=0 $Y2=0
cc_639 N_Q_M1034_s N_VGND_c_1192_n 0.0023218f $X=6.58 $Y=0.235 $X2=0 $Y2=0
cc_640 N_Q_c_1096_n N_VGND_c_1192_n 0.012508f $X=6.725 $Y=0.43 $X2=0 $Y2=0
cc_641 N_Q_c_1097_n A_1403_47# 0.00366293f $X=7.805 $Y=1.01 $X2=-0.19 $Y2=-0.245
cc_642 N_Q_c_1097_n A_1584_131# 0.00412065f $X=7.805 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_643 N_Q_N_c_1164_n N_VGND_c_1183_n 0.0288715f $X=9.8 $Y=0.43 $X2=0 $Y2=0
cc_644 N_Q_N_c_1164_n N_VGND_c_1191_n 0.0207694f $X=9.8 $Y=0.43 $X2=0 $Y2=0
cc_645 N_Q_N_c_1164_n N_VGND_c_1192_n 0.0131509f $X=9.8 $Y=0.43 $X2=0 $Y2=0
cc_646 N_VGND_c_1192_n A_556_47# 0.00346804f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_647 N_VGND_c_1192_n A_720_47# 0.00345315f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_648 N_VGND_c_1192_n A_900_47# 0.00316843f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_649 N_VGND_c_1192_n A_1133_47# 0.00899413f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_650 N_VGND_c_1192_n A_1403_47# 0.00899413f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
