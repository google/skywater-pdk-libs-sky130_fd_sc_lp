* File: sky130_fd_sc_lp__o211a_1.spice
* Created: Fri Aug 28 11:01:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211a_1.pex.spice"
.subckt sky130_fd_sc_lp__o211a_1  VNB VPB A1 A2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_237#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_266_49#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1974 AS=0.2226 PD=1.31 PS=2.21 NRD=13.56 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1005 N_A_266_49#_M1005_d N_A2_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1974 PD=1.23 PS=1.31 NRD=7.848 NRS=13.56 M=1 R=5.6 SA=75000.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1008 A_581_49# N_B1_M1008_g N_A_266_49#_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1638 PD=1.05 PS=1.23 NRD=7.14 NRS=7.848 M=1 R=5.6 SA=75001.3
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_80_237#_M1009_d N_C1_M1009_g A_581_49# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_80_237#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.3339 PD=1.88 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1000 A_365_367# N_A1_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3906 PD=1.47 PS=1.88 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_80_237#_M1001_d N_A2_M1001_g A_365_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1323 PD=1.65 PS=1.47 NRD=8.5892 NRS=7.8012 M=1 R=8.4 SA=75001.3
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_A_80_237#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=7.8012 NRS=8.5892 M=1 R=8.4 SA=75001.9
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1006 N_A_80_237#_M1006_d N_C1_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=9.3772 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o211a_1.pxi.spice"
*
.ends
*
*
