* File: sky130_fd_sc_lp__sdlclkp_4.pxi.spice
* Created: Wed Sep  2 10:37:18 2020
* 
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%SCE N_SCE_M1022_g N_SCE_M1014_g N_SCE_c_181_n
+ N_SCE_c_182_n SCE SCE SCE SCE SCE N_SCE_c_184_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%SCE
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%GATE N_GATE_M1019_g N_GATE_M1012_g
+ N_GATE_c_215_n GATE GATE GATE N_GATE_c_217_n N_GATE_c_218_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%GATE
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%A_252_361# N_A_252_361#_M1017_s
+ N_A_252_361#_M1026_s N_A_252_361#_c_286_n N_A_252_361#_c_287_n
+ N_A_252_361#_c_288_n N_A_252_361#_c_289_n N_A_252_361#_c_290_n
+ N_A_252_361#_M1027_g N_A_252_361#_c_272_n N_A_252_361#_c_273_n
+ N_A_252_361#_c_274_n N_A_252_361#_c_292_n N_A_252_361#_M1015_g
+ N_A_252_361#_c_275_n N_A_252_361#_c_276_n N_A_252_361#_c_277_n
+ N_A_252_361#_M1011_g N_A_252_361#_M1025_g N_A_252_361#_c_278_n
+ N_A_252_361#_c_294_n N_A_252_361#_c_279_n N_A_252_361#_c_280_n
+ N_A_252_361#_c_281_n N_A_252_361#_c_282_n N_A_252_361#_c_283_n
+ N_A_252_361#_c_296_n N_A_252_361#_c_297_n N_A_252_361#_c_284_n
+ N_A_252_361#_c_285_n PM_SKY130_FD_SC_LP__SDLCLKP_4%A_252_361#
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%A_335_70# N_A_335_70#_M1027_d
+ N_A_335_70#_M1015_d N_A_335_70#_c_419_n N_A_335_70#_M1020_g
+ N_A_335_70#_c_420_n N_A_335_70#_c_421_n N_A_335_70#_M1016_g
+ N_A_335_70#_c_423_n N_A_335_70#_c_424_n N_A_335_70#_c_425_n
+ N_A_335_70#_c_426_n N_A_335_70#_c_434_n N_A_335_70#_c_427_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%A_335_70#
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%A_762_107# N_A_762_107#_M1004_d
+ N_A_762_107#_M1005_d N_A_762_107#_M1009_g N_A_762_107#_M1000_g
+ N_A_762_107#_c_495_n N_A_762_107#_M1003_g N_A_762_107#_c_496_n
+ N_A_762_107#_M1007_g N_A_762_107#_c_506_n N_A_762_107#_c_520_n
+ N_A_762_107#_c_497_n N_A_762_107#_c_508_n N_A_762_107#_c_563_p
+ N_A_762_107#_c_564_p N_A_762_107#_c_569_p N_A_762_107#_c_509_n
+ N_A_762_107#_c_498_n N_A_762_107#_c_511_n N_A_762_107#_c_499_n
+ N_A_762_107#_c_512_n N_A_762_107#_c_513_n N_A_762_107#_c_500_n
+ N_A_762_107#_c_501_n N_A_762_107#_c_502_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%A_762_107#
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%A_634_133# N_A_634_133#_M1011_d
+ N_A_634_133#_M1020_d N_A_634_133#_c_635_n N_A_634_133#_M1004_g
+ N_A_634_133#_M1005_g N_A_634_133#_c_636_n N_A_634_133#_c_637_n
+ N_A_634_133#_c_638_n N_A_634_133#_c_639_n N_A_634_133#_c_640_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%A_634_133#
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%CLK N_CLK_M1017_g N_CLK_c_706_n N_CLK_M1026_g
+ N_CLK_M1002_g N_CLK_c_707_n N_CLK_M1018_g CLK CLK N_CLK_c_705_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%CLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%A_1275_367# N_A_1275_367#_M1003_d
+ N_A_1275_367#_M1018_d N_A_1275_367#_M1001_g N_A_1275_367#_c_758_n
+ N_A_1275_367#_M1006_g N_A_1275_367#_M1008_g N_A_1275_367#_c_760_n
+ N_A_1275_367#_M1010_g N_A_1275_367#_M1013_g N_A_1275_367#_c_762_n
+ N_A_1275_367#_M1021_g N_A_1275_367#_M1023_g N_A_1275_367#_c_764_n
+ N_A_1275_367#_M1024_g N_A_1275_367#_c_779_n N_A_1275_367#_c_765_n
+ N_A_1275_367#_c_766_n N_A_1275_367#_c_785_n N_A_1275_367#_c_788_n
+ N_A_1275_367#_c_767_n N_A_1275_367#_c_828_p N_A_1275_367#_c_793_n
+ N_A_1275_367#_c_796_n N_A_1275_367#_c_768_n N_A_1275_367#_c_769_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%A_1275_367#
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%VPWR N_VPWR_M1022_s N_VPWR_M1015_s
+ N_VPWR_M1000_d N_VPWR_M1026_d N_VPWR_M1007_d N_VPWR_M1008_s N_VPWR_M1023_s
+ N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n N_VPWR_c_883_n N_VPWR_c_926_n
+ N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n N_VPWR_c_888_n
+ N_VPWR_c_889_n N_VPWR_c_914_n VPWR N_VPWR_c_890_n N_VPWR_c_891_n
+ N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n
+ N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_899_n N_VPWR_c_879_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%VPWR
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%A_134_70# N_A_134_70#_M1014_d
+ N_A_134_70#_M1011_s N_A_134_70#_M1019_d N_A_134_70#_M1020_s
+ N_A_134_70#_c_995_n N_A_134_70#_c_998_n N_A_134_70#_c_999_n
+ N_A_134_70#_c_1000_n N_A_134_70#_c_1001_n N_A_134_70#_c_1002_n
+ N_A_134_70#_c_996_n N_A_134_70#_c_1068_p N_A_134_70#_c_1004_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%A_134_70#
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%GCLK N_GCLK_M1006_d N_GCLK_M1021_d
+ N_GCLK_M1001_d N_GCLK_M1013_d N_GCLK_c_1074_n N_GCLK_c_1117_p N_GCLK_c_1070_n
+ N_GCLK_c_1071_n N_GCLK_c_1089_n N_GCLK_c_1093_n N_GCLK_c_1095_n GCLK GCLK GCLK
+ GCLK GCLK PM_SKY130_FD_SC_LP__SDLCLKP_4%GCLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_4%VGND N_VGND_M1014_s N_VGND_M1012_d
+ N_VGND_M1009_d N_VGND_M1017_d N_VGND_M1006_s N_VGND_M1010_s N_VGND_M1024_s
+ N_VGND_c_1124_n N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n
+ N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n N_VGND_c_1131_n
+ N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n VGND N_VGND_c_1135_n
+ N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n N_VGND_c_1139_n
+ N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n N_VGND_c_1143_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_4%VGND
cc_1 VNB N_SCE_M1022_g 0.00176214f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_2 VNB N_SCE_M1014_g 0.0256345f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.56
cc_3 VNB N_SCE_c_181_n 0.0354816f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.105
cc_4 VNB N_SCE_c_182_n 0.0229255f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.625
cc_5 VNB SCE 0.0358644f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_SCE_c_184_n 0.0358859f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_7 VNB N_GATE_M1019_g 0.0028449f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_8 VNB N_GATE_M1012_g 0.0215869f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.56
cc_9 VNB N_GATE_c_215_n 0.0590441f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.475
cc_10 VNB GATE 0.015038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_GATE_c_217_n 0.0166166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_GATE_c_218_n 0.00159914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_252_361#_M1027_g 0.0380805f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_14 VNB N_A_252_361#_c_272_n 0.0151917f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_A_252_361#_c_273_n 0.00679905f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_16 VNB N_A_252_361#_c_274_n 0.0177835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_252_361#_c_275_n 0.00917919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_252_361#_c_276_n 0.0295676f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_19 VNB N_A_252_361#_c_277_n 0.0175098f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.925
cc_20 VNB N_A_252_361#_c_278_n 0.0066402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_252_361#_c_279_n 0.0115749f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=2.405
cc_22 VNB N_A_252_361#_c_280_n 0.0358268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_252_361#_c_281_n 0.0974324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_252_361#_c_282_n 0.0124782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_252_361#_c_283_n 0.0190108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_252_361#_c_284_n 0.00979406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_252_361#_c_285_n 0.0111148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_335_70#_c_419_n 0.00719266f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.56
cc_29 VNB N_A_335_70#_c_420_n 0.00876873f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.475
cc_30 VNB N_A_335_70#_c_421_n 0.0177961f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_31 VNB N_A_335_70#_M1016_g 0.0232939f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_A_335_70#_c_423_n 0.0038743f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_33 VNB N_A_335_70#_c_424_n 0.00945614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_335_70#_c_425_n 0.00644325f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.925
cc_35 VNB N_A_335_70#_c_426_n 0.00634008f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.12
cc_36 VNB N_A_335_70#_c_427_n 0.00913795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_762_107#_M1009_g 0.038498f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.105
cc_38 VNB N_A_762_107#_c_495_n 0.0195656f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_39 VNB N_A_762_107#_c_496_n 0.0323047f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_40 VNB N_A_762_107#_c_497_n 0.00618598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_762_107#_c_498_n 0.00165104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_762_107#_c_499_n 0.00243007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_762_107#_c_500_n 0.00478538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_762_107#_c_501_n 0.0125011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_762_107#_c_502_n 0.00996867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_634_133#_c_635_n 0.0228858f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.56
cc_47 VNB N_A_634_133#_c_636_n 0.00135804f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_48 VNB N_A_634_133#_c_637_n 0.00108343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_634_133#_c_638_n 0.0181636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_634_133#_c_639_n 0.00192145f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_51 VNB N_A_634_133#_c_640_n 0.0382634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_CLK_M1017_g 0.0539035f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_53 VNB N_CLK_M1002_g 0.0236372f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=0.955
cc_54 VNB CLK 0.00916617f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_55 VNB N_CLK_c_705_n 0.056442f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.925
cc_56 VNB N_A_1275_367#_M1001_g 0.00645296f $X=-0.19 $Y=-0.245 $X2=0.312
+ $Y2=1.105
cc_57 VNB N_A_1275_367#_c_758_n 0.0184016f $X=-0.19 $Y=-0.245 $X2=0.387
+ $Y2=1.105
cc_58 VNB N_A_1275_367#_M1008_g 0.00663333f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_59 VNB N_A_1275_367#_c_760_n 0.0159966f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_60 VNB N_A_1275_367#_M1013_g 0.00661601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1275_367#_c_762_n 0.0159715f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.12
cc_62 VNB N_A_1275_367#_M1023_g 0.0105915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1275_367#_c_764_n 0.0209288f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.295
cc_64 VNB N_A_1275_367#_c_765_n 0.0136391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1275_367#_c_766_n 0.0016618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1275_367#_c_767_n 0.00128304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1275_367#_c_768_n 0.00337696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1275_367#_c_769_n 0.100316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VPWR_c_879_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_134_70#_c_995_n 0.0140121f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.625
cc_71 VNB N_A_134_70#_c_996_n 0.00478567f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_72 VNB N_GCLK_c_1070_n 0.00244579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_GCLK_c_1071_n 0.00235275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB GCLK 0.00280469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB GCLK 0.00124196f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=2.035
cc_76 VNB N_VGND_c_1124_n 0.0147631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1125_n 0.0211201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1126_n 0.017937f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_79 VNB N_VGND_c_1127_n 0.00833135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1128_n 0.00658906f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.665
cc_81 VNB N_VGND_c_1129_n 0.00902309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1130_n 3.10897e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1131_n 0.0111894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1132_n 0.047921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1133_n 0.0325448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1134_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1135_n 0.0617961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1136_n 0.0277446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1137_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1138_n 0.0136917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1139_n 0.00596278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1140_n 0.0127525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1141_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1142_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1143_n 0.467455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VPB N_SCE_M1022_g 0.0538209f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_97 VPB SCE 0.0348193f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_98 VPB N_GATE_M1019_g 0.0426537f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_99 VPB GATE 0.0111206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_GATE_c_218_n 0.00302686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_252_361#_c_286_n 0.0636605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_252_361#_c_287_n 0.029045f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.105
cc_103 VPB N_A_252_361#_c_288_n 0.00906035f $X=-0.19 $Y=1.655 $X2=0.387
+ $Y2=0.955
cc_104 VPB N_A_252_361#_c_289_n 0.159597f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.105
cc_105 VPB N_A_252_361#_c_290_n 0.0120406f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.475
cc_106 VPB N_A_252_361#_c_274_n 0.00591872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_252_361#_c_292_n 0.0179455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_252_361#_M1025_g 0.0307837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_252_361#_c_294_n 0.00566813f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=2.035
cc_110 VPB N_A_252_361#_c_283_n 0.0077153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_252_361#_c_296_n 0.00430241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_252_361#_c_297_n 0.0085966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_335_70#_c_419_n 0.0147646f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.56
cc_114 VPB N_A_335_70#_M1020_g 0.0462049f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.105
cc_115 VPB N_A_335_70#_c_420_n 0.00902132f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.475
cc_116 VPB N_A_335_70#_c_421_n 0.00661778f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_117 VPB N_A_335_70#_c_423_n 0.00127355f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_118 VPB N_A_335_70#_c_425_n 0.00228088f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.925
cc_119 VPB N_A_335_70#_c_434_n 0.0140016f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=2.035
cc_120 VPB N_A_335_70#_c_427_n 0.0271984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_762_107#_M1009_g 0.00583724f $X=-0.19 $Y=1.655 $X2=0.312
+ $Y2=1.105
cc_122 VPB N_A_762_107#_M1000_g 0.0261812f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.475
cc_123 VPB N_A_762_107#_M1007_g 0.0203812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_762_107#_c_506_n 0.00581722f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.925
cc_125 VPB N_A_762_107#_c_497_n 8.50551e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_762_107#_c_508_n 0.0207819f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=2.035
cc_127 VPB N_A_762_107#_c_509_n 0.0016742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_762_107#_c_498_n 0.00658622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_762_107#_c_511_n 0.0373665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_762_107#_c_512_n 4.79266e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_762_107#_c_513_n 0.0167636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_762_107#_c_500_n 0.00261149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_762_107#_c_502_n 0.00607421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_634_133#_M1005_g 0.0273298f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.475
cc_135 VPB N_A_634_133#_c_637_n 0.00942226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_634_133#_c_640_n 0.0100674f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_CLK_c_706_n 0.0210344f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.955
cc_138 VPB N_CLK_c_707_n 0.0188193f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.475
cc_139 VPB CLK 0.00591693f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_140 VPB N_CLK_c_705_n 0.0222106f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.925
cc_141 VPB N_A_1275_367#_M1001_g 0.0198811f $X=-0.19 $Y=1.655 $X2=0.312
+ $Y2=1.105
cc_142 VPB N_A_1275_367#_M1008_g 0.0187631f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_143 VPB N_A_1275_367#_M1013_g 0.0187631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_1275_367#_M1023_g 0.0264961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_1275_367#_c_767_n 0.00166092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_880_n 0.0103988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_881_n 0.0239601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_882_n 0.0118836f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.925
cc_149 VPB N_VPWR_c_883_n 0.0152644f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.12
cc_150 VPB N_VPWR_c_884_n 0.00495479f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=2.405
cc_151 VPB N_VPWR_c_885_n 0.0215328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_886_n 0.00236429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_887_n 0.00403269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_888_n 0.0130773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_889_n 0.0629959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_890_n 0.0292103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_891_n 0.0578293f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_892_n 0.0437554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_893_n 0.0152066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_894_n 0.0179513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_895_n 0.0034365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_896_n 0.0114188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_897_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_898_n 0.00349565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_899_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_879_n 0.0877722f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_134_70#_c_995_n 0.00211561f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.625
cc_168 VPB N_A_134_70#_c_998_n 0.0115886f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_169 VPB N_A_134_70#_c_999_n 0.0077251f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_170 VPB N_A_134_70#_c_1000_n 0.00294365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_134_70#_c_1001_n 0.0260029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_134_70#_c_1002_n 0.00192191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_134_70#_c_996_n 0.016955f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_174 VPB N_A_134_70#_c_1004_n 0.00431027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_GCLK_c_1074_n 9.46915e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_176 VPB N_GCLK_c_1070_n 0.00373964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_GCLK_c_1071_n 9.90345e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB GCLK 4.69342e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 N_SCE_M1022_g N_GATE_M1019_g 0.0486569f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_180 N_SCE_M1014_g N_GATE_M1012_g 0.00825767f $X=0.595 $Y=0.56 $X2=0 $Y2=0
cc_181 N_SCE_c_182_n N_GATE_c_215_n 0.0486569f $X=0.327 $Y=1.625 $X2=0 $Y2=0
cc_182 SCE N_GATE_c_215_n 0.00102444f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_183 N_SCE_c_184_n N_GATE_c_215_n 0.00806755f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_184 N_SCE_c_181_n N_GATE_c_217_n 0.00825767f $X=0.387 $Y=1.105 $X2=0 $Y2=0
cc_185 SCE N_VPWR_M1022_s 0.00297624f $X=0.155 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_186 N_SCE_M1022_g N_VPWR_c_881_n 0.00511835f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_187 SCE N_VPWR_c_881_n 0.0218679f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_188 N_SCE_M1022_g N_VPWR_c_890_n 0.00478016f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_189 N_SCE_M1022_g N_VPWR_c_879_n 0.008524f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_190 SCE N_VPWR_c_879_n 0.00386786f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_191 N_SCE_M1014_g N_A_134_70#_c_995_n 0.00457031f $X=0.595 $Y=0.56 $X2=0
+ $Y2=0
cc_192 N_SCE_c_182_n N_A_134_70#_c_995_n 0.00310251f $X=0.327 $Y=1.625 $X2=0
+ $Y2=0
cc_193 SCE N_A_134_70#_c_995_n 0.0607268f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_194 N_SCE_c_184_n N_A_134_70#_c_995_n 0.00348569f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_195 N_SCE_M1022_g N_A_134_70#_c_998_n 0.00324876f $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_196 SCE N_A_134_70#_c_998_n 0.0161137f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_197 N_SCE_M1022_g N_A_134_70#_c_1004_n 0.00126524f $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_198 SCE N_A_134_70#_c_1004_n 0.0101929f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_199 N_SCE_M1014_g N_VGND_c_1125_n 0.00928596f $X=0.595 $Y=0.56 $X2=0 $Y2=0
cc_200 N_SCE_c_181_n N_VGND_c_1125_n 0.00380198f $X=0.387 $Y=1.105 $X2=0 $Y2=0
cc_201 SCE N_VGND_c_1125_n 0.0205137f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_202 N_SCE_M1014_g N_VGND_c_1126_n 0.00428763f $X=0.595 $Y=0.56 $X2=0 $Y2=0
cc_203 N_SCE_M1014_g N_VGND_c_1143_n 0.00834303f $X=0.595 $Y=0.56 $X2=0 $Y2=0
cc_204 SCE N_VGND_c_1143_n 0.00556143f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_205 GATE N_A_252_361#_c_287_n 0.00611062f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_206 N_GATE_M1019_g N_A_252_361#_c_288_n 0.0313196f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_207 N_GATE_c_215_n N_A_252_361#_c_288_n 0.00360431f $X=1.15 $Y=1.445 $X2=0
+ $Y2=0
cc_208 N_GATE_c_218_n N_A_252_361#_c_288_n 0.00611062f $X=1.315 $Y=1.357 $X2=0
+ $Y2=0
cc_209 N_GATE_M1012_g N_A_252_361#_M1027_g 0.0131449f $X=1.06 $Y=0.56 $X2=0
+ $Y2=0
cc_210 GATE N_A_252_361#_M1027_g 0.0131671f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_211 N_GATE_c_217_n N_A_252_361#_M1027_g 0.013273f $X=1.15 $Y=1.09 $X2=0 $Y2=0
cc_212 N_GATE_c_218_n N_A_252_361#_M1027_g 7.98902e-19 $X=1.315 $Y=1.357 $X2=0
+ $Y2=0
cc_213 GATE N_A_252_361#_c_272_n 0.011602f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_214 N_GATE_c_215_n N_A_252_361#_c_273_n 0.013273f $X=1.15 $Y=1.445 $X2=0
+ $Y2=0
cc_215 GATE N_A_252_361#_c_273_n 0.00586843f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_216 N_GATE_c_215_n N_A_252_361#_c_274_n 0.00189696f $X=1.15 $Y=1.445 $X2=0
+ $Y2=0
cc_217 GATE N_A_252_361#_c_274_n 0.0220038f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_218 GATE N_A_252_361#_c_275_n 0.00845535f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_219 GATE N_A_252_361#_c_278_n 0.00470257f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_220 GATE N_A_252_361#_c_281_n 0.00213552f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_221 GATE N_A_335_70#_c_424_n 0.016583f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_222 GATE N_A_335_70#_c_425_n 0.0578055f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_223 N_GATE_M1012_g N_A_335_70#_c_426_n 3.48559e-19 $X=1.06 $Y=0.56 $X2=0
+ $Y2=0
cc_224 GATE N_A_335_70#_c_426_n 0.0216059f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_225 GATE N_A_335_70#_c_434_n 0.00133334f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_226 GATE N_A_335_70#_c_427_n 0.00176797f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_227 N_GATE_M1019_g N_VPWR_c_882_n 0.00151517f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_228 N_GATE_M1019_g N_VPWR_c_890_n 0.0030129f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_229 N_GATE_M1019_g N_VPWR_c_879_n 0.00394749f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_230 N_GATE_M1019_g N_A_134_70#_c_995_n 0.0094168f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_231 N_GATE_M1012_g N_A_134_70#_c_995_n 0.00936345f $X=1.06 $Y=0.56 $X2=0
+ $Y2=0
cc_232 N_GATE_c_215_n N_A_134_70#_c_995_n 0.00778453f $X=1.15 $Y=1.445 $X2=0
+ $Y2=0
cc_233 N_GATE_c_218_n N_A_134_70#_c_995_n 0.0682607f $X=1.315 $Y=1.357 $X2=0
+ $Y2=0
cc_234 N_GATE_M1019_g N_A_134_70#_c_998_n 0.0186933f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_235 N_GATE_c_215_n N_A_134_70#_c_999_n 2.34978e-19 $X=1.15 $Y=1.445 $X2=0
+ $Y2=0
cc_236 GATE N_A_134_70#_c_999_n 0.015044f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_237 N_GATE_c_218_n N_A_134_70#_c_999_n 0.0547947f $X=1.315 $Y=1.357 $X2=0
+ $Y2=0
cc_238 N_GATE_M1019_g N_A_134_70#_c_1004_n 0.00600965f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_239 N_GATE_c_215_n N_A_134_70#_c_1004_n 0.00640233f $X=1.15 $Y=1.445 $X2=0
+ $Y2=0
cc_240 N_GATE_c_218_n N_A_134_70#_c_1004_n 0.0139953f $X=1.315 $Y=1.357 $X2=0
+ $Y2=0
cc_241 N_GATE_M1012_g N_VGND_c_1125_n 5.40789e-19 $X=1.06 $Y=0.56 $X2=0 $Y2=0
cc_242 N_GATE_M1012_g N_VGND_c_1126_n 0.00478016f $X=1.06 $Y=0.56 $X2=0 $Y2=0
cc_243 N_GATE_M1012_g N_VGND_c_1127_n 0.00418155f $X=1.06 $Y=0.56 $X2=0 $Y2=0
cc_244 GATE N_VGND_c_1127_n 0.00920231f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_245 N_GATE_c_217_n N_VGND_c_1127_n 0.00372849f $X=1.15 $Y=1.09 $X2=0 $Y2=0
cc_246 N_GATE_c_218_n N_VGND_c_1127_n 0.0102124f $X=1.315 $Y=1.357 $X2=0 $Y2=0
cc_247 N_GATE_M1012_g N_VGND_c_1143_n 0.00945541f $X=1.06 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_252_361#_c_276_n N_A_335_70#_c_419_n 0.030465f $X=3.02 $Y=1.27 $X2=0
+ $Y2=0
cc_249 N_A_252_361#_c_289_n N_A_335_70#_M1020_g 0.0104164f $X=3.45 $Y=3.15 $X2=0
+ $Y2=0
cc_250 N_A_252_361#_M1025_g N_A_335_70#_M1020_g 0.0124191f $X=3.525 $Y=2.525
+ $X2=0 $Y2=0
cc_251 N_A_252_361#_M1025_g N_A_335_70#_c_421_n 0.00532637f $X=3.525 $Y=2.525
+ $X2=0 $Y2=0
cc_252 N_A_252_361#_c_277_n N_A_335_70#_M1016_g 0.0184335f $X=3.095 $Y=1.195
+ $X2=0 $Y2=0
cc_253 N_A_252_361#_c_280_n N_A_335_70#_M1016_g 0.00649445f $X=3.7 $Y=0.35 $X2=0
+ $Y2=0
cc_254 N_A_252_361#_c_284_n N_A_335_70#_M1016_g 0.00346756f $X=3.785 $Y=0.35
+ $X2=0 $Y2=0
cc_255 N_A_252_361#_c_277_n N_A_335_70#_c_424_n 0.00205835f $X=3.095 $Y=1.195
+ $X2=0 $Y2=0
cc_256 N_A_252_361#_c_278_n N_A_335_70#_c_424_n 9.22109e-19 $X=2.03 $Y=1.27
+ $X2=0 $Y2=0
cc_257 N_A_252_361#_c_280_n N_A_335_70#_c_424_n 0.0233726f $X=3.7 $Y=0.35 $X2=0
+ $Y2=0
cc_258 N_A_252_361#_c_281_n N_A_335_70#_c_424_n 0.0201666f $X=2.43 $Y=0.35 $X2=0
+ $Y2=0
cc_259 N_A_252_361#_c_274_n N_A_335_70#_c_425_n 0.00207743f $X=2.03 $Y=1.805
+ $X2=0 $Y2=0
cc_260 N_A_252_361#_c_276_n N_A_335_70#_c_425_n 0.00225155f $X=3.02 $Y=1.27
+ $X2=0 $Y2=0
cc_261 N_A_252_361#_c_294_n N_A_335_70#_c_425_n 0.00342394f $X=2.03 $Y=1.88
+ $X2=0 $Y2=0
cc_262 N_A_252_361#_c_279_n N_A_335_70#_c_425_n 0.00619503f $X=2.43 $Y=1.27
+ $X2=0 $Y2=0
cc_263 N_A_252_361#_c_281_n N_A_335_70#_c_425_n 0.0204781f $X=2.43 $Y=0.35 $X2=0
+ $Y2=0
cc_264 N_A_252_361#_M1027_g N_A_335_70#_c_426_n 0.00575819f $X=1.6 $Y=0.56 $X2=0
+ $Y2=0
cc_265 N_A_252_361#_c_272_n N_A_335_70#_c_426_n 0.0011181f $X=1.955 $Y=1.27
+ $X2=0 $Y2=0
cc_266 N_A_252_361#_c_280_n N_A_335_70#_c_426_n 0.00279077f $X=3.7 $Y=0.35 $X2=0
+ $Y2=0
cc_267 N_A_252_361#_c_281_n N_A_335_70#_c_426_n 0.00454373f $X=2.43 $Y=0.35
+ $X2=0 $Y2=0
cc_268 N_A_252_361#_c_292_n N_A_335_70#_c_434_n 0.0140096f $X=2.03 $Y=1.955
+ $X2=0 $Y2=0
cc_269 N_A_252_361#_c_275_n N_A_335_70#_c_434_n 0.00295973f $X=2.265 $Y=1.27
+ $X2=0 $Y2=0
cc_270 N_A_252_361#_c_274_n N_A_335_70#_c_427_n 0.0188921f $X=2.03 $Y=1.805
+ $X2=0 $Y2=0
cc_271 N_A_252_361#_c_279_n N_A_335_70#_c_427_n 0.0211693f $X=2.43 $Y=1.27 $X2=0
+ $Y2=0
cc_272 N_A_252_361#_c_282_n N_A_762_107#_M1004_d 0.00678554f $X=5.085 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_273 N_A_252_361#_c_282_n N_A_762_107#_M1009_g 0.00814169f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_274 N_A_252_361#_c_284_n N_A_762_107#_M1009_g 0.00489652f $X=3.785 $Y=0.35
+ $X2=0 $Y2=0
cc_275 N_A_252_361#_M1025_g N_A_762_107#_M1000_g 0.0401089f $X=3.525 $Y=2.525
+ $X2=0 $Y2=0
cc_276 N_A_252_361#_c_283_n N_A_762_107#_c_520_n 0.00929968f $X=5.17 $Y=1.93
+ $X2=0 $Y2=0
cc_277 N_A_252_361#_c_296_n N_A_762_107#_c_520_n 0.0175863f $X=5.255 $Y=2.035
+ $X2=0 $Y2=0
cc_278 N_A_252_361#_c_283_n N_A_762_107#_c_497_n 0.0421926f $X=5.17 $Y=1.93
+ $X2=0 $Y2=0
cc_279 N_A_252_361#_M1026_s N_A_762_107#_c_508_n 0.00281919f $X=5.435 $Y=1.835
+ $X2=0 $Y2=0
cc_280 N_A_252_361#_c_296_n N_A_762_107#_c_508_n 0.0143211f $X=5.255 $Y=2.035
+ $X2=0 $Y2=0
cc_281 N_A_252_361#_c_297_n N_A_762_107#_c_508_n 0.0309065f $X=5.56 $Y=2.035
+ $X2=0 $Y2=0
cc_282 N_A_252_361#_c_282_n N_A_762_107#_c_499_n 0.0219977f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_283 N_A_252_361#_c_283_n N_A_762_107#_c_499_n 0.0170646f $X=5.17 $Y=1.93
+ $X2=0 $Y2=0
cc_284 N_A_252_361#_c_283_n N_A_762_107#_c_512_n 0.0141629f $X=5.17 $Y=1.93
+ $X2=0 $Y2=0
cc_285 N_A_252_361#_c_282_n N_A_634_133#_c_635_n 0.0159414f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_286 N_A_252_361#_c_284_n N_A_634_133#_c_635_n 0.00408944f $X=3.785 $Y=0.35
+ $X2=0 $Y2=0
cc_287 N_A_252_361#_c_285_n N_A_634_133#_c_635_n 0.0100969f $X=5.265 $Y=0.445
+ $X2=0 $Y2=0
cc_288 N_A_252_361#_c_296_n N_A_634_133#_M1005_g 0.00109359f $X=5.255 $Y=2.035
+ $X2=0 $Y2=0
cc_289 N_A_252_361#_c_277_n N_A_634_133#_c_636_n 0.00150364f $X=3.095 $Y=1.195
+ $X2=0 $Y2=0
cc_290 N_A_252_361#_c_280_n N_A_634_133#_c_636_n 0.0131174f $X=3.7 $Y=0.35 $X2=0
+ $Y2=0
cc_291 N_A_252_361#_c_289_n N_A_634_133#_c_637_n 0.00320139f $X=3.45 $Y=3.15
+ $X2=0 $Y2=0
cc_292 N_A_252_361#_M1025_g N_A_634_133#_c_637_n 0.0107526f $X=3.525 $Y=2.525
+ $X2=0 $Y2=0
cc_293 N_A_252_361#_c_282_n N_A_634_133#_c_638_n 0.0178105f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_294 N_A_252_361#_c_284_n N_A_634_133#_c_638_n 0.00444167f $X=3.785 $Y=0.35
+ $X2=0 $Y2=0
cc_295 N_A_252_361#_c_276_n N_A_634_133#_c_639_n 0.00103365f $X=3.02 $Y=1.27
+ $X2=0 $Y2=0
cc_296 N_A_252_361#_c_282_n N_A_634_133#_c_640_n 0.00380096f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_297 N_A_252_361#_c_283_n N_A_634_133#_c_640_n 0.00199436f $X=5.17 $Y=1.93
+ $X2=0 $Y2=0
cc_298 N_A_252_361#_c_283_n N_CLK_M1017_g 0.0207f $X=5.17 $Y=1.93 $X2=0 $Y2=0
cc_299 N_A_252_361#_c_285_n N_CLK_M1017_g 0.00711079f $X=5.265 $Y=0.445 $X2=0
+ $Y2=0
cc_300 N_A_252_361#_c_283_n N_CLK_c_706_n 0.00323014f $X=5.17 $Y=1.93 $X2=0
+ $Y2=0
cc_301 N_A_252_361#_c_297_n N_CLK_c_706_n 0.00284228f $X=5.56 $Y=2.035 $X2=0
+ $Y2=0
cc_302 N_A_252_361#_c_283_n CLK 0.0421211f $X=5.17 $Y=1.93 $X2=0 $Y2=0
cc_303 N_A_252_361#_c_297_n CLK 0.0215698f $X=5.56 $Y=2.035 $X2=0 $Y2=0
cc_304 N_A_252_361#_c_283_n N_CLK_c_705_n 3.23951e-19 $X=5.17 $Y=1.93 $X2=0
+ $Y2=0
cc_305 N_A_252_361#_c_297_n N_CLK_c_705_n 0.00255472f $X=5.56 $Y=2.035 $X2=0
+ $Y2=0
cc_306 N_A_252_361#_c_286_n N_VPWR_c_882_n 0.00989746f $X=1.335 $Y=3.075 $X2=0
+ $Y2=0
cc_307 N_A_252_361#_c_289_n N_VPWR_c_882_n 0.0200829f $X=3.45 $Y=3.15 $X2=0
+ $Y2=0
cc_308 N_A_252_361#_c_292_n N_VPWR_c_882_n 0.00179401f $X=2.03 $Y=1.955 $X2=0
+ $Y2=0
cc_309 N_A_252_361#_M1025_g N_VPWR_c_883_n 0.0108077f $X=3.525 $Y=2.525 $X2=0
+ $Y2=0
cc_310 N_A_252_361#_M1025_g N_VPWR_c_914_n 0.00175164f $X=3.525 $Y=2.525 $X2=0
+ $Y2=0
cc_311 N_A_252_361#_c_290_n N_VPWR_c_890_n 0.00718072f $X=1.41 $Y=3.15 $X2=0
+ $Y2=0
cc_312 N_A_252_361#_c_289_n N_VPWR_c_891_n 0.0473923f $X=3.45 $Y=3.15 $X2=0
+ $Y2=0
cc_313 N_A_252_361#_c_289_n N_VPWR_c_879_n 0.061746f $X=3.45 $Y=3.15 $X2=0 $Y2=0
cc_314 N_A_252_361#_c_290_n N_VPWR_c_879_n 0.0112037f $X=1.41 $Y=3.15 $X2=0
+ $Y2=0
cc_315 N_A_252_361#_c_288_n N_A_134_70#_c_995_n 0.00108411f $X=1.41 $Y=1.88
+ $X2=0 $Y2=0
cc_316 N_A_252_361#_c_286_n N_A_134_70#_c_998_n 0.00974115f $X=1.335 $Y=3.075
+ $X2=0 $Y2=0
cc_317 N_A_252_361#_c_286_n N_A_134_70#_c_999_n 0.0143104f $X=1.335 $Y=3.075
+ $X2=0 $Y2=0
cc_318 N_A_252_361#_c_287_n N_A_134_70#_c_999_n 0.00851796f $X=1.955 $Y=1.88
+ $X2=0 $Y2=0
cc_319 N_A_252_361#_c_292_n N_A_134_70#_c_999_n 0.0080095f $X=2.03 $Y=1.955
+ $X2=0 $Y2=0
cc_320 N_A_252_361#_c_286_n N_A_134_70#_c_1000_n 0.00205036f $X=1.335 $Y=3.075
+ $X2=0 $Y2=0
cc_321 N_A_252_361#_c_292_n N_A_134_70#_c_1000_n 0.0226067f $X=2.03 $Y=1.955
+ $X2=0 $Y2=0
cc_322 N_A_252_361#_c_289_n N_A_134_70#_c_1001_n 0.022032f $X=3.45 $Y=3.15 $X2=0
+ $Y2=0
cc_323 N_A_252_361#_c_292_n N_A_134_70#_c_1001_n 0.00151465f $X=2.03 $Y=1.955
+ $X2=0 $Y2=0
cc_324 N_A_252_361#_M1025_g N_A_134_70#_c_1001_n 0.005862f $X=3.525 $Y=2.525
+ $X2=0 $Y2=0
cc_325 N_A_252_361#_c_289_n N_A_134_70#_c_1002_n 0.00274093f $X=3.45 $Y=3.15
+ $X2=0 $Y2=0
cc_326 N_A_252_361#_c_292_n N_A_134_70#_c_996_n 0.00333577f $X=2.03 $Y=1.955
+ $X2=0 $Y2=0
cc_327 N_A_252_361#_c_276_n N_A_134_70#_c_996_n 0.0125313f $X=3.02 $Y=1.27 $X2=0
+ $Y2=0
cc_328 N_A_252_361#_c_277_n N_A_134_70#_c_996_n 0.00117603f $X=3.095 $Y=1.195
+ $X2=0 $Y2=0
cc_329 N_A_252_361#_M1025_g N_A_134_70#_c_996_n 8.05738e-19 $X=3.525 $Y=2.525
+ $X2=0 $Y2=0
cc_330 N_A_252_361#_c_280_n N_A_134_70#_c_996_n 0.0114272f $X=3.7 $Y=0.35 $X2=0
+ $Y2=0
cc_331 N_A_252_361#_c_281_n N_A_134_70#_c_996_n 0.00176924f $X=2.43 $Y=0.35
+ $X2=0 $Y2=0
cc_332 N_A_252_361#_c_282_n N_VGND_M1009_d 0.0105055f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_333 N_A_252_361#_M1027_g N_VGND_c_1127_n 0.00364048f $X=1.6 $Y=0.56 $X2=0
+ $Y2=0
cc_334 N_A_252_361#_c_283_n N_VGND_c_1128_n 0.0158929f $X=5.17 $Y=1.93 $X2=0
+ $Y2=0
cc_335 N_A_252_361#_c_285_n N_VGND_c_1128_n 0.0298413f $X=5.265 $Y=0.445 $X2=0
+ $Y2=0
cc_336 N_A_252_361#_c_282_n N_VGND_c_1133_n 0.0149155f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_337 N_A_252_361#_c_285_n N_VGND_c_1133_n 0.0199466f $X=5.265 $Y=0.445 $X2=0
+ $Y2=0
cc_338 N_A_252_361#_M1027_g N_VGND_c_1135_n 0.00450978f $X=1.6 $Y=0.56 $X2=0
+ $Y2=0
cc_339 N_A_252_361#_c_280_n N_VGND_c_1135_n 0.0921784f $X=3.7 $Y=0.35 $X2=0
+ $Y2=0
cc_340 N_A_252_361#_c_281_n N_VGND_c_1135_n 0.00677996f $X=2.43 $Y=0.35 $X2=0
+ $Y2=0
cc_341 N_A_252_361#_c_282_n N_VGND_c_1135_n 0.00422649f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_342 N_A_252_361#_c_284_n N_VGND_c_1135_n 0.011658f $X=3.785 $Y=0.35 $X2=0
+ $Y2=0
cc_343 N_A_252_361#_c_282_n N_VGND_c_1140_n 0.0240258f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_344 N_A_252_361#_c_284_n N_VGND_c_1140_n 0.00761546f $X=3.785 $Y=0.35 $X2=0
+ $Y2=0
cc_345 N_A_252_361#_M1017_s N_VGND_c_1143_n 0.00216397f $X=5.14 $Y=0.235 $X2=0
+ $Y2=0
cc_346 N_A_252_361#_M1027_g N_VGND_c_1143_n 0.00869169f $X=1.6 $Y=0.56 $X2=0
+ $Y2=0
cc_347 N_A_252_361#_c_280_n N_VGND_c_1143_n 0.0525782f $X=3.7 $Y=0.35 $X2=0
+ $Y2=0
cc_348 N_A_252_361#_c_281_n N_VGND_c_1143_n 0.0101713f $X=2.43 $Y=0.35 $X2=0
+ $Y2=0
cc_349 N_A_252_361#_c_282_n N_VGND_c_1143_n 0.0286515f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_350 N_A_252_361#_c_284_n N_VGND_c_1143_n 0.00645941f $X=3.785 $Y=0.35 $X2=0
+ $Y2=0
cc_351 N_A_252_361#_c_285_n N_VGND_c_1143_n 0.0130351f $X=5.265 $Y=0.445 $X2=0
+ $Y2=0
cc_352 N_A_252_361#_c_284_n A_720_133# 0.00136037f $X=3.785 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_353 N_A_335_70#_M1020_g N_A_762_107#_M1009_g 0.00474587f $X=3.095 $Y=2.525
+ $X2=0 $Y2=0
cc_354 N_A_335_70#_c_421_n N_A_762_107#_M1009_g 0.0113266f $X=3.525 $Y=1.375
+ $X2=0 $Y2=0
cc_355 N_A_335_70#_M1016_g N_A_762_107#_M1009_g 0.0609898f $X=3.525 $Y=0.875
+ $X2=0 $Y2=0
cc_356 N_A_335_70#_c_421_n N_A_762_107#_c_498_n 7.77066e-19 $X=3.525 $Y=1.375
+ $X2=0 $Y2=0
cc_357 N_A_335_70#_M1016_g N_A_634_133#_c_636_n 0.0112748f $X=3.525 $Y=0.875
+ $X2=0 $Y2=0
cc_358 N_A_335_70#_M1020_g N_A_634_133#_c_637_n 0.00676697f $X=3.095 $Y=2.525
+ $X2=0 $Y2=0
cc_359 N_A_335_70#_c_420_n N_A_634_133#_c_637_n 0.0163086f $X=3.41 $Y=1.66 $X2=0
+ $Y2=0
cc_360 N_A_335_70#_c_421_n N_A_634_133#_c_637_n 0.00879229f $X=3.525 $Y=1.375
+ $X2=0 $Y2=0
cc_361 N_A_335_70#_c_421_n N_A_634_133#_c_638_n 0.0068014f $X=3.525 $Y=1.375
+ $X2=0 $Y2=0
cc_362 N_A_335_70#_M1016_g N_A_634_133#_c_638_n 0.00817362f $X=3.525 $Y=0.875
+ $X2=0 $Y2=0
cc_363 N_A_335_70#_c_421_n N_A_634_133#_c_639_n 0.00320147f $X=3.525 $Y=1.375
+ $X2=0 $Y2=0
cc_364 N_A_335_70#_M1016_g N_A_634_133#_c_639_n 0.00180242f $X=3.525 $Y=0.875
+ $X2=0 $Y2=0
cc_365 N_A_335_70#_M1020_g N_VPWR_c_879_n 9.39239e-19 $X=3.095 $Y=2.525 $X2=0
+ $Y2=0
cc_366 N_A_335_70#_c_425_n N_A_134_70#_c_999_n 0.00370107f $X=2.51 $Y=1.74 $X2=0
+ $Y2=0
cc_367 N_A_335_70#_c_434_n N_A_134_70#_c_999_n 0.00680086f $X=2.31 $Y=2.21 $X2=0
+ $Y2=0
cc_368 N_A_335_70#_c_434_n N_A_134_70#_c_1000_n 0.0418436f $X=2.31 $Y=2.21 $X2=0
+ $Y2=0
cc_369 N_A_335_70#_c_434_n N_A_134_70#_c_1001_n 0.0302168f $X=2.31 $Y=2.21 $X2=0
+ $Y2=0
cc_370 N_A_335_70#_c_419_n N_A_134_70#_c_996_n 0.0153888f $X=3.02 $Y=1.66 $X2=0
+ $Y2=0
cc_371 N_A_335_70#_M1020_g N_A_134_70#_c_996_n 0.017191f $X=3.095 $Y=2.525 $X2=0
+ $Y2=0
cc_372 N_A_335_70#_c_421_n N_A_134_70#_c_996_n 9.16865e-19 $X=3.525 $Y=1.375
+ $X2=0 $Y2=0
cc_373 N_A_335_70#_M1016_g N_A_134_70#_c_996_n 2.203e-19 $X=3.525 $Y=0.875 $X2=0
+ $Y2=0
cc_374 N_A_335_70#_c_424_n N_A_134_70#_c_996_n 0.00632692f $X=2.425 $Y=0.7 $X2=0
+ $Y2=0
cc_375 N_A_335_70#_c_425_n N_A_134_70#_c_996_n 0.148556f $X=2.51 $Y=1.74 $X2=0
+ $Y2=0
cc_376 N_A_335_70#_c_427_n N_A_134_70#_c_996_n 0.00164622f $X=2.675 $Y=1.74
+ $X2=0 $Y2=0
cc_377 N_A_335_70#_c_424_n N_VGND_c_1135_n 0.00542523f $X=2.425 $Y=0.7 $X2=0
+ $Y2=0
cc_378 N_A_335_70#_c_426_n N_VGND_c_1135_n 0.0106668f $X=1.815 $Y=0.56 $X2=0
+ $Y2=0
cc_379 N_A_335_70#_c_424_n N_VGND_c_1143_n 0.00853284f $X=2.425 $Y=0.7 $X2=0
+ $Y2=0
cc_380 N_A_335_70#_c_426_n N_VGND_c_1143_n 0.011421f $X=1.815 $Y=0.56 $X2=0
+ $Y2=0
cc_381 N_A_762_107#_M1009_g N_A_634_133#_c_635_n 0.0180232f $X=3.885 $Y=0.875
+ $X2=0 $Y2=0
cc_382 N_A_762_107#_c_497_n N_A_634_133#_c_635_n 0.00930102f $X=4.817 $Y=1.635
+ $X2=0 $Y2=0
cc_383 N_A_762_107#_c_499_n N_A_634_133#_c_635_n 0.00545514f $X=4.817 $Y=0.972
+ $X2=0 $Y2=0
cc_384 N_A_762_107#_M1009_g N_A_634_133#_M1005_g 0.00427078f $X=3.885 $Y=0.875
+ $X2=0 $Y2=0
cc_385 N_A_762_107#_c_506_n N_A_634_133#_M1005_g 0.0129653f $X=4.71 $Y=1.72
+ $X2=0 $Y2=0
cc_386 N_A_762_107#_c_520_n N_A_634_133#_M1005_g 0.0145374f $X=4.812 $Y=2.31
+ $X2=0 $Y2=0
cc_387 N_A_762_107#_c_497_n N_A_634_133#_M1005_g 0.00589026f $X=4.817 $Y=1.635
+ $X2=0 $Y2=0
cc_388 N_A_762_107#_c_498_n N_A_634_133#_M1005_g 7.623e-19 $X=3.972 $Y=1.72
+ $X2=0 $Y2=0
cc_389 N_A_762_107#_c_511_n N_A_634_133#_M1005_g 0.00608333f $X=3.975 $Y=1.93
+ $X2=0 $Y2=0
cc_390 N_A_762_107#_c_512_n N_A_634_133#_M1005_g 0.00352045f $X=4.812 $Y=1.72
+ $X2=0 $Y2=0
cc_391 N_A_762_107#_c_513_n N_A_634_133#_M1005_g 0.00704016f $X=4.875 $Y=2.425
+ $X2=0 $Y2=0
cc_392 N_A_762_107#_M1009_g N_A_634_133#_c_636_n 0.00271009f $X=3.885 $Y=0.875
+ $X2=0 $Y2=0
cc_393 N_A_762_107#_M1009_g N_A_634_133#_c_637_n 0.00259401f $X=3.885 $Y=0.875
+ $X2=0 $Y2=0
cc_394 N_A_762_107#_M1000_g N_A_634_133#_c_637_n 0.00372176f $X=3.885 $Y=2.525
+ $X2=0 $Y2=0
cc_395 N_A_762_107#_c_498_n N_A_634_133#_c_637_n 0.0235973f $X=3.972 $Y=1.72
+ $X2=0 $Y2=0
cc_396 N_A_762_107#_M1009_g N_A_634_133#_c_638_n 0.0131655f $X=3.885 $Y=0.875
+ $X2=0 $Y2=0
cc_397 N_A_762_107#_c_506_n N_A_634_133#_c_638_n 0.0293792f $X=4.71 $Y=1.72
+ $X2=0 $Y2=0
cc_398 N_A_762_107#_c_497_n N_A_634_133#_c_638_n 0.0161179f $X=4.817 $Y=1.635
+ $X2=0 $Y2=0
cc_399 N_A_762_107#_c_498_n N_A_634_133#_c_638_n 0.0263935f $X=3.972 $Y=1.72
+ $X2=0 $Y2=0
cc_400 N_A_762_107#_c_511_n N_A_634_133#_c_638_n 9.2809e-19 $X=3.975 $Y=1.93
+ $X2=0 $Y2=0
cc_401 N_A_762_107#_M1009_g N_A_634_133#_c_640_n 0.0182872f $X=3.885 $Y=0.875
+ $X2=0 $Y2=0
cc_402 N_A_762_107#_c_506_n N_A_634_133#_c_640_n 0.0100862f $X=4.71 $Y=1.72
+ $X2=0 $Y2=0
cc_403 N_A_762_107#_c_497_n N_A_634_133#_c_640_n 0.00648556f $X=4.817 $Y=1.635
+ $X2=0 $Y2=0
cc_404 N_A_762_107#_c_499_n N_A_634_133#_c_640_n 0.00334255f $X=4.817 $Y=0.972
+ $X2=0 $Y2=0
cc_405 N_A_762_107#_c_508_n N_CLK_c_706_n 0.0155071f $X=5.905 $Y=2.4 $X2=0 $Y2=0
cc_406 N_A_762_107#_c_509_n N_CLK_c_706_n 9.61374e-19 $X=6.35 $Y=1.93 $X2=0
+ $Y2=0
cc_407 N_A_762_107#_c_513_n N_CLK_c_706_n 0.0025612f $X=4.875 $Y=2.425 $X2=0
+ $Y2=0
cc_408 N_A_762_107#_c_495_n N_CLK_M1002_g 0.0737082f $X=6.365 $Y=1.185 $X2=0
+ $Y2=0
cc_409 N_A_762_107#_c_501_n N_CLK_M1002_g 0.00228216f $X=6.75 $Y=1.51 $X2=0
+ $Y2=0
cc_410 N_A_762_107#_c_508_n N_CLK_c_707_n 0.00186123f $X=5.905 $Y=2.4 $X2=0
+ $Y2=0
cc_411 N_A_762_107#_c_563_p N_CLK_c_707_n 0.00218198f $X=5.99 $Y=2.31 $X2=0
+ $Y2=0
cc_412 N_A_762_107#_c_564_p N_CLK_c_707_n 0.0140207f $X=6.265 $Y=2.015 $X2=0
+ $Y2=0
cc_413 N_A_762_107#_c_509_n N_CLK_c_707_n 0.0057478f $X=6.35 $Y=1.93 $X2=0 $Y2=0
cc_414 N_A_762_107#_c_496_n CLK 0.00323546f $X=6.75 $Y=1.335 $X2=0 $Y2=0
cc_415 N_A_762_107#_c_508_n CLK 0.00465993f $X=5.905 $Y=2.4 $X2=0 $Y2=0
cc_416 N_A_762_107#_c_564_p CLK 7.76592e-19 $X=6.265 $Y=2.015 $X2=0 $Y2=0
cc_417 N_A_762_107#_c_569_p CLK 0.0150037f $X=6.075 $Y=2.015 $X2=0 $Y2=0
cc_418 N_A_762_107#_c_509_n CLK 0.00620842f $X=6.35 $Y=1.93 $X2=0 $Y2=0
cc_419 N_A_762_107#_c_500_n CLK 0.0281951f $X=6.75 $Y=1.51 $X2=0 $Y2=0
cc_420 N_A_762_107#_c_501_n CLK 7.45196e-19 $X=6.75 $Y=1.51 $X2=0 $Y2=0
cc_421 N_A_762_107#_c_496_n N_CLK_c_705_n 0.00468597f $X=6.75 $Y=1.335 $X2=0
+ $Y2=0
cc_422 N_A_762_107#_M1007_g N_CLK_c_705_n 0.0360984f $X=6.73 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_762_107#_c_564_p N_CLK_c_705_n 0.00171045f $X=6.265 $Y=2.015 $X2=0
+ $Y2=0
cc_424 N_A_762_107#_c_569_p N_CLK_c_705_n 9.40339e-19 $X=6.075 $Y=2.015 $X2=0
+ $Y2=0
cc_425 N_A_762_107#_c_509_n N_CLK_c_705_n 0.00178854f $X=6.35 $Y=1.93 $X2=0
+ $Y2=0
cc_426 N_A_762_107#_c_500_n N_CLK_c_705_n 0.00592777f $X=6.75 $Y=1.51 $X2=0
+ $Y2=0
cc_427 N_A_762_107#_c_502_n N_CLK_c_705_n 0.00881075f $X=6.75 $Y=1.675 $X2=0
+ $Y2=0
cc_428 N_A_762_107#_c_564_p N_A_1275_367#_M1018_d 0.00152788f $X=6.265 $Y=2.015
+ $X2=0 $Y2=0
cc_429 N_A_762_107#_c_509_n N_A_1275_367#_M1018_d 8.73614e-19 $X=6.35 $Y=1.93
+ $X2=0 $Y2=0
cc_430 N_A_762_107#_M1007_g N_A_1275_367#_M1001_g 0.0315106f $X=6.73 $Y=2.465
+ $X2=0 $Y2=0
cc_431 N_A_762_107#_c_502_n N_A_1275_367#_M1001_g 0.00693383f $X=6.75 $Y=1.675
+ $X2=0 $Y2=0
cc_432 N_A_762_107#_c_495_n N_A_1275_367#_c_779_n 0.0142765f $X=6.365 $Y=1.185
+ $X2=0 $Y2=0
cc_433 N_A_762_107#_c_496_n N_A_1275_367#_c_765_n 0.00746469f $X=6.75 $Y=1.335
+ $X2=0 $Y2=0
cc_434 N_A_762_107#_c_500_n N_A_1275_367#_c_765_n 0.0127925f $X=6.75 $Y=1.51
+ $X2=0 $Y2=0
cc_435 N_A_762_107#_c_495_n N_A_1275_367#_c_766_n 0.00569877f $X=6.365 $Y=1.185
+ $X2=0 $Y2=0
cc_436 N_A_762_107#_c_496_n N_A_1275_367#_c_766_n 0.00667673f $X=6.75 $Y=1.335
+ $X2=0 $Y2=0
cc_437 N_A_762_107#_c_500_n N_A_1275_367#_c_766_n 0.023347f $X=6.75 $Y=1.51
+ $X2=0 $Y2=0
cc_438 N_A_762_107#_M1007_g N_A_1275_367#_c_785_n 0.00390528f $X=6.73 $Y=2.465
+ $X2=0 $Y2=0
cc_439 N_A_762_107#_c_500_n N_A_1275_367#_c_785_n 0.00327048f $X=6.75 $Y=1.51
+ $X2=0 $Y2=0
cc_440 N_A_762_107#_c_502_n N_A_1275_367#_c_785_n 0.00281217f $X=6.75 $Y=1.675
+ $X2=0 $Y2=0
cc_441 N_A_762_107#_M1007_g N_A_1275_367#_c_788_n 0.00468614f $X=6.73 $Y=2.465
+ $X2=0 $Y2=0
cc_442 N_A_762_107#_c_500_n N_A_1275_367#_c_788_n 0.0118852f $X=6.75 $Y=1.51
+ $X2=0 $Y2=0
cc_443 N_A_762_107#_M1007_g N_A_1275_367#_c_767_n 0.001674f $X=6.73 $Y=2.465
+ $X2=0 $Y2=0
cc_444 N_A_762_107#_c_509_n N_A_1275_367#_c_767_n 0.00529673f $X=6.35 $Y=1.93
+ $X2=0 $Y2=0
cc_445 N_A_762_107#_c_501_n N_A_1275_367#_c_767_n 0.002867f $X=6.75 $Y=1.51
+ $X2=0 $Y2=0
cc_446 N_A_762_107#_M1007_g N_A_1275_367#_c_793_n 0.0132505f $X=6.73 $Y=2.465
+ $X2=0 $Y2=0
cc_447 N_A_762_107#_c_500_n N_A_1275_367#_c_793_n 0.00581388f $X=6.75 $Y=1.51
+ $X2=0 $Y2=0
cc_448 N_A_762_107#_c_502_n N_A_1275_367#_c_793_n 4.7932e-19 $X=6.75 $Y=1.675
+ $X2=0 $Y2=0
cc_449 N_A_762_107#_M1007_g N_A_1275_367#_c_796_n 0.00694987f $X=6.73 $Y=2.465
+ $X2=0 $Y2=0
cc_450 N_A_762_107#_c_495_n N_A_1275_367#_c_768_n 4.36514e-19 $X=6.365 $Y=1.185
+ $X2=0 $Y2=0
cc_451 N_A_762_107#_c_496_n N_A_1275_367#_c_768_n 0.002867f $X=6.75 $Y=1.335
+ $X2=0 $Y2=0
cc_452 N_A_762_107#_c_500_n N_A_1275_367#_c_768_n 0.0258362f $X=6.75 $Y=1.51
+ $X2=0 $Y2=0
cc_453 N_A_762_107#_c_496_n N_A_1275_367#_c_769_n 0.0209471f $X=6.75 $Y=1.335
+ $X2=0 $Y2=0
cc_454 N_A_762_107#_c_506_n N_VPWR_M1000_d 0.00331815f $X=4.71 $Y=1.72 $X2=0
+ $Y2=0
cc_455 N_A_762_107#_c_508_n N_VPWR_M1026_d 0.00430824f $X=5.905 $Y=2.4 $X2=0
+ $Y2=0
cc_456 N_A_762_107#_c_563_p N_VPWR_M1026_d 0.00315349f $X=5.99 $Y=2.31 $X2=0
+ $Y2=0
cc_457 N_A_762_107#_c_564_p N_VPWR_M1026_d 0.00544015f $X=6.265 $Y=2.015 $X2=0
+ $Y2=0
cc_458 N_A_762_107#_c_569_p N_VPWR_M1026_d 0.00278484f $X=6.075 $Y=2.015 $X2=0
+ $Y2=0
cc_459 N_A_762_107#_M1000_g N_VPWR_c_883_n 0.00704662f $X=3.885 $Y=2.525 $X2=0
+ $Y2=0
cc_460 N_A_762_107#_M1000_g N_VPWR_c_926_n 0.00481866f $X=3.885 $Y=2.525 $X2=0
+ $Y2=0
cc_461 N_A_762_107#_c_506_n N_VPWR_c_926_n 0.0145773f $X=4.71 $Y=1.72 $X2=0
+ $Y2=0
cc_462 N_A_762_107#_c_498_n N_VPWR_c_926_n 0.00723326f $X=3.972 $Y=1.72 $X2=0
+ $Y2=0
cc_463 N_A_762_107#_c_511_n N_VPWR_c_926_n 8.91891e-19 $X=3.975 $Y=1.93 $X2=0
+ $Y2=0
cc_464 N_A_762_107#_c_508_n N_VPWR_c_884_n 0.00504147f $X=5.905 $Y=2.4 $X2=0
+ $Y2=0
cc_465 N_A_762_107#_M1007_g N_VPWR_c_885_n 0.00410857f $X=6.73 $Y=2.465 $X2=0
+ $Y2=0
cc_466 N_A_762_107#_M1007_g N_VPWR_c_886_n 0.011194f $X=6.73 $Y=2.465 $X2=0
+ $Y2=0
cc_467 N_A_762_107#_M1000_g N_VPWR_c_914_n 0.00515094f $X=3.885 $Y=2.525 $X2=0
+ $Y2=0
cc_468 N_A_762_107#_c_506_n N_VPWR_c_914_n 0.00696881f $X=4.71 $Y=1.72 $X2=0
+ $Y2=0
cc_469 N_A_762_107#_c_498_n N_VPWR_c_914_n 0.0102924f $X=3.972 $Y=1.72 $X2=0
+ $Y2=0
cc_470 N_A_762_107#_c_511_n N_VPWR_c_914_n 0.0011259f $X=3.975 $Y=1.93 $X2=0
+ $Y2=0
cc_471 N_A_762_107#_M1000_g N_VPWR_c_891_n 0.0035863f $X=3.885 $Y=2.525 $X2=0
+ $Y2=0
cc_472 N_A_762_107#_c_513_n N_VPWR_c_892_n 0.0108158f $X=4.875 $Y=2.425 $X2=0
+ $Y2=0
cc_473 N_A_762_107#_M1000_g N_VPWR_c_879_n 0.00401353f $X=3.885 $Y=2.525 $X2=0
+ $Y2=0
cc_474 N_A_762_107#_M1007_g N_VPWR_c_879_n 0.00658318f $X=6.73 $Y=2.465 $X2=0
+ $Y2=0
cc_475 N_A_762_107#_c_508_n N_VPWR_c_879_n 0.0328891f $X=5.905 $Y=2.4 $X2=0
+ $Y2=0
cc_476 N_A_762_107#_c_513_n N_VPWR_c_879_n 0.0115959f $X=4.875 $Y=2.425 $X2=0
+ $Y2=0
cc_477 N_A_762_107#_c_495_n N_VGND_c_1128_n 0.0033684f $X=6.365 $Y=1.185 $X2=0
+ $Y2=0
cc_478 N_A_762_107#_c_495_n N_VGND_c_1129_n 0.00370278f $X=6.365 $Y=1.185 $X2=0
+ $Y2=0
cc_479 N_A_762_107#_M1009_g N_VGND_c_1135_n 5.92631e-19 $X=3.885 $Y=0.875 $X2=0
+ $Y2=0
cc_480 N_A_762_107#_c_495_n N_VGND_c_1136_n 0.0054895f $X=6.365 $Y=1.185 $X2=0
+ $Y2=0
cc_481 N_A_762_107#_M1004_d N_VGND_c_1143_n 0.00288526f $X=4.585 $Y=0.245 $X2=0
+ $Y2=0
cc_482 N_A_762_107#_c_495_n N_VGND_c_1143_n 0.0111524f $X=6.365 $Y=1.185 $X2=0
+ $Y2=0
cc_483 N_A_634_133#_c_640_n N_CLK_c_705_n 0.00331872f $X=4.51 $Y=1.36 $X2=0
+ $Y2=0
cc_484 N_A_634_133#_M1005_g N_VPWR_c_883_n 0.0058712f $X=4.66 $Y=2.325 $X2=0
+ $Y2=0
cc_485 N_A_634_133#_c_637_n N_VPWR_c_914_n 0.011623f $X=3.31 $Y=2.53 $X2=0 $Y2=0
cc_486 N_A_634_133#_c_637_n N_VPWR_c_891_n 0.00463078f $X=3.31 $Y=2.53 $X2=0
+ $Y2=0
cc_487 N_A_634_133#_M1005_g N_VPWR_c_892_n 0.00431485f $X=4.66 $Y=2.325 $X2=0
+ $Y2=0
cc_488 N_A_634_133#_M1005_g N_VPWR_c_879_n 0.00544287f $X=4.66 $Y=2.325 $X2=0
+ $Y2=0
cc_489 N_A_634_133#_c_637_n N_VPWR_c_879_n 0.00767749f $X=3.31 $Y=2.53 $X2=0
+ $Y2=0
cc_490 N_A_634_133#_c_636_n N_A_134_70#_c_996_n 0.012934f $X=3.31 $Y=0.875 $X2=0
+ $Y2=0
cc_491 N_A_634_133#_c_637_n N_A_134_70#_c_996_n 0.0670572f $X=3.31 $Y=2.53 $X2=0
+ $Y2=0
cc_492 N_A_634_133#_c_639_n N_A_134_70#_c_996_n 0.0181924f $X=3.327 $Y=1.357
+ $X2=0 $Y2=0
cc_493 N_A_634_133#_c_635_n N_VGND_c_1133_n 0.00400062f $X=4.51 $Y=1.195 $X2=0
+ $Y2=0
cc_494 N_A_634_133#_c_635_n N_VGND_c_1140_n 0.00659856f $X=4.51 $Y=1.195 $X2=0
+ $Y2=0
cc_495 N_A_634_133#_c_635_n N_VGND_c_1143_n 0.00814141f $X=4.51 $Y=1.195 $X2=0
+ $Y2=0
cc_496 N_CLK_M1002_g N_A_1275_367#_c_779_n 0.00201647f $X=6.005 $Y=0.655 $X2=0
+ $Y2=0
cc_497 N_CLK_M1002_g N_A_1275_367#_c_766_n 7.94034e-19 $X=6.005 $Y=0.655 $X2=0
+ $Y2=0
cc_498 N_CLK_c_707_n N_VPWR_c_884_n 0.00460896f $X=6.3 $Y=1.725 $X2=0 $Y2=0
cc_499 N_CLK_c_707_n N_VPWR_c_885_n 0.00585385f $X=6.3 $Y=1.725 $X2=0 $Y2=0
cc_500 N_CLK_c_706_n N_VPWR_c_892_n 0.00312414f $X=5.775 $Y=1.725 $X2=0 $Y2=0
cc_501 N_CLK_c_706_n N_VPWR_c_879_n 0.00410284f $X=5.775 $Y=1.725 $X2=0 $Y2=0
cc_502 N_CLK_c_707_n N_VPWR_c_879_n 0.0120255f $X=6.3 $Y=1.725 $X2=0 $Y2=0
cc_503 N_CLK_M1017_g N_VGND_c_1128_n 0.011502f $X=5.48 $Y=0.445 $X2=0 $Y2=0
cc_504 N_CLK_M1002_g N_VGND_c_1128_n 0.020081f $X=6.005 $Y=0.655 $X2=0 $Y2=0
cc_505 CLK N_VGND_c_1128_n 0.0268314f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_506 N_CLK_c_705_n N_VGND_c_1128_n 0.00110431f $X=6.005 $Y=1.535 $X2=0 $Y2=0
cc_507 N_CLK_M1017_g N_VGND_c_1133_n 0.0054945f $X=5.48 $Y=0.445 $X2=0 $Y2=0
cc_508 N_CLK_M1002_g N_VGND_c_1136_n 0.00486043f $X=6.005 $Y=0.655 $X2=0 $Y2=0
cc_509 N_CLK_M1017_g N_VGND_c_1143_n 0.0116565f $X=5.48 $Y=0.445 $X2=0 $Y2=0
cc_510 N_CLK_M1002_g N_VGND_c_1143_n 0.00818711f $X=6.005 $Y=0.655 $X2=0 $Y2=0
cc_511 N_A_1275_367#_c_785_n N_VPWR_M1007_d 0.00864242f $X=7.025 $Y=1.93 $X2=0
+ $Y2=0
cc_512 N_A_1275_367#_c_793_n N_VPWR_c_885_n 0.0127325f $X=6.515 $Y=2.445 $X2=0
+ $Y2=0
cc_513 N_A_1275_367#_M1001_g N_VPWR_c_886_n 0.0138164f $X=7.265 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_1275_367#_M1008_g N_VPWR_c_886_n 6.82636e-19 $X=7.695 $Y=2.465 $X2=0
+ $Y2=0
cc_515 N_A_1275_367#_c_785_n N_VPWR_c_886_n 0.0155659f $X=7.025 $Y=1.93 $X2=0
+ $Y2=0
cc_516 N_A_1275_367#_c_796_n N_VPWR_c_886_n 0.0580378f $X=6.597 $Y=2.28 $X2=0
+ $Y2=0
cc_517 N_A_1275_367#_M1008_g N_VPWR_c_887_n 0.00189108f $X=7.695 $Y=2.465 $X2=0
+ $Y2=0
cc_518 N_A_1275_367#_M1013_g N_VPWR_c_887_n 0.00195866f $X=8.125 $Y=2.465 $X2=0
+ $Y2=0
cc_519 N_A_1275_367#_M1023_g N_VPWR_c_889_n 0.00658071f $X=8.555 $Y=2.465 $X2=0
+ $Y2=0
cc_520 N_A_1275_367#_c_769_n N_VPWR_c_889_n 5.89537e-19 $X=8.615 $Y=1.35 $X2=0
+ $Y2=0
cc_521 N_A_1275_367#_M1001_g N_VPWR_c_893_n 0.00564095f $X=7.265 $Y=2.465 $X2=0
+ $Y2=0
cc_522 N_A_1275_367#_M1008_g N_VPWR_c_893_n 0.00585385f $X=7.695 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A_1275_367#_M1013_g N_VPWR_c_894_n 0.00585385f $X=8.125 $Y=2.465 $X2=0
+ $Y2=0
cc_524 N_A_1275_367#_M1023_g N_VPWR_c_894_n 0.00585385f $X=8.555 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A_1275_367#_M1018_d N_VPWR_c_879_n 0.00363622f $X=6.375 $Y=1.835 $X2=0
+ $Y2=0
cc_526 N_A_1275_367#_M1001_g N_VPWR_c_879_n 0.00948291f $X=7.265 $Y=2.465 $X2=0
+ $Y2=0
cc_527 N_A_1275_367#_M1008_g N_VPWR_c_879_n 0.0105224f $X=7.695 $Y=2.465 $X2=0
+ $Y2=0
cc_528 N_A_1275_367#_M1013_g N_VPWR_c_879_n 0.0105224f $X=8.125 $Y=2.465 $X2=0
+ $Y2=0
cc_529 N_A_1275_367#_M1023_g N_VPWR_c_879_n 0.0109507f $X=8.555 $Y=2.465 $X2=0
+ $Y2=0
cc_530 N_A_1275_367#_c_793_n N_VPWR_c_879_n 0.0128642f $X=6.515 $Y=2.445 $X2=0
+ $Y2=0
cc_531 N_A_1275_367#_M1001_g N_GCLK_c_1074_n 0.00112786f $X=7.265 $Y=2.465 $X2=0
+ $Y2=0
cc_532 N_A_1275_367#_M1008_g N_GCLK_c_1074_n 0.00153102f $X=7.695 $Y=2.465 $X2=0
+ $Y2=0
cc_533 N_A_1275_367#_c_767_n N_GCLK_c_1074_n 0.00464507f $X=7.11 $Y=1.845 $X2=0
+ $Y2=0
cc_534 N_A_1275_367#_M1008_g N_GCLK_c_1070_n 0.0146866f $X=7.695 $Y=2.465 $X2=0
+ $Y2=0
cc_535 N_A_1275_367#_M1013_g N_GCLK_c_1070_n 0.0158565f $X=8.125 $Y=2.465 $X2=0
+ $Y2=0
cc_536 N_A_1275_367#_c_828_p N_GCLK_c_1070_n 0.0377215f $X=7.97 $Y=1.35 $X2=0
+ $Y2=0
cc_537 N_A_1275_367#_c_769_n N_GCLK_c_1070_n 0.00272261f $X=8.615 $Y=1.35 $X2=0
+ $Y2=0
cc_538 N_A_1275_367#_M1001_g N_GCLK_c_1071_n 0.001463f $X=7.265 $Y=2.465 $X2=0
+ $Y2=0
cc_539 N_A_1275_367#_c_767_n N_GCLK_c_1071_n 0.0137139f $X=7.11 $Y=1.845 $X2=0
+ $Y2=0
cc_540 N_A_1275_367#_c_828_p N_GCLK_c_1071_n 0.0202789f $X=7.97 $Y=1.35 $X2=0
+ $Y2=0
cc_541 N_A_1275_367#_c_769_n N_GCLK_c_1071_n 0.00282576f $X=8.615 $Y=1.35 $X2=0
+ $Y2=0
cc_542 N_A_1275_367#_c_760_n N_GCLK_c_1089_n 0.0097033f $X=7.755 $Y=1.185 $X2=0
+ $Y2=0
cc_543 N_A_1275_367#_c_762_n N_GCLK_c_1089_n 0.0112704f $X=8.185 $Y=1.185 $X2=0
+ $Y2=0
cc_544 N_A_1275_367#_c_828_p N_GCLK_c_1089_n 0.029905f $X=7.97 $Y=1.35 $X2=0
+ $Y2=0
cc_545 N_A_1275_367#_c_769_n N_GCLK_c_1089_n 0.00247845f $X=8.615 $Y=1.35 $X2=0
+ $Y2=0
cc_546 N_A_1275_367#_c_828_p N_GCLK_c_1093_n 0.014315f $X=7.97 $Y=1.35 $X2=0
+ $Y2=0
cc_547 N_A_1275_367#_c_769_n N_GCLK_c_1093_n 0.00256622f $X=8.615 $Y=1.35 $X2=0
+ $Y2=0
cc_548 N_A_1275_367#_M1023_g N_GCLK_c_1095_n 0.0022257f $X=8.555 $Y=2.465 $X2=0
+ $Y2=0
cc_549 N_A_1275_367#_M1013_g GCLK 0.00205756f $X=8.125 $Y=2.465 $X2=0 $Y2=0
cc_550 N_A_1275_367#_c_762_n GCLK 0.00271741f $X=8.185 $Y=1.185 $X2=0 $Y2=0
cc_551 N_A_1275_367#_M1023_g GCLK 0.00431939f $X=8.555 $Y=2.465 $X2=0 $Y2=0
cc_552 N_A_1275_367#_c_764_n GCLK 0.00250231f $X=8.615 $Y=1.185 $X2=0 $Y2=0
cc_553 N_A_1275_367#_c_828_p GCLK 0.0191053f $X=7.97 $Y=1.35 $X2=0 $Y2=0
cc_554 N_A_1275_367#_c_769_n GCLK 0.0308491f $X=8.615 $Y=1.35 $X2=0 $Y2=0
cc_555 N_A_1275_367#_M1023_g GCLK 0.0100493f $X=8.555 $Y=2.465 $X2=0 $Y2=0
cc_556 N_A_1275_367#_c_769_n GCLK 5.52796e-19 $X=8.615 $Y=1.35 $X2=0 $Y2=0
cc_557 N_A_1275_367#_M1013_g GCLK 0.00155543f $X=8.125 $Y=2.465 $X2=0 $Y2=0
cc_558 N_A_1275_367#_M1023_g GCLK 0.00829792f $X=8.555 $Y=2.465 $X2=0 $Y2=0
cc_559 N_A_1275_367#_c_765_n N_VGND_M1006_s 6.37779e-19 $X=7.025 $Y=1.085 $X2=0
+ $Y2=0
cc_560 N_A_1275_367#_c_768_n N_VGND_M1006_s 0.00209042f $X=7.11 $Y=1.085 $X2=0
+ $Y2=0
cc_561 N_A_1275_367#_c_779_n N_VGND_c_1128_n 0.0243674f $X=6.58 $Y=0.42 $X2=0
+ $Y2=0
cc_562 N_A_1275_367#_c_766_n N_VGND_c_1128_n 0.00158338f $X=6.685 $Y=1.085 $X2=0
+ $Y2=0
cc_563 N_A_1275_367#_c_758_n N_VGND_c_1129_n 0.0113101f $X=7.325 $Y=1.185 $X2=0
+ $Y2=0
cc_564 N_A_1275_367#_c_760_n N_VGND_c_1129_n 6.11179e-19 $X=7.755 $Y=1.185 $X2=0
+ $Y2=0
cc_565 N_A_1275_367#_c_779_n N_VGND_c_1129_n 0.0338805f $X=6.58 $Y=0.42 $X2=0
+ $Y2=0
cc_566 N_A_1275_367#_c_765_n N_VGND_c_1129_n 0.00657374f $X=7.025 $Y=1.085 $X2=0
+ $Y2=0
cc_567 N_A_1275_367#_c_828_p N_VGND_c_1129_n 0.00208825f $X=7.97 $Y=1.35 $X2=0
+ $Y2=0
cc_568 N_A_1275_367#_c_768_n N_VGND_c_1129_n 0.015057f $X=7.11 $Y=1.085 $X2=0
+ $Y2=0
cc_569 N_A_1275_367#_c_769_n N_VGND_c_1129_n 3.48823e-19 $X=8.615 $Y=1.35 $X2=0
+ $Y2=0
cc_570 N_A_1275_367#_c_758_n N_VGND_c_1130_n 5.68743e-19 $X=7.325 $Y=1.185 $X2=0
+ $Y2=0
cc_571 N_A_1275_367#_c_760_n N_VGND_c_1130_n 0.00989638f $X=7.755 $Y=1.185 $X2=0
+ $Y2=0
cc_572 N_A_1275_367#_c_762_n N_VGND_c_1130_n 0.0111959f $X=8.185 $Y=1.185 $X2=0
+ $Y2=0
cc_573 N_A_1275_367#_c_764_n N_VGND_c_1130_n 9.98661e-19 $X=8.615 $Y=1.185 $X2=0
+ $Y2=0
cc_574 N_A_1275_367#_c_762_n N_VGND_c_1132_n 0.0010228f $X=8.185 $Y=1.185 $X2=0
+ $Y2=0
cc_575 N_A_1275_367#_c_764_n N_VGND_c_1132_n 0.0180051f $X=8.615 $Y=1.185 $X2=0
+ $Y2=0
cc_576 N_A_1275_367#_c_779_n N_VGND_c_1136_n 0.0167743f $X=6.58 $Y=0.42 $X2=0
+ $Y2=0
cc_577 N_A_1275_367#_c_758_n N_VGND_c_1137_n 0.00486043f $X=7.325 $Y=1.185 $X2=0
+ $Y2=0
cc_578 N_A_1275_367#_c_760_n N_VGND_c_1137_n 0.00486043f $X=7.755 $Y=1.185 $X2=0
+ $Y2=0
cc_579 N_A_1275_367#_c_762_n N_VGND_c_1138_n 0.00486043f $X=8.185 $Y=1.185 $X2=0
+ $Y2=0
cc_580 N_A_1275_367#_c_764_n N_VGND_c_1138_n 0.00525069f $X=8.615 $Y=1.185 $X2=0
+ $Y2=0
cc_581 N_A_1275_367#_M1003_d N_VGND_c_1143_n 0.00288212f $X=6.44 $Y=0.235 $X2=0
+ $Y2=0
cc_582 N_A_1275_367#_c_758_n N_VGND_c_1143_n 0.00824727f $X=7.325 $Y=1.185 $X2=0
+ $Y2=0
cc_583 N_A_1275_367#_c_760_n N_VGND_c_1143_n 0.00455156f $X=7.755 $Y=1.185 $X2=0
+ $Y2=0
cc_584 N_A_1275_367#_c_762_n N_VGND_c_1143_n 0.00462979f $X=8.185 $Y=1.185 $X2=0
+ $Y2=0
cc_585 N_A_1275_367#_c_764_n N_VGND_c_1143_n 0.00897288f $X=8.615 $Y=1.185 $X2=0
+ $Y2=0
cc_586 N_A_1275_367#_c_779_n N_VGND_c_1143_n 0.0102362f $X=6.58 $Y=0.42 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_881_n N_A_134_70#_c_998_n 4.71234e-19 $X=0.26 $Y=2.825 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_882_n N_A_134_70#_c_998_n 0.0472087f $X=1.61 $Y=2.465 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_890_n N_A_134_70#_c_998_n 0.023158f $X=1.445 $Y=3.33 $X2=0 $Y2=0
cc_590 N_VPWR_c_879_n N_A_134_70#_c_998_n 0.0181539f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_591 N_VPWR_M1015_s N_A_134_70#_c_999_n 0.0094698f $X=1.485 $Y=2.065 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_882_n N_A_134_70#_c_999_n 0.0211114f $X=1.61 $Y=2.465 $X2=0
+ $Y2=0
cc_593 N_VPWR_M1015_s N_A_134_70#_c_1000_n 0.00650699f $X=1.485 $Y=2.065 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_882_n N_A_134_70#_c_1000_n 0.0443491f $X=1.61 $Y=2.465 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_891_n N_A_134_70#_c_1001_n 0.0633334f $X=3.935 $Y=3.33 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_879_n N_A_134_70#_c_1001_n 0.0326554f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_882_n N_A_134_70#_c_1002_n 0.016526f $X=1.61 $Y=2.465 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_891_n N_A_134_70#_c_1002_n 0.0115893f $X=3.935 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_VPWR_c_879_n N_A_134_70#_c_1002_n 0.00583135f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_879_n N_GCLK_M1001_d 0.00345315f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_601 N_VPWR_c_879_n N_GCLK_M1013_d 0.00281059f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_602 N_VPWR_c_893_n N_GCLK_c_1074_n 0.0144039f $X=7.78 $Y=3.33 $X2=0 $Y2=0
cc_603 N_VPWR_c_879_n N_GCLK_c_1074_n 0.00944728f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_604 N_VPWR_c_887_n N_GCLK_c_1070_n 0.0172048f $X=7.91 $Y=2.11 $X2=0 $Y2=0
cc_605 N_VPWR_c_894_n N_GCLK_c_1095_n 0.0140491f $X=8.675 $Y=3.33 $X2=0 $Y2=0
cc_606 N_VPWR_c_879_n N_GCLK_c_1095_n 0.0110907f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_607 N_VPWR_c_889_n GCLK 0.0248843f $X=8.77 $Y=1.98 $X2=0 $Y2=0
cc_608 N_A_134_70#_c_1068_p N_VGND_c_1126_n 0.00861831f $X=0.81 $Y=0.56 $X2=0
+ $Y2=0
cc_609 N_A_134_70#_c_1068_p N_VGND_c_1143_n 0.00955401f $X=0.81 $Y=0.56 $X2=0
+ $Y2=0
cc_610 N_GCLK_c_1089_n N_VGND_M1010_s 0.00328155f $X=8.305 $Y=0.93 $X2=0 $Y2=0
cc_611 N_GCLK_c_1089_n N_VGND_c_1130_n 0.016709f $X=8.305 $Y=0.93 $X2=0 $Y2=0
cc_612 GCLK N_VGND_c_1132_n 0.00334085f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_613 N_GCLK_c_1117_p N_VGND_c_1137_n 0.0124525f $X=7.54 $Y=0.42 $X2=0 $Y2=0
cc_614 GCLK N_VGND_c_1138_n 0.00607f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_615 N_GCLK_M1006_d N_VGND_c_1143_n 0.00408812f $X=7.4 $Y=0.235 $X2=0 $Y2=0
cc_616 N_GCLK_M1021_d N_VGND_c_1143_n 0.00398295f $X=8.26 $Y=0.235 $X2=0 $Y2=0
cc_617 N_GCLK_c_1117_p N_VGND_c_1143_n 0.00730901f $X=7.54 $Y=0.42 $X2=0 $Y2=0
cc_618 N_GCLK_c_1089_n N_VGND_c_1143_n 0.0108725f $X=8.305 $Y=0.93 $X2=0 $Y2=0
cc_619 GCLK N_VGND_c_1143_n 0.0069731f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_620 N_VGND_c_1143_n A_1216_47# 0.00899413f $X=8.88 $Y=0 $X2=-0.19 $Y2=-0.245
