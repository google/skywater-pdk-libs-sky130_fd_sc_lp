# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__xor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 1.180000 1.300000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.729000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.260000 1.180000 5.635000 1.515000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.220000 1.180000 7.535000 1.715000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.040000 0.265000 9.475000 1.125000 ;
        RECT 9.190000 1.125000 9.475000 3.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.090000  0.565000 2.000000 0.735000 ;
      RECT 0.090000  0.735000 0.605000 1.245000 ;
      RECT 0.090000  1.245000 0.260000 2.035000 ;
      RECT 0.090000  2.035000 0.440000 3.065000 ;
      RECT 0.440000  1.525000 0.790000 1.845000 ;
      RECT 0.440000  1.845000 1.650000 1.855000 ;
      RECT 0.620000  1.855000 1.650000 2.015000 ;
      RECT 0.620000  2.195000 0.950000 3.245000 ;
      RECT 0.785000  0.085000 1.115000 0.385000 ;
      RECT 1.440000  2.015000 1.770000 2.895000 ;
      RECT 1.440000  2.895000 4.060000 3.065000 ;
      RECT 1.480000  0.915000 1.650000 1.845000 ;
      RECT 1.830000  0.735000 2.000000 1.425000 ;
      RECT 1.830000  1.425000 2.825000 1.595000 ;
      RECT 1.985000  2.035000 2.315000 2.545000 ;
      RECT 1.985000  2.545000 3.710000 2.715000 ;
      RECT 2.180000  0.265000 3.360000 0.435000 ;
      RECT 2.180000  0.435000 2.430000 1.245000 ;
      RECT 2.495000  1.595000 2.825000 2.365000 ;
      RECT 2.655000  0.615000 3.010000 1.245000 ;
      RECT 2.655000  1.245000 2.825000 1.425000 ;
      RECT 3.005000  1.865000 3.360000 2.365000 ;
      RECT 3.190000  0.435000 3.360000 1.865000 ;
      RECT 3.540000  0.265000 5.430000 0.435000 ;
      RECT 3.540000  0.435000 3.710000 2.545000 ;
      RECT 3.890000  0.615000 5.080000 0.785000 ;
      RECT 3.890000  0.785000 4.060000 1.395000 ;
      RECT 3.890000  1.395000 4.160000 1.725000 ;
      RECT 3.890000  1.905000 4.570000 2.745000 ;
      RECT 3.890000  2.745000 4.060000 2.895000 ;
      RECT 4.240000  0.965000 4.570000 1.215000 ;
      RECT 4.400000  1.215000 4.570000 1.905000 ;
      RECT 4.830000  0.785000 5.080000 3.065000 ;
      RECT 5.260000  0.435000 5.430000 0.775000 ;
      RECT 5.260000  0.775000 6.340000 0.945000 ;
      RECT 5.260000  1.765000 5.590000 3.245000 ;
      RECT 5.610000  0.085000 5.860000 0.595000 ;
      RECT 5.885000  1.125000 6.690000 1.295000 ;
      RECT 5.885000  1.295000 6.135000 2.825000 ;
      RECT 6.090000  0.265000 7.885000 0.435000 ;
      RECT 6.090000  0.435000 6.340000 0.775000 ;
      RECT 6.315000  1.475000 6.645000 2.895000 ;
      RECT 6.315000  2.895000 8.235000 3.065000 ;
      RECT 6.520000  0.615000 7.470000 0.785000 ;
      RECT 6.520000  0.785000 6.690000 1.125000 ;
      RECT 6.825000  1.920000 7.155000 2.715000 ;
      RECT 6.870000  0.965000 7.040000 1.920000 ;
      RECT 7.220000  0.785000 7.470000 1.000000 ;
      RECT 7.335000  1.895000 7.885000 2.065000 ;
      RECT 7.335000  2.065000 7.715000 2.715000 ;
      RECT 7.715000  0.435000 7.885000 1.895000 ;
      RECT 7.895000  2.245000 8.235000 2.895000 ;
      RECT 8.065000  0.665000 8.315000 1.125000 ;
      RECT 8.065000  1.125000 8.235000 2.245000 ;
      RECT 8.440000  1.815000 8.610000 3.245000 ;
      RECT 8.530000  0.085000 8.860000 1.125000 ;
      RECT 8.680000  1.305000 9.010000 1.635000 ;
      RECT 8.790000  1.635000 9.010000 2.150000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  1.950000 3.205000 2.120000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  1.950000 6.085000 2.120000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  1.950000 7.045000 2.120000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  1.950000 8.965000 2.120000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
    LAYER met1 ;
      RECT 2.975000 1.920000 3.265000 1.965000 ;
      RECT 2.975000 1.965000 6.145000 2.105000 ;
      RECT 2.975000 2.105000 3.265000 2.150000 ;
      RECT 5.855000 1.920000 6.145000 1.965000 ;
      RECT 5.855000 2.105000 6.145000 2.150000 ;
      RECT 6.815000 1.920000 7.105000 1.965000 ;
      RECT 6.815000 1.965000 9.025000 2.105000 ;
      RECT 6.815000 2.105000 7.105000 2.150000 ;
      RECT 8.735000 1.920000 9.025000 1.965000 ;
      RECT 8.735000 2.105000 9.025000 2.150000 ;
  END
END sky130_fd_sc_lp__xor3_1
