* File: sky130_fd_sc_lp__dlxtp_lp.spice
* Created: Wed Sep  2 09:48:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxtp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dlxtp_lp  VNB VPB GATE D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1010 A_114_102# N_GATE_M1010_g N_A_27_102#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_GATE_M1001_g A_114_102# VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0441 PD=0.73 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1012 A_278_102# N_D_M1012_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0651 PD=0.63 PS=0.73 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1020 N_A_350_102#_M1020_d N_D_M1020_g A_278_102# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_584_47# N_A_27_102#_M1003_g N_A_463_491#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_27_102#_M1002_g A_584_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1029 AS=0.0504 PD=0.91 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1023 A_790_47# N_A_350_102#_M1023_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1029 PD=0.66 PS=0.91 NRD=18.564 NRS=59.988 M=1 R=2.8 SA=75001.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_824_491#_M1004_d N_A_463_491#_M1004_g A_790_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1009 A_982_47# N_A_27_102#_M1009_g N_A_824_491#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1027_407#_M1005_g A_982_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1106 AS=0.0504 PD=0.92 PS=0.66 NRD=1.428 NRS=18.564 M=1 R=2.8 SA=75002.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1025 A_1198_47# N_A_824_491#_M1025_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2212 PD=1.08 PS=1.84 NRD=9.276 NRS=36.42 M=1 R=5.6 SA=75001.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1026 N_A_1027_407#_M1026_d N_A_824_491#_M1026_g A_1198_47# VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1008 PD=2.25 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6
+ SA=75002.1 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 A_1474_53# N_A_1027_407#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1018 N_Q_M1018_d N_A_1027_407#_M1018_g A_1474_53# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 A_114_470# N_GATE_M1022_g N_A_27_102#_M1022_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_GATE_M1000_g A_114_470# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1019 A_278_470# N_D_M1019_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75001 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1017 N_A_350_102#_M1017_d N_D_M1017_g A_278_470# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1021 A_550_491# N_A_27_102#_M1021_g N_A_463_491#_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=19.9955 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1024 N_VPWR_M1024_d N_A_27_102#_M1024_g A_550_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1466 AS=0.0768 PD=1.12 PS=0.88 NRD=24.6053 NRS=19.9955 M=1 R=4.26667
+ SA=75000.6 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1014 A_746_491# N_A_350_102#_M1014_g N_VPWR_M1024_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1466 PD=0.88 PS=1.12 NRD=19.9955 NRS=24.6053 M=1 R=4.26667
+ SA=75001.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1016 N_A_824_491#_M1016_d N_A_27_102#_M1016_g A_746_491# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.138023 AS=0.0768 PD=1.24981 PS=0.88 NRD=0 NRS=19.9955 M=1
+ R=4.26667 SA=75001.6 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1008 A_933_535# N_A_463_491#_M1008_g N_A_824_491#_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0987 AS=0.0905774 PD=0.89 PS=0.820189 NRD=84.4145 NRS=53.9386 M=1
+ R=2.8 SA=75002.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_A_1027_407#_M1027_g A_933_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.121275 AS=0.0987 PD=0.9225 PS=0.89 NRD=143.042 NRS=84.4145 M=1 R=2.8
+ SA=75002.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1011 A_1204_367# N_A_824_491#_M1011_g N_VPWR_M1027_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.363825 PD=1.47 PS=2.7675 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_A_1027_407#_M1013_d N_A_824_491#_M1013_g A_1204_367# VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 A_1474_367# N_A_1027_407#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.3591 PD=1.47 PS=3.09 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1007 N_Q_M1007_d N_A_1027_407#_M1007_g A_1474_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.9271 P=20.81
*
.include "sky130_fd_sc_lp__dlxtp_lp.pxi.spice"
*
.ends
*
*
