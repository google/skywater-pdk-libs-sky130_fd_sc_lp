* File: sky130_fd_sc_lp__a2111oi_1.spice
* Created: Fri Aug 28 09:46:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a2111oi_1  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_D1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1659 AS=0.2478 PD=1.235 PS=2.27 NRD=8.568 NRS=1.428 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_C1_M1008_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2646 AS=0.1659 PD=1.47 PS=1.235 NRD=24.996 NRS=7.848 M=1 R=5.6 SA=75000.8
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.2646 PD=1.26 PS=1.47 NRD=9.276 NRS=24.996 M=1 R=5.6 SA=75001.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1006 A_499_47# N_A1_M1006_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.1764 PD=1.05 PS=1.26 NRD=7.14 NRS=10.704 M=1 R=5.6 SA=75002.1 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g A_499_47# VNB NSHORT L=0.15 W=0.84 AD=0.2352
+ AS=0.0882 PD=2.24 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75002.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1005 A_157_367# N_D1_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26 AD=0.2079
+ AS=0.6048 PD=1.59 PS=3.48 NRD=17.1981 NRS=33.6082 M=1 R=8.4 SA=75000.4
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1000 A_253_367# N_C1_M1000_g A_157_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.2079 PD=1.56 PS=1.59 NRD=14.8341 NRS=17.1981 M=1 R=8.4 SA=75000.9
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1004 N_A_343_367#_M1004_d N_B1_M1004_g A_253_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.189 PD=1.68 PS=1.56 NRD=11.7215 NRS=14.8341 M=1 R=8.4
+ SA=75001.3 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_343_367#_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2646 AS=0.2646 PD=1.68 PS=1.68 NRD=10.1455 NRS=10.1455 M=1 R=8.4
+ SA=75001.9 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1007 N_A_343_367#_M1007_d N_A2_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2646 PD=3.05 PS=1.68 NRD=0 NRS=11.7215 M=1 R=8.4
+ SA=75002.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a2111oi_1.pxi.spice"
*
.ends
*
*
