* File: sky130_fd_sc_lp__invlp_0.spice
* Created: Fri Aug 28 10:39:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__invlp_0.pex.spice"
.subckt sky130_fd_sc_lp__invlp_0  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 A_124_92# N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_124_92# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 A_124_468# N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1824 PD=0.88 PS=1.85 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g A_124_468# VPB PHIGHVT L=0.15 W=0.64 AD=0.1824
+ AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__invlp_0.pxi.spice"
*
.ends
*
*
