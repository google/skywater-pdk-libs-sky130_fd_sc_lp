* File: sky130_fd_sc_lp__a22o_4.pxi.spice
* Created: Wed Sep  2 09:22:40 2020
* 
x_PM_SKY130_FD_SC_LP__A22O_4%A_103_263# N_A_103_263#_M1001_d
+ N_A_103_263#_M1007_s N_A_103_263#_M1005_s N_A_103_263#_M1019_s
+ N_A_103_263#_M1000_g N_A_103_263#_M1008_g N_A_103_263#_M1003_g
+ N_A_103_263#_M1011_g N_A_103_263#_M1010_g N_A_103_263#_M1014_g
+ N_A_103_263#_M1021_g N_A_103_263#_M1022_g N_A_103_263#_c_122_n
+ N_A_103_263#_c_123_n N_A_103_263#_c_124_n N_A_103_263#_c_135_p
+ N_A_103_263#_c_236_p N_A_103_263#_c_137_p N_A_103_263#_c_132_n
+ N_A_103_263#_c_140_p N_A_103_263#_c_125_n N_A_103_263#_c_141_p
+ N_A_103_263#_c_142_p N_A_103_263#_c_173_p N_A_103_263#_c_126_n
+ PM_SKY130_FD_SC_LP__A22O_4%A_103_263#
x_PM_SKY130_FD_SC_LP__A22O_4%B2 N_B2_M1015_g N_B2_M1005_g N_B2_M1020_g
+ N_B2_M1023_g N_B2_c_272_n N_B2_c_273_n N_B2_c_274_n B2 N_B2_c_275_n
+ N_B2_c_276_n PM_SKY130_FD_SC_LP__A22O_4%B2
x_PM_SKY130_FD_SC_LP__A22O_4%B1 N_B1_c_358_n N_B1_M1001_g N_B1_M1004_g
+ N_B1_c_360_n N_B1_M1006_g N_B1_M1019_g B1 N_B1_c_362_n N_B1_c_363_n
+ PM_SKY130_FD_SC_LP__A22O_4%B1
x_PM_SKY130_FD_SC_LP__A22O_4%A2 N_A2_M1012_g N_A2_M1013_g N_A2_M1016_g
+ N_A2_M1017_g N_A2_c_412_n N_A2_c_413_n N_A2_c_414_n A2 A2 N_A2_c_416_n
+ N_A2_c_417_n PM_SKY130_FD_SC_LP__A22O_4%A2
x_PM_SKY130_FD_SC_LP__A22O_4%A1 N_A1_c_478_n N_A1_M1007_g N_A1_M1002_g
+ N_A1_c_480_n N_A1_M1018_g N_A1_M1009_g A1 A1 N_A1_c_483_n
+ PM_SKY130_FD_SC_LP__A22O_4%A1
x_PM_SKY130_FD_SC_LP__A22O_4%VPWR N_VPWR_M1000_s N_VPWR_M1008_s N_VPWR_M1014_s
+ N_VPWR_M1012_d N_VPWR_M1009_d N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n
+ N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n VPWR N_VPWR_c_539_n
+ N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_527_n N_VPWR_c_543_n N_VPWR_c_544_n
+ PM_SKY130_FD_SC_LP__A22O_4%VPWR
x_PM_SKY130_FD_SC_LP__A22O_4%X N_X_M1003_s N_X_M1021_s N_X_M1000_d N_X_M1011_d
+ N_X_c_628_n N_X_c_629_n N_X_c_622_n N_X_c_662_n N_X_c_630_n N_X_c_676_p
+ N_X_c_623_n N_X_c_667_n N_X_c_674_p N_X_c_631_n N_X_c_624_n X X X X X
+ PM_SKY130_FD_SC_LP__A22O_4%X
x_PM_SKY130_FD_SC_LP__A22O_4%A_549_367# N_A_549_367#_M1005_d
+ N_A_549_367#_M1004_d N_A_549_367#_M1023_d N_A_549_367#_M1002_s
+ N_A_549_367#_M1017_s N_A_549_367#_c_682_n N_A_549_367#_c_692_n
+ N_A_549_367#_c_683_n N_A_549_367#_c_694_n N_A_549_367#_c_695_n
+ N_A_549_367#_c_703_n N_A_549_367#_c_712_n N_A_549_367#_c_739_n
+ N_A_549_367#_c_716_n N_A_549_367#_c_684_n N_A_549_367#_c_685_n
+ N_A_549_367#_c_710_n N_A_549_367#_c_721_n
+ PM_SKY130_FD_SC_LP__A22O_4%A_549_367#
x_PM_SKY130_FD_SC_LP__A22O_4%VGND N_VGND_M1003_d N_VGND_M1010_d N_VGND_M1022_d
+ N_VGND_M1020_d N_VGND_M1016_s N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n
+ N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n N_VGND_c_753_n N_VGND_c_754_n
+ N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n VGND N_VGND_c_758_n
+ N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ PM_SKY130_FD_SC_LP__A22O_4%VGND
x_PM_SKY130_FD_SC_LP__A22O_4%A_632_47# N_A_632_47#_M1015_s N_A_632_47#_M1006_s
+ N_A_632_47#_c_839_n PM_SKY130_FD_SC_LP__A22O_4%A_632_47#
x_PM_SKY130_FD_SC_LP__A22O_4%A_1006_47# N_A_1006_47#_M1013_d
+ N_A_1006_47#_M1018_d N_A_1006_47#_c_849_n N_A_1006_47#_c_862_n
+ N_A_1006_47#_c_857_n N_A_1006_47#_c_852_n
+ PM_SKY130_FD_SC_LP__A22O_4%A_1006_47#
cc_1 VNB N_A_103_263#_M1000_g 5.40282e-19 $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.465
cc_2 VNB N_A_103_263#_M1008_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=2.465
cc_3 VNB N_A_103_263#_M1003_g 0.0284736f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.655
cc_4 VNB N_A_103_263#_M1011_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.7 $Y2=2.465
cc_5 VNB N_A_103_263#_M1010_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=0.655
cc_6 VNB N_A_103_263#_M1014_g 5.76584e-19 $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=2.465
cc_7 VNB N_A_103_263#_M1021_g 0.0214055f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=0.655
cc_8 VNB N_A_103_263#_M1022_g 0.0226113f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=0.655
cc_9 VNB N_A_103_263#_c_122_n 0.00185932f $X=-0.19 $Y=-0.245 $X2=2.63 $Y2=1.485
cc_10 VNB N_A_103_263#_c_123_n 0.00286818f $X=-0.19 $Y=-0.245 $X2=2.715
+ $Y2=1.385
cc_11 VNB N_A_103_263#_c_124_n 5.23438e-19 $X=-0.19 $Y=-0.245 $X2=2.715
+ $Y2=1.955
cc_12 VNB N_A_103_263#_c_125_n 0.001196f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=1.485
cc_13 VNB N_A_103_263#_c_126_n 0.142259f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=1.48
cc_14 VNB N_B2_M1015_g 0.0263308f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=1.835
cc_15 VNB N_B2_M1020_g 0.0271536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B2_c_272_n 0.00856386f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=1.645
cc_17 VNB N_B2_c_273_n 0.00211183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B2_c_274_n 0.0260103f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.315
cc_19 VNB N_B2_c_275_n 0.0264402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_c_276_n 0.00128133f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.315
cc_21 VNB N_B1_c_358_n 0.0164422f $X=-0.19 $Y=-0.245 $X2=3.59 $Y2=0.235
cc_22 VNB N_B1_M1004_g 0.00649785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_360_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_M1019_g 0.00649785f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.645
cc_25 VNB N_B1_c_362_n 0.00523549f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.315
cc_26 VNB N_B1_c_363_n 0.0339238f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.655
cc_27 VNB N_A2_M1013_g 0.0274163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_M1016_g 0.0243714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A2_M1017_g 0.00700975f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.465
cc_30 VNB N_A2_c_412_n 0.00856256f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=1.645
cc_31 VNB N_A2_c_413_n 0.00211183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_c_414_n 0.0260063f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.315
cc_33 VNB A2 0.00604556f $X=-0.19 $Y=-0.245 $X2=1.7 $Y2=1.645
cc_34 VNB N_A2_c_416_n 0.0562023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_417_n 0.0016291f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=0.655
cc_36 VNB N_A1_c_478_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=3.59 $Y2=0.235
cc_37 VNB N_A1_M1002_g 0.00649923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_c_480_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A1_M1009_g 0.00688674f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.645
cc_40 VNB A1 0.00873741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A1_c_483_n 0.0344458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_527_n 0.283096f $X=-0.19 $Y=-0.245 $X2=5.6 $Y2=0.865
cc_43 VNB N_X_c_622_n 0.0262098f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.465
cc_44 VNB N_X_c_623_n 0.00561181f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.315
cc_45 VNB N_X_c_624_n 0.00134924f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=0.655
cc_46 VNB X 0.0522398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB X 0.00999519f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.485
cc_48 VNB X 0.0257759f $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=2.045
cc_49 VNB N_VGND_c_747_n 0.0150313f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=2.465
cc_50 VNB N_VGND_c_748_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.655
cc_51 VNB N_VGND_c_749_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_750_n 0.00269342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_751_n 0.00295613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_752_n 0.0108094f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=2.465
cc_55 VNB N_VGND_c_753_n 0.0360654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_754_n 0.0284514f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=0.655
cc_57 VNB N_VGND_c_755_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_756_n 0.0130339f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=1.315
cc_59 VNB N_VGND_c_757_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=0.655
cc_60 VNB N_VGND_c_758_n 0.0350279f $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=1.48
cc_61 VNB N_VGND_c_759_n 0.0383148f $X=-0.19 $Y=-0.245 $X2=3.73 $Y2=0.925
cc_62 VNB N_VGND_c_760_n 0.00513098f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=1.485
cc_63 VNB N_VGND_c_761_n 0.00525267f $X=-0.19 $Y=-0.245 $X2=4.18 $Y2=2.045
cc_64 VNB N_VGND_c_762_n 0.350343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VPB N_A_103_263#_M1000_g 0.0229919f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.465
cc_66 VPB N_A_103_263#_M1008_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.27 $Y2=2.465
cc_67 VPB N_A_103_263#_M1011_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.7 $Y2=2.465
cc_68 VPB N_A_103_263#_M1014_g 0.024074f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.465
cc_69 VPB N_A_103_263#_c_124_n 0.00464921f $X=-0.19 $Y=1.655 $X2=2.715 $Y2=1.955
cc_70 VPB N_A_103_263#_c_132_n 0.00545378f $X=-0.19 $Y=1.655 $X2=2.8 $Y2=2.045
cc_71 VPB N_B2_M1005_g 0.0225593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B2_M1023_g 0.0188534f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.465
cc_73 VPB N_B2_c_272_n 0.00683345f $X=-0.19 $Y=1.655 $X2=1.27 $Y2=1.645
cc_74 VPB N_B2_c_273_n 0.00319037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_B2_c_274_n 0.00632477f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.315
cc_76 VPB N_B2_c_275_n 0.00643987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_B2_c_276_n 0.00223935f $X=-0.19 $Y=1.655 $X2=1.72 $Y2=1.315
cc_78 VPB N_B1_M1004_g 0.0188227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_B1_M1019_g 0.0188234f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.645
cc_80 VPB N_A2_M1012_g 0.0197033f $X=-0.19 $Y=1.655 $X2=3.16 $Y2=1.835
cc_81 VPB N_A2_M1017_g 0.0247639f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.465
cc_82 VPB N_A2_c_412_n 0.00727897f $X=-0.19 $Y=1.655 $X2=1.27 $Y2=1.645
cc_83 VPB N_A2_c_413_n 0.00264042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A2_c_414_n 0.00632078f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.315
cc_85 VPB N_A2_c_417_n 0.00831934f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=0.655
cc_86 VPB N_A1_M1002_g 0.0196793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A1_M1009_g 0.0186439f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.645
cc_88 VPB N_VPWR_c_528_n 0.0415892f $X=-0.19 $Y=1.655 $X2=1.27 $Y2=2.465
cc_89 VPB N_VPWR_c_529_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_530_n 0.00652077f $X=-0.19 $Y=1.655 $X2=1.72 $Y2=0.655
cc_91 VPB N_VPWR_c_531_n 0.00496764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_532_n 4.06069e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_533_n 0.0167814f $X=-0.19 $Y=1.655 $X2=2.58 $Y2=0.655
cc_94 VPB N_VPWR_c_534_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_535_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.485
cc_96 VPB N_VPWR_c_536_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.48
cc_97 VPB N_VPWR_c_537_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_538_n 0.00459045f $X=-0.19 $Y=1.655 $X2=2.38 $Y2=1.485
cc_99 VPB N_VPWR_c_539_n 0.0594369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_540_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_541_n 0.0153759f $X=-0.19 $Y=1.655 $X2=5.625 $Y2=0.865
cc_102 VPB N_VPWR_c_527_n 0.0698314f $X=-0.19 $Y=1.655 $X2=5.6 $Y2=0.865
cc_103 VPB N_VPWR_c_543_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_544_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.48
cc_105 VPB N_X_c_628_n 0.00955059f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.645
cc_106 VPB N_X_c_629_n 0.0183576f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.465
cc_107 VPB N_X_c_630_n 0.00578283f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=0.655
cc_108 VPB N_X_c_631_n 0.00144499f $X=-0.19 $Y=1.655 $X2=2.58 $Y2=0.655
cc_109 VPB X 0.00564837f $X=-0.19 $Y=1.655 $X2=3.205 $Y2=2.045
cc_110 VPB N_A_549_367#_c_682_n 0.00613424f $X=-0.19 $Y=1.655 $X2=1.27 $Y2=2.465
cc_111 VPB N_A_549_367#_c_683_n 0.00195038f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.315
cc_112 VPB N_A_549_367#_c_684_n 0.00778529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_549_367#_c_685_n 0.0360021f $X=-0.19 $Y=1.655 $X2=2.58 $Y2=0.655
cc_114 N_A_103_263#_M1022_g N_B2_M1015_g 0.0321433f $X=2.58 $Y=0.655 $X2=0 $Y2=0
cc_115 N_A_103_263#_c_123_n N_B2_M1015_g 0.004895f $X=2.715 $Y=1.385 $X2=0 $Y2=0
cc_116 N_A_103_263#_c_135_p N_B2_M1015_g 0.0145055f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_117 N_A_103_263#_c_124_n N_B2_M1005_g 0.00625793f $X=2.715 $Y=1.955 $X2=0
+ $Y2=0
cc_118 N_A_103_263#_c_137_p N_B2_M1005_g 0.0142117f $X=3.205 $Y=2.045 $X2=0
+ $Y2=0
cc_119 N_A_103_263#_c_135_p N_B2_M1020_g 0.0150564f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_120 N_A_103_263#_c_135_p N_B2_c_272_n 0.0106244f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_121 N_A_103_263#_c_140_p N_B2_c_272_n 0.0403667f $X=4.065 $Y=2.045 $X2=0
+ $Y2=0
cc_122 N_A_103_263#_c_141_p N_B2_c_272_n 0.0131052f $X=3.3 $Y=2.12 $X2=0 $Y2=0
cc_123 N_A_103_263#_c_142_p N_B2_c_272_n 0.0131052f $X=4.16 $Y=2.13 $X2=0 $Y2=0
cc_124 N_A_103_263#_c_135_p N_B2_c_273_n 0.0126184f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_125 N_A_103_263#_c_142_p N_B2_c_273_n 0.00334932f $X=4.16 $Y=2.13 $X2=0 $Y2=0
cc_126 N_A_103_263#_c_135_p N_B2_c_274_n 7.78777e-19 $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_127 N_A_103_263#_c_142_p N_B2_c_274_n 2.57653e-19 $X=4.16 $Y=2.13 $X2=0 $Y2=0
cc_128 N_A_103_263#_M1014_g N_B2_c_275_n 2.92549e-19 $X=2.13 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_103_263#_c_123_n N_B2_c_275_n 2.61744e-19 $X=2.715 $Y=1.385 $X2=0
+ $Y2=0
cc_130 N_A_103_263#_c_124_n N_B2_c_275_n 7.60368e-19 $X=2.715 $Y=1.955 $X2=0
+ $Y2=0
cc_131 N_A_103_263#_c_135_p N_B2_c_275_n 0.00231963f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_132 N_A_103_263#_c_137_p N_B2_c_275_n 0.00210436f $X=3.205 $Y=2.045 $X2=0
+ $Y2=0
cc_133 N_A_103_263#_c_125_n N_B2_c_275_n 0.0015198f $X=2.715 $Y=1.485 $X2=0
+ $Y2=0
cc_134 N_A_103_263#_c_126_n N_B2_c_275_n 0.0153025f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_135 N_A_103_263#_c_123_n N_B2_c_276_n 0.00291453f $X=2.715 $Y=1.385 $X2=0
+ $Y2=0
cc_136 N_A_103_263#_c_124_n N_B2_c_276_n 0.0151624f $X=2.715 $Y=1.955 $X2=0
+ $Y2=0
cc_137 N_A_103_263#_c_135_p N_B2_c_276_n 0.00969601f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_138 N_A_103_263#_c_137_p N_B2_c_276_n 0.0147026f $X=3.205 $Y=2.045 $X2=0
+ $Y2=0
cc_139 N_A_103_263#_c_125_n N_B2_c_276_n 0.0165945f $X=2.715 $Y=1.485 $X2=0
+ $Y2=0
cc_140 N_A_103_263#_c_141_p N_B2_c_276_n 0.0015941f $X=3.3 $Y=2.12 $X2=0 $Y2=0
cc_141 N_A_103_263#_c_126_n N_B2_c_276_n 2.65372e-19 $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_142 N_A_103_263#_c_135_p N_B1_c_358_n 0.00945519f $X=5.485 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_103_263#_c_140_p N_B1_M1004_g 0.0125125f $X=4.065 $Y=2.045 $X2=0
+ $Y2=0
cc_144 N_A_103_263#_c_135_p N_B1_c_360_n 0.00945519f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_145 N_A_103_263#_c_140_p N_B1_M1019_g 0.0125619f $X=4.065 $Y=2.045 $X2=0
+ $Y2=0
cc_146 N_A_103_263#_c_123_n N_B1_c_362_n 0.00495798f $X=2.715 $Y=1.385 $X2=0
+ $Y2=0
cc_147 N_A_103_263#_c_135_p N_B1_c_362_n 0.0390392f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_148 N_A_103_263#_c_135_p N_B1_c_363_n 0.00229312f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_149 N_A_103_263#_c_135_p N_A2_M1013_g 0.0149687f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_150 N_A_103_263#_c_135_p N_A2_c_412_n 0.00563137f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_151 N_A_103_263#_c_135_p N_A2_c_413_n 0.0126184f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_152 N_A_103_263#_c_135_p N_A2_c_414_n 7.73704e-19 $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_153 N_A_103_263#_c_135_p N_A1_c_478_n 0.0101105f $X=5.485 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_103_263#_c_173_p N_A1_c_480_n 0.00397842f $X=5.6 $Y=0.865 $X2=0 $Y2=0
cc_155 N_A_103_263#_c_135_p A1 0.0114899f $X=5.485 $Y=0.925 $X2=0 $Y2=0
cc_156 N_A_103_263#_c_173_p A1 0.0175737f $X=5.6 $Y=0.865 $X2=0 $Y2=0
cc_157 N_A_103_263#_c_173_p N_A1_c_483_n 0.0023208f $X=5.6 $Y=0.865 $X2=0 $Y2=0
cc_158 N_A_103_263#_M1000_g N_VPWR_c_528_n 0.0160937f $X=0.84 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_103_263#_M1008_g N_VPWR_c_528_n 7.27171e-19 $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_103_263#_M1000_g N_VPWR_c_529_n 7.27171e-19 $X=0.84 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_103_263#_M1008_g N_VPWR_c_529_n 0.0147004f $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_103_263#_M1011_g N_VPWR_c_529_n 0.0147923f $X=1.7 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_103_263#_M1014_g N_VPWR_c_529_n 7.43396e-19 $X=2.13 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_103_263#_M1014_g N_VPWR_c_530_n 0.00760043f $X=2.13 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_103_263#_c_122_n N_VPWR_c_530_n 0.0154892f $X=2.63 $Y=1.485 $X2=0
+ $Y2=0
cc_166 N_A_103_263#_c_124_n N_VPWR_c_530_n 0.0106157f $X=2.715 $Y=1.955 $X2=0
+ $Y2=0
cc_167 N_A_103_263#_c_132_n N_VPWR_c_530_n 0.015311f $X=2.8 $Y=2.045 $X2=0 $Y2=0
cc_168 N_A_103_263#_c_126_n N_VPWR_c_530_n 0.00632085f $X=2.58 $Y=1.48 $X2=0
+ $Y2=0
cc_169 N_A_103_263#_M1000_g N_VPWR_c_535_n 0.00486043f $X=0.84 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_103_263#_M1008_g N_VPWR_c_535_n 0.00486043f $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_103_263#_M1011_g N_VPWR_c_537_n 0.00486043f $X=1.7 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_103_263#_M1014_g N_VPWR_c_537_n 0.00585385f $X=2.13 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_103_263#_M1005_s N_VPWR_c_527_n 0.00225186f $X=3.16 $Y=1.835 $X2=0
+ $Y2=0
cc_174 N_A_103_263#_M1019_s N_VPWR_c_527_n 0.00225186f $X=4.02 $Y=1.835 $X2=0
+ $Y2=0
cc_175 N_A_103_263#_M1000_g N_VPWR_c_527_n 0.00824727f $X=0.84 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_103_263#_M1008_g N_VPWR_c_527_n 0.00824727f $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_103_263#_M1011_g N_VPWR_c_527_n 0.00824727f $X=1.7 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_103_263#_M1014_g N_VPWR_c_527_n 0.0118358f $X=2.13 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_103_263#_M1000_g N_X_c_628_n 0.015176f $X=0.84 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_103_263#_c_122_n N_X_c_628_n 0.0316102f $X=2.63 $Y=1.485 $X2=0 $Y2=0
cc_181 N_A_103_263#_c_126_n N_X_c_628_n 0.00601639f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_182 N_A_103_263#_M1003_g N_X_c_622_n 0.0159751f $X=1.29 $Y=0.655 $X2=0 $Y2=0
cc_183 N_A_103_263#_c_122_n N_X_c_622_n 0.064179f $X=2.63 $Y=1.485 $X2=0 $Y2=0
cc_184 N_A_103_263#_c_126_n N_X_c_622_n 0.0185359f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_185 N_A_103_263#_M1008_g N_X_c_630_n 0.0131657f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_103_263#_M1011_g N_X_c_630_n 0.0130597f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_103_263#_M1014_g N_X_c_630_n 0.00118751f $X=2.13 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_103_263#_c_122_n N_X_c_630_n 0.0660589f $X=2.63 $Y=1.485 $X2=0 $Y2=0
cc_189 N_A_103_263#_c_124_n N_X_c_630_n 0.00213368f $X=2.715 $Y=1.955 $X2=0
+ $Y2=0
cc_190 N_A_103_263#_c_126_n N_X_c_630_n 0.00508014f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_191 N_A_103_263#_M1010_g N_X_c_623_n 0.0138978f $X=1.72 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_103_263#_M1021_g N_X_c_623_n 0.0135203f $X=2.15 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A_103_263#_M1022_g N_X_c_623_n 0.00115089f $X=2.58 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A_103_263#_c_122_n N_X_c_623_n 0.0635201f $X=2.63 $Y=1.485 $X2=0 $Y2=0
cc_195 N_A_103_263#_c_123_n N_X_c_623_n 0.0122688f $X=2.715 $Y=1.385 $X2=0 $Y2=0
cc_196 N_A_103_263#_c_126_n N_X_c_623_n 0.00505664f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_197 N_A_103_263#_c_122_n N_X_c_631_n 0.0154948f $X=2.63 $Y=1.485 $X2=0 $Y2=0
cc_198 N_A_103_263#_c_126_n N_X_c_631_n 0.00250529f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_199 N_A_103_263#_c_122_n N_X_c_624_n 0.014679f $X=2.63 $Y=1.485 $X2=0 $Y2=0
cc_200 N_A_103_263#_c_126_n N_X_c_624_n 0.00262131f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_201 N_A_103_263#_M1000_g X 0.00299292f $X=0.84 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A_103_263#_c_122_n X 0.0162503f $X=2.63 $Y=1.485 $X2=0 $Y2=0
cc_203 N_A_103_263#_c_126_n X 0.00709498f $X=2.58 $Y=1.48 $X2=0 $Y2=0
cc_204 N_A_103_263#_c_124_n N_A_549_367#_M1005_d 0.00176694f $X=2.715 $Y=1.955
+ $X2=-0.19 $Y2=-0.245
cc_205 N_A_103_263#_c_137_p N_A_549_367#_M1005_d 0.00638241f $X=3.205 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_206 N_A_103_263#_c_132_n N_A_549_367#_M1005_d 0.00114555f $X=2.8 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_207 N_A_103_263#_c_140_p N_A_549_367#_M1004_d 0.00340214f $X=4.065 $Y=2.045
+ $X2=0 $Y2=0
cc_208 N_A_103_263#_c_137_p N_A_549_367#_c_682_n 0.0142524f $X=3.205 $Y=2.045
+ $X2=0 $Y2=0
cc_209 N_A_103_263#_c_132_n N_A_549_367#_c_682_n 0.00856802f $X=2.8 $Y=2.045
+ $X2=0 $Y2=0
cc_210 N_A_103_263#_M1005_s N_A_549_367#_c_692_n 0.00332344f $X=3.16 $Y=1.835
+ $X2=0 $Y2=0
cc_211 N_A_103_263#_c_141_p N_A_549_367#_c_692_n 0.0126348f $X=3.3 $Y=2.12 $X2=0
+ $Y2=0
cc_212 N_A_103_263#_c_140_p N_A_549_367#_c_694_n 0.0171443f $X=4.065 $Y=2.045
+ $X2=0 $Y2=0
cc_213 N_A_103_263#_M1019_s N_A_549_367#_c_695_n 0.00332344f $X=4.02 $Y=1.835
+ $X2=0 $Y2=0
cc_214 N_A_103_263#_c_142_p N_A_549_367#_c_695_n 0.0126348f $X=4.16 $Y=2.13
+ $X2=0 $Y2=0
cc_215 N_A_103_263#_c_123_n N_VGND_M1022_d 5.25086e-19 $X=2.715 $Y=1.385 $X2=0
+ $Y2=0
cc_216 N_A_103_263#_c_135_p N_VGND_M1022_d 0.00618567f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_217 N_A_103_263#_c_236_p N_VGND_M1022_d 9.59089e-19 $X=2.8 $Y=0.925 $X2=0
+ $Y2=0
cc_218 N_A_103_263#_c_135_p N_VGND_M1020_d 0.0140727f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_219 N_A_103_263#_M1003_g N_VGND_c_747_n 0.0120503f $X=1.29 $Y=0.655 $X2=0
+ $Y2=0
cc_220 N_A_103_263#_M1010_g N_VGND_c_747_n 6.25324e-19 $X=1.72 $Y=0.655 $X2=0
+ $Y2=0
cc_221 N_A_103_263#_M1003_g N_VGND_c_748_n 6.31957e-19 $X=1.29 $Y=0.655 $X2=0
+ $Y2=0
cc_222 N_A_103_263#_M1010_g N_VGND_c_748_n 0.0109915f $X=1.72 $Y=0.655 $X2=0
+ $Y2=0
cc_223 N_A_103_263#_M1021_g N_VGND_c_748_n 0.0108513f $X=2.15 $Y=0.655 $X2=0
+ $Y2=0
cc_224 N_A_103_263#_M1022_g N_VGND_c_748_n 6.22495e-19 $X=2.58 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_A_103_263#_M1021_g N_VGND_c_749_n 0.00486043f $X=2.15 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_A_103_263#_M1022_g N_VGND_c_749_n 0.00486043f $X=2.58 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_A_103_263#_M1021_g N_VGND_c_750_n 5.6167e-19 $X=2.15 $Y=0.655 $X2=0
+ $Y2=0
cc_228 N_A_103_263#_M1022_g N_VGND_c_750_n 0.00998635f $X=2.58 $Y=0.655 $X2=0
+ $Y2=0
cc_229 N_A_103_263#_c_135_p N_VGND_c_750_n 0.012288f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_230 N_A_103_263#_c_236_p N_VGND_c_750_n 0.00966429f $X=2.8 $Y=0.925 $X2=0
+ $Y2=0
cc_231 N_A_103_263#_c_135_p N_VGND_c_751_n 0.0217657f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_232 N_A_103_263#_M1003_g N_VGND_c_756_n 0.00486043f $X=1.29 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_103_263#_M1010_g N_VGND_c_756_n 0.00486043f $X=1.72 $Y=0.655 $X2=0
+ $Y2=0
cc_234 N_A_103_263#_M1001_d N_VGND_c_762_n 0.00225186f $X=3.59 $Y=0.235 $X2=0
+ $Y2=0
cc_235 N_A_103_263#_M1007_s N_VGND_c_762_n 0.00224381f $X=5.46 $Y=0.235 $X2=0
+ $Y2=0
cc_236 N_A_103_263#_M1003_g N_VGND_c_762_n 0.00824727f $X=1.29 $Y=0.655 $X2=0
+ $Y2=0
cc_237 N_A_103_263#_M1010_g N_VGND_c_762_n 0.00824727f $X=1.72 $Y=0.655 $X2=0
+ $Y2=0
cc_238 N_A_103_263#_M1021_g N_VGND_c_762_n 0.00824727f $X=2.15 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_103_263#_M1022_g N_VGND_c_762_n 0.00824727f $X=2.58 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_103_263#_c_135_p N_VGND_c_762_n 0.0217134f $X=5.485 $Y=0.925 $X2=0
+ $Y2=0
cc_241 N_A_103_263#_c_236_p N_VGND_c_762_n 6.25088e-19 $X=2.8 $Y=0.925 $X2=0
+ $Y2=0
cc_242 N_A_103_263#_c_135_p N_A_632_47#_M1015_s 0.00491906f $X=5.485 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_243 N_A_103_263#_c_135_p N_A_632_47#_M1006_s 0.00491906f $X=5.485 $Y=0.925
+ $X2=0 $Y2=0
cc_244 N_A_103_263#_M1001_d N_A_632_47#_c_839_n 0.00330393f $X=3.59 $Y=0.235
+ $X2=0 $Y2=0
cc_245 N_A_103_263#_c_135_p N_A_632_47#_c_839_n 0.0616608f $X=5.485 $Y=0.925
+ $X2=0 $Y2=0
cc_246 N_A_103_263#_c_135_p N_A_1006_47#_M1013_d 0.00491906f $X=5.485 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_247 N_A_103_263#_M1007_s N_A_1006_47#_c_849_n 0.00329373f $X=5.46 $Y=0.235
+ $X2=0 $Y2=0
cc_248 N_A_103_263#_c_135_p N_A_1006_47#_c_849_n 0.00613089f $X=5.485 $Y=0.925
+ $X2=0 $Y2=0
cc_249 N_A_103_263#_c_173_p N_A_1006_47#_c_849_n 0.0143265f $X=5.6 $Y=0.865
+ $X2=0 $Y2=0
cc_250 N_A_103_263#_c_135_p N_A_1006_47#_c_852_n 0.0148011f $X=5.485 $Y=0.925
+ $X2=0 $Y2=0
cc_251 N_B2_M1015_g N_B1_c_358_n 0.0398136f $X=3.085 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_252 N_B2_M1005_g N_B1_M1004_g 0.0345661f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_253 N_B2_c_272_n N_B1_M1004_g 0.00992403f $X=4.23 $Y=1.7 $X2=0 $Y2=0
cc_254 N_B2_M1020_g N_B1_c_360_n 0.0402416f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_255 N_B2_M1023_g N_B1_M1019_g 0.0352257f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B2_c_272_n N_B1_M1019_g 0.00992403f $X=4.23 $Y=1.7 $X2=0 $Y2=0
cc_257 N_B2_M1015_g N_B1_c_362_n 0.00153558f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_258 N_B2_M1020_g N_B1_c_362_n 8.93616e-19 $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_259 N_B2_c_272_n N_B1_c_362_n 0.0445968f $X=4.23 $Y=1.7 $X2=0 $Y2=0
cc_260 N_B2_c_273_n N_B1_c_362_n 0.00661829f $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_261 N_B2_c_274_n N_B1_c_362_n 3.44327e-19 $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_262 N_B2_c_275_n N_B1_c_362_n 5.97007e-19 $X=3.065 $Y=1.51 $X2=0 $Y2=0
cc_263 N_B2_c_276_n N_B1_c_362_n 0.00815143f $X=3.065 $Y=1.51 $X2=0 $Y2=0
cc_264 N_B2_c_272_n N_B1_c_363_n 0.00243542f $X=4.23 $Y=1.7 $X2=0 $Y2=0
cc_265 N_B2_c_273_n N_B1_c_363_n 0.00132951f $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_266 N_B2_c_274_n N_B1_c_363_n 0.0215098f $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_267 N_B2_c_275_n N_B1_c_363_n 0.0214703f $X=3.065 $Y=1.51 $X2=0 $Y2=0
cc_268 N_B2_c_276_n N_B1_c_363_n 0.00132315f $X=3.065 $Y=1.51 $X2=0 $Y2=0
cc_269 N_B2_M1023_g N_A2_M1012_g 0.0134965f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_270 N_B2_c_273_n N_A2_M1012_g 3.97293e-19 $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_271 N_B2_M1020_g N_A2_M1013_g 0.0295522f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_272 N_B2_M1023_g N_A2_c_413_n 3.33163e-19 $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_273 N_B2_c_273_n N_A2_c_413_n 0.0288097f $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_274 N_B2_c_274_n N_A2_c_413_n 0.00114936f $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_275 N_B2_c_273_n N_A2_c_414_n 0.00114936f $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_276 N_B2_c_274_n N_A2_c_414_n 0.0201104f $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_277 N_B2_M1005_g N_VPWR_c_530_n 0.00721315f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_278 N_B2_M1005_g N_VPWR_c_539_n 0.00357842f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_279 N_B2_M1023_g N_VPWR_c_539_n 0.00357877f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_280 N_B2_M1005_g N_VPWR_c_527_n 0.00667816f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_281 N_B2_M1023_g N_VPWR_c_527_n 0.00556347f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_282 N_B2_M1005_g N_A_549_367#_c_682_n 0.0102639f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_B2_M1005_g N_A_549_367#_c_692_n 0.010474f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_284 N_B2_M1005_g N_A_549_367#_c_683_n 5.89773e-19 $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_B2_M1005_g N_A_549_367#_c_694_n 5.565e-19 $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_286 N_B2_M1023_g N_A_549_367#_c_694_n 5.6475e-19 $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_B2_M1023_g N_A_549_367#_c_695_n 0.0121905f $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_B2_c_273_n N_A_549_367#_c_703_n 0.00646895f $X=4.395 $Y=1.51 $X2=0
+ $Y2=0
cc_289 N_B2_c_274_n N_A_549_367#_c_703_n 4.62566e-19 $X=4.395 $Y=1.51 $X2=0
+ $Y2=0
cc_290 N_B2_M1015_g N_VGND_c_750_n 0.00520786f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_291 N_B2_M1020_g N_VGND_c_751_n 0.00896145f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_292 N_B2_M1015_g N_VGND_c_758_n 0.00539883f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_293 N_B2_M1020_g N_VGND_c_758_n 0.00564095f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_294 N_B2_M1015_g N_VGND_c_762_n 0.0063753f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_295 N_B2_M1020_g N_VGND_c_762_n 0.00524073f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_296 N_B2_M1015_g N_A_632_47#_c_839_n 0.00524047f $X=3.085 $Y=0.655 $X2=0
+ $Y2=0
cc_297 N_B1_M1004_g N_VPWR_c_539_n 0.00357842f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_298 N_B1_M1019_g N_VPWR_c_539_n 0.00357842f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_299 N_B1_M1004_g N_VPWR_c_527_n 0.00537847f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_300 N_B1_M1019_g N_VPWR_c_527_n 0.00537847f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_301 N_B1_M1004_g N_A_549_367#_c_682_n 5.565e-19 $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_302 N_B1_M1004_g N_A_549_367#_c_692_n 0.010474f $X=3.515 $Y=2.465 $X2=0 $Y2=0
cc_303 N_B1_M1004_g N_A_549_367#_c_694_n 0.00919214f $X=3.515 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_B1_M1019_g N_A_549_367#_c_694_n 0.00930067f $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_B1_M1019_g N_A_549_367#_c_695_n 0.010474f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_306 N_B1_M1004_g N_A_549_367#_c_710_n 5.89773e-19 $X=3.515 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_B1_M1019_g N_A_549_367#_c_710_n 5.89773e-19 $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_B1_c_360_n N_VGND_c_751_n 0.00121f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_309 N_B1_c_358_n N_VGND_c_758_n 0.00357877f $X=3.515 $Y=1.185 $X2=0 $Y2=0
cc_310 N_B1_c_360_n N_VGND_c_758_n 0.00357877f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_311 N_B1_c_358_n N_VGND_c_762_n 0.00544922f $X=3.515 $Y=1.185 $X2=0 $Y2=0
cc_312 N_B1_c_360_n N_VGND_c_762_n 0.00544922f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_313 N_B1_c_358_n N_A_632_47#_c_839_n 0.0139064f $X=3.515 $Y=1.185 $X2=0 $Y2=0
cc_314 N_B1_c_360_n N_A_632_47#_c_839_n 0.0139464f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_315 N_A2_M1013_g N_A1_c_478_n 0.039855f $X=4.955 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_316 N_A2_M1012_g N_A1_M1002_g 0.0269976f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A2_c_412_n N_A1_M1002_g 0.0101589f $X=6.285 $Y=1.7 $X2=0 $Y2=0
cc_318 N_A2_M1016_g N_A1_c_480_n 0.0250392f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_319 N_A2_M1017_g N_A1_M1009_g 0.0250392f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A2_c_412_n N_A1_M1009_g 0.0103994f $X=6.285 $Y=1.7 $X2=0 $Y2=0
cc_321 N_A2_M1013_g A1 8.91727e-19 $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_322 N_A2_M1016_g A1 0.0024485f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_323 N_A2_c_412_n A1 0.0589249f $X=6.285 $Y=1.7 $X2=0 $Y2=0
cc_324 N_A2_c_413_n A1 0.0066674f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_325 N_A2_c_414_n A1 3.44095e-19 $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_326 A2 A1 0.0197311f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_327 N_A2_c_412_n N_A1_c_483_n 0.00243542f $X=6.285 $Y=1.7 $X2=0 $Y2=0
cc_328 N_A2_c_413_n N_A1_c_483_n 0.00132951f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_329 N_A2_c_414_n N_A1_c_483_n 0.0215098f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_330 A2 N_A1_c_483_n 0.0010715f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_331 N_A2_c_416_n N_A1_c_483_n 0.0250392f $X=6.45 $Y=1.375 $X2=0 $Y2=0
cc_332 N_A2_M1012_g N_VPWR_c_531_n 0.00429274f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A2_M1017_g N_VPWR_c_532_n 0.0161499f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_M1012_g N_VPWR_c_539_n 0.00585385f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_335 N_A2_M1017_g N_VPWR_c_541_n 0.00486043f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_336 N_A2_M1012_g N_VPWR_c_527_n 0.0109272f $X=4.875 $Y=2.465 $X2=0 $Y2=0
cc_337 N_A2_M1017_g N_VPWR_c_527_n 0.00917987f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_338 N_A2_M1012_g N_A_549_367#_c_712_n 0.0133686f $X=4.875 $Y=2.465 $X2=0
+ $Y2=0
cc_339 N_A2_c_412_n N_A_549_367#_c_712_n 0.0237845f $X=6.285 $Y=1.7 $X2=0 $Y2=0
cc_340 N_A2_c_413_n N_A_549_367#_c_712_n 0.0210724f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_341 N_A2_c_414_n N_A_549_367#_c_712_n 6.86827e-19 $X=4.935 $Y=1.51 $X2=0
+ $Y2=0
cc_342 N_A2_M1017_g N_A_549_367#_c_716_n 0.0121978f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_343 N_A2_c_412_n N_A_549_367#_c_716_n 0.036159f $X=6.285 $Y=1.7 $X2=0 $Y2=0
cc_344 N_A2_c_417_n N_A_549_367#_c_716_n 0.00460096f $X=6.45 $Y=1.615 $X2=0
+ $Y2=0
cc_345 N_A2_c_416_n N_A_549_367#_c_684_n 0.00111724f $X=6.45 $Y=1.375 $X2=0
+ $Y2=0
cc_346 N_A2_c_417_n N_A_549_367#_c_684_n 0.0222039f $X=6.45 $Y=1.615 $X2=0 $Y2=0
cc_347 N_A2_c_412_n N_A_549_367#_c_721_n 0.0161462f $X=6.285 $Y=1.7 $X2=0 $Y2=0
cc_348 N_A2_M1013_g N_VGND_c_751_n 0.00695429f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A2_M1016_g N_VGND_c_753_n 0.00677718f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_350 A2 N_VGND_c_753_n 0.0212353f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_351 N_A2_c_416_n N_VGND_c_753_n 0.00205546f $X=6.45 $Y=1.375 $X2=0 $Y2=0
cc_352 N_A2_M1013_g N_VGND_c_759_n 0.00547467f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_353 N_A2_M1016_g N_VGND_c_759_n 0.00585385f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_354 N_A2_M1013_g N_VGND_c_762_n 0.00670468f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_355 N_A2_M1016_g N_VGND_c_762_n 0.011494f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_356 N_A2_M1013_g N_A_1006_47#_c_852_n 0.00559844f $X=4.955 $Y=0.655 $X2=0
+ $Y2=0
cc_357 N_A1_M1002_g N_VPWR_c_531_n 0.0027519f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A1_M1002_g N_VPWR_c_532_n 6.86814e-19 $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_359 N_A1_M1009_g N_VPWR_c_532_n 0.014371f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_360 N_A1_M1002_g N_VPWR_c_540_n 0.00585385f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A1_M1009_g N_VPWR_c_540_n 0.00486043f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A1_M1002_g N_VPWR_c_527_n 0.0107422f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A1_M1009_g N_VPWR_c_527_n 0.00824727f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A1_M1002_g N_A_549_367#_c_712_n 0.0133747f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A1_M1009_g N_A_549_367#_c_716_n 0.0122129f $X=5.815 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_A1_c_478_n N_VGND_c_759_n 0.00357877f $X=5.385 $Y=1.185 $X2=0 $Y2=0
cc_367 N_A1_c_480_n N_VGND_c_759_n 0.00357877f $X=5.815 $Y=1.185 $X2=0 $Y2=0
cc_368 N_A1_c_478_n N_VGND_c_762_n 0.00544922f $X=5.385 $Y=1.185 $X2=0 $Y2=0
cc_369 N_A1_c_480_n N_VGND_c_762_n 0.00537654f $X=5.815 $Y=1.185 $X2=0 $Y2=0
cc_370 N_A1_c_478_n N_A_1006_47#_c_849_n 0.010814f $X=5.385 $Y=1.185 $X2=0 $Y2=0
cc_371 N_A1_c_480_n N_A_1006_47#_c_849_n 0.0124008f $X=5.815 $Y=1.185 $X2=0
+ $Y2=0
cc_372 A1 N_A_1006_47#_c_849_n 0.00358314f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_373 A1 N_A_1006_47#_c_857_n 0.0146042f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_374 N_A1_c_478_n N_A_1006_47#_c_852_n 0.00263296f $X=5.385 $Y=1.185 $X2=0
+ $Y2=0
cc_375 N_A1_c_480_n N_A_1006_47#_c_852_n 3.49705e-19 $X=5.815 $Y=1.185 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_527_n N_X_M1000_d 0.00536646f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPWR_c_527_n N_X_M1011_d 0.00397496f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_378 N_VPWR_M1000_s N_X_c_628_n 0.00262981f $X=0.5 $Y=1.835 $X2=0 $Y2=0
cc_379 N_VPWR_c_528_n N_X_c_628_n 0.0220026f $X=0.625 $Y=2.18 $X2=0 $Y2=0
cc_380 N_VPWR_c_535_n N_X_c_662_n 0.0124525f $X=1.32 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_527_n N_X_c_662_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_382 N_VPWR_M1008_s N_X_c_630_n 0.00176461f $X=1.345 $Y=1.835 $X2=0 $Y2=0
cc_383 N_VPWR_c_529_n N_X_c_630_n 0.0170777f $X=1.485 $Y=2.18 $X2=0 $Y2=0
cc_384 N_VPWR_c_530_n N_X_c_630_n 0.00164217f $X=2.345 $Y=1.98 $X2=0 $Y2=0
cc_385 N_VPWR_c_537_n N_X_c_667_n 0.0138717f $X=2.22 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_c_527_n N_X_c_667_n 0.00886411f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_387 N_VPWR_c_527_n N_A_549_367#_M1005_d 0.00215158f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_388 N_VPWR_c_527_n N_A_549_367#_M1004_d 0.00223559f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_527_n N_A_549_367#_M1023_d 0.00276635f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_527_n N_A_549_367#_M1002_s 0.00397496f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_527_n N_A_549_367#_M1017_s 0.00371702f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_530_n N_A_549_367#_c_682_n 0.036855f $X=2.345 $Y=1.98 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_539_n N_A_549_367#_c_692_n 0.0298674f $X=4.965 $Y=3.33 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_527_n N_A_549_367#_c_692_n 0.0187823f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_530_n N_A_549_367#_c_683_n 0.0111191f $X=2.345 $Y=1.98 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_539_n N_A_549_367#_c_683_n 0.0211865f $X=4.965 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_527_n N_A_549_367#_c_683_n 0.0126421f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_539_n N_A_549_367#_c_695_n 0.0518631f $X=4.965 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_527_n N_A_549_367#_c_695_n 0.0329308f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_M1012_d N_A_549_367#_c_712_n 0.00504637f $X=4.95 $Y=1.835 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_531_n N_A_549_367#_c_712_n 0.0200142f $X=5.13 $Y=2.38 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_540_n N_A_549_367#_c_739_n 0.0138717f $X=5.865 $Y=3.33 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_527_n N_A_549_367#_c_739_n 0.00886411f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_M1009_d N_A_549_367#_c_716_n 0.00353353f $X=5.89 $Y=1.835 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_532_n N_A_549_367#_c_716_n 0.0170777f $X=6.03 $Y=2.38 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_541_n N_A_549_367#_c_685_n 0.0178111f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_527_n N_A_549_367#_c_685_n 0.0100304f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_539_n N_A_549_367#_c_710_n 0.01906f $X=4.965 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_c_527_n N_A_549_367#_c_710_n 0.0124545f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_X_c_622_n N_VGND_M1003_d 0.00234752f $X=1.41 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_411 N_X_c_623_n N_VGND_M1010_d 0.00180746f $X=2.27 $Y=1.13 $X2=0 $Y2=0
cc_412 N_X_c_622_n N_VGND_c_747_n 0.0220025f $X=1.41 $Y=1.13 $X2=0 $Y2=0
cc_413 X N_VGND_c_747_n 0.0221568f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_414 N_X_c_623_n N_VGND_c_748_n 0.0163515f $X=2.27 $Y=1.13 $X2=0 $Y2=0
cc_415 N_X_c_674_p N_VGND_c_749_n 0.0124525f $X=2.365 $Y=0.42 $X2=0 $Y2=0
cc_416 X N_VGND_c_754_n 0.0160151f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_417 N_X_c_676_p N_VGND_c_756_n 0.0120977f $X=1.505 $Y=0.42 $X2=0 $Y2=0
cc_418 N_X_M1003_s N_VGND_c_762_n 0.00571434f $X=1.365 $Y=0.235 $X2=0 $Y2=0
cc_419 N_X_M1021_s N_VGND_c_762_n 0.00536646f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_420 N_X_c_676_p N_VGND_c_762_n 0.00691495f $X=1.505 $Y=0.42 $X2=0 $Y2=0
cc_421 N_X_c_674_p N_VGND_c_762_n 0.00730901f $X=2.365 $Y=0.42 $X2=0 $Y2=0
cc_422 X N_VGND_c_762_n 0.0121058f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_423 N_VGND_c_762_n N_A_632_47#_M1015_s 0.00225186f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_424 N_VGND_c_762_n N_A_632_47#_M1006_s 0.00241018f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_758_n N_A_632_47#_c_839_n 0.0661207f $X=4.445 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_762_n N_A_632_47#_c_839_n 0.0423718f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_762_n N_A_1006_47#_M1013_d 0.00225186f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_428 N_VGND_c_762_n N_A_1006_47#_M1018_d 0.00220345f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_759_n N_A_1006_47#_c_862_n 0.0139427f $X=6.335 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_762_n N_A_1006_47#_c_862_n 0.00894187f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_751_n N_A_1006_47#_c_852_n 0.0251888f $X=4.61 $Y=0.485 $X2=0
+ $Y2=0
cc_432 N_VGND_c_759_n N_A_1006_47#_c_852_n 0.0522841f $X=6.335 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_c_762_n N_A_1006_47#_c_852_n 0.0338756f $X=6.48 $Y=0 $X2=0 $Y2=0
