* NGSPICE file created from sky130_fd_sc_lp__a21boi_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21boi_m A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR A1 a_306_395# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1001 VGND A2 a_310_47# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.827e+11p ps=1.71e+06u
M1002 VGND B1_N a_27_535# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 Y a_27_535# VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1004 a_306_395# a_27_535# Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VPWR B1_N a_27_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 a_306_395# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_310_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

