# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o2bb2ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.905000 1.210000 6.565000 1.425000 ;
        RECT 5.905000 1.425000 7.935000 1.595000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.170000 8.975000 1.425000 ;
        RECT 8.285000 1.425000 9.635000 1.595000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.405000 1.425000 1.415000 1.645000 ;
        RECT 1.055000 1.645000 1.415000 1.950000 ;
        RECT 1.055000 1.950000 3.810000 2.130000 ;
        RECT 3.480000 1.425000 3.810000 1.950000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 1.425000 3.205000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.965600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 2.300000 4.405000 2.630000 ;
        RECT 3.995000 1.075000 5.515000 1.245000 ;
        RECT 3.995000 1.245000 4.165000 1.775000 ;
        RECT 3.995000 1.775000 5.265000 1.945000 ;
        RECT 3.995000 1.945000 4.405000 2.300000 ;
        RECT 4.165000 0.605000 4.495000 1.075000 ;
        RECT 4.215000 2.630000 4.405000 3.075000 ;
        RECT 5.075000 1.945000 5.265000 3.075000 ;
        RECT 5.185000 0.615000 5.515000 1.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.135000  0.305000  0.385000 1.075000 ;
      RECT 0.135000  1.075000  2.975000 1.085000 ;
      RECT 0.135000  1.085000  3.825000 1.255000 ;
      RECT 0.265000  1.815000  0.475000 3.245000 ;
      RECT 0.565000  0.085000  0.895000 0.905000 ;
      RECT 0.695000  1.815000  0.885000 2.350000 ;
      RECT 0.695000  2.350000  1.785000 2.520000 ;
      RECT 0.695000  2.520000  0.895000 3.075000 ;
      RECT 1.065000  0.305000  1.255000 1.075000 ;
      RECT 1.065000  2.690000  1.395000 3.245000 ;
      RECT 1.425000  0.085000  1.755000 0.905000 ;
      RECT 1.575000  2.520000  1.785000 2.800000 ;
      RECT 1.575000  2.800000  3.575000 3.075000 ;
      RECT 1.925000  0.305000  2.115000 1.075000 ;
      RECT 2.285000  0.085000  2.615000 0.905000 ;
      RECT 2.785000  0.305000  2.975000 1.075000 ;
      RECT 3.145000  0.085000  3.485000 0.915000 ;
      RECT 3.655000  0.265000  5.945000 0.435000 ;
      RECT 3.655000  0.435000  3.985000 0.905000 ;
      RECT 3.655000  0.905000  3.825000 1.085000 ;
      RECT 3.745000  2.800000  4.045000 3.245000 ;
      RECT 4.345000  1.425000  5.725000 1.595000 ;
      RECT 4.575000  2.115000  4.905000 3.245000 ;
      RECT 4.675000  0.435000  5.005000 0.895000 ;
      RECT 5.435000  2.125000  6.110000 3.245000 ;
      RECT 5.555000  1.595000  5.725000 1.765000 ;
      RECT 5.555000  1.765000  9.995000 1.945000 ;
      RECT 5.685000  0.435000  5.945000 1.040000 ;
      RECT 6.135000  0.305000  6.395000 0.870000 ;
      RECT 6.135000  0.870000  7.255000 1.040000 ;
      RECT 6.280000  1.945000  6.470000 3.075000 ;
      RECT 6.565000  0.085000  6.895000 0.700000 ;
      RECT 6.640000  2.125000  6.970000 3.245000 ;
      RECT 7.055000  1.040000  7.255000 1.075000 ;
      RECT 7.055000  1.075000  8.115000 1.245000 ;
      RECT 7.065000  0.305000  7.255000 0.870000 ;
      RECT 7.140000  1.945000  7.330000 3.075000 ;
      RECT 7.425000  0.085000  7.755000 0.905000 ;
      RECT 7.500000  2.125000  8.170000 3.245000 ;
      RECT 7.925000  0.265000  9.985000 0.435000 ;
      RECT 7.925000  0.435000  8.115000 1.075000 ;
      RECT 8.285000  0.605000  8.585000 0.815000 ;
      RECT 8.285000  0.815000  9.475000 1.000000 ;
      RECT 8.340000  1.945000  8.530000 3.075000 ;
      RECT 8.700000  2.125000  9.030000 3.245000 ;
      RECT 8.755000  0.435000  8.975000 0.635000 ;
      RECT 9.145000  0.605000  9.475000 0.815000 ;
      RECT 9.145000  1.000000  9.475000 1.075000 ;
      RECT 9.145000  1.075000  9.995000 1.255000 ;
      RECT 9.210000  1.945000  9.390000 3.075000 ;
      RECT 9.560000  2.115000  9.890000 3.245000 ;
      RECT 9.655000  0.435000  9.985000 0.905000 ;
      RECT 9.815000  1.255000  9.995000 1.765000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__o2bb2ai_4
END LIBRARY
