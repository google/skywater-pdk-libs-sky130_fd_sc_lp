* File: sky130_fd_sc_lp__a2111oi_4.pxi.spice
* Created: Wed Sep  2 09:17:02 2020
* 
x_PM_SKY130_FD_SC_LP__A2111OI_4%D1 N_D1_c_153_n N_D1_M1014_g N_D1_M1000_g
+ N_D1_c_155_n N_D1_M1022_g N_D1_M1016_g N_D1_c_157_n N_D1_M1023_g N_D1_M1027_g
+ N_D1_c_159_n N_D1_M1039_g N_D1_M1038_g D1 D1 D1 N_D1_c_162_n
+ PM_SKY130_FD_SC_LP__A2111OI_4%D1
x_PM_SKY130_FD_SC_LP__A2111OI_4%C1 N_C1_M1009_g N_C1_M1006_g N_C1_M1018_g
+ N_C1_M1010_g N_C1_M1031_g N_C1_M1030_g N_C1_M1034_g N_C1_M1032_g C1 C1 C1 C1
+ N_C1_c_245_n PM_SKY130_FD_SC_LP__A2111OI_4%C1
x_PM_SKY130_FD_SC_LP__A2111OI_4%B1 N_B1_M1001_g N_B1_M1007_g N_B1_M1003_g
+ N_B1_M1011_g N_B1_M1019_g N_B1_M1033_g N_B1_M1025_g N_B1_M1035_g B1 B1 B1 B1
+ N_B1_c_345_n PM_SKY130_FD_SC_LP__A2111OI_4%B1
x_PM_SKY130_FD_SC_LP__A2111OI_4%A1 N_A1_M1008_g N_A1_c_438_n N_A1_M1002_g
+ N_A1_M1020_g N_A1_c_440_n N_A1_M1013_g N_A1_M1024_g N_A1_c_442_n N_A1_M1015_g
+ N_A1_M1028_g N_A1_c_444_n N_A1_M1029_g A1 A1 A1 A1 N_A1_c_445_n N_A1_c_446_n
+ PM_SKY130_FD_SC_LP__A2111OI_4%A1
x_PM_SKY130_FD_SC_LP__A2111OI_4%A2 N_A2_M1012_g N_A2_M1004_g N_A2_M1017_g
+ N_A2_M1005_g N_A2_M1036_g N_A2_M1021_g N_A2_M1037_g N_A2_M1026_g N_A2_c_535_n
+ N_A2_c_536_n A2 N_A2_c_537_n N_A2_c_542_n PM_SKY130_FD_SC_LP__A2111OI_4%A2
x_PM_SKY130_FD_SC_LP__A2111OI_4%A_27_367# N_A_27_367#_M1000_s
+ N_A_27_367#_M1016_s N_A_27_367#_M1038_s N_A_27_367#_M1010_s
+ N_A_27_367#_M1032_s N_A_27_367#_c_609_n N_A_27_367#_c_610_n
+ N_A_27_367#_c_616_n N_A_27_367#_c_618_n N_A_27_367#_c_622_n
+ N_A_27_367#_c_624_n N_A_27_367#_c_634_n N_A_27_367#_c_636_n
+ N_A_27_367#_c_611_n N_A_27_367#_c_612_n N_A_27_367#_c_627_n
+ N_A_27_367#_c_629_n N_A_27_367#_c_645_n
+ PM_SKY130_FD_SC_LP__A2111OI_4%A_27_367#
x_PM_SKY130_FD_SC_LP__A2111OI_4%Y N_Y_M1014_d N_Y_M1023_d N_Y_M1009_s
+ N_Y_M1031_s N_Y_M1001_d N_Y_M1019_d N_Y_M1002_d N_Y_M1015_d N_Y_M1000_d
+ N_Y_M1027_d N_Y_c_689_n N_Y_c_705_n N_Y_c_797_p N_Y_c_699_n N_Y_c_700_n
+ N_Y_c_813_p N_Y_c_788_n N_Y_c_709_n N_Y_c_701_n N_Y_c_811_p N_Y_c_791_n
+ N_Y_c_718_n N_Y_c_812_p N_Y_c_690_n N_Y_c_735_n N_Y_c_691_n N_Y_c_740_n
+ N_Y_c_692_n N_Y_c_693_n N_Y_c_833_p N_Y_c_772_n N_Y_c_720_n N_Y_c_702_n
+ N_Y_c_724_n N_Y_c_694_n N_Y_c_695_n N_Y_c_696_n N_Y_c_776_n N_Y_c_778_n Y Y
+ N_Y_c_763_n Y N_Y_c_697_n PM_SKY130_FD_SC_LP__A2111OI_4%Y
x_PM_SKY130_FD_SC_LP__A2111OI_4%A_454_367# N_A_454_367#_M1006_d
+ N_A_454_367#_M1030_d N_A_454_367#_M1007_d N_A_454_367#_M1033_d
+ N_A_454_367#_c_843_n N_A_454_367#_c_842_n N_A_454_367#_c_857_n
+ N_A_454_367#_c_850_n N_A_454_367#_c_852_n N_A_454_367#_c_861_n
+ N_A_454_367#_c_863_n PM_SKY130_FD_SC_LP__A2111OI_4%A_454_367#
x_PM_SKY130_FD_SC_LP__A2111OI_4%A_819_367# N_A_819_367#_M1007_s
+ N_A_819_367#_M1011_s N_A_819_367#_M1035_s N_A_819_367#_M1020_d
+ N_A_819_367#_M1028_d N_A_819_367#_M1017_s N_A_819_367#_M1037_s
+ N_A_819_367#_c_893_n N_A_819_367#_c_907_n N_A_819_367#_c_894_n
+ N_A_819_367#_c_954_n N_A_819_367#_c_910_n N_A_819_367#_c_966_p
+ N_A_819_367#_c_895_n N_A_819_367#_c_889_n N_A_819_367#_c_890_n
+ N_A_819_367#_c_898_n N_A_819_367#_c_891_n N_A_819_367#_c_900_n
+ N_A_819_367#_c_969_p N_A_819_367#_c_934_n N_A_819_367#_c_901_n
+ N_A_819_367#_c_970_p N_A_819_367#_c_902_n N_A_819_367#_c_903_n
+ N_A_819_367#_c_967_p N_A_819_367#_c_892_n
+ PM_SKY130_FD_SC_LP__A2111OI_4%A_819_367#
x_PM_SKY130_FD_SC_LP__A2111OI_4%VPWR N_VPWR_M1008_s N_VPWR_M1024_s
+ N_VPWR_M1012_d N_VPWR_M1036_d N_VPWR_c_989_n N_VPWR_c_990_n N_VPWR_c_991_n
+ N_VPWR_c_992_n N_VPWR_c_993_n N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_996_n
+ N_VPWR_c_997_n N_VPWR_c_998_n N_VPWR_c_999_n N_VPWR_c_1000_n VPWR
+ N_VPWR_c_1001_n N_VPWR_c_988_n PM_SKY130_FD_SC_LP__A2111OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A2111OI_4%VGND N_VGND_M1014_s N_VGND_M1022_s
+ N_VGND_M1039_s N_VGND_M1018_d N_VGND_M1034_d N_VGND_M1003_s N_VGND_M1025_s
+ N_VGND_M1004_s N_VGND_M1021_s N_VGND_c_1116_n N_VGND_c_1117_n N_VGND_c_1118_n
+ N_VGND_c_1119_n N_VGND_c_1120_n N_VGND_c_1121_n N_VGND_c_1122_n
+ N_VGND_c_1123_n N_VGND_c_1124_n N_VGND_c_1125_n N_VGND_c_1126_n
+ N_VGND_c_1127_n N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n
+ N_VGND_c_1131_n N_VGND_c_1132_n N_VGND_c_1133_n VGND N_VGND_c_1134_n
+ N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n
+ N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n
+ N_VGND_c_1143_n PM_SKY130_FD_SC_LP__A2111OI_4%VGND
x_PM_SKY130_FD_SC_LP__A2111OI_4%A_1201_47# N_A_1201_47#_M1002_s
+ N_A_1201_47#_M1013_s N_A_1201_47#_M1029_s N_A_1201_47#_M1005_d
+ N_A_1201_47#_M1026_d N_A_1201_47#_c_1278_n N_A_1201_47#_c_1303_n
+ N_A_1201_47#_c_1280_n N_A_1201_47#_c_1319_n N_A_1201_47#_c_1282_n
+ N_A_1201_47#_c_1271_n N_A_1201_47#_c_1272_n N_A_1201_47#_c_1323_n
+ N_A_1201_47#_c_1273_n N_A_1201_47#_c_1274_n N_A_1201_47#_c_1275_n
+ N_A_1201_47#_c_1332_n N_A_1201_47#_c_1276_n
+ PM_SKY130_FD_SC_LP__A2111OI_4%A_1201_47#
cc_1 VNB N_D1_c_153_n 0.0184169f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_D1_M1000_g 0.00761757f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_D1_c_155_n 0.0160024f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.185
cc_4 VNB N_D1_M1016_g 0.00706401f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_5 VNB N_D1_c_157_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_6 VNB N_D1_M1027_g 0.0070671f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_7 VNB N_D1_c_159_n 0.0161951f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_8 VNB N_D1_M1038_g 0.00689767f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_9 VNB D1 0.00252193f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_10 VNB N_D1_c_162_n 0.0777785f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.35
cc_11 VNB N_C1_M1009_g 0.0245129f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_12 VNB N_C1_M1018_g 0.0227171f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.515
cc_13 VNB N_C1_M1031_g 0.0227174f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_14 VNB N_C1_M1034_g 0.0246415f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_15 VNB C1 0.00416985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_c_245_n 0.0760402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_M1001_g 0.0246425f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_18 VNB N_B1_M1003_g 0.0226997f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.515
cc_19 VNB N_B1_M1019_g 0.0228546f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_20 VNB N_B1_M1025_g 0.0312008f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_21 VNB B1 0.00323207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_345_n 0.0867462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_M1008_g 0.00685677f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_24 VNB N_A1_c_438_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_25 VNB N_A1_M1020_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_26 VNB N_A1_c_440_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_27 VNB N_A1_M1024_g 0.00677278f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_28 VNB N_A1_c_442_n 0.0162029f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_29 VNB N_A1_M1028_g 0.00750138f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_30 VNB N_A1_c_444_n 0.0172087f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_31 VNB N_A1_c_445_n 0.00588109f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.322
cc_32 VNB N_A1_c_446_n 0.10306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_M1012_g 0.00150975f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_34 VNB N_A2_M1004_g 0.0218807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_M1017_g 0.00145535f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.515
cc_36 VNB N_A2_M1005_g 0.0204793f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.185
cc_37 VNB N_A2_M1036_g 0.00157222f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_38 VNB N_A2_M1021_g 0.0204793f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_39 VNB N_A2_M1037_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_40 VNB N_A2_M1026_g 0.0277576f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_41 VNB N_A2_c_535_n 0.00684221f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.35
cc_42 VNB N_A2_c_536_n 0.0577683f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.35
cc_43 VNB N_A2_c_537_n 0.0863888f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.35
cc_44 VNB N_Y_c_689_n 0.0273694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_690_n 0.00901485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_691_n 0.00990539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_692_n 0.0076266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Y_c_693_n 0.016978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_Y_c_694_n 0.00357956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Y_c_695_n 0.00186402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Y_c_696_n 0.00186402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_Y_c_697_n 0.00368581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_819_367#_c_889_n 0.00289786f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.35
cc_54 VNB N_A_819_367#_c_890_n 0.00206162f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.35
cc_55 VNB N_A_819_367#_c_891_n 0.00622705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_819_367#_c_892_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_988_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1116_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1117_n 0.0221009f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_60 VNB N_VGND_c_1118_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1119_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.35
cc_62 VNB N_VGND_c_1120_n 3.19317e-19 $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.35
cc_63 VNB N_VGND_c_1121_n 0.0152106f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.35
cc_64 VNB N_VGND_c_1122_n 0.00427232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1123_n 0.0149762f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.322
cc_66 VNB N_VGND_c_1124_n 0.00175469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1125_n 0.00792815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1126_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1127_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1128_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1129_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1130_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1131_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1132_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1133_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1134_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1135_n 0.0152106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1136_n 0.0593468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1137_n 0.0196718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1138_n 0.484703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1139_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1140_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1141_n 0.0039769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1142_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1143_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1201_47#_c_1271_n 0.00289786f $X=-0.19 $Y=-0.245 $X2=1.765
+ $Y2=2.465
cc_87 VNB N_A_1201_47#_c_1272_n 0.00524313f $X=-0.19 $Y=-0.245 $X2=1.765
+ $Y2=2.465
cc_88 VNB N_A_1201_47#_c_1273_n 0.0119905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1201_47#_c_1274_n 0.0296037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1201_47#_c_1275_n 0.00526146f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=1.35
cc_91 VNB N_A_1201_47#_c_1276_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VPB N_D1_M1000_g 0.0234875f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_93 VPB N_D1_M1016_g 0.0186758f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_94 VPB N_D1_M1027_g 0.0186943f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_95 VPB N_D1_M1038_g 0.0200559f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_96 VPB N_C1_M1006_g 0.0182386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_C1_M1010_g 0.0180542f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.185
cc_98 VPB N_C1_M1030_g 0.0180542f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.655
cc_99 VPB N_C1_M1032_g 0.024227f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_100 VPB C1 0.0132503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_C1_c_245_n 0.019717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_B1_M1007_g 0.024227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_B1_M1011_g 0.0180542f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.185
cc_104 VPB N_B1_M1033_g 0.0180507f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.655
cc_105 VPB N_B1_M1035_g 0.0186689f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_106 VPB B1 0.0123631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_B1_c_345_n 0.0248041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A1_M1008_g 0.018727f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_109 VPB N_A1_M1020_g 0.0185652f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.655
cc_110 VPB N_A1_M1024_g 0.0188161f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.655
cc_111 VPB N_A1_M1028_g 0.0202673f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=0.655
cc_112 VPB N_A2_M1012_g 0.020758f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_113 VPB N_A2_M1017_g 0.0201993f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.515
cc_114 VPB N_A2_M1036_g 0.0196247f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_115 VPB N_A2_M1037_g 0.0248454f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_116 VPB N_A2_c_542_n 0.00260877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_27_367#_c_609_n 0.00746637f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.655
cc_118 VPB N_A_27_367#_c_610_n 0.0348412f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.515
cc_119 VPB N_A_27_367#_c_611_n 0.0018268f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.35
cc_120 VPB N_A_27_367#_c_612_n 0.006028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_Y_c_689_n 0.00229001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_Y_c_699_n 0.00167596f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_123 VPB N_Y_c_700_n 0.00567923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_Y_c_701_n 0.00683765f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.322
cc_125 VPB N_Y_c_702_n 0.00172998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_454_367#_c_842_n 0.0120055f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_127 VPB N_A_819_367#_c_893_n 0.00596005f $X=-0.19 $Y=1.655 $X2=1.765
+ $Y2=0.655
cc_128 VPB N_A_819_367#_c_894_n 0.0018268f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_129 VPB N_A_819_367#_c_895_n 0.00112894f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.35
cc_130 VPB N_A_819_367#_c_889_n 0.00559032f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.35
cc_131 VPB N_A_819_367#_c_890_n 9.84893e-19 $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.35
cc_132 VPB N_A_819_367#_c_898_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.35
cc_133 VPB N_A_819_367#_c_891_n 0.00609925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_819_367#_c_900_n 0.00116335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_819_367#_c_901_n 0.00247465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_819_367#_c_902_n 0.0119591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_819_367#_c_903_n 0.0450352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_989_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.185
cc_139 VPB N_VPWR_c_990_n 3.31161e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_991_n 3.46032e-19 $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_141 VPB N_VPWR_c_992_n 4.14e-19 $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_142 VPB N_VPWR_c_993_n 0.142827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_994_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.35
cc_144 VPB N_VPWR_c_995_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.35
cc_145 VPB N_VPWR_c_996_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.35
cc_146 VPB N_VPWR_c_997_n 0.0160778f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.35
cc_147 VPB N_VPWR_c_998_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=1.35
cc_148 VPB N_VPWR_c_999_n 0.0149571f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.35
cc_149 VPB N_VPWR_c_1000_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_1001_n 0.0220585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_988_n 0.0632693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 N_D1_c_159_n N_C1_M1009_g 0.0378259f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_153 D1 N_C1_M1009_g 7.19099e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_D1_M1038_g N_C1_M1006_g 0.0181962f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_155 N_D1_M1038_g C1 0.00128594f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_156 D1 C1 5.70818e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_157 N_D1_c_162_n C1 0.00168126f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_158 D1 N_C1_c_245_n 6.27594e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_D1_c_162_n N_C1_c_245_n 0.0209053f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_160 N_D1_M1000_g N_A_27_367#_c_609_n 5.81207e-19 $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_D1_M1000_g N_A_27_367#_c_610_n 0.0110657f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_162 N_D1_M1016_g N_A_27_367#_c_610_n 6.30056e-19 $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_D1_M1000_g N_A_27_367#_c_616_n 0.0105205f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_164 N_D1_M1016_g N_A_27_367#_c_616_n 0.0105205f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_165 N_D1_M1000_g N_A_27_367#_c_618_n 6.30056e-19 $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_D1_M1016_g N_A_27_367#_c_618_n 0.0103748f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_167 N_D1_M1027_g N_A_27_367#_c_618_n 0.0103748f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_168 N_D1_M1038_g N_A_27_367#_c_618_n 6.30056e-19 $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_D1_M1027_g N_A_27_367#_c_622_n 0.0105205f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_170 N_D1_M1038_g N_A_27_367#_c_622_n 0.0105205f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_171 N_D1_M1027_g N_A_27_367#_c_624_n 6.62591e-19 $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_D1_M1038_g N_A_27_367#_c_624_n 0.0129208f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_173 D1 N_A_27_367#_c_624_n 7.60446e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_174 N_D1_M1016_g N_A_27_367#_c_627_n 5.81207e-19 $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_D1_M1027_g N_A_27_367#_c_627_n 5.81207e-19 $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_D1_M1038_g N_A_27_367#_c_629_n 5.81207e-19 $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_D1_c_153_n N_Y_c_689_n 0.0241205f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_178 D1 N_Y_c_689_n 0.0178929f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_179 N_D1_c_153_n N_Y_c_705_n 0.014841f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_180 D1 N_Y_c_705_n 0.0057147f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_181 N_D1_M1000_g N_Y_c_699_n 0.0166275f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_182 D1 N_Y_c_699_n 0.00517328f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_183 N_D1_c_155_n N_Y_c_709_n 0.0122595f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_184 N_D1_c_157_n N_Y_c_709_n 0.0122595f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_185 D1 N_Y_c_709_n 0.039834f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_186 N_D1_c_162_n N_Y_c_709_n 0.00230884f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_187 N_D1_M1016_g N_Y_c_701_n 0.0143115f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_188 N_D1_M1027_g N_Y_c_701_n 0.014051f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_189 N_D1_M1038_g N_Y_c_701_n 0.00309561f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_190 D1 N_Y_c_701_n 0.0445191f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_191 N_D1_c_162_n N_Y_c_701_n 0.00472934f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_192 N_D1_c_159_n N_Y_c_718_n 0.0122129f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_193 D1 N_Y_c_718_n 0.0119493f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_194 D1 N_Y_c_720_n 0.0142048f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_195 N_D1_c_162_n N_Y_c_720_n 0.00240082f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_196 D1 N_Y_c_702_n 0.011071f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_197 N_D1_c_162_n N_Y_c_702_n 0.00242866f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_198 D1 N_Y_c_724_n 0.0142048f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_199 N_D1_c_162_n N_Y_c_724_n 0.00240082f $X=1.765 $Y=1.35 $X2=0 $Y2=0
cc_200 D1 N_Y_c_694_n 0.00165708f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_201 N_D1_M1000_g N_VPWR_c_993_n 0.00357842f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_202 N_D1_M1016_g N_VPWR_c_993_n 0.00357842f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_203 N_D1_M1027_g N_VPWR_c_993_n 0.00357842f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_204 N_D1_M1038_g N_VPWR_c_993_n 0.00357842f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_205 N_D1_M1000_g N_VPWR_c_988_n 0.00628379f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_206 N_D1_M1016_g N_VPWR_c_988_n 0.00535118f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_207 N_D1_M1027_g N_VPWR_c_988_n 0.00535118f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_208 N_D1_M1038_g N_VPWR_c_988_n 0.00537652f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_209 N_D1_c_153_n N_VGND_c_1117_n 0.0128375f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_210 N_D1_c_155_n N_VGND_c_1117_n 5.75816e-19 $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_211 N_D1_c_153_n N_VGND_c_1118_n 5.75816e-19 $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_212 N_D1_c_155_n N_VGND_c_1118_n 0.0105703f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_213 N_D1_c_157_n N_VGND_c_1118_n 0.0105703f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_214 N_D1_c_159_n N_VGND_c_1118_n 5.75816e-19 $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_215 N_D1_c_157_n N_VGND_c_1119_n 5.75816e-19 $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_216 N_D1_c_159_n N_VGND_c_1119_n 0.0104941f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_217 N_D1_c_157_n N_VGND_c_1128_n 0.00486043f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_218 N_D1_c_159_n N_VGND_c_1128_n 0.00486043f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_219 N_D1_c_153_n N_VGND_c_1134_n 0.00486043f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_220 N_D1_c_155_n N_VGND_c_1134_n 0.00486043f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_221 N_D1_c_153_n N_VGND_c_1138_n 0.00824727f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_222 N_D1_c_155_n N_VGND_c_1138_n 0.00824727f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_223 N_D1_c_157_n N_VGND_c_1138_n 0.00824727f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_224 N_D1_c_159_n N_VGND_c_1138_n 0.00824727f $X=1.765 $Y=1.185 $X2=0 $Y2=0
cc_225 N_C1_M1034_g N_B1_M1001_g 0.0238448f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_226 C1 N_B1_M1007_g 2.966e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_227 N_C1_M1032_g B1 4.41967e-19 $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_228 C1 B1 0.0245421f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_229 N_C1_c_245_n B1 3.08904e-19 $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_230 C1 N_B1_c_345_n 3.08904e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_231 N_C1_c_245_n N_B1_c_345_n 0.0230593f $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_232 N_C1_M1006_g N_A_27_367#_c_624_n 0.0126317f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_233 N_C1_M1010_g N_A_27_367#_c_624_n 6.14778e-19 $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_234 C1 N_A_27_367#_c_624_n 0.0053925f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_235 N_C1_c_245_n N_A_27_367#_c_624_n 2.9941e-19 $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_236 N_C1_M1006_g N_A_27_367#_c_634_n 0.0105205f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_237 N_C1_M1010_g N_A_27_367#_c_634_n 0.0105205f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_238 N_C1_M1006_g N_A_27_367#_c_636_n 5.66402e-19 $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_C1_M1010_g N_A_27_367#_c_636_n 0.00948562f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_C1_M1030_g N_A_27_367#_c_636_n 0.00948562f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_C1_M1032_g N_A_27_367#_c_636_n 5.66402e-19 $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_242 N_C1_M1030_g N_A_27_367#_c_611_n 0.0105205f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_243 N_C1_M1032_g N_A_27_367#_c_611_n 0.0111103f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_244 N_C1_M1030_g N_A_27_367#_c_612_n 5.66402e-19 $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_245 N_C1_M1032_g N_A_27_367#_c_612_n 0.0102119f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_246 N_C1_M1006_g N_A_27_367#_c_629_n 5.81207e-19 $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_C1_M1010_g N_A_27_367#_c_645_n 5.81207e-19 $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_248 N_C1_M1030_g N_A_27_367#_c_645_n 5.81207e-19 $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_249 C1 N_Y_c_701_n 0.00275099f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_250 N_C1_M1009_g N_Y_c_718_n 0.0133654f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_251 C1 N_Y_c_718_n 0.00784313f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_252 N_C1_c_245_n N_Y_c_718_n 0.00127178f $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_253 N_C1_M1018_g N_Y_c_690_n 0.0130736f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_254 N_C1_M1031_g N_Y_c_690_n 0.0142932f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_255 C1 N_Y_c_690_n 0.0492556f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_256 N_C1_c_245_n N_Y_c_690_n 0.00246472f $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_257 N_C1_M1031_g N_Y_c_735_n 6.15713e-19 $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_258 N_C1_M1034_g N_Y_c_735_n 0.0108881f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_259 N_C1_M1034_g N_Y_c_691_n 0.0124074f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_260 C1 N_Y_c_691_n 0.0231609f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_261 N_C1_c_245_n N_Y_c_691_n 0.0044365f $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_262 N_C1_M1034_g N_Y_c_740_n 6.50401e-19 $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_263 N_C1_M1009_g N_Y_c_694_n 0.0039223f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_264 N_C1_M1018_g N_Y_c_694_n 0.00101535f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_265 C1 N_Y_c_694_n 0.0166818f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_266 N_C1_c_245_n N_Y_c_694_n 0.00256759f $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_267 N_C1_M1034_g N_Y_c_695_n 0.00248804f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_268 C1 N_Y_c_695_n 0.0210392f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_269 N_C1_c_245_n N_Y_c_695_n 0.00256759f $X=3.575 $Y=1.51 $X2=0 $Y2=0
cc_270 N_C1_M1010_g N_A_454_367#_c_843_n 0.0122595f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_C1_M1030_g N_A_454_367#_c_843_n 0.0122129f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_272 C1 N_A_454_367#_c_843_n 0.0428505f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_273 N_C1_c_245_n N_A_454_367#_c_843_n 5.64665e-19 $X=3.575 $Y=1.51 $X2=0
+ $Y2=0
cc_274 N_C1_M1032_g N_A_454_367#_c_842_n 0.0143f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_275 C1 N_A_454_367#_c_842_n 0.024547f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_276 N_C1_c_245_n N_A_454_367#_c_842_n 9.10462e-19 $X=3.575 $Y=1.51 $X2=0
+ $Y2=0
cc_277 C1 N_A_454_367#_c_850_n 0.0154121f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_278 N_C1_c_245_n N_A_454_367#_c_850_n 6.37898e-19 $X=3.575 $Y=1.51 $X2=0
+ $Y2=0
cc_279 C1 N_A_454_367#_c_852_n 0.0154121f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_280 N_C1_c_245_n N_A_454_367#_c_852_n 6.37898e-19 $X=3.575 $Y=1.51 $X2=0
+ $Y2=0
cc_281 N_C1_M1032_g N_A_819_367#_c_893_n 0.00124397f $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_282 N_C1_M1006_g N_VPWR_c_993_n 0.00357842f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_283 N_C1_M1010_g N_VPWR_c_993_n 0.00357842f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_284 N_C1_M1030_g N_VPWR_c_993_n 0.00357842f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_285 N_C1_M1032_g N_VPWR_c_993_n 0.00357842f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_286 N_C1_M1006_g N_VPWR_c_988_n 0.00537652f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_287 N_C1_M1010_g N_VPWR_c_988_n 0.00535118f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_288 N_C1_M1030_g N_VPWR_c_988_n 0.00535118f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_289 N_C1_M1032_g N_VPWR_c_988_n 0.00682158f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_290 N_C1_M1009_g N_VGND_c_1119_n 0.0104941f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_291 N_C1_M1018_g N_VGND_c_1119_n 5.75816e-19 $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_292 N_C1_M1009_g N_VGND_c_1120_n 6.24193e-19 $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_293 N_C1_M1018_g N_VGND_c_1120_n 0.0117077f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_294 N_C1_M1031_g N_VGND_c_1120_n 0.011844f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_295 N_C1_M1034_g N_VGND_c_1120_n 7.13044e-19 $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_296 N_C1_M1031_g N_VGND_c_1121_n 0.00486043f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_297 N_C1_M1034_g N_VGND_c_1121_n 0.00564131f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_298 N_C1_M1034_g N_VGND_c_1122_n 0.00566589f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_299 N_C1_M1009_g N_VGND_c_1130_n 0.00486043f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_300 N_C1_M1018_g N_VGND_c_1130_n 0.00486043f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_301 N_C1_M1009_g N_VGND_c_1138_n 0.00824727f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_302 N_C1_M1018_g N_VGND_c_1138_n 0.00824727f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_303 N_C1_M1031_g N_VGND_c_1138_n 0.00824727f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_304 N_C1_M1034_g N_VGND_c_1138_n 0.0105044f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_305 B1 N_A1_M1008_g 7.18297e-19 $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_306 N_B1_c_345_n N_A1_M1008_g 0.0253841f $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_307 N_B1_M1025_g N_A1_c_445_n 0.00240464f $X=5.315 $Y=0.655 $X2=0 $Y2=0
cc_308 B1 N_A1_c_445_n 7.49417e-19 $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_309 N_B1_c_345_n N_A1_c_445_n 0.00238131f $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_310 N_B1_M1025_g N_A1_c_446_n 0.00244607f $X=5.315 $Y=0.655 $X2=0 $Y2=0
cc_311 B1 N_A1_c_446_n 0.00203151f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_312 N_B1_c_345_n N_A1_c_446_n 0.00542003f $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_313 N_B1_M1007_g N_A_27_367#_c_612_n 0.00126742f $X=4.435 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_B1_M1001_g N_Y_c_735_n 4.01631e-19 $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_315 N_B1_M1001_g N_Y_c_691_n 0.0131448f $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_316 B1 N_Y_c_691_n 0.0103335f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_317 N_B1_M1001_g N_Y_c_740_n 0.0102042f $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_318 N_B1_M1003_g N_Y_c_740_n 6.09683e-19 $X=4.455 $Y=0.655 $X2=0 $Y2=0
cc_319 N_B1_M1003_g N_Y_c_692_n 0.0142932f $X=4.455 $Y=0.655 $X2=0 $Y2=0
cc_320 N_B1_M1019_g N_Y_c_692_n 0.0118874f $X=4.885 $Y=0.655 $X2=0 $Y2=0
cc_321 B1 N_Y_c_692_n 0.0447626f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_322 N_B1_c_345_n N_Y_c_692_n 0.00255068f $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_323 N_B1_M1025_g N_Y_c_693_n 0.0154623f $X=5.315 $Y=0.655 $X2=0 $Y2=0
cc_324 B1 N_Y_c_693_n 0.016683f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_325 N_B1_c_345_n N_Y_c_693_n 0.00947039f $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_326 N_B1_M1001_g N_Y_c_696_n 0.002183f $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_327 B1 N_Y_c_696_n 0.0202401f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_328 N_B1_c_345_n N_Y_c_696_n 0.00256759f $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_329 N_B1_M1019_g N_Y_c_763_n 0.00701455f $X=4.885 $Y=0.655 $X2=0 $Y2=0
cc_330 N_B1_M1003_g N_Y_c_697_n 4.41847e-19 $X=4.455 $Y=0.655 $X2=0 $Y2=0
cc_331 N_B1_M1019_g N_Y_c_697_n 0.00558076f $X=4.885 $Y=0.655 $X2=0 $Y2=0
cc_332 N_B1_M1025_g N_Y_c_697_n 0.0049417f $X=5.315 $Y=0.655 $X2=0 $Y2=0
cc_333 B1 N_Y_c_697_n 0.0201948f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_334 N_B1_c_345_n N_Y_c_697_n 0.00265365f $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_335 N_B1_M1007_g N_A_454_367#_c_842_n 0.0143f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_336 B1 N_A_454_367#_c_842_n 0.0426898f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_337 N_B1_c_345_n N_A_454_367#_c_842_n 0.00218648f $X=5.475 $Y=1.51 $X2=0
+ $Y2=0
cc_338 N_B1_M1011_g N_A_454_367#_c_857_n 0.0136084f $X=4.865 $Y=2.465 $X2=0
+ $Y2=0
cc_339 N_B1_M1033_g N_A_454_367#_c_857_n 0.0116966f $X=5.295 $Y=2.465 $X2=0
+ $Y2=0
cc_340 B1 N_A_454_367#_c_857_n 0.0377771f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_341 N_B1_c_345_n N_A_454_367#_c_857_n 5.6803e-19 $X=5.475 $Y=1.51 $X2=0 $Y2=0
cc_342 B1 N_A_454_367#_c_861_n 0.0170883f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_343 N_B1_c_345_n N_A_454_367#_c_861_n 6.36429e-19 $X=5.475 $Y=1.51 $X2=0
+ $Y2=0
cc_344 N_B1_M1011_g N_A_454_367#_c_863_n 6.07415e-19 $X=4.865 $Y=2.465 $X2=0
+ $Y2=0
cc_345 N_B1_M1033_g N_A_454_367#_c_863_n 0.0102551f $X=5.295 $Y=2.465 $X2=0
+ $Y2=0
cc_346 N_B1_M1035_g N_A_454_367#_c_863_n 0.0103139f $X=5.725 $Y=2.465 $X2=0
+ $Y2=0
cc_347 B1 N_A_454_367#_c_863_n 0.0230948f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_348 N_B1_c_345_n N_A_454_367#_c_863_n 6.37898e-19 $X=5.475 $Y=1.51 $X2=0
+ $Y2=0
cc_349 N_B1_M1007_g N_A_819_367#_c_893_n 0.0105232f $X=4.435 $Y=2.465 $X2=0
+ $Y2=0
cc_350 N_B1_M1011_g N_A_819_367#_c_893_n 5.74651e-19 $X=4.865 $Y=2.465 $X2=0
+ $Y2=0
cc_351 N_B1_M1007_g N_A_819_367#_c_907_n 0.0105205f $X=4.435 $Y=2.465 $X2=0
+ $Y2=0
cc_352 N_B1_M1011_g N_A_819_367#_c_907_n 0.012237f $X=4.865 $Y=2.465 $X2=0 $Y2=0
cc_353 N_B1_M1007_g N_A_819_367#_c_894_n 5.89773e-19 $X=4.435 $Y=2.465 $X2=0
+ $Y2=0
cc_354 N_B1_M1033_g N_A_819_367#_c_910_n 0.0114565f $X=5.295 $Y=2.465 $X2=0
+ $Y2=0
cc_355 N_B1_M1035_g N_A_819_367#_c_910_n 0.0114588f $X=5.725 $Y=2.465 $X2=0
+ $Y2=0
cc_356 N_B1_M1035_g N_A_819_367#_c_895_n 0.00208503f $X=5.725 $Y=2.465 $X2=0
+ $Y2=0
cc_357 B1 N_A_819_367#_c_890_n 0.0136855f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_358 N_B1_c_345_n N_A_819_367#_c_890_n 0.00190497f $X=5.475 $Y=1.51 $X2=0
+ $Y2=0
cc_359 N_B1_M1035_g N_VPWR_c_989_n 0.00109252f $X=5.725 $Y=2.465 $X2=0 $Y2=0
cc_360 N_B1_M1007_g N_VPWR_c_993_n 0.00357842f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_361 N_B1_M1011_g N_VPWR_c_993_n 0.00357877f $X=4.865 $Y=2.465 $X2=0 $Y2=0
cc_362 N_B1_M1033_g N_VPWR_c_993_n 0.00357877f $X=5.295 $Y=2.465 $X2=0 $Y2=0
cc_363 N_B1_M1035_g N_VPWR_c_993_n 0.00357877f $X=5.725 $Y=2.465 $X2=0 $Y2=0
cc_364 N_B1_M1007_g N_VPWR_c_988_n 0.00673168f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_365 N_B1_M1011_g N_VPWR_c_988_n 0.0053512f $X=4.865 $Y=2.465 $X2=0 $Y2=0
cc_366 N_B1_M1033_g N_VPWR_c_988_n 0.0053512f $X=5.295 $Y=2.465 $X2=0 $Y2=0
cc_367 N_B1_M1035_g N_VPWR_c_988_n 0.00537654f $X=5.725 $Y=2.465 $X2=0 $Y2=0
cc_368 N_B1_M1001_g N_VGND_c_1122_n 0.00209888f $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_369 N_B1_M1001_g N_VGND_c_1123_n 0.00579312f $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_370 N_B1_M1003_g N_VGND_c_1123_n 0.00486043f $X=4.455 $Y=0.655 $X2=0 $Y2=0
cc_371 N_B1_M1001_g N_VGND_c_1124_n 7.05142e-19 $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_372 N_B1_M1003_g N_VGND_c_1124_n 0.0107763f $X=4.455 $Y=0.655 $X2=0 $Y2=0
cc_373 N_B1_M1019_g N_VGND_c_1124_n 0.00152071f $X=4.885 $Y=0.655 $X2=0 $Y2=0
cc_374 N_B1_M1019_g N_VGND_c_1125_n 6.31226e-19 $X=4.885 $Y=0.655 $X2=0 $Y2=0
cc_375 N_B1_M1025_g N_VGND_c_1125_n 0.0126799f $X=5.315 $Y=0.655 $X2=0 $Y2=0
cc_376 N_B1_M1019_g N_VGND_c_1135_n 0.00564131f $X=4.885 $Y=0.655 $X2=0 $Y2=0
cc_377 N_B1_M1025_g N_VGND_c_1135_n 0.00486043f $X=5.315 $Y=0.655 $X2=0 $Y2=0
cc_378 N_B1_M1001_g N_VGND_c_1138_n 0.0106925f $X=4.025 $Y=0.655 $X2=0 $Y2=0
cc_379 N_B1_M1003_g N_VGND_c_1138_n 0.00824727f $X=4.455 $Y=0.655 $X2=0 $Y2=0
cc_380 N_B1_M1019_g N_VGND_c_1138_n 0.0101089f $X=4.885 $Y=0.655 $X2=0 $Y2=0
cc_381 N_B1_M1025_g N_VGND_c_1138_n 0.00824727f $X=5.315 $Y=0.655 $X2=0 $Y2=0
cc_382 N_B1_M1025_g N_A_1201_47#_c_1275_n 0.00105173f $X=5.315 $Y=0.655 $X2=0
+ $Y2=0
cc_383 N_A1_c_444_n N_A2_M1004_g 0.0235382f $X=7.655 $Y=1.185 $X2=0 $Y2=0
cc_384 N_A1_c_445_n N_A2_M1004_g 4.57746e-19 $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_385 N_A1_M1028_g N_A2_c_537_n 0.0288051f $X=7.465 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A1_c_445_n N_A2_c_537_n 7.98138e-19 $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_387 N_A1_c_446_n N_A2_c_537_n 0.0163596f $X=7.655 $Y=1.35 $X2=0 $Y2=0
cc_388 N_A1_M1028_g N_A2_c_542_n 6.47733e-19 $X=7.465 $Y=2.465 $X2=0 $Y2=0
cc_389 N_A1_c_445_n N_A2_c_542_n 0.00365558f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_390 N_A1_c_446_n N_A2_c_542_n 8.46471e-19 $X=7.655 $Y=1.35 $X2=0 $Y2=0
cc_391 N_A1_c_438_n N_Y_c_693_n 0.0129296f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_392 N_A1_c_445_n N_Y_c_693_n 0.0417922f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_393 N_A1_c_446_n N_Y_c_693_n 0.00718335f $X=7.655 $Y=1.35 $X2=0 $Y2=0
cc_394 N_A1_c_440_n N_Y_c_772_n 0.0108425f $X=6.795 $Y=1.185 $X2=0 $Y2=0
cc_395 N_A1_c_442_n N_Y_c_772_n 0.01014f $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_396 N_A1_c_445_n N_Y_c_772_n 0.0376019f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_397 N_A1_c_446_n N_Y_c_772_n 0.00271364f $X=7.655 $Y=1.35 $X2=0 $Y2=0
cc_398 N_A1_c_445_n N_Y_c_776_n 0.015706f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_399 N_A1_c_446_n N_Y_c_776_n 0.00277275f $X=7.655 $Y=1.35 $X2=0 $Y2=0
cc_400 N_A1_c_444_n N_Y_c_778_n 0.00701021f $X=7.655 $Y=1.185 $X2=0 $Y2=0
cc_401 N_A1_c_445_n N_Y_c_778_n 0.0183602f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_402 N_A1_c_446_n N_Y_c_778_n 0.00277275f $X=7.655 $Y=1.35 $X2=0 $Y2=0
cc_403 N_A1_c_445_n N_Y_c_697_n 0.00157043f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_404 N_A1_M1008_g N_A_819_367#_c_895_n 0.0014373f $X=6.155 $Y=2.465 $X2=0
+ $Y2=0
cc_405 N_A1_M1008_g N_A_819_367#_c_889_n 0.0138902f $X=6.155 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_A1_M1020_g N_A_819_367#_c_889_n 0.0142932f $X=6.585 $Y=2.465 $X2=0
+ $Y2=0
cc_407 N_A1_c_445_n N_A_819_367#_c_889_n 0.0477254f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_408 N_A1_c_446_n N_A_819_367#_c_889_n 0.00400107f $X=7.655 $Y=1.35 $X2=0
+ $Y2=0
cc_409 N_A1_c_445_n N_A_819_367#_c_890_n 0.0162617f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_410 N_A1_c_446_n N_A_819_367#_c_890_n 6.41898e-19 $X=7.655 $Y=1.35 $X2=0
+ $Y2=0
cc_411 N_A1_M1020_g N_A_819_367#_c_898_n 0.0014373f $X=6.585 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A1_M1024_g N_A_819_367#_c_898_n 0.0014373f $X=7.015 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A1_M1024_g N_A_819_367#_c_891_n 0.0144087f $X=7.015 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_A1_M1028_g N_A_819_367#_c_891_n 0.0149854f $X=7.465 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_A1_c_445_n N_A_819_367#_c_891_n 0.0588189f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_416 N_A1_c_446_n N_A_819_367#_c_891_n 0.00982516f $X=7.655 $Y=1.35 $X2=0
+ $Y2=0
cc_417 N_A1_M1028_g N_A_819_367#_c_900_n 9.33414e-19 $X=7.465 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A1_c_445_n N_A_819_367#_c_892_n 0.0156157f $X=7.535 $Y=1.35 $X2=0 $Y2=0
cc_419 N_A1_c_446_n N_A_819_367#_c_892_n 0.00299787f $X=7.655 $Y=1.35 $X2=0
+ $Y2=0
cc_420 N_A1_M1008_g N_VPWR_c_989_n 0.0185929f $X=6.155 $Y=2.465 $X2=0 $Y2=0
cc_421 N_A1_M1020_g N_VPWR_c_989_n 0.01742f $X=6.585 $Y=2.465 $X2=0 $Y2=0
cc_422 N_A1_M1024_g N_VPWR_c_989_n 7.69607e-19 $X=7.015 $Y=2.465 $X2=0 $Y2=0
cc_423 N_A1_M1020_g N_VPWR_c_990_n 7.69607e-19 $X=6.585 $Y=2.465 $X2=0 $Y2=0
cc_424 N_A1_M1024_g N_VPWR_c_990_n 0.0176121f $X=7.015 $Y=2.465 $X2=0 $Y2=0
cc_425 N_A1_M1028_g N_VPWR_c_990_n 0.0155689f $X=7.465 $Y=2.465 $X2=0 $Y2=0
cc_426 N_A1_M1028_g N_VPWR_c_991_n 5.99575e-19 $X=7.465 $Y=2.465 $X2=0 $Y2=0
cc_427 N_A1_M1008_g N_VPWR_c_993_n 0.00486043f $X=6.155 $Y=2.465 $X2=0 $Y2=0
cc_428 N_A1_M1020_g N_VPWR_c_995_n 0.00486043f $X=6.585 $Y=2.465 $X2=0 $Y2=0
cc_429 N_A1_M1024_g N_VPWR_c_995_n 0.00486043f $X=7.015 $Y=2.465 $X2=0 $Y2=0
cc_430 N_A1_M1028_g N_VPWR_c_997_n 0.00564095f $X=7.465 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A1_M1008_g N_VPWR_c_988_n 0.0082726f $X=6.155 $Y=2.465 $X2=0 $Y2=0
cc_432 N_A1_M1020_g N_VPWR_c_988_n 0.00824727f $X=6.585 $Y=2.465 $X2=0 $Y2=0
cc_433 N_A1_M1024_g N_VPWR_c_988_n 0.00824727f $X=7.015 $Y=2.465 $X2=0 $Y2=0
cc_434 N_A1_M1028_g N_VPWR_c_988_n 0.00977012f $X=7.465 $Y=2.465 $X2=0 $Y2=0
cc_435 N_A1_c_438_n N_VGND_c_1125_n 0.00212298f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_436 N_A1_c_444_n N_VGND_c_1126_n 0.00121435f $X=7.655 $Y=1.185 $X2=0 $Y2=0
cc_437 N_A1_c_438_n N_VGND_c_1136_n 0.00357877f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_438 N_A1_c_440_n N_VGND_c_1136_n 0.00357877f $X=6.795 $Y=1.185 $X2=0 $Y2=0
cc_439 N_A1_c_442_n N_VGND_c_1136_n 0.00357877f $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_440 N_A1_c_444_n N_VGND_c_1136_n 0.00357877f $X=7.655 $Y=1.185 $X2=0 $Y2=0
cc_441 N_A1_c_438_n N_VGND_c_1138_n 0.0068216f $X=6.365 $Y=1.185 $X2=0 $Y2=0
cc_442 N_A1_c_440_n N_VGND_c_1138_n 0.00542194f $X=6.795 $Y=1.185 $X2=0 $Y2=0
cc_443 N_A1_c_442_n N_VGND_c_1138_n 0.00542194f $X=7.225 $Y=1.185 $X2=0 $Y2=0
cc_444 N_A1_c_444_n N_VGND_c_1138_n 0.00567744f $X=7.655 $Y=1.185 $X2=0 $Y2=0
cc_445 N_A1_c_438_n N_A_1201_47#_c_1278_n 0.00912428f $X=6.365 $Y=1.185 $X2=0
+ $Y2=0
cc_446 N_A1_c_440_n N_A_1201_47#_c_1278_n 0.0101276f $X=6.795 $Y=1.185 $X2=0
+ $Y2=0
cc_447 N_A1_c_442_n N_A_1201_47#_c_1280_n 0.0101276f $X=7.225 $Y=1.185 $X2=0
+ $Y2=0
cc_448 N_A1_c_444_n N_A_1201_47#_c_1280_n 0.013738f $X=7.655 $Y=1.185 $X2=0
+ $Y2=0
cc_449 N_A1_c_444_n N_A_1201_47#_c_1282_n 0.00746521f $X=7.655 $Y=1.185 $X2=0
+ $Y2=0
cc_450 N_A1_c_444_n N_A_1201_47#_c_1272_n 0.00496179f $X=7.655 $Y=1.185 $X2=0
+ $Y2=0
cc_451 N_A2_c_537_n N_A_819_367#_c_891_n 0.00167992f $X=9.545 $Y=1.46 $X2=0
+ $Y2=0
cc_452 N_A2_c_542_n N_A_819_367#_c_891_n 0.0134641f $X=8.485 $Y=1.567 $X2=0
+ $Y2=0
cc_453 N_A2_M1012_g N_A_819_367#_c_900_n 0.00351422f $X=8.015 $Y=2.465 $X2=0
+ $Y2=0
cc_454 N_A2_M1012_g N_A_819_367#_c_934_n 0.0148275f $X=8.015 $Y=2.465 $X2=0
+ $Y2=0
cc_455 N_A2_M1017_g N_A_819_367#_c_934_n 0.0147415f $X=8.445 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A2_c_535_n N_A_819_367#_c_934_n 0.00200155f $X=9.81 $Y=1.46 $X2=0 $Y2=0
cc_457 N_A2_c_537_n N_A_819_367#_c_934_n 4.97995e-19 $X=9.545 $Y=1.46 $X2=0
+ $Y2=0
cc_458 N_A2_c_542_n N_A_819_367#_c_934_n 0.0367614f $X=8.485 $Y=1.567 $X2=0
+ $Y2=0
cc_459 N_A2_M1017_g N_A_819_367#_c_901_n 0.00512717f $X=8.445 $Y=2.465 $X2=0
+ $Y2=0
cc_460 N_A2_c_535_n N_A_819_367#_c_901_n 0.0188266f $X=9.81 $Y=1.46 $X2=0 $Y2=0
cc_461 N_A2_c_537_n N_A_819_367#_c_901_n 0.0054037f $X=9.545 $Y=1.46 $X2=0 $Y2=0
cc_462 N_A2_c_542_n N_A_819_367#_c_901_n 0.00385841f $X=8.485 $Y=1.567 $X2=0
+ $Y2=0
cc_463 N_A2_M1036_g N_A_819_367#_c_902_n 0.0136053f $X=8.965 $Y=2.465 $X2=0
+ $Y2=0
cc_464 N_A2_M1037_g N_A_819_367#_c_902_n 0.0146218f $X=9.395 $Y=2.465 $X2=0
+ $Y2=0
cc_465 N_A2_c_535_n N_A_819_367#_c_902_n 0.0676667f $X=9.81 $Y=1.46 $X2=0 $Y2=0
cc_466 N_A2_c_537_n N_A_819_367#_c_902_n 0.0108698f $X=9.545 $Y=1.46 $X2=0 $Y2=0
cc_467 N_A2_M1012_g N_VPWR_c_990_n 7.44587e-19 $X=8.015 $Y=2.465 $X2=0 $Y2=0
cc_468 N_A2_M1012_g N_VPWR_c_991_n 0.0150766f $X=8.015 $Y=2.465 $X2=0 $Y2=0
cc_469 N_A2_M1017_g N_VPWR_c_991_n 0.0149385f $X=8.445 $Y=2.465 $X2=0 $Y2=0
cc_470 N_A2_M1036_g N_VPWR_c_991_n 6.14576e-19 $X=8.965 $Y=2.465 $X2=0 $Y2=0
cc_471 N_A2_M1017_g N_VPWR_c_992_n 6.85582e-19 $X=8.445 $Y=2.465 $X2=0 $Y2=0
cc_472 N_A2_M1036_g N_VPWR_c_992_n 0.0153268f $X=8.965 $Y=2.465 $X2=0 $Y2=0
cc_473 N_A2_M1037_g N_VPWR_c_992_n 0.0169864f $X=9.395 $Y=2.465 $X2=0 $Y2=0
cc_474 N_A2_M1012_g N_VPWR_c_997_n 0.00486043f $X=8.015 $Y=2.465 $X2=0 $Y2=0
cc_475 N_A2_M1017_g N_VPWR_c_999_n 0.00486043f $X=8.445 $Y=2.465 $X2=0 $Y2=0
cc_476 N_A2_M1036_g N_VPWR_c_999_n 0.00486043f $X=8.965 $Y=2.465 $X2=0 $Y2=0
cc_477 N_A2_M1037_g N_VPWR_c_1001_n 0.00486043f $X=9.395 $Y=2.465 $X2=0 $Y2=0
cc_478 N_A2_M1012_g N_VPWR_c_988_n 0.00866436f $X=8.015 $Y=2.465 $X2=0 $Y2=0
cc_479 N_A2_M1017_g N_VPWR_c_988_n 0.0084632f $X=8.445 $Y=2.465 $X2=0 $Y2=0
cc_480 N_A2_M1036_g N_VPWR_c_988_n 0.0084632f $X=8.965 $Y=2.465 $X2=0 $Y2=0
cc_481 N_A2_M1037_g N_VPWR_c_988_n 0.0093271f $X=9.395 $Y=2.465 $X2=0 $Y2=0
cc_482 N_A2_M1004_g N_VGND_c_1126_n 0.0118784f $X=8.18 $Y=0.655 $X2=0 $Y2=0
cc_483 N_A2_M1005_g N_VGND_c_1126_n 0.0106005f $X=8.61 $Y=0.655 $X2=0 $Y2=0
cc_484 N_A2_M1021_g N_VGND_c_1126_n 6.22495e-19 $X=9.04 $Y=0.655 $X2=0 $Y2=0
cc_485 N_A2_M1005_g N_VGND_c_1127_n 6.22495e-19 $X=8.61 $Y=0.655 $X2=0 $Y2=0
cc_486 N_A2_M1021_g N_VGND_c_1127_n 0.0106005f $X=9.04 $Y=0.655 $X2=0 $Y2=0
cc_487 N_A2_M1026_g N_VGND_c_1127_n 0.0123781f $X=9.47 $Y=0.655 $X2=0 $Y2=0
cc_488 N_A2_M1005_g N_VGND_c_1132_n 0.00486043f $X=8.61 $Y=0.655 $X2=0 $Y2=0
cc_489 N_A2_M1021_g N_VGND_c_1132_n 0.00486043f $X=9.04 $Y=0.655 $X2=0 $Y2=0
cc_490 N_A2_M1004_g N_VGND_c_1136_n 0.00486043f $X=8.18 $Y=0.655 $X2=0 $Y2=0
cc_491 N_A2_M1026_g N_VGND_c_1137_n 0.00486043f $X=9.47 $Y=0.655 $X2=0 $Y2=0
cc_492 N_A2_M1004_g N_VGND_c_1138_n 0.00848452f $X=8.18 $Y=0.655 $X2=0 $Y2=0
cc_493 N_A2_M1005_g N_VGND_c_1138_n 0.00824727f $X=8.61 $Y=0.655 $X2=0 $Y2=0
cc_494 N_A2_M1021_g N_VGND_c_1138_n 0.00824727f $X=9.04 $Y=0.655 $X2=0 $Y2=0
cc_495 N_A2_M1026_g N_VGND_c_1138_n 0.00928491f $X=9.47 $Y=0.655 $X2=0 $Y2=0
cc_496 N_A2_M1004_g N_A_1201_47#_c_1271_n 0.0137305f $X=8.18 $Y=0.655 $X2=0
+ $Y2=0
cc_497 N_A2_M1005_g N_A_1201_47#_c_1271_n 0.0137676f $X=8.61 $Y=0.655 $X2=0
+ $Y2=0
cc_498 N_A2_c_537_n N_A_1201_47#_c_1271_n 0.00419449f $X=9.545 $Y=1.46 $X2=0
+ $Y2=0
cc_499 N_A2_c_542_n N_A_1201_47#_c_1271_n 0.0486159f $X=8.485 $Y=1.567 $X2=0
+ $Y2=0
cc_500 N_A2_c_537_n N_A_1201_47#_c_1272_n 0.00371147f $X=9.545 $Y=1.46 $X2=0
+ $Y2=0
cc_501 N_A2_c_542_n N_A_1201_47#_c_1272_n 0.00980074f $X=8.485 $Y=1.567 $X2=0
+ $Y2=0
cc_502 N_A2_M1021_g N_A_1201_47#_c_1273_n 0.0138141f $X=9.04 $Y=0.655 $X2=0
+ $Y2=0
cc_503 N_A2_M1026_g N_A_1201_47#_c_1273_n 0.0148713f $X=9.47 $Y=0.655 $X2=0
+ $Y2=0
cc_504 N_A2_c_535_n N_A_1201_47#_c_1273_n 0.0676669f $X=9.81 $Y=1.46 $X2=0 $Y2=0
cc_505 N_A2_c_536_n N_A_1201_47#_c_1273_n 0.00776021f $X=9.81 $Y=1.46 $X2=0
+ $Y2=0
cc_506 N_A2_c_537_n N_A_1201_47#_c_1273_n 0.00278708f $X=9.545 $Y=1.46 $X2=0
+ $Y2=0
cc_507 N_A2_c_535_n N_A_1201_47#_c_1276_n 0.0153308f $X=9.81 $Y=1.46 $X2=0 $Y2=0
cc_508 N_A2_c_537_n N_A_1201_47#_c_1276_n 0.0028903f $X=9.545 $Y=1.46 $X2=0
+ $Y2=0
cc_509 N_A_27_367#_c_616_n N_Y_M1000_d 0.00332344f $X=0.955 $Y=2.99 $X2=0 $Y2=0
cc_510 N_A_27_367#_c_622_n N_Y_M1027_d 0.00332344f $X=1.815 $Y=2.99 $X2=0 $Y2=0
cc_511 N_A_27_367#_M1000_s N_Y_c_699_n 2.33864e-19 $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_512 N_A_27_367#_c_610_n N_Y_c_699_n 0.00362085f $X=0.26 $Y=2.13 $X2=0 $Y2=0
cc_513 N_A_27_367#_M1000_s N_Y_c_700_n 0.00397347f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_514 N_A_27_367#_c_610_n N_Y_c_700_n 0.0162291f $X=0.26 $Y=2.13 $X2=0 $Y2=0
cc_515 N_A_27_367#_c_616_n N_Y_c_788_n 0.0126348f $X=0.955 $Y=2.99 $X2=0 $Y2=0
cc_516 N_A_27_367#_M1016_s N_Y_c_701_n 0.00176461f $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_517 N_A_27_367#_c_618_n N_Y_c_701_n 0.0170777f $X=1.12 $Y=2.13 $X2=0 $Y2=0
cc_518 N_A_27_367#_c_622_n N_Y_c_791_n 0.0126348f $X=1.815 $Y=2.99 $X2=0 $Y2=0
cc_519 N_A_27_367#_c_634_n N_A_454_367#_M1006_d 0.00332344f $X=2.675 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_520 N_A_27_367#_c_611_n N_A_454_367#_M1030_d 0.00332344f $X=3.535 $Y=2.99
+ $X2=0 $Y2=0
cc_521 N_A_27_367#_M1010_s N_A_454_367#_c_843_n 0.00333177f $X=2.7 $Y=1.835
+ $X2=0 $Y2=0
cc_522 N_A_27_367#_c_636_n N_A_454_367#_c_843_n 0.0170777f $X=2.84 $Y=2.385
+ $X2=0 $Y2=0
cc_523 N_A_27_367#_M1032_s N_A_454_367#_c_842_n 0.00586493f $X=3.56 $Y=1.835
+ $X2=0 $Y2=0
cc_524 N_A_27_367#_c_612_n N_A_454_367#_c_842_n 0.0220026f $X=3.7 $Y=2.385 $X2=0
+ $Y2=0
cc_525 N_A_27_367#_c_634_n N_A_454_367#_c_850_n 0.0126348f $X=2.675 $Y=2.99
+ $X2=0 $Y2=0
cc_526 N_A_27_367#_c_611_n N_A_454_367#_c_852_n 0.0126348f $X=3.535 $Y=2.99
+ $X2=0 $Y2=0
cc_527 N_A_27_367#_c_612_n N_A_819_367#_c_893_n 0.0488195f $X=3.7 $Y=2.385 $X2=0
+ $Y2=0
cc_528 N_A_27_367#_c_611_n N_A_819_367#_c_894_n 0.0147157f $X=3.535 $Y=2.99
+ $X2=0 $Y2=0
cc_529 N_A_27_367#_c_609_n N_VPWR_c_993_n 0.0211538f $X=0.26 $Y=2.905 $X2=0
+ $Y2=0
cc_530 N_A_27_367#_c_616_n N_VPWR_c_993_n 0.0298674f $X=0.955 $Y=2.99 $X2=0
+ $Y2=0
cc_531 N_A_27_367#_c_622_n N_VPWR_c_993_n 0.0298674f $X=1.815 $Y=2.99 $X2=0
+ $Y2=0
cc_532 N_A_27_367#_c_634_n N_VPWR_c_993_n 0.0298674f $X=2.675 $Y=2.99 $X2=0
+ $Y2=0
cc_533 N_A_27_367#_c_611_n N_VPWR_c_993_n 0.0510539f $X=3.535 $Y=2.99 $X2=0
+ $Y2=0
cc_534 N_A_27_367#_c_627_n N_VPWR_c_993_n 0.0189946f $X=1.12 $Y=2.99 $X2=0 $Y2=0
cc_535 N_A_27_367#_c_629_n N_VPWR_c_993_n 0.0189946f $X=1.98 $Y=2.99 $X2=0 $Y2=0
cc_536 N_A_27_367#_c_645_n N_VPWR_c_993_n 0.0189946f $X=2.84 $Y=2.99 $X2=0 $Y2=0
cc_537 N_A_27_367#_M1000_s N_VPWR_c_988_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_538 N_A_27_367#_M1016_s N_VPWR_c_988_n 0.00223559f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_539 N_A_27_367#_M1038_s N_VPWR_c_988_n 0.00223559f $X=1.84 $Y=1.835 $X2=0
+ $Y2=0
cc_540 N_A_27_367#_M1010_s N_VPWR_c_988_n 0.00223559f $X=2.7 $Y=1.835 $X2=0
+ $Y2=0
cc_541 N_A_27_367#_M1032_s N_VPWR_c_988_n 0.00215962f $X=3.56 $Y=1.835 $X2=0
+ $Y2=0
cc_542 N_A_27_367#_c_609_n N_VPWR_c_988_n 0.0126374f $X=0.26 $Y=2.905 $X2=0
+ $Y2=0
cc_543 N_A_27_367#_c_616_n N_VPWR_c_988_n 0.0187823f $X=0.955 $Y=2.99 $X2=0
+ $Y2=0
cc_544 N_A_27_367#_c_622_n N_VPWR_c_988_n 0.0187823f $X=1.815 $Y=2.99 $X2=0
+ $Y2=0
cc_545 N_A_27_367#_c_634_n N_VPWR_c_988_n 0.0187823f $X=2.675 $Y=2.99 $X2=0
+ $Y2=0
cc_546 N_A_27_367#_c_611_n N_VPWR_c_988_n 0.0314875f $X=3.535 $Y=2.99 $X2=0
+ $Y2=0
cc_547 N_A_27_367#_c_627_n N_VPWR_c_988_n 0.0124451f $X=1.12 $Y=2.99 $X2=0 $Y2=0
cc_548 N_A_27_367#_c_629_n N_VPWR_c_988_n 0.0124451f $X=1.98 $Y=2.99 $X2=0 $Y2=0
cc_549 N_A_27_367#_c_645_n N_VPWR_c_988_n 0.0124451f $X=2.84 $Y=2.99 $X2=0 $Y2=0
cc_550 N_Y_c_691_n N_A_454_367#_c_842_n 0.00590406f $X=4.095 $Y=1.17 $X2=0 $Y2=0
cc_551 N_Y_M1000_d N_VPWR_c_988_n 0.00225186f $X=0.55 $Y=1.835 $X2=0 $Y2=0
cc_552 N_Y_M1027_d N_VPWR_c_988_n 0.00225186f $X=1.41 $Y=1.835 $X2=0 $Y2=0
cc_553 N_Y_c_689_n N_VGND_M1014_s 0.00183394f $X=0.23 $Y=1.705 $X2=-0.19
+ $Y2=-0.245
cc_554 N_Y_c_705_n N_VGND_M1014_s 6.72674e-19 $X=0.595 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_555 N_Y_c_797_p N_VGND_M1014_s 0.0104135f $X=0.32 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_556 N_Y_c_709_n N_VGND_M1022_s 0.00329816f $X=1.455 $Y=0.955 $X2=0 $Y2=0
cc_557 N_Y_c_718_n N_VGND_M1039_s 0.0077642f $X=2.305 $Y=0.955 $X2=0 $Y2=0
cc_558 N_Y_c_693_n N_VGND_M1025_s 0.00565861f $X=6.46 $Y=0.955 $X2=0 $Y2=0
cc_559 N_Y_c_705_n N_VGND_c_1117_n 0.00362085f $X=0.595 $Y=0.955 $X2=0 $Y2=0
cc_560 N_Y_c_797_p N_VGND_c_1117_n 0.0162291f $X=0.32 $Y=0.955 $X2=0 $Y2=0
cc_561 N_Y_c_709_n N_VGND_c_1118_n 0.0170777f $X=1.455 $Y=0.955 $X2=0 $Y2=0
cc_562 N_Y_c_718_n N_VGND_c_1119_n 0.0170777f $X=2.305 $Y=0.955 $X2=0 $Y2=0
cc_563 N_Y_c_690_n N_VGND_c_1120_n 0.0216087f $X=3.175 $Y=1.17 $X2=0 $Y2=0
cc_564 N_Y_c_735_n N_VGND_c_1121_n 0.0150063f $X=3.27 $Y=0.42 $X2=0 $Y2=0
cc_565 N_Y_c_691_n N_VGND_c_1122_n 0.0247883f $X=4.095 $Y=1.17 $X2=0 $Y2=0
cc_566 N_Y_c_740_n N_VGND_c_1123_n 0.0143246f $X=4.24 $Y=0.42 $X2=0 $Y2=0
cc_567 N_Y_c_692_n N_VGND_c_1124_n 0.0184616f $X=4.945 $Y=1.17 $X2=0 $Y2=0
cc_568 N_Y_c_693_n N_VGND_c_1125_n 0.021083f $X=6.46 $Y=0.955 $X2=0 $Y2=0
cc_569 N_Y_c_811_p N_VGND_c_1128_n 0.0124525f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_570 N_Y_c_812_p N_VGND_c_1130_n 0.0124525f $X=2.41 $Y=0.42 $X2=0 $Y2=0
cc_571 N_Y_c_813_p N_VGND_c_1134_n 0.0124525f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_572 N_Y_c_763_n N_VGND_c_1135_n 0.0150063f $X=5.1 $Y=0.42 $X2=0 $Y2=0
cc_573 N_Y_M1014_d N_VGND_c_1138_n 0.00536646f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_574 N_Y_M1023_d N_VGND_c_1138_n 0.00536646f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_575 N_Y_M1009_s N_VGND_c_1138_n 0.00536646f $X=2.27 $Y=0.235 $X2=0 $Y2=0
cc_576 N_Y_M1031_s N_VGND_c_1138_n 0.00380103f $X=3.13 $Y=0.235 $X2=0 $Y2=0
cc_577 N_Y_M1001_d N_VGND_c_1138_n 0.00380103f $X=4.1 $Y=0.235 $X2=0 $Y2=0
cc_578 N_Y_M1019_d N_VGND_c_1138_n 0.00380103f $X=4.96 $Y=0.235 $X2=0 $Y2=0
cc_579 N_Y_M1002_d N_VGND_c_1138_n 0.00225186f $X=6.44 $Y=0.235 $X2=0 $Y2=0
cc_580 N_Y_M1015_d N_VGND_c_1138_n 0.00225186f $X=7.3 $Y=0.235 $X2=0 $Y2=0
cc_581 N_Y_c_813_p N_VGND_c_1138_n 0.00730901f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_582 N_Y_c_811_p N_VGND_c_1138_n 0.00730901f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_583 N_Y_c_812_p N_VGND_c_1138_n 0.00730901f $X=2.41 $Y=0.42 $X2=0 $Y2=0
cc_584 N_Y_c_735_n N_VGND_c_1138_n 0.00950443f $X=3.27 $Y=0.42 $X2=0 $Y2=0
cc_585 N_Y_c_740_n N_VGND_c_1138_n 0.00916141f $X=4.24 $Y=0.42 $X2=0 $Y2=0
cc_586 N_Y_c_763_n N_VGND_c_1138_n 0.00950443f $X=5.1 $Y=0.42 $X2=0 $Y2=0
cc_587 N_Y_c_693_n N_A_1201_47#_M1002_s 0.00525829f $X=6.46 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_588 N_Y_c_772_n N_A_1201_47#_M1013_s 0.00329816f $X=7.31 $Y=0.955 $X2=0 $Y2=0
cc_589 N_Y_M1002_d N_A_1201_47#_c_1278_n 0.00332344f $X=6.44 $Y=0.235 $X2=0
+ $Y2=0
cc_590 N_Y_c_693_n N_A_1201_47#_c_1278_n 0.0046334f $X=6.46 $Y=0.955 $X2=0 $Y2=0
cc_591 N_Y_c_833_p N_A_1201_47#_c_1278_n 0.0122337f $X=6.58 $Y=0.76 $X2=0 $Y2=0
cc_592 N_Y_c_772_n N_A_1201_47#_c_1278_n 0.0046334f $X=7.31 $Y=0.955 $X2=0 $Y2=0
cc_593 N_Y_c_772_n N_A_1201_47#_c_1303_n 0.0130514f $X=7.31 $Y=0.955 $X2=0 $Y2=0
cc_594 N_Y_M1015_d N_A_1201_47#_c_1280_n 0.00332344f $X=7.3 $Y=0.235 $X2=0 $Y2=0
cc_595 N_Y_c_772_n N_A_1201_47#_c_1280_n 0.0046334f $X=7.31 $Y=0.955 $X2=0 $Y2=0
cc_596 N_Y_c_778_n N_A_1201_47#_c_1280_n 0.0138531f $X=7.44 $Y=0.76 $X2=0 $Y2=0
cc_597 N_Y_c_778_n N_A_1201_47#_c_1282_n 0.0230705f $X=7.44 $Y=0.76 $X2=0 $Y2=0
cc_598 N_Y_c_778_n N_A_1201_47#_c_1272_n 2.9127e-19 $X=7.44 $Y=0.76 $X2=0 $Y2=0
cc_599 N_Y_c_693_n N_A_1201_47#_c_1275_n 0.0211076f $X=6.46 $Y=0.955 $X2=0 $Y2=0
cc_600 N_A_454_367#_c_842_n N_A_819_367#_M1007_s 0.00479831f $X=4.555 $Y=2.015
+ $X2=-0.19 $Y2=1.655
cc_601 N_A_454_367#_c_857_n N_A_819_367#_M1011_s 0.00340761f $X=5.345 $Y=2.025
+ $X2=0 $Y2=0
cc_602 N_A_454_367#_c_842_n N_A_819_367#_c_893_n 0.0220026f $X=4.555 $Y=2.015
+ $X2=0 $Y2=0
cc_603 N_A_454_367#_M1007_d N_A_819_367#_c_907_n 0.00332344f $X=4.51 $Y=1.835
+ $X2=0 $Y2=0
cc_604 N_A_454_367#_c_861_n N_A_819_367#_c_907_n 0.0126348f $X=4.65 $Y=2.095
+ $X2=0 $Y2=0
cc_605 N_A_454_367#_c_857_n N_A_819_367#_c_954_n 0.0127742f $X=5.345 $Y=2.025
+ $X2=0 $Y2=0
cc_606 N_A_454_367#_M1033_d N_A_819_367#_c_910_n 0.00332344f $X=5.37 $Y=1.835
+ $X2=0 $Y2=0
cc_607 N_A_454_367#_c_863_n N_A_819_367#_c_910_n 0.0159805f $X=5.51 $Y=2.095
+ $X2=0 $Y2=0
cc_608 N_A_454_367#_M1006_d N_VPWR_c_988_n 0.00225186f $X=2.27 $Y=1.835 $X2=0
+ $Y2=0
cc_609 N_A_454_367#_M1030_d N_VPWR_c_988_n 0.00225186f $X=3.13 $Y=1.835 $X2=0
+ $Y2=0
cc_610 N_A_454_367#_M1007_d N_VPWR_c_988_n 0.00225186f $X=4.51 $Y=1.835 $X2=0
+ $Y2=0
cc_611 N_A_454_367#_M1033_d N_VPWR_c_988_n 0.00225186f $X=5.37 $Y=1.835 $X2=0
+ $Y2=0
cc_612 N_A_819_367#_c_934_n N_VPWR_M1012_d 0.00334931f $X=8.565 $Y=2.015 $X2=0
+ $Y2=0
cc_613 N_A_819_367#_c_902_n N_VPWR_M1036_d 0.00176461f $X=9.515 $Y=1.8 $X2=0
+ $Y2=0
cc_614 N_A_819_367#_c_889_n N_VPWR_c_989_n 0.0216087f $X=6.705 $Y=1.69 $X2=0
+ $Y2=0
cc_615 N_A_819_367#_c_891_n N_VPWR_c_990_n 0.021739f $X=7.565 $Y=1.69 $X2=0
+ $Y2=0
cc_616 N_A_819_367#_c_934_n N_VPWR_c_991_n 0.0170777f $X=8.565 $Y=2.015 $X2=0
+ $Y2=0
cc_617 N_A_819_367#_c_902_n N_VPWR_c_992_n 0.0170777f $X=9.515 $Y=1.8 $X2=0
+ $Y2=0
cc_618 N_A_819_367#_c_907_n N_VPWR_c_993_n 0.0319341f $X=4.955 $Y=2.99 $X2=0
+ $Y2=0
cc_619 N_A_819_367#_c_894_n N_VPWR_c_993_n 0.0211865f $X=4.385 $Y=2.99 $X2=0
+ $Y2=0
cc_620 N_A_819_367#_c_910_n N_VPWR_c_993_n 0.0361172f $X=5.845 $Y=2.99 $X2=0
+ $Y2=0
cc_621 N_A_819_367#_c_966_p N_VPWR_c_993_n 0.0125234f $X=5.94 $Y=2.905 $X2=0
+ $Y2=0
cc_622 N_A_819_367#_c_967_p N_VPWR_c_993_n 0.0135879f $X=5.065 $Y=2.99 $X2=0
+ $Y2=0
cc_623 N_A_819_367#_c_898_n N_VPWR_c_995_n 0.0124525f $X=6.8 $Y=1.98 $X2=0 $Y2=0
cc_624 N_A_819_367#_c_969_p N_VPWR_c_997_n 0.0215996f $X=7.73 $Y=2.475 $X2=0
+ $Y2=0
cc_625 N_A_819_367#_c_970_p N_VPWR_c_999_n 0.0187806f $X=8.705 $Y=2.455 $X2=0
+ $Y2=0
cc_626 N_A_819_367#_c_903_n N_VPWR_c_1001_n 0.0178111f $X=9.61 $Y=1.98 $X2=0
+ $Y2=0
cc_627 N_A_819_367#_M1007_s N_VPWR_c_988_n 0.00215158f $X=4.095 $Y=1.835 $X2=0
+ $Y2=0
cc_628 N_A_819_367#_M1011_s N_VPWR_c_988_n 0.00223563f $X=4.94 $Y=1.835 $X2=0
+ $Y2=0
cc_629 N_A_819_367#_M1035_s N_VPWR_c_988_n 0.00376627f $X=5.8 $Y=1.835 $X2=0
+ $Y2=0
cc_630 N_A_819_367#_M1020_d N_VPWR_c_988_n 0.00536646f $X=6.66 $Y=1.835 $X2=0
+ $Y2=0
cc_631 N_A_819_367#_M1028_d N_VPWR_c_988_n 0.00569199f $X=7.54 $Y=1.835 $X2=0
+ $Y2=0
cc_632 N_A_819_367#_M1017_s N_VPWR_c_988_n 0.00609022f $X=8.52 $Y=1.835 $X2=0
+ $Y2=0
cc_633 N_A_819_367#_M1037_s N_VPWR_c_988_n 0.00371702f $X=9.47 $Y=1.835 $X2=0
+ $Y2=0
cc_634 N_A_819_367#_c_907_n N_VPWR_c_988_n 0.0201012f $X=4.955 $Y=2.99 $X2=0
+ $Y2=0
cc_635 N_A_819_367#_c_894_n N_VPWR_c_988_n 0.0126421f $X=4.385 $Y=2.99 $X2=0
+ $Y2=0
cc_636 N_A_819_367#_c_910_n N_VPWR_c_988_n 0.023676f $X=5.845 $Y=2.99 $X2=0
+ $Y2=0
cc_637 N_A_819_367#_c_966_p N_VPWR_c_988_n 0.0073762f $X=5.94 $Y=2.905 $X2=0
+ $Y2=0
cc_638 N_A_819_367#_c_898_n N_VPWR_c_988_n 0.00730901f $X=6.8 $Y=1.98 $X2=0
+ $Y2=0
cc_639 N_A_819_367#_c_969_p N_VPWR_c_988_n 0.0127519f $X=7.73 $Y=2.475 $X2=0
+ $Y2=0
cc_640 N_A_819_367#_c_970_p N_VPWR_c_988_n 0.010808f $X=8.705 $Y=2.455 $X2=0
+ $Y2=0
cc_641 N_A_819_367#_c_903_n N_VPWR_c_988_n 0.0100304f $X=9.61 $Y=1.98 $X2=0
+ $Y2=0
cc_642 N_A_819_367#_c_967_p N_VPWR_c_988_n 0.00855309f $X=5.065 $Y=2.99 $X2=0
+ $Y2=0
cc_643 N_VGND_c_1138_n N_A_1201_47#_M1002_s 0.00231914f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_644 N_VGND_c_1138_n N_A_1201_47#_M1013_s 0.00225168f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_645 N_VGND_c_1138_n N_A_1201_47#_M1029_s 0.00453833f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_646 N_VGND_c_1138_n N_A_1201_47#_M1005_d 0.00536646f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_647 N_VGND_c_1138_n N_A_1201_47#_M1026_d 0.00371702f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_648 N_VGND_c_1136_n N_A_1201_47#_c_1278_n 0.0331715f $X=8.23 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1138_n N_A_1201_47#_c_1278_n 0.0206255f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_650 N_VGND_c_1136_n N_A_1201_47#_c_1280_n 0.0405913f $X=8.23 $Y=0 $X2=0 $Y2=0
cc_651 N_VGND_c_1138_n N_A_1201_47#_c_1280_n 0.0260732f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_c_1136_n N_A_1201_47#_c_1319_n 0.0129414f $X=8.23 $Y=0 $X2=0 $Y2=0
cc_653 N_VGND_c_1138_n N_A_1201_47#_c_1319_n 0.00738676f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_654 N_VGND_M1004_s N_A_1201_47#_c_1271_n 0.00176461f $X=8.255 $Y=0.235 $X2=0
+ $Y2=0
cc_655 N_VGND_c_1126_n N_A_1201_47#_c_1271_n 0.0170777f $X=8.395 $Y=0.38 $X2=0
+ $Y2=0
cc_656 N_VGND_c_1132_n N_A_1201_47#_c_1323_n 0.0124525f $X=9.09 $Y=0 $X2=0 $Y2=0
cc_657 N_VGND_c_1138_n N_A_1201_47#_c_1323_n 0.00730901f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_658 N_VGND_M1021_s N_A_1201_47#_c_1273_n 0.00176461f $X=9.115 $Y=0.235 $X2=0
+ $Y2=0
cc_659 N_VGND_c_1127_n N_A_1201_47#_c_1273_n 0.0170777f $X=9.255 $Y=0.38 $X2=0
+ $Y2=0
cc_660 N_VGND_c_1137_n N_A_1201_47#_c_1274_n 0.0178111f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_661 N_VGND_c_1138_n N_A_1201_47#_c_1274_n 0.0100304f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_662 N_VGND_c_1125_n N_A_1201_47#_c_1275_n 0.0262305f $X=5.53 $Y=0.565 $X2=0
+ $Y2=0
cc_663 N_VGND_c_1136_n N_A_1201_47#_c_1275_n 0.0202427f $X=8.23 $Y=0 $X2=0 $Y2=0
cc_664 N_VGND_c_1138_n N_A_1201_47#_c_1275_n 0.0124224f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1136_n N_A_1201_47#_c_1332_n 0.0148321f $X=8.23 $Y=0 $X2=0 $Y2=0
cc_666 N_VGND_c_1138_n N_A_1201_47#_c_1332_n 0.0101926f $X=9.84 $Y=0 $X2=0 $Y2=0
