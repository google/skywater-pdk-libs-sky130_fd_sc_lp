* NGSPICE file created from sky130_fd_sc_lp__a311o_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a311o_lp A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_257_414# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.6e+11p pd=5.12e+06u as=6.65e+11p ps=5.33e+06u
M1001 a_372_47# A2 a_294_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1002 a_85_21# A1 a_372_47# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1003 a_257_414# A3 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_294_47# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.793e+11p ps=3.01e+06u
M1005 VGND B1 a_536_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 VPWR a_85_21# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1007 VGND a_85_21# a_115_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1008 VPWR A2 a_257_414# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_85_21# C1 a_596_414# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=5.25e+11p ps=3.05e+06u
M1010 a_536_47# B1 a_85_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_596_414# B1 a_257_414# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_694_47# C1 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 a_85_21# C1 a_694_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_115_47# a_85_21# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

