# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o221ai_m
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o221ai_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535000 1.885000 3.205000 2.120000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.995000 1.795000 1.505000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895000 1.210000 1.285000 1.405000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 0.840000 2.905000 1.355000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.950000 0.835000 2.120000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.441250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.345000 0.555000 0.675000 ;
        RECT 0.155000 0.675000 0.325000 2.300000 ;
        RECT 0.155000 2.300000 1.925000 2.470000 ;
        RECT 0.155000 2.470000 0.490000 2.860000 ;
        RECT 1.715000 2.470000 1.925000 2.630000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.545000  0.860000 0.985000 1.030000 ;
      RECT 0.545000  1.030000 0.715000 1.585000 ;
      RECT 0.545000  1.585000 1.185000 1.685000 ;
      RECT 0.545000  1.685000 3.255000 1.705000 ;
      RECT 0.545000  1.705000 2.145000 1.755000 ;
      RECT 0.710000  2.650000 1.040000 3.245000 ;
      RECT 0.775000  0.345000 0.985000 0.860000 ;
      RECT 1.015000  1.755000 2.145000 1.855000 ;
      RECT 1.220000  0.345000 1.430000 0.645000 ;
      RECT 1.220000  0.645000 2.430000 0.660000 ;
      RECT 1.220000  0.660000 2.375000 0.815000 ;
      RECT 1.610000  0.085000 1.940000 0.465000 ;
      RECT 1.975000  1.535000 3.255000 1.685000 ;
      RECT 2.205000  0.330000 2.430000 0.645000 ;
      RECT 2.540000  2.485000 2.870000 3.245000 ;
      RECT 2.650000  0.330000 3.255000 0.660000 ;
      RECT 3.085000  0.660000 3.255000 1.535000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__o221ai_m
END LIBRARY
