* NGSPICE file created from sky130_fd_sc_lp__sregsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sregsbp_1 ASYNC CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_264_531# SCE VPWR VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.70875e+12p ps=2.163e+07u
M1001 VGND a_1273_393# a_1319_119# VNB nshort w=420000u l=150000u
+  ad=1.864e+12p pd=1.682e+07u as=8.82e+10p ps=1.26e+06u
M1002 a_1825_125# a_1273_393# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1003 a_2083_65# ASYNC a_2222_47# VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.344e+11p ps=1.7e+06u
M1004 VGND a_2083_65# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1005 VPWR CLK a_761_357# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.591e+11p ps=3.09e+06u
M1006 VGND a_2083_65# a_2035_91# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_2042_451# a_934_357# a_1903_125# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.856e+11p ps=2.47e+06u
M1008 VPWR a_2083_65# a_2042_451# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1139_463# a_934_357# a_342_531# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.373e+11p ps=2.81e+06u
M1010 a_1273_393# ASYNC a_1501_119# VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.536e+11p ps=1.76e+06u
M1011 VPWR a_2083_65# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.591e+11p ps=3.09e+06u
M1012 a_312_47# a_75_531# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1013 a_342_531# D a_312_47# VNB nshort w=420000u l=150000u
+  ad=2.583e+11p pd=2.91e+06u as=0p ps=0u
M1014 Q a_2456_451# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1015 a_2083_65# a_1903_125# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 Q a_2456_451# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1017 a_1225_463# a_761_357# a_1139_463# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_1831_373# a_1273_393# VPWR VPB phighvt w=840000u l=150000u
+  ad=3.276e+11p pd=2.76e+06u as=0p ps=0u
M1019 VPWR a_1139_463# a_1273_393# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=4.788e+11p ps=4.5e+06u
M1020 a_342_531# D a_264_531# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_2035_91# a_761_357# a_1903_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.515e+11p ps=2.64e+06u
M1022 a_75_531# SCE VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1023 a_2456_451# a_2083_65# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1024 a_486_47# SCE a_342_531# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1025 VGND SCD a_486_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_2456_451# a_2083_65# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1027 a_1903_125# a_934_357# a_1825_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR SCD a_428_531# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.596e+11p ps=1.6e+06u
M1029 a_934_357# a_761_357# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1030 a_428_531# a_75_531# a_342_531# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_636_531# a_342_531# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1032 a_1139_463# a_761_357# a_342_531# VNB nshort w=420000u l=150000u
+  ad=1.827e+11p pd=1.71e+06u as=0p ps=0u
M1033 VPWR a_1273_393# a_1225_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1273_393# ASYNC VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR ASYNC a_2083_65# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_636_531# a_342_531# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1037 a_1319_119# a_934_357# a_1139_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1501_119# a_1139_463# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND CLK a_761_357# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1040 a_2222_47# a_1903_125# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR SCE a_75_531# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1042 a_1903_125# a_761_357# a_1831_373# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_934_357# a_761_357# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
.ends

