* File: sky130_fd_sc_lp__or3_m.spice
* Created: Fri Aug 28 11:23:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3_m.pex.spice"
.subckt sky130_fd_sc_lp__or3_m  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_C_M1002_g N_A_43_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1386 AS=0.1113 PD=1.08 PS=1.37 NRD=108.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1001 N_A_43_47#_M1001_d N_B_M1001_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1386 PD=0.7 PS=1.08 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_43_47#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_43_47#_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=11.424 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_216_397# N_C_M1005_g N_A_43_47#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 A_288_397# N_B_M1007_g A_216_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_288_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=14.0658 NRS=23.443 M=1 R=2.8 SA=75000.9
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_43_47#_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=37.5088 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__or3_m.pxi.spice"
*
.ends
*
*
