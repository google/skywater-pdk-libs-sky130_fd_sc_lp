* File: sky130_fd_sc_lp__dfxbp_1.spice
* Created: Wed Sep  2 09:44:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfxbp_1.pex.spice"
.subckt sky130_fd_sc_lp__dfxbp_1  VNB VPB CLK D VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1004 N_A_110_82#_M1004_d N_CLK_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1113 PD=1.41 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_110_82#_M1008_g N_A_217_463#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1365 AS=0.1113 PD=1.07 PS=1.37 NRD=47.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75005.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_440_463#_M1022_d N_D_M1022_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1365 PD=0.7 PS=1.07 NRD=0 NRS=58.56 M=1 R=2.8 SA=75001
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1010 N_A_526_463#_M1010_d N_A_110_82#_M1010_g N_A_440_463#_M1022_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1014 A_655_119# N_A_217_463#_M1014_g N_A_526_463#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_697_93#_M1005_g A_655_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.13543 AS=0.0441 PD=1.04208 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1024 N_A_697_93#_M1024_d N_A_526_463#_M1024_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.64 AD=0.130294 AS=0.20637 PD=1.22566 PS=1.58792 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1018 N_A_997_119#_M1018_d N_A_217_463#_M1018_g N_A_697_93#_M1024_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0819 AS=0.0855057 PD=0.81 PS=0.80434 NRD=14.28 NRS=27.852
+ M=1 R=2.8 SA=75003.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 A_1105_119# N_A_110_82#_M1000_g N_A_997_119#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0462 AS=0.0819 PD=0.64 PS=0.81 NRD=15.708 NRS=17.136 M=1 R=2.8
+ SA=75004.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_1149_93#_M1009_g A_1105_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.119938 AS=0.0462 PD=0.935094 PS=0.64 NRD=52.14 NRS=15.708 M=1 R=2.8
+ SA=75004.5 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1006 N_A_1149_93#_M1006_d N_A_997_119#_M1006_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.182762 PD=1.81 PS=1.42491 NRD=0 NRS=14.988 M=1
+ R=4.26667 SA=75003.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_A_1149_93#_M1011_g N_A_1401_22#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0952 AS=0.1113 PD=0.823333 PS=1.37 NRD=21.42 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_Q_N_M1012_d N_A_1401_22#_M1012_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1904 PD=2.21 PS=1.64667 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_Q_M1015_d N_A_1149_93#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1026 N_A_110_82#_M1026_d N_CLK_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A_110_82#_M1002_g N_A_217_463#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.177328 AS=0.1696 PD=1.43698 PS=1.81 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1023 N_A_440_463#_M1023_d N_D_M1023_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.116372 PD=0.7 PS=0.943019 NRD=0 NRS=104.154 M=1 R=2.8
+ SA=75000.9 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1027 N_A_526_463#_M1027_d N_A_217_463#_M1027_g N_A_440_463#_M1023_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1212 AS=0.0588 PD=1.07 PS=0.7 NRD=44.5417 NRS=0 M=1
+ R=2.8 SA=75001.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1016 A_650_499# N_A_110_82#_M1016_g N_A_526_463#_M1027_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0882 AS=0.1212 PD=0.96 PS=1.07 NRD=72.693 NRS=46.886 M=1 R=2.8
+ SA=75001.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_697_93#_M1001_g A_650_499# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.144167 AS=0.0882 PD=1.1 PS=0.96 NRD=135.201 NRS=72.693 M=1 R=2.8
+ SA=75001.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_697_93#_M1013_d N_A_526_463#_M1013_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.231 AS=0.288333 PD=1.39 PS=2.2 NRD=0 NRS=67.5907 M=1 R=5.6
+ SA=75001.2 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1025 N_A_997_119#_M1025_d N_A_110_82#_M1025_g N_A_697_93#_M1013_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1792 AS=0.231 PD=1.62 PS=1.39 NRD=0 NRS=63.3158 M=1 R=5.6
+ SA=75001.9 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1019 A_1137_379# N_A_217_463#_M1019_g N_A_997_119#_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=44.5417 M=1 R=2.8
+ SA=75001.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_1149_93#_M1003_g A_1137_379# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0917 AS=0.0441 PD=0.82 PS=0.63 NRD=28.1316 NRS=23.443 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1020 N_A_1149_93#_M1020_d N_A_997_119#_M1020_g N_VPWR_M1003_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1834 PD=2.21 PS=1.64 NRD=0 NRS=5.8509 M=1 R=5.6
+ SA=75001.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_VPWR_M1021_d N_A_1149_93#_M1021_g N_A_1401_22#_M1021_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.136185 AS=0.1696 PD=1.10147 PS=1.81 NRD=48.5605 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1007 N_Q_N_M1007_d N_A_1401_22#_M1007_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.268115 PD=3.05 PS=2.16853 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1017 N_Q_M1017_d N_A_1149_93#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.6127 P=23.69
c_94 VNB 0 6.36774e-20 $X=0 $Y=0
c_180 VPB 0 4.113e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dfxbp_1.pxi.spice"
*
.ends
*
*
