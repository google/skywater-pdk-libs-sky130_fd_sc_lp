* File: sky130_fd_sc_lp__and3b_2.pxi.spice
* Created: Fri Aug 28 10:06:44 2020
* 
x_PM_SKY130_FD_SC_LP__AND3B_2%A_N N_A_N_M1005_g N_A_N_M1008_g A_N A_N
+ N_A_N_c_67_n N_A_N_c_68_n PM_SKY130_FD_SC_LP__AND3B_2%A_N
x_PM_SKY130_FD_SC_LP__AND3B_2%A_204_27# N_A_204_27#_M1007_d N_A_204_27#_M1000_d
+ N_A_204_27#_M1002_d N_A_204_27#_M1009_g N_A_204_27#_M1001_g
+ N_A_204_27#_M1010_g N_A_204_27#_M1011_g N_A_204_27#_c_96_n N_A_204_27#_c_97_n
+ N_A_204_27#_c_98_n N_A_204_27#_c_105_n N_A_204_27#_c_106_n N_A_204_27#_c_107_n
+ N_A_204_27#_c_99_n N_A_204_27#_c_108_n N_A_204_27#_c_100_n N_A_204_27#_c_110_n
+ N_A_204_27#_c_101_n PM_SKY130_FD_SC_LP__AND3B_2%A_204_27#
x_PM_SKY130_FD_SC_LP__AND3B_2%C N_C_M1000_g N_C_M1003_g C N_C_c_179_n
+ N_C_c_180_n N_C_c_181_n PM_SKY130_FD_SC_LP__AND3B_2%C
x_PM_SKY130_FD_SC_LP__AND3B_2%B N_B_M1006_g N_B_M1004_g B B N_B_c_213_n
+ N_B_c_214_n PM_SKY130_FD_SC_LP__AND3B_2%B
x_PM_SKY130_FD_SC_LP__AND3B_2%A_27_137# N_A_27_137#_M1005_s N_A_27_137#_M1008_s
+ N_A_27_137#_M1007_g N_A_27_137#_M1002_g N_A_27_137#_c_247_n
+ N_A_27_137#_c_248_n N_A_27_137#_c_249_n N_A_27_137#_c_272_n
+ N_A_27_137#_c_250_n N_A_27_137#_c_256_n N_A_27_137#_c_251_n
+ N_A_27_137#_c_252_n N_A_27_137#_c_253_n PM_SKY130_FD_SC_LP__AND3B_2%A_27_137#
x_PM_SKY130_FD_SC_LP__AND3B_2%VPWR N_VPWR_M1008_d N_VPWR_M1011_d N_VPWR_M1004_d
+ N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n VPWR
+ N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_316_n N_VPWR_c_324_n N_VPWR_c_325_n
+ N_VPWR_c_326_n PM_SKY130_FD_SC_LP__AND3B_2%VPWR
x_PM_SKY130_FD_SC_LP__AND3B_2%X N_X_M1009_d N_X_M1001_s X X X X X N_X_c_350_n
+ PM_SKY130_FD_SC_LP__AND3B_2%X
x_PM_SKY130_FD_SC_LP__AND3B_2%VGND N_VGND_M1005_d N_VGND_M1010_s N_VGND_c_370_n
+ N_VGND_c_371_n VGND N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n
+ N_VGND_c_375_n PM_SKY130_FD_SC_LP__AND3B_2%VGND
cc_1 VNB N_A_N_M1008_g 0.00607065f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.045
cc_2 VNB A_N 0.00821029f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_67_n 0.0361605f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.38
cc_4 VNB N_A_N_c_68_n 0.0192586f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.215
cc_5 VNB N_A_204_27#_M1009_g 0.0314456f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.38
cc_6 VNB N_A_204_27#_M1001_g 0.00151548f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.545
cc_7 VNB N_A_204_27#_M1010_g 0.0241405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_204_27#_M1011_g 0.00168812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_204_27#_c_96_n 0.00565983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_204_27#_c_97_n 0.0034009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_204_27#_c_98_n 0.0427295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_204_27#_c_99_n 0.042938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_204_27#_c_100_n 0.00135772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_204_27#_c_101_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C_M1000_g 0.00650873f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.895
cc_16 VNB N_C_c_179_n 0.030727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_c_180_n 0.00704771f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.38
cc_18 VNB N_C_c_181_n 0.0170007f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.38
cc_19 VNB N_B_M1004_g 0.00624219f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.045
cc_20 VNB B 0.0106641f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_21 VNB N_B_c_213_n 0.0287671f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.38
cc_22 VNB N_B_c_214_n 0.0148077f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.215
cc_23 VNB N_A_27_137#_M1007_g 0.01482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_137#_M1002_g 0.0156119f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.38
cc_25 VNB N_A_27_137#_c_247_n 0.00933124f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.545
cc_26 VNB N_A_27_137#_c_248_n 0.0298368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_137#_c_249_n 0.0125711f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.665
cc_28 VNB N_A_27_137#_c_250_n 0.0234584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_137#_c_251_n 0.00255626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_137#_c_252_n 0.0222427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_137#_c_253_n 0.0472449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_316_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_370_n 0.0167433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_371_n 0.0196181f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_35 VNB N_VGND_c_372_n 0.0191092f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.545
cc_36 VNB N_VGND_c_373_n 0.0503259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_374_n 0.23589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_375_n 0.0169876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_N_M1008_g 0.0299267f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.045
cc_40 VPB A_N 0.00509921f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_41 VPB N_A_204_27#_M1001_g 0.0227463f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.545
cc_42 VPB N_A_204_27#_M1011_g 0.0237715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_204_27#_c_97_n 0.00106735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_204_27#_c_105_n 0.00698625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_204_27#_c_106_n 9.25944e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_204_27#_c_107_n 0.00877719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_204_27#_c_108_n 0.0152238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_204_27#_c_100_n 0.00580392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_204_27#_c_110_n 0.00805403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_C_M1000_g 0.0269322f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.895
cc_51 VPB N_B_M1004_g 0.0239158f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.045
cc_52 VPB N_A_27_137#_M1002_g 0.0301547f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.38
cc_53 VPB N_A_27_137#_c_248_n 0.0131866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_27_137#_c_256_n 0.0150746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_317_n 0.0345324f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.38
cc_56 VPB N_VPWR_c_318_n 0.0186115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_319_n 0.0337645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_320_n 0.0707922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_321_n 0.0308037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_322_n 0.0217138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_316_n 0.12861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_324_n 0.0285356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_325_n 0.00535651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_326_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 A_N N_A_204_27#_M1009_g 0.00460341f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A_N_c_67_n N_A_204_27#_M1009_g 0.0146649f $X=0.59 $Y=1.38 $X2=0 $Y2=0
cc_67 N_A_N_c_68_n N_A_204_27#_M1009_g 0.0152427f $X=0.577 $Y=1.215 $X2=0 $Y2=0
cc_68 N_A_N_M1008_g N_A_204_27#_c_96_n 0.0144444f $X=0.535 $Y=2.045 $X2=0 $Y2=0
cc_69 N_A_N_M1008_g N_A_27_137#_c_248_n 0.00901421f $X=0.535 $Y=2.045 $X2=0
+ $Y2=0
cc_70 A_N N_A_27_137#_c_248_n 0.0411522f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_N_c_68_n N_A_27_137#_c_248_n 0.0143426f $X=0.577 $Y=1.215 $X2=0 $Y2=0
cc_72 N_A_N_c_68_n N_A_27_137#_c_250_n 0.0120797f $X=0.577 $Y=1.215 $X2=0 $Y2=0
cc_73 N_A_N_M1008_g N_A_27_137#_c_256_n 0.00487555f $X=0.535 $Y=2.045 $X2=0
+ $Y2=0
cc_74 N_A_N_c_67_n N_A_27_137#_c_256_n 0.00120052f $X=0.59 $Y=1.38 $X2=0 $Y2=0
cc_75 A_N N_A_27_137#_c_251_n 0.0144571f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_N_c_67_n N_A_27_137#_c_251_n 9.28324e-19 $X=0.59 $Y=1.38 $X2=0 $Y2=0
cc_77 N_A_N_c_68_n N_A_27_137#_c_251_n 0.0114782f $X=0.577 $Y=1.215 $X2=0 $Y2=0
cc_78 N_A_N_M1008_g N_VPWR_c_317_n 0.00367322f $X=0.535 $Y=2.045 $X2=0 $Y2=0
cc_79 A_N N_VPWR_c_317_n 0.0232947f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A_N_c_67_n N_VPWR_c_317_n 4.57668e-19 $X=0.59 $Y=1.38 $X2=0 $Y2=0
cc_81 N_A_N_M1008_g N_X_c_350_n 0.00100129f $X=0.535 $Y=2.045 $X2=0 $Y2=0
cc_82 A_N N_X_c_350_n 0.0401797f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_N_c_67_n N_X_c_350_n 2.77461e-19 $X=0.59 $Y=1.38 $X2=0 $Y2=0
cc_84 N_A_N_c_68_n N_X_c_350_n 0.00151683f $X=0.577 $Y=1.215 $X2=0 $Y2=0
cc_85 N_A_N_c_68_n N_VGND_c_372_n 6.44673e-19 $X=0.577 $Y=1.215 $X2=0 $Y2=0
cc_86 N_A_204_27#_M1011_g N_C_M1000_g 0.00780503f $X=1.525 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_204_27#_c_97_n N_C_M1000_g 0.00206816f $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_88 N_A_204_27#_c_98_n N_C_M1000_g 0.00306095f $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_89 N_A_204_27#_c_105_n N_C_M1000_g 0.0148173f $X=2.405 $Y=1.82 $X2=0 $Y2=0
cc_90 N_A_204_27#_c_100_n N_C_M1000_g 0.0152807f $X=2.56 $Y=1.82 $X2=0 $Y2=0
cc_91 N_A_204_27#_M1010_g N_C_c_179_n 0.00140984f $X=1.525 $Y=0.685 $X2=0 $Y2=0
cc_92 N_A_204_27#_c_97_n N_C_c_179_n 2.40702e-19 $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_93 N_A_204_27#_c_98_n N_C_c_179_n 0.0160603f $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_94 N_A_204_27#_c_105_n N_C_c_179_n 0.00371746f $X=2.405 $Y=1.82 $X2=0 $Y2=0
cc_95 N_A_204_27#_c_100_n N_C_c_179_n 6.94505e-19 $X=2.56 $Y=1.82 $X2=0 $Y2=0
cc_96 N_A_204_27#_M1010_g N_C_c_180_n 0.00141685f $X=1.525 $Y=0.685 $X2=0 $Y2=0
cc_97 N_A_204_27#_c_97_n N_C_c_180_n 0.0192198f $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_98 N_A_204_27#_c_98_n N_C_c_180_n 0.00164917f $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_99 N_A_204_27#_c_105_n N_C_c_180_n 0.0264819f $X=2.405 $Y=1.82 $X2=0 $Y2=0
cc_100 N_A_204_27#_M1010_g N_C_c_181_n 0.00952856f $X=1.525 $Y=0.685 $X2=0 $Y2=0
cc_101 N_A_204_27#_c_107_n N_B_M1004_g 0.0127377f $X=3.4 $Y=1.74 $X2=0 $Y2=0
cc_102 N_A_204_27#_c_100_n N_B_M1004_g 0.00718378f $X=2.56 $Y=1.82 $X2=0 $Y2=0
cc_103 N_A_204_27#_c_107_n B 0.0393271f $X=3.4 $Y=1.74 $X2=0 $Y2=0
cc_104 N_A_204_27#_c_99_n B 0.0291415f $X=3.505 $Y=0.895 $X2=0 $Y2=0
cc_105 N_A_204_27#_c_100_n B 0.015286f $X=2.56 $Y=1.82 $X2=0 $Y2=0
cc_106 N_A_204_27#_c_107_n N_B_c_213_n 0.0030082f $X=3.4 $Y=1.74 $X2=0 $Y2=0
cc_107 N_A_204_27#_c_100_n N_B_c_213_n 0.0015978f $X=2.56 $Y=1.82 $X2=0 $Y2=0
cc_108 N_A_204_27#_c_99_n N_A_27_137#_M1007_g 0.00318013f $X=3.505 $Y=0.895
+ $X2=0 $Y2=0
cc_109 N_A_204_27#_c_107_n N_A_27_137#_M1002_g 0.0208768f $X=3.4 $Y=1.74 $X2=0
+ $Y2=0
cc_110 N_A_204_27#_c_108_n N_A_27_137#_M1002_g 4.71016e-19 $X=3.515 $Y=2.035
+ $X2=0 $Y2=0
cc_111 N_A_204_27#_c_100_n N_A_27_137#_M1002_g 6.30804e-19 $X=2.56 $Y=1.82 $X2=0
+ $Y2=0
cc_112 N_A_204_27#_c_99_n N_A_27_137#_c_247_n 0.0135423f $X=3.505 $Y=0.895 $X2=0
+ $Y2=0
cc_113 N_A_204_27#_c_98_n N_A_27_137#_c_249_n 0.00157216f $X=1.74 $Y=1.46 $X2=0
+ $Y2=0
cc_114 N_A_204_27#_c_97_n N_A_27_137#_c_272_n 0.00811825f $X=1.74 $Y=1.46 $X2=0
+ $Y2=0
cc_115 N_A_204_27#_c_98_n N_A_27_137#_c_272_n 0.00125237f $X=1.74 $Y=1.46 $X2=0
+ $Y2=0
cc_116 N_A_204_27#_M1009_g N_A_27_137#_c_250_n 0.00153848f $X=1.095 $Y=0.685
+ $X2=0 $Y2=0
cc_117 N_A_204_27#_M1009_g N_A_27_137#_c_251_n 0.0152237f $X=1.095 $Y=0.685
+ $X2=0 $Y2=0
cc_118 N_A_204_27#_M1010_g N_A_27_137#_c_251_n 0.0167292f $X=1.525 $Y=0.685
+ $X2=0 $Y2=0
cc_119 N_A_204_27#_c_105_n N_VPWR_M1011_d 0.0136337f $X=2.405 $Y=1.82 $X2=0
+ $Y2=0
cc_120 N_A_204_27#_c_106_n N_VPWR_M1011_d 0.00316132f $X=1.855 $Y=1.82 $X2=0
+ $Y2=0
cc_121 N_A_204_27#_M1001_g N_VPWR_c_317_n 0.0112428f $X=1.095 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_204_27#_M1001_g N_VPWR_c_318_n 0.00503406f $X=1.095 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_204_27#_M1011_g N_VPWR_c_318_n 0.0054895f $X=1.525 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_204_27#_M1011_g N_VPWR_c_319_n 0.0046137f $X=1.525 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_204_27#_c_98_n N_VPWR_c_319_n 9.46278e-19 $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_126 N_A_204_27#_c_105_n N_VPWR_c_319_n 0.00565709f $X=2.405 $Y=1.82 $X2=0
+ $Y2=0
cc_127 N_A_204_27#_c_106_n N_VPWR_c_319_n 0.017752f $X=1.855 $Y=1.82 $X2=0 $Y2=0
cc_128 N_A_204_27#_c_100_n N_VPWR_c_319_n 0.00359104f $X=2.56 $Y=1.82 $X2=0
+ $Y2=0
cc_129 N_A_204_27#_c_107_n N_VPWR_c_320_n 0.0236663f $X=3.4 $Y=1.74 $X2=0 $Y2=0
cc_130 N_A_204_27#_M1001_g N_VPWR_c_316_n 0.0100356f $X=1.095 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_204_27#_M1011_g N_VPWR_c_316_n 0.0110654f $X=1.525 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_204_27#_M1009_g N_X_c_350_n 0.0161835f $X=1.095 $Y=0.685 $X2=0 $Y2=0
cc_133 N_A_204_27#_M1001_g N_X_c_350_n 0.0246882f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_204_27#_M1010_g N_X_c_350_n 0.0165159f $X=1.525 $Y=0.685 $X2=0 $Y2=0
cc_135 N_A_204_27#_M1011_g N_X_c_350_n 0.0255656f $X=1.525 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_204_27#_c_96_n N_X_c_350_n 0.00193569f $X=1.095 $Y=1.55 $X2=0 $Y2=0
cc_137 N_A_204_27#_c_97_n N_X_c_350_n 0.0309436f $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_138 N_A_204_27#_c_98_n N_X_c_350_n 0.00746429f $X=1.74 $Y=1.46 $X2=0 $Y2=0
cc_139 N_A_204_27#_c_106_n N_X_c_350_n 0.013571f $X=1.855 $Y=1.82 $X2=0 $Y2=0
cc_140 N_A_204_27#_c_101_n N_X_c_350_n 0.00865625f $X=1.45 $Y=1.46 $X2=0 $Y2=0
cc_141 N_A_204_27#_M1010_g N_VGND_c_370_n 0.00884127f $X=1.525 $Y=0.685 $X2=0
+ $Y2=0
cc_142 N_A_204_27#_M1009_g N_VGND_c_371_n 0.00387708f $X=1.095 $Y=0.685 $X2=0
+ $Y2=0
cc_143 N_A_204_27#_M1010_g N_VGND_c_371_n 0.00387708f $X=1.525 $Y=0.685 $X2=0
+ $Y2=0
cc_144 N_A_204_27#_c_99_n N_VGND_c_373_n 0.00428109f $X=3.505 $Y=0.895 $X2=0
+ $Y2=0
cc_145 N_A_204_27#_M1009_g N_VGND_c_374_n 0.00650542f $X=1.095 $Y=0.685 $X2=0
+ $Y2=0
cc_146 N_A_204_27#_M1010_g N_VGND_c_374_n 0.00656008f $X=1.525 $Y=0.685 $X2=0
+ $Y2=0
cc_147 N_A_204_27#_c_99_n N_VGND_c_374_n 0.00757309f $X=3.505 $Y=0.895 $X2=0
+ $Y2=0
cc_148 N_A_204_27#_M1009_g N_VGND_c_375_n 0.00908632f $X=1.095 $Y=0.685 $X2=0
+ $Y2=0
cc_149 N_C_M1000_g N_B_M1004_g 0.0207358f $X=2.355 $Y=2.045 $X2=0 $Y2=0
cc_150 N_C_c_180_n B 0.0299888f $X=2.28 $Y=1.38 $X2=0 $Y2=0
cc_151 N_C_c_181_n B 0.00247611f $X=2.28 $Y=1.215 $X2=0 $Y2=0
cc_152 N_C_c_179_n N_B_c_213_n 0.0315823f $X=2.28 $Y=1.38 $X2=0 $Y2=0
cc_153 N_C_c_180_n N_B_c_213_n 3.55724e-19 $X=2.28 $Y=1.38 $X2=0 $Y2=0
cc_154 N_C_c_180_n N_B_c_214_n 3.07604e-19 $X=2.28 $Y=1.38 $X2=0 $Y2=0
cc_155 N_C_c_181_n N_B_c_214_n 0.0315823f $X=2.28 $Y=1.215 $X2=0 $Y2=0
cc_156 N_C_c_179_n N_A_27_137#_c_249_n 8.83138e-19 $X=2.28 $Y=1.38 $X2=0 $Y2=0
cc_157 N_C_c_180_n N_A_27_137#_c_249_n 0.0186953f $X=2.28 $Y=1.38 $X2=0 $Y2=0
cc_158 N_C_c_181_n N_A_27_137#_c_249_n 0.0207968f $X=2.28 $Y=1.215 $X2=0 $Y2=0
cc_159 N_C_M1000_g N_VPWR_c_319_n 0.00488195f $X=2.355 $Y=2.045 $X2=0 $Y2=0
cc_160 N_C_c_180_n N_X_c_350_n 0.00540608f $X=2.28 $Y=1.38 $X2=0 $Y2=0
cc_161 N_C_c_181_n N_VGND_c_373_n 6.49089e-19 $X=2.28 $Y=1.215 $X2=0 $Y2=0
cc_162 B N_A_27_137#_M1007_g 0.00282055f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_163 N_B_c_214_n N_A_27_137#_M1007_g 0.0194762f $X=2.82 $Y=1.215 $X2=0 $Y2=0
cc_164 N_B_M1004_g N_A_27_137#_M1002_g 0.0192878f $X=2.785 $Y=2.045 $X2=0 $Y2=0
cc_165 B N_A_27_137#_M1002_g 0.00238178f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B_c_213_n N_A_27_137#_M1002_g 0.0099726f $X=2.82 $Y=1.38 $X2=0 $Y2=0
cc_167 B N_A_27_137#_c_247_n 0.00366582f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_168 N_B_c_213_n N_A_27_137#_c_247_n 0.00970271f $X=2.82 $Y=1.38 $X2=0 $Y2=0
cc_169 B N_A_27_137#_c_249_n 0.0264975f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_170 N_B_c_213_n N_A_27_137#_c_249_n 8.80764e-19 $X=2.82 $Y=1.38 $X2=0 $Y2=0
cc_171 N_B_c_214_n N_A_27_137#_c_249_n 0.0166202f $X=2.82 $Y=1.215 $X2=0 $Y2=0
cc_172 B N_A_27_137#_c_252_n 0.00969428f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 B N_A_27_137#_c_253_n 5.96983e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_174 N_B_c_214_n N_A_27_137#_c_253_n 0.00109563f $X=2.82 $Y=1.215 $X2=0 $Y2=0
cc_175 N_B_M1004_g N_VPWR_c_320_n 0.00517002f $X=2.785 $Y=2.045 $X2=0 $Y2=0
cc_176 N_B_c_214_n N_VGND_c_373_n 6.49089e-19 $X=2.82 $Y=1.215 $X2=0 $Y2=0
cc_177 N_A_27_137#_M1002_g N_VPWR_c_320_n 0.0039037f $X=3.3 $Y=2.045 $X2=0 $Y2=0
cc_178 N_A_27_137#_c_251_n N_X_M1009_d 0.0043453f $X=1.645 $Y=0.707 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_27_137#_c_251_n N_X_c_350_n 0.0193629f $X=1.645 $Y=0.707 $X2=0 $Y2=0
cc_180 N_A_27_137#_c_251_n N_VGND_M1005_d 0.0109834f $X=1.645 $Y=0.707 $X2=-0.19
+ $Y2=-0.245
cc_181 N_A_27_137#_c_249_n N_VGND_M1010_s 0.0154775f $X=3.045 $Y=0.707 $X2=0
+ $Y2=0
cc_182 N_A_27_137#_c_272_n N_VGND_M1010_s 0.00429335f $X=1.807 $Y=0.707 $X2=0
+ $Y2=0
cc_183 N_A_27_137#_c_272_n N_VGND_c_370_n 0.0253077f $X=1.807 $Y=0.707 $X2=0
+ $Y2=0
cc_184 N_A_27_137#_c_251_n N_VGND_c_371_n 0.0135517f $X=1.645 $Y=0.707 $X2=0
+ $Y2=0
cc_185 N_A_27_137#_c_250_n N_VGND_c_372_n 0.00805322f $X=0.26 $Y=0.63 $X2=0
+ $Y2=0
cc_186 N_A_27_137#_c_251_n N_VGND_c_372_n 0.00435866f $X=1.645 $Y=0.707 $X2=0
+ $Y2=0
cc_187 N_A_27_137#_c_249_n N_VGND_c_373_n 0.0239469f $X=3.045 $Y=0.707 $X2=0
+ $Y2=0
cc_188 N_A_27_137#_c_252_n N_VGND_c_373_n 0.0218606f $X=3.21 $Y=0.41 $X2=0 $Y2=0
cc_189 N_A_27_137#_c_253_n N_VGND_c_373_n 0.00578905f $X=3.21 $Y=0.41 $X2=0
+ $Y2=0
cc_190 N_A_27_137#_c_249_n N_VGND_c_374_n 0.032215f $X=3.045 $Y=0.707 $X2=0
+ $Y2=0
cc_191 N_A_27_137#_c_272_n N_VGND_c_374_n 0.00185211f $X=1.807 $Y=0.707 $X2=0
+ $Y2=0
cc_192 N_A_27_137#_c_250_n N_VGND_c_374_n 0.0105845f $X=0.26 $Y=0.63 $X2=0 $Y2=0
cc_193 N_A_27_137#_c_251_n N_VGND_c_374_n 0.0290646f $X=1.645 $Y=0.707 $X2=0
+ $Y2=0
cc_194 N_A_27_137#_c_252_n N_VGND_c_374_n 0.0111921f $X=3.21 $Y=0.41 $X2=0 $Y2=0
cc_195 N_A_27_137#_c_253_n N_VGND_c_374_n 0.0112336f $X=3.21 $Y=0.41 $X2=0 $Y2=0
cc_196 N_A_27_137#_c_251_n N_VGND_c_375_n 0.0243422f $X=1.645 $Y=0.707 $X2=0
+ $Y2=0
cc_197 N_A_27_137#_c_249_n A_489_137# 0.00219103f $X=3.045 $Y=0.707 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_27_137#_c_249_n A_561_137# 0.00230327f $X=3.045 $Y=0.707 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_27_137#_c_252_n A_561_137# 0.00124702f $X=3.21 $Y=0.41 $X2=-0.19
+ $Y2=-0.245
cc_200 N_VPWR_c_316_n N_X_M1001_s 0.00223559f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_317_n N_X_c_350_n 0.088579f $X=0.75 $Y=2.095 $X2=0 $Y2=0
cc_202 N_VPWR_c_318_n N_X_c_350_n 0.0209688f $X=1.645 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_316_n N_X_c_350_n 0.013415f $X=3.6 $Y=3.33 $X2=0 $Y2=0
