* File: sky130_fd_sc_lp__nand3b_m.pex.spice
* Created: Wed Sep  2 10:05:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3B_M%A_N 3 7 11 12 13 14 15 20
r42 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.545
+ $Y=1.005 $X2=0.545 $Y2=1.005
r43 14 15 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.632 $Y=1.295
+ $X2=0.632 $Y2=1.665
r44 14 21 9.6872 $w=3.43e-07 $l=2.9e-07 $layer=LI1_cond $X=0.632 $Y=1.295
+ $X2=0.632 $Y2=1.005
r45 13 21 2.67233 $w=3.43e-07 $l=8e-08 $layer=LI1_cond $X=0.632 $Y=0.925
+ $X2=0.632 $Y2=1.005
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.545 $Y=1.345
+ $X2=0.545 $Y2=1.005
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.345
+ $X2=0.545 $Y2=1.51
r48 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=0.84
+ $X2=0.545 $Y2=1.005
r49 7 12 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.635 $Y=2.165
+ $X2=0.635 $Y2=1.51
r50 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.525 $Y=0.445
+ $X2=0.525 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_M%C 3 7 9 10 11 12 13 14 19
c42 9 0 7.5703e-20 $X=1.09 $Y=0.765
c43 3 0 9.76249e-20 $X=1.065 $Y=2.165
r44 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09
+ $Y=0.93 $X2=1.09 $Y2=0.93
r45 14 20 15.0229 $w=2.78e-07 $l=3.65e-07 $layer=LI1_cond $X=1.145 $Y=1.295
+ $X2=1.145 $Y2=0.93
r46 13 20 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=1.145 $Y=0.925
+ $X2=1.145 $Y2=0.93
r47 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.145 $Y=0.555
+ $X2=1.145 $Y2=0.925
r48 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.09 $Y=1.27
+ $X2=1.09 $Y2=0.93
r49 10 11 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.27
+ $X2=1.09 $Y2=1.435
r50 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=0.765
+ $X2=1.09 $Y2=0.93
r51 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.18 $Y=0.445 $X2=1.18
+ $Y2=0.765
r52 3 11 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.065 $Y=2.165
+ $X2=1.065 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_M%B 3 7 11 12 13 14 15 20
r39 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.29
+ $X2=1.63 $Y2=1.455
r40 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.29
+ $X2=1.63 $Y2=1.125
r41 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.29 $X2=1.63 $Y2=1.29
r42 14 15 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.63 $Y=0.925
+ $X2=1.63 $Y2=1.29
r43 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=0.555
+ $X2=1.63 $Y2=0.925
r44 11 12 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=1.517 $Y=1.675
+ $X2=1.517 $Y2=1.825
r45 11 23 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.54 $Y=1.675
+ $X2=1.54 $Y2=1.455
r46 7 22 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.54 $Y=0.445
+ $X2=1.54 $Y2=1.125
r47 3 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.495 $Y=2.165
+ $X2=1.495 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_M%A_37_47# 1 2 7 9 11 15 17 20 24 33 36 37 40
+ 41 42
c67 42 0 9.76249e-20 $X=0.477 $Y=2.715
c68 33 0 7.5703e-20 $X=0.31 $Y=0.51
c69 20 0 2.12886e-20 $X=2.11 $Y=0.84
r70 41 46 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.575 $Y=2.88
+ $X2=0.575 $Y2=2.97
r71 40 42 5.06676 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.477 $Y=2.88
+ $X2=0.477 $Y2=2.715
r72 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=2.88 $X2=0.575 $Y2=2.88
r73 38 42 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.42 $Y=2.335
+ $X2=0.42 $Y2=2.715
r74 36 38 3.77045 $w=4.73e-07 $l=1.05e-07 $layer=LI1_cond $X=0.347 $Y=2.23
+ $X2=0.347 $Y2=2.335
r75 36 37 7.85596 $w=4.73e-07 $l=1.05e-07 $layer=LI1_cond $X=0.347 $Y=2.23
+ $X2=0.347 $Y2=2.125
r76 30 33 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=0.195 $Y=0.51
+ $X2=0.31 $Y2=0.51
r77 26 30 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.195 $Y=0.615
+ $X2=0.195 $Y2=0.51
r78 26 37 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=0.195 $Y=0.615
+ $X2=0.195 $Y2=2.125
r79 22 24 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.925 $Y=1.77
+ $X2=2.11 $Y2=1.77
r80 18 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.9 $Y=0.84 $X2=2.11
+ $Y2=0.84
r81 17 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.11 $Y=1.695
+ $X2=2.11 $Y2=1.77
r82 16 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.11 $Y=0.915
+ $X2=2.11 $Y2=0.84
r83 16 17 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.11 $Y=0.915
+ $X2=2.11 $Y2=1.695
r84 13 15 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.925 $Y=2.895
+ $X2=1.925 $Y2=2.165
r85 12 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=1.845
+ $X2=1.925 $Y2=1.77
r86 12 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=1.845
+ $X2=1.925 $Y2=2.165
r87 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.9 $Y=0.765 $X2=1.9
+ $Y2=0.84
r88 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.9 $Y=0.765 $X2=1.9
+ $Y2=0.445
r89 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=2.97
+ $X2=0.575 $Y2=2.97
r90 7 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.85 $Y=2.97
+ $X2=1.925 $Y2=2.895
r91 7 8 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.85 $Y=2.97 $X2=0.74
+ $Y2=2.97
r92 2 36 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.295
+ $Y=1.955 $X2=0.42 $Y2=2.23
r93 1 33 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_M%VPWR 1 2 9 12 13 15 19 22 23 24 25 26 27 35
+ 36 39
r37 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 36 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 33 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.71 $Y2=3.33
r41 33 35 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 27 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 27 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 24 30 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.87 $Y=3.33 $X2=0.72
+ $Y2=3.33
r46 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.33
+ $X2=0.955 $Y2=3.33
r47 22 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=3.33
r48 21 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.545
+ $X2=1.71 $Y2=2.46
r49 21 22 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.71 $Y=2.545 $X2=1.71
+ $Y2=3.245
r50 17 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.375
+ $X2=1.71 $Y2=2.46
r51 17 19 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.71 $Y=2.375
+ $X2=1.71 $Y2=2.23
r52 16 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.955 $Y2=3.33
r53 15 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=1.71 $Y2=3.33
r54 15 16 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=1.04 $Y2=3.33
r55 14 23 1.34256 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.04 $Y=2.46
+ $X2=0.902 $Y2=2.46
r56 13 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.46
+ $X2=1.71 $Y2=2.46
r57 13 14 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.625 $Y=2.46
+ $X2=1.04 $Y2=2.46
r58 12 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=3.245
+ $X2=0.955 $Y2=3.33
r59 11 23 5.16603 $w=1.7e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.955 $Y=2.545
+ $X2=0.902 $Y2=2.46
r60 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.955 $Y=2.545
+ $X2=0.955 $Y2=3.245
r61 7 23 5.16603 $w=1.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.85 $Y=2.375
+ $X2=0.902 $Y2=2.46
r62 7 9 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.85 $Y=2.375
+ $X2=0.85 $Y2=2.23
r63 2 19 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.955 $X2=1.71 $Y2=2.23
r64 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.955 $X2=0.85 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_M%Y 1 2 3 10 11 17 23 27
r29 25 27 0.570093 $w=4.28e-07 $l=2e-08 $layer=LI1_cond $X=2.14 $Y=1.885
+ $X2=2.16 $Y2=1.885
r30 23 25 13.1121 $w=4.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.68 $Y=1.885
+ $X2=2.14 $Y2=1.885
r31 21 23 11.4019 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=1.885 $X2=1.68
+ $Y2=1.885
r32 11 27 6.19161 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.885
r33 11 25 2.26247 $w=3.3e-07 $l=3.05e-07 $layer=LI1_cond $X=2.14 $Y=1.58
+ $X2=2.14 $Y2=1.885
r34 11 17 26.9798 $w=4.98e-07 $l=1.07e-06 $layer=LI1_cond $X=2.14 $Y=1.58
+ $X2=2.14 $Y2=0.51
r35 10 23 6.19161 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.885
r36 3 25 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.955 $X2=2.14 $Y2=2.1
r37 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.955 $X2=1.28 $Y2=2.1
r38 1 17 182 $w=1.7e-07 $l=3.47851e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.14 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_M%VGND 1 8 10 17 18 21
c34 18 0 2.12886e-20 $X=2.16 $Y=0
r35 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r37 14 17 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r38 12 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.74
+ $Y2=0
r39 12 14 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=1.2
+ $Y2=0
r40 10 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r41 10 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r42 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 6 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r44 6 8 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0.38
r45 1 8 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.38
.ends

