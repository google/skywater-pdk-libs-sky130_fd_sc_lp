* File: sky130_fd_sc_lp__dfstp_2.pxi.spice
* Created: Wed Sep  2 09:44:27 2020
* 
x_PM_SKY130_FD_SC_LP__DFSTP_2%CLK N_CLK_c_246_n N_CLK_c_251_n N_CLK_M1009_g
+ N_CLK_M1007_g N_CLK_c_252_n CLK CLK N_CLK_c_249_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%CLK
x_PM_SKY130_FD_SC_LP__DFSTP_2%D N_D_c_289_n N_D_c_290_n N_D_c_293_n N_D_c_294_n
+ N_D_c_291_n N_D_M1006_g N_D_c_295_n N_D_M1011_g D N_D_c_292_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%D
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_196_465# N_A_196_465#_M1015_d
+ N_A_196_465#_M1024_d N_A_196_465#_M1002_g N_A_196_465#_c_345_n
+ N_A_196_465#_c_346_n N_A_196_465#_M1031_g N_A_196_465#_M1030_g
+ N_A_196_465#_M1014_g N_A_196_465#_c_349_n N_A_196_465#_c_350_n
+ N_A_196_465#_c_367_n N_A_196_465#_c_368_n N_A_196_465#_c_351_n
+ N_A_196_465#_c_352_n N_A_196_465#_c_353_n N_A_196_465#_c_354_n
+ N_A_196_465#_c_369_n N_A_196_465#_c_355_n N_A_196_465#_c_356_n
+ N_A_196_465#_c_374_n N_A_196_465#_c_357_n N_A_196_465#_c_358_n
+ N_A_196_465#_c_359_n N_A_196_465#_c_360_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%A_196_465#
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_614_93# N_A_614_93#_M1020_s N_A_614_93#_M1003_d
+ N_A_614_93#_M1021_g N_A_614_93#_M1023_g N_A_614_93#_c_534_n
+ N_A_614_93#_c_535_n N_A_614_93#_c_526_n N_A_614_93#_c_536_n
+ N_A_614_93#_c_527_n N_A_614_93#_c_528_n N_A_614_93#_c_529_n
+ N_A_614_93#_c_553_p N_A_614_93#_c_530_n N_A_614_93#_c_531_n
+ N_A_614_93#_c_532_n PM_SKY130_FD_SC_LP__DFSTP_2%A_614_93#
x_PM_SKY130_FD_SC_LP__DFSTP_2%SET_B N_SET_B_M1025_g N_SET_B_M1010_g
+ N_SET_B_c_611_n N_SET_B_M1013_g N_SET_B_c_620_n N_SET_B_c_621_n
+ N_SET_B_M1033_g N_SET_B_c_612_n N_SET_B_c_613_n N_SET_B_c_614_n
+ N_SET_B_c_615_n N_SET_B_c_616_n N_SET_B_c_625_n N_SET_B_c_626_n SET_B SET_B
+ SET_B SET_B N_SET_B_c_629_n PM_SKY130_FD_SC_LP__DFSTP_2%SET_B
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_486_119# N_A_486_119#_M1029_d
+ N_A_486_119#_M1002_d N_A_486_119#_M1003_g N_A_486_119#_M1020_g
+ N_A_486_119#_c_734_n N_A_486_119#_M1000_g N_A_486_119#_c_736_n
+ N_A_486_119#_c_737_n N_A_486_119#_M1027_g N_A_486_119#_c_738_n
+ N_A_486_119#_c_739_n N_A_486_119#_c_740_n N_A_486_119#_c_741_n
+ N_A_486_119#_c_742_n N_A_486_119#_c_743_n N_A_486_119#_c_748_n
+ N_A_486_119#_c_744_n N_A_486_119#_c_775_n N_A_486_119#_c_750_n
+ N_A_486_119#_c_745_n PM_SKY130_FD_SC_LP__DFSTP_2%A_486_119#
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_27_465# N_A_27_465#_M1007_s N_A_27_465#_M1009_s
+ N_A_27_465#_M1024_g N_A_27_465#_M1015_g N_A_27_465#_c_891_n
+ N_A_27_465#_c_892_n N_A_27_465#_c_881_n N_A_27_465#_c_882_n
+ N_A_27_465#_M1029_g N_A_27_465#_M1019_g N_A_27_465#_c_894_n
+ N_A_27_465#_M1032_g N_A_27_465#_M1026_g N_A_27_465#_c_897_n
+ N_A_27_465#_c_898_n N_A_27_465#_c_885_n N_A_27_465#_c_899_n
+ N_A_27_465#_c_886_n N_A_27_465#_c_887_n N_A_27_465#_c_888_n
+ N_A_27_465#_c_889_n PM_SKY130_FD_SC_LP__DFSTP_2%A_27_465#
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_1309_65# N_A_1309_65#_M1017_d
+ N_A_1309_65#_M1004_d N_A_1309_65#_M1001_g N_A_1309_65#_c_1024_n
+ N_A_1309_65#_c_1030_n N_A_1309_65#_c_1031_n N_A_1309_65#_c_1032_n
+ N_A_1309_65#_M1008_g N_A_1309_65#_c_1034_n N_A_1309_65#_c_1025_n
+ N_A_1309_65#_c_1035_n N_A_1309_65#_c_1036_n N_A_1309_65#_c_1026_n
+ N_A_1309_65#_c_1027_n N_A_1309_65#_c_1038_n N_A_1309_65#_c_1028_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%A_1309_65#
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_1158_47# N_A_1158_47#_M1030_d
+ N_A_1158_47#_M1014_d N_A_1158_47#_M1033_d N_A_1158_47#_c_1117_n
+ N_A_1158_47#_M1017_g N_A_1158_47#_c_1118_n N_A_1158_47#_c_1119_n
+ N_A_1158_47#_M1004_g N_A_1158_47#_c_1120_n N_A_1158_47#_c_1121_n
+ N_A_1158_47#_c_1122_n N_A_1158_47#_c_1123_n N_A_1158_47#_c_1124_n
+ N_A_1158_47#_c_1137_n N_A_1158_47#_c_1138_n N_A_1158_47#_M1018_g
+ N_A_1158_47#_c_1139_n N_A_1158_47#_M1005_g N_A_1158_47#_c_1126_n
+ N_A_1158_47#_c_1127_n N_A_1158_47#_c_1128_n N_A_1158_47#_c_1129_n
+ N_A_1158_47#_c_1130_n N_A_1158_47#_c_1142_n N_A_1158_47#_c_1143_n
+ N_A_1158_47#_c_1131_n N_A_1158_47#_c_1132_n N_A_1158_47#_c_1146_n
+ N_A_1158_47#_c_1147_n N_A_1158_47#_c_1148_n N_A_1158_47#_c_1133_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%A_1158_47#
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_1855_47# N_A_1855_47#_M1018_s
+ N_A_1855_47#_M1005_s N_A_1855_47#_M1016_g N_A_1855_47#_M1012_g
+ N_A_1855_47#_c_1260_n N_A_1855_47#_c_1261_n N_A_1855_47#_M1028_g
+ N_A_1855_47#_M1022_g N_A_1855_47#_c_1263_n N_A_1855_47#_c_1264_n
+ N_A_1855_47#_c_1265_n N_A_1855_47#_c_1266_n N_A_1855_47#_c_1267_n
+ N_A_1855_47#_c_1268_n N_A_1855_47#_c_1269_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%A_1855_47#
x_PM_SKY130_FD_SC_LP__DFSTP_2%VPWR N_VPWR_M1009_d N_VPWR_M1011_s N_VPWR_M1023_d
+ N_VPWR_M1025_d N_VPWR_M1008_d N_VPWR_M1004_s N_VPWR_M1005_d N_VPWR_M1022_s
+ N_VPWR_c_1328_n N_VPWR_c_1329_n N_VPWR_c_1330_n N_VPWR_c_1331_n
+ N_VPWR_c_1332_n N_VPWR_c_1333_n N_VPWR_c_1334_n N_VPWR_c_1335_n
+ N_VPWR_c_1336_n N_VPWR_c_1337_n N_VPWR_c_1338_n N_VPWR_c_1339_n
+ N_VPWR_c_1340_n N_VPWR_c_1341_n N_VPWR_c_1342_n N_VPWR_c_1343_n
+ N_VPWR_c_1344_n VPWR N_VPWR_c_1345_n N_VPWR_c_1346_n N_VPWR_c_1347_n
+ N_VPWR_c_1348_n N_VPWR_c_1349_n N_VPWR_c_1350_n N_VPWR_c_1351_n
+ N_VPWR_c_1352_n N_VPWR_c_1327_n PM_SKY130_FD_SC_LP__DFSTP_2%VPWR
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_400_119# N_A_400_119#_M1006_d
+ N_A_400_119#_M1011_d N_A_400_119#_c_1502_n N_A_400_119#_c_1468_n
+ N_A_400_119#_c_1466_n N_A_400_119#_c_1467_n N_A_400_119#_c_1470_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%A_400_119#
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_988_379# N_A_988_379#_M1000_d
+ N_A_988_379#_M1026_d N_A_988_379#_c_1511_n N_A_988_379#_c_1512_n
+ N_A_988_379#_c_1513_n PM_SKY130_FD_SC_LP__DFSTP_2%A_988_379#
x_PM_SKY130_FD_SC_LP__DFSTP_2%A_1095_425# N_A_1095_425#_M1014_s
+ N_A_1095_425#_M1008_s N_A_1095_425#_c_1538_n N_A_1095_425#_c_1539_n
+ N_A_1095_425#_c_1540_n N_A_1095_425#_c_1541_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%A_1095_425#
x_PM_SKY130_FD_SC_LP__DFSTP_2%Q N_Q_M1016_d N_Q_M1012_d Q Q Q Q Q Q Q
+ N_Q_c_1563_n PM_SKY130_FD_SC_LP__DFSTP_2%Q
x_PM_SKY130_FD_SC_LP__DFSTP_2%VGND N_VGND_M1007_d N_VGND_M1006_s N_VGND_M1021_d
+ N_VGND_M1010_d N_VGND_M1013_d N_VGND_M1018_d N_VGND_M1028_s N_VGND_c_1579_n
+ N_VGND_c_1580_n N_VGND_c_1581_n N_VGND_c_1582_n N_VGND_c_1583_n
+ N_VGND_c_1584_n N_VGND_c_1585_n N_VGND_c_1586_n N_VGND_c_1587_n
+ N_VGND_c_1588_n N_VGND_c_1589_n N_VGND_c_1590_n N_VGND_c_1591_n
+ N_VGND_c_1681_n VGND N_VGND_c_1592_n N_VGND_c_1593_n N_VGND_c_1594_n
+ N_VGND_c_1595_n N_VGND_c_1596_n N_VGND_c_1597_n N_VGND_c_1598_n
+ N_VGND_c_1599_n N_VGND_c_1600_n N_VGND_c_1601_n
+ PM_SKY130_FD_SC_LP__DFSTP_2%VGND
cc_1 VNB N_CLK_c_246_n 0.0241377f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=2.065
cc_2 VNB N_CLK_M1007_g 0.0223853f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.58
cc_3 VNB CLK 0.00944533f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_CLK_c_249_n 0.0456256f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.09
cc_5 VNB N_D_c_289_n 0.0227927f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.255
cc_6 VNB N_D_c_290_n 0.0214855f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=2.065
cc_7 VNB N_D_c_291_n 0.0167212f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.645
cc_8 VNB N_D_c_292_n 0.0246504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_196_465#_c_345_n 0.0109044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_196_465#_c_346_n 0.0116158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_196_465#_M1031_g 0.0332932f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_A_196_465#_M1030_g 0.0388755f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.09
cc_13 VNB N_A_196_465#_c_349_n 0.0169862f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.09
cc_14 VNB N_A_196_465#_c_350_n 0.00482332f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.295
cc_15 VNB N_A_196_465#_c_351_n 0.00473498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_196_465#_c_352_n 0.00356451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_196_465#_c_353_n 0.00238975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_196_465#_c_354_n 0.00430364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_196_465#_c_355_n 0.00182226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_196_465#_c_356_n 0.0441677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_196_465#_c_357_n 0.00144207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_196_465#_c_358_n 0.0100823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_196_465#_c_359_n 0.00469572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_196_465#_c_360_n 0.0357034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_614_93#_c_526_n 0.0170454f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.09
cc_26 VNB N_A_614_93#_c_527_n 0.0102505f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.295
cc_27 VNB N_A_614_93#_c_528_n 3.11212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_614_93#_c_529_n 0.0331874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_614_93#_c_530_n 0.00510864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_614_93#_c_531_n 0.0189682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_614_93#_c_532_n 0.00991981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_SET_B_M1010_g 0.0270317f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.58
cc_33 VNB N_SET_B_c_611_n 0.0689014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_SET_B_c_612_n 0.0185226f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.09
cc_35 VNB N_SET_B_c_613_n 0.00587103f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.925
cc_36 VNB N_SET_B_c_614_n 0.00446596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_SET_B_c_615_n 0.011017f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.295
cc_38 VNB N_SET_B_c_616_n 0.0330707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB SET_B 0.00553878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB SET_B 0.0127543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_486_119#_M1003_g 0.00241197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_486_119#_M1020_g 0.0485266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_486_119#_c_734_n 0.0250304f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_44 VNB N_A_486_119#_M1000_g 0.00270324f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.09
cc_45 VNB N_A_486_119#_c_736_n 0.0222871f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.09
cc_46 VNB N_A_486_119#_c_737_n 0.0181083f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.925
cc_47 VNB N_A_486_119#_c_738_n 0.016213f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.295
cc_48 VNB N_A_486_119#_c_739_n 0.0326349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_486_119#_c_740_n 0.0119037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_486_119#_c_741_n 0.0203167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_486_119#_c_742_n 0.0265093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_486_119#_c_743_n 0.00333276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_486_119#_c_744_n 0.00538172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_486_119#_c_745_n 3.86187e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_465#_M1015_g 0.0461578f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_56 VNB N_A_27_465#_c_881_n 0.102619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_465#_c_882_n 0.0113962f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.255
cc_58 VNB N_A_27_465#_M1029_g 0.0338535f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.09
cc_59 VNB N_A_27_465#_M1032_g 0.047494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_465#_c_885_n 0.0318268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_465#_c_886_n 0.00128424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_27_465#_c_887_n 0.0135009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_465#_c_888_n 0.00402994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_27_465#_c_889_n 0.0228015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1309_65#_M1001_g 0.0374712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1309_65#_c_1024_n 0.00128857f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=2.14
cc_67 VNB N_A_1309_65#_c_1025_n 0.0210821f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.09
cc_68 VNB N_A_1309_65#_c_1026_n 0.0182097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1309_65#_c_1027_n 0.015128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1309_65#_c_1028_n 0.00401544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1158_47#_c_1117_n 0.0189711f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=2.14
cc_72 VNB N_A_1158_47#_c_1118_n 0.0647042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1158_47#_c_1119_n 0.0117256f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_74 VNB N_A_1158_47#_c_1120_n 0.0117856f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.09
cc_75 VNB N_A_1158_47#_c_1121_n 0.021098f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.09
cc_76 VNB N_A_1158_47#_c_1122_n 0.00476428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1158_47#_c_1123_n 0.0325494f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.09
cc_78 VNB N_A_1158_47#_c_1124_n 0.0121868f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.295
cc_79 VNB N_A_1158_47#_M1018_g 0.0216454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1158_47#_c_1126_n 0.011701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1158_47#_c_1127_n 0.00642107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1158_47#_c_1128_n 0.00446755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1158_47#_c_1129_n 0.0204053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1158_47#_c_1130_n 0.00444991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1158_47#_c_1131_n 0.0171068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1158_47#_c_1132_n 0.00267605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1158_47#_c_1133_n 0.0842395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1855_47#_M1012_g 0.00864382f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.14
cc_89 VNB N_A_1855_47#_c_1260_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_90 VNB N_A_1855_47#_c_1261_n 0.0215271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1855_47#_M1022_g 0.0255673f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.09
cc_92 VNB N_A_1855_47#_c_1263_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=0.925
cc_93 VNB N_A_1855_47#_c_1264_n 0.0123107f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.295
cc_94 VNB N_A_1855_47#_c_1265_n 0.00307852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1855_47#_c_1266_n 0.00897222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1855_47#_c_1267_n 0.00536819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1855_47#_c_1268_n 0.0397206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1855_47#_c_1269_n 0.0176094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VPWR_c_1327_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_400_119#_c_1466_n 0.00624608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_400_119#_c_1467_n 0.00458034f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.09
cc_102 VNB N_Q_c_1563_n 0.00854714f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.09
cc_103 VNB N_VGND_c_1579_n 0.00215472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1580_n 0.0127903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1581_n 0.0223226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1582_n 0.00790143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1583_n 0.0113054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1584_n 4.07942e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1585_n 0.00296085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1586_n 0.0113208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1587_n 0.0499388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1588_n 0.03913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1589_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1590_n 0.0541549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1591_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1592_n 0.0180939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1593_n 0.0162973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1594_n 0.040712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1595_n 0.0609401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1596_n 0.0150561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1597_n 0.00511859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1598_n 0.00392849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1599_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1600_n 0.00491384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1601_n 0.579035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VPB N_CLK_c_246_n 0.023017f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=2.065
cc_127 VPB N_CLK_c_251_n 0.0214245f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_128 VPB N_CLK_c_252_n 0.0274802f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.14
cc_129 VPB N_D_c_293_n 0.0207919f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_130 VPB N_D_c_294_n 0.0236031f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.645
cc_131 VPB N_D_c_295_n 0.0177986f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.58
cc_132 VPB D 0.00337299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_D_c_292_n 0.0278198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_196_465#_M1002_g 0.0368518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_196_465#_c_345_n 0.0104077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_196_465#_c_346_n 0.00358714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_196_465#_M1014_g 0.0436231f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.925
cc_138 VPB N_A_196_465#_c_349_n 0.0209334f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.09
cc_139 VPB N_A_196_465#_c_350_n 0.00713954f $X=-0.19 $Y=1.655 $X2=0.642
+ $Y2=1.295
cc_140 VPB N_A_196_465#_c_367_n 8.58732e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_196_465#_c_368_n 0.00174455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_196_465#_c_369_n 0.0118493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_196_465#_c_355_n 0.00314045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_196_465#_c_360_n 0.00995148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_614_93#_M1023_g 0.0179283f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_146 VPB N_A_614_93#_c_534_n 0.0120162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_614_93#_c_535_n 0.0314616f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.09
cc_148 VPB N_A_614_93#_c_536_n 0.00159259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_614_93#_c_532_n 0.0105327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_SET_B_M1025_g 0.0198438f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_151 VPB N_SET_B_c_620_n 0.0404207f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.14
cc_152 VPB N_SET_B_c_621_n 0.0148087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_SET_B_M1033_g 0.0404857f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_SET_B_c_612_n 0.0080427f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.09
cc_155 VPB N_SET_B_c_613_n 0.00230423f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.925
cc_156 VPB N_SET_B_c_625_n 0.0080889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_SET_B_c_626_n 0.0315859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB SET_B 0.00321223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB SET_B 0.00711893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_SET_B_c_629_n 0.0242891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_486_119#_M1003_g 0.0421051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_486_119#_M1000_g 0.0300986f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.09
cc_163 VPB N_A_486_119#_c_748_n 0.00866941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_486_119#_c_744_n 0.0108085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_486_119#_c_750_n 3.83052e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_486_119#_c_745_n 0.00340515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_27_465#_M1024_g 0.0367512f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=2.14
cc_168 VPB N_A_27_465#_c_891_n 0.129924f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_169 VPB N_A_27_465#_c_892_n 0.0122479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_27_465#_M1019_g 0.0344581f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.09
cc_171 VPB N_A_27_465#_c_894_n 0.258192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_27_465#_M1032_g 0.0100737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_27_465#_M1026_g 0.0134488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_27_465#_c_897_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_27_465#_c_898_n 0.014887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_27_465#_c_899_n 0.049176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_27_465#_c_886_n 0.0015813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_27_465#_c_888_n 0.00692367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_27_465#_c_889_n 0.0274459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1309_65#_c_1024_n 0.0300032f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.14
cc_181 VPB N_A_1309_65#_c_1030_n 0.0443363f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_182 VPB N_A_1309_65#_c_1031_n 0.0210104f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_183 VPB N_A_1309_65#_c_1032_n 0.0104278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1309_65#_M1008_g 0.0272589f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.09
cc_185 VPB N_A_1309_65#_c_1034_n 0.112616f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.09
cc_186 VPB N_A_1309_65#_c_1035_n 0.0156203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1309_65#_c_1036_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1309_65#_c_1027_n 0.010684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1309_65#_c_1038_n 0.0661619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1158_47#_M1004_g 0.0266334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1158_47#_c_1120_n 0.00529972f $X=-0.19 $Y=1.655 $X2=0.505
+ $Y2=1.09
cc_192 VPB N_A_1158_47#_c_1122_n 0.00820206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_1158_47#_c_1137_n 0.0330002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_1158_47#_c_1138_n 0.0135842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1158_47#_c_1139_n 0.0195532f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1158_47#_c_1126_n 0.0108831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_1158_47#_c_1127_n 2.22871e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1158_47#_c_1142_n 0.0180063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_1158_47#_c_1143_n 0.00103876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1158_47#_c_1131_n 0.00859512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1158_47#_c_1132_n 0.0114297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1158_47#_c_1146_n 0.0031333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1158_47#_c_1147_n 2.99451e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1158_47#_c_1148_n 0.00263254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1855_47#_M1012_g 0.0237211f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.14
cc_206 VPB N_A_1855_47#_M1022_g 0.0272176f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.09
cc_207 VPB N_A_1855_47#_c_1265_n 0.0129687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1328_n 0.0108006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1329_n 0.0169133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1330_n 0.012206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1331_n 0.00269989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1332_n 0.0143757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1333_n 0.00883621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1334_n 0.0151993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1335_n 0.022426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1336_n 0.0130585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1337_n 0.0112949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1338_n 0.0666542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1339_n 0.0186345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1340_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1341_n 0.0371424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1342_n 0.00356967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1343_n 0.0675247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1344_n 0.00303699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1345_n 0.0211152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1346_n 0.0185345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1347_n 0.0314979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1348_n 0.0199215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1349_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1350_n 0.00769791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1351_n 0.00263749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1352_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1327_n 0.0686901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_400_119#_c_1468_n 0.00133479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_400_119#_c_1466_n 0.00337844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_400_119#_c_1470_n 0.00757078f $X=-0.19 $Y=1.655 $X2=0.642
+ $Y2=0.925
cc_237 VPB N_A_988_379#_c_1511_n 0.0128879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_988_379#_c_1512_n 0.00433569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_988_379#_c_1513_n 0.0260717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1095_425#_c_1538_n 0.00337954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_1095_425#_c_1539_n 0.00366833f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=2.14
cc_242 VPB N_A_1095_425#_c_1540_n 0.00167045f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=0.84
cc_243 VPB N_A_1095_425#_c_1541_n 0.00386885f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.21
cc_244 VPB N_Q_c_1563_n 0.00487158f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.09
cc_245 CLK N_A_196_465#_c_353_n 0.0439115f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_246 N_CLK_c_249_n N_A_196_465#_c_353_n 2.493e-19 $X=0.505 $Y=1.09 $X2=0 $Y2=0
cc_247 CLK N_A_196_465#_c_374_n 0.00165478f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_248 N_CLK_c_246_n N_A_27_465#_M1024_g 0.00259742f $X=0.23 $Y=2.065 $X2=0
+ $Y2=0
cc_249 N_CLK_c_252_n N_A_27_465#_M1024_g 0.00798027f $X=0.475 $Y=2.14 $X2=0
+ $Y2=0
cc_250 N_CLK_c_246_n N_A_27_465#_M1015_g 0.00249896f $X=0.23 $Y=2.065 $X2=0
+ $Y2=0
cc_251 CLK N_A_27_465#_M1015_g 0.00569036f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_252 N_CLK_c_249_n N_A_27_465#_M1015_g 0.0192996f $X=0.505 $Y=1.09 $X2=0 $Y2=0
cc_253 N_CLK_c_251_n N_A_27_465#_c_892_n 0.00798027f $X=0.475 $Y=2.215 $X2=0
+ $Y2=0
cc_254 N_CLK_M1007_g N_A_27_465#_c_882_n 0.0113757f $X=0.505 $Y=0.58 $X2=0 $Y2=0
cc_255 N_CLK_c_246_n N_A_27_465#_c_885_n 0.0121407f $X=0.23 $Y=2.065 $X2=0 $Y2=0
cc_256 N_CLK_M1007_g N_A_27_465#_c_885_n 0.00463299f $X=0.505 $Y=0.58 $X2=0
+ $Y2=0
cc_257 CLK N_A_27_465#_c_885_n 0.0407542f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_258 N_CLK_c_249_n N_A_27_465#_c_885_n 0.0123365f $X=0.505 $Y=1.09 $X2=0 $Y2=0
cc_259 N_CLK_c_246_n N_A_27_465#_c_899_n 0.00842207f $X=0.23 $Y=2.065 $X2=0
+ $Y2=0
cc_260 N_CLK_c_251_n N_A_27_465#_c_899_n 0.00341644f $X=0.475 $Y=2.215 $X2=0
+ $Y2=0
cc_261 N_CLK_c_252_n N_A_27_465#_c_899_n 0.0145886f $X=0.475 $Y=2.14 $X2=0 $Y2=0
cc_262 N_CLK_c_252_n N_A_27_465#_c_886_n 0.00601154f $X=0.475 $Y=2.14 $X2=0
+ $Y2=0
cc_263 CLK N_A_27_465#_c_886_n 0.0340232f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_264 N_CLK_c_249_n N_A_27_465#_c_886_n 0.00272476f $X=0.505 $Y=1.09 $X2=0
+ $Y2=0
cc_265 N_CLK_c_249_n N_A_27_465#_c_887_n 0.00477279f $X=0.505 $Y=1.09 $X2=0
+ $Y2=0
cc_266 N_CLK_c_246_n N_A_27_465#_c_888_n 0.0118065f $X=0.23 $Y=2.065 $X2=0 $Y2=0
cc_267 N_CLK_c_249_n N_A_27_465#_c_888_n 0.00211599f $X=0.505 $Y=1.09 $X2=0
+ $Y2=0
cc_268 N_CLK_c_246_n N_A_27_465#_c_889_n 0.0215144f $X=0.23 $Y=2.065 $X2=0 $Y2=0
cc_269 N_CLK_c_252_n N_A_27_465#_c_889_n 0.00217096f $X=0.475 $Y=2.14 $X2=0
+ $Y2=0
cc_270 CLK N_A_27_465#_c_889_n 0.00583462f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_271 N_CLK_c_249_n N_A_27_465#_c_889_n 0.00913195f $X=0.505 $Y=1.09 $X2=0
+ $Y2=0
cc_272 N_CLK_c_251_n N_VPWR_c_1328_n 0.0031763f $X=0.475 $Y=2.215 $X2=0 $Y2=0
cc_273 N_CLK_c_251_n N_VPWR_c_1339_n 0.00465548f $X=0.475 $Y=2.215 $X2=0 $Y2=0
cc_274 N_CLK_c_251_n N_VPWR_c_1327_n 0.00922874f $X=0.475 $Y=2.215 $X2=0 $Y2=0
cc_275 N_CLK_M1007_g N_VGND_c_1579_n 0.0111078f $X=0.505 $Y=0.58 $X2=0 $Y2=0
cc_276 CLK N_VGND_c_1579_n 0.0214959f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_277 N_CLK_c_249_n N_VGND_c_1579_n 5.53818e-19 $X=0.505 $Y=1.09 $X2=0 $Y2=0
cc_278 N_CLK_M1007_g N_VGND_c_1592_n 0.00444681f $X=0.505 $Y=0.58 $X2=0 $Y2=0
cc_279 N_CLK_M1007_g N_VGND_c_1601_n 0.00789248f $X=0.505 $Y=0.58 $X2=0 $Y2=0
cc_280 CLK N_VGND_c_1601_n 0.00195932f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_281 N_D_c_293_n N_A_196_465#_M1002_g 0.0179675f $X=1.85 $Y=2.13 $X2=0 $Y2=0
cc_282 D N_A_196_465#_M1002_g 0.00251079f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_283 N_D_c_292_n N_A_196_465#_M1002_g 0.00154541f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_284 N_D_c_289_n N_A_196_465#_M1031_g 0.00142137f $X=1.85 $Y=1.2 $X2=0 $Y2=0
cc_285 N_D_c_289_n N_A_196_465#_c_349_n 0.00793962f $X=1.85 $Y=1.2 $X2=0 $Y2=0
cc_286 N_D_c_293_n N_A_196_465#_c_349_n 0.00958063f $X=1.85 $Y=2.13 $X2=0 $Y2=0
cc_287 D N_A_196_465#_c_349_n 2.82918e-19 $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_288 N_D_c_292_n N_A_196_465#_c_349_n 0.0222378f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_289 N_D_c_295_n N_A_196_465#_c_367_n 0.00186412f $X=1.925 $Y=2.205 $X2=0
+ $Y2=0
cc_290 N_D_c_291_n N_A_196_465#_c_351_n 0.00296912f $X=1.925 $Y=1.125 $X2=0
+ $Y2=0
cc_291 N_D_c_289_n N_A_196_465#_c_352_n 0.00586102f $X=1.85 $Y=1.2 $X2=0 $Y2=0
cc_292 N_D_c_293_n N_A_196_465#_c_352_n 0.00333834f $X=1.85 $Y=2.13 $X2=0 $Y2=0
cc_293 D N_A_196_465#_c_352_n 0.0293043f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_294 N_D_c_292_n N_A_196_465#_c_352_n 0.0161606f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_295 N_D_c_292_n N_A_196_465#_c_354_n 0.004033f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_296 N_D_c_295_n N_A_196_465#_c_369_n 0.00226217f $X=1.925 $Y=2.205 $X2=0
+ $Y2=0
cc_297 D N_A_196_465#_c_369_n 0.0293717f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_298 N_D_c_292_n N_A_196_465#_c_369_n 0.00728054f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_299 N_D_c_289_n N_A_196_465#_c_355_n 0.00127169f $X=1.85 $Y=1.2 $X2=0 $Y2=0
cc_300 N_D_c_293_n N_A_196_465#_c_355_n 4.15302e-19 $X=1.85 $Y=2.13 $X2=0 $Y2=0
cc_301 D N_A_196_465#_c_355_n 0.00302485f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_302 N_D_c_292_n N_A_196_465#_c_355_n 0.00132419f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_303 N_D_c_289_n N_A_196_465#_c_356_n 0.0115246f $X=1.85 $Y=1.2 $X2=0 $Y2=0
cc_304 N_D_c_290_n N_A_196_465#_c_356_n 0.00823671f $X=1.655 $Y=1.2 $X2=0 $Y2=0
cc_305 N_D_c_292_n N_A_196_465#_c_356_n 0.00330439f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_306 N_D_c_290_n N_A_196_465#_c_357_n 0.00769135f $X=1.655 $Y=1.2 $X2=0 $Y2=0
cc_307 N_D_c_292_n N_A_196_465#_c_357_n 0.00854552f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_308 N_D_c_292_n N_A_27_465#_M1024_g 0.0108953f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_309 N_D_c_290_n N_A_27_465#_M1015_g 0.0159907f $X=1.655 $Y=1.2 $X2=0 $Y2=0
cc_310 N_D_c_295_n N_A_27_465#_c_891_n 0.0103107f $X=1.925 $Y=2.205 $X2=0 $Y2=0
cc_311 N_D_c_291_n N_A_27_465#_c_881_n 0.0104164f $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_312 N_D_c_291_n N_A_27_465#_M1029_g 0.0125031f $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_313 N_D_c_292_n N_A_27_465#_c_889_n 0.0159907f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_314 N_D_c_294_n N_VPWR_c_1329_n 0.00715989f $X=1.655 $Y=2.13 $X2=0 $Y2=0
cc_315 N_D_c_295_n N_VPWR_c_1329_n 0.0105172f $X=1.925 $Y=2.205 $X2=0 $Y2=0
cc_316 D N_VPWR_c_1329_n 0.0191467f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_317 N_D_c_295_n N_VPWR_c_1327_n 7.88961e-19 $X=1.925 $Y=2.205 $X2=0 $Y2=0
cc_318 N_D_c_295_n N_A_400_119#_c_1468_n 0.00127846f $X=1.925 $Y=2.205 $X2=0
+ $Y2=0
cc_319 N_D_c_289_n N_A_400_119#_c_1466_n 0.00196889f $X=1.85 $Y=1.2 $X2=0 $Y2=0
cc_320 D N_A_400_119#_c_1466_n 0.00818219f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_321 N_D_c_292_n N_A_400_119#_c_1466_n 0.00221535f $X=1.49 $Y=1.97 $X2=0 $Y2=0
cc_322 N_D_c_291_n N_A_400_119#_c_1467_n 0.00295457f $X=1.925 $Y=1.125 $X2=0
+ $Y2=0
cc_323 N_D_c_293_n N_A_400_119#_c_1470_n 0.0032408f $X=1.85 $Y=2.13 $X2=0 $Y2=0
cc_324 D N_A_400_119#_c_1470_n 0.00543178f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_325 N_D_c_290_n N_VGND_c_1580_n 0.00778068f $X=1.655 $Y=1.2 $X2=0 $Y2=0
cc_326 N_D_c_291_n N_VGND_c_1580_n 0.00594441f $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_327 N_D_c_291_n N_VGND_c_1601_n 9.39239e-19 $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_328 N_A_196_465#_c_356_n N_A_614_93#_c_534_n 0.00108751f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_329 N_A_196_465#_M1002_g N_A_614_93#_c_535_n 0.00303994f $X=2.355 $Y=2.525
+ $X2=0 $Y2=0
cc_330 N_A_196_465#_c_356_n N_A_614_93#_c_526_n 0.0175568f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_331 N_A_196_465#_M1031_g N_A_614_93#_c_528_n 0.00120255f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_332 N_A_196_465#_c_356_n N_A_614_93#_c_528_n 0.022835f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_333 N_A_196_465#_c_346_n N_A_614_93#_c_529_n 0.0339593f $X=2.785 $Y=1.435
+ $X2=0 $Y2=0
cc_334 N_A_196_465#_c_356_n N_A_614_93#_c_529_n 0.00207561f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_335 N_A_196_465#_c_356_n N_A_614_93#_c_530_n 0.00467942f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_336 N_A_196_465#_M1031_g N_A_614_93#_c_531_n 0.0339593f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_337 N_A_196_465#_c_346_n N_A_614_93#_c_532_n 0.00418355f $X=2.785 $Y=1.435
+ $X2=0 $Y2=0
cc_338 N_A_196_465#_c_350_n N_A_614_93#_c_532_n 0.00303994f $X=2.355 $Y=1.68
+ $X2=0 $Y2=0
cc_339 N_A_196_465#_c_356_n N_SET_B_c_613_n 0.0147904f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_340 N_A_196_465#_c_356_n N_SET_B_c_614_n 0.0082435f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_341 N_A_196_465#_c_356_n N_SET_B_c_615_n 0.0315835f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_342 N_A_196_465#_c_358_n N_SET_B_c_615_n 0.00133684f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_343 N_A_196_465#_c_359_n N_SET_B_c_615_n 4.94263e-19 $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_344 N_A_196_465#_c_356_n N_SET_B_c_616_n 3.42511e-19 $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_345 N_A_196_465#_c_356_n N_SET_B_c_625_n 0.00426613f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_346 N_A_196_465#_c_356_n N_SET_B_c_626_n 6.93625e-19 $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_347 N_A_196_465#_M1030_g SET_B 0.00256559f $X=5.715 $Y=0.555 $X2=0 $Y2=0
cc_348 N_A_196_465#_c_358_n SET_B 0.00113403f $X=5.52 $Y=1.295 $X2=0 $Y2=0
cc_349 N_A_196_465#_c_359_n SET_B 0.0281662f $X=5.52 $Y=1.295 $X2=0 $Y2=0
cc_350 N_A_196_465#_c_360_n SET_B 0.00653544f $X=5.715 $Y=1.51 $X2=0 $Y2=0
cc_351 N_A_196_465#_M1014_g N_SET_B_c_629_n 0.0185793f $X=5.815 $Y=2.335 $X2=0
+ $Y2=0
cc_352 N_A_196_465#_c_356_n N_SET_B_c_629_n 0.0310327f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_353 N_A_196_465#_c_358_n N_SET_B_c_629_n 0.00248956f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_354 N_A_196_465#_c_359_n N_SET_B_c_629_n 0.0239669f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_355 N_A_196_465#_c_360_n N_SET_B_c_629_n 0.00879639f $X=5.715 $Y=1.51 $X2=0
+ $Y2=0
cc_356 N_A_196_465#_c_356_n N_A_486_119#_M1020_g 9.50914e-19 $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_357 N_A_196_465#_c_356_n N_A_486_119#_c_734_n 0.0105044f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_358 N_A_196_465#_c_360_n N_A_486_119#_M1000_g 0.00209279f $X=5.715 $Y=1.51
+ $X2=0 $Y2=0
cc_359 N_A_196_465#_M1030_g N_A_486_119#_c_736_n 0.00558481f $X=5.715 $Y=0.555
+ $X2=0 $Y2=0
cc_360 N_A_196_465#_c_356_n N_A_486_119#_c_736_n 0.00742566f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_361 N_A_196_465#_c_358_n N_A_486_119#_c_736_n 0.00138257f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_362 N_A_196_465#_c_359_n N_A_486_119#_c_736_n 0.00424282f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_363 N_A_196_465#_c_360_n N_A_486_119#_c_736_n 0.0179862f $X=5.715 $Y=1.51
+ $X2=0 $Y2=0
cc_364 N_A_196_465#_M1030_g N_A_486_119#_c_737_n 0.0634169f $X=5.715 $Y=0.555
+ $X2=0 $Y2=0
cc_365 N_A_196_465#_c_356_n N_A_486_119#_c_738_n 0.00179429f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_366 N_A_196_465#_c_356_n N_A_486_119#_c_739_n 0.00640737f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_367 N_A_196_465#_c_356_n N_A_486_119#_c_742_n 0.00487384f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_368 N_A_196_465#_c_358_n N_A_486_119#_c_742_n 0.0013652f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_369 N_A_196_465#_c_359_n N_A_486_119#_c_742_n 5.42335e-19 $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_370 N_A_196_465#_c_360_n N_A_486_119#_c_742_n 0.00164743f $X=5.715 $Y=1.51
+ $X2=0 $Y2=0
cc_371 N_A_196_465#_c_345_n N_A_486_119#_c_743_n 0.00117947f $X=2.67 $Y=1.59
+ $X2=0 $Y2=0
cc_372 N_A_196_465#_c_346_n N_A_486_119#_c_743_n 0.00520506f $X=2.785 $Y=1.435
+ $X2=0 $Y2=0
cc_373 N_A_196_465#_M1031_g N_A_486_119#_c_743_n 0.0166293f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_374 N_A_196_465#_c_356_n N_A_486_119#_c_743_n 0.0157931f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_375 N_A_196_465#_M1002_g N_A_486_119#_c_748_n 0.00520166f $X=2.355 $Y=2.525
+ $X2=0 $Y2=0
cc_376 N_A_196_465#_c_350_n N_A_486_119#_c_748_n 0.00138292f $X=2.355 $Y=1.68
+ $X2=0 $Y2=0
cc_377 N_A_196_465#_c_346_n N_A_486_119#_c_744_n 0.00248916f $X=2.785 $Y=1.435
+ $X2=0 $Y2=0
cc_378 N_A_196_465#_c_356_n N_A_486_119#_c_744_n 0.0192808f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_379 N_A_196_465#_c_345_n N_A_486_119#_c_775_n 0.00359004f $X=2.67 $Y=1.59
+ $X2=0 $Y2=0
cc_380 N_A_196_465#_M1031_g N_A_486_119#_c_775_n 0.00641939f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_381 N_A_196_465#_c_356_n N_A_486_119#_c_775_n 0.00729496f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_382 N_A_196_465#_c_345_n N_A_486_119#_c_750_n 0.00246931f $X=2.67 $Y=1.59
+ $X2=0 $Y2=0
cc_383 N_A_196_465#_c_346_n N_A_486_119#_c_750_n 0.00441098f $X=2.785 $Y=1.435
+ $X2=0 $Y2=0
cc_384 N_A_196_465#_c_350_n N_A_486_119#_c_750_n 2.72469e-19 $X=2.355 $Y=1.68
+ $X2=0 $Y2=0
cc_385 N_A_196_465#_c_356_n N_A_486_119#_c_745_n 0.0125814f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_386 N_A_196_465#_c_369_n N_A_27_465#_M1024_g 0.00912067f $X=1.13 $Y=2.315
+ $X2=0 $Y2=0
cc_387 N_A_196_465#_c_351_n N_A_27_465#_M1015_g 0.00238098f $X=1.19 $Y=0.58
+ $X2=0 $Y2=0
cc_388 N_A_196_465#_c_353_n N_A_27_465#_M1015_g 0.00568267f $X=1.19 $Y=1.005
+ $X2=0 $Y2=0
cc_389 N_A_196_465#_c_354_n N_A_27_465#_M1015_g 0.00228769f $X=1.19 $Y=1.545
+ $X2=0 $Y2=0
cc_390 N_A_196_465#_c_357_n N_A_27_465#_M1015_g 0.0124206f $X=1.2 $Y=1.295 $X2=0
+ $Y2=0
cc_391 N_A_196_465#_M1002_g N_A_27_465#_c_891_n 0.0103073f $X=2.355 $Y=2.525
+ $X2=0 $Y2=0
cc_392 N_A_196_465#_c_368_n N_A_27_465#_c_891_n 0.00388788f $X=1.13 $Y=2.48
+ $X2=0 $Y2=0
cc_393 N_A_196_465#_c_351_n N_A_27_465#_c_881_n 0.00487016f $X=1.19 $Y=0.58
+ $X2=0 $Y2=0
cc_394 N_A_196_465#_M1031_g N_A_27_465#_M1029_g 0.0159729f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_395 N_A_196_465#_c_350_n N_A_27_465#_M1029_g 0.00474437f $X=2.355 $Y=1.68
+ $X2=0 $Y2=0
cc_396 N_A_196_465#_M1002_g N_A_27_465#_M1019_g 0.0136812f $X=2.355 $Y=2.525
+ $X2=0 $Y2=0
cc_397 N_A_196_465#_c_346_n N_A_27_465#_M1019_g 0.00265396f $X=2.785 $Y=1.435
+ $X2=0 $Y2=0
cc_398 N_A_196_465#_M1014_g N_A_27_465#_c_894_n 0.00363882f $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_399 N_A_196_465#_M1030_g N_A_27_465#_M1032_g 0.025054f $X=5.715 $Y=0.555
+ $X2=0 $Y2=0
cc_400 N_A_196_465#_c_359_n N_A_27_465#_M1032_g 4.84017e-19 $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_401 N_A_196_465#_c_360_n N_A_27_465#_M1032_g 0.0102558f $X=5.715 $Y=1.51
+ $X2=0 $Y2=0
cc_402 N_A_196_465#_M1014_g N_A_27_465#_M1026_g 0.014683f $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_403 N_A_196_465#_M1014_g N_A_27_465#_c_898_n 0.0102558f $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_404 N_A_196_465#_c_369_n N_A_27_465#_c_899_n 0.0140367f $X=1.13 $Y=2.315
+ $X2=0 $Y2=0
cc_405 N_A_196_465#_c_354_n N_A_27_465#_c_886_n 0.00476801f $X=1.19 $Y=1.545
+ $X2=0 $Y2=0
cc_406 N_A_196_465#_c_369_n N_A_27_465#_c_886_n 0.0137158f $X=1.13 $Y=2.315
+ $X2=0 $Y2=0
cc_407 N_A_196_465#_c_354_n N_A_27_465#_c_889_n 0.00680892f $X=1.19 $Y=1.545
+ $X2=0 $Y2=0
cc_408 N_A_196_465#_c_369_n N_A_27_465#_c_889_n 0.00502547f $X=1.13 $Y=2.315
+ $X2=0 $Y2=0
cc_409 N_A_196_465#_M1030_g N_A_1158_47#_c_1128_n 0.00983419f $X=5.715 $Y=0.555
+ $X2=0 $Y2=0
cc_410 N_A_196_465#_M1030_g N_A_1158_47#_c_1130_n 0.00561444f $X=5.715 $Y=0.555
+ $X2=0 $Y2=0
cc_411 N_A_196_465#_c_360_n N_A_1158_47#_c_1130_n 0.00345798f $X=5.715 $Y=1.51
+ $X2=0 $Y2=0
cc_412 N_A_196_465#_M1014_g N_A_1158_47#_c_1146_n 0.0019096f $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_413 N_A_196_465#_M1014_g N_A_1158_47#_c_1147_n 2.05438e-19 $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_414 N_A_196_465#_c_367_n N_VPWR_c_1328_n 0.00176027f $X=1.13 $Y=2.42 $X2=0
+ $Y2=0
cc_415 N_A_196_465#_M1002_g N_VPWR_c_1329_n 8.45149e-19 $X=2.355 $Y=2.525 $X2=0
+ $Y2=0
cc_416 N_A_196_465#_c_367_n N_VPWR_c_1329_n 0.0322318f $X=1.13 $Y=2.42 $X2=0
+ $Y2=0
cc_417 N_A_196_465#_c_368_n N_VPWR_c_1345_n 0.00946276f $X=1.13 $Y=2.48 $X2=0
+ $Y2=0
cc_418 N_A_196_465#_M1002_g N_VPWR_c_1327_n 9.39239e-19 $X=2.355 $Y=2.525 $X2=0
+ $Y2=0
cc_419 N_A_196_465#_c_368_n N_VPWR_c_1327_n 0.00687052f $X=1.13 $Y=2.48 $X2=0
+ $Y2=0
cc_420 N_A_196_465#_M1002_g N_A_400_119#_c_1468_n 5.87696e-19 $X=2.355 $Y=2.525
+ $X2=0 $Y2=0
cc_421 N_A_196_465#_M1002_g N_A_400_119#_c_1466_n 0.00938663f $X=2.355 $Y=2.525
+ $X2=0 $Y2=0
cc_422 N_A_196_465#_c_345_n N_A_400_119#_c_1466_n 0.0038976f $X=2.67 $Y=1.59
+ $X2=0 $Y2=0
cc_423 N_A_196_465#_c_346_n N_A_400_119#_c_1466_n 5.25656e-19 $X=2.785 $Y=1.435
+ $X2=0 $Y2=0
cc_424 N_A_196_465#_M1031_g N_A_400_119#_c_1466_n 0.00124016f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_425 N_A_196_465#_c_350_n N_A_400_119#_c_1466_n 0.0121057f $X=2.355 $Y=1.68
+ $X2=0 $Y2=0
cc_426 N_A_196_465#_c_355_n N_A_400_119#_c_1466_n 0.0270041f $X=2.035 $Y=1.545
+ $X2=0 $Y2=0
cc_427 N_A_196_465#_c_356_n N_A_400_119#_c_1466_n 0.0149103f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_428 N_A_196_465#_M1031_g N_A_400_119#_c_1467_n 5.44279e-19 $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_429 N_A_196_465#_c_349_n N_A_400_119#_c_1467_n 0.00581449f $X=2.28 $Y=1.68
+ $X2=0 $Y2=0
cc_430 N_A_196_465#_c_355_n N_A_400_119#_c_1467_n 0.00393626f $X=2.035 $Y=1.545
+ $X2=0 $Y2=0
cc_431 N_A_196_465#_c_356_n N_A_400_119#_c_1467_n 0.0141352f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_432 N_A_196_465#_c_357_n N_A_400_119#_c_1467_n 0.00517047f $X=1.2 $Y=1.295
+ $X2=0 $Y2=0
cc_433 N_A_196_465#_M1002_g N_A_400_119#_c_1470_n 0.0119027f $X=2.355 $Y=2.525
+ $X2=0 $Y2=0
cc_434 N_A_196_465#_c_349_n N_A_400_119#_c_1470_n 0.00587315f $X=2.28 $Y=1.68
+ $X2=0 $Y2=0
cc_435 N_A_196_465#_c_355_n N_A_400_119#_c_1470_n 0.00452194f $X=2.035 $Y=1.545
+ $X2=0 $Y2=0
cc_436 N_A_196_465#_M1014_g N_A_988_379#_c_1511_n 0.00247834f $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_437 N_A_196_465#_M1014_g N_A_988_379#_c_1513_n 5.20259e-19 $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_438 N_A_196_465#_M1014_g N_A_1095_425#_c_1541_n 0.0124267f $X=5.815 $Y=2.335
+ $X2=0 $Y2=0
cc_439 N_A_196_465#_c_351_n N_VGND_c_1580_n 0.0419374f $X=1.19 $Y=0.58 $X2=0
+ $Y2=0
cc_440 N_A_196_465#_c_352_n N_VGND_c_1580_n 0.00456279f $X=1.945 $Y=1.545 $X2=0
+ $Y2=0
cc_441 N_A_196_465#_c_356_n N_VGND_c_1580_n 0.00736547f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_442 N_A_196_465#_M1031_g N_VGND_c_1581_n 0.00135348f $X=2.785 $Y=0.805 $X2=0
+ $Y2=0
cc_443 N_A_196_465#_c_356_n N_VGND_c_1581_n 0.0010845f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_444 N_A_196_465#_c_356_n N_VGND_c_1582_n 0.0131412f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_445 N_A_196_465#_M1031_g N_VGND_c_1588_n 0.00361554f $X=2.785 $Y=0.805 $X2=0
+ $Y2=0
cc_446 N_A_196_465#_M1030_g N_VGND_c_1590_n 0.00579312f $X=5.715 $Y=0.555 $X2=0
+ $Y2=0
cc_447 N_A_196_465#_c_351_n N_VGND_c_1593_n 0.00906443f $X=1.19 $Y=0.58 $X2=0
+ $Y2=0
cc_448 N_A_196_465#_M1031_g N_VGND_c_1601_n 0.00477801f $X=2.785 $Y=0.805 $X2=0
+ $Y2=0
cc_449 N_A_196_465#_M1030_g N_VGND_c_1601_n 0.0118663f $X=5.715 $Y=0.555 $X2=0
+ $Y2=0
cc_450 N_A_196_465#_c_351_n N_VGND_c_1601_n 0.0087406f $X=1.19 $Y=0.58 $X2=0
+ $Y2=0
cc_451 N_A_196_465#_c_353_n N_VGND_c_1601_n 0.00163715f $X=1.19 $Y=1.005 $X2=0
+ $Y2=0
cc_452 N_A_614_93#_c_536_n N_SET_B_M1025_g 0.00306762f $X=3.72 $Y=2.36 $X2=0
+ $Y2=0
cc_453 N_A_614_93#_c_526_n N_SET_B_c_614_n 0.0142998f $X=3.785 $Y=1.1 $X2=0
+ $Y2=0
cc_454 N_A_614_93#_c_527_n N_SET_B_c_614_n 0.00226176f $X=3.87 $Y=1.015 $X2=0
+ $Y2=0
cc_455 N_A_614_93#_c_534_n N_SET_B_c_625_n 0.02221f $X=3.635 $Y=2.025 $X2=0
+ $Y2=0
cc_456 N_A_614_93#_c_553_p N_SET_B_c_625_n 9.0634e-19 $X=3.9 $Y=2.525 $X2=0
+ $Y2=0
cc_457 N_A_614_93#_c_534_n N_SET_B_c_626_n 9.85655e-19 $X=3.635 $Y=2.025 $X2=0
+ $Y2=0
cc_458 N_A_614_93#_M1023_g N_A_486_119#_M1003_g 0.0137271f $X=3.145 $Y=2.525
+ $X2=0 $Y2=0
cc_459 N_A_614_93#_c_534_n N_A_486_119#_M1003_g 0.0098221f $X=3.635 $Y=2.025
+ $X2=0 $Y2=0
cc_460 N_A_614_93#_c_535_n N_A_486_119#_M1003_g 0.0217225f $X=3.235 $Y=1.99
+ $X2=0 $Y2=0
cc_461 N_A_614_93#_c_536_n N_A_486_119#_M1003_g 0.00684915f $X=3.72 $Y=2.36
+ $X2=0 $Y2=0
cc_462 N_A_614_93#_c_553_p N_A_486_119#_M1003_g 0.00788693f $X=3.9 $Y=2.525
+ $X2=0 $Y2=0
cc_463 N_A_614_93#_c_526_n N_A_486_119#_M1020_g 0.00132115f $X=3.785 $Y=1.1
+ $X2=0 $Y2=0
cc_464 N_A_614_93#_c_527_n N_A_486_119#_M1020_g 0.0124088f $X=3.87 $Y=1.015
+ $X2=0 $Y2=0
cc_465 N_A_614_93#_c_526_n N_A_486_119#_c_738_n 0.00367835f $X=3.785 $Y=1.1
+ $X2=0 $Y2=0
cc_466 N_A_614_93#_c_528_n N_A_486_119#_c_738_n 9.04406e-19 $X=3.235 $Y=1.1
+ $X2=0 $Y2=0
cc_467 N_A_614_93#_c_529_n N_A_486_119#_c_738_n 0.0120604f $X=3.235 $Y=1.29
+ $X2=0 $Y2=0
cc_468 N_A_614_93#_c_532_n N_A_486_119#_c_738_n 0.0122872f $X=3.235 $Y=1.825
+ $X2=0 $Y2=0
cc_469 N_A_614_93#_c_526_n N_A_486_119#_c_739_n 0.00376802f $X=3.785 $Y=1.1
+ $X2=0 $Y2=0
cc_470 N_A_614_93#_c_530_n N_A_486_119#_c_739_n 0.00238493f $X=3.995 $Y=0.445
+ $X2=0 $Y2=0
cc_471 N_A_614_93#_c_528_n N_A_486_119#_c_743_n 0.0176274f $X=3.235 $Y=1.1 $X2=0
+ $Y2=0
cc_472 N_A_614_93#_c_531_n N_A_486_119#_c_743_n 0.00324367f $X=3.235 $Y=1.125
+ $X2=0 $Y2=0
cc_473 N_A_614_93#_M1023_g N_A_486_119#_c_748_n 0.00213576f $X=3.145 $Y=2.525
+ $X2=0 $Y2=0
cc_474 N_A_614_93#_c_534_n N_A_486_119#_c_748_n 0.0151879f $X=3.635 $Y=2.025
+ $X2=0 $Y2=0
cc_475 N_A_614_93#_c_535_n N_A_486_119#_c_748_n 0.00171987f $X=3.235 $Y=1.99
+ $X2=0 $Y2=0
cc_476 N_A_614_93#_c_532_n N_A_486_119#_c_748_n 0.00374574f $X=3.235 $Y=1.825
+ $X2=0 $Y2=0
cc_477 N_A_614_93#_c_534_n N_A_486_119#_c_744_n 0.0391835f $X=3.635 $Y=2.025
+ $X2=0 $Y2=0
cc_478 N_A_614_93#_c_535_n N_A_486_119#_c_744_n 0.00150916f $X=3.235 $Y=1.99
+ $X2=0 $Y2=0
cc_479 N_A_614_93#_c_526_n N_A_486_119#_c_744_n 0.00493245f $X=3.785 $Y=1.1
+ $X2=0 $Y2=0
cc_480 N_A_614_93#_c_528_n N_A_486_119#_c_744_n 0.0223028f $X=3.235 $Y=1.1 $X2=0
+ $Y2=0
cc_481 N_A_614_93#_c_529_n N_A_486_119#_c_744_n 0.0015229f $X=3.235 $Y=1.29
+ $X2=0 $Y2=0
cc_482 N_A_614_93#_c_532_n N_A_486_119#_c_744_n 0.0110778f $X=3.235 $Y=1.825
+ $X2=0 $Y2=0
cc_483 N_A_614_93#_c_531_n N_A_486_119#_c_775_n 6.75672e-19 $X=3.235 $Y=1.125
+ $X2=0 $Y2=0
cc_484 N_A_614_93#_c_534_n N_A_486_119#_c_745_n 0.0146482f $X=3.635 $Y=2.025
+ $X2=0 $Y2=0
cc_485 N_A_614_93#_c_526_n N_A_486_119#_c_745_n 0.0214261f $X=3.785 $Y=1.1 $X2=0
+ $Y2=0
cc_486 N_A_614_93#_c_528_n N_A_486_119#_c_745_n 0.00174661f $X=3.235 $Y=1.1
+ $X2=0 $Y2=0
cc_487 N_A_614_93#_c_529_n N_A_486_119#_c_745_n 5.95896e-19 $X=3.235 $Y=1.29
+ $X2=0 $Y2=0
cc_488 N_A_614_93#_c_553_p N_A_486_119#_c_745_n 0.00426527f $X=3.9 $Y=2.525
+ $X2=0 $Y2=0
cc_489 N_A_614_93#_c_532_n N_A_486_119#_c_745_n 6.81521e-19 $X=3.235 $Y=1.825
+ $X2=0 $Y2=0
cc_490 N_A_614_93#_M1023_g N_A_27_465#_M1019_g 0.0396153f $X=3.145 $Y=2.525
+ $X2=0 $Y2=0
cc_491 N_A_614_93#_M1023_g N_A_27_465#_c_894_n 0.0103107f $X=3.145 $Y=2.525
+ $X2=0 $Y2=0
cc_492 N_A_614_93#_c_553_p N_A_27_465#_c_894_n 0.00429322f $X=3.9 $Y=2.525 $X2=0
+ $Y2=0
cc_493 N_A_614_93#_M1023_g N_VPWR_c_1330_n 0.00997303f $X=3.145 $Y=2.525 $X2=0
+ $Y2=0
cc_494 N_A_614_93#_c_534_n N_VPWR_c_1330_n 0.0167735f $X=3.635 $Y=2.025 $X2=0
+ $Y2=0
cc_495 N_A_614_93#_c_535_n N_VPWR_c_1330_n 0.00392572f $X=3.235 $Y=1.99 $X2=0
+ $Y2=0
cc_496 N_A_614_93#_c_553_p N_VPWR_c_1330_n 0.025364f $X=3.9 $Y=2.525 $X2=0 $Y2=0
cc_497 N_A_614_93#_c_553_p N_VPWR_c_1346_n 0.0057608f $X=3.9 $Y=2.525 $X2=0
+ $Y2=0
cc_498 N_A_614_93#_M1023_g N_VPWR_c_1327_n 7.88961e-19 $X=3.145 $Y=2.525 $X2=0
+ $Y2=0
cc_499 N_A_614_93#_c_553_p N_VPWR_c_1327_n 0.0089445f $X=3.9 $Y=2.525 $X2=0
+ $Y2=0
cc_500 N_A_614_93#_c_532_n N_A_400_119#_c_1466_n 3.36115e-19 $X=3.235 $Y=1.825
+ $X2=0 $Y2=0
cc_501 N_A_614_93#_c_528_n N_VGND_M1021_d 0.00194443f $X=3.235 $Y=1.1 $X2=0
+ $Y2=0
cc_502 N_A_614_93#_c_526_n N_VGND_c_1581_n 0.00972467f $X=3.785 $Y=1.1 $X2=0
+ $Y2=0
cc_503 N_A_614_93#_c_527_n N_VGND_c_1581_n 0.0138628f $X=3.87 $Y=1.015 $X2=0
+ $Y2=0
cc_504 N_A_614_93#_c_528_n N_VGND_c_1581_n 0.0140943f $X=3.235 $Y=1.1 $X2=0
+ $Y2=0
cc_505 N_A_614_93#_c_529_n N_VGND_c_1581_n 9.37087e-19 $X=3.235 $Y=1.29 $X2=0
+ $Y2=0
cc_506 N_A_614_93#_c_530_n N_VGND_c_1581_n 0.0203137f $X=3.995 $Y=0.445 $X2=0
+ $Y2=0
cc_507 N_A_614_93#_c_531_n N_VGND_c_1581_n 0.00939839f $X=3.235 $Y=1.125 $X2=0
+ $Y2=0
cc_508 N_A_614_93#_c_531_n N_VGND_c_1588_n 0.0035863f $X=3.235 $Y=1.125 $X2=0
+ $Y2=0
cc_509 N_A_614_93#_c_530_n N_VGND_c_1594_n 0.0175354f $X=3.995 $Y=0.445 $X2=0
+ $Y2=0
cc_510 N_A_614_93#_M1020_s N_VGND_c_1601_n 0.00338576f $X=3.87 $Y=0.235 $X2=0
+ $Y2=0
cc_511 N_A_614_93#_c_530_n N_VGND_c_1601_n 0.0118544f $X=3.995 $Y=0.445 $X2=0
+ $Y2=0
cc_512 N_A_614_93#_c_531_n N_VGND_c_1601_n 0.00401353f $X=3.235 $Y=1.125 $X2=0
+ $Y2=0
cc_513 N_SET_B_M1025_g N_A_486_119#_M1003_g 0.0132585f $X=4.115 $Y=2.525 $X2=0
+ $Y2=0
cc_514 N_SET_B_c_613_n N_A_486_119#_M1003_g 0.00158966f $X=4.22 $Y=1.765 $X2=0
+ $Y2=0
cc_515 N_SET_B_c_625_n N_A_486_119#_M1003_g 0.00260812f $X=4.14 $Y=1.85 $X2=0
+ $Y2=0
cc_516 N_SET_B_c_626_n N_A_486_119#_M1003_g 0.0208161f $X=4.14 $Y=1.99 $X2=0
+ $Y2=0
cc_517 N_SET_B_M1010_g N_A_486_119#_M1020_g 0.0712652f $X=4.57 $Y=0.445 $X2=0
+ $Y2=0
cc_518 N_SET_B_c_613_n N_A_486_119#_M1020_g 0.0021502f $X=4.22 $Y=1.765 $X2=0
+ $Y2=0
cc_519 N_SET_B_c_614_n N_A_486_119#_M1020_g 0.0142452f $X=4.305 $Y=1.11 $X2=0
+ $Y2=0
cc_520 N_SET_B_c_613_n N_A_486_119#_c_734_n 0.00705388f $X=4.22 $Y=1.765 $X2=0
+ $Y2=0
cc_521 N_SET_B_c_615_n N_A_486_119#_c_734_n 0.00427031f $X=4.66 $Y=1.07 $X2=0
+ $Y2=0
cc_522 N_SET_B_c_616_n N_A_486_119#_c_734_n 0.0194496f $X=4.66 $Y=1.07 $X2=0
+ $Y2=0
cc_523 N_SET_B_c_629_n N_A_486_119#_c_734_n 0.0097655f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_524 N_SET_B_M1025_g N_A_486_119#_M1000_g 0.00413416f $X=4.115 $Y=2.525 $X2=0
+ $Y2=0
cc_525 N_SET_B_c_613_n N_A_486_119#_M1000_g 0.00366457f $X=4.22 $Y=1.765 $X2=0
+ $Y2=0
cc_526 N_SET_B_c_625_n N_A_486_119#_M1000_g 8.41149e-19 $X=4.14 $Y=1.85 $X2=0
+ $Y2=0
cc_527 N_SET_B_c_626_n N_A_486_119#_M1000_g 0.00585973f $X=4.14 $Y=1.99 $X2=0
+ $Y2=0
cc_528 N_SET_B_c_629_n N_A_486_119#_M1000_g 0.0183151f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_529 N_SET_B_M1010_g N_A_486_119#_c_737_n 0.010362f $X=4.57 $Y=0.445 $X2=0
+ $Y2=0
cc_530 N_SET_B_c_616_n N_A_486_119#_c_737_n 0.00276406f $X=4.66 $Y=1.07 $X2=0
+ $Y2=0
cc_531 N_SET_B_c_625_n N_A_486_119#_c_739_n 9.70937e-19 $X=4.14 $Y=1.85 $X2=0
+ $Y2=0
cc_532 N_SET_B_c_626_n N_A_486_119#_c_739_n 0.0222405f $X=4.14 $Y=1.99 $X2=0
+ $Y2=0
cc_533 N_SET_B_c_613_n N_A_486_119#_c_740_n 0.0138811f $X=4.22 $Y=1.765 $X2=0
+ $Y2=0
cc_534 N_SET_B_c_629_n N_A_486_119#_c_741_n 0.0102433f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_535 N_SET_B_c_615_n N_A_486_119#_c_742_n 0.00165723f $X=4.66 $Y=1.07 $X2=0
+ $Y2=0
cc_536 N_SET_B_c_616_n N_A_486_119#_c_742_n 0.0155743f $X=4.66 $Y=1.07 $X2=0
+ $Y2=0
cc_537 N_SET_B_c_629_n N_A_486_119#_c_742_n 0.0052455f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_538 N_SET_B_c_613_n N_A_486_119#_c_745_n 0.0249711f $X=4.22 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_SET_B_M1025_g N_A_27_465#_c_894_n 0.0103107f $X=4.115 $Y=2.525 $X2=0
+ $Y2=0
cc_540 SET_B N_A_27_465#_M1032_g 0.0255555f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_541 SET_B N_A_27_465#_c_898_n 5.81983e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_542 SET_B N_A_27_465#_c_898_n 0.00781572f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_543 N_SET_B_c_611_n N_A_1309_65#_M1001_g 0.0616632f $X=6.98 $Y=0.985 $X2=0
+ $Y2=0
cc_544 SET_B N_A_1309_65#_M1001_g 0.0113292f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_545 N_SET_B_c_621_n N_A_1309_65#_c_1024_n 0.0142318f $X=7.45 $Y=1.84 $X2=0
+ $Y2=0
cc_546 SET_B N_A_1309_65#_c_1024_n 0.0133433f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_547 N_SET_B_c_621_n N_A_1309_65#_M1008_g 0.00687352f $X=7.45 $Y=1.84 $X2=0
+ $Y2=0
cc_548 N_SET_B_M1033_g N_A_1309_65#_M1008_g 0.0145768f $X=7.865 $Y=2.525 $X2=0
+ $Y2=0
cc_549 N_SET_B_M1033_g N_A_1309_65#_c_1034_n 0.0104164f $X=7.865 $Y=2.525 $X2=0
+ $Y2=0
cc_550 N_SET_B_c_612_n N_A_1309_65#_c_1025_n 0.0142318f $X=7.285 $Y=1.765 $X2=0
+ $Y2=0
cc_551 SET_B N_A_1309_65#_c_1025_n 0.0161978f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_552 SET_B N_A_1309_65#_c_1035_n 7.29045e-19 $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_553 N_SET_B_c_611_n N_A_1158_47#_c_1117_n 0.00129316f $X=6.98 $Y=0.985 $X2=0
+ $Y2=0
cc_554 SET_B N_A_1158_47#_c_1117_n 0.0010573f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_555 N_SET_B_c_611_n N_A_1158_47#_c_1119_n 0.0129783f $X=6.98 $Y=0.985 $X2=0
+ $Y2=0
cc_556 N_SET_B_c_620_n N_A_1158_47#_M1004_g 0.00281367f $X=7.79 $Y=1.84 $X2=0
+ $Y2=0
cc_557 N_SET_B_c_611_n N_A_1158_47#_c_1129_n 0.0256118f $X=6.98 $Y=0.985 $X2=0
+ $Y2=0
cc_558 SET_B N_A_1158_47#_c_1129_n 0.104553f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_559 SET_B N_A_1158_47#_c_1130_n 0.0168526f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_560 N_SET_B_c_621_n N_A_1158_47#_c_1142_n 0.0147811f $X=7.45 $Y=1.84 $X2=0
+ $Y2=0
cc_561 N_SET_B_M1033_g N_A_1158_47#_c_1142_n 0.0208212f $X=7.865 $Y=2.525 $X2=0
+ $Y2=0
cc_562 N_SET_B_M1033_g N_A_1158_47#_c_1143_n 0.00236895f $X=7.865 $Y=2.525 $X2=0
+ $Y2=0
cc_563 N_SET_B_c_611_n N_A_1158_47#_c_1131_n 0.00109841f $X=6.98 $Y=0.985 $X2=0
+ $Y2=0
cc_564 SET_B N_A_1158_47#_c_1131_n 0.0124658f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_565 N_SET_B_c_620_n N_A_1158_47#_c_1132_n 0.0081128f $X=7.79 $Y=1.84 $X2=0
+ $Y2=0
cc_566 N_SET_B_c_612_n N_A_1158_47#_c_1132_n 0.00133781f $X=7.285 $Y=1.765 $X2=0
+ $Y2=0
cc_567 SET_B N_A_1158_47#_c_1132_n 0.0231056f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_568 SET_B N_A_1158_47#_c_1146_n 0.0137944f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_569 SET_B N_A_1158_47#_c_1146_n 0.0131177f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_570 SET_B N_A_1158_47#_c_1147_n 0.106437f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_571 SET_B N_A_1158_47#_c_1133_n 9.21238e-19 $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_572 N_SET_B_c_629_n N_VPWR_M1025_d 0.00239457f $X=5.905 $Y=1.59 $X2=0 $Y2=0
cc_573 N_SET_B_M1025_g N_VPWR_c_1331_n 0.00771243f $X=4.115 $Y=2.525 $X2=0 $Y2=0
cc_574 N_SET_B_c_625_n N_VPWR_c_1331_n 0.0119932f $X=4.14 $Y=1.85 $X2=0 $Y2=0
cc_575 N_SET_B_c_626_n N_VPWR_c_1331_n 8.95726e-19 $X=4.14 $Y=1.99 $X2=0 $Y2=0
cc_576 N_SET_B_c_629_n N_VPWR_c_1331_n 0.0279874f $X=5.905 $Y=1.59 $X2=0 $Y2=0
cc_577 N_SET_B_M1025_g N_VPWR_c_1332_n 0.00643939f $X=4.115 $Y=2.525 $X2=0 $Y2=0
cc_578 N_SET_B_M1033_g N_VPWR_c_1333_n 0.001816f $X=7.865 $Y=2.525 $X2=0 $Y2=0
cc_579 N_SET_B_M1033_g N_VPWR_c_1335_n 0.00423915f $X=7.865 $Y=2.525 $X2=0 $Y2=0
cc_580 N_SET_B_M1025_g N_VPWR_c_1327_n 7.88961e-19 $X=4.115 $Y=2.525 $X2=0 $Y2=0
cc_581 N_SET_B_M1033_g N_VPWR_c_1327_n 9.39239e-19 $X=7.865 $Y=2.525 $X2=0 $Y2=0
cc_582 N_SET_B_c_629_n N_A_988_379#_M1000_d 0.00239457f $X=5.905 $Y=1.59
+ $X2=-0.19 $Y2=-0.245
cc_583 N_SET_B_c_629_n N_A_988_379#_c_1511_n 0.0220026f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_584 N_SET_B_c_629_n N_A_1095_425#_c_1538_n 0.0166593f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_585 N_SET_B_c_629_n N_A_1095_425#_c_1541_n 0.00478688f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_586 N_SET_B_M1010_g N_VGND_c_1582_n 0.0162508f $X=4.57 $Y=0.445 $X2=0 $Y2=0
cc_587 N_SET_B_c_611_n N_VGND_c_1583_n 0.00961495f $X=6.98 $Y=0.985 $X2=0 $Y2=0
cc_588 N_SET_B_c_611_n N_VGND_c_1590_n 0.00429764f $X=6.98 $Y=0.985 $X2=0 $Y2=0
cc_589 N_SET_B_M1010_g N_VGND_c_1594_n 0.00585385f $X=4.57 $Y=0.445 $X2=0 $Y2=0
cc_590 N_SET_B_M1010_g N_VGND_c_1601_n 0.0115242f $X=4.57 $Y=0.445 $X2=0 $Y2=0
cc_591 N_SET_B_c_611_n N_VGND_c_1601_n 0.00435987f $X=6.98 $Y=0.985 $X2=0 $Y2=0
cc_592 N_A_486_119#_c_748_n N_A_27_465#_c_891_n 0.00330098f $X=2.73 $Y=2.435
+ $X2=0 $Y2=0
cc_593 N_A_486_119#_c_743_n N_A_27_465#_M1029_g 0.00140517f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_594 N_A_486_119#_c_775_n N_A_27_465#_M1029_g 0.00325747f $X=2.73 $Y=0.725
+ $X2=0 $Y2=0
cc_595 N_A_486_119#_c_748_n N_A_27_465#_M1019_g 0.0165265f $X=2.73 $Y=2.435
+ $X2=0 $Y2=0
cc_596 N_A_486_119#_c_744_n N_A_27_465#_M1019_g 8.05699e-19 $X=3.615 $Y=1.64
+ $X2=0 $Y2=0
cc_597 N_A_486_119#_M1003_g N_A_27_465#_c_894_n 0.00989604f $X=3.685 $Y=2.525
+ $X2=0 $Y2=0
cc_598 N_A_486_119#_M1000_g N_A_27_465#_c_894_n 0.0101459f $X=4.865 $Y=2.315
+ $X2=0 $Y2=0
cc_599 N_A_486_119#_c_737_n N_A_1158_47#_c_1128_n 0.00177792f $X=5.355 $Y=0.985
+ $X2=0 $Y2=0
cc_600 N_A_486_119#_c_737_n N_A_1158_47#_c_1130_n 8.31149e-19 $X=5.355 $Y=0.985
+ $X2=0 $Y2=0
cc_601 N_A_486_119#_c_748_n N_VPWR_c_1329_n 5.72484e-19 $X=2.73 $Y=2.435 $X2=0
+ $Y2=0
cc_602 N_A_486_119#_M1003_g N_VPWR_c_1330_n 0.00671009f $X=3.685 $Y=2.525 $X2=0
+ $Y2=0
cc_603 N_A_486_119#_c_748_n N_VPWR_c_1330_n 0.0135336f $X=2.73 $Y=2.435 $X2=0
+ $Y2=0
cc_604 N_A_486_119#_M1003_g N_VPWR_c_1332_n 7.84513e-19 $X=3.685 $Y=2.525 $X2=0
+ $Y2=0
cc_605 N_A_486_119#_M1000_g N_VPWR_c_1332_n 0.00221662f $X=4.865 $Y=2.315 $X2=0
+ $Y2=0
cc_606 N_A_486_119#_c_748_n N_VPWR_c_1341_n 0.00649869f $X=2.73 $Y=2.435 $X2=0
+ $Y2=0
cc_607 N_A_486_119#_M1003_g N_VPWR_c_1327_n 9.39239e-19 $X=3.685 $Y=2.525 $X2=0
+ $Y2=0
cc_608 N_A_486_119#_M1000_g N_VPWR_c_1327_n 7.82699e-19 $X=4.865 $Y=2.315 $X2=0
+ $Y2=0
cc_609 N_A_486_119#_c_748_n N_VPWR_c_1327_n 0.0102727f $X=2.73 $Y=2.435 $X2=0
+ $Y2=0
cc_610 N_A_486_119#_c_748_n N_A_400_119#_c_1468_n 0.00431258f $X=2.73 $Y=2.435
+ $X2=0 $Y2=0
cc_611 N_A_486_119#_c_743_n N_A_400_119#_c_1466_n 0.0263494f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_612 N_A_486_119#_c_748_n N_A_400_119#_c_1466_n 0.0267202f $X=2.73 $Y=2.435
+ $X2=0 $Y2=0
cc_613 N_A_486_119#_c_750_n N_A_400_119#_c_1466_n 0.012867f $X=2.73 $Y=1.64
+ $X2=0 $Y2=0
cc_614 N_A_486_119#_c_743_n N_A_400_119#_c_1467_n 0.0127469f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_615 N_A_486_119#_c_775_n N_A_400_119#_c_1467_n 0.00160576f $X=2.73 $Y=0.725
+ $X2=0 $Y2=0
cc_616 N_A_486_119#_c_748_n N_A_400_119#_c_1470_n 0.0161373f $X=2.73 $Y=2.435
+ $X2=0 $Y2=0
cc_617 N_A_486_119#_M1000_g N_A_988_379#_c_1511_n 0.0108812f $X=4.865 $Y=2.315
+ $X2=0 $Y2=0
cc_618 N_A_486_119#_M1000_g N_A_988_379#_c_1512_n 5.13126e-19 $X=4.865 $Y=2.315
+ $X2=0 $Y2=0
cc_619 N_A_486_119#_M1000_g N_A_1095_425#_c_1538_n 5.36524e-19 $X=4.865 $Y=2.315
+ $X2=0 $Y2=0
cc_620 N_A_486_119#_M1020_g N_VGND_c_1581_n 0.00331497f $X=4.21 $Y=0.445 $X2=0
+ $Y2=0
cc_621 N_A_486_119#_c_743_n N_VGND_c_1581_n 3.7393e-19 $X=2.73 $Y=1.555 $X2=0
+ $Y2=0
cc_622 N_A_486_119#_c_775_n N_VGND_c_1581_n 0.00873321f $X=2.73 $Y=0.725 $X2=0
+ $Y2=0
cc_623 N_A_486_119#_c_737_n N_VGND_c_1582_n 0.00813089f $X=5.355 $Y=0.985 $X2=0
+ $Y2=0
cc_624 N_A_486_119#_c_741_n N_VGND_c_1582_n 0.00142195f $X=5.11 $Y=1.54 $X2=0
+ $Y2=0
cc_625 N_A_486_119#_c_742_n N_VGND_c_1582_n 0.00872797f $X=5.355 $Y=1.06 $X2=0
+ $Y2=0
cc_626 N_A_486_119#_c_775_n N_VGND_c_1588_n 0.00650647f $X=2.73 $Y=0.725 $X2=0
+ $Y2=0
cc_627 N_A_486_119#_c_737_n N_VGND_c_1590_n 0.00585385f $X=5.355 $Y=0.985 $X2=0
+ $Y2=0
cc_628 N_A_486_119#_M1020_g N_VGND_c_1594_n 0.00585385f $X=4.21 $Y=0.445 $X2=0
+ $Y2=0
cc_629 N_A_486_119#_M1020_g N_VGND_c_1601_n 0.0122126f $X=4.21 $Y=0.445 $X2=0
+ $Y2=0
cc_630 N_A_486_119#_c_737_n N_VGND_c_1601_n 0.0114039f $X=5.355 $Y=0.985 $X2=0
+ $Y2=0
cc_631 N_A_486_119#_c_775_n N_VGND_c_1601_n 0.0117564f $X=2.73 $Y=0.725 $X2=0
+ $Y2=0
cc_632 N_A_27_465#_M1032_g N_A_1309_65#_M1001_g 0.0822724f $X=6.26 $Y=0.665
+ $X2=0 $Y2=0
cc_633 N_A_27_465#_M1032_g N_A_1309_65#_c_1024_n 0.00602247f $X=6.26 $Y=0.665
+ $X2=0 $Y2=0
cc_634 N_A_27_465#_c_898_n N_A_1309_65#_c_1024_n 0.00893821f $X=6.36 $Y=1.94
+ $X2=0 $Y2=0
cc_635 N_A_27_465#_M1026_g N_A_1309_65#_c_1030_n 0.0131346f $X=6.36 $Y=2.545
+ $X2=0 $Y2=0
cc_636 N_A_27_465#_c_894_n N_A_1309_65#_c_1032_n 0.0131346f $X=6.285 $Y=3.15
+ $X2=0 $Y2=0
cc_637 N_A_27_465#_M1026_g N_A_1309_65#_c_1035_n 0.00893821f $X=6.36 $Y=2.545
+ $X2=0 $Y2=0
cc_638 N_A_27_465#_M1032_g N_A_1158_47#_c_1128_n 0.0151038f $X=6.26 $Y=0.665
+ $X2=0 $Y2=0
cc_639 N_A_27_465#_M1032_g N_A_1158_47#_c_1129_n 0.0150297f $X=6.26 $Y=0.665
+ $X2=0 $Y2=0
cc_640 N_A_27_465#_M1026_g N_A_1158_47#_c_1142_n 0.00613732f $X=6.36 $Y=2.545
+ $X2=0 $Y2=0
cc_641 N_A_27_465#_c_898_n N_A_1158_47#_c_1146_n 0.00205897f $X=6.36 $Y=1.94
+ $X2=0 $Y2=0
cc_642 N_A_27_465#_M1026_g N_A_1158_47#_c_1147_n 0.00498662f $X=6.36 $Y=2.545
+ $X2=0 $Y2=0
cc_643 N_A_27_465#_c_898_n N_A_1158_47#_c_1147_n 8.90692e-19 $X=6.36 $Y=1.94
+ $X2=0 $Y2=0
cc_644 N_A_27_465#_M1024_g N_VPWR_c_1328_n 0.00803159f $X=0.905 $Y=2.645 $X2=0
+ $Y2=0
cc_645 N_A_27_465#_c_899_n N_VPWR_c_1328_n 0.00119148f $X=0.26 $Y=2.47 $X2=0
+ $Y2=0
cc_646 N_A_27_465#_c_886_n N_VPWR_c_1328_n 0.00781344f $X=0.68 $Y=1.66 $X2=0
+ $Y2=0
cc_647 N_A_27_465#_c_889_n N_VPWR_c_1328_n 0.0039271f $X=0.975 $Y=1.66 $X2=0
+ $Y2=0
cc_648 N_A_27_465#_M1024_g N_VPWR_c_1329_n 0.00355852f $X=0.905 $Y=2.645 $X2=0
+ $Y2=0
cc_649 N_A_27_465#_c_891_n N_VPWR_c_1329_n 0.0257254f $X=2.71 $Y=3.15 $X2=0
+ $Y2=0
cc_650 N_A_27_465#_M1019_g N_VPWR_c_1330_n 0.00805374f $X=2.785 $Y=2.525 $X2=0
+ $Y2=0
cc_651 N_A_27_465#_c_894_n N_VPWR_c_1330_n 0.0223422f $X=6.285 $Y=3.15 $X2=0
+ $Y2=0
cc_652 N_A_27_465#_c_894_n N_VPWR_c_1332_n 0.0398672f $X=6.285 $Y=3.15 $X2=0
+ $Y2=0
cc_653 N_A_27_465#_c_899_n N_VPWR_c_1339_n 0.0119419f $X=0.26 $Y=2.47 $X2=0
+ $Y2=0
cc_654 N_A_27_465#_c_891_n N_VPWR_c_1341_n 0.0413023f $X=2.71 $Y=3.15 $X2=0
+ $Y2=0
cc_655 N_A_27_465#_c_894_n N_VPWR_c_1343_n 0.0378727f $X=6.285 $Y=3.15 $X2=0
+ $Y2=0
cc_656 N_A_27_465#_c_892_n N_VPWR_c_1345_n 0.0231877f $X=0.98 $Y=3.15 $X2=0
+ $Y2=0
cc_657 N_A_27_465#_c_894_n N_VPWR_c_1346_n 0.0208443f $X=6.285 $Y=3.15 $X2=0
+ $Y2=0
cc_658 N_A_27_465#_c_891_n N_VPWR_c_1327_n 0.0507022f $X=2.71 $Y=3.15 $X2=0
+ $Y2=0
cc_659 N_A_27_465#_c_892_n N_VPWR_c_1327_n 0.0113264f $X=0.98 $Y=3.15 $X2=0
+ $Y2=0
cc_660 N_A_27_465#_c_894_n N_VPWR_c_1327_n 0.0836632f $X=6.285 $Y=3.15 $X2=0
+ $Y2=0
cc_661 N_A_27_465#_c_897_n N_VPWR_c_1327_n 0.00577283f $X=2.785 $Y=3.15 $X2=0
+ $Y2=0
cc_662 N_A_27_465#_c_899_n N_VPWR_c_1327_n 0.0100524f $X=0.26 $Y=2.47 $X2=0
+ $Y2=0
cc_663 N_A_27_465#_c_881_n N_A_400_119#_c_1502_n 0.0030764f $X=2.28 $Y=0.18
+ $X2=0 $Y2=0
cc_664 N_A_27_465#_c_891_n N_A_400_119#_c_1468_n 0.00339216f $X=2.71 $Y=3.15
+ $X2=0 $Y2=0
cc_665 N_A_27_465#_M1029_g N_A_400_119#_c_1466_n 4.46536e-19 $X=2.355 $Y=0.805
+ $X2=0 $Y2=0
cc_666 N_A_27_465#_M1029_g N_A_400_119#_c_1467_n 0.0106397f $X=2.355 $Y=0.805
+ $X2=0 $Y2=0
cc_667 N_A_27_465#_M1019_g N_A_400_119#_c_1470_n 2.52175e-19 $X=2.785 $Y=2.525
+ $X2=0 $Y2=0
cc_668 N_A_27_465#_c_894_n N_A_988_379#_c_1512_n 0.0076867f $X=6.285 $Y=3.15
+ $X2=0 $Y2=0
cc_669 N_A_27_465#_c_894_n N_A_988_379#_c_1513_n 0.0201126f $X=6.285 $Y=3.15
+ $X2=0 $Y2=0
cc_670 N_A_27_465#_M1026_g N_A_988_379#_c_1513_n 0.0140139f $X=6.36 $Y=2.545
+ $X2=0 $Y2=0
cc_671 N_A_27_465#_M1026_g N_A_1095_425#_c_1541_n 0.012067f $X=6.36 $Y=2.545
+ $X2=0 $Y2=0
cc_672 N_A_27_465#_M1015_g N_VGND_c_1579_n 0.00707758f $X=0.975 $Y=0.58 $X2=0
+ $Y2=0
cc_673 N_A_27_465#_c_882_n N_VGND_c_1579_n 0.00606728f $X=1.05 $Y=0.18 $X2=0
+ $Y2=0
cc_674 N_A_27_465#_M1015_g N_VGND_c_1580_n 0.00340903f $X=0.975 $Y=0.58 $X2=0
+ $Y2=0
cc_675 N_A_27_465#_c_881_n N_VGND_c_1580_n 0.023215f $X=2.28 $Y=0.18 $X2=0 $Y2=0
cc_676 N_A_27_465#_M1029_g N_VGND_c_1580_n 0.00606057f $X=2.355 $Y=0.805 $X2=0
+ $Y2=0
cc_677 N_A_27_465#_c_881_n N_VGND_c_1588_n 0.0190354f $X=2.28 $Y=0.18 $X2=0
+ $Y2=0
cc_678 N_A_27_465#_M1032_g N_VGND_c_1590_n 0.00517164f $X=6.26 $Y=0.665 $X2=0
+ $Y2=0
cc_679 N_A_27_465#_c_887_n N_VGND_c_1592_n 0.00999822f $X=0.27 $Y=0.575 $X2=0
+ $Y2=0
cc_680 N_A_27_465#_c_882_n N_VGND_c_1593_n 0.0197685f $X=1.05 $Y=0.18 $X2=0
+ $Y2=0
cc_681 N_A_27_465#_c_881_n N_VGND_c_1601_n 0.0432072f $X=2.28 $Y=0.18 $X2=0
+ $Y2=0
cc_682 N_A_27_465#_c_882_n N_VGND_c_1601_n 0.008022f $X=1.05 $Y=0.18 $X2=0 $Y2=0
cc_683 N_A_27_465#_M1032_g N_VGND_c_1601_n 0.00519032f $X=6.26 $Y=0.665 $X2=0
+ $Y2=0
cc_684 N_A_27_465#_c_887_n N_VGND_c_1601_n 0.0109072f $X=0.27 $Y=0.575 $X2=0
+ $Y2=0
cc_685 N_A_1309_65#_c_1028_n N_A_1158_47#_c_1117_n 0.00326045f $X=7.955 $Y=0.57
+ $X2=0 $Y2=0
cc_686 N_A_1309_65#_c_1028_n N_A_1158_47#_c_1118_n 0.0111034f $X=7.955 $Y=0.57
+ $X2=0 $Y2=0
cc_687 N_A_1309_65#_c_1027_n N_A_1158_47#_M1004_g 0.0135177f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_688 N_A_1309_65#_c_1038_n N_A_1158_47#_M1004_g 2.69703e-19 $X=8.9 $Y=2.6
+ $X2=0 $Y2=0
cc_689 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1120_n 0.0159235f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_690 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1122_n 0.00416624f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_691 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1124_n 0.00612735f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_692 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1139_n 5.09626e-19 $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_693 N_A_1309_65#_c_1038_n N_A_1158_47#_c_1139_n 0.00463249f $X=8.9 $Y=2.6
+ $X2=0 $Y2=0
cc_694 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1126_n 0.00235108f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_695 N_A_1309_65#_M1017_d N_A_1158_47#_c_1129_n 0.00226217f $X=7.63 $Y=0.455
+ $X2=0 $Y2=0
cc_696 N_A_1309_65#_M1001_g N_A_1158_47#_c_1129_n 0.0139858f $X=6.62 $Y=0.665
+ $X2=0 $Y2=0
cc_697 N_A_1309_65#_c_1025_n N_A_1158_47#_c_1129_n 8.72004e-19 $X=6.835 $Y=1.55
+ $X2=0 $Y2=0
cc_698 N_A_1309_65#_c_1026_n N_A_1158_47#_c_1129_n 0.00109361f $X=8.735 $Y=0.53
+ $X2=0 $Y2=0
cc_699 N_A_1309_65#_c_1028_n N_A_1158_47#_c_1129_n 0.0204689f $X=7.955 $Y=0.57
+ $X2=0 $Y2=0
cc_700 N_A_1309_65#_c_1024_n N_A_1158_47#_c_1142_n 0.00509456f $X=6.835 $Y=2.155
+ $X2=0 $Y2=0
cc_701 N_A_1309_65#_M1008_g N_A_1158_47#_c_1142_n 0.00984479f $X=7.435 $Y=2.525
+ $X2=0 $Y2=0
cc_702 N_A_1309_65#_c_1025_n N_A_1158_47#_c_1142_n 7.97866e-19 $X=6.835 $Y=1.55
+ $X2=0 $Y2=0
cc_703 N_A_1309_65#_c_1035_n N_A_1158_47#_c_1142_n 0.0110533f $X=6.945 $Y=2.23
+ $X2=0 $Y2=0
cc_704 N_A_1309_65#_c_1034_n N_A_1158_47#_c_1143_n 0.00435665f $X=8.735 $Y=3.15
+ $X2=0 $Y2=0
cc_705 N_A_1309_65#_c_1026_n N_A_1158_47#_c_1131_n 0.0360871f $X=8.735 $Y=0.53
+ $X2=0 $Y2=0
cc_706 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1131_n 0.0482279f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_707 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1132_n 0.00654345f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_708 N_A_1309_65#_c_1035_n N_A_1158_47#_c_1147_n 2.18456e-19 $X=6.945 $Y=2.23
+ $X2=0 $Y2=0
cc_709 N_A_1309_65#_c_1026_n N_A_1158_47#_c_1133_n 0.0244218f $X=8.735 $Y=0.53
+ $X2=0 $Y2=0
cc_710 N_A_1309_65#_c_1027_n N_A_1158_47#_c_1133_n 0.0128966f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_711 N_A_1309_65#_c_1028_n N_A_1158_47#_c_1133_n 0.00183408f $X=7.955 $Y=0.57
+ $X2=0 $Y2=0
cc_712 N_A_1309_65#_c_1026_n N_A_1855_47#_c_1264_n 0.0148637f $X=8.735 $Y=0.53
+ $X2=0 $Y2=0
cc_713 N_A_1309_65#_c_1027_n N_A_1855_47#_c_1264_n 0.0461786f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_714 N_A_1309_65#_c_1027_n N_A_1855_47#_c_1265_n 0.0903849f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_715 N_A_1309_65#_c_1038_n N_A_1855_47#_c_1265_n 0.00174916f $X=8.9 $Y=2.6
+ $X2=0 $Y2=0
cc_716 N_A_1309_65#_c_1027_n N_A_1855_47#_c_1267_n 0.0285593f $X=8.88 $Y=1.835
+ $X2=0 $Y2=0
cc_717 N_A_1309_65#_M1008_g N_VPWR_c_1333_n 0.0118298f $X=7.435 $Y=2.525 $X2=0
+ $Y2=0
cc_718 N_A_1309_65#_c_1034_n N_VPWR_c_1333_n 0.0184263f $X=8.735 $Y=3.15 $X2=0
+ $Y2=0
cc_719 N_A_1309_65#_c_1034_n N_VPWR_c_1334_n 0.0179038f $X=8.735 $Y=3.15 $X2=0
+ $Y2=0
cc_720 N_A_1309_65#_c_1034_n N_VPWR_c_1335_n 0.017719f $X=8.735 $Y=3.15 $X2=0
+ $Y2=0
cc_721 N_A_1309_65#_c_1027_n N_VPWR_c_1335_n 0.0934478f $X=8.88 $Y=1.835 $X2=0
+ $Y2=0
cc_722 N_A_1309_65#_c_1038_n N_VPWR_c_1335_n 0.0143825f $X=8.9 $Y=2.6 $X2=0
+ $Y2=0
cc_723 N_A_1309_65#_c_1027_n N_VPWR_c_1336_n 0.0119031f $X=8.88 $Y=1.835 $X2=0
+ $Y2=0
cc_724 N_A_1309_65#_c_1038_n N_VPWR_c_1336_n 0.00730807f $X=8.9 $Y=2.6 $X2=0
+ $Y2=0
cc_725 N_A_1309_65#_c_1032_n N_VPWR_c_1343_n 0.0206019f $X=7.02 $Y=3.15 $X2=0
+ $Y2=0
cc_726 N_A_1309_65#_c_1034_n N_VPWR_c_1347_n 0.0141962f $X=8.735 $Y=3.15 $X2=0
+ $Y2=0
cc_727 N_A_1309_65#_c_1027_n N_VPWR_c_1347_n 0.0223605f $X=8.88 $Y=1.835 $X2=0
+ $Y2=0
cc_728 N_A_1309_65#_c_1031_n N_VPWR_c_1327_n 0.00943716f $X=7.36 $Y=3.15 $X2=0
+ $Y2=0
cc_729 N_A_1309_65#_c_1032_n N_VPWR_c_1327_n 0.00559553f $X=7.02 $Y=3.15 $X2=0
+ $Y2=0
cc_730 N_A_1309_65#_c_1034_n N_VPWR_c_1327_n 0.0440439f $X=8.735 $Y=3.15 $X2=0
+ $Y2=0
cc_731 N_A_1309_65#_c_1036_n N_VPWR_c_1327_n 0.00829772f $X=7.435 $Y=3.15 $X2=0
+ $Y2=0
cc_732 N_A_1309_65#_c_1027_n N_VPWR_c_1327_n 0.0112511f $X=8.88 $Y=1.835 $X2=0
+ $Y2=0
cc_733 N_A_1309_65#_c_1030_n N_A_988_379#_c_1513_n 0.00681689f $X=6.945 $Y=3.075
+ $X2=0 $Y2=0
cc_734 N_A_1309_65#_c_1030_n N_A_1095_425#_c_1540_n 0.00226483f $X=6.945
+ $Y=3.075 $X2=0 $Y2=0
cc_735 N_A_1309_65#_c_1031_n N_A_1095_425#_c_1540_n 0.00287373f $X=7.36 $Y=3.15
+ $X2=0 $Y2=0
cc_736 N_A_1309_65#_M1008_g N_A_1095_425#_c_1540_n 0.00339238f $X=7.435 $Y=2.525
+ $X2=0 $Y2=0
cc_737 N_A_1309_65#_c_1030_n N_A_1095_425#_c_1541_n 0.0134316f $X=6.945 $Y=3.075
+ $X2=0 $Y2=0
cc_738 N_A_1309_65#_c_1035_n N_A_1095_425#_c_1541_n 0.0028635f $X=6.945 $Y=2.23
+ $X2=0 $Y2=0
cc_739 N_A_1309_65#_M1001_g N_VGND_c_1583_n 0.00170531f $X=6.62 $Y=0.665 $X2=0
+ $Y2=0
cc_740 N_A_1309_65#_c_1028_n N_VGND_c_1583_n 0.0126699f $X=7.955 $Y=0.57 $X2=0
+ $Y2=0
cc_741 N_A_1309_65#_M1001_g N_VGND_c_1590_n 0.00517164f $X=6.62 $Y=0.665 $X2=0
+ $Y2=0
cc_742 N_A_1309_65#_c_1026_n N_VGND_c_1595_n 0.010631f $X=8.735 $Y=0.53 $X2=0
+ $Y2=0
cc_743 N_A_1309_65#_c_1028_n N_VGND_c_1595_n 0.0318702f $X=7.955 $Y=0.57 $X2=0
+ $Y2=0
cc_744 N_A_1309_65#_M1001_g N_VGND_c_1601_n 0.00519032f $X=6.62 $Y=0.665 $X2=0
+ $Y2=0
cc_745 N_A_1309_65#_c_1026_n N_VGND_c_1601_n 0.0114673f $X=8.735 $Y=0.53 $X2=0
+ $Y2=0
cc_746 N_A_1309_65#_c_1028_n N_VGND_c_1601_n 0.0324821f $X=7.955 $Y=0.57 $X2=0
+ $Y2=0
cc_747 N_A_1158_47#_c_1137_n N_A_1855_47#_M1012_g 0.0195057f $X=9.54 $Y=1.8
+ $X2=0 $Y2=0
cc_748 N_A_1158_47#_c_1118_n N_A_1855_47#_c_1264_n 0.00495346f $X=8.285 $Y=0.27
+ $X2=0 $Y2=0
cc_749 N_A_1158_47#_c_1121_n N_A_1855_47#_c_1264_n 0.00355357f $X=9.155 $Y=1.315
+ $X2=0 $Y2=0
cc_750 N_A_1158_47#_c_1123_n N_A_1855_47#_c_1264_n 0.0199166f $X=9.54 $Y=0.87
+ $X2=0 $Y2=0
cc_751 N_A_1158_47#_M1018_g N_A_1855_47#_c_1264_n 0.00415083f $X=9.615 $Y=0.445
+ $X2=0 $Y2=0
cc_752 N_A_1158_47#_c_1133_n N_A_1855_47#_c_1264_n 7.0734e-19 $X=8.45 $Y=0.96
+ $X2=0 $Y2=0
cc_753 N_A_1158_47#_M1004_g N_A_1855_47#_c_1265_n 9.15784e-19 $X=8.665 $Y=1.835
+ $X2=0 $Y2=0
cc_754 N_A_1158_47#_c_1122_n N_A_1855_47#_c_1265_n 0.00283872f $X=9.155 $Y=1.725
+ $X2=0 $Y2=0
cc_755 N_A_1158_47#_c_1137_n N_A_1855_47#_c_1265_n 0.0207299f $X=9.54 $Y=1.8
+ $X2=0 $Y2=0
cc_756 N_A_1158_47#_c_1139_n N_A_1855_47#_c_1265_n 0.00451162f $X=9.615 $Y=1.875
+ $X2=0 $Y2=0
cc_757 N_A_1158_47#_c_1123_n N_A_1855_47#_c_1266_n 0.00695185f $X=9.54 $Y=0.87
+ $X2=0 $Y2=0
cc_758 N_A_1158_47#_c_1137_n N_A_1855_47#_c_1266_n 0.00722699f $X=9.54 $Y=1.8
+ $X2=0 $Y2=0
cc_759 N_A_1158_47#_c_1121_n N_A_1855_47#_c_1267_n 0.00473669f $X=9.155 $Y=1.315
+ $X2=0 $Y2=0
cc_760 N_A_1158_47#_c_1137_n N_A_1855_47#_c_1267_n 3.93747e-19 $X=9.54 $Y=1.8
+ $X2=0 $Y2=0
cc_761 N_A_1158_47#_c_1121_n N_A_1855_47#_c_1268_n 0.00456568f $X=9.155 $Y=1.315
+ $X2=0 $Y2=0
cc_762 N_A_1158_47#_M1018_g N_A_1855_47#_c_1269_n 0.015838f $X=9.615 $Y=0.445
+ $X2=0 $Y2=0
cc_763 N_A_1158_47#_c_1142_n N_VPWR_c_1333_n 0.0160706f $X=7.955 $Y=2.18 $X2=0
+ $Y2=0
cc_764 N_A_1158_47#_c_1143_n N_VPWR_c_1334_n 0.00415128f $X=8.08 $Y=2.525 $X2=0
+ $Y2=0
cc_765 N_A_1158_47#_M1004_g N_VPWR_c_1335_n 0.00168517f $X=8.665 $Y=1.835 $X2=0
+ $Y2=0
cc_766 N_A_1158_47#_c_1126_n N_VPWR_c_1335_n 0.00128552f $X=8.512 $Y=1.39 $X2=0
+ $Y2=0
cc_767 N_A_1158_47#_c_1143_n N_VPWR_c_1335_n 0.0326859f $X=8.08 $Y=2.525 $X2=0
+ $Y2=0
cc_768 N_A_1158_47#_c_1131_n N_VPWR_c_1335_n 0.0126768f $X=8.085 $Y=1.465 $X2=0
+ $Y2=0
cc_769 N_A_1158_47#_c_1132_n N_VPWR_c_1335_n 0.0324848f $X=8.085 $Y=2.095 $X2=0
+ $Y2=0
cc_770 N_A_1158_47#_c_1148_n N_VPWR_c_1335_n 0.0145186f $X=8.075 $Y=2.18 $X2=0
+ $Y2=0
cc_771 N_A_1158_47#_c_1139_n N_VPWR_c_1336_n 0.00197417f $X=9.615 $Y=1.875 $X2=0
+ $Y2=0
cc_772 N_A_1158_47#_c_1139_n N_VPWR_c_1347_n 0.00375548f $X=9.615 $Y=1.875 $X2=0
+ $Y2=0
cc_773 N_A_1158_47#_c_1139_n N_VPWR_c_1327_n 0.00447875f $X=9.615 $Y=1.875 $X2=0
+ $Y2=0
cc_774 N_A_1158_47#_c_1143_n N_VPWR_c_1327_n 0.00625693f $X=8.08 $Y=2.525 $X2=0
+ $Y2=0
cc_775 N_A_1158_47#_c_1142_n N_A_988_379#_M1026_d 0.00244268f $X=7.955 $Y=2.18
+ $X2=0 $Y2=0
cc_776 N_A_1158_47#_M1014_d N_A_988_379#_c_1513_n 0.00307529f $X=5.89 $Y=2.125
+ $X2=0 $Y2=0
cc_777 N_A_1158_47#_c_1142_n N_A_1095_425#_c_1540_n 0.0227936f $X=7.955 $Y=2.18
+ $X2=0 $Y2=0
cc_778 N_A_1158_47#_M1014_d N_A_1095_425#_c_1541_n 0.00531861f $X=5.89 $Y=2.125
+ $X2=0 $Y2=0
cc_779 N_A_1158_47#_c_1142_n N_A_1095_425#_c_1541_n 0.0342763f $X=7.955 $Y=2.18
+ $X2=0 $Y2=0
cc_780 N_A_1158_47#_c_1146_n N_A_1095_425#_c_1541_n 0.0254553f $X=6.255 $Y=2.22
+ $X2=0 $Y2=0
cc_781 N_A_1158_47#_c_1129_n N_VGND_M1013_d 0.00525719f $X=7.975 $Y=0.95 $X2=0
+ $Y2=0
cc_782 N_A_1158_47#_c_1119_n N_VGND_c_1583_n 0.0107868f $X=7.63 $Y=0.27 $X2=0
+ $Y2=0
cc_783 N_A_1158_47#_c_1129_n N_VGND_c_1583_n 0.01937f $X=7.975 $Y=0.95 $X2=0
+ $Y2=0
cc_784 N_A_1158_47#_M1018_g N_VGND_c_1584_n 0.00601949f $X=9.615 $Y=0.445 $X2=0
+ $Y2=0
cc_785 N_A_1158_47#_M1018_g N_VGND_c_1585_n 0.00343843f $X=9.615 $Y=0.445 $X2=0
+ $Y2=0
cc_786 N_A_1158_47#_c_1128_n N_VGND_c_1590_n 0.0210895f $X=5.95 $Y=0.39 $X2=0
+ $Y2=0
cc_787 N_A_1158_47#_M1018_g N_VGND_c_1681_n 0.00171458f $X=9.615 $Y=0.445 $X2=0
+ $Y2=0
cc_788 N_A_1158_47#_c_1119_n N_VGND_c_1595_n 0.0251559f $X=7.63 $Y=0.27 $X2=0
+ $Y2=0
cc_789 N_A_1158_47#_M1018_g N_VGND_c_1595_n 0.00564095f $X=9.615 $Y=0.445 $X2=0
+ $Y2=0
cc_790 N_A_1158_47#_M1030_d N_VGND_c_1601_n 0.00231914f $X=5.79 $Y=0.235 $X2=0
+ $Y2=0
cc_791 N_A_1158_47#_c_1118_n N_VGND_c_1601_n 0.0258528f $X=8.285 $Y=0.27 $X2=0
+ $Y2=0
cc_792 N_A_1158_47#_c_1119_n N_VGND_c_1601_n 0.00994933f $X=7.63 $Y=0.27 $X2=0
+ $Y2=0
cc_793 N_A_1158_47#_c_1124_n N_VGND_c_1601_n 0.00457926f $X=9.23 $Y=0.87 $X2=0
+ $Y2=0
cc_794 N_A_1158_47#_M1018_g N_VGND_c_1601_n 0.0107826f $X=9.615 $Y=0.445 $X2=0
+ $Y2=0
cc_795 N_A_1158_47#_c_1128_n N_VGND_c_1601_n 0.0126604f $X=5.95 $Y=0.39 $X2=0
+ $Y2=0
cc_796 N_A_1158_47#_c_1129_n A_1267_91# 0.00366293f $X=7.975 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_797 N_A_1158_47#_c_1129_n A_1339_91# 0.00366293f $X=7.975 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_798 N_A_1855_47#_M1012_g N_VPWR_c_1336_n 0.0185472f $X=10.125 $Y=2.465 $X2=0
+ $Y2=0
cc_799 N_A_1855_47#_c_1265_n N_VPWR_c_1336_n 0.0011898f $X=9.4 $Y=2.13 $X2=0
+ $Y2=0
cc_800 N_A_1855_47#_c_1266_n N_VPWR_c_1336_n 0.00842408f $X=9.97 $Y=1.35 $X2=0
+ $Y2=0
cc_801 N_A_1855_47#_c_1268_n N_VPWR_c_1336_n 0.00249114f $X=10.002 $Y=1.26 $X2=0
+ $Y2=0
cc_802 N_A_1855_47#_M1022_g N_VPWR_c_1338_n 0.00929098f $X=10.555 $Y=2.465 $X2=0
+ $Y2=0
cc_803 N_A_1855_47#_c_1265_n N_VPWR_c_1347_n 0.0048157f $X=9.4 $Y=2.13 $X2=0
+ $Y2=0
cc_804 N_A_1855_47#_M1012_g N_VPWR_c_1348_n 0.00585385f $X=10.125 $Y=2.465 $X2=0
+ $Y2=0
cc_805 N_A_1855_47#_M1022_g N_VPWR_c_1348_n 0.00585385f $X=10.555 $Y=2.465 $X2=0
+ $Y2=0
cc_806 N_A_1855_47#_M1012_g N_VPWR_c_1327_n 0.0122727f $X=10.125 $Y=2.465 $X2=0
+ $Y2=0
cc_807 N_A_1855_47#_M1022_g N_VPWR_c_1327_n 0.0114507f $X=10.555 $Y=2.465 $X2=0
+ $Y2=0
cc_808 N_A_1855_47#_c_1265_n N_VPWR_c_1327_n 0.00777987f $X=9.4 $Y=2.13 $X2=0
+ $Y2=0
cc_809 N_A_1855_47#_c_1260_n N_Q_c_1563_n 0.0162686f $X=10.48 $Y=1.26 $X2=0
+ $Y2=0
cc_810 N_A_1855_47#_c_1261_n N_Q_c_1563_n 0.00311209f $X=10.555 $Y=1.185 $X2=0
+ $Y2=0
cc_811 N_A_1855_47#_M1022_g N_Q_c_1563_n 0.0135487f $X=10.555 $Y=2.465 $X2=0
+ $Y2=0
cc_812 N_A_1855_47#_c_1266_n N_Q_c_1563_n 0.0262928f $X=9.97 $Y=1.35 $X2=0 $Y2=0
cc_813 N_A_1855_47#_c_1268_n N_Q_c_1563_n 0.010561f $X=10.002 $Y=1.26 $X2=0
+ $Y2=0
cc_814 N_A_1855_47#_c_1269_n N_Q_c_1563_n 0.00342387f $X=10.002 $Y=1.185 $X2=0
+ $Y2=0
cc_815 N_A_1855_47#_c_1261_n N_VGND_c_1584_n 6.5348e-19 $X=10.555 $Y=1.185 $X2=0
+ $Y2=0
cc_816 N_A_1855_47#_c_1269_n N_VGND_c_1584_n 0.00643439f $X=10.002 $Y=1.185
+ $X2=0 $Y2=0
cc_817 N_A_1855_47#_c_1264_n N_VGND_c_1585_n 0.0231505f $X=9.4 $Y=0.42 $X2=0
+ $Y2=0
cc_818 N_A_1855_47#_c_1266_n N_VGND_c_1585_n 0.0230997f $X=9.97 $Y=1.35 $X2=0
+ $Y2=0
cc_819 N_A_1855_47#_c_1268_n N_VGND_c_1585_n 0.00553375f $X=10.002 $Y=1.26 $X2=0
+ $Y2=0
cc_820 N_A_1855_47#_c_1269_n N_VGND_c_1585_n 0.00543223f $X=10.002 $Y=1.185
+ $X2=0 $Y2=0
cc_821 N_A_1855_47#_c_1261_n N_VGND_c_1587_n 0.00715777f $X=10.555 $Y=1.185
+ $X2=0 $Y2=0
cc_822 N_A_1855_47#_c_1266_n N_VGND_c_1681_n 0.00101671f $X=9.97 $Y=1.35 $X2=0
+ $Y2=0
cc_823 N_A_1855_47#_c_1269_n N_VGND_c_1681_n 0.00426092f $X=10.002 $Y=1.185
+ $X2=0 $Y2=0
cc_824 N_A_1855_47#_c_1264_n N_VGND_c_1595_n 0.0185207f $X=9.4 $Y=0.42 $X2=0
+ $Y2=0
cc_825 N_A_1855_47#_c_1261_n N_VGND_c_1596_n 0.00585385f $X=10.555 $Y=1.185
+ $X2=0 $Y2=0
cc_826 N_A_1855_47#_c_1269_n N_VGND_c_1596_n 0.00564095f $X=10.002 $Y=1.185
+ $X2=0 $Y2=0
cc_827 N_A_1855_47#_M1018_s N_VGND_c_1601_n 0.00245057f $X=9.275 $Y=0.235 $X2=0
+ $Y2=0
cc_828 N_A_1855_47#_c_1261_n N_VGND_c_1601_n 0.0114507f $X=10.555 $Y=1.185 $X2=0
+ $Y2=0
cc_829 N_A_1855_47#_c_1264_n N_VGND_c_1601_n 0.010808f $X=9.4 $Y=0.42 $X2=0
+ $Y2=0
cc_830 N_A_1855_47#_c_1269_n N_VGND_c_1601_n 0.00948291f $X=10.002 $Y=1.185
+ $X2=0 $Y2=0
cc_831 N_VPWR_c_1341_n N_A_400_119#_c_1468_n 0.00327175f $X=3.195 $Y=3.33 $X2=0
+ $Y2=0
cc_832 N_VPWR_c_1327_n N_A_400_119#_c_1468_n 0.00482454f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_833 N_VPWR_c_1327_n N_A_988_379#_M1026_d 0.00204235f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_834 N_VPWR_c_1332_n N_A_988_379#_c_1511_n 0.0130458f $X=4.455 $Y=3.245 $X2=0
+ $Y2=0
cc_835 N_VPWR_c_1332_n N_A_988_379#_c_1512_n 0.0183902f $X=4.455 $Y=3.245 $X2=0
+ $Y2=0
cc_836 N_VPWR_c_1343_n N_A_988_379#_c_1512_n 0.0209882f $X=7.555 $Y=3.33 $X2=0
+ $Y2=0
cc_837 N_VPWR_c_1327_n N_A_988_379#_c_1512_n 0.0113884f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_838 N_VPWR_c_1343_n N_A_988_379#_c_1513_n 0.0913304f $X=7.555 $Y=3.33 $X2=0
+ $Y2=0
cc_839 N_VPWR_c_1327_n N_A_988_379#_c_1513_n 0.0544045f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_840 N_VPWR_c_1343_n N_A_1095_425#_c_1541_n 0.00895986f $X=7.555 $Y=3.33 $X2=0
+ $Y2=0
cc_841 N_VPWR_c_1327_n N_A_1095_425#_c_1541_n 0.0155888f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_842 N_VPWR_c_1327_n N_Q_M1012_d 0.00362709f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_843 N_VPWR_c_1338_n N_Q_c_1563_n 0.00153242f $X=10.77 $Y=1.98 $X2=0 $Y2=0
cc_844 N_VPWR_c_1348_n N_Q_c_1563_n 0.0142265f $X=10.635 $Y=3.33 $X2=0 $Y2=0
cc_845 N_VPWR_c_1327_n N_Q_c_1563_n 0.00925289f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_846 N_A_400_119#_c_1502_n N_VGND_c_1588_n 0.00357861f $X=2.14 $Y=0.805 $X2=0
+ $Y2=0
cc_847 N_A_400_119#_c_1502_n N_VGND_c_1601_n 0.00567908f $X=2.14 $Y=0.805 $X2=0
+ $Y2=0
cc_848 N_A_988_379#_c_1511_n N_A_1095_425#_c_1538_n 0.0261668f $X=5.08 $Y=2.19
+ $X2=0 $Y2=0
cc_849 N_A_988_379#_c_1511_n N_A_1095_425#_c_1539_n 0.0139f $X=5.08 $Y=2.19
+ $X2=0 $Y2=0
cc_850 N_A_988_379#_c_1513_n N_A_1095_425#_c_1539_n 0.0217425f $X=6.67 $Y=2.95
+ $X2=0 $Y2=0
cc_851 N_A_988_379#_M1026_d N_A_1095_425#_c_1541_n 0.00754474f $X=6.435 $Y=2.125
+ $X2=0 $Y2=0
cc_852 N_A_988_379#_c_1513_n N_A_1095_425#_c_1541_n 0.0707721f $X=6.67 $Y=2.95
+ $X2=0 $Y2=0
cc_853 N_Q_c_1563_n N_VGND_c_1587_n 0.00153242f $X=10.34 $Y=0.42 $X2=0 $Y2=0
cc_854 N_Q_c_1563_n N_VGND_c_1596_n 0.0142265f $X=10.34 $Y=0.42 $X2=0 $Y2=0
cc_855 N_Q_M1016_d N_VGND_c_1601_n 0.00362709f $X=10.2 $Y=0.235 $X2=0 $Y2=0
cc_856 N_Q_c_1563_n N_VGND_c_1601_n 0.00925289f $X=10.34 $Y=0.42 $X2=0 $Y2=0
cc_857 N_VGND_c_1601_n A_857_47# 0.00899413f $X=10.8 $Y=0 $X2=-0.19 $Y2=-0.245
cc_858 N_VGND_c_1601_n A_1086_47# 0.00899413f $X=10.8 $Y=0 $X2=-0.19 $Y2=-0.245
