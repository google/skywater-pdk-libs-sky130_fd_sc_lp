* File: sky130_fd_sc_lp__a311o_1.pex.spice
* Created: Wed Sep  2 09:25:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311O_1%A_80_21# 1 2 3 10 12 15 20 23 24 25 26 27 30
+ 32 36 40 44 45 49
r106 40 42 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=3.545 $Y=1.98
+ $X2=3.545 $Y2=2.95
r107 38 40 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.545 $Y=1.865
+ $X2=3.545 $Y2=1.98
r108 34 36 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.545 $Y=0.855
+ $X2=3.545 $Y2=0.38
r109 33 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0.94
+ $X2=2.49 $Y2=0.94
r110 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.38 $Y=0.94
+ $X2=3.545 $Y2=0.855
r111 32 33 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.38 $Y=0.94
+ $X2=2.655 $Y2=0.94
r112 28 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.855
+ $X2=2.49 $Y2=0.94
r113 28 30 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.49 $Y=0.855
+ $X2=2.49 $Y2=0.42
r114 26 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.38 $Y=1.78
+ $X2=3.545 $Y2=1.865
r115 26 27 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=3.38 $Y=1.78
+ $X2=0.84 $Y2=1.78
r116 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0.94
+ $X2=2.49 $Y2=0.94
r117 24 25 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=2.325 $Y=0.94
+ $X2=0.84 $Y2=0.94
r118 23 27 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.722 $Y=1.695
+ $X2=0.84 $Y2=1.78
r119 23 44 8.82722 $w=2.33e-07 $l=1.8e-07 $layer=LI1_cond $X=0.722 $Y=1.695
+ $X2=0.722 $Y2=1.515
r120 21 49 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.61 $Y=1.35
+ $X2=0.72 $Y2=1.35
r121 21 46 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.61 $Y=1.35
+ $X2=0.475 $Y2=1.35
r122 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.35 $X2=0.61 $Y2=1.35
r123 18 44 6.51225 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=0.682 $Y=1.358
+ $X2=0.682 $Y2=1.515
r124 18 20 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=0.682 $Y=1.358
+ $X2=0.682 $Y2=1.35
r125 17 25 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=0.682 $Y=1.025
+ $X2=0.84 $Y2=0.94
r126 17 20 11.8903 $w=3.13e-07 $l=3.25e-07 $layer=LI1_cond $X=0.682 $Y=1.025
+ $X2=0.682 $Y2=1.35
r127 13 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.515
+ $X2=0.72 $Y2=1.35
r128 13 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.72 $Y=1.515
+ $X2=0.72 $Y2=2.465
r129 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=1.35
r130 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
r131 3 42 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.835 $X2=3.545 $Y2=2.95
r132 3 40 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.835 $X2=3.545 $Y2=1.98
r133 2 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.235 $X2=3.545 $Y2=0.38
r134 1 30 91 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.235 $X2=2.49 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%A3 3 7 8 11 13
r36 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.36 $X2=1.2
+ $Y2=1.525
r37 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.36 $X2=1.2
+ $Y2=1.195
r38 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2 $Y=1.36
+ $X2=1.2 $Y2=1.36
r39 7 13 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.29 $Y=0.655 $X2=1.29
+ $Y2=1.195
r40 3 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.22 $Y=2.465 $X2=1.22
+ $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%A2 3 5 7 8 11
c32 3 0 2.14203e-20 $X=1.65 $Y=2.465
r33 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.35
+ $X2=1.74 $Y2=1.515
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.35 $X2=1.74 $Y2=1.35
r35 5 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.185
+ $X2=1.74 $Y2=1.35
r36 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.74 $Y=1.185 $X2=1.74
+ $Y2=0.655
r37 3 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.65 $Y=2.465
+ $X2=1.65 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%A1 1 3 6 8 14 15
c32 14 0 2.68576e-20 $X=2.28 $Y=1.36
r33 13 15 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.28 $Y=1.36
+ $X2=2.43 $Y2=1.36
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.36 $X2=2.28 $Y2=1.36
r35 10 13 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.19 $Y=1.36 $X2=2.28
+ $Y2=1.36
r36 8 14 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.16 $Y=1.36 $X2=2.28
+ $Y2=1.36
r37 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.525
+ $X2=2.43 $Y2=1.36
r38 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.43 $Y=1.525 $X2=2.43
+ $Y2=2.465
r39 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.195
+ $X2=2.19 $Y2=1.36
r40 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.19 $Y=1.195 $X2=2.19
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%B1 3 6 8 9 13 15
c33 6 0 5.43728e-21 $X=2.97 $Y=2.465
r34 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.35
+ $X2=2.88 $Y2=1.515
r35 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.35
+ $X2=2.88 $Y2=1.185
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.35 $X2=2.88 $Y2=1.35
r37 9 14 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.36 $X2=2.88
+ $Y2=1.36
r38 8 14 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.64 $Y=1.36 $X2=2.88
+ $Y2=1.36
r39 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.97 $Y=2.465
+ $X2=2.97 $Y2=1.515
r40 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.79 $Y=0.655
+ $X2=2.79 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%C1 1 3 6 8 13
r24 10 13 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.33 $Y=1.36
+ $X2=3.57 $Y2=1.36
r25 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.36 $X2=3.57 $Y2=1.36
r26 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.525
+ $X2=3.33 $Y2=1.36
r27 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.33 $Y=1.525 $X2=3.33
+ $Y2=2.465
r28 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.195
+ $X2=3.33 $Y2=1.36
r29 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.33 $Y=1.195 $X2=3.33
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%X 1 2 7 8 9 10 11 12 13 25 37 40
r20 38 40 1.59477 $w=5.83e-07 $l=7.8e-08 $layer=LI1_cond $X=0.377 $Y=2.327
+ $X2=0.377 $Y2=2.405
r21 13 45 2.76018 $w=5.83e-07 $l=1.35e-07 $layer=LI1_cond $X=0.377 $Y=2.775
+ $X2=0.377 $Y2=2.91
r22 12 38 0.0817831 $w=5.83e-07 $l=4e-09 $layer=LI1_cond $X=0.377 $Y=2.323
+ $X2=0.377 $Y2=2.327
r23 12 52 4.15049 $w=5.83e-07 $l=2.03e-07 $layer=LI1_cond $X=0.377 $Y=2.323
+ $X2=0.377 $Y2=2.12
r24 12 13 7.5036 $w=5.83e-07 $l=3.67e-07 $layer=LI1_cond $X=0.377 $Y=2.408
+ $X2=0.377 $Y2=2.775
r25 12 40 0.0613374 $w=5.83e-07 $l=3e-09 $layer=LI1_cond $X=0.377 $Y=2.408
+ $X2=0.377 $Y2=2.405
r26 11 52 0.879169 $w=5.83e-07 $l=4.3e-08 $layer=LI1_cond $X=0.377 $Y=2.077
+ $X2=0.377 $Y2=2.12
r27 11 37 0.858723 $w=5.83e-07 $l=4.2e-08 $layer=LI1_cond $X=0.377 $Y=2.077
+ $X2=0.377 $Y2=2.035
r28 11 37 1.83537 $w=2.68e-07 $l=4.3e-08 $layer=LI1_cond $X=0.22 $Y=1.992
+ $X2=0.22 $Y2=2.035
r29 10 11 13.9574 $w=2.68e-07 $l=3.27e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=1.992
r30 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.665
r31 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.925 $X2=0.22
+ $Y2=1.295
r32 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.555 $X2=0.22
+ $Y2=0.925
r33 7 25 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=0.555
+ $X2=0.22 $Y2=0.42
r34 2 52 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=1.835 $X2=0.505 $Y2=2.12
r35 2 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=1.835 $X2=0.505 $Y2=2.91
r36 1 25 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%VPWR 1 2 9 15 18 19 20 26 35 36 39
r45 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 30 39 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=2.38 $Y=3.33 $X2=2.04
+ $Y2=3.33
r52 30 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 26 39 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=1.7 $Y=3.33 $X2=2.04
+ $Y2=3.33
r55 26 28 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.7 $Y=3.33 $X2=1.68
+ $Y2=3.33
r56 24 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 20 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 20 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 18 23 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 18 19 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.84 $Y=3.33 $X2=0.97
+ $Y2=3.33
r62 17 28 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.68
+ $Y2=3.33
r63 17 19 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=0.97
+ $Y2=3.33
r64 13 39 2.80049 $w=6.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=3.245
+ $X2=2.04 $Y2=3.33
r65 13 15 13.4559 $w=6.78e-07 $l=7.65e-07 $layer=LI1_cond $X=2.04 $Y=3.245
+ $X2=2.04 $Y2=2.48
r66 9 12 33.2435 $w=2.58e-07 $l=7.5e-07 $layer=LI1_cond $X=0.97 $Y=2.2 $X2=0.97
+ $Y2=2.95
r67 7 19 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=3.245
+ $X2=0.97 $Y2=3.33
r68 7 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.97 $Y=3.245
+ $X2=0.97 $Y2=2.95
r69 2 15 150 $w=1.7e-07 $l=8.55614e-07 $layer=licon1_PDIFF $count=4 $X=1.725
+ $Y=1.835 $X2=2.215 $Y2=2.48
r70 1 12 400 $w=1.7e-07 $l=1.20163e-06 $layer=licon1_PDIFF $count=1 $X=0.795
+ $Y=1.835 $X2=0.975 $Y2=2.95
r71 1 9 400 $w=1.7e-07 $l=4.4601e-07 $layer=licon1_PDIFF $count=1 $X=0.795
+ $Y=1.835 $X2=0.975 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%A_259_367# 1 2 7 9 11 13 15
r17 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=2.205
+ $X2=2.715 $Y2=2.12
r18 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.715 $Y=2.205
+ $X2=2.715 $Y2=2.56
r19 12 18 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.53 $Y=2.12 $X2=1.4
+ $Y2=2.12
r20 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=2.12
+ $X2=2.715 $Y2=2.12
r21 11 12 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.55 $Y=2.12
+ $X2=1.53 $Y2=2.12
r22 7 18 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=2.205 $X2=1.4
+ $Y2=2.12
r23 7 9 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=1.4 $Y=2.205 $X2=1.4
+ $Y2=2.525
r24 2 20 600 $w=1.7e-07 $l=3.756e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.835 $X2=2.715 $Y2=2.12
r25 2 15 300 $w=1.7e-07 $l=8.23332e-07 $layer=licon1_PDIFF $count=2 $X=2.505
+ $Y=1.835 $X2=2.715 $Y2=2.56
r26 1 18 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=1.295
+ $Y=1.835 $X2=1.435 $Y2=2.12
r27 1 9 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.295
+ $Y=1.835 $X2=1.435 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_1%VGND 1 2 9 11 13 18 25 26 38
r44 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 31 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r46 26 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r47 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r48 23 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.045
+ $Y2=0
r49 23 25 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.6
+ $Y2=0
r50 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r51 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r52 19 21 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.24 $Y=0 $X2=2.64
+ $Y2=0
r53 18 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.045
+ $Y2=0
r54 18 21 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r55 16 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 13 35 9.2006 $w=7.13e-07 $l=5.5e-07 $layer=LI1_cond $X=0.882 $Y=0 $X2=0.882
+ $Y2=0.55
r58 13 19 9.46138 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=0.882 $Y=0 $X2=1.24
+ $Y2=0
r59 13 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r60 13 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r62 11 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r63 11 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r64 7 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=0.085
+ $X2=3.045 $Y2=0
r65 7 9 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.045 $Y=0.085
+ $X2=3.045 $Y2=0.56
r66 2 9 182 $w=1.7e-07 $l=4.05123e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3.045 $Y2=0.56
r67 1 35 91 $w=1.7e-07 $l=6.64078e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=1.075 $Y2=0.55
.ends

