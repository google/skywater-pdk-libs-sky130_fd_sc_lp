* File: sky130_fd_sc_lp__a32oi_2.pex.spice
* Created: Fri Aug 28 10:01:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32OI_2%B2 1 3 6 8 10 13 17 20 21 30
c48 8 0 1.03418e-19 $X=0.985 $Y=1.275
r49 25 28 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.4 $Y=1.44
+ $X2=0.555 $Y2=1.44
r50 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.4
+ $Y=1.44 $X2=0.4 $Y2=1.44
r51 21 26 8.55291 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=0.285 $Y=1.665
+ $X2=0.285 $Y2=1.4
r52 20 26 3.38889 $w=3.78e-07 $l=1.05e-07 $layer=LI1_cond $X=0.285 $Y=1.295
+ $X2=0.285 $Y2=1.4
r53 18 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.895 $Y=1.44
+ $X2=0.985 $Y2=1.44
r54 18 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.895 $Y=1.44
+ $X2=0.555 $Y2=1.44
r55 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=1.44 $X2=0.895 $Y2=1.44
r56 15 26 3.157 $w=2.5e-07 $l=2e-07 $layer=LI1_cond $X=0.485 $Y=1.4 $X2=0.285
+ $Y2=1.4
r57 15 17 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.485 $Y=1.4
+ $X2=0.895 $Y2=1.4
r58 11 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.605
+ $X2=0.985 $Y2=1.44
r59 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.985 $Y=1.605
+ $X2=0.985 $Y2=2.465
r60 8 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.275
+ $X2=0.985 $Y2=1.44
r61 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.985 $Y=1.275
+ $X2=0.985 $Y2=0.745
r62 4 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.605
+ $X2=0.555 $Y2=1.44
r63 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.555 $Y=1.605
+ $X2=0.555 $Y2=2.465
r64 1 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.275
+ $X2=0.555 $Y2=1.44
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.555 $Y=1.275
+ $X2=0.555 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%B1 3 7 13 17 19 20 23 25 26
c56 17 0 5.96051e-20 $X=1.845 $Y=2.465
r57 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.51 $X2=2.06 $Y2=1.51
r58 22 25 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.845 $Y=1.51
+ $X2=2.06 $Y2=1.51
r59 22 23 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.51
+ $X2=1.77 $Y2=1.51
r60 20 26 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.08 $Y=1.665
+ $X2=2.08 $Y2=1.51
r61 15 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.675
+ $X2=1.845 $Y2=1.51
r62 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.845 $Y=1.675
+ $X2=1.845 $Y2=2.465
r63 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.345
+ $X2=1.845 $Y2=1.51
r64 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.845 $Y=1.345
+ $X2=1.845 $Y2=0.745
r65 10 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.49 $Y=1.42
+ $X2=1.415 $Y2=1.42
r66 10 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.49 $Y=1.42
+ $X2=1.77 $Y2=1.42
r67 5 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.415 $Y=1.495
+ $X2=1.415 $Y2=1.42
r68 5 7 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.415 $Y=1.495
+ $X2=1.415 $Y2=2.465
r69 1 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.415 $Y=1.345
+ $X2=1.415 $Y2=1.42
r70 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.415 $Y=1.345 $X2=1.415
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%A1 3 7 11 15 17 23 25
c54 23 0 5.96051e-20 $X=2.6 $Y=1.51
c55 11 0 1.53238e-19 $X=3.385 $Y=0.745
r56 24 25 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.955 $Y=1.51
+ $X2=3.385 $Y2=1.51
r57 22 24 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.6 $Y=1.51
+ $X2=2.955 $Y2=1.51
r58 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.51 $X2=2.6 $Y2=1.51
r59 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.51 $Y=1.51 $X2=2.6
+ $Y2=1.51
r60 17 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.6 $Y=1.665
+ $X2=2.6 $Y2=1.51
r61 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.385 $Y=1.675
+ $X2=3.385 $Y2=1.51
r62 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.385 $Y=1.675
+ $X2=3.385 $Y2=2.465
r63 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.385 $Y=1.345
+ $X2=3.385 $Y2=1.51
r64 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.385 $Y=1.345 $X2=3.385
+ $Y2=0.745
r65 5 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.345
+ $X2=2.955 $Y2=1.51
r66 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.955 $Y=1.345 $X2=2.955
+ $Y2=0.745
r67 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.675
+ $X2=2.51 $Y2=1.51
r68 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.51 $Y=1.675 $X2=2.51
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%A2 3 7 11 15 17 18 19 30
c50 30 0 3.76971e-19 $X=4.695 $Y=1.51
c51 3 0 1.53238e-19 $X=3.815 $Y=0.745
r52 28 30 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.49 $Y=1.51
+ $X2=4.695 $Y2=1.51
r53 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.49
+ $Y=1.51 $X2=4.49 $Y2=1.51
r54 26 28 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=4.245 $Y=1.51
+ $X2=4.49 $Y2=1.51
r55 25 26 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.895 $Y=1.51
+ $X2=4.245 $Y2=1.51
r56 23 25 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.815 $Y=1.51
+ $X2=3.895 $Y2=1.51
r57 19 29 2.48218 $w=3.23e-07 $l=7e-08 $layer=LI1_cond $X=4.56 $Y=1.587 $X2=4.49
+ $Y2=1.587
r58 18 29 14.5385 $w=3.23e-07 $l=4.1e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.49 $Y2=1.587
r59 17 18 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.587
+ $X2=4.08 $Y2=1.587
r60 13 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=1.675
+ $X2=4.695 $Y2=1.51
r61 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.695 $Y=1.675
+ $X2=4.695 $Y2=2.465
r62 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.345
+ $X2=4.245 $Y2=1.51
r63 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.245 $Y=1.345 $X2=4.245
+ $Y2=0.745
r64 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.895 $Y=1.675
+ $X2=3.895 $Y2=1.51
r65 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.895 $Y=1.675
+ $X2=3.895 $Y2=2.465
r66 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.345
+ $X2=3.815 $Y2=1.51
r67 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.815 $Y=1.345 $X2=3.815
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%A3 3 5 7 10 12 14 15 23
r38 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.36 $X2=5.84 $Y2=1.36
r39 21 23 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.705 $Y=1.36
+ $X2=5.84 $Y2=1.36
r40 20 21 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.555 $Y=1.36
+ $X2=5.705 $Y2=1.36
r41 19 20 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=5.275 $Y=1.36
+ $X2=5.555 $Y2=1.36
r42 17 19 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.125 $Y=1.36
+ $X2=5.275 $Y2=1.36
r43 15 24 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=6 $Y=1.36 $X2=5.84
+ $Y2=1.36
r44 12 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.705 $Y=1.195
+ $X2=5.705 $Y2=1.36
r45 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.705 $Y=1.195
+ $X2=5.705 $Y2=0.665
r46 8 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.555 $Y=1.525
+ $X2=5.555 $Y2=1.36
r47 8 10 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=5.555 $Y=1.525 $X2=5.555
+ $Y2=2.465
r48 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=1.195
+ $X2=5.275 $Y2=1.36
r49 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.275 $Y=1.195
+ $X2=5.275 $Y2=0.665
r50 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.525
+ $X2=5.125 $Y2=1.36
r51 1 3 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=5.125 $Y=1.525 $X2=5.125
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%A_43_367# 1 2 3 4 5 6 19 21 23 27 31 33 34
+ 35 39 41 43 45 47 49 53 59
c71 41 0 1.94336e-19 $X=3.645 $Y=2.09
r72 67 68 1.64865 $w=1.85e-07 $l=2.5e-08 $layer=LI1_cond $X=4.91 $Y=1.98
+ $X2=4.91 $Y2=2.005
r73 65 67 9.23243 $w=1.85e-07 $l=1.4e-07 $layer=LI1_cond $X=4.91 $Y=1.84
+ $X2=4.91 $Y2=1.98
r74 53 55 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=5.805 $Y=1.98
+ $X2=5.805 $Y2=2.91
r75 51 53 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=5.805 $Y=1.925
+ $X2=5.805 $Y2=1.98
r76 50 65 1.22693 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.005 $Y=1.84
+ $X2=4.91 $Y2=1.84
r77 49 51 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.675 $Y=1.84
+ $X2=5.805 $Y2=1.925
r78 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.675 $Y=1.84
+ $X2=5.005 $Y2=1.84
r79 45 68 5.45789 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=2.09 $X2=4.91
+ $Y2=2.005
r80 45 47 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=4.91 $Y=2.09
+ $X2=4.91 $Y2=2.445
r81 44 64 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.775 $Y=2.005
+ $X2=3.645 $Y2=2.005
r82 43 68 1.22693 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.815 $Y=2.005
+ $X2=4.91 $Y2=2.005
r83 43 44 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.815 $Y=2.005
+ $X2=3.775 $Y2=2.005
r84 42 62 3.52026 $w=2.65e-07 $l=8.74643e-08 $layer=LI1_cond $X=3.645 $Y=2.29
+ $X2=3.64 $Y2=2.375
r85 41 64 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=2.09
+ $X2=3.645 $Y2=2.005
r86 41 42 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=3.645 $Y=2.09
+ $X2=3.645 $Y2=2.29
r87 37 62 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.46
+ $X2=3.64 $Y2=2.375
r88 37 39 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.64 $Y=2.46
+ $X2=3.64 $Y2=2.485
r89 36 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.375
+ $X2=2.18 $Y2=2.375
r90 35 62 2.98021 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.505 $Y=2.375
+ $X2=3.64 $Y2=2.375
r91 35 36 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.505 $Y=2.375
+ $X2=2.345 $Y2=2.375
r92 33 61 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.46 $X2=2.18
+ $Y2=2.375
r93 33 34 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.18 $Y=2.46
+ $X2=2.18 $Y2=2.905
r94 32 59 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.295 $Y=2.99 $X2=1.2
+ $Y2=2.99
r95 31 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=2.18 $Y2=2.905
r96 31 32 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=1.295 $Y2=2.99
r97 27 30 40.8612 $w=1.88e-07 $l=7e-07 $layer=LI1_cond $X=1.2 $Y=2.2 $X2=1.2
+ $Y2=2.9
r98 25 59 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.905 $X2=1.2
+ $Y2=2.99
r99 25 30 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=2.905 $X2=1.2
+ $Y2=2.9
r100 24 58 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.435 $Y=2.99
+ $X2=0.305 $Y2=2.99
r101 23 59 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.105 $Y=2.99
+ $X2=1.2 $Y2=2.99
r102 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=2.99
+ $X2=0.435 $Y2=2.99
r103 19 58 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=2.905
+ $X2=0.305 $Y2=2.99
r104 19 21 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.305 $Y=2.905
+ $X2=0.305 $Y2=2.095
r105 6 55 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.63
+ $Y=1.835 $X2=5.77 $Y2=2.91
r106 6 53 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.63
+ $Y=1.835 $X2=5.77 $Y2=1.98
r107 5 67 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.77
+ $Y=1.835 $X2=4.91 $Y2=1.98
r108 5 47 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=4.77
+ $Y=1.835 $X2=4.91 $Y2=2.445
r109 4 64 600 $w=1.7e-07 $l=3.27872e-07 $layer=licon1_PDIFF $count=1 $X=3.46
+ $Y=1.835 $X2=3.64 $Y2=2.085
r110 4 39 300 $w=1.7e-07 $l=7.34507e-07 $layer=licon1_PDIFF $count=2 $X=3.46
+ $Y=1.835 $X2=3.64 $Y2=2.485
r111 3 61 300 $w=1.7e-07 $l=6.87823e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.835 $X2=2.18 $Y2=2.405
r112 2 30 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=2.9
r113 2 27 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=2.2
r114 1 58 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.91
r115 1 21 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%Y 1 2 3 4 15 19 20 23 25 27 29 30 31 37 38
+ 39 40 48 53 55
c87 55 0 1.82635e-19 $X=3.12 $Y=1.295
c88 38 0 1.53238e-19 $X=3.035 $Y=1.21
c89 23 0 1.03418e-19 $X=1.63 $Y=0.69
r90 52 55 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=1.245 $X2=3.17
+ $Y2=1.295
r91 40 53 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=3.17 $Y=2.02 $X2=3.17
+ $Y2=1.92
r92 39 53 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.17 $Y=1.665
+ $X2=3.17 $Y2=1.92
r93 38 46 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=1.16 $X2=3.17
+ $Y2=1.075
r94 38 52 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=1.16 $X2=3.17
+ $Y2=1.245
r95 38 39 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=3.17 $Y=1.312
+ $X2=3.17 $Y2=1.665
r96 38 55 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=3.17 $Y=1.312
+ $X2=3.17 $Y2=1.295
r97 37 46 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.17 $Y=0.925
+ $X2=3.17 $Y2=1.075
r98 37 48 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.17 $Y=0.925
+ $X2=3.17 $Y2=0.69
r99 35 36 2.08904 $w=2.92e-07 $l=5e-08 $layer=LI1_cond $X=1.63 $Y=1.97 $X2=1.63
+ $Y2=2.02
r100 33 35 7.93836 $w=2.92e-07 $l=1.9e-07 $layer=LI1_cond $X=1.63 $Y=1.78
+ $X2=1.63 $Y2=1.97
r101 32 36 2.95306 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=2.02
+ $X2=1.63 $Y2=2.02
r102 31 40 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=2.02
+ $X2=3.17 $Y2=2.02
r103 31 32 67.1 $w=1.98e-07 $l=1.21e-06 $layer=LI1_cond $X=3.005 $Y=2.02
+ $X2=1.795 $Y2=2.02
r104 29 38 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=1.16
+ $X2=3.17 $Y2=1.16
r105 29 30 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.005 $Y=1.16
+ $X2=1.795 $Y2=1.16
r106 25 36 3.88869 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=1.63 $Y=2.12 $X2=1.63
+ $Y2=2.02
r107 25 27 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.31
r108 21 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.63 $Y=1.075
+ $X2=1.795 $Y2=1.16
r109 21 23 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.63 $Y=1.075
+ $X2=1.63 $Y2=0.69
r110 19 33 3.90229 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=1.78
+ $X2=1.63 $Y2=1.78
r111 19 20 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.465 $Y=1.78
+ $X2=0.935 $Y2=1.78
r112 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.77 $Y=1.97
+ $X2=0.77 $Y2=2.65
r113 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.77 $Y=1.865
+ $X2=0.935 $Y2=1.78
r114 13 15 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.77 $Y=1.865
+ $X2=0.77 $Y2=1.97
r115 4 35 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.835 $X2=1.63 $Y2=1.97
r116 4 27 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=1.49
+ $Y=1.835 $X2=1.63 $Y2=2.31
r117 3 17 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=2.65
r118 3 15 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=1.97
r119 2 48 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=3.03
+ $Y=0.325 $X2=3.17 $Y2=0.69
r120 1 23 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=1.49
+ $Y=0.325 $X2=1.63 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%VPWR 1 2 3 12 16 21 22 23 30 40 41 46 52 54
r75 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 51 52 11.3415 $w=7.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=3.022
+ $X2=3.335 $Y2=3.022
r77 48 51 0.761833 $w=7.83e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=3.022
+ $X2=3.17 $Y2=3.022
r78 44 48 7.3136 $w=7.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=3.022
+ $X2=3.12 $Y2=3.022
r79 44 46 10.0464 $w=7.83e-07 $l=8e-08 $layer=LI1_cond $X=2.64 $Y=3.022 $X2=2.56
+ $Y2=3.022
r80 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r82 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r83 38 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 35 54 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.295 $Y2=3.33
r86 35 37 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 34 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 33 52 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=3.335 $Y2=3.33
r89 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r90 30 54 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.295 $Y2=3.33
r91 30 33 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r92 28 45 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 27 46 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.56 $Y2=3.33
r94 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r96 23 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 23 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 21 37 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.175 $Y=3.33
+ $X2=5.04 $Y2=3.33
r99 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=3.33
+ $X2=5.34 $Y2=3.33
r100 20 40 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=6 $Y2=3.33
r101 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=5.34 $Y2=3.33
r102 16 19 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=5.34 $Y=2.18
+ $X2=5.34 $Y2=2.95
r103 14 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=3.245
+ $X2=5.34 $Y2=3.33
r104 14 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.34 $Y=3.245
+ $X2=5.34 $Y2=2.95
r105 10 54 2.86223 $w=7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=3.245
+ $X2=4.295 $Y2=3.33
r106 10 12 14.6947 $w=6.98e-07 $l=8.6e-07 $layer=LI1_cond $X=4.295 $Y=3.245
+ $X2=4.295 $Y2=2.385
r107 3 19 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.835 $X2=5.34 $Y2=2.95
r108 3 16 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.835 $X2=5.34 $Y2=2.18
r109 2 12 150 $w=1.7e-07 $l=7.63544e-07 $layer=licon1_PDIFF $count=4 $X=3.97
+ $Y=1.835 $X2=4.48 $Y2=2.385
r110 1 51 300 $w=1.7e-07 $l=1.18184e-06 $layer=licon1_PDIFF $count=2 $X=2.585
+ $Y=1.835 $X2=3.17 $Y2=2.76
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%A_43_65# 1 2 3 12 14 15 20 21 24
r35 22 24 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.13 $Y=0.435
+ $X2=2.13 $Y2=0.47
r36 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.965 $Y=0.35
+ $X2=2.13 $Y2=0.435
r37 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.965 $Y=0.35
+ $X2=1.295 $Y2=0.35
r38 17 19 23.3493 $w=1.88e-07 $l=4e-07 $layer=LI1_cond $X=1.2 $Y=0.87 $X2=1.2
+ $Y2=0.47
r39 16 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.2 $Y=0.435
+ $X2=1.295 $Y2=0.35
r40 16 19 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=1.2 $Y=0.435 $X2=1.2
+ $Y2=0.47
r41 14 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.105 $Y=0.955
+ $X2=1.2 $Y2=0.87
r42 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=0.955
+ $X2=0.435 $Y2=0.955
r43 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.305 $Y=0.87
+ $X2=0.435 $Y2=0.955
r44 10 12 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.305 $Y=0.87
+ $X2=0.305 $Y2=0.48
r45 3 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.92
+ $Y=0.325 $X2=2.13 $Y2=0.47
r46 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.325 $X2=1.2 $Y2=0.47
r47 1 12 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.325 $X2=0.34 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%VGND 1 2 3 12 16 18 20 22 24 29 37 43 46 50
r66 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r67 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r68 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r70 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r71 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r72 38 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.06
+ $Y2=0
r73 38 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.52
+ $Y2=0
r74 37 49 4.65202 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.997
+ $Y2=0
r75 37 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.52
+ $Y2=0
r76 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r77 35 36 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r78 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r79 32 35 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r80 32 33 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r81 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.77
+ $Y2=0
r82 30 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.2
+ $Y2=0
r83 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=0 $X2=5.06
+ $Y2=0
r84 29 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.56
+ $Y2=0
r85 27 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r86 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r87 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.77
+ $Y2=0
r88 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r89 22 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r90 22 33 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=1.2
+ $Y2=0
r91 18 49 3.11416 $w=3.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.997 $Y2=0
r92 18 20 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.39
r93 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0
r94 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0.39
r95 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0
r96 10 12 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0.575
r97 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.78
+ $Y=0.245 $X2=5.92 $Y2=0.39
r98 2 16 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.935
+ $Y=0.245 $X2=5.06 $Y2=0.39
r99 1 12 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.325 $X2=0.77 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%A_509_65# 1 2 3 12 14 15 18 20 24 26
r40 22 24 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=4.53 $Y=0.435
+ $X2=4.53 $Y2=0.47
r41 21 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.695 $Y=0.35 $X2=3.6
+ $Y2=0.35
r42 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.365 $Y=0.35
+ $X2=4.53 $Y2=0.435
r43 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.365 $Y=0.35
+ $X2=3.695 $Y2=0.35
r44 16 26 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.435 $X2=3.6
+ $Y2=0.35
r45 16 18 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.6 $Y=0.435 $X2=3.6
+ $Y2=0.47
r46 14 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.505 $Y=0.35 $X2=3.6
+ $Y2=0.35
r47 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.505 $Y=0.35
+ $X2=2.835 $Y2=0.35
r48 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.67 $Y=0.435
+ $X2=2.835 $Y2=0.35
r49 10 12 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.67 $Y=0.435
+ $X2=2.67 $Y2=0.47
r50 3 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.32
+ $Y=0.325 $X2=4.53 $Y2=0.47
r51 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.46
+ $Y=0.325 $X2=3.6 $Y2=0.47
r52 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.545
+ $Y=0.325 $X2=2.67 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_2%A_778_65# 1 2 9 11 12 15
c30 12 0 1.53238e-19 $X=4.195 $Y=1.16
r31 13 15 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=5.49 $Y=1.075
+ $X2=5.49 $Y2=0.42
r32 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.395 $Y=1.16
+ $X2=5.49 $Y2=1.075
r33 11 12 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=5.395 $Y=1.16
+ $X2=4.195 $Y2=1.16
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.03 $Y=1.075
+ $X2=4.195 $Y2=1.16
r35 7 9 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.03 $Y=1.075
+ $X2=4.03 $Y2=0.69
r36 2 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=5.35
+ $Y=0.245 $X2=5.49 $Y2=0.42
r37 1 9 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=3.89
+ $Y=0.325 $X2=4.03 $Y2=0.69
.ends

