* File: sky130_fd_sc_lp__or3b_1.pxi.spice
* Created: Fri Aug 28 11:23:55 2020
* 
x_PM_SKY130_FD_SC_LP__OR3B_1%C_N N_C_N_c_68_n N_C_N_M1003_g N_C_N_M1006_g
+ N_C_N_c_70_n C_N C_N C_N C_N C_N N_C_N_c_72_n N_C_N_c_73_n
+ PM_SKY130_FD_SC_LP__OR3B_1%C_N
x_PM_SKY130_FD_SC_LP__OR3B_1%A_110_70# N_A_110_70#_M1003_d N_A_110_70#_M1006_d
+ N_A_110_70#_M1008_g N_A_110_70#_M1009_g N_A_110_70#_c_94_n N_A_110_70#_c_98_n
+ N_A_110_70#_c_95_n N_A_110_70#_c_96_n PM_SKY130_FD_SC_LP__OR3B_1%A_110_70#
x_PM_SKY130_FD_SC_LP__OR3B_1%B N_B_M1000_g N_B_M1007_g N_B_c_138_n N_B_c_139_n
+ N_B_c_140_n B B B B N_B_c_142_n PM_SKY130_FD_SC_LP__OR3B_1%B
x_PM_SKY130_FD_SC_LP__OR3B_1%A N_A_M1002_g N_A_M1004_g A A N_A_c_185_n
+ PM_SKY130_FD_SC_LP__OR3B_1%A
x_PM_SKY130_FD_SC_LP__OR3B_1%A_220_74# N_A_220_74#_M1008_s N_A_220_74#_M1007_d
+ N_A_220_74#_M1009_s N_A_220_74#_M1005_g N_A_220_74#_M1001_g
+ N_A_220_74#_c_221_n N_A_220_74#_c_222_n N_A_220_74#_c_223_n
+ N_A_220_74#_c_224_n N_A_220_74#_c_213_n N_A_220_74#_c_225_n
+ N_A_220_74#_c_214_n N_A_220_74#_c_215_n N_A_220_74#_c_216_n
+ N_A_220_74#_c_217_n N_A_220_74#_c_256_n N_A_220_74#_c_218_n
+ N_A_220_74#_c_219_n PM_SKY130_FD_SC_LP__OR3B_1%A_220_74#
x_PM_SKY130_FD_SC_LP__OR3B_1%VPWR N_VPWR_M1006_s N_VPWR_M1004_d N_VPWR_c_302_n
+ N_VPWR_c_303_n N_VPWR_c_304_n VPWR N_VPWR_c_305_n N_VPWR_c_306_n
+ N_VPWR_c_301_n N_VPWR_c_308_n PM_SKY130_FD_SC_LP__OR3B_1%VPWR
x_PM_SKY130_FD_SC_LP__OR3B_1%X N_X_M1005_d N_X_M1001_d N_X_c_338_n X X X X X X
+ N_X_c_340_n PM_SKY130_FD_SC_LP__OR3B_1%X
x_PM_SKY130_FD_SC_LP__OR3B_1%VGND N_VGND_M1003_s N_VGND_M1008_d N_VGND_M1002_d
+ N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n VGND
+ N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n
+ N_VGND_c_367_n PM_SKY130_FD_SC_LP__OR3B_1%VGND
cc_1 VNB N_C_N_c_68_n 0.0241988f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.353
cc_2 VNB N_C_N_M1006_g 0.00643698f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_3 VNB N_C_N_c_70_n 0.0243916f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.55
cc_4 VNB C_N 0.0331722f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_C_N_c_72_n 0.0250662f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_6 VNB N_C_N_c_73_n 0.0249498f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_7 VNB N_A_110_70#_M1008_g 0.0289549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_110_70#_c_94_n 0.00852841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_110_70#_c_95_n 0.0122087f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_10 VNB N_A_110_70#_c_96_n 0.0855188f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=0.925
cc_11 VNB N_B_M1000_g 0.003646f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.88
cc_12 VNB N_B_c_138_n 0.0179399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_139_n 0.0208672f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.55
cc_14 VNB N_B_c_140_n 0.0174606f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_15 VNB B 0.00830752f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_B_c_142_n 0.0152145f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.045
cc_17 VNB N_A_M1002_g 0.0515707f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.88
cc_18 VNB N_A_220_74#_c_213_n 0.00334016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_220_74#_c_214_n 0.00898668f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=1.665
cc_20 VNB N_A_220_74#_c_215_n 0.0356387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_220_74#_c_216_n 0.00383113f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=2.405
cc_22 VNB N_A_220_74#_c_217_n 0.00203784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_220_74#_c_218_n 0.00205003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_220_74#_c_219_n 0.0221229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_301_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_338_n 0.00536733f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.55
cc_27 VNB X 0.0283215f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_28 VNB N_X_c_340_n 0.0231719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_358_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.55
cc_30 VNB N_VGND_c_359_n 0.0216486f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_VGND_c_360_n 0.00871714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_361_n 0.0117205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_362_n 0.0316861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_363_n 0.0197343f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=1.665
cc_35 VNB N_VGND_c_364_n 0.0192239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_365_n 0.215618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_366_n 0.00442399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_367_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_C_N_M1006_g 0.0772608f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_40 VPB C_N 0.0376815f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_41 VPB N_A_110_70#_M1009_g 0.0213894f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_42 VPB N_A_110_70#_c_98_n 0.0310618f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.045
cc_43 VPB N_A_110_70#_c_95_n 0.0079781f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.88
cc_44 VPB N_A_110_70#_c_96_n 0.0179728f $X=-0.19 $Y=1.655 $X2=0.245 $Y2=0.925
cc_45 VPB N_B_M1000_g 0.0181855f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.88
cc_46 VPB B 0.00223979f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_47 VPB N_A_M1002_g 0.0405263f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.88
cc_48 VPB A 0.0250734f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_49 VPB N_A_c_185_n 0.0501255f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_50 VPB N_A_220_74#_M1001_g 0.0280578f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_51 VPB N_A_220_74#_c_221_n 0.00246007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_220_74#_c_222_n 0.00196285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_220_74#_c_223_n 0.017587f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.045
cc_54 VPB N_A_220_74#_c_224_n 0.00889213f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.88
cc_55 VPB N_A_220_74#_c_225_n 0.00162532f $X=-0.19 $Y=1.655 $X2=0.245 $Y2=1.045
cc_56 VPB N_A_220_74#_c_217_n 0.00163027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_302_n 0.0112117f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_58 VPB N_VPWR_c_303_n 0.0216486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_304_n 0.01575f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_60 VPB N_VPWR_c_305_n 0.0561264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_306_n 0.0187803f $X=-0.19 $Y=1.655 $X2=0.245 $Y2=1.295
cc_62 VPB N_VPWR_c_301_n 0.0748358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_308_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB X 0.00719036f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_65 VPB X 0.043257f $X=-0.19 $Y=1.655 $X2=0.245 $Y2=1.665
cc_66 VPB N_X_c_340_n 0.00780156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 C_N N_A_110_70#_c_94_n 0.119573f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_68 N_C_N_c_73_n N_A_110_70#_c_94_n 0.0116283f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_69 N_C_N_c_70_n N_A_110_70#_c_98_n 0.0116283f $X=0.352 $Y=1.55 $X2=0 $Y2=0
cc_70 N_C_N_c_72_n N_A_110_70#_c_95_n 0.0116283f $X=0.32 $Y=1.045 $X2=0 $Y2=0
cc_71 C_N N_A_110_70#_c_96_n 4.89329e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_72 N_C_N_c_72_n N_A_110_70#_c_96_n 0.0349035f $X=0.32 $Y=1.045 $X2=0 $Y2=0
cc_73 N_C_N_M1006_g N_VPWR_c_303_n 0.0144309f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_74 C_N N_VPWR_c_303_n 0.0250477f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_C_N_M1006_g N_VPWR_c_305_n 0.00396895f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_76 N_C_N_M1006_g N_VPWR_c_301_n 0.00796233f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_77 C_N N_VPWR_c_301_n 0.00151387f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_78 C_N N_VGND_c_359_n 0.0250475f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_79 N_C_N_c_72_n N_VGND_c_359_n 0.00156152f $X=0.32 $Y=1.045 $X2=0 $Y2=0
cc_80 N_C_N_c_73_n N_VGND_c_359_n 0.0144309f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_81 N_C_N_c_73_n N_VGND_c_362_n 0.00396895f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_82 C_N N_VGND_c_365_n 0.00151387f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_83 N_C_N_c_73_n N_VGND_c_365_n 0.00796233f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_84 N_A_110_70#_M1008_g N_B_c_138_n 0.0108435f $X=1.44 $Y=0.58 $X2=0 $Y2=0
cc_85 N_A_110_70#_c_96_n N_B_c_139_n 0.0305825f $X=0.955 $Y=1.165 $X2=0 $Y2=0
cc_86 N_A_110_70#_M1009_g N_B_c_140_n 0.0305825f $X=1.44 $Y=2.045 $X2=0 $Y2=0
cc_87 N_A_110_70#_M1008_g B 0.00878976f $X=1.44 $Y=0.58 $X2=0 $Y2=0
cc_88 N_A_110_70#_M1008_g N_B_c_142_n 0.0305825f $X=1.44 $Y=0.58 $X2=0 $Y2=0
cc_89 N_A_110_70#_M1009_g A 5.05838e-19 $X=1.44 $Y=2.045 $X2=0 $Y2=0
cc_90 N_A_110_70#_c_98_n A 0.0109423f $X=0.69 $Y=2.77 $X2=0 $Y2=0
cc_91 N_A_110_70#_M1009_g N_A_220_74#_c_221_n 0.00495656f $X=1.44 $Y=2.045 $X2=0
+ $Y2=0
cc_92 N_A_110_70#_M1009_g N_A_220_74#_c_222_n 0.00164598f $X=1.44 $Y=2.045 $X2=0
+ $Y2=0
cc_93 N_A_110_70#_c_98_n N_A_220_74#_c_222_n 0.0300528f $X=0.69 $Y=2.77 $X2=0
+ $Y2=0
cc_94 N_A_110_70#_c_96_n N_A_220_74#_c_222_n 0.00714526f $X=0.955 $Y=1.165 $X2=0
+ $Y2=0
cc_95 N_A_110_70#_M1009_g N_A_220_74#_c_223_n 0.00918486f $X=1.44 $Y=2.045 $X2=0
+ $Y2=0
cc_96 N_A_110_70#_M1009_g N_A_220_74#_c_224_n 0.0023146f $X=1.44 $Y=2.045 $X2=0
+ $Y2=0
cc_97 N_A_110_70#_c_98_n N_A_220_74#_c_224_n 0.012957f $X=0.69 $Y=2.77 $X2=0
+ $Y2=0
cc_98 N_A_110_70#_M1008_g N_A_220_74#_c_216_n 0.00434514f $X=1.44 $Y=0.58 $X2=0
+ $Y2=0
cc_99 N_A_110_70#_c_94_n N_A_220_74#_c_216_n 0.0236703f $X=0.69 $Y=0.56 $X2=0
+ $Y2=0
cc_100 N_A_110_70#_c_96_n N_A_220_74#_c_216_n 0.00642725f $X=0.955 $Y=1.165
+ $X2=0 $Y2=0
cc_101 N_A_110_70#_M1008_g N_A_220_74#_c_217_n 0.00723064f $X=1.44 $Y=0.58 $X2=0
+ $Y2=0
cc_102 N_A_110_70#_M1009_g N_A_220_74#_c_217_n 0.00521738f $X=1.44 $Y=2.045
+ $X2=0 $Y2=0
cc_103 N_A_110_70#_c_94_n N_A_220_74#_c_217_n 0.00915199f $X=0.69 $Y=0.56 $X2=0
+ $Y2=0
cc_104 N_A_110_70#_c_98_n N_A_220_74#_c_217_n 0.00731686f $X=0.69 $Y=2.77 $X2=0
+ $Y2=0
cc_105 N_A_110_70#_c_95_n N_A_220_74#_c_217_n 0.0491125f $X=0.955 $Y=1.165 $X2=0
+ $Y2=0
cc_106 N_A_110_70#_c_96_n N_A_220_74#_c_217_n 0.0317193f $X=0.955 $Y=1.165 $X2=0
+ $Y2=0
cc_107 N_A_110_70#_c_98_n N_VPWR_c_305_n 0.00930971f $X=0.69 $Y=2.77 $X2=0 $Y2=0
cc_108 N_A_110_70#_c_98_n N_VPWR_c_301_n 0.00926582f $X=0.69 $Y=2.77 $X2=0 $Y2=0
cc_109 N_A_110_70#_M1008_g N_VGND_c_360_n 0.00335484f $X=1.44 $Y=0.58 $X2=0
+ $Y2=0
cc_110 N_A_110_70#_M1008_g N_VGND_c_362_n 0.0043575f $X=1.44 $Y=0.58 $X2=0 $Y2=0
cc_111 N_A_110_70#_c_94_n N_VGND_c_362_n 0.00930971f $X=0.69 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A_110_70#_M1008_g N_VGND_c_365_n 0.00827011f $X=1.44 $Y=0.58 $X2=0
+ $Y2=0
cc_113 N_A_110_70#_c_94_n N_VGND_c_365_n 0.00926582f $X=0.69 $Y=0.56 $X2=0 $Y2=0
cc_114 N_B_M1000_g N_A_M1002_g 0.0229668f $X=1.8 $Y=2.045 $X2=0 $Y2=0
cc_115 N_B_c_138_n N_A_M1002_g 0.0115764f $X=1.89 $Y=0.9 $X2=0 $Y2=0
cc_116 B N_A_M1002_g 0.00240625f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_117 N_B_c_142_n N_A_M1002_g 0.0412718f $X=1.89 $Y=1.065 $X2=0 $Y2=0
cc_118 N_B_M1000_g A 8.92655e-19 $X=1.8 $Y=2.045 $X2=0 $Y2=0
cc_119 N_B_M1000_g N_A_220_74#_c_221_n 8.4952e-19 $X=1.8 $Y=2.045 $X2=0 $Y2=0
cc_120 N_B_c_140_n N_A_220_74#_c_221_n 3.1423e-19 $X=1.89 $Y=1.57 $X2=0 $Y2=0
cc_121 N_B_c_139_n N_A_220_74#_c_222_n 3.1423e-19 $X=1.89 $Y=1.405 $X2=0 $Y2=0
cc_122 N_B_M1000_g N_A_220_74#_c_223_n 0.0076289f $X=1.8 $Y=2.045 $X2=0 $Y2=0
cc_123 B N_A_220_74#_c_223_n 0.0275634f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_124 N_B_c_138_n N_A_220_74#_c_213_n 0.00358411f $X=1.89 $Y=0.9 $X2=0 $Y2=0
cc_125 B N_A_220_74#_c_213_n 0.0350544f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_126 N_B_c_142_n N_A_220_74#_c_213_n 0.00260225f $X=1.89 $Y=1.065 $X2=0 $Y2=0
cc_127 N_B_M1000_g N_A_220_74#_c_225_n 0.00453918f $X=1.8 $Y=2.045 $X2=0 $Y2=0
cc_128 B N_A_220_74#_c_225_n 0.0363108f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_129 N_B_c_138_n N_A_220_74#_c_216_n 8.06752e-19 $X=1.89 $Y=0.9 $X2=0 $Y2=0
cc_130 B N_A_220_74#_c_217_n 0.0876944f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_131 N_B_c_142_n N_A_220_74#_c_217_n 3.1423e-19 $X=1.89 $Y=1.065 $X2=0 $Y2=0
cc_132 N_B_c_138_n N_A_220_74#_c_256_n 0.00378744f $X=1.89 $Y=0.9 $X2=0 $Y2=0
cc_133 B N_A_220_74#_c_256_n 0.0010755f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_134 N_B_c_142_n N_A_220_74#_c_256_n 0.00179723f $X=1.89 $Y=1.065 $X2=0 $Y2=0
cc_135 N_B_M1000_g N_A_220_74#_c_218_n 2.77264e-19 $X=1.8 $Y=2.045 $X2=0 $Y2=0
cc_136 N_B_c_139_n N_A_220_74#_c_218_n 0.00181041f $X=1.89 $Y=1.405 $X2=0 $Y2=0
cc_137 B N_A_220_74#_c_218_n 0.0273841f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_138 B A_303_367# 0.00106497f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_139 B A_375_367# 0.00318116f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_140 N_B_c_138_n N_VGND_c_360_n 0.00335484f $X=1.89 $Y=0.9 $X2=0 $Y2=0
cc_141 B N_VGND_c_360_n 0.0194534f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_142 N_B_c_142_n N_VGND_c_360_n 3.97629e-19 $X=1.89 $Y=1.065 $X2=0 $Y2=0
cc_143 N_B_c_138_n N_VGND_c_363_n 0.00434051f $X=1.89 $Y=0.9 $X2=0 $Y2=0
cc_144 N_B_c_138_n N_VGND_c_365_n 0.00446966f $X=1.89 $Y=0.9 $X2=0 $Y2=0
cc_145 B N_VGND_c_365_n 0.00663019f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_A_220_74#_M1001_g 0.0178327f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_147 N_A_M1002_g N_A_220_74#_c_223_n 0.00636162f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_148 A N_A_220_74#_c_223_n 0.0711098f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_149 N_A_c_185_n N_A_220_74#_c_223_n 0.00174302f $X=2.34 $Y=2.855 $X2=0 $Y2=0
cc_150 N_A_M1002_g N_A_220_74#_c_213_n 0.012905f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_151 N_A_M1002_g N_A_220_74#_c_225_n 0.0152305f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_152 N_A_M1002_g N_A_220_74#_c_214_n 0.0145879f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_A_220_74#_c_215_n 0.0180878f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_A_220_74#_c_256_n 0.00439829f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_A_220_74#_c_218_n 0.00371475f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_156 N_A_M1002_g N_A_220_74#_c_219_n 0.0137189f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_157 N_A_M1002_g N_VPWR_c_304_n 0.0114547f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_158 A N_VPWR_c_304_n 0.0311145f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_159 A N_VPWR_c_305_n 0.0443668f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_160 N_A_c_185_n N_VPWR_c_305_n 0.0103159f $X=2.34 $Y=2.855 $X2=0 $Y2=0
cc_161 A N_VPWR_c_301_n 0.0329853f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_162 N_A_c_185_n N_VPWR_c_301_n 0.0135938f $X=2.34 $Y=2.855 $X2=0 $Y2=0
cc_163 N_A_M1002_g N_VGND_c_361_n 0.00831486f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_164 N_A_M1002_g N_VGND_c_363_n 0.00395672f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_165 N_A_M1002_g N_VGND_c_365_n 0.00690805f $X=2.34 $Y=0.58 $X2=0 $Y2=0
cc_166 N_A_220_74#_M1001_g N_VPWR_c_304_n 0.00585774f $X=2.865 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_220_74#_c_223_n N_VPWR_c_304_n 0.0140122f $X=2.155 $Y=2.385 $X2=0
+ $Y2=0
cc_168 N_A_220_74#_c_225_n N_VPWR_c_304_n 0.0348952f $X=2.24 $Y=2.3 $X2=0 $Y2=0
cc_169 N_A_220_74#_c_214_n N_VPWR_c_304_n 0.0224144f $X=2.82 $Y=1.485 $X2=0
+ $Y2=0
cc_170 N_A_220_74#_c_215_n N_VPWR_c_304_n 0.00230627f $X=2.82 $Y=1.485 $X2=0
+ $Y2=0
cc_171 N_A_220_74#_M1001_g N_VPWR_c_306_n 0.00585385f $X=2.865 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_220_74#_M1001_g N_VPWR_c_301_n 0.0128414f $X=2.865 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_220_74#_c_223_n N_VPWR_c_301_n 0.00233445f $X=2.155 $Y=2.385 $X2=0
+ $Y2=0
cc_174 N_A_220_74#_c_224_n N_VPWR_c_301_n 0.0127005f $X=1.39 $Y=2.385 $X2=0
+ $Y2=0
cc_175 N_A_220_74#_c_225_n A_375_367# 0.00421038f $X=2.24 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_220_74#_c_219_n X 0.00223205f $X=2.82 $Y=1.32 $X2=0 $Y2=0
cc_177 N_A_220_74#_M1001_g X 0.00343671f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_220_74#_c_215_n X 2.71753e-19 $X=2.82 $Y=1.485 $X2=0 $Y2=0
cc_179 N_A_220_74#_M1001_g N_X_c_340_n 0.00402789f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_220_74#_c_214_n N_X_c_340_n 0.0250942f $X=2.82 $Y=1.485 $X2=0 $Y2=0
cc_181 N_A_220_74#_c_215_n N_X_c_340_n 0.00810943f $X=2.82 $Y=1.485 $X2=0 $Y2=0
cc_182 N_A_220_74#_c_219_n N_X_c_340_n 0.00385201f $X=2.82 $Y=1.32 $X2=0 $Y2=0
cc_183 N_A_220_74#_c_213_n N_VGND_c_361_n 0.035359f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_184 N_A_220_74#_c_214_n N_VGND_c_361_n 0.0210682f $X=2.82 $Y=1.485 $X2=0
+ $Y2=0
cc_185 N_A_220_74#_c_215_n N_VGND_c_361_n 0.00224228f $X=2.82 $Y=1.485 $X2=0
+ $Y2=0
cc_186 N_A_220_74#_c_256_n N_VGND_c_361_n 0.0214585f $X=2.24 $Y=0.53 $X2=0 $Y2=0
cc_187 N_A_220_74#_c_219_n N_VGND_c_361_n 0.00367574f $X=2.82 $Y=1.32 $X2=0
+ $Y2=0
cc_188 N_A_220_74#_c_216_n N_VGND_c_362_n 0.0098881f $X=1.225 $Y=0.585 $X2=0
+ $Y2=0
cc_189 N_A_220_74#_c_256_n N_VGND_c_363_n 0.010891f $X=2.24 $Y=0.53 $X2=0 $Y2=0
cc_190 N_A_220_74#_c_219_n N_VGND_c_364_n 0.00461464f $X=2.82 $Y=1.32 $X2=0
+ $Y2=0
cc_191 N_A_220_74#_c_216_n N_VGND_c_365_n 0.0113119f $X=1.225 $Y=0.585 $X2=0
+ $Y2=0
cc_192 N_A_220_74#_c_256_n N_VGND_c_365_n 0.0123102f $X=2.24 $Y=0.53 $X2=0 $Y2=0
cc_193 N_A_220_74#_c_219_n N_VGND_c_365_n 0.00912455f $X=2.82 $Y=1.32 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_301_n N_X_M1001_d 0.00336915f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_304_n X 9.42942e-19 $X=2.605 $Y=1.985 $X2=0 $Y2=0
cc_196 N_VPWR_c_306_n X 0.0188828f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_301_n X 0.010808f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_198 X N_VGND_c_361_n 0.00127971f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_199 X N_VGND_c_364_n 0.0124046f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_200 X N_VGND_c_365_n 0.0102675f $X=3.035 $Y=0.47 $X2=0 $Y2=0
