# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 0.840000 0.915000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.350000 0.255000 5.665000 1.095000 ;
        RECT 5.350000 1.815000 5.665000 3.075000 ;
        RECT 5.495000 1.095000 5.665000 1.815000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325000 0.375000 7.595000 3.075000 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.255000 1.775000 1.115000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 0.660000  0.085000 0.915000 0.670000 ;
        RECT 2.340000  0.085000 2.670000 0.575000 ;
        RECT 4.075000  0.085000 4.530000 0.805000 ;
        RECT 5.835000  0.085000 6.135000 1.170000 ;
        RECT 6.825000  0.085000 7.155000 1.175000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.725000 2.075000 0.985000 3.245000 ;
        RECT 2.295000 2.765000 2.555000 3.245000 ;
        RECT 4.020000 2.355000 4.730000 3.245000 ;
        RECT 4.400000 2.115000 4.730000 2.355000 ;
        RECT 5.835000 1.815000 6.135000 3.245000 ;
        RECT 6.825000 1.845000 7.155000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.340000 0.490000 0.670000 ;
      RECT 0.085000 0.670000 0.285000 1.705000 ;
      RECT 0.085000 1.705000 2.680000 1.905000 ;
      RECT 0.260000 1.905000 0.555000 2.755000 ;
      RECT 1.085000 0.365000 1.360000 1.285000 ;
      RECT 1.085000 1.285000 2.320000 1.365000 ;
      RECT 1.085000 1.365000 3.140000 1.535000 ;
      RECT 1.155000 2.075000 3.140000 2.255000 ;
      RECT 1.155000 2.255000 1.450000 2.755000 ;
      RECT 1.795000 2.425000 3.510000 2.595000 ;
      RECT 1.795000 2.595000 2.125000 3.075000 ;
      RECT 1.945000 0.280000 2.135000 0.745000 ;
      RECT 1.945000 0.745000 3.310000 0.915000 ;
      RECT 1.990000 1.085000 2.320000 1.285000 ;
      RECT 2.890000 1.535000 3.140000 2.075000 ;
      RECT 3.015000 2.765000 3.850000 3.075000 ;
      RECT 3.050000 0.915000 3.310000 1.015000 ;
      RECT 3.050000 1.015000 3.510000 1.185000 ;
      RECT 3.225000 0.275000 3.650000 0.575000 ;
      RECT 3.310000 1.185000 3.510000 2.425000 ;
      RECT 3.480000 0.575000 3.650000 0.665000 ;
      RECT 3.480000 0.665000 3.850000 0.835000 ;
      RECT 3.680000 0.835000 3.850000 0.975000 ;
      RECT 3.680000 0.975000 4.550000 1.145000 ;
      RECT 3.680000 1.145000 3.850000 2.765000 ;
      RECT 4.020000 1.315000 4.210000 1.775000 ;
      RECT 4.020000 1.775000 5.160000 1.945000 ;
      RECT 4.020000 1.945000 4.210000 1.985000 ;
      RECT 4.380000 1.145000 4.550000 1.185000 ;
      RECT 4.380000 1.185000 4.755000 1.515000 ;
      RECT 4.720000 0.255000 5.105000 1.005000 ;
      RECT 4.900000 1.945000 5.160000 3.055000 ;
      RECT 4.935000 1.005000 5.105000 1.265000 ;
      RECT 4.935000 1.265000 5.315000 1.595000 ;
      RECT 4.935000 1.595000 5.160000 1.775000 ;
      RECT 6.305000 0.790000 6.635000 1.345000 ;
      RECT 6.305000 1.345000 7.155000 1.675000 ;
      RECT 6.305000 1.675000 6.635000 2.495000 ;
  END
END sky130_fd_sc_lp__dlxbp_1
