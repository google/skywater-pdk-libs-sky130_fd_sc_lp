* File: sky130_fd_sc_lp__einvn_0.pex.spice
* Created: Wed Sep  2 09:51:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVN_0%A_28_141# 1 2 7 9 12 16 18 23
c35 18 0 1.54446e-20 $X=0.93 $Y=0.43
r36 19 23 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=0.93 $Y=0.43
+ $X2=1.045 $Y2=0.43
r37 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=0.43 $X2=0.93 $Y2=0.43
r38 16 18 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.43 $Y=0.43 $X2=0.93
+ $Y2=0.43
r39 12 14 59.3683 $w=3.28e-07 $l=1.7e-06 $layer=LI1_cond $X=0.265 $Y=0.915
+ $X2=0.265 $Y2=2.615
r40 10 16 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=0.265 $Y=0.595
+ $X2=0.43 $Y2=0.43
r41 10 12 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.265 $Y=0.595
+ $X2=0.265 $Y2=0.915
r42 7 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=0.595
+ $X2=1.045 $Y2=0.43
r43 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.045 $Y=0.595
+ $X2=1.045 $Y2=0.915
r44 2 14 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.405 $X2=0.305 $Y2=2.615
r45 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.705 $X2=0.265 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_0%TE_B 3 6 9 13 18 20 21 22 27
r44 27 29 47.4991 $w=4.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.71
+ $X2=0.64 $Y2=1.545
r45 21 22 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.737 $Y=1.665
+ $X2=0.737 $Y2=2.035
r46 21 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=1.71 $X2=0.71 $Y2=1.71
r47 20 21 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.737 $Y=1.295
+ $X2=0.737 $Y2=1.665
r48 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.045 $Y=2.215
+ $X2=1.045 $Y2=2.14
r49 11 13 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.045 $Y=2.215
+ $X2=1.045 $Y2=2.725
r50 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=2.215
+ $X2=0.52 $Y2=2.14
r51 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.52 $Y=2.215 $X2=0.52
+ $Y2=2.615
r52 6 18 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.64 $Y=2.14
+ $X2=1.045 $Y2=2.14
r53 6 15 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=0.64 $Y=2.14 $X2=0.52
+ $Y2=2.14
r54 5 27 8.28314 $w=4.7e-07 $l=7e-08 $layer=POLY_cond $X=0.64 $Y=1.78 $X2=0.64
+ $Y2=1.71
r55 5 6 33.7242 $w=4.7e-07 $l=2.85e-07 $layer=POLY_cond $X=0.64 $Y=1.78 $X2=0.64
+ $Y2=2.065
r56 3 29 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.48 $Y=0.915
+ $X2=0.48 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_0%A 3 7 9 10 11 12 13 20
c37 3 0 1.54446e-20 $X=1.435 $Y=0.915
r38 20 23 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.312 $Y=1.66
+ $X2=1.312 $Y2=1.825
r39 20 22 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.312 $Y=1.66
+ $X2=1.312 $Y2=1.495
r40 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.24 $Y=2.405
+ $X2=1.24 $Y2=2.775
r41 11 12 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.24 $Y=2.035
+ $X2=1.24 $Y2=2.405
r42 10 11 16.0062 $w=2.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.24 $Y=1.66
+ $X2=1.24 $Y2=2.035
r43 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.66 $X2=1.28 $Y2=1.66
r44 9 10 15.5793 $w=2.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.24 $Y=1.295
+ $X2=1.24 $Y2=1.66
r45 7 23 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.435 $Y=2.725
+ $X2=1.435 $Y2=1.825
r46 3 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.435 $Y=0.915
+ $X2=1.435 $Y2=1.495
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_0%VPWR 1 6 8 10 17 18 21
r25 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 15 21 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.767 $Y2=3.33
r28 15 17 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 21 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.767 $Y2=3.33
r32 10 12 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33 $X2=0.24
+ $Y2=3.33
r33 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 4 21 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.767 $Y=3.245
+ $X2=0.767 $Y2=3.33
r36 4 6 24.0809 $w=3.33e-07 $l=7e-07 $layer=LI1_cond $X=0.767 $Y=3.245 $X2=0.767
+ $Y2=2.545
r37 1 6 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.405 $X2=0.765 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_0%Z 1 2 7 8 9 10 11 12
r10 12 32 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.69 $Y=2.775
+ $X2=1.69 $Y2=2.55
r11 11 32 5.76222 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.69 $Y=2.405
+ $X2=1.69 $Y2=2.55
r12 10 11 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=2.035
+ $X2=1.69 $Y2=2.405
r13 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=1.665
+ $X2=1.69 $Y2=2.035
r14 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=1.295 $X2=1.69
+ $Y2=1.665
r15 7 8 15.101 $w=2.88e-07 $l=3.8e-07 $layer=LI1_cond $X=1.69 $Y=0.915 $X2=1.69
+ $Y2=1.295
r16 2 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=2.405 $X2=1.65 $Y2=2.55
r17 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.705 $X2=1.65 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_0%VGND 1 4 9 10 12 19 20 23
r30 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r31 20 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r32 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r33 17 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.28
+ $Y2=0
r34 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.68
+ $Y2=0
r35 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 12 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.28
+ $Y2=0
r37 12 14 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=0.24
+ $Y2=0
r38 10 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r39 10 15 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r40 8 23 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085 $X2=1.28
+ $Y2=0
r41 8 9 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.28 $Y=0.085 $X2=1.28
+ $Y2=0.775
r42 4 9 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=1.195 $Y=0.907
+ $X2=1.28 $Y2=0.775
r43 4 6 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=1.195 $Y=0.907 $X2=0.765
+ $Y2=0.907
r44 1 6 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.705 $X2=0.765 $Y2=0.9
.ends

