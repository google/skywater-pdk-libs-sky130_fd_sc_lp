* File: sky130_fd_sc_lp__a2bb2oi_2.pex.spice
* Created: Wed Sep  2 09:24:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%B1 3 7 11 15 17 20 23 25 27 28 31 32 33
c86 23 0 1.73586e-19 $X=0.64 $Y=1.92
c87 15 0 2.55454e-19 $X=1.94 $Y=2.465
r88 32 33 14.7198 $w=3.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.2 $Y=2.02
+ $X2=1.595 $Y2=2.02
r89 31 46 3.24051 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=0.64 $Y=2.02 $X2=0.73
+ $Y2=2.02
r90 31 32 24.0118 $w=1.98e-07 $l=4.33e-07 $layer=LI1_cond $X=0.767 $Y=2.02
+ $X2=1.2 $Y2=2.02
r91 31 46 2.05182 $w=1.98e-07 $l=3.7e-08 $layer=LI1_cond $X=0.767 $Y=2.02
+ $X2=0.73 $Y2=2.02
r92 28 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.51
+ $X2=1.85 $Y2=1.675
r93 28 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.51
+ $X2=1.85 $Y2=1.345
r94 27 30 5.17595 $w=4.18e-07 $l=1.45e-07 $layer=LI1_cond $X=1.805 $Y=1.51
+ $X2=1.805 $Y2=1.655
r95 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.51 $X2=1.85 $Y2=1.51
r96 25 33 2.93074 $w=2.85e-07 $l=1e-07 $layer=LI1_cond $X=1.737 $Y=1.92
+ $X2=1.737 $Y2=2.02
r97 25 30 10.7157 $w=2.83e-07 $l=2.65e-07 $layer=LI1_cond $X=1.737 $Y=1.92
+ $X2=1.737 $Y2=1.655
r98 23 31 3.60057 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=0.64 $Y=1.92 $X2=0.64
+ $Y2=2.02
r99 22 23 18.1768 $w=1.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.64 $Y=1.625
+ $X2=0.64 $Y2=1.92
r100 20 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.4 $Y=1.46
+ $X2=0.4 $Y2=1.625
r101 20 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.4 $Y=1.46
+ $X2=0.4 $Y2=1.295
r102 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.4
+ $Y=1.46 $X2=0.4 $Y2=1.46
r103 17 22 7.0541 $w=2.5e-07 $l=1.63936e-07 $layer=LI1_cond $X=0.55 $Y=1.5
+ $X2=0.64 $Y2=1.625
r104 17 19 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=0.55 $Y=1.5 $X2=0.4
+ $Y2=1.5
r105 15 44 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.94 $Y=2.465
+ $X2=1.94 $Y2=1.675
r106 11 43 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.86 $Y=0.745 $X2=1.86
+ $Y2=1.345
r107 7 41 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.49 $Y=2.465
+ $X2=0.49 $Y2=1.625
r108 3 40 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.49 $Y=0.745
+ $X2=0.49 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%B2 3 7 11 15 17 23 24
c50 23 0 6.47804e-20 $X=1.075 $Y=1.51
r51 22 24 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=1.075 $Y=1.51
+ $X2=1.35 $Y2=1.51
r52 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.51 $X2=1.075 $Y2=1.51
r53 19 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.92 $Y=1.51
+ $X2=1.075 $Y2=1.51
r54 17 23 3.59985 $w=5.13e-07 $l=1.55e-07 $layer=LI1_cond $X=1.167 $Y=1.665
+ $X2=1.167 $Y2=1.51
r55 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.675
+ $X2=1.35 $Y2=1.51
r56 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.35 $Y=1.675
+ $X2=1.35 $Y2=2.465
r57 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.345
+ $X2=1.35 $Y2=1.51
r58 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.35 $Y=1.345 $X2=1.35
+ $Y2=0.745
r59 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.675
+ $X2=0.92 $Y2=1.51
r60 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.92 $Y=1.675 $X2=0.92
+ $Y2=2.465
r61 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.345
+ $X2=0.92 $Y2=1.51
r62 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.92 $Y=1.345 $X2=0.92
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%A_459_39# 1 2 3 12 16 18 20 22 25 27 29 30
+ 34 37 38 41 44 45 46 47 48 51 55 59
c118 44 0 2.64564e-19 $X=4.22 $Y=1.705
c119 12 0 6.78225e-20 $X=2.37 $Y=0.745
r120 57 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.05 $Y=1.16
+ $X2=4.22 $Y2=1.16
r121 53 55 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.91 $Y=1.075
+ $X2=4.91 $Y2=0.47
r122 49 51 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=4.895 $Y=1.875
+ $X2=4.895 $Y2=1.98
r123 47 49 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.785 $Y=1.79
+ $X2=4.895 $Y2=1.875
r124 47 48 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.785 $Y=1.79
+ $X2=4.305 $Y2=1.79
r125 46 58 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=1.16
+ $X2=4.22 $Y2=1.16
r126 45 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.825 $Y=1.16
+ $X2=4.91 $Y2=1.075
r127 45 46 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.825 $Y=1.16
+ $X2=4.305 $Y2=1.16
r128 44 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.22 $Y=1.705
+ $X2=4.305 $Y2=1.79
r129 43 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.22 $Y=1.245
+ $X2=4.22 $Y2=1.16
r130 43 44 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.22 $Y=1.245
+ $X2=4.22 $Y2=1.705
r131 39 57 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=1.075
+ $X2=4.05 $Y2=1.16
r132 39 41 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=4.05 $Y=1.075
+ $X2=4.05 $Y2=0.47
r133 37 57 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.955 $Y=1.16
+ $X2=4.05 $Y2=1.16
r134 37 38 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.955 $Y=1.16
+ $X2=3.335 $Y2=1.16
r135 35 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.25 $Y=1.44 $X2=3.25
+ $Y2=1.35
r136 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.44 $X2=3.25 $Y2=1.44
r137 32 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.21 $Y=1.245
+ $X2=3.335 $Y2=1.16
r138 32 34 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=3.21 $Y=1.245
+ $X2=3.21 $Y2=1.44
r139 30 31 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.8 $Y=1.35 $X2=2.8
+ $Y2=1.5
r140 28 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=1.35
+ $X2=2.8 $Y2=1.35
r141 27 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.35
+ $X2=3.25 $Y2=1.35
r142 27 28 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.085 $Y=1.35
+ $X2=2.875 $Y2=1.35
r143 23 31 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.8 $Y=1.575
+ $X2=2.8 $Y2=1.5
r144 23 25 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.8 $Y=1.575
+ $X2=2.8 $Y2=2.465
r145 20 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.8 $Y=1.275
+ $X2=2.8 $Y2=1.35
r146 20 22 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.8 $Y=1.275
+ $X2=2.8 $Y2=0.745
r147 19 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.5
+ $X2=2.37 $Y2=1.5
r148 18 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.725 $Y=1.5
+ $X2=2.8 $Y2=1.5
r149 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.725 $Y=1.5
+ $X2=2.445 $Y2=1.5
r150 14 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.575
+ $X2=2.37 $Y2=1.5
r151 14 16 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.37 $Y=1.575
+ $X2=2.37 $Y2=2.465
r152 10 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.425
+ $X2=2.37 $Y2=1.5
r153 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.37 $Y=1.425
+ $X2=2.37 $Y2=0.745
r154 3 51 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.77
+ $Y=1.835 $X2=4.91 $Y2=1.98
r155 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.77
+ $Y=0.325 $X2=4.91 $Y2=0.47
r156 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.91
+ $Y=0.325 $X2=4.05 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%A1_N 3 7 11 15 17 21 24
c58 7 0 8.27999e-20 $X=3.835 $Y=2.465
r59 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.835 $Y=1.51
+ $X2=4.265 $Y2=1.51
r60 20 23 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.79 $Y=1.51
+ $X2=3.835 $Y2=1.51
r61 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.79
+ $Y=1.51 $X2=3.79 $Y2=1.51
r62 17 21 4.94032 $w=4.58e-07 $l=1.9e-07 $layer=LI1_cond $X=3.6 $Y=1.645
+ $X2=3.79 $Y2=1.645
r63 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.675
+ $X2=4.265 $Y2=1.51
r64 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.265 $Y=1.675
+ $X2=4.265 $Y2=2.465
r65 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.345
+ $X2=4.265 $Y2=1.51
r66 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.265 $Y=1.345 $X2=4.265
+ $Y2=0.745
r67 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.675
+ $X2=3.835 $Y2=1.51
r68 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.835 $Y=1.675
+ $X2=3.835 $Y2=2.465
r69 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.345
+ $X2=3.835 $Y2=1.51
r70 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.835 $Y=1.345 $X2=3.835
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%A2_N 1 3 6 8 12 15 17 18 19 23
r46 25 27 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=5.237 $Y=1.44
+ $X2=5.237 $Y2=1.605
r47 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.26
+ $Y=1.44 $X2=5.26 $Y2=1.44
r48 19 26 5.38235 $w=4.98e-07 $l=2.25e-07 $layer=LI1_cond $X=5.425 $Y=1.665
+ $X2=5.425 $Y2=1.44
r49 18 26 3.46863 $w=4.98e-07 $l=1.45e-07 $layer=LI1_cond $X=5.425 $Y=1.295
+ $X2=5.425 $Y2=1.44
r50 15 27 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.125 $Y=2.465
+ $X2=5.125 $Y2=1.605
r51 12 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.125 $Y=0.745
+ $X2=5.125 $Y2=1.275
r52 9 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.77 $Y=1.35
+ $X2=4.695 $Y2=1.35
r53 8 25 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=5.237 $Y=1.35
+ $X2=5.237 $Y2=1.44
r54 8 23 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=5.237 $Y=1.35
+ $X2=5.237 $Y2=1.275
r55 8 9 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.05 $Y=1.35 $X2=4.77
+ $Y2=1.35
r56 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.695 $Y=1.425
+ $X2=4.695 $Y2=1.35
r57 4 6 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.695 $Y=1.425
+ $X2=4.695 $Y2=2.465
r58 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.695 $Y=1.275
+ $X2=4.695 $Y2=1.35
r59 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.695 $Y=1.275
+ $X2=4.695 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%A_30_367# 1 2 3 4 15 19 21 25 29 33 34 35
+ 37 39 41
r61 35 45 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=2.99
r62 35 37 40.5571 $w=2.58e-07 $l=9.15e-07 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=1.99
r63 33 45 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.92 $Y=2.99 $X2=3.05
+ $Y2=2.99
r64 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.92 $Y=2.99
+ $X2=2.25 $Y2=2.99
r65 32 34 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.25 $Y2=2.99
r66 31 43 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=2.46 $X2=2.15
+ $Y2=2.375
r67 31 32 24.6773 $w=1.98e-07 $l=4.45e-07 $layer=LI1_cond $X=2.15 $Y=2.46
+ $X2=2.15 $Y2=2.905
r68 27 43 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=2.29 $X2=2.15
+ $Y2=2.375
r69 27 29 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=2.15 $Y=2.29 $X2=2.15
+ $Y2=1.99
r70 26 41 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.24 $Y=2.375 $X2=1.14
+ $Y2=2.375
r71 25 43 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.05 $Y=2.375 $X2=2.15
+ $Y2=2.375
r72 25 26 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.05 $Y=2.375
+ $X2=1.24 $Y2=2.375
r73 22 39 2.98021 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.38 $Y=2.375
+ $X2=0.245 $Y2=2.375
r74 21 41 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.04 $Y=2.375 $X2=1.14
+ $Y2=2.375
r75 21 22 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.04 $Y=2.375
+ $X2=0.38 $Y2=2.375
r76 17 39 3.52026 $w=2.65e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.245 $Y2=2.375
r77 17 19 0.443247 $w=2.58e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=2.46 $X2=0.24
+ $Y2=2.47
r78 13 39 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.29
+ $X2=0.245 $Y2=2.375
r79 13 15 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.245 $Y=2.29
+ $X2=0.245 $Y2=1.98
r80 4 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.835 $X2=3.015 $Y2=2.91
r81 4 37 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.835 $X2=3.015 $Y2=1.99
r82 3 43 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.835 $X2=2.155 $Y2=2.44
r83 3 29 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.835 $X2=2.155 $Y2=1.99
r84 2 41 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.455
r85 1 19 300 $w=1.7e-07 $l=6.94694e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.47
r86 1 15 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%VPWR 1 2 3 12 16 20 22 24 29 34 47 48 51
+ 54 57
r77 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r82 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r83 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=5.52
+ $Y2=3.33
r84 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r85 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.05 $Y2=3.33
r86 42 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 41 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r89 38 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r90 37 40 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r91 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r92 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=1.655 $Y2=3.33
r93 35 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 34 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=4.05 $Y2=3.33
r95 34 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=3.6 $Y2=3.33
r96 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r97 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r99 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=3.33
+ $X2=0.705 $Y2=3.33
r100 30 32 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.87 $Y=3.33
+ $X2=1.2 $Y2=3.33
r101 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.655 $Y2=3.33
r102 29 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 27 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 24 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=3.33
+ $X2=0.705 $Y2=3.33
r106 24 26 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.54 $Y=3.33 $X2=0.24
+ $Y2=3.33
r107 22 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 22 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 18 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=3.245
+ $X2=4.05 $Y2=3.33
r110 18 20 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=4.05 $Y=3.245
+ $X2=4.05 $Y2=2.49
r111 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=3.245
+ $X2=1.655 $Y2=3.33
r112 14 16 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.655 $Y=3.245
+ $X2=1.655 $Y2=2.775
r113 10 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=3.245
+ $X2=0.705 $Y2=3.33
r114 10 12 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.705 $Y=3.245
+ $X2=0.705 $Y2=2.775
r115 3 20 300 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=2 $X=3.91
+ $Y=1.835 $X2=4.05 $Y2=2.49
r116 2 16 600 $w=1.7e-07 $l=1.04871e-06 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.655 $Y2=2.775
r117 1 12 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%Y 1 2 3 12 14 15 18 20 24 26 27 28 32
c58 26 0 1.3523e-19 $X=2.62 $Y=1.16
c59 18 0 1.90673e-19 $X=2.585 $Y=1.97
r60 27 28 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=0.555
+ $X2=2.62 $Y2=0.925
r61 27 32 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.62 $Y=0.555
+ $X2=2.62 $Y2=0.45
r62 25 28 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=2.62 $Y=1.075
+ $X2=2.62 $Y2=0.925
r63 25 26 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.075
+ $X2=2.62 $Y2=1.16
r64 22 26 3.64284 $w=2.55e-07 $l=8.74643e-08 $layer=LI1_cond $X=2.625 $Y=1.245
+ $X2=2.62 $Y2=1.16
r65 22 24 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=2.625 $Y=1.245
+ $X2=2.625 $Y2=1.805
r66 18 24 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=1.97
+ $X2=2.585 $Y2=1.805
r67 18 20 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.585 $Y=1.97
+ $X2=2.585 $Y2=2.65
r68 14 26 2.83584 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.49 $Y=1.16 $X2=2.62
+ $Y2=1.16
r69 14 15 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.49 $Y=1.16
+ $X2=1.3 $Y2=1.16
r70 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.135 $Y=1.075
+ $X2=1.3 $Y2=1.16
r71 10 12 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.135 $Y=1.075
+ $X2=1.135 $Y2=0.7
r72 3 20 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.835 $X2=2.585 $Y2=2.65
r73 3 18 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.835 $X2=2.585 $Y2=1.97
r74 2 32 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.325 $X2=2.585 $Y2=0.45
r75 1 12 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.325 $X2=1.135 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%A_699_367# 1 2 3 10 12 14 16 17 18 20 22
r40 20 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=2.905 $X2=5.34
+ $Y2=2.99
r41 20 22 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=5.34 $Y=2.905
+ $X2=5.34 $Y2=2.085
r42 19 29 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.615 $Y=2.99
+ $X2=4.5 $Y2=2.99
r43 18 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=2.99
+ $X2=5.34 $Y2=2.99
r44 18 19 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.175 $Y=2.99
+ $X2=4.615 $Y2=2.99
r45 17 29 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=2.905 $X2=4.5
+ $Y2=2.99
r46 16 27 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=2.215 $X2=4.5
+ $Y2=2.13
r47 16 17 34.5733 $w=2.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4.5 $Y=2.215 $X2=4.5
+ $Y2=2.905
r48 15 25 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.715 $Y=2.13
+ $X2=3.585 $Y2=2.13
r49 14 27 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.385 $Y=2.13
+ $X2=4.5 $Y2=2.13
r50 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.385 $Y=2.13
+ $X2=3.715 $Y2=2.13
r51 10 25 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=2.215
+ $X2=3.585 $Y2=2.13
r52 10 12 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=3.585 $Y=2.215
+ $X2=3.585 $Y2=2.91
r53 3 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.835 $X2=5.34 $Y2=2.91
r54 3 22 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.835 $X2=5.34 $Y2=2.085
r55 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.835 $X2=4.48 $Y2=2.91
r56 2 27 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.835 $X2=4.48 $Y2=2.21
r57 1 25 400 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.835 $X2=3.62 $Y2=2.21
r58 1 12 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.835 $X2=3.62 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%VGND 1 2 3 4 5 16 18 22 26 28 30 32 34 42
+ 47 52 61 73 77
r78 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r79 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r80 66 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r81 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r82 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 56 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r84 56 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r85 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r86 53 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=0 $X2=4.48
+ $Y2=0
r87 53 55 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=0 $X2=5.04
+ $Y2=0
r88 52 76 4.49945 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.467
+ $Y2=0
r89 52 55 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.04
+ $Y2=0
r90 51 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r91 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r92 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r93 48 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=4.08
+ $Y2=0
r94 47 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.48
+ $Y2=0
r95 47 50 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.08
+ $Y2=0
r96 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r97 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r98 43 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.155
+ $Y2=0
r99 43 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.64
+ $Y2=0
r100 42 70 6.34682 $w=8.63e-07 $l=4.5e-07 $layer=LI1_cond $X=3.352 $Y=0
+ $X2=3.352 $Y2=0.45
r101 42 48 10.735 $w=1.7e-07 $l=4.33e-07 $layer=LI1_cond $X=3.352 $Y=0 $X2=3.785
+ $Y2=0
r102 42 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r103 42 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r104 42 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.64
+ $Y2=0
r105 41 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r106 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r107 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r108 38 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r109 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r110 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r111 35 58 4.42547 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.202 $Y2=0
r112 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.72 $Y2=0
r113 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=0 $X2=2.155
+ $Y2=0
r114 34 40 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.99 $Y=0 $X2=1.68
+ $Y2=0
r115 32 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r116 32 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r117 28 76 3.26672 $w=3.3e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.467 $Y2=0
r118 28 30 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0.47
r119 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0
r120 24 26 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0.45
r121 20 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0
r122 20 22 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0.45
r123 16 58 3.05205 $w=2.95e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.202 $Y2=0
r124 16 18 15.0404 $w=2.93e-07 $l=3.85e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.47
r125 5 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.2
+ $Y=0.325 $X2=5.34 $Y2=0.47
r126 4 26 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.34
+ $Y=0.325 $X2=4.48 $Y2=0.45
r127 3 70 45.5 $w=1.7e-07 $l=8.05078e-07 $layer=licon1_NDIFF $count=4 $X=2.875
+ $Y=0.325 $X2=3.62 $Y2=0.45
r128 2 22 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=1.935
+ $Y=0.325 $X2=2.155 $Y2=0.45
r129 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.325 $X2=0.275 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_2%A_113_65# 1 2 9 11 12 15
c24 11 0 6.78225e-20 $X=1.47 $Y=0.35
r25 13 15 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.645 $Y=0.435
+ $X2=1.645 $Y2=0.45
r26 11 13 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=1.47 $Y=0.35
+ $X2=1.645 $Y2=0.435
r27 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=0.35 $X2=0.8
+ $Y2=0.35
r28 7 12 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.687 $Y=0.435
+ $X2=0.8 $Y2=0.35
r29 7 9 1.79269 $w=2.23e-07 $l=3.5e-08 $layer=LI1_cond $X=0.687 $Y=0.435
+ $X2=0.687 $Y2=0.47
r30 2 15 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=1.425
+ $Y=0.325 $X2=1.645 $Y2=0.45
r31 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.325 $X2=0.705 $Y2=0.47
.ends

