* NGSPICE file created from sky130_fd_sc_lp__bufbuf_16.ext - technology: sky130A

.subckt sky130_fd_sc_lp__bufbuf_16 A VGND VNB VPB VPWR X
M1000 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.8224e+12p pd=2.464e+07u as=4.9014e+12p ps=4.306e+07u
M1001 VPWR a_27_49# a_196_49# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=6.867e+11p ps=6.13e+06u
M1002 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=1.8816e+12p pd=1.792e+07u as=3.2676e+12p ps=3.13e+07u
M1003 a_610_47# a_196_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0584e+12p pd=9.24e+06u as=0p ps=0u
M1004 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_196_49# a_610_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.72e+06u
M1009 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_196_49# a_610_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A a_27_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1019 a_610_47# a_196_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_196_49# a_27_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_610_47# a_196_49# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_196_49# a_610_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_196_49# a_27_49# VGND VNB nshort w=840000u l=150000u
+  ad=4.578e+11p pd=4.45e+06u as=0p ps=0u
M1028 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_610_47# a_196_49# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_196_49# a_27_49# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_610_47# a_196_49# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_196_49# a_610_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_196_49# a_27_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_610_47# a_196_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_196_49# a_610_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR a_196_49# a_610_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VGND a_610_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 X a_610_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VGND a_27_49# a_196_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 X a_610_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VPWR a_610_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VPWR A a_27_49# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

