* File: sky130_fd_sc_lp__clkbuf_8.spice
* Created: Wed Sep  2 09:38:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkbuf_8.pex.spice"
.subckt sky130_fd_sc_lp__clkbuf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_A_110_47#_M1005_d N_A_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75004.1
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_110_47#_M1005_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75003.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1011_s N_A_110_47#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75003.2
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_110_47#_M1008_g N_X_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1008_d N_A_110_47#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_110_47#_M1010_g N_X_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1010_d N_A_110_47#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_110_47#_M1015_g N_X_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1015_d N_A_110_47#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_110_47#_M1019_g N_X_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0588 PD=1.38 PS=0.7 NRD=1.428 NRS=0 M=1 R=2.8 SA=75004.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_110_47#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g N_A_110_47#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1000 N_X_M1000_d N_A_110_47#_M1000_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1001 N_X_M1000_d N_A_110_47#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1002 N_X_M1002_d N_A_110_47#_M1002_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1004 N_X_M1002_d N_A_110_47#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_X_M1007_d N_A_110_47#_M1007_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1012 N_X_M1007_d N_A_110_47#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_X_M1013_d N_A_110_47#_M1013_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_X_M1013_d N_A_110_47#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.5559 P=15.05
*
.include "sky130_fd_sc_lp__clkbuf_8.pxi.spice"
*
.ends
*
*
