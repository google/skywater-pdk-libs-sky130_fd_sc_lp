* File: sky130_fd_sc_lp__or4_lp.pex.spice
* Created: Wed Sep  2 10:32:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4_LP%D 1 3 7 10 12 14 16 17 18 19 22 23 24
r52 22 24 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.37
+ $X2=0.595 $Y2=1.205
r53 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.37 $X2=0.605 $Y2=1.37
r54 19 23 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.635 $Y=1.665
+ $X2=0.635 $Y2=1.37
r55 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=0.855 $Y2=0.445
r56 13 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=0.805
+ $X2=0.495 $Y2=0.805
r57 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.855 $Y2=0.73
r58 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.57 $Y2=0.805
r59 10 18 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.645 $Y=2.595
+ $X2=0.645 $Y2=1.875
r60 7 18 33.6482 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.7
+ $X2=0.595 $Y2=1.875
r61 6 22 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.595 $Y=1.38 $X2=0.595
+ $Y2=1.37
r62 6 7 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.595 $Y=1.38
+ $X2=0.595 $Y2=1.7
r63 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=0.805
r64 4 24 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=1.205
r65 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.805
r66 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.73 $X2=0.495
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_LP%C 3 7 9 10 12 14 16 17 18 19 20 21 22 23 29
+ 30
r68 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.175
+ $Y=1.43 $X2=1.175 $Y2=1.43
r69 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=2.405
+ $X2=1.175 $Y2=2.775
r70 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=2.035
+ $X2=1.175 $Y2=2.405
r71 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.665
+ $X2=1.175 $Y2=2.035
r72 20 30 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.175 $Y=1.665
+ $X2=1.175 $Y2=1.43
r73 17 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.175 $Y=1.77
+ $X2=1.175 $Y2=1.43
r74 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.77
+ $X2=1.175 $Y2=1.935
r75 16 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.265
+ $X2=1.175 $Y2=1.43
r76 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.645 $Y=0.73
+ $X2=1.645 $Y2=0.445
r77 11 19 5.30422 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.36 $Y=0.805
+ $X2=1.275 $Y2=0.805
r78 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.57 $Y=0.805
+ $X2=1.645 $Y2=0.73
r79 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.57 $Y=0.805
+ $X2=1.36 $Y2=0.805
r80 7 19 20.4101 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=1.285 $Y=0.73
+ $X2=1.275 $Y2=0.805
r81 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.285 $Y=0.73 $X2=1.285
+ $Y2=0.445
r82 5 19 20.4101 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=1.265 $Y=0.88
+ $X2=1.275 $Y2=0.805
r83 5 16 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.265 $Y=0.88
+ $X2=1.265 $Y2=1.265
r84 3 18 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.135 $Y=2.595
+ $X2=1.135 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_LP%B 3 5 9 11 15 17 18 19 20 30 34
r49 33 35 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=1.77
+ $X2=1.745 $Y2=1.935
r50 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.745
+ $Y=1.77 $X2=1.745 $Y2=1.77
r51 30 33 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.745 $Y=1.68
+ $X2=1.745 $Y2=1.77
r52 19 20 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.405
+ $X2=1.92 $Y2=2.775
r53 18 19 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.92 $Y2=2.405
r54 18 34 4.46424 $w=7.08e-07 $l=2.65e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.92 $Y2=1.77
r55 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.725 $Y=1.605
+ $X2=2.725 $Y2=1.045
r56 12 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.325 $Y=1.68
+ $X2=2.25 $Y2=1.68
r57 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.65 $Y=1.68
+ $X2=2.725 $Y2=1.605
r58 11 12 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.65 $Y=1.68
+ $X2=2.325 $Y2=1.68
r59 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=1.605
+ $X2=2.25 $Y2=1.68
r60 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.25 $Y=1.605 $X2=2.25
+ $Y2=1.135
r61 6 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.68
+ $X2=1.745 $Y2=1.68
r62 5 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.175 $Y=1.68
+ $X2=2.25 $Y2=1.68
r63 5 6 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.175 $Y=1.68
+ $X2=1.91 $Y2=1.68
r64 3 35 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.705 $Y=2.595
+ $X2=1.705 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_LP%A 3 7 11 13 14 15 28 29
c45 29 0 5.86521e-20 $X=3.205 $Y=1.77
r46 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.77 $X2=3.205 $Y2=1.77
r47 26 28 7.47287 $w=2.58e-07 $l=4e-08 $layer=POLY_cond $X=3.165 $Y=1.77
+ $X2=3.205 $Y2=1.77
r48 25 26 1.86822 $w=2.58e-07 $l=1e-08 $layer=POLY_cond $X=3.155 $Y=1.77
+ $X2=3.165 $Y2=1.77
r49 14 15 5.23727 $w=8.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.947 $Y=2.405
+ $X2=2.947 $Y2=2.775
r50 13 14 5.23727 $w=8.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.947 $Y=2.035
+ $X2=2.947 $Y2=2.405
r51 13 29 3.75102 $w=8.43e-07 $l=2.65e-07 $layer=LI1_cond $X=2.947 $Y=2.035
+ $X2=2.947 $Y2=1.77
r52 9 28 57.9147 $w=2.58e-07 $l=3.83732e-07 $layer=POLY_cond $X=3.515 $Y=1.605
+ $X2=3.205 $Y2=1.77
r53 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.515 $Y=1.605
+ $X2=3.515 $Y2=1.045
r54 5 25 15.449 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=1.605
+ $X2=3.155 $Y2=1.77
r55 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.155 $Y=1.605
+ $X2=3.155 $Y2=1.045
r56 1 26 3.5867 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.935
+ $X2=3.165 $Y2=1.77
r57 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.165 $Y=1.935
+ $X2=3.165 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_LP%A_27_47# 1 2 3 4 15 17 19 20 22 24 29 32 34
+ 35 36 39 41 44 47 49 50 54 56 57 58 68
c133 68 0 1.22683e-19 $X=4.305 $Y=1.53
r134 64 66 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.945 $Y=1.53
+ $X2=3.98 $Y2=1.53
r135 62 68 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=4.01 $Y=1.53
+ $X2=4.305 $Y2=1.53
r136 62 66 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.01 $Y=1.53 $X2=3.98
+ $Y2=1.53
r137 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.53 $X2=4.01 $Y2=1.53
r138 58 61 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.01 $Y=1.41
+ $X2=4.01 $Y2=1.53
r139 51 54 9.4163 $w=4.08e-07 $l=3.35e-07 $layer=LI1_cond $X=1.605 $Y=0.47
+ $X2=1.94 $Y2=0.47
r140 49 50 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.317 $Y=2.24
+ $X2=0.317 $Y2=2.075
r141 44 46 9.79758 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=0.267 $Y=0.47
+ $X2=0.267 $Y2=0.675
r142 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=1.41
+ $X2=2.94 $Y2=1.41
r143 41 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=1.41
+ $X2=4.01 $Y2=1.41
r144 41 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.845 $Y=1.41
+ $X2=3.105 $Y2=1.41
r145 37 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=1.325
+ $X2=2.94 $Y2=1.41
r146 37 39 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.94 $Y=1.325
+ $X2=2.94 $Y2=1.045
r147 35 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=1.41
+ $X2=2.94 $Y2=1.41
r148 35 36 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=2.775 $Y=1.41
+ $X2=1.69 $Y2=1.41
r149 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.605 $Y=1.325
+ $X2=1.69 $Y2=1.41
r150 33 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.025
+ $X2=1.605 $Y2=0.94
r151 33 34 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.605 $Y=1.025
+ $X2=1.605 $Y2=1.325
r152 32 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.855
+ $X2=1.605 $Y2=0.94
r153 31 51 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.605 $Y=0.675
+ $X2=1.605 $Y2=0.47
r154 31 32 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.605 $Y=0.675
+ $X2=1.605 $Y2=0.855
r155 30 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.94
+ $X2=0.175 $Y2=0.94
r156 29 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.94
+ $X2=1.605 $Y2=0.94
r157 29 30 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.52 $Y=0.94
+ $X2=0.26 $Y2=0.94
r158 25 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=1.025
+ $X2=0.175 $Y2=0.94
r159 25 50 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=0.175 $Y=1.025
+ $X2=0.175 $Y2=2.075
r160 24 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=0.855
+ $X2=0.175 $Y2=0.94
r161 24 46 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.175 $Y=0.855
+ $X2=0.175 $Y2=0.675
r162 20 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.365
+ $X2=4.305 $Y2=1.53
r163 20 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.305 $Y=1.365
+ $X2=4.305 $Y2=1.045
r164 17 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.365
+ $X2=3.945 $Y2=1.53
r165 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.945 $Y=1.365
+ $X2=3.945 $Y2=1.045
r166 13 66 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.695
+ $X2=3.98 $Y2=1.53
r167 13 15 223.608 $w=2.5e-07 $l=9e-07 $layer=POLY_cond $X=3.98 $Y=1.695
+ $X2=3.98 $Y2=2.595
r168 4 49 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.235
+ $Y=2.095 $X2=0.38 $Y2=2.24
r169 3 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.835 $X2=2.94 $Y2=1.045
r170 2 54 182 $w=1.7e-07 $l=3.26994e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.235 $X2=1.94 $Y2=0.47
r171 1 44 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_LP%VPWR 1 6 10 12 19 20 23
c39 6 0 6.40308e-20 $X=3.715 $Y=2.24
r40 23 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r41 20 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r43 17 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=3.715 $Y2=3.33
r44 17 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r45 14 15 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 12 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=3.715 $Y2=3.33
r47 12 14 215.947 $w=1.68e-07 $l=3.31e-06 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 10 24 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 10 15 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 6 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.715 $Y=2.24 $X2=3.715
+ $Y2=2.95
r51 4 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=3.245
+ $X2=3.715 $Y2=3.33
r52 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.715 $Y=3.245
+ $X2=3.715 $Y2=2.95
r53 1 9 400 $w=1.7e-07 $l=1.04614e-06 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=2.095 $X2=3.715 $Y2=2.95
r54 1 6 400 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=2.095 $X2=3.715 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_LP%X 1 2 7 8 9 10 11 12 13 36
r18 22 36 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=4.52 $Y=2.075 $X2=4.52
+ $Y2=2.035
r19 12 13 8.1187 $w=5.56e-07 $l=3.7e-07 $layer=LI1_cond $X=4.382 $Y=2.405
+ $X2=4.382 $Y2=2.775
r20 12 39 3.6205 $w=5.56e-07 $l=1.65e-07 $layer=LI1_cond $X=4.382 $Y=2.405
+ $X2=4.382 $Y2=2.24
r21 11 39 3.13777 $w=5.56e-07 $l=1.43e-07 $layer=LI1_cond $X=4.382 $Y=2.097
+ $X2=4.382 $Y2=2.24
r22 11 22 2.48216 $w=5.56e-07 $l=1.48593e-07 $layer=LI1_cond $X=4.382 $Y=2.097
+ $X2=4.52 $Y2=2.075
r23 11 36 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=4.52 $Y=2.012
+ $X2=4.52 $Y2=2.035
r24 10 11 12.1181 $w=3.28e-07 $l=3.47e-07 $layer=LI1_cond $X=4.52 $Y=1.665
+ $X2=4.52 $Y2=2.012
r25 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=1.295
+ $X2=4.52 $Y2=1.665
r26 9 29 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.52 $Y=1.295
+ $X2=4.52 $Y2=1.045
r27 8 29 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.52 $Y=0.925 $X2=4.52
+ $Y2=1.045
r28 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=0.555 $X2=4.52
+ $Y2=0.925
r29 2 39 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.105
+ $Y=2.095 $X2=4.245 $Y2=2.24
r30 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.835 $X2=4.52 $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_LP%VGND 1 2 3 12 14 19 22 25 26 27 29 38 44 45
+ 48 51
r82 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r83 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r84 45 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r85 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r86 42 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=3.73
+ $Y2=0
r87 42 44 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.56
+ $Y2=0
r88 41 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r89 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r90 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=0 $X2=3.73
+ $Y2=0
r91 38 40 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.565 $Y=0 $X2=2.64
+ $Y2=0
r92 37 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r93 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r94 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r95 34 36 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=2.16
+ $Y2=0
r96 32 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r97 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r98 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r99 29 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r100 27 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r101 27 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r102 25 36 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=0
+ $X2=2.16 $Y2=0
r103 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.37
+ $Y2=0
r104 24 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.455 $Y=0
+ $X2=2.64 $Y2=0
r105 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.37
+ $Y2=0
r106 20 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0
r107 20 22 31.2557 $w=3.28e-07 $l=8.95e-07 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0.98
r108 18 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=0.085
+ $X2=2.37 $Y2=0
r109 18 19 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.37 $Y=0.085
+ $X2=2.37 $Y2=0.895
r110 14 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.285 $Y=1.02
+ $X2=2.37 $Y2=0.895
r111 14 16 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.285 $Y=1.02
+ $X2=2.035 $Y2=1.02
r112 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r113 10 12 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.445
r114 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.835 $X2=3.73 $Y2=0.98
r115 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.925 $X2=2.035 $Y2=1.06
r116 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.445
.ends

