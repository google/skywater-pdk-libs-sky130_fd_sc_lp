* NGSPICE file created from sky130_fd_sc_lp__clkbuflp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__clkbuflp_2 A VGND VNB VPB VPWR X
M1000 VGND A a_110_47# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR A a_27_47# VPB phighvt w=1e+06u l=250000u
+  ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u
M1002 VPWR a_27_47# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1003 a_110_47# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 X a_27_47# a_268_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_268_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_426_47# a_27_47# X VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 VGND a_27_47# a_426_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_27_47# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

