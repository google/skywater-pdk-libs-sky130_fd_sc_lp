* File: sky130_fd_sc_lp__a211o_1.pxi.spice
* Created: Fri Aug 28 09:47:25 2020
* 
x_PM_SKY130_FD_SC_LP__A211O_1%A_80_237# N_A_80_237#_M1001_d N_A_80_237#_M1007_d
+ N_A_80_237#_M1000_d N_A_80_237#_M1008_g N_A_80_237#_c_53_n N_A_80_237#_M1009_g
+ N_A_80_237#_c_54_n N_A_80_237#_c_55_n N_A_80_237#_c_65_p N_A_80_237#_c_120_p
+ N_A_80_237#_c_60_n N_A_80_237#_c_61_n N_A_80_237#_c_123_p N_A_80_237#_c_56_n
+ N_A_80_237#_c_62_n N_A_80_237#_c_57_n N_A_80_237#_c_78_p
+ PM_SKY130_FD_SC_LP__A211O_1%A_80_237#
x_PM_SKY130_FD_SC_LP__A211O_1%A2 N_A2_c_139_n N_A2_M1002_g N_A2_c_140_n
+ N_A2_M1003_g A2 N_A2_c_142_n PM_SKY130_FD_SC_LP__A211O_1%A2
x_PM_SKY130_FD_SC_LP__A211O_1%A1 N_A1_M1001_g N_A1_M1004_g A1 N_A1_c_172_n
+ N_A1_c_173_n N_A1_c_174_n PM_SKY130_FD_SC_LP__A211O_1%A1
x_PM_SKY130_FD_SC_LP__A211O_1%B1 N_B1_M1006_g N_B1_M1005_g B1 N_B1_c_204_n
+ N_B1_c_205_n PM_SKY130_FD_SC_LP__A211O_1%B1
x_PM_SKY130_FD_SC_LP__A211O_1%C1 N_C1_c_231_n N_C1_M1007_g N_C1_M1000_g C1
+ N_C1_c_234_n PM_SKY130_FD_SC_LP__A211O_1%C1
x_PM_SKY130_FD_SC_LP__A211O_1%X N_X_M1009_s N_X_M1008_s X X X X X X X
+ N_X_c_254_n PM_SKY130_FD_SC_LP__A211O_1%X
x_PM_SKY130_FD_SC_LP__A211O_1%VPWR N_VPWR_M1008_d N_VPWR_M1003_d N_VPWR_c_269_n
+ N_VPWR_c_270_n VPWR N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n
+ N_VPWR_c_268_n N_VPWR_c_275_n N_VPWR_c_276_n PM_SKY130_FD_SC_LP__A211O_1%VPWR
x_PM_SKY130_FD_SC_LP__A211O_1%A_217_367# N_A_217_367#_M1003_s
+ N_A_217_367#_M1004_d N_A_217_367#_c_312_n N_A_217_367#_c_313_n
+ N_A_217_367#_c_317_n N_A_217_367#_c_318_n N_A_217_367#_c_330_n
+ PM_SKY130_FD_SC_LP__A211O_1%A_217_367#
x_PM_SKY130_FD_SC_LP__A211O_1%VGND N_VGND_M1009_d N_VGND_M1006_d N_VGND_c_334_n
+ VGND N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n
+ N_VGND_c_339_n N_VGND_c_340_n PM_SKY130_FD_SC_LP__A211O_1%VGND
cc_1 VNB N_A_80_237#_M1008_g 0.00916818f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_A_80_237#_c_53_n 0.0223136f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.185
cc_3 VNB N_A_80_237#_c_54_n 0.00399475f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.35
cc_4 VNB N_A_80_237#_c_55_n 0.0555507f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.35
cc_5 VNB N_A_80_237#_c_56_n 0.00750854f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=0.94
cc_6 VNB N_A_80_237#_c_57_n 0.0232127f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.42
cc_7 VNB N_A2_c_139_n 0.0194062f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.235
cc_8 VNB N_A2_c_140_n 0.0318015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_M1003_g 0.00837672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_142_n 0.00302018f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_11 VNB N_A1_M1004_g 0.00825767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_c_172_n 0.0286403f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_13 VNB N_A1_c_173_n 0.00842565f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_14 VNB N_A1_c_174_n 0.0174643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1005_g 0.00779945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB B1 0.00851237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_204_n 0.0282606f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_18 VNB N_B1_c_205_n 0.0185525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C1_c_231_n 0.0230209f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.235
cc_20 VNB N_C1_M1000_g 0.0112001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB C1 0.00309203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C1_c_234_n 0.0539447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_254_n 0.0580557f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.94
cc_24 VNB N_VPWR_c_268_n 0.143779f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=2.91
cc_25 VNB N_VGND_c_334_n 0.00561478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_335_n 0.0308022f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.695
cc_27 VNB N_VGND_c_336_n 0.0179557f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.78
cc_28 VNB N_VGND_c_337_n 0.189715f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=0.855
cc_29 VNB N_VGND_c_338_n 0.0164907f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=0.94
cc_30 VNB N_VGND_c_339_n 0.0149858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_340_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.42
cc_32 VPB N_A_80_237#_M1008_g 0.0277639f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_33 VPB N_A_80_237#_c_54_n 7.43006e-19 $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.35
cc_34 VPB N_A_80_237#_c_60_n 0.0300651f $X=-0.19 $Y=1.655 $X2=2.915 $Y2=1.78
cc_35 VPB N_A_80_237#_c_61_n 0.00546974f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.78
cc_36 VPB N_A_80_237#_c_62_n 0.0470856f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.98
cc_37 VPB N_A2_M1003_g 0.0247846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A1_M1004_g 0.0207025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_B1_M1005_g 0.0196641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_C1_M1000_g 0.0245806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_X_c_254_n 0.0554157f $X=-0.19 $Y=1.655 $X2=1.905 $Y2=0.94
cc_42 VPB N_VPWR_c_269_n 0.0144541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_270_n 0.0050746f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.655
cc_44 VPB N_VPWR_c_271_n 0.0174123f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.35
cc_45 VPB N_VPWR_c_272_n 0.0181354f $X=-0.19 $Y=1.655 $X2=2.915 $Y2=1.78
cc_46 VPB N_VPWR_c_273_n 0.0440547f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.98
cc_47 VPB N_VPWR_c_268_n 0.0537813f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=2.91
cc_48 VPB N_VPWR_c_275_n 0.00535651f $X=-0.19 $Y=1.655 $X2=3.095 $Y2=0.855
cc_49 VPB N_VPWR_c_276_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_217_367#_c_312_n 0.00195979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_217_367#_c_313_n 0.00803344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 N_A_80_237#_c_54_n N_A2_c_139_n 0.00466704f $X=0.75 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_53 N_A_80_237#_c_55_n N_A2_c_139_n 3.28199e-19 $X=0.75 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_54 N_A_80_237#_c_65_p N_A2_c_139_n 0.014749f $X=1.905 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_55 N_A_80_237#_c_54_n N_A2_c_140_n 3.92978e-19 $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_56 N_A_80_237#_c_55_n N_A2_c_140_n 0.0189439f $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_57 N_A_80_237#_c_65_p N_A2_c_140_n 0.00391065f $X=1.905 $Y=0.94 $X2=0 $Y2=0
cc_58 N_A_80_237#_c_60_n N_A2_c_140_n 0.00482651f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_59 N_A_80_237#_c_54_n N_A2_M1003_g 0.00473994f $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_60 N_A_80_237#_c_60_n N_A2_M1003_g 0.0143976f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_61 N_A_80_237#_c_54_n N_A2_c_142_n 0.0259612f $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_80_237#_c_55_n N_A2_c_142_n 0.00195965f $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_63 N_A_80_237#_c_65_p N_A2_c_142_n 0.020507f $X=1.905 $Y=0.94 $X2=0 $Y2=0
cc_64 N_A_80_237#_c_60_n N_A2_c_142_n 0.0230001f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_65 N_A_80_237#_c_60_n N_A1_M1004_g 0.0112552f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_66 N_A_80_237#_c_60_n N_A1_c_172_n 0.00122069f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_67 N_A_80_237#_c_78_p N_A1_c_172_n 0.00359541f $X=2.07 $Y=0.94 $X2=0 $Y2=0
cc_68 N_A_80_237#_c_65_p N_A1_c_173_n 0.0205542f $X=1.905 $Y=0.94 $X2=0 $Y2=0
cc_69 N_A_80_237#_c_60_n N_A1_c_173_n 0.036737f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_70 N_A_80_237#_c_78_p N_A1_c_173_n 0.00990255f $X=2.07 $Y=0.94 $X2=0 $Y2=0
cc_71 N_A_80_237#_c_65_p N_A1_c_174_n 0.0125368f $X=1.905 $Y=0.94 $X2=0 $Y2=0
cc_72 N_A_80_237#_c_60_n N_B1_M1005_g 0.0153485f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_73 N_A_80_237#_c_62_n N_B1_M1005_g 0.00391071f $X=3.08 $Y=1.98 $X2=0 $Y2=0
cc_74 N_A_80_237#_c_60_n B1 0.037132f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_75 N_A_80_237#_c_56_n B1 0.0306669f $X=2.945 $Y=0.94 $X2=0 $Y2=0
cc_76 N_A_80_237#_c_60_n N_B1_c_204_n 0.00122615f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_77 N_A_80_237#_c_56_n N_B1_c_204_n 0.00365043f $X=2.945 $Y=0.94 $X2=0 $Y2=0
cc_78 N_A_80_237#_c_56_n N_B1_c_205_n 0.0132146f $X=2.945 $Y=0.94 $X2=0 $Y2=0
cc_79 N_A_80_237#_c_56_n N_C1_c_231_n 0.0121429f $X=2.945 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_80_237#_c_60_n N_C1_M1000_g 0.01632f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_81 N_A_80_237#_c_62_n N_C1_M1000_g 0.0248121f $X=3.08 $Y=1.98 $X2=0 $Y2=0
cc_82 N_A_80_237#_c_60_n C1 0.0286458f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_83 N_A_80_237#_c_56_n C1 0.0226511f $X=2.945 $Y=0.94 $X2=0 $Y2=0
cc_84 N_A_80_237#_c_60_n N_C1_c_234_n 0.00226177f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_85 N_A_80_237#_c_56_n N_C1_c_234_n 0.00673878f $X=2.945 $Y=0.94 $X2=0 $Y2=0
cc_86 N_A_80_237#_M1008_g N_X_c_254_n 0.0288921f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_80_237#_c_53_n N_X_c_254_n 0.00486661f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_88 N_A_80_237#_c_54_n N_X_c_254_n 0.0470269f $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_89 N_A_80_237#_c_55_n N_X_c_254_n 0.0115619f $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_80_237#_c_61_n N_X_c_254_n 0.012284f $X=0.915 $Y=1.78 $X2=0 $Y2=0
cc_91 N_A_80_237#_c_61_n N_VPWR_M1008_d 0.00270358f $X=0.915 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_80_237#_c_60_n N_VPWR_M1003_d 0.0026214f $X=2.915 $Y=1.78 $X2=0 $Y2=0
cc_93 N_A_80_237#_M1008_g N_VPWR_c_269_n 0.00477918f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_A_80_237#_c_55_n N_VPWR_c_269_n 9.88813e-19 $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_95 N_A_80_237#_c_61_n N_VPWR_c_269_n 0.0214721f $X=0.915 $Y=1.78 $X2=0 $Y2=0
cc_96 N_A_80_237#_M1008_g N_VPWR_c_271_n 0.00579312f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_97 N_A_80_237#_c_62_n N_VPWR_c_273_n 0.0210467f $X=3.08 $Y=1.98 $X2=0 $Y2=0
cc_98 N_A_80_237#_M1000_d N_VPWR_c_268_n 0.00215158f $X=2.94 $Y=1.835 $X2=0
+ $Y2=0
cc_99 N_A_80_237#_M1008_g N_VPWR_c_268_n 0.0126572f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_100 N_A_80_237#_c_62_n N_VPWR_c_268_n 0.0125689f $X=3.08 $Y=1.98 $X2=0 $Y2=0
cc_101 N_A_80_237#_c_60_n N_A_217_367#_M1003_s 0.00234752f $X=2.915 $Y=1.78
+ $X2=-0.19 $Y2=-0.245
cc_102 N_A_80_237#_c_60_n N_A_217_367#_M1004_d 0.00261503f $X=2.915 $Y=1.78
+ $X2=0 $Y2=0
cc_103 N_A_80_237#_c_60_n N_A_217_367#_c_312_n 0.020301f $X=2.915 $Y=1.78 $X2=0
+ $Y2=0
cc_104 N_A_80_237#_c_60_n N_A_217_367#_c_317_n 0.0381341f $X=2.915 $Y=1.78 $X2=0
+ $Y2=0
cc_105 N_A_80_237#_c_60_n N_A_217_367#_c_318_n 0.0200142f $X=2.915 $Y=1.78 $X2=0
+ $Y2=0
cc_106 N_A_80_237#_c_60_n A_504_367# 0.00595227f $X=2.915 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_80_237#_c_54_n N_VGND_M1009_d 7.50871e-19 $X=0.75 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_108 N_A_80_237#_c_65_p N_VGND_M1009_d 0.0105286f $X=1.905 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_80_237#_c_120_p N_VGND_M1009_d 0.00413959f $X=0.915 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_80_237#_c_56_n N_VGND_M1006_d 0.00507283f $X=2.945 $Y=0.94 $X2=0
+ $Y2=0
cc_111 N_A_80_237#_c_56_n N_VGND_c_334_n 0.0196002f $X=2.945 $Y=0.94 $X2=0 $Y2=0
cc_112 N_A_80_237#_c_123_p N_VGND_c_335_n 0.0222962f $X=2.07 $Y=0.375 $X2=0
+ $Y2=0
cc_113 N_A_80_237#_c_57_n N_VGND_c_336_n 0.0192303f $X=3.08 $Y=0.42 $X2=0 $Y2=0
cc_114 N_A_80_237#_M1001_d N_VGND_c_337_n 0.00399873f $X=1.86 $Y=0.235 $X2=0
+ $Y2=0
cc_115 N_A_80_237#_M1007_d N_VGND_c_337_n 0.00211137f $X=2.94 $Y=0.235 $X2=0
+ $Y2=0
cc_116 N_A_80_237#_c_53_n N_VGND_c_337_n 0.00978457f $X=0.515 $Y=1.185 $X2=0
+ $Y2=0
cc_117 N_A_80_237#_c_65_p N_VGND_c_337_n 0.0184645f $X=1.905 $Y=0.94 $X2=0 $Y2=0
cc_118 N_A_80_237#_c_120_p N_VGND_c_337_n 0.00117642f $X=0.915 $Y=0.94 $X2=0
+ $Y2=0
cc_119 N_A_80_237#_c_123_p N_VGND_c_337_n 0.0127519f $X=2.07 $Y=0.375 $X2=0
+ $Y2=0
cc_120 N_A_80_237#_c_56_n N_VGND_c_337_n 0.0117491f $X=2.945 $Y=0.94 $X2=0 $Y2=0
cc_121 N_A_80_237#_c_57_n N_VGND_c_337_n 0.0115856f $X=3.08 $Y=0.42 $X2=0 $Y2=0
cc_122 N_A_80_237#_c_53_n N_VGND_c_338_n 0.00525069f $X=0.515 $Y=1.185 $X2=0
+ $Y2=0
cc_123 N_A_80_237#_c_53_n N_VGND_c_339_n 0.0147439f $X=0.515 $Y=1.185 $X2=0
+ $Y2=0
cc_124 N_A_80_237#_c_55_n N_VGND_c_339_n 0.00117978f $X=0.75 $Y=1.35 $X2=0 $Y2=0
cc_125 N_A_80_237#_c_65_p N_VGND_c_339_n 0.029374f $X=1.905 $Y=0.94 $X2=0 $Y2=0
cc_126 N_A_80_237#_c_120_p N_VGND_c_339_n 0.023869f $X=0.915 $Y=0.94 $X2=0 $Y2=0
cc_127 N_A_80_237#_c_65_p A_294_47# 0.00425358f $X=1.905 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A2_c_140_n N_A1_M1004_g 0.0344703f $X=1.425 $Y=1.525 $X2=0 $Y2=0
cc_129 N_A2_c_140_n N_A1_c_172_n 0.0426567f $X=1.425 $Y=1.525 $X2=0 $Y2=0
cc_130 N_A2_c_142_n N_A1_c_172_n 3.39157e-19 $X=1.305 $Y=1.36 $X2=0 $Y2=0
cc_131 N_A2_c_140_n N_A1_c_173_n 0.00232902f $X=1.425 $Y=1.525 $X2=0 $Y2=0
cc_132 N_A2_c_142_n N_A1_c_173_n 0.0256327f $X=1.305 $Y=1.36 $X2=0 $Y2=0
cc_133 N_A2_c_139_n N_A1_c_174_n 0.0339574f $X=1.395 $Y=1.195 $X2=0 $Y2=0
cc_134 N_A2_M1003_g N_VPWR_c_269_n 0.00271044f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A2_M1003_g N_VPWR_c_270_n 0.00219364f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_M1003_g N_VPWR_c_272_n 0.00585385f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A2_M1003_g N_VPWR_c_268_n 0.0120419f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A2_M1003_g N_A_217_367#_c_317_n 0.0133747f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A2_c_139_n N_VGND_c_335_n 0.00486043f $X=1.395 $Y=1.195 $X2=0 $Y2=0
cc_140 N_A2_c_139_n N_VGND_c_337_n 0.00455001f $X=1.395 $Y=1.195 $X2=0 $Y2=0
cc_141 N_A2_c_139_n N_VGND_c_339_n 0.017921f $X=1.395 $Y=1.195 $X2=0 $Y2=0
cc_142 N_A1_M1004_g N_B1_M1005_g 0.0212379f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A1_c_172_n B1 3.8273e-19 $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_144 N_A1_c_173_n B1 0.0212768f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_145 N_A1_c_172_n N_B1_c_204_n 0.0216574f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_146 N_A1_c_173_n N_B1_c_204_n 3.82779e-19 $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_147 N_A1_c_174_n N_B1_c_205_n 0.0260728f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_VPWR_c_270_n 0.00361115f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A1_M1004_g N_VPWR_c_273_n 0.00585385f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A1_M1004_g N_VPWR_c_268_n 0.0109484f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A1_M1004_g N_A_217_367#_c_317_n 0.0133747f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A1_c_174_n N_VGND_c_335_n 0.00585385f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A1_c_174_n N_VGND_c_337_n 0.00684023f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_154 N_A1_c_174_n N_VGND_c_339_n 0.00250933f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_155 N_B1_c_205_n N_C1_c_231_n 0.0232095f $X=2.415 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_156 N_B1_M1005_g N_C1_M1000_g 0.0774782f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_157 B1 C1 0.0256318f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_158 N_B1_c_204_n C1 2.3766e-19 $X=2.415 $Y=1.35 $X2=0 $Y2=0
cc_159 B1 N_C1_c_234_n 0.00240641f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_160 N_B1_c_204_n N_C1_c_234_n 0.0211546f $X=2.415 $Y=1.35 $X2=0 $Y2=0
cc_161 N_B1_M1005_g N_VPWR_c_273_n 0.00585385f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_162 N_B1_M1005_g N_VPWR_c_268_n 0.0110801f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B1_c_205_n N_VGND_c_334_n 0.00400211f $X=2.415 $Y=1.185 $X2=0 $Y2=0
cc_164 N_B1_c_205_n N_VGND_c_335_n 0.00585385f $X=2.415 $Y=1.185 $X2=0 $Y2=0
cc_165 N_B1_c_205_n N_VGND_c_337_n 0.00691388f $X=2.415 $Y=1.185 $X2=0 $Y2=0
cc_166 N_C1_M1000_g N_VPWR_c_273_n 0.0054895f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_167 N_C1_M1000_g N_VPWR_c_268_n 0.0109725f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_168 N_C1_c_231_n N_VGND_c_334_n 0.00400211f $X=2.865 $Y=1.185 $X2=0 $Y2=0
cc_169 N_C1_c_231_n N_VGND_c_336_n 0.00585385f $X=2.865 $Y=1.185 $X2=0 $Y2=0
cc_170 N_C1_c_231_n N_VGND_c_337_n 0.00743588f $X=2.865 $Y=1.185 $X2=0 $Y2=0
cc_171 N_X_c_254_n N_VPWR_c_271_n 0.0196832f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_172 N_X_M1008_s N_VPWR_c_268_n 0.00215158f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_173 N_X_c_254_n N_VPWR_c_268_n 0.0118828f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_174 N_X_c_254_n N_A_217_367#_c_312_n 3.07662e-19 $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_175 N_X_M1009_s N_VGND_c_337_n 0.00336915f $X=0.175 $Y=0.235 $X2=0 $Y2=0
cc_176 N_X_c_254_n N_VGND_c_337_n 0.0119743f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_177 N_X_c_254_n N_VGND_c_338_n 0.0210334f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_178 N_VPWR_c_268_n N_A_217_367#_M1003_s 0.00232552f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_179 N_VPWR_c_268_n N_A_217_367#_M1004_d 0.00392255f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_269_n N_A_217_367#_c_312_n 0.0129305f $X=0.69 $Y=2.21 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_269_n N_A_217_367#_c_313_n 0.0656518f $X=0.69 $Y=2.21 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_272_n N_A_217_367#_c_313_n 0.0192303f $X=1.515 $Y=3.33 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_268_n N_A_217_367#_c_313_n 0.0115856f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_184 N_VPWR_M1003_d N_A_217_367#_c_317_n 0.00509967f $X=1.5 $Y=1.835 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_270_n N_A_217_367#_c_317_n 0.0200142f $X=1.68 $Y=2.5 $X2=0 $Y2=0
cc_186 N_VPWR_c_273_n N_A_217_367#_c_330_n 0.0202063f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_268_n N_A_217_367#_c_330_n 0.0127519f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_268_n A_504_367# 0.0115639f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_189 N_VGND_c_337_n A_294_47# 0.00357568f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
