* File: sky130_fd_sc_lp__a2bb2o_2.spice
* Created: Fri Aug 28 09:55:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2o_2.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2o_2  VNB VPB B1 B2 A2_N A1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1013 A_146_131# N_B1_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.3
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_218_131#_M1010_d N_B2_M1010_g A_146_131# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_260_341#_M1011_g N_A_218_131#_M1010_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.175925 AS=0.0588 PD=1.315 PS=0.7 NRD=103.956 NRS=0 M=1
+ R=2.8 SA=75001 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1006 N_A_260_341#_M1006_d N_A2_N_M1006_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.175925 PD=0.7 PS=1.315 NRD=0 NRS=103.956 M=1 R=2.8
+ SA=75001.8 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A1_N_M1007_g N_A_260_341#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0896 AS=0.0588 PD=0.81 PS=0.7 NRD=28.56 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_218_131#_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1012 N_X_M1004_d N_A_218_131#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.315 PD=1.12 PS=2.43 NRD=0 NRS=12.852 M=1 R=5.6 SA=75001.9
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_A_27_481#_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1024 AS=0.1696 PD=0.96 PS=1.81 NRD=6.1464 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 N_A_27_481#_M1008_d N_B2_M1008_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=6.1464 M=1 R=4.26667 SA=75000.7
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_218_131#_M1002_d N_A_260_341#_M1002_g N_A_27_481#_M1008_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 A_480_367# N_A2_N_M1005_g N_A_260_341#_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A1_N_M1009_g A_480_367# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.146964 AS=0.0672 PD=1.13516 PS=0.85 NRD=53.7416 NRS=15.3857 M=1 R=4.26667
+ SA=75000.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1009_d N_A_218_131#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.289336 AS=0.1764 PD=2.23484 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_218_131#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4725 AS=0.1764 PD=3.27 PS=1.54 NRD=14.0658 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.3 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a2bb2o_2.pxi.spice"
*
.ends
*
*
