* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand3_4 A B C VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_33_57# B a_460_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND C a_460_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_33_57# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_460_57# B a_33_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Y A a_33_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_460_57# B a_33_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_460_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VGND C a_460_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_33_57# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_460_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 Y A a_33_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_33_57# B a_460_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
