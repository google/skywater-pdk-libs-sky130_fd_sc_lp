* File: sky130_fd_sc_lp__o2bb2ai_1.spice
* Created: Wed Sep  2 10:22:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2ai_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1003 A_115_52# N_A1_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_115_367#_M1009_d N_A2_N_M1009_g A_115_52# VNB NSHORT L=0.15 W=0.84
+ AD=0.2856 AS=0.0882 PD=2.36 PS=1.05 NRD=10.704 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1004 N_A_396_47#_M1004_d N_A_115_367#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_B2_M1006_g N_A_396_47#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.1176 PD=1.22 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_A_396_47#_M1008_d N_B1_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1596 PD=2.21 PS=1.22 NRD=0 NRS=4.284 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_115_367#_M1005_d N_A1_N_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A2_N_M1007_g N_A_115_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.53865 AS=0.1764 PD=2.115 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_115_367#_M1001_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.53865 PD=1.62 PS=2.115 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1002 A_504_367# N_B2_M1002_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1701
+ AS=0.2268 PD=1.53 PS=1.62 NRD=12.4898 NRS=9.3772 M=1 R=8.4 SA=75002.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g A_504_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1701 PD=3.05 PS=1.53 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75002.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o2bb2ai_1.pxi.spice"
*
.ends
*
*
