* File: sky130_fd_sc_lp__maj3_2.pxi.spice
* Created: Fri Aug 28 10:43:01 2020
* 
x_PM_SKY130_FD_SC_LP__MAJ3_2%C N_C_M1008_g N_C_M1002_g N_C_M1011_g N_C_M1015_g
+ N_C_c_82_n N_C_c_89_n N_C_c_83_n N_C_c_84_n N_C_c_91_n C C N_C_c_93_n
+ N_C_c_94_n N_C_c_95_n C PM_SKY130_FD_SC_LP__MAJ3_2%C
x_PM_SKY130_FD_SC_LP__MAJ3_2%A N_A_M1009_g N_A_M1003_g N_A_M1000_g N_A_M1006_g
+ N_A_c_175_n N_A_c_176_n A A N_A_c_172_n PM_SKY130_FD_SC_LP__MAJ3_2%A
x_PM_SKY130_FD_SC_LP__MAJ3_2%B N_B_c_230_n N_B_M1010_g N_B_M1007_g N_B_M1004_g
+ N_B_M1014_g N_B_c_227_n B N_B_c_228_n N_B_c_229_n PM_SKY130_FD_SC_LP__MAJ3_2%B
x_PM_SKY130_FD_SC_LP__MAJ3_2%A_59_491# N_A_59_491#_M1002_s N_A_59_491#_M1007_d
+ N_A_59_491#_M1008_s N_A_59_491#_M1010_d N_A_59_491#_M1001_g
+ N_A_59_491#_M1005_g N_A_59_491#_M1012_g N_A_59_491#_M1013_g
+ N_A_59_491#_c_285_n N_A_59_491#_c_286_n N_A_59_491#_c_297_n
+ N_A_59_491#_c_287_n N_A_59_491#_c_288_n N_A_59_491#_c_317_n
+ N_A_59_491#_c_318_n N_A_59_491#_c_289_n N_A_59_491#_c_290_n
+ N_A_59_491#_c_298_n N_A_59_491#_c_291_n N_A_59_491#_c_292_n
+ N_A_59_491#_c_293_n PM_SKY130_FD_SC_LP__MAJ3_2%A_59_491#
x_PM_SKY130_FD_SC_LP__MAJ3_2%VPWR N_VPWR_M1009_d N_VPWR_M1011_d N_VPWR_M1013_d
+ N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n
+ N_VPWR_c_423_n VPWR N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n
+ N_VPWR_c_417_n PM_SKY130_FD_SC_LP__MAJ3_2%VPWR
x_PM_SKY130_FD_SC_LP__MAJ3_2%X N_X_M1001_d N_X_M1005_s N_X_c_483_n N_X_c_488_n
+ N_X_c_481_n X X N_X_c_489_n X PM_SKY130_FD_SC_LP__MAJ3_2%X
x_PM_SKY130_FD_SC_LP__MAJ3_2%VGND N_VGND_M1003_d N_VGND_M1015_d N_VGND_M1012_s
+ N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n N_VGND_c_522_n
+ N_VGND_c_523_n VGND N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n
+ N_VGND_c_527_n PM_SKY130_FD_SC_LP__MAJ3_2%VGND
cc_1 VNB N_C_M1002_g 0.0485366f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.455
cc_2 VNB N_C_M1015_g 0.0631207f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.455
cc_3 VNB N_C_c_82_n 0.0172986f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.77
cc_4 VNB N_C_c_83_n 0.00187656f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_5 VNB N_C_c_84_n 0.0178514f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_6 VNB N_A_M1003_g 0.0364539f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.455
cc_7 VNB N_A_M1006_g 0.0364539f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_8 VNB A 0.00495415f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_9 VNB N_A_c_172_n 0.0431779f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=2.15
cc_10 VNB N_B_M1007_g 0.0359094f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.455
cc_11 VNB N_B_M1014_g 0.0358876f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.455
cc_12 VNB N_B_c_227_n 0.019703f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_13 VNB N_B_c_228_n 0.0279441f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=2.15
cc_14 VNB N_B_c_229_n 9.55467e-19 $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.15
cc_15 VNB N_A_59_491#_M1001_g 0.0219059f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.455
cc_16 VNB N_A_59_491#_M1005_g 0.00234668f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.77
cc_17 VNB N_A_59_491#_M1012_g 0.0254753f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_18 VNB N_A_59_491#_M1013_g 0.0167082f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.15
cc_19 VNB N_A_59_491#_c_285_n 0.0306178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_59_491#_c_286_n 0.0244471f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_21 VNB N_A_59_491#_c_287_n 0.0327739f $X=-0.19 $Y=-0.245 $X2=2.745 $Y2=1.905
cc_22 VNB N_A_59_491#_c_288_n 0.0255986f $X=-0.19 $Y=-0.245 $X2=2.745 $Y2=2.235
cc_23 VNB N_A_59_491#_c_289_n 0.0212968f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=2.035
cc_24 VNB N_A_59_491#_c_290_n 0.00410597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_59_491#_c_291_n 0.00233723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_59_491#_c_292_n 0.00546493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_59_491#_c_293_n 0.0610246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_417_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_481_n 0.00792293f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.455
cc_30 VNB X 0.0057241f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.95
cc_31 VNB N_VGND_c_518_n 0.00322653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_519_n 0.00418963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_520_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.265
cc_34 VNB N_VGND_c_521_n 0.0475212f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.935
cc_35 VNB N_VGND_c_522_n 0.0366353f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_36 VNB N_VGND_c_523_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.43
cc_37 VNB N_VGND_c_524_n 0.0342543f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.15
cc_38 VNB N_VGND_c_525_n 0.0224829f $X=-0.19 $Y=-0.245 $X2=2.69 $Y2=2.07
cc_39 VNB N_VGND_c_526_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=2.622 $Y2=2.07
cc_40 VNB N_VGND_c_527_n 0.237655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_C_M1008_g 0.0429679f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.775
cc_42 VPB N_C_M1011_g 0.0245518f $X=-0.19 $Y=1.655 $X2=2.685 $Y2=2.775
cc_43 VPB N_C_M1015_g 0.0154343f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=0.455
cc_44 VPB N_C_c_82_n 0.00880373f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.77
cc_45 VPB N_C_c_89_n 0.01781f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.935
cc_46 VPB N_C_c_83_n 0.0026386f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.43
cc_47 VPB N_C_c_91_n 0.00335145f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.15
cc_48 VPB C 0.00413871f $X=-0.19 $Y=1.655 $X2=3.035 $Y2=1.95
cc_49 VPB N_C_c_93_n 0.0353619f $X=-0.19 $Y=1.655 $X2=2.745 $Y2=2.07
cc_50 VPB N_C_c_94_n 0.00589938f $X=-0.19 $Y=1.655 $X2=2.69 $Y2=2.07
cc_51 VPB N_C_c_95_n 0.0353904f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=2.07
cc_52 VPB N_A_M1009_g 0.0164406f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.775
cc_53 VPB N_A_M1000_g 0.0363928f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=1.905
cc_54 VPB N_A_c_175_n 0.0134308f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.77
cc_55 VPB N_A_c_176_n 0.00958703f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.935
cc_56 VPB A 0.00278654f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.43
cc_57 VPB N_A_c_172_n 0.0217025f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=2.15
cc_58 VPB N_B_c_230_n 0.0188791f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.935
cc_59 VPB N_B_M1010_g 0.0373077f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.775
cc_60 VPB N_B_M1004_g 0.037134f $X=-0.19 $Y=1.655 $X2=2.685 $Y2=2.775
cc_61 VPB N_B_c_228_n 0.00764058f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=2.15
cc_62 VPB N_B_c_229_n 9.57312e-19 $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.15
cc_63 VPB N_A_59_491#_M1005_g 0.0225058f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.77
cc_64 VPB N_A_59_491#_M1013_g 0.0259807f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.15
cc_65 VPB N_A_59_491#_c_285_n 0.0369678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_59_491#_c_297_n 0.00924704f $X=-0.19 $Y=1.655 $X2=2.745 $Y2=2.07
cc_67 VPB N_A_59_491#_c_298_n 0.0411538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_418_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_419_n 0.00578219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_420_n 0.0106521f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.265
cc_71 VPB N_VPWR_c_421_n 0.0633614f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.935
cc_72 VPB N_VPWR_c_422_n 0.0347463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_423_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=2.15
cc_74 VPB N_VPWR_c_424_n 0.0294516f $X=-0.19 $Y=1.655 $X2=3.035 $Y2=1.95
cc_75 VPB N_VPWR_c_425_n 0.0252319f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=2.07
cc_76 VPB N_VPWR_c_426_n 0.00436716f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=2.07
cc_77 VPB N_VPWR_c_417_n 0.0462347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_X_c_483_n 0.00426611f $X=-0.19 $Y=1.655 $X2=2.685 $Y2=2.235
cc_79 VPB N_X_c_481_n 8.45165e-19 $X=-0.19 $Y=1.655 $X2=2.725 $Y2=0.455
cc_80 N_C_M1002_g N_A_M1003_g 0.0327071f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_81 N_C_c_95_n N_A_M1000_g 0.0100586f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_82 N_C_M1008_g N_A_c_175_n 0.0102625f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_83 N_C_c_82_n N_A_c_175_n 0.0327071f $X=0.605 $Y=1.77 $X2=0 $Y2=0
cc_84 N_C_c_83_n N_A_c_175_n 0.00279641f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_85 N_C_c_95_n N_A_c_175_n 0.00828264f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_86 N_C_M1008_g N_A_c_176_n 0.0567159f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_87 N_C_c_95_n N_A_c_176_n 0.00535682f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_88 N_C_M1002_g A 0.00228675f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_89 N_C_c_83_n A 0.0301543f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_90 N_C_c_95_n A 0.0542554f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_91 N_C_c_83_n N_A_c_172_n 0.00294342f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_92 N_C_c_84_n N_A_c_172_n 0.0327071f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_93 N_C_c_95_n N_A_c_172_n 0.00154709f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_94 N_C_c_95_n N_B_c_230_n 6.87623e-19 $X=2.525 $Y=2.07 $X2=-0.19 $Y2=-0.245
cc_95 N_C_c_95_n N_B_M1010_g 0.0145507f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_96 N_C_M1011_g N_B_M1004_g 0.0513974f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_97 N_C_c_93_n N_B_M1004_g 0.0204443f $X=2.745 $Y=2.07 $X2=0 $Y2=0
cc_98 N_C_c_94_n N_B_M1004_g 0.00431937f $X=2.69 $Y=2.07 $X2=0 $Y2=0
cc_99 N_C_c_95_n N_B_M1004_g 0.0157135f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_100 N_C_M1015_g N_B_M1014_g 0.0662722f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_101 N_C_M1015_g N_B_c_228_n 0.0260349f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_102 N_C_M1015_g N_B_c_229_n 0.0028429f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_103 N_C_c_95_n N_B_c_229_n 0.0247338f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_104 N_C_M1015_g N_A_59_491#_M1001_g 0.0278986f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_105 N_C_M1011_g N_A_59_491#_M1005_g 0.0112553f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_106 N_C_M1015_g N_A_59_491#_M1005_g 0.00783231f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_107 C N_A_59_491#_M1005_g 0.00324614f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_108 N_C_c_93_n N_A_59_491#_M1005_g 0.00773957f $X=2.745 $Y=2.07 $X2=0 $Y2=0
cc_109 N_C_M1008_g N_A_59_491#_c_285_n 0.00676992f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_110 N_C_M1002_g N_A_59_491#_c_285_n 0.00642101f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_111 N_C_c_83_n N_A_59_491#_c_285_n 0.05802f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_112 N_C_c_84_n N_A_59_491#_c_285_n 0.0148853f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_113 N_C_c_91_n N_A_59_491#_c_285_n 0.013787f $X=0.77 $Y=2.15 $X2=0 $Y2=0
cc_114 N_C_M1002_g N_A_59_491#_c_286_n 0.0147765f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_115 N_C_M1008_g N_A_59_491#_c_297_n 0.00861729f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_116 N_C_M1011_g N_A_59_491#_c_297_n 4.79243e-19 $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_117 N_C_c_95_n N_A_59_491#_c_297_n 0.105619f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_118 N_C_M1002_g N_A_59_491#_c_287_n 0.0111275f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_119 N_C_M1002_g N_A_59_491#_c_288_n 0.00469762f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_120 N_C_c_83_n N_A_59_491#_c_288_n 0.0202605f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_121 N_C_c_84_n N_A_59_491#_c_288_n 0.00117077f $X=0.605 $Y=1.43 $X2=0 $Y2=0
cc_122 N_C_M1011_g N_A_59_491#_c_317_n 0.00135784f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_123 N_C_M1015_g N_A_59_491#_c_318_n 0.00207813f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_124 N_C_M1015_g N_A_59_491#_c_289_n 0.0186808f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_125 N_C_M1015_g N_A_59_491#_c_290_n 0.00484273f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_126 N_C_M1008_g N_A_59_491#_c_298_n 0.0151155f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_127 N_C_c_89_n N_A_59_491#_c_298_n 5.67461e-19 $X=0.605 $Y=1.935 $X2=0 $Y2=0
cc_128 N_C_c_91_n N_A_59_491#_c_298_n 0.0268068f $X=0.77 $Y=2.15 $X2=0 $Y2=0
cc_129 N_C_M1015_g N_A_59_491#_c_292_n 0.00424902f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_130 C N_A_59_491#_c_292_n 0.016374f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_131 N_C_M1015_g N_A_59_491#_c_293_n 0.0125301f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_132 C N_A_59_491#_c_293_n 0.00321274f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_133 C N_VPWR_M1011_d 0.0143944f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_134 N_C_M1008_g N_VPWR_c_418_n 0.00208736f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_135 N_C_M1011_g N_VPWR_c_419_n 0.0175306f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_136 C N_VPWR_c_419_n 0.0270284f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_137 N_C_c_93_n N_VPWR_c_419_n 0.0036332f $X=2.745 $Y=2.07 $X2=0 $Y2=0
cc_138 N_C_M1011_g N_VPWR_c_422_n 0.00486043f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_139 N_C_M1008_g N_VPWR_c_424_n 0.00427116f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_140 N_C_M1008_g N_VPWR_c_417_n 0.00721535f $X=0.655 $Y=2.775 $X2=0 $Y2=0
cc_141 N_C_M1011_g N_VPWR_c_417_n 0.00827383f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_142 N_C_M1015_g N_X_c_483_n 4.72317e-19 $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_143 C N_X_c_483_n 0.0230175f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_144 N_C_c_93_n N_X_c_483_n 2.2968e-19 $X=2.745 $Y=2.07 $X2=0 $Y2=0
cc_145 N_C_M1011_g N_X_c_488_n 9.72613e-19 $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_146 N_C_M1015_g N_X_c_489_n 9.59835e-19 $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_147 N_C_M1002_g N_VGND_c_518_n 0.00234408f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_148 N_C_M1015_g N_VGND_c_519_n 0.0131192f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_149 N_C_M1015_g N_VGND_c_522_n 0.00477554f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_150 N_C_M1002_g N_VGND_c_524_n 0.00539624f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_151 N_C_M1002_g N_VGND_c_527_n 0.0109911f $X=0.695 $Y=0.455 $X2=0 $Y2=0
cc_152 N_C_M1015_g N_VGND_c_527_n 0.00822887f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_153 A N_B_c_230_n 0.00406885f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_154 N_A_c_172_n N_B_c_230_n 0.0407093f $X=1.25 $Y=1.38 $X2=-0.19 $Y2=-0.245
cc_155 N_A_M1000_g N_B_M1010_g 0.0407093f $X=1.475 $Y=2.775 $X2=0 $Y2=0
cc_156 N_A_M1006_g N_B_M1007_g 0.0333401f $X=1.515 $Y=0.455 $X2=0 $Y2=0
cc_157 A N_B_c_227_n 0.00519684f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A_c_172_n N_B_c_227_n 0.0333401f $X=1.25 $Y=1.38 $X2=0 $Y2=0
cc_159 N_A_c_172_n N_B_c_228_n 0.0162234f $X=1.25 $Y=1.38 $X2=0 $Y2=0
cc_160 A N_B_c_229_n 0.0522891f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_161 N_A_c_172_n N_B_c_229_n 4.59271e-19 $X=1.25 $Y=1.38 $X2=0 $Y2=0
cc_162 N_A_M1003_g N_A_59_491#_c_286_n 0.00208107f $X=1.085 $Y=0.455 $X2=0 $Y2=0
cc_163 N_A_M1009_g N_A_59_491#_c_297_n 0.011768f $X=1.045 $Y=2.775 $X2=0 $Y2=0
cc_164 N_A_M1000_g N_A_59_491#_c_297_n 0.011768f $X=1.475 $Y=2.775 $X2=0 $Y2=0
cc_165 N_A_c_176_n N_A_59_491#_c_297_n 0.00116336f $X=1.065 $Y=2.325 $X2=0 $Y2=0
cc_166 N_A_M1003_g N_A_59_491#_c_287_n 0.0163744f $X=1.085 $Y=0.455 $X2=0 $Y2=0
cc_167 N_A_M1006_g N_A_59_491#_c_287_n 0.0141145f $X=1.515 $Y=0.455 $X2=0 $Y2=0
cc_168 A N_A_59_491#_c_287_n 0.0541139f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A_c_172_n N_A_59_491#_c_287_n 0.00259406f $X=1.25 $Y=1.38 $X2=0 $Y2=0
cc_170 N_A_M1000_g N_A_59_491#_c_317_n 0.00173846f $X=1.475 $Y=2.775 $X2=0 $Y2=0
cc_171 N_A_M1006_g N_A_59_491#_c_318_n 0.00207813f $X=1.515 $Y=0.455 $X2=0 $Y2=0
cc_172 N_A_M1009_g N_A_59_491#_c_298_n 0.00173296f $X=1.045 $Y=2.775 $X2=0 $Y2=0
cc_173 N_A_M1009_g N_VPWR_c_418_n 0.0106592f $X=1.045 $Y=2.775 $X2=0 $Y2=0
cc_174 N_A_M1000_g N_VPWR_c_418_n 0.0106632f $X=1.475 $Y=2.775 $X2=0 $Y2=0
cc_175 N_A_M1000_g N_VPWR_c_422_n 0.00366311f $X=1.475 $Y=2.775 $X2=0 $Y2=0
cc_176 N_A_M1009_g N_VPWR_c_424_n 0.00366311f $X=1.045 $Y=2.775 $X2=0 $Y2=0
cc_177 N_A_M1009_g N_VPWR_c_417_n 0.00433859f $X=1.045 $Y=2.775 $X2=0 $Y2=0
cc_178 N_A_M1000_g N_VPWR_c_417_n 0.00433859f $X=1.475 $Y=2.775 $X2=0 $Y2=0
cc_179 N_A_M1003_g N_VGND_c_518_n 0.0130723f $X=1.085 $Y=0.455 $X2=0 $Y2=0
cc_180 N_A_M1006_g N_VGND_c_518_n 0.0130723f $X=1.515 $Y=0.455 $X2=0 $Y2=0
cc_181 N_A_M1006_g N_VGND_c_522_n 0.00477554f $X=1.515 $Y=0.455 $X2=0 $Y2=0
cc_182 N_A_M1003_g N_VGND_c_524_n 0.00477554f $X=1.085 $Y=0.455 $X2=0 $Y2=0
cc_183 N_A_M1003_g N_VGND_c_527_n 0.00822887f $X=1.085 $Y=0.455 $X2=0 $Y2=0
cc_184 N_A_M1006_g N_VGND_c_527_n 0.00822887f $X=1.515 $Y=0.455 $X2=0 $Y2=0
cc_185 N_B_M1010_g N_A_59_491#_c_297_n 0.0109292f $X=1.865 $Y=2.775 $X2=0 $Y2=0
cc_186 N_B_M1004_g N_A_59_491#_c_297_n 0.00474967f $X=2.295 $Y=2.775 $X2=0 $Y2=0
cc_187 N_B_M1007_g N_A_59_491#_c_287_n 0.0146407f $X=1.905 $Y=0.455 $X2=0 $Y2=0
cc_188 N_B_M1010_g N_A_59_491#_c_317_n 0.00992358f $X=1.865 $Y=2.775 $X2=0 $Y2=0
cc_189 N_B_M1004_g N_A_59_491#_c_317_n 0.00972272f $X=2.295 $Y=2.775 $X2=0 $Y2=0
cc_190 N_B_M1007_g N_A_59_491#_c_318_n 0.0129069f $X=1.905 $Y=0.455 $X2=0 $Y2=0
cc_191 N_B_M1014_g N_A_59_491#_c_318_n 0.0129069f $X=2.335 $Y=0.455 $X2=0 $Y2=0
cc_192 N_B_M1014_g N_A_59_491#_c_289_n 0.013791f $X=2.335 $Y=0.455 $X2=0 $Y2=0
cc_193 N_B_c_229_n N_A_59_491#_c_289_n 0.00171113f $X=2.145 $Y=1.38 $X2=0 $Y2=0
cc_194 N_B_c_229_n N_A_59_491#_c_290_n 0.00193777f $X=2.145 $Y=1.38 $X2=0 $Y2=0
cc_195 N_B_M1007_g N_A_59_491#_c_291_n 0.00372856f $X=1.905 $Y=0.455 $X2=0 $Y2=0
cc_196 N_B_M1014_g N_A_59_491#_c_291_n 0.0028029f $X=2.335 $Y=0.455 $X2=0 $Y2=0
cc_197 N_B_c_227_n N_A_59_491#_c_291_n 7.76954e-19 $X=2.12 $Y=1.365 $X2=0 $Y2=0
cc_198 N_B_c_229_n N_A_59_491#_c_291_n 0.0258126f $X=2.145 $Y=1.38 $X2=0 $Y2=0
cc_199 N_B_c_229_n N_A_59_491#_c_292_n 0.00993782f $X=2.145 $Y=1.38 $X2=0 $Y2=0
cc_200 N_B_M1010_g N_VPWR_c_418_n 0.00208565f $X=1.865 $Y=2.775 $X2=0 $Y2=0
cc_201 N_B_M1004_g N_VPWR_c_419_n 0.0030761f $X=2.295 $Y=2.775 $X2=0 $Y2=0
cc_202 N_B_M1010_g N_VPWR_c_422_n 0.00428586f $X=1.865 $Y=2.775 $X2=0 $Y2=0
cc_203 N_B_M1004_g N_VPWR_c_422_n 0.00549284f $X=2.295 $Y=2.775 $X2=0 $Y2=0
cc_204 N_B_M1010_g N_VPWR_c_417_n 0.00606026f $X=1.865 $Y=2.775 $X2=0 $Y2=0
cc_205 N_B_M1004_g N_VPWR_c_417_n 0.0100104f $X=2.295 $Y=2.775 $X2=0 $Y2=0
cc_206 N_B_M1007_g N_VGND_c_518_n 0.00234408f $X=1.905 $Y=0.455 $X2=0 $Y2=0
cc_207 N_B_M1014_g N_VGND_c_519_n 0.00234408f $X=2.335 $Y=0.455 $X2=0 $Y2=0
cc_208 N_B_M1007_g N_VGND_c_522_n 0.00539624f $X=1.905 $Y=0.455 $X2=0 $Y2=0
cc_209 N_B_M1014_g N_VGND_c_522_n 0.00539624f $X=2.335 $Y=0.455 $X2=0 $Y2=0
cc_210 N_B_M1007_g N_VGND_c_527_n 0.00990635f $X=1.905 $Y=0.455 $X2=0 $Y2=0
cc_211 N_B_M1014_g N_VGND_c_527_n 0.00990635f $X=2.335 $Y=0.455 $X2=0 $Y2=0
cc_212 N_A_59_491#_c_297_n A_146_491# 0.0024629f $X=1.915 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_59_491#_c_297_n N_VPWR_M1009_d 0.00176557f $X=1.915 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_59_491#_c_297_n N_VPWR_c_418_n 0.0156967f $X=1.915 $Y=2.5 $X2=0 $Y2=0
cc_215 N_A_59_491#_c_317_n N_VPWR_c_418_n 0.0095042f $X=2.08 $Y=2.74 $X2=0 $Y2=0
cc_216 N_A_59_491#_c_298_n N_VPWR_c_418_n 0.00982657f $X=0.605 $Y=2.74 $X2=0
+ $Y2=0
cc_217 N_A_59_491#_M1005_g N_VPWR_c_419_n 0.00905242f $X=3.395 $Y=2.465 $X2=0
+ $Y2=0
cc_218 N_A_59_491#_c_297_n N_VPWR_c_419_n 0.00571183f $X=1.915 $Y=2.5 $X2=0
+ $Y2=0
cc_219 N_A_59_491#_c_317_n N_VPWR_c_419_n 0.0151909f $X=2.08 $Y=2.74 $X2=0 $Y2=0
cc_220 N_A_59_491#_M1013_g N_VPWR_c_421_n 0.00903023f $X=3.825 $Y=2.465 $X2=0
+ $Y2=0
cc_221 N_A_59_491#_c_297_n N_VPWR_c_422_n 0.00577798f $X=1.915 $Y=2.5 $X2=0
+ $Y2=0
cc_222 N_A_59_491#_c_317_n N_VPWR_c_422_n 0.01781f $X=2.08 $Y=2.74 $X2=0 $Y2=0
cc_223 N_A_59_491#_c_297_n N_VPWR_c_424_n 0.00577798f $X=1.915 $Y=2.5 $X2=0
+ $Y2=0
cc_224 N_A_59_491#_c_298_n N_VPWR_c_424_n 0.0320591f $X=0.605 $Y=2.74 $X2=0
+ $Y2=0
cc_225 N_A_59_491#_M1005_g N_VPWR_c_425_n 0.00549284f $X=3.395 $Y=2.465 $X2=0
+ $Y2=0
cc_226 N_A_59_491#_M1013_g N_VPWR_c_425_n 0.00549284f $X=3.825 $Y=2.465 $X2=0
+ $Y2=0
cc_227 N_A_59_491#_M1008_s N_VPWR_c_417_n 0.00233022f $X=0.295 $Y=2.455 $X2=0
+ $Y2=0
cc_228 N_A_59_491#_M1010_d N_VPWR_c_417_n 0.0022543f $X=1.94 $Y=2.455 $X2=0
+ $Y2=0
cc_229 N_A_59_491#_M1005_g N_VPWR_c_417_n 0.0106221f $X=3.395 $Y=2.465 $X2=0
+ $Y2=0
cc_230 N_A_59_491#_M1013_g N_VPWR_c_417_n 0.0107443f $X=3.825 $Y=2.465 $X2=0
+ $Y2=0
cc_231 N_A_59_491#_c_297_n N_VPWR_c_417_n 0.0244981f $X=1.915 $Y=2.5 $X2=0 $Y2=0
cc_232 N_A_59_491#_c_317_n N_VPWR_c_417_n 0.0124547f $X=2.08 $Y=2.74 $X2=0 $Y2=0
cc_233 N_A_59_491#_c_298_n N_VPWR_c_417_n 0.0197704f $X=0.605 $Y=2.74 $X2=0
+ $Y2=0
cc_234 N_A_59_491#_c_297_n A_310_491# 0.0024629f $X=1.915 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_59_491#_M1005_g N_X_c_483_n 0.00465717f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_59_491#_M1013_g N_X_c_483_n 0.00226992f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_59_491#_c_293_n N_X_c_483_n 0.00177921f $X=3.665 $Y=1.435 $X2=0 $Y2=0
cc_238 N_A_59_491#_M1005_g N_X_c_488_n 0.0193059f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A_59_491#_M1013_g N_X_c_488_n 0.0141675f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_59_491#_M1001_g N_X_c_481_n 4.73407e-19 $X=3.235 $Y=0.665 $X2=0 $Y2=0
cc_241 N_A_59_491#_M1012_g N_X_c_481_n 0.00634628f $X=3.665 $Y=0.665 $X2=0 $Y2=0
cc_242 N_A_59_491#_M1013_g N_X_c_481_n 0.0176122f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A_59_491#_c_290_n N_X_c_481_n 0.00410914f $X=3.02 $Y=1.285 $X2=0 $Y2=0
cc_244 N_A_59_491#_c_292_n N_X_c_481_n 0.0238922f $X=3.26 $Y=1.45 $X2=0 $Y2=0
cc_245 N_A_59_491#_c_293_n N_X_c_481_n 0.0164514f $X=3.665 $Y=1.435 $X2=0 $Y2=0
cc_246 N_A_59_491#_M1001_g N_X_c_489_n 0.00953732f $X=3.235 $Y=0.665 $X2=0 $Y2=0
cc_247 N_A_59_491#_M1012_g N_X_c_489_n 0.0197729f $X=3.665 $Y=0.665 $X2=0 $Y2=0
cc_248 N_A_59_491#_M1001_g X 0.00317517f $X=3.235 $Y=0.665 $X2=0 $Y2=0
cc_249 N_A_59_491#_M1012_g X 0.00795695f $X=3.665 $Y=0.665 $X2=0 $Y2=0
cc_250 N_A_59_491#_c_290_n X 0.00335182f $X=3.02 $Y=1.285 $X2=0 $Y2=0
cc_251 N_A_59_491#_c_292_n X 0.0111211f $X=3.26 $Y=1.45 $X2=0 $Y2=0
cc_252 N_A_59_491#_c_293_n X 0.004267f $X=3.665 $Y=1.435 $X2=0 $Y2=0
cc_253 N_A_59_491#_c_289_n N_VGND_M1015_d 0.00417717f $X=2.935 $Y=0.95 $X2=0
+ $Y2=0
cc_254 N_A_59_491#_c_290_n N_VGND_M1015_d 8.89872e-19 $X=3.02 $Y=1.285 $X2=0
+ $Y2=0
cc_255 N_A_59_491#_c_286_n N_VGND_c_518_n 0.0133059f $X=0.48 $Y=0.475 $X2=0
+ $Y2=0
cc_256 N_A_59_491#_c_287_n N_VGND_c_518_n 0.026201f $X=1.955 $Y=0.95 $X2=0 $Y2=0
cc_257 N_A_59_491#_c_318_n N_VGND_c_518_n 0.0133059f $X=2.12 $Y=0.475 $X2=0
+ $Y2=0
cc_258 N_A_59_491#_M1001_g N_VGND_c_519_n 0.00523621f $X=3.235 $Y=0.665 $X2=0
+ $Y2=0
cc_259 N_A_59_491#_c_318_n N_VGND_c_519_n 0.0133059f $X=2.12 $Y=0.475 $X2=0
+ $Y2=0
cc_260 N_A_59_491#_c_289_n N_VGND_c_519_n 0.0262415f $X=2.935 $Y=0.95 $X2=0
+ $Y2=0
cc_261 N_A_59_491#_M1012_g N_VGND_c_521_n 0.00959302f $X=3.665 $Y=0.665 $X2=0
+ $Y2=0
cc_262 N_A_59_491#_c_318_n N_VGND_c_522_n 0.0178561f $X=2.12 $Y=0.475 $X2=0
+ $Y2=0
cc_263 N_A_59_491#_c_286_n N_VGND_c_524_n 0.0196261f $X=0.48 $Y=0.475 $X2=0
+ $Y2=0
cc_264 N_A_59_491#_M1001_g N_VGND_c_525_n 0.00539624f $X=3.235 $Y=0.665 $X2=0
+ $Y2=0
cc_265 N_A_59_491#_M1012_g N_VGND_c_525_n 0.00353054f $X=3.665 $Y=0.665 $X2=0
+ $Y2=0
cc_266 N_A_59_491#_M1002_s N_VGND_c_527_n 0.00229455f $X=0.335 $Y=0.245 $X2=0
+ $Y2=0
cc_267 N_A_59_491#_M1007_d N_VGND_c_527_n 0.0022543f $X=1.98 $Y=0.245 $X2=0
+ $Y2=0
cc_268 N_A_59_491#_M1001_g N_VGND_c_527_n 0.0100586f $X=3.235 $Y=0.665 $X2=0
+ $Y2=0
cc_269 N_A_59_491#_M1012_g N_VGND_c_527_n 0.00636855f $X=3.665 $Y=0.665 $X2=0
+ $Y2=0
cc_270 N_A_59_491#_c_286_n N_VGND_c_527_n 0.0125379f $X=0.48 $Y=0.475 $X2=0
+ $Y2=0
cc_271 N_A_59_491#_c_318_n N_VGND_c_527_n 0.0124703f $X=2.12 $Y=0.475 $X2=0
+ $Y2=0
cc_272 N_A_59_491#_c_289_n N_VGND_c_527_n 5.7995e-19 $X=2.935 $Y=0.95 $X2=0
+ $Y2=0
cc_273 A_146_491# N_VPWR_c_417_n 0.00318022f $X=0.73 $Y=2.455 $X2=3.02 $Y2=1.285
cc_274 N_VPWR_c_417_n A_310_491# 0.00318022f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_275 N_VPWR_c_417_n A_474_491# 0.010279f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_276 N_VPWR_c_417_n N_X_M1005_s 0.00223819f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_277 N_VPWR_c_421_n N_X_c_483_n 0.0469769f $X=4.04 $Y=1.96 $X2=0 $Y2=0
cc_278 N_VPWR_c_419_n N_X_c_488_n 0.0272566f $X=2.9 $Y=2.58 $X2=0 $Y2=0
cc_279 N_VPWR_c_425_n N_X_c_488_n 0.0177952f $X=3.955 $Y=3.33 $X2=0 $Y2=0
cc_280 N_VPWR_c_417_n N_X_c_488_n 0.0123247f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_281 X N_VGND_c_521_n 0.03181f $X=3.6 $Y=0.925 $X2=0 $Y2=0
cc_282 N_X_c_489_n N_VGND_c_525_n 0.0269934f $X=3.45 $Y=0.43 $X2=0 $Y2=0
cc_283 N_X_M1001_d N_VGND_c_527_n 0.00223819f $X=3.31 $Y=0.245 $X2=0 $Y2=0
cc_284 N_X_c_489_n N_VGND_c_527_n 0.0179352f $X=3.45 $Y=0.43 $X2=0 $Y2=0
cc_285 A_154_49# N_VGND_c_527_n 0.010279f $X=0.77 $Y=0.245 $X2=4.08 $Y2=0
cc_286 N_VGND_c_527_n A_318_49# 0.010279f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_287 N_VGND_c_527_n A_482_49# 0.010279f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
