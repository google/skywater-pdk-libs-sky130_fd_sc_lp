* File: sky130_fd_sc_lp__mux4_1.spice
* Created: Fri Aug 28 10:46:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux4_1.pex.spice"
.subckt sky130_fd_sc_lp__mux4_1  VNB VPB A1 A0 S0 A3 A2 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A2	A2
* A3	A3
* S0	S0
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_A1_M1014_g N_A_33_81#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.1113 PD=0.75 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1008 A_212_81# N_A0_M1008_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0693 PD=0.63 PS=0.75 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_284_81#_M1009_d N_A_254_55#_M1009_g A_212_81# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_A_33_81#_M1018_d N_S0_M1018_g N_A_284_81#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1407 AS=0.0588 PD=1.51 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_S0_M1011_g N_A_254_55#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.110925 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_A_793_117#_M1016_d N_S0_M1016_g N_A_710_117#_M1016_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_879_117#_M1007_d N_A_254_55#_M1007_g N_A_793_117#_M1016_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A3_M1012_g N_A_710_117#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_879_117#_M1015_d N_A2_M1015_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0756 PD=1.37 PS=0.78 NRD=0 NRS=2.856 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_1245_21#_M1004_d N_S1_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_1635_149#_M1001_d N_S1_M1001_g N_A_793_117#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.2247 PD=0.7 PS=1.91 NRD=0 NRS=77.136 M=1 R=2.8
+ SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_284_81#_M1006_d N_A_1245_21#_M1006_g N_A_1635_149#_M1001_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_X_M1020_d N_A_1635_149#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_27_519#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1013 N_A_196_519#_M1013_d N_A0_M1013_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_284_81#_M1005_d N_A_254_55#_M1005_g N_A_27_519#_M1005_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_A_196_519#_M1023_d N_S0_M1023_g N_A_284_81#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.0588 PD=1.43 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_S0_M1021_g N_A_254_55#_M1021_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_793_117#_M1003_d N_S0_M1003_g N_A_799_501#_M1003_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1024 A_968_501# N_A_254_55#_M1024_g N_A_793_117#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A3_M1019_g A_968_501# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=21.0987 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1025 N_A_799_501#_M1025_d N_A2_M1025_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0735 PD=1.37 PS=0.77 NRD=0 NRS=11.7215 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_1245_21#_M1010_d N_S1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1449 PD=1.37 PS=1.53 NRD=0 NRS=32.8202 M=1 R=2.8
+ SA=75000.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_A_1635_149#_M1017_d N_S1_M1017_g N_A_284_81#_M1017_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_793_117#_M1022_d N_A_1245_21#_M1022_g N_A_1635_149#_M1017_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_1635_149#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=19.5079 P=24.65
c_112 VNB 0 3.62571e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__mux4_1.pxi.spice"
*
.ends
*
*
