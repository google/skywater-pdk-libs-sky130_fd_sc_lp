* File: sky130_fd_sc_lp__o41a_4.pxi.spice
* Created: Wed Sep  2 10:27:41 2020
* 
x_PM_SKY130_FD_SC_LP__O41A_4%A_83_23# N_A_83_23#_M1013_s N_A_83_23#_M1004_d
+ N_A_83_23#_M1002_d N_A_83_23#_M1000_g N_A_83_23#_M1006_g N_A_83_23#_M1010_g
+ N_A_83_23#_M1009_g N_A_83_23#_M1011_g N_A_83_23#_M1019_g N_A_83_23#_M1016_g
+ N_A_83_23#_M1020_g N_A_83_23#_c_127_n N_A_83_23#_c_128_n N_A_83_23#_c_129_n
+ N_A_83_23#_c_138_n N_A_83_23#_c_149_p N_A_83_23#_c_130_n N_A_83_23#_c_131_n
+ N_A_83_23#_c_215_p N_A_83_23#_c_150_p N_A_83_23#_c_132_n
+ PM_SKY130_FD_SC_LP__O41A_4%A_83_23#
x_PM_SKY130_FD_SC_LP__O41A_4%B1 N_B1_M1004_g N_B1_M1017_g N_B1_c_253_n
+ N_B1_M1013_g N_B1_c_254_n N_B1_M1026_g B1 N_B1_c_256_n
+ PM_SKY130_FD_SC_LP__O41A_4%B1
x_PM_SKY130_FD_SC_LP__O41A_4%A4 N_A4_c_305_n N_A4_M1024_g N_A4_M1002_g
+ N_A4_c_307_n N_A4_M1025_g N_A4_M1008_g A4 N_A4_c_310_n
+ PM_SKY130_FD_SC_LP__O41A_4%A4
x_PM_SKY130_FD_SC_LP__O41A_4%A3 N_A3_c_351_n N_A3_M1012_g N_A3_M1014_g
+ N_A3_c_353_n N_A3_M1023_g N_A3_M1027_g A3 A3 A3 N_A3_c_356_n
+ PM_SKY130_FD_SC_LP__O41A_4%A3
x_PM_SKY130_FD_SC_LP__O41A_4%A2 N_A2_c_403_n N_A2_M1003_g N_A2_c_404_n
+ N_A2_c_405_n N_A2_M1015_g N_A2_c_407_n N_A2_M1007_g N_A2_M1021_g A2 A2
+ N_A2_c_409_n PM_SKY130_FD_SC_LP__O41A_4%A2
x_PM_SKY130_FD_SC_LP__O41A_4%A1 N_A1_c_452_n N_A1_M1001_g N_A1_M1005_g
+ N_A1_c_454_n N_A1_M1018_g N_A1_M1022_g A1 A1 A1 N_A1_c_457_n
+ PM_SKY130_FD_SC_LP__O41A_4%A1
x_PM_SKY130_FD_SC_LP__O41A_4%VPWR N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_M1020_d
+ N_VPWR_M1017_s N_VPWR_M1005_d N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n
+ N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n
+ N_VPWR_c_498_n N_VPWR_c_499_n VPWR N_VPWR_c_500_n N_VPWR_c_501_n
+ N_VPWR_c_502_n N_VPWR_c_489_n N_VPWR_c_504_n N_VPWR_c_505_n
+ PM_SKY130_FD_SC_LP__O41A_4%VPWR
x_PM_SKY130_FD_SC_LP__O41A_4%X N_X_M1000_d N_X_M1011_d N_X_M1006_s N_X_M1019_s
+ N_X_c_591_n N_X_c_596_n N_X_c_597_n N_X_c_644_p N_X_c_629_n N_X_c_592_n
+ N_X_c_598_n N_X_c_643_p N_X_c_634_n N_X_c_593_n N_X_c_599_n X X N_X_c_594_n X
+ PM_SKY130_FD_SC_LP__O41A_4%X
x_PM_SKY130_FD_SC_LP__O41A_4%A_652_345# N_A_652_345#_M1002_s
+ N_A_652_345#_M1008_s N_A_652_345#_M1027_d N_A_652_345#_c_649_n
+ N_A_652_345#_c_650_n N_A_652_345#_c_651_n N_A_652_345#_c_665_n
+ N_A_652_345#_c_652_n N_A_652_345#_c_653_n N_A_652_345#_c_678_n
+ PM_SKY130_FD_SC_LP__O41A_4%A_652_345#
x_PM_SKY130_FD_SC_LP__O41A_4%A_907_345# N_A_907_345#_M1014_s
+ N_A_907_345#_M1015_s N_A_907_345#_c_716_n N_A_907_345#_c_699_n
+ N_A_907_345#_c_700_n N_A_907_345#_c_704_n N_A_907_345#_c_706_n
+ PM_SKY130_FD_SC_LP__O41A_4%A_907_345#
x_PM_SKY130_FD_SC_LP__O41A_4%A_1108_367# N_A_1108_367#_M1015_d
+ N_A_1108_367#_M1021_d N_A_1108_367#_M1022_s N_A_1108_367#_c_724_n
+ N_A_1108_367#_c_725_n N_A_1108_367#_c_726_n N_A_1108_367#_c_748_n
+ N_A_1108_367#_c_727_n N_A_1108_367#_c_752_n N_A_1108_367#_c_728_n
+ PM_SKY130_FD_SC_LP__O41A_4%A_1108_367#
x_PM_SKY130_FD_SC_LP__O41A_4%VGND N_VGND_M1000_s N_VGND_M1010_s N_VGND_M1016_s
+ N_VGND_M1024_d N_VGND_M1012_d N_VGND_M1003_s N_VGND_M1001_s N_VGND_c_763_n
+ N_VGND_c_764_n N_VGND_c_765_n N_VGND_c_766_n N_VGND_c_767_n N_VGND_c_768_n
+ N_VGND_c_769_n N_VGND_c_770_n N_VGND_c_771_n N_VGND_c_772_n N_VGND_c_773_n
+ N_VGND_c_774_n N_VGND_c_775_n N_VGND_c_776_n VGND N_VGND_c_777_n
+ N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n
+ N_VGND_c_783_n PM_SKY130_FD_SC_LP__O41A_4%VGND
x_PM_SKY130_FD_SC_LP__O41A_4%A_480_47# N_A_480_47#_M1013_d N_A_480_47#_M1026_d
+ N_A_480_47#_M1025_s N_A_480_47#_M1023_s N_A_480_47#_M1007_d
+ N_A_480_47#_M1018_d N_A_480_47#_c_883_n N_A_480_47#_c_886_n
+ N_A_480_47#_c_887_n N_A_480_47#_c_932_n N_A_480_47#_c_900_n
+ N_A_480_47#_c_936_n N_A_480_47#_c_908_n N_A_480_47#_c_940_n
+ N_A_480_47#_c_877_n N_A_480_47#_c_878_n N_A_480_47#_c_879_n
+ N_A_480_47#_c_904_n N_A_480_47#_c_906_n N_A_480_47#_c_912_n
+ PM_SKY130_FD_SC_LP__O41A_4%A_480_47#
cc_1 VNB N_A_83_23#_M1000_g 0.025885f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.665
cc_2 VNB N_A_83_23#_M1010_g 0.0213918f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.665
cc_3 VNB N_A_83_23#_M1011_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.665
cc_4 VNB N_A_83_23#_M1016_g 0.0257797f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.665
cc_5 VNB N_A_83_23#_c_127_n 0.00720617f $X=-0.19 $Y=-0.245 $X2=2.32 $Y2=1.49
cc_6 VNB N_A_83_23#_c_128_n 0.00245458f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.395
cc_7 VNB N_A_83_23#_c_129_n 0.00219973f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=1.815
cc_8 VNB N_A_83_23#_c_130_n 0.00290207f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=0.95
cc_9 VNB N_A_83_23#_c_131_n 0.00301164f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=1.71
cc_10 VNB N_A_83_23#_c_132_n 0.0710376f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.49
cc_11 VNB N_B1_M1004_g 0.00658622f $X=-0.19 $Y=-0.245 $X2=3.675 $Y2=1.725
cc_12 VNB N_B1_M1017_g 0.0100315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_253_n 0.0193592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_254_n 0.0164415f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.665
cc_15 VNB B1 0.00317705f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_16 VNB N_B1_c_256_n 0.0868823f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_17 VNB N_A4_c_305_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.235
cc_18 VNB N_A4_M1002_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A4_c_307_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A4_M1008_g 0.00152414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A4 0.00191494f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_22 VNB N_A4_c_310_n 0.0369038f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.655
cc_23 VNB N_A3_c_351_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.235
cc_24 VNB N_A3_M1014_g 0.00152414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A3_c_353_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A3_M1027_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A3 0.00777036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A3_c_356_n 0.0447126f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.325
cc_29 VNB N_A2_c_403_n 0.0223198f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.235
cc_30 VNB N_A2_c_404_n 0.03501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_405_n 0.0183903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_M1015_g 0.0102769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_c_407_n 0.0223198f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.325
cc_34 VNB N_A2_M1021_g 0.00728015f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_35 VNB N_A2_c_409_n 0.0372146f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.325
cc_36 VNB N_A1_c_452_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.235
cc_37 VNB N_A1_M1005_g 0.00677981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_c_454_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A1_M1022_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB A1 0.0274896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A1_c_457_n 0.0500903f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_42 VNB N_VPWR_c_489_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_591_n 0.00143767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_592_n 0.00599427f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.665
cc_45 VNB N_X_c_593_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=2.32 $Y2=1.49
cc_46 VNB N_X_c_594_n 0.00919693f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.49
cc_47 VNB X 0.0218021f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.395
cc_48 VNB N_VGND_c_763_n 0.01092f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.655
cc_49 VNB N_VGND_c_764_n 0.0281524f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_50 VNB N_VGND_c_765_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.665
cc_51 VNB N_VGND_c_766_n 0.0146034f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_52 VNB N_VGND_c_767_n 0.00461568f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.665
cc_53 VNB N_VGND_c_768_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.655
cc_54 VNB N_VGND_c_769_n 0.00398746f $X=-0.19 $Y=-0.245 $X2=2.32 $Y2=1.49
cc_55 VNB N_VGND_c_770_n 0.00462055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_771_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.49
cc_57 VNB N_VGND_c_772_n 0.00501779f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.04
cc_58 VNB N_VGND_c_773_n 0.0376577f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.395
cc_59 VNB N_VGND_c_774_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=1.815
cc_60 VNB N_VGND_c_775_n 0.0167145f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=1.98
cc_61 VNB N_VGND_c_776_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=2.91
cc_62 VNB N_VGND_c_777_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=2.79 $Y2=0.95
cc_63 VNB N_VGND_c_778_n 0.0204173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_779_n 0.379781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_780_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_781_n 0.00490486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_782_n 0.0167145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_783_n 0.0210511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_480_47#_c_877_n 0.0075508f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.49
cc_70 VNB N_A_480_47#_c_878_n 0.0235425f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.49
cc_71 VNB N_A_480_47#_c_879_n 0.00456063f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.49
cc_72 VPB N_A_83_23#_M1006_g 0.0224142f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_73 VPB N_A_83_23#_M1009_g 0.0188421f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_74 VPB N_A_83_23#_M1019_g 0.0188632f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_75 VPB N_A_83_23#_M1020_g 0.019714f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_76 VPB N_A_83_23#_c_129_n 0.00174831f $X=-0.19 $Y=1.655 $X2=2.425 $Y2=1.815
cc_77 VPB N_A_83_23#_c_138_n 3.01779e-19 $X=-0.19 $Y=1.655 $X2=2.425 $Y2=1.98
cc_78 VPB N_A_83_23#_c_131_n 0.022366f $X=-0.19 $Y=1.655 $X2=3.72 $Y2=1.71
cc_79 VPB N_A_83_23#_c_132_n 0.00700947f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.49
cc_80 VPB N_B1_M1004_g 0.0197397f $X=-0.19 $Y=1.655 $X2=3.675 $Y2=1.725
cc_81 VPB N_B1_M1017_g 0.023307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A4_M1002_g 0.0245012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A4_M1008_g 0.0194248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A3_M1014_g 0.019309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A3_M1027_g 0.0246887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A2_M1015_g 0.023891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A2_M1021_g 0.0188441f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_88 VPB N_A1_M1005_g 0.018645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A1_M1022_g 0.0246191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_490_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_91 VPB N_VPWR_c_491_n 0.0415885f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.325
cc_92 VPB N_VPWR_c_492_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_93 VPB N_VPWR_c_493_n 0.00324451f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.655
cc_94 VPB N_VPWR_c_494_n 0.0132456f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.665
cc_95 VPB N_VPWR_c_495_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=2.32 $Y2=1.49
cc_96 VPB N_VPWR_c_496_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.49
cc_97 VPB N_VPWR_c_497_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.49
cc_98 VPB N_VPWR_c_498_n 0.012927f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.04
cc_99 VPB N_VPWR_c_499_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.395
cc_100 VPB N_VPWR_c_500_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.425 $Y2=1.98
cc_101 VPB N_VPWR_c_501_n 0.0892952f $X=-0.19 $Y=1.655 $X2=3.815 $Y2=2.57
cc_102 VPB N_VPWR_c_502_n 0.0170541f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.49
cc_103 VPB N_VPWR_c_489_n 0.0707231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_504_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_505_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_X_c_596_n 0.00143767f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_107 VPB N_X_c_597_n 0.00896757f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_108 VPB N_X_c_598_n 0.00531071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_X_c_599_n 0.00144314f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.49
cc_110 VPB X 0.00506177f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.395
cc_111 VPB N_A_652_345#_c_649_n 0.00867198f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.665
cc_112 VPB N_A_652_345#_c_650_n 0.00403194f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_113 VPB N_A_652_345#_c_651_n 0.0040695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_652_345#_c_652_n 0.00795953f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_115 VPB N_A_652_345#_c_653_n 0.00238942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_907_345#_c_699_n 0.0149504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_907_345#_c_700_n 0.00205773f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.655
cc_118 VPB N_A_1108_367#_c_724_n 0.00843415f $X=-0.19 $Y=1.655 $X2=0.49
+ $Y2=0.665
cc_119 VPB N_A_1108_367#_c_725_n 0.00357895f $X=-0.19 $Y=1.655 $X2=0.49
+ $Y2=1.655
cc_120 VPB N_A_1108_367#_c_726_n 0.00393881f $X=-0.19 $Y=1.655 $X2=0.49
+ $Y2=2.465
cc_121 VPB N_A_1108_367#_c_727_n 0.0112291f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.655
cc_122 VPB N_A_1108_367#_c_728_n 0.00202614f $X=-0.19 $Y=1.655 $X2=1.35
+ $Y2=1.655
cc_123 N_A_83_23#_c_127_n N_B1_M1004_g 0.0084026f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_124 N_A_83_23#_c_129_n N_B1_M1004_g 0.00630562f $X=2.425 $Y=1.815 $X2=0 $Y2=0
cc_125 N_A_83_23#_c_138_n N_B1_M1004_g 7.82894e-19 $X=2.425 $Y=1.98 $X2=0 $Y2=0
cc_126 N_A_83_23#_c_132_n N_B1_M1004_g 0.0229909f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_127 N_A_83_23#_c_129_n N_B1_M1017_g 0.00269499f $X=2.425 $Y=1.815 $X2=0 $Y2=0
cc_128 N_A_83_23#_c_138_n N_B1_M1017_g 0.00109751f $X=2.425 $Y=1.98 $X2=0 $Y2=0
cc_129 N_A_83_23#_c_131_n N_B1_M1017_g 0.0192202f $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_130 N_A_83_23#_c_128_n N_B1_c_253_n 0.0050767f $X=2.415 $Y=1.395 $X2=0 $Y2=0
cc_131 N_A_83_23#_c_149_p N_B1_c_253_n 0.0116765f $X=2.79 $Y=0.95 $X2=0 $Y2=0
cc_132 N_A_83_23#_c_150_p N_B1_c_253_n 0.00767008f $X=2.955 $Y=0.735 $X2=0 $Y2=0
cc_133 N_A_83_23#_c_150_p N_B1_c_254_n 0.00645311f $X=2.955 $Y=0.735 $X2=0 $Y2=0
cc_134 N_A_83_23#_c_128_n B1 0.013306f $X=2.415 $Y=1.395 $X2=0 $Y2=0
cc_135 N_A_83_23#_c_129_n B1 0.00312004f $X=2.425 $Y=1.815 $X2=0 $Y2=0
cc_136 N_A_83_23#_c_149_p B1 0.00695724f $X=2.79 $Y=0.95 $X2=0 $Y2=0
cc_137 N_A_83_23#_c_131_n B1 0.0442322f $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_138 N_A_83_23#_c_150_p B1 0.0205523f $X=2.955 $Y=0.735 $X2=0 $Y2=0
cc_139 N_A_83_23#_M1016_g N_B1_c_256_n 0.0229909f $X=1.78 $Y=0.665 $X2=0 $Y2=0
cc_140 N_A_83_23#_c_127_n N_B1_c_256_n 0.0104076f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_141 N_A_83_23#_c_128_n N_B1_c_256_n 0.0147955f $X=2.415 $Y=1.395 $X2=0 $Y2=0
cc_142 N_A_83_23#_c_129_n N_B1_c_256_n 0.00939386f $X=2.425 $Y=1.815 $X2=0 $Y2=0
cc_143 N_A_83_23#_c_149_p N_B1_c_256_n 0.00449095f $X=2.79 $Y=0.95 $X2=0 $Y2=0
cc_144 N_A_83_23#_c_131_n N_B1_c_256_n 0.0149795f $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_145 N_A_83_23#_c_150_p N_B1_c_256_n 0.00236751f $X=2.955 $Y=0.735 $X2=0 $Y2=0
cc_146 N_A_83_23#_c_131_n N_A4_M1002_g 0.0170961f $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_147 N_A_83_23#_c_131_n N_A4_M1008_g 9.83373e-19 $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_148 N_A_83_23#_c_131_n A4 0.0269632f $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_149 N_A_83_23#_c_131_n N_A4_c_310_n 0.00389015f $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_150 N_A_83_23#_M1006_g N_VPWR_c_491_n 0.0153838f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_83_23#_M1009_g N_VPWR_c_491_n 7.27171e-19 $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_83_23#_M1006_g N_VPWR_c_492_n 7.24342e-19 $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_83_23#_M1009_g N_VPWR_c_492_n 0.0141279f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_83_23#_M1019_g N_VPWR_c_492_n 0.0141279f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_83_23#_M1020_g N_VPWR_c_492_n 7.24342e-19 $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_83_23#_M1019_g N_VPWR_c_493_n 8.15296e-19 $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_83_23#_M1020_g N_VPWR_c_493_n 0.0195356f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_83_23#_c_127_n N_VPWR_c_493_n 0.0221617f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_159 N_A_83_23#_c_138_n N_VPWR_c_493_n 0.047967f $X=2.425 $Y=1.98 $X2=0 $Y2=0
cc_160 N_A_83_23#_c_131_n N_VPWR_c_494_n 0.0248366f $X=3.72 $Y=1.71 $X2=0 $Y2=0
cc_161 N_A_83_23#_M1019_g N_VPWR_c_496_n 0.00486043f $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_83_23#_M1020_g N_VPWR_c_496_n 0.00486043f $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_83_23#_c_138_n N_VPWR_c_498_n 0.0124525f $X=2.425 $Y=1.98 $X2=0 $Y2=0
cc_164 N_A_83_23#_M1006_g N_VPWR_c_500_n 0.00486043f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_83_23#_M1009_g N_VPWR_c_500_n 0.00486043f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_83_23#_M1004_d N_VPWR_c_489_n 0.00536646f $X=2.285 $Y=1.835 $X2=0
+ $Y2=0
cc_167 N_A_83_23#_M1006_g N_VPWR_c_489_n 0.00824727f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_83_23#_M1009_g N_VPWR_c_489_n 0.00824727f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_83_23#_M1019_g N_VPWR_c_489_n 0.00824727f $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_83_23#_M1020_g N_VPWR_c_489_n 0.00824727f $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_83_23#_c_138_n N_VPWR_c_489_n 0.00730901f $X=2.425 $Y=1.98 $X2=0
+ $Y2=0
cc_172 N_A_83_23#_M1000_g N_X_c_591_n 0.0163859f $X=0.49 $Y=0.665 $X2=0 $Y2=0
cc_173 N_A_83_23#_c_127_n N_X_c_591_n 0.00730993f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_174 N_A_83_23#_M1006_g N_X_c_596_n 0.0156636f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_83_23#_c_127_n N_X_c_596_n 0.00730993f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_176 N_A_83_23#_M1010_g N_X_c_592_n 0.0138879f $X=0.92 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A_83_23#_M1011_g N_X_c_592_n 0.0135652f $X=1.35 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A_83_23#_M1016_g N_X_c_592_n 0.00216603f $X=1.78 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_83_23#_c_127_n N_X_c_592_n 0.0625611f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_180 N_A_83_23#_c_128_n N_X_c_592_n 0.00375066f $X=2.415 $Y=1.395 $X2=0 $Y2=0
cc_181 N_A_83_23#_c_132_n N_X_c_592_n 0.00497162f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_182 N_A_83_23#_M1009_g N_X_c_598_n 0.0131755f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_83_23#_M1019_g N_X_c_598_n 0.0130133f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_83_23#_M1020_g N_X_c_598_n 0.00117092f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_83_23#_c_127_n N_X_c_598_n 0.0625611f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_186 N_A_83_23#_c_129_n N_X_c_598_n 0.00209731f $X=2.425 $Y=1.815 $X2=0 $Y2=0
cc_187 N_A_83_23#_c_132_n N_X_c_598_n 0.00497162f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_188 N_A_83_23#_c_127_n N_X_c_593_n 0.0154426f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_189 N_A_83_23#_c_132_n N_X_c_593_n 0.00253619f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_190 N_A_83_23#_c_127_n N_X_c_599_n 0.0154426f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_191 N_A_83_23#_c_132_n N_X_c_599_n 0.00253619f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_192 N_A_83_23#_M1000_g X 0.0201308f $X=0.49 $Y=0.665 $X2=0 $Y2=0
cc_193 N_A_83_23#_c_127_n X 0.015451f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_194 N_A_83_23#_c_131_n N_A_652_345#_M1002_s 0.00264426f $X=3.72 $Y=1.71
+ $X2=-0.19 $Y2=-0.245
cc_195 N_A_83_23#_c_131_n N_A_652_345#_c_649_n 0.0223219f $X=3.72 $Y=1.71 $X2=0
+ $Y2=0
cc_196 N_A_83_23#_M1002_d N_A_652_345#_c_650_n 0.00176461f $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_197 N_A_83_23#_c_215_p N_A_652_345#_c_650_n 0.0126348f $X=3.815 $Y=1.85 $X2=0
+ $Y2=0
cc_198 N_A_83_23#_c_131_n N_A_652_345#_c_653_n 0.0127664f $X=3.72 $Y=1.71 $X2=0
+ $Y2=0
cc_199 N_A_83_23#_M1000_g N_VGND_c_764_n 0.0117219f $X=0.49 $Y=0.665 $X2=0 $Y2=0
cc_200 N_A_83_23#_M1010_g N_VGND_c_764_n 6.10117e-19 $X=0.92 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_83_23#_M1000_g N_VGND_c_765_n 6.10117e-19 $X=0.49 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_83_23#_M1010_g N_VGND_c_765_n 0.0109182f $X=0.92 $Y=0.665 $X2=0 $Y2=0
cc_203 N_A_83_23#_M1011_g N_VGND_c_765_n 0.0109182f $X=1.35 $Y=0.665 $X2=0 $Y2=0
cc_204 N_A_83_23#_M1016_g N_VGND_c_765_n 6.10117e-19 $X=1.78 $Y=0.665 $X2=0
+ $Y2=0
cc_205 N_A_83_23#_M1011_g N_VGND_c_766_n 6.80895e-19 $X=1.35 $Y=0.665 $X2=0
+ $Y2=0
cc_206 N_A_83_23#_M1016_g N_VGND_c_766_n 0.0175492f $X=1.78 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A_83_23#_c_127_n N_VGND_c_766_n 0.0183854f $X=2.32 $Y=1.49 $X2=0 $Y2=0
cc_208 N_A_83_23#_c_128_n N_VGND_c_766_n 0.00514434f $X=2.415 $Y=1.395 $X2=0
+ $Y2=0
cc_209 N_A_83_23#_c_130_n N_VGND_c_766_n 0.0154392f $X=2.51 $Y=0.95 $X2=0 $Y2=0
cc_210 N_A_83_23#_c_150_p N_VGND_c_766_n 0.00493189f $X=2.955 $Y=0.735 $X2=0
+ $Y2=0
cc_211 N_A_83_23#_M1011_g N_VGND_c_771_n 0.00477554f $X=1.35 $Y=0.665 $X2=0
+ $Y2=0
cc_212 N_A_83_23#_M1016_g N_VGND_c_771_n 0.00477554f $X=1.78 $Y=0.665 $X2=0
+ $Y2=0
cc_213 N_A_83_23#_M1000_g N_VGND_c_777_n 0.00477554f $X=0.49 $Y=0.665 $X2=0
+ $Y2=0
cc_214 N_A_83_23#_M1010_g N_VGND_c_777_n 0.00477554f $X=0.92 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_83_23#_M1013_s N_VGND_c_779_n 0.00225186f $X=2.815 $Y=0.235 $X2=0
+ $Y2=0
cc_216 N_A_83_23#_M1000_g N_VGND_c_779_n 0.00825815f $X=0.49 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_83_23#_M1010_g N_VGND_c_779_n 0.00825815f $X=0.92 $Y=0.665 $X2=0
+ $Y2=0
cc_218 N_A_83_23#_M1011_g N_VGND_c_779_n 0.00825815f $X=1.35 $Y=0.665 $X2=0
+ $Y2=0
cc_219 N_A_83_23#_M1016_g N_VGND_c_779_n 0.00825815f $X=1.78 $Y=0.665 $X2=0
+ $Y2=0
cc_220 N_A_83_23#_c_149_p N_VGND_c_779_n 6.50149e-19 $X=2.79 $Y=0.95 $X2=0 $Y2=0
cc_221 N_A_83_23#_c_130_n N_VGND_c_779_n 0.00185388f $X=2.51 $Y=0.95 $X2=0 $Y2=0
cc_222 N_A_83_23#_c_128_n N_A_480_47#_M1013_d 3.95862e-19 $X=2.415 $Y=1.395
+ $X2=-0.19 $Y2=-0.245
cc_223 N_A_83_23#_c_149_p N_A_480_47#_M1013_d 0.00226064f $X=2.79 $Y=0.95
+ $X2=-0.19 $Y2=-0.245
cc_224 N_A_83_23#_c_130_n N_A_480_47#_M1013_d 0.00188466f $X=2.51 $Y=0.95
+ $X2=-0.19 $Y2=-0.245
cc_225 N_A_83_23#_M1013_s N_A_480_47#_c_883_n 0.00332344f $X=2.815 $Y=0.235
+ $X2=0 $Y2=0
cc_226 N_A_83_23#_c_149_p N_A_480_47#_c_883_n 0.00336912f $X=2.79 $Y=0.95 $X2=0
+ $Y2=0
cc_227 N_A_83_23#_c_150_p N_A_480_47#_c_883_n 0.0154725f $X=2.955 $Y=0.735 $X2=0
+ $Y2=0
cc_228 N_A_83_23#_c_131_n N_A_480_47#_c_886_n 0.00317151f $X=3.72 $Y=1.71 $X2=0
+ $Y2=0
cc_229 N_A_83_23#_c_131_n N_A_480_47#_c_887_n 0.00562534f $X=3.72 $Y=1.71 $X2=0
+ $Y2=0
cc_230 N_A_83_23#_M1016_g N_A_480_47#_c_879_n 9.33115e-19 $X=1.78 $Y=0.665 $X2=0
+ $Y2=0
cc_231 N_A_83_23#_c_149_p N_A_480_47#_c_879_n 0.00752362f $X=2.79 $Y=0.95 $X2=0
+ $Y2=0
cc_232 N_A_83_23#_c_130_n N_A_480_47#_c_879_n 0.0128326f $X=2.51 $Y=0.95 $X2=0
+ $Y2=0
cc_233 N_B1_c_254_n N_A4_c_305_n 0.0142501f $X=3.17 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_234 B1 A4 0.019637f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_235 N_B1_c_256_n A4 6.90096e-19 $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_236 B1 N_A4_c_310_n 7.76196e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_237 N_B1_c_256_n N_A4_c_310_n 0.0201725f $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_238 N_B1_M1004_g N_VPWR_c_493_n 0.019546f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1017_g N_VPWR_c_493_n 8.06385e-19 $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_M1004_g N_VPWR_c_494_n 7.58291e-19 $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B1_M1017_g N_VPWR_c_494_n 0.0184222f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B1_M1004_g N_VPWR_c_498_n 0.00486043f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1017_g N_VPWR_c_498_n 0.00486043f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B1_M1004_g N_VPWR_c_489_n 0.00824727f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_M1017_g N_VPWR_c_489_n 0.00824727f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B1_M1017_g N_A_652_345#_c_649_n 0.00170434f $X=2.64 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_B1_c_253_n N_VGND_c_766_n 0.00600791f $X=2.74 $Y=1.185 $X2=0 $Y2=0
cc_248 N_B1_c_256_n N_VGND_c_766_n 4.56546e-19 $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_249 N_B1_c_253_n N_VGND_c_773_n 0.00357877f $X=2.74 $Y=1.185 $X2=0 $Y2=0
cc_250 N_B1_c_254_n N_VGND_c_773_n 0.00357877f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_251 N_B1_c_253_n N_VGND_c_779_n 0.00681251f $X=2.74 $Y=1.185 $X2=0 $Y2=0
cc_252 N_B1_c_254_n N_VGND_c_779_n 0.00537654f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_253 N_B1_c_253_n N_A_480_47#_c_883_n 0.00989015f $X=2.74 $Y=1.185 $X2=0 $Y2=0
cc_254 N_B1_c_254_n N_A_480_47#_c_883_n 0.0114565f $X=3.17 $Y=1.185 $X2=0 $Y2=0
cc_255 N_B1_c_256_n N_A_480_47#_c_879_n 7.2246e-19 $X=3.17 $Y=1.35 $X2=0 $Y2=0
cc_256 N_A4_c_307_n N_A3_c_351_n 0.0145954f $X=4.03 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_257 N_A4_M1008_g N_A3_M1014_g 0.0245462f $X=4.03 $Y=2.355 $X2=0 $Y2=0
cc_258 A4 A3 0.0179136f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_259 N_A4_c_310_n A3 0.0141431f $X=4.03 $Y=1.35 $X2=0 $Y2=0
cc_260 N_A4_c_310_n N_A3_c_356_n 0.0234213f $X=4.03 $Y=1.35 $X2=0 $Y2=0
cc_261 N_A4_M1002_g N_VPWR_c_494_n 0.00269693f $X=3.6 $Y=2.355 $X2=0 $Y2=0
cc_262 N_A4_M1002_g N_VPWR_c_501_n 0.00291444f $X=3.6 $Y=2.355 $X2=0 $Y2=0
cc_263 N_A4_M1008_g N_VPWR_c_501_n 0.00291444f $X=4.03 $Y=2.355 $X2=0 $Y2=0
cc_264 N_A4_M1002_g N_VPWR_c_489_n 0.00428623f $X=3.6 $Y=2.355 $X2=0 $Y2=0
cc_265 N_A4_M1008_g N_VPWR_c_489_n 0.00399215f $X=4.03 $Y=2.355 $X2=0 $Y2=0
cc_266 N_A4_M1002_g N_A_652_345#_c_649_n 0.0109621f $X=3.6 $Y=2.355 $X2=0 $Y2=0
cc_267 N_A4_M1008_g N_A_652_345#_c_649_n 6.47031e-19 $X=4.03 $Y=2.355 $X2=0
+ $Y2=0
cc_268 N_A4_M1002_g N_A_652_345#_c_650_n 0.0101655f $X=3.6 $Y=2.355 $X2=0 $Y2=0
cc_269 N_A4_M1008_g N_A_652_345#_c_650_n 0.0117389f $X=4.03 $Y=2.355 $X2=0 $Y2=0
cc_270 N_A4_M1002_g N_A_652_345#_c_651_n 0.00233316f $X=3.6 $Y=2.355 $X2=0 $Y2=0
cc_271 N_A4_M1002_g N_A_652_345#_c_665_n 6.95406e-19 $X=3.6 $Y=2.355 $X2=0 $Y2=0
cc_272 N_A4_M1008_g N_A_652_345#_c_665_n 0.014865f $X=4.03 $Y=2.355 $X2=0 $Y2=0
cc_273 N_A4_M1008_g N_A_652_345#_c_653_n 0.00347585f $X=4.03 $Y=2.355 $X2=0
+ $Y2=0
cc_274 N_A4_c_305_n N_VGND_c_767_n 0.00357769f $X=3.6 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A4_c_307_n N_VGND_c_767_n 0.00211454f $X=4.03 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A4_c_307_n N_VGND_c_768_n 0.00585385f $X=4.03 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A4_c_305_n N_VGND_c_773_n 0.00585385f $X=3.6 $Y=1.185 $X2=0 $Y2=0
cc_278 N_A4_c_305_n N_VGND_c_779_n 0.0106551f $X=3.6 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A4_c_307_n N_VGND_c_779_n 0.0106551f $X=4.03 $Y=1.185 $X2=0 $Y2=0
cc_280 N_A4_c_305_n N_A_480_47#_c_886_n 0.0129873f $X=3.6 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A4_c_307_n N_A_480_47#_c_886_n 0.0138631f $X=4.03 $Y=1.185 $X2=0 $Y2=0
cc_282 A4 N_A_480_47#_c_886_n 0.0187087f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_283 N_A4_c_310_n N_A_480_47#_c_886_n 0.00252346f $X=4.03 $Y=1.35 $X2=0 $Y2=0
cc_284 A4 N_A_480_47#_c_887_n 0.00276452f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_285 N_A3_c_353_n N_A2_c_403_n 0.0145953f $X=4.89 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_286 A3 N_A2_c_405_n 0.00183669f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_287 N_A3_c_356_n N_A2_c_405_n 0.0236035f $X=4.89 $Y=1.35 $X2=0 $Y2=0
cc_288 A3 A2 0.019879f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_289 N_A3_M1014_g N_VPWR_c_501_n 0.00450424f $X=4.46 $Y=2.355 $X2=0 $Y2=0
cc_290 N_A3_M1027_g N_VPWR_c_501_n 0.0029147f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_291 N_A3_M1014_g N_VPWR_c_489_n 0.00862457f $X=4.46 $Y=2.355 $X2=0 $Y2=0
cc_292 N_A3_M1027_g N_VPWR_c_489_n 0.00428625f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_293 N_A3_M1014_g N_A_652_345#_c_650_n 0.00290301f $X=4.46 $Y=2.355 $X2=0
+ $Y2=0
cc_294 N_A3_M1014_g N_A_652_345#_c_665_n 0.0148657f $X=4.46 $Y=2.355 $X2=0 $Y2=0
cc_295 N_A3_M1027_g N_A_652_345#_c_665_n 7.03894e-19 $X=4.89 $Y=2.355 $X2=0
+ $Y2=0
cc_296 N_A3_M1014_g N_A_652_345#_c_652_n 0.01115f $X=4.46 $Y=2.355 $X2=0 $Y2=0
cc_297 N_A3_M1027_g N_A_652_345#_c_652_n 0.0143121f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_298 A3 N_A_652_345#_c_652_n 0.0574461f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_299 N_A3_c_356_n N_A_652_345#_c_652_n 0.00426203f $X=4.89 $Y=1.35 $X2=0 $Y2=0
cc_300 N_A3_M1014_g N_A_652_345#_c_653_n 0.00214624f $X=4.46 $Y=2.355 $X2=0
+ $Y2=0
cc_301 A3 N_A_652_345#_c_653_n 0.027718f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_302 N_A3_c_356_n N_A_652_345#_c_653_n 0.00179731f $X=4.89 $Y=1.35 $X2=0 $Y2=0
cc_303 N_A3_M1014_g N_A_652_345#_c_678_n 6.55518e-19 $X=4.46 $Y=2.355 $X2=0
+ $Y2=0
cc_304 N_A3_M1027_g N_A_652_345#_c_678_n 0.0113619f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_305 N_A3_M1027_g N_A_907_345#_c_699_n 0.0143655f $X=4.89 $Y=2.355 $X2=0 $Y2=0
cc_306 N_A3_M1014_g N_A_907_345#_c_700_n 7.3655e-19 $X=4.46 $Y=2.355 $X2=0 $Y2=0
cc_307 N_A3_M1027_g N_A_1108_367#_c_724_n 0.00141706f $X=4.89 $Y=2.355 $X2=0
+ $Y2=0
cc_308 N_A3_M1027_g N_A_1108_367#_c_726_n 3.95484e-19 $X=4.89 $Y=2.355 $X2=0
+ $Y2=0
cc_309 N_A3_c_351_n N_VGND_c_768_n 0.00585385f $X=4.46 $Y=1.185 $X2=0 $Y2=0
cc_310 N_A3_c_351_n N_VGND_c_769_n 0.00211189f $X=4.46 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A3_c_353_n N_VGND_c_769_n 0.00209041f $X=4.89 $Y=1.185 $X2=0 $Y2=0
cc_312 N_A3_c_351_n N_VGND_c_779_n 0.0106551f $X=4.46 $Y=1.185 $X2=0 $Y2=0
cc_313 N_A3_c_353_n N_VGND_c_779_n 0.0106687f $X=4.89 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A3_c_353_n N_VGND_c_782_n 0.00585385f $X=4.89 $Y=1.185 $X2=0 $Y2=0
cc_315 A3 N_A_480_47#_c_886_n 0.00867174f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_316 N_A3_c_351_n N_A_480_47#_c_900_n 0.0129934f $X=4.46 $Y=1.185 $X2=0 $Y2=0
cc_317 N_A3_c_353_n N_A_480_47#_c_900_n 0.0129934f $X=4.89 $Y=1.185 $X2=0 $Y2=0
cc_318 A3 N_A_480_47#_c_900_n 0.0371803f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_319 N_A3_c_356_n N_A_480_47#_c_900_n 0.00230884f $X=4.89 $Y=1.35 $X2=0 $Y2=0
cc_320 A3 N_A_480_47#_c_904_n 0.0174739f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_321 N_A3_c_356_n N_A_480_47#_c_904_n 0.00128991f $X=4.89 $Y=1.35 $X2=0 $Y2=0
cc_322 A3 N_A_480_47#_c_906_n 0.014701f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_323 N_A3_c_356_n N_A_480_47#_c_906_n 0.00139393f $X=4.89 $Y=1.35 $X2=0 $Y2=0
cc_324 N_A2_c_407_n N_A1_c_452_n 0.0145953f $X=6.24 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A2_M1021_g N_A1_M1005_g 0.0274522f $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_326 A2 A1 0.0198783f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_327 N_A2_c_409_n A1 0.00208709f $X=6.31 $Y=1.35 $X2=0 $Y2=0
cc_328 N_A2_c_409_n N_A1_c_457_n 0.0241566f $X=6.31 $Y=1.35 $X2=0 $Y2=0
cc_329 N_A2_M1021_g N_VPWR_c_495_n 0.00136666f $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A2_M1015_g N_VPWR_c_501_n 0.00357842f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A2_M1021_g N_VPWR_c_501_n 0.00547432f $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A2_M1015_g N_VPWR_c_489_n 0.00675085f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A2_M1021_g N_VPWR_c_489_n 0.00990114f $X=6.31 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_c_405_n N_A_652_345#_c_652_n 9.12731e-19 $X=5.395 $Y=1.35 $X2=0
+ $Y2=0
cc_335 N_A2_M1015_g N_A_652_345#_c_652_n 0.00311437f $X=5.88 $Y=2.465 $X2=0
+ $Y2=0
cc_336 N_A2_M1015_g N_A_652_345#_c_678_n 3.00735e-19 $X=5.88 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_A2_M1015_g N_A_907_345#_c_699_n 0.0129552f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_338 N_A2_M1015_g N_A_907_345#_c_704_n 6.12373e-19 $X=5.88 $Y=2.465 $X2=0
+ $Y2=0
cc_339 N_A2_M1021_g N_A_907_345#_c_704_n 0.00203265f $X=6.31 $Y=2.465 $X2=0
+ $Y2=0
cc_340 N_A2_M1015_g N_A_907_345#_c_706_n 0.0148052f $X=5.88 $Y=2.465 $X2=0 $Y2=0
cc_341 N_A2_M1021_g N_A_907_345#_c_706_n 0.00882136f $X=6.31 $Y=2.465 $X2=0
+ $Y2=0
cc_342 N_A2_c_404_n N_A_1108_367#_c_725_n 0.0010123f $X=5.805 $Y=1.35 $X2=0
+ $Y2=0
cc_343 N_A2_M1015_g N_A_1108_367#_c_725_n 0.0154606f $X=5.88 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A2_M1021_g N_A_1108_367#_c_725_n 0.0158554f $X=6.31 $Y=2.465 $X2=0
+ $Y2=0
cc_345 A2 N_A_1108_367#_c_725_n 0.0234234f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_346 N_A2_c_409_n N_A_1108_367#_c_725_n 0.00257059f $X=6.31 $Y=1.35 $X2=0
+ $Y2=0
cc_347 N_A2_c_404_n N_A_1108_367#_c_726_n 0.00631451f $X=5.805 $Y=1.35 $X2=0
+ $Y2=0
cc_348 A2 N_A_1108_367#_c_726_n 0.0151447f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_349 N_A2_c_407_n N_VGND_c_775_n 0.00585385f $X=6.24 $Y=1.185 $X2=0 $Y2=0
cc_350 N_A2_c_403_n N_VGND_c_779_n 0.0120521f $X=5.32 $Y=1.185 $X2=0 $Y2=0
cc_351 N_A2_c_407_n N_VGND_c_779_n 0.0120657f $X=6.24 $Y=1.185 $X2=0 $Y2=0
cc_352 N_A2_c_403_n N_VGND_c_782_n 0.00585385f $X=5.32 $Y=1.185 $X2=0 $Y2=0
cc_353 N_A2_c_403_n N_VGND_c_783_n 0.00567529f $X=5.32 $Y=1.185 $X2=0 $Y2=0
cc_354 N_A2_c_407_n N_VGND_c_783_n 0.00562637f $X=6.24 $Y=1.185 $X2=0 $Y2=0
cc_355 N_A2_c_403_n N_A_480_47#_c_908_n 0.0173661f $X=5.32 $Y=1.185 $X2=0 $Y2=0
cc_356 N_A2_c_404_n N_A_480_47#_c_908_n 0.0145729f $X=5.805 $Y=1.35 $X2=0 $Y2=0
cc_357 N_A2_c_407_n N_A_480_47#_c_908_n 0.0163763f $X=6.24 $Y=1.185 $X2=0 $Y2=0
cc_358 A2 N_A_480_47#_c_908_n 0.0586165f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_359 N_A2_c_409_n N_A_480_47#_c_912_n 0.00175003f $X=6.31 $Y=1.35 $X2=0 $Y2=0
cc_360 N_A1_M1005_g N_VPWR_c_495_n 0.0153689f $X=6.74 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A1_M1022_g N_VPWR_c_495_n 0.016151f $X=7.17 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A1_M1005_g N_VPWR_c_501_n 0.00486043f $X=6.74 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A1_M1022_g N_VPWR_c_502_n 0.00486043f $X=7.17 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A1_M1005_g N_VPWR_c_489_n 0.0082726f $X=6.74 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A1_M1022_g N_VPWR_c_489_n 0.00921135f $X=7.17 $Y=2.465 $X2=0 $Y2=0
cc_366 A1 N_A_1108_367#_c_725_n 0.00192505f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_367 N_A1_M1005_g N_A_1108_367#_c_727_n 0.0143687f $X=6.74 $Y=2.465 $X2=0
+ $Y2=0
cc_368 N_A1_M1022_g N_A_1108_367#_c_727_n 0.0153816f $X=7.17 $Y=2.465 $X2=0
+ $Y2=0
cc_369 A1 N_A_1108_367#_c_727_n 0.0460118f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_370 N_A1_c_457_n N_A_1108_367#_c_727_n 0.00425064f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_371 A1 N_A_1108_367#_c_728_n 0.0117399f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_372 N_A1_c_457_n N_A_1108_367#_c_728_n 7.12273e-19 $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_373 N_A1_c_452_n N_VGND_c_770_n 0.00211999f $X=6.67 $Y=1.185 $X2=0 $Y2=0
cc_374 N_A1_c_454_n N_VGND_c_770_n 0.00357769f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_375 N_A1_c_452_n N_VGND_c_775_n 0.00585385f $X=6.67 $Y=1.185 $X2=0 $Y2=0
cc_376 N_A1_c_454_n N_VGND_c_778_n 0.00585385f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_377 N_A1_c_452_n N_VGND_c_779_n 0.0106551f $X=6.67 $Y=1.185 $X2=0 $Y2=0
cc_378 N_A1_c_454_n N_VGND_c_779_n 0.0116476f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_379 N_A1_c_452_n N_A_480_47#_c_877_n 0.0129934f $X=6.67 $Y=1.185 $X2=0 $Y2=0
cc_380 N_A1_c_454_n N_A_480_47#_c_877_n 0.0129934f $X=7.1 $Y=1.185 $X2=0 $Y2=0
cc_381 A1 N_A_480_47#_c_877_n 0.0616108f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_382 N_A1_c_457_n N_A_480_47#_c_877_n 0.00460541f $X=7.1 $Y=1.35 $X2=0 $Y2=0
cc_383 A1 N_A_480_47#_c_912_n 0.0139141f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_384 N_VPWR_c_489_n N_X_M1006_s 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_489_n N_X_M1019_s 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_M1006_d N_X_c_596_n 2.33864e-19 $X=0.15 $Y=1.835 $X2=0 $Y2=0
cc_387 N_VPWR_c_491_n N_X_c_596_n 0.00362085f $X=0.275 $Y=2.18 $X2=0 $Y2=0
cc_388 N_VPWR_M1006_d N_X_c_597_n 0.00247068f $X=0.15 $Y=1.835 $X2=0 $Y2=0
cc_389 N_VPWR_c_491_n N_X_c_597_n 0.0203341f $X=0.275 $Y=2.18 $X2=0 $Y2=0
cc_390 N_VPWR_c_500_n N_X_c_629_n 0.0124525f $X=0.97 $Y=3.33 $X2=0 $Y2=0
cc_391 N_VPWR_c_489_n N_X_c_629_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_M1009_d N_X_c_598_n 0.00180746f $X=0.995 $Y=1.835 $X2=0 $Y2=0
cc_393 N_VPWR_c_492_n N_X_c_598_n 0.0163515f $X=1.135 $Y=2.19 $X2=0 $Y2=0
cc_394 N_VPWR_c_493_n N_X_c_598_n 0.00503283f $X=1.995 $Y=1.98 $X2=0 $Y2=0
cc_395 N_VPWR_c_496_n N_X_c_634_n 0.0124525f $X=1.83 $Y=3.33 $X2=0 $Y2=0
cc_396 N_VPWR_c_489_n N_X_c_634_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_397 N_VPWR_c_494_n N_A_652_345#_c_649_n 0.06831f $X=2.855 $Y=2.07 $X2=0 $Y2=0
cc_398 N_VPWR_c_501_n N_A_652_345#_c_650_n 0.0568424f $X=6.79 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_489_n N_A_652_345#_c_650_n 0.0313831f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_494_n N_A_652_345#_c_651_n 0.0134078f $X=2.855 $Y=2.07 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_501_n N_A_652_345#_c_651_n 0.0235688f $X=6.79 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_489_n N_A_652_345#_c_651_n 0.0127152f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_489_n N_A_907_345#_M1015_s 0.00223559f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_501_n N_A_907_345#_c_699_n 0.0722646f $X=6.79 $Y=3.33 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_489_n N_A_907_345#_c_699_n 0.042407f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_406 N_VPWR_c_501_n N_A_907_345#_c_700_n 0.0136205f $X=6.79 $Y=3.33 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_489_n N_A_907_345#_c_700_n 0.00738676f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_501_n N_A_907_345#_c_704_n 0.01906f $X=6.79 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_c_489_n N_A_907_345#_c_704_n 0.0124545f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_489_n N_A_1108_367#_M1015_d 0.0021598f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_411 N_VPWR_c_489_n N_A_1108_367#_M1021_d 0.00536646f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_489_n N_A_1108_367#_M1022_s 0.00444756f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_501_n N_A_1108_367#_c_748_n 0.0124525f $X=6.79 $Y=3.33 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_489_n N_A_1108_367#_c_748_n 0.00730901f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_415 N_VPWR_M1005_d N_A_1108_367#_c_727_n 0.00201607f $X=6.815 $Y=1.835 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_495_n N_A_1108_367#_c_727_n 0.013593f $X=6.955 $Y=2.19 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_502_n N_A_1108_367#_c_752_n 0.0135387f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_489_n N_A_1108_367#_c_752_n 0.00769778f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_419 N_X_c_591_n N_VGND_M1000_s 2.33864e-19 $X=0.61 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_420 N_X_c_594_n N_VGND_M1000_s 0.0021884f $X=0.21 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_421 N_X_c_592_n N_VGND_M1010_s 0.00176461f $X=1.47 $Y=1.14 $X2=0 $Y2=0
cc_422 N_X_c_591_n N_VGND_c_764_n 0.00362085f $X=0.61 $Y=1.14 $X2=0 $Y2=0
cc_423 N_X_c_594_n N_VGND_c_764_n 0.0203341f $X=0.21 $Y=1.225 $X2=0 $Y2=0
cc_424 N_X_c_592_n N_VGND_c_765_n 0.0170777f $X=1.47 $Y=1.14 $X2=0 $Y2=0
cc_425 N_X_c_592_n N_VGND_c_766_n 0.00276194f $X=1.47 $Y=1.14 $X2=0 $Y2=0
cc_426 N_X_c_643_p N_VGND_c_771_n 0.0124525f $X=1.565 $Y=0.42 $X2=0 $Y2=0
cc_427 N_X_c_644_p N_VGND_c_777_n 0.0124525f $X=0.705 $Y=0.42 $X2=0 $Y2=0
cc_428 N_X_M1000_d N_VGND_c_779_n 0.00536646f $X=0.565 $Y=0.245 $X2=0 $Y2=0
cc_429 N_X_M1011_d N_VGND_c_779_n 0.00536646f $X=1.425 $Y=0.245 $X2=0 $Y2=0
cc_430 N_X_c_644_p N_VGND_c_779_n 0.00730901f $X=0.705 $Y=0.42 $X2=0 $Y2=0
cc_431 N_X_c_643_p N_VGND_c_779_n 0.00730901f $X=1.565 $Y=0.42 $X2=0 $Y2=0
cc_432 N_A_652_345#_c_652_n N_A_907_345#_M1014_s 0.00176461f $X=4.94 $Y=1.69
+ $X2=-0.19 $Y2=1.655
cc_433 N_A_652_345#_c_652_n N_A_907_345#_c_716_n 0.0135055f $X=4.94 $Y=1.69
+ $X2=0 $Y2=0
cc_434 N_A_652_345#_M1027_d N_A_907_345#_c_699_n 0.00324607f $X=4.965 $Y=1.725
+ $X2=0 $Y2=0
cc_435 N_A_652_345#_c_678_n N_A_907_345#_c_699_n 0.0206016f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_436 N_A_652_345#_c_650_n N_A_907_345#_c_700_n 0.011362f $X=4.08 $Y=2.99 $X2=0
+ $Y2=0
cc_437 N_A_652_345#_c_678_n N_A_1108_367#_c_724_n 0.0548751f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_438 N_A_652_345#_c_652_n N_A_1108_367#_c_726_n 0.00520465f $X=4.94 $Y=1.69
+ $X2=0 $Y2=0
cc_439 N_A_652_345#_c_678_n N_A_1108_367#_c_726_n 0.00695919f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_440 N_A_652_345#_c_652_n N_A_480_47#_c_908_n 0.00100413f $X=4.94 $Y=1.69
+ $X2=0 $Y2=0
cc_441 N_A_652_345#_c_652_n N_A_480_47#_c_906_n 0.00145268f $X=4.94 $Y=1.69
+ $X2=0 $Y2=0
cc_442 N_A_907_345#_c_699_n N_A_1108_367#_M1015_d 0.00500911f $X=5.93 $Y=2.985
+ $X2=-0.19 $Y2=1.655
cc_443 N_A_907_345#_c_699_n N_A_1108_367#_c_724_n 0.0190318f $X=5.93 $Y=2.985
+ $X2=0 $Y2=0
cc_444 N_A_907_345#_M1015_s N_A_1108_367#_c_725_n 0.00180746f $X=5.955 $Y=1.835
+ $X2=0 $Y2=0
cc_445 N_A_907_345#_c_706_n N_A_1108_367#_c_725_n 0.0163515f $X=6.095 $Y=2.14
+ $X2=0 $Y2=0
cc_446 N_A_1108_367#_c_725_n N_A_480_47#_c_908_n 0.0020325f $X=6.43 $Y=1.79
+ $X2=0 $Y2=0
cc_447 N_A_1108_367#_c_725_n N_A_480_47#_c_912_n 0.0012179f $X=6.43 $Y=1.79
+ $X2=0 $Y2=0
cc_448 N_VGND_c_779_n N_A_480_47#_M1013_d 0.00215161f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_449 N_VGND_c_779_n N_A_480_47#_M1026_d 0.00254871f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_779_n N_A_480_47#_M1025_s 0.00293134f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_779_n N_A_480_47#_M1023_s 0.0027574f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_779_n N_A_480_47#_M1007_d 0.0027574f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_c_779_n N_A_480_47#_M1018_d 0.00266958f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_773_n N_A_480_47#_c_883_n 0.0499087f $X=3.685 $Y=0 $X2=0 $Y2=0
cc_455 N_VGND_c_779_n N_A_480_47#_c_883_n 0.0324982f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_456 N_VGND_M1024_d N_A_480_47#_c_886_n 0.00385462f $X=3.675 $Y=0.235 $X2=0
+ $Y2=0
cc_457 N_VGND_c_767_n N_A_480_47#_c_886_n 0.0135055f $X=3.815 $Y=0.535 $X2=0
+ $Y2=0
cc_458 N_VGND_c_768_n N_A_480_47#_c_932_n 0.0149362f $X=4.545 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_779_n N_A_480_47#_c_932_n 0.0100304f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_460 N_VGND_M1012_d N_A_480_47#_c_900_n 0.00329816f $X=4.535 $Y=0.235 $X2=0
+ $Y2=0
cc_461 N_VGND_c_769_n N_A_480_47#_c_900_n 0.0135055f $X=4.675 $Y=0.535 $X2=0
+ $Y2=0
cc_462 N_VGND_c_779_n N_A_480_47#_c_936_n 0.0102248f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_c_782_n N_A_480_47#_c_936_n 0.0151136f $X=5.405 $Y=0.307 $X2=0
+ $Y2=0
cc_464 N_VGND_M1003_s N_A_480_47#_c_908_n 0.0162231f $X=5.395 $Y=0.235 $X2=0
+ $Y2=0
cc_465 N_VGND_c_783_n N_A_480_47#_c_908_n 0.0531371f $X=6.15 $Y=0.307 $X2=0
+ $Y2=0
cc_466 N_VGND_c_775_n N_A_480_47#_c_940_n 0.0151136f $X=6.755 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_c_779_n N_A_480_47#_c_940_n 0.0102248f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_468 N_VGND_M1001_s N_A_480_47#_c_877_n 0.00329816f $X=6.745 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_VGND_c_770_n N_A_480_47#_c_877_n 0.0135055f $X=6.885 $Y=0.535 $X2=0
+ $Y2=0
cc_470 N_VGND_c_778_n N_A_480_47#_c_878_n 0.0192334f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_779_n N_A_480_47#_c_878_n 0.012111f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_766_n N_A_480_47#_c_879_n 0.0306103f $X=1.995 $Y=0.39 $X2=0
+ $Y2=0
cc_473 N_VGND_c_773_n N_A_480_47#_c_879_n 0.0172549f $X=3.685 $Y=0 $X2=0 $Y2=0
cc_474 N_VGND_c_779_n N_A_480_47#_c_879_n 0.00991703f $X=7.44 $Y=0 $X2=0 $Y2=0
