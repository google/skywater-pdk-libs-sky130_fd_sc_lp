* NGSPICE file created from sky130_fd_sc_lp__o221ai_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o221ai_m A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_148_47# C1 Y VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.113e+11p ps=1.37e+06u
M1001 VPWR A1 a_441_463# VPB phighvt w=420000u l=150000u
+  ad=2.943e+11p pd=3.13e+06u as=8.82e+10p ps=1.26e+06u
M1002 Y B2 a_245_480# VPB phighvt w=420000u l=150000u
+  ad=3.2995e+11p pd=3.32e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_234_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=2.415e+11p pd=2.83e+06u as=1.764e+11p ps=1.68e+06u
M1004 a_148_47# B2 a_234_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_234_47# B1 a_148_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C1 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_441_463# A2 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_234_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_245_480# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

