* File: sky130_fd_sc_lp__fa_0.spice
* Created: Fri Aug 28 10:34:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fa_0.pex.spice"
.subckt sky130_fd_sc_lp__fa_0  VNB VPB A B CIN COUT VPWR SUM VGND
* 
* VGND	VGND
* SUM	SUM
* VPWR	VPWR
* COUT	COUT
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1026 N_VGND_M1026_d N_A_80_225#_M1026_g N_COUT_M1026_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1003 A_224_119# N_A_M1003_g N_VGND_M1026_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002 A=0.063
+ P=1.14 MULT=1
MM1020 N_A_80_225#_M1020_d N_B_M1020_g A_224_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_382_119#_M1022_d N_CIN_M1022_g N_A_80_225#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=8.568 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_B_M1027_g N_A_382_119#_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.102125 AS=0.0672 PD=0.965 PS=0.74 NRD=18.564 NRS=2.856 M=1 R=2.8
+ SA=75001.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1023 N_A_382_119#_M1023_d N_A_M1023_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.102125 PD=1.37 PS=0.965 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_781_119#_M1002_d N_CIN_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_B_M1017_g N_A_781_119#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0588 PD=0.8 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1013 N_A_781_119#_M1013_d N_A_M1013_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0798 PD=0.7 PS=0.8 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1011 N_A_1059_119#_M1011_d N_A_80_225#_M1011_g N_A_781_119#_M1013_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 A_1145_119# N_CIN_M1012_g N_A_1059_119#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75002 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1014 A_1239_119# N_B_M1014_g A_1145_119# VNB NSHORT L=0.15 W=0.42 AD=0.09945
+ AS=0.0672 PD=1.08 PS=0.74 NRD=51.936 NRS=30 M=1 R=2.8 SA=75002.5 SB=75000.5
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g A_1239_119# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.09945 PD=0.7 PS=1.08 NRD=0 NRS=51.936 M=1 R=2.8 SA=75001.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_SUM_M1006_d N_A_1059_119#_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_80_225#_M1007_g N_COUT_M1007_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.1696 PD=1.24377 PS=1.81 NRD=16.9223 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1010 A_218_532# N_A_M1010_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.0880019 PD=0.66 PS=0.816226 NRD=30.4759 NRS=25.7873 M=1 R=2.8 SA=75000.7
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1025 N_A_80_225#_M1025_d N_B_M1025_g A_218_532# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=30.4759 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_404_532#_M1005_d N_CIN_M1005_g N_A_80_225#_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=21.0987 M=1 R=2.8
+ SA=75001.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_B_M1021_g N_A_404_532#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_404_532#_M1016_d N_A_M1016_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_781_457#_M1004_d N_CIN_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_B_M1018_g N_A_781_457#_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0588 PD=0.8 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1008 N_A_781_457#_M1008_d N_A_M1008_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0798 PD=0.7 PS=0.8 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_1059_119#_M1024_d N_A_80_225#_M1024_g N_A_781_457#_M1008_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=21.0987 NRS=0 M=1
+ R=2.8 SA=75001.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1019 A_1161_457# N_CIN_M1019_g N_A_1059_119#_M1024_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=30.4759 NRS=16.4101 M=1 R=2.8
+ SA=75002.1 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1009 A_1239_457# N_B_M1009_g A_1161_457# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0504 PD=0.81 PS=0.66 NRD=65.6601 NRS=30.4759 M=1 R=2.8 SA=75002.5
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g A_1239_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0905774 AS=0.0819 PD=0.820189 PS=0.81 NRD=46.886 NRS=65.6601 M=1 R=2.8
+ SA=75003 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_SUM_M1000_d N_A_1059_119#_M1000_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.138023 PD=1.81 PS=1.24981 NRD=0 NRS=6.1464 M=1 R=4.26667
+ SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.0319 P=19.85
c_80 VNB 0 8.70569e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__fa_0.pxi.spice"
*
.ends
*
*
