* NGSPICE file created from sky130_fd_sc_lp__dlxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
M1000 Q_N a_1266_147# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=1.6405e+12p ps=1.405e+07u
M1001 VGND a_758_359# a_748_47# VNB nshort w=420000u l=150000u
+  ad=1.0458e+12p pd=1.011e+07u as=8.82e+10p ps=1.26e+06u
M1002 VPWR D a_46_62# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1003 a_608_491# a_367_491# a_568_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=8.82e+10p ps=1.26e+06u
M1004 VGND a_758_359# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1005 a_536_491# a_46_62# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1006 VPWR a_758_359# a_713_491# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=9.45e+10p ps=1.29e+06u
M1007 a_568_47# a_46_62# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_215_62# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1009 a_758_359# a_608_491# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1010 VPWR a_215_62# a_367_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1011 a_713_491# a_367_491# a_608_491# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.158e+11p ps=2.03e+06u
M1012 a_1266_147# a_758_359# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1013 VGND a_215_62# a_367_491# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1014 Q_N a_1266_147# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1015 a_748_47# a_215_62# a_608_491# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1266_147# a_758_359# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1017 VPWR a_758_359# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1018 a_758_359# a_608_491# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1019 a_608_491# a_215_62# a_536_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_215_62# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1021 VGND D a_46_62# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

