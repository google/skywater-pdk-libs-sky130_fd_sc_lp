* File: sky130_fd_sc_lp__o311a_m.spice
* Created: Wed Sep  2 10:23:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311a_m.pex.spice"
.subckt sky130_fd_sc_lp__o311a_m  VNB VPB A1 A2 A3 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_93_153#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_250_47#_M1003_d N_A1_M1003_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_250_47#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_250_47#_M1010_d N_A3_M1010_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0588 PD=0.81 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1007 A_530_47# N_B1_M1007_g N_A_250_47#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=31.428 M=1 R=2.8 SA=75002
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_93_153#_M1001_d N_C1_M1001_g A_530_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_93_153#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09345 AS=0.1197 PD=0.865 PS=1.41 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1004 A_242_397# N_A1_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.09345 PD=0.63 PS=0.865 NRD=23.443 NRS=77.3816 M=1 R=2.8
+ SA=75000.8 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1000 A_314_397# N_A2_M1000_g A_242_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=65.6601 NRS=23.443 M=1 R=2.8 SA=75001.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_93_153#_M1005_d N_A3_M1005_g A_314_397# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=0 NRS=65.6601 M=1 R=2.8 SA=75001.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_A_93_153#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=51.5943 M=1 R=2.8 SA=75002.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_93_153#_M1006_d N_C1_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_84 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o311a_m.pxi.spice"
*
.ends
*
*
