# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux2_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__mux2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.815000 1.565000 5.145000 1.895000 ;
        RECT 4.975000 1.025000 7.095000 1.195000 ;
        RECT 4.975000 1.195000 5.145000 1.565000 ;
        RECT 6.765000 1.195000 7.095000 1.395000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.025000 4.805000 1.355000 ;
        RECT 4.475000 1.355000 4.645000 1.780000 ;
        RECT 6.355000 1.550000 6.595000 1.565000 ;
        RECT 6.355000 1.565000 7.095000 1.925000 ;
      LAYER mcon ;
        RECT 4.475000 1.580000 4.645000 1.750000 ;
        RECT 6.395000 1.580000 6.565000 1.750000 ;
      LAYER met1 ;
        RECT 4.415000 1.550000 4.705000 1.595000 ;
        RECT 4.415000 1.595000 6.625000 1.735000 ;
        RECT 4.415000 1.735000 4.705000 1.780000 ;
        RECT 6.335000 1.550000 6.625000 1.595000 ;
        RECT 6.335000 1.735000 6.625000 1.780000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.807000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.605000 4.305000 1.980000 ;
        RECT 3.965000 1.980000 4.565000 2.065000 ;
        RECT 3.965000 2.065000 5.685000 2.150000 ;
        RECT 4.395000 2.150000 5.685000 2.235000 ;
        RECT 5.355000 1.555000 5.685000 2.065000 ;
        RECT 7.805000 1.920000 8.035000 2.150000 ;
        RECT 7.865000 1.345000 8.370000 1.675000 ;
        RECT 7.865000 1.675000 8.035000 1.920000 ;
      LAYER mcon ;
        RECT 5.435000 1.950000 5.605000 2.120000 ;
        RECT 7.835000 1.950000 8.005000 2.120000 ;
      LAYER met1 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 1.965000 8.065000 2.105000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.295000 0.875000 0.925000 ;
        RECT 0.545000 0.925000 3.525000 1.095000 ;
        RECT 0.545000 1.095000 0.875000 1.815000 ;
        RECT 0.545000 1.815000 3.375000 1.985000 ;
        RECT 0.545000 1.985000 0.875000 3.075000 ;
        RECT 1.405000 0.295000 1.735000 0.925000 ;
        RECT 1.405000 1.985000 1.735000 3.075000 ;
        RECT 2.265000 0.295000 2.595000 0.925000 ;
        RECT 2.265000 1.985000 2.595000 3.075000 ;
        RECT 3.125000 1.985000 3.375000 3.075000 ;
        RECT 3.195000 0.295000 3.525000 0.925000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.640000 0.085000 ;
        RECT 0.115000  0.085000 0.375000 1.115000 ;
        RECT 1.055000  0.085000 1.225000 0.755000 ;
        RECT 1.915000  0.085000 2.085000 0.755000 ;
        RECT 2.775000  0.085000 3.025000 0.755000 ;
        RECT 3.705000  0.085000 3.955000 1.095000 ;
        RECT 5.680000  0.085000 6.010000 0.515000 ;
        RECT 7.665000  0.085000 7.995000 0.835000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.640000 3.415000 ;
        RECT 0.115000 1.795000 0.365000 3.245000 ;
        RECT 1.055000 2.155000 1.225000 3.245000 ;
        RECT 1.915000 2.155000 2.085000 3.245000 ;
        RECT 2.775000 2.155000 2.945000 3.245000 ;
        RECT 3.555000 2.660000 3.885000 3.245000 ;
        RECT 5.690000 2.775000 6.020000 3.245000 ;
        RECT 7.745000 2.660000 8.075000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.120000 1.265000 4.305000 1.435000 ;
      RECT 1.120000 1.435000 3.795000 1.595000 ;
      RECT 3.625000 1.595000 3.795000 2.320000 ;
      RECT 3.625000 2.320000 4.225000 2.405000 ;
      RECT 3.625000 2.405000 5.860000 2.435000 ;
      RECT 3.625000 2.435000 7.020000 2.490000 ;
      RECT 4.055000 2.490000 7.020000 2.575000 ;
      RECT 4.135000 0.685000 6.950000 0.855000 ;
      RECT 4.135000 0.855000 4.305000 1.265000 ;
      RECT 4.170000 0.255000 5.500000 0.425000 ;
      RECT 4.170000 0.425000 4.500000 0.515000 ;
      RECT 4.190000 2.745000 4.520000 2.905000 ;
      RECT 4.190000 2.905000 5.520000 3.075000 ;
      RECT 4.670000 0.595000 5.000000 0.685000 ;
      RECT 4.690000 2.575000 5.020000 2.735000 ;
      RECT 5.170000 0.425000 5.500000 0.515000 ;
      RECT 5.190000 2.745000 5.520000 2.905000 ;
      RECT 5.690000 2.575000 7.020000 2.605000 ;
      RECT 5.895000 1.555000 6.185000 2.095000 ;
      RECT 5.895000 2.095000 7.535000 2.235000 ;
      RECT 6.030000 2.235000 7.535000 2.265000 ;
      RECT 6.190000 0.295000 7.450000 0.465000 ;
      RECT 6.190000 2.775000 6.520000 2.905000 ;
      RECT 6.190000 2.905000 7.520000 3.075000 ;
      RECT 6.620000 0.635000 6.950000 0.685000 ;
      RECT 6.690000 2.605000 7.020000 2.735000 ;
      RECT 7.120000 0.465000 7.450000 0.835000 ;
      RECT 7.190000 2.660000 7.520000 2.905000 ;
      RECT 7.365000 1.005000 8.495000 1.175000 ;
      RECT 7.365000 1.175000 7.695000 1.515000 ;
      RECT 7.365000 1.515000 7.535000 2.095000 ;
      RECT 7.365000 2.265000 7.535000 2.320000 ;
      RECT 7.365000 2.320000 8.505000 2.490000 ;
      RECT 8.165000 0.255000 8.495000 1.005000 ;
      RECT 8.255000 1.845000 8.505000 2.320000 ;
      RECT 8.255000 2.490000 8.505000 3.075000 ;
  END
END sky130_fd_sc_lp__mux2_8
