* File: sky130_fd_sc_lp__nor3b_1.spice
* Created: Fri Aug 28 10:56:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor3b_1.pex.spice"
.subckt sky130_fd_sc_lp__nor3b_1  VNB VPB C_N A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_C_N_M1000_g N_A_82_131#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0931 AS=0.1113 PD=0.826667 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84 AD=0.1323
+ AS=0.1862 PD=1.155 PS=1.65333 NRD=4.992 NRS=8.568 M=1 R=5.6 SA=75000.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.84 AD=0.1197
+ AS=0.1323 PD=1.125 PS=1.155 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_82_131#_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1197 PD=2.21 PS=1.125 NRD=0 NRS=0.708 M=1 R=5.6 SA=75001.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_C_N_M1004_g N_A_82_131#_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09765 AS=0.1113 PD=0.83 PS=1.37 NRD=83.2522 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1006 A_275_367# N_A_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.29295 PD=1.47 PS=2.49 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.4 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1007 A_347_367# N_B_M1007_g A_275_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75000.7
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_82_131#_M1001_g A_347_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3528 AS=0.2457 PD=3.08 PS=1.65 NRD=2.3443 NRS=21.8867 M=1 R=8.4
+ SA=75001.3 SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__nor3b_1.pxi.spice"
*
.ends
*
*
