* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
X0 a_531_423# a_587_350# a_286_423# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1789_141# a_872_324# a_1865_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND DE a_120_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_902_396# a_1067_65# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 VPWR a_120_179# a_459_423# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_286_423# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_231_53# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_872_324# a_958_290# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_120_179# a_404_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1865_367# a_958_290# a_1971_388# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1986_57# a_1067_65# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_1781_367# a_872_324# a_1865_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_902_396# a_958_290# a_1004_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1865_367# a_958_290# a_1986_57# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VGND a_587_350# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_531_423# a_587_350# a_404_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_459_423# D a_531_423# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VGND a_587_350# a_1789_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_902_396# a_958_290# a_531_423# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_761_396# a_872_324# a_902_396# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VPWR a_587_350# a_1971_388# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR a_587_350# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_761_396# a_1067_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_872_324# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_587_350# a_1865_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_231_53# D a_531_423# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_531_423# a_872_324# a_902_396# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VGND a_902_396# a_1067_65# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 VGND a_1865_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 VPWR DE a_120_179# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 VPWR a_1865_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 VPWR a_872_324# a_958_290# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 a_1781_367# a_1067_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_872_324# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_587_350# a_1865_367# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1004_91# a_1067_65# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
