* NGSPICE file created from sky130_fd_sc_lp__mux2i_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__mux2i_m A0 A1 S VGND VNB VPB VPWR Y
M1000 VGND S a_416_125# VNB nshort w=420000u l=150000u
+  ad=2.751e+11p pd=2.99e+06u as=1.659e+11p ps=1.63e+06u
M1001 Y A1 a_256_497# VPB phighvt w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=8.82e+10p ps=1.26e+06u
M1002 a_452_497# A0 Y VPB phighvt w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1003 VPWR S a_452_497# VPB phighvt w=420000u l=150000u
+  ad=3.024e+11p pd=3.12e+06u as=0p ps=0u
M1004 VGND S a_55_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1005 VPWR S a_55_125# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 a_256_497# a_55_125# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A0 a_250_125# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=8.82e+10p ps=1.26e+06u
M1008 a_250_125# a_55_125# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_416_125# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

