* File: sky130_fd_sc_lp__and4_2.pex.spice
* Created: Fri Aug 28 10:07:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4_2%A 2 5 9 11 12 13 17 18
r31 17 19 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.17
+ $X2=0.597 $Y2=1.005
r32 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.17 $X2=0.585 $Y2=1.17
r33 12 13 7.56494 $w=5.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.377 $Y=1.295
+ $X2=0.377 $Y2=1.665
r34 12 18 2.55572 $w=5.83e-07 $l=1.25e-07 $layer=LI1_cond $X=0.377 $Y=1.295
+ $X2=0.377 $Y2=1.17
r35 9 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.7 $Y=2.045 $X2=0.7
+ $Y2=1.675
r36 5 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.7 $Y=0.455 $X2=0.7
+ $Y2=1.005
r37 2 11 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.597 $Y=1.498
+ $X2=0.597 $Y2=1.675
r38 1 17 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.597 $Y=1.182
+ $X2=0.597 $Y2=1.17
r39 1 2 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.597 $Y=1.182
+ $X2=0.597 $Y2=1.498
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_2%B 3 7 11 12 13 16
r40 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.09 $X2=1.15 $Y2=1.09
r41 13 17 1.17263 $w=5.08e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.26 $X2=1.15
+ $Y2=1.26
r42 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.15 $Y=1.43
+ $X2=1.15 $Y2=1.09
r43 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.43
+ $X2=1.15 $Y2=1.595
r44 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=0.925
+ $X2=1.15 $Y2=1.09
r45 7 12 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.13 $Y=2.045
+ $X2=1.13 $Y2=1.595
r46 3 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.06 $Y=0.455 $X2=1.06
+ $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_2%C 3 7 11 12 13 16 17
r36 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.09 $X2=1.69 $Y2=1.09
r37 13 17 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.69 $Y=1.295
+ $X2=1.69 $Y2=1.09
r38 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=1.43
+ $X2=1.69 $Y2=1.09
r39 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.43
+ $X2=1.69 $Y2=1.595
r40 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=0.925
+ $X2=1.69 $Y2=1.09
r41 7 12 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.78 $Y=2.045
+ $X2=1.78 $Y2=1.595
r42 3 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.6 $Y=0.455 $X2=1.6
+ $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_2%D 3 7 11 12 13 16 17
r40 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.09 $X2=2.23 $Y2=1.09
r41 13 17 1.64168 $w=5.08e-07 $l=7e-08 $layer=LI1_cond $X=2.16 $Y=1.26 $X2=2.23
+ $Y2=1.26
r42 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=1.43
+ $X2=2.23 $Y2=1.09
r43 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.43
+ $X2=2.23 $Y2=1.595
r44 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=0.925
+ $X2=2.23 $Y2=1.09
r45 7 12 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.21 $Y=2.045
+ $X2=2.21 $Y2=1.595
r46 3 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.14 $Y=0.455 $X2=2.14
+ $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_2%A_72_49# 1 2 3 12 16 20 24 28 30 31 32 36 38
+ 43 45 48 52
c101 43 0 1.0248e-19 $X=2.77 $Y=1.51
r102 51 52 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.905 $Y=1.51
+ $X2=3.335 $Y2=1.51
r103 45 47 15.3108 $w=2.51e-07 $l=3.15e-07 $layer=LI1_cond $X=0.95 $Y=1.77
+ $X2=0.95 $Y2=2.085
r104 44 51 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.77 $Y=1.51
+ $X2=2.905 $Y2=1.51
r105 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.51 $X2=2.77 $Y2=1.51
r106 41 43 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=2.73 $Y=1.685
+ $X2=2.73 $Y2=1.51
r107 40 43 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.73 $Y=0.835
+ $X2=2.73 $Y2=1.51
r108 39 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.09 $Y=1.77
+ $X2=1.96 $Y2=1.77
r109 38 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.605 $Y=1.77
+ $X2=2.73 $Y2=1.685
r110 38 39 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.605 $Y=1.77
+ $X2=2.09 $Y2=1.77
r111 34 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=1.855
+ $X2=1.96 $Y2=1.77
r112 34 36 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=1.96 $Y=1.855
+ $X2=1.96 $Y2=2.045
r113 33 45 3.01842 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.08 $Y=1.77
+ $X2=0.95 $Y2=1.77
r114 32 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.83 $Y=1.77
+ $X2=1.96 $Y2=1.77
r115 32 33 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.83 $Y=1.77
+ $X2=1.08 $Y2=1.77
r116 30 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.605 $Y=0.75
+ $X2=2.73 $Y2=0.835
r117 30 31 127.545 $w=1.68e-07 $l=1.955e-06 $layer=LI1_cond $X=2.605 $Y=0.75
+ $X2=0.65 $Y2=0.75
r118 26 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.485 $Y=0.665
+ $X2=0.65 $Y2=0.75
r119 26 28 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.485 $Y=0.665
+ $X2=0.485 $Y2=0.455
r120 22 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=1.675
+ $X2=3.335 $Y2=1.51
r121 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.335 $Y=1.675
+ $X2=3.335 $Y2=2.465
r122 18 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=1.345
+ $X2=3.335 $Y2=1.51
r123 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.335 $Y=1.345
+ $X2=3.335 $Y2=0.665
r124 14 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.675
+ $X2=2.905 $Y2=1.51
r125 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.905 $Y=1.675
+ $X2=2.905 $Y2=2.465
r126 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.345
+ $X2=2.905 $Y2=1.51
r127 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.905 $Y=1.345
+ $X2=2.905 $Y2=0.665
r128 3 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=2.045
r129 2 47 600 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.775
+ $Y=1.835 $X2=0.915 $Y2=2.085
r130 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.36
+ $Y=0.245 $X2=0.485 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_2%VPWR 1 2 3 4 15 19 23 27 29 34 35 37 38 39 48
+ 52 58 62
r41 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 56 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 56 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 53 58 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.557 $Y2=3.33
r47 53 55 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 52 61 4.34925 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.632 $Y2=3.33
r49 52 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 51 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 48 58 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.557 $Y2=3.33
r53 48 50 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.26 $Y=3.33 $X2=2.16
+ $Y2=3.33
r54 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 43 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 39 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 39 47 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 37 46 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.28 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=3.33
+ $X2=1.445 $Y2=3.33
r61 36 50 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.445 $Y2=3.33
r63 34 42 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.32 $Y=3.33 $X2=0.24
+ $Y2=3.33
r64 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=3.33
+ $X2=0.485 $Y2=3.33
r65 33 46 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.65 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=3.33
+ $X2=0.485 $Y2=3.33
r67 29 32 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=3.57 $Y=1.98
+ $X2=3.57 $Y2=2.95
r68 27 61 3.0886 $w=2.9e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.632 $Y2=3.33
r69 27 32 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=2.95
r70 23 26 7.73933 $w=5.93e-07 $l=3.85e-07 $layer=LI1_cond $X=2.557 $Y=2.11
+ $X2=2.557 $Y2=2.495
r71 21 58 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.557 $Y=3.245
+ $X2=2.557 $Y2=3.33
r72 21 26 15.0766 $w=5.93e-07 $l=7.5e-07 $layer=LI1_cond $X=2.557 $Y=3.245
+ $X2=2.557 $Y2=2.495
r73 17 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=3.245
+ $X2=1.445 $Y2=3.33
r74 17 19 39.6371 $w=3.28e-07 $l=1.135e-06 $layer=LI1_cond $X=1.445 $Y=3.245
+ $X2=1.445 $Y2=2.11
r75 13 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.485 $Y=3.245
+ $X2=0.485 $Y2=3.33
r76 13 15 41.907 $w=3.28e-07 $l=1.2e-06 $layer=LI1_cond $X=0.485 $Y=3.245
+ $X2=0.485 $Y2=2.045
r77 4 32 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.835 $X2=3.55 $Y2=2.95
r78 4 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.835 $X2=3.55 $Y2=1.98
r79 3 26 300 $w=1.7e-07 $l=8.38391e-07 $layer=licon1_PDIFF $count=2 $X=2.285
+ $Y=1.835 $X2=2.69 $Y2=2.495
r80 3 23 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.425 $Y2=2.11
r81 2 19 600 $w=1.7e-07 $l=3.76331e-07 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.835 $X2=1.445 $Y2=2.11
r82 1 15 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.36
+ $Y=1.835 $X2=0.485 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_2%X 1 2 7 8 9 10 11 12 13 22
r17 13 40 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.14 $Y=2.775
+ $X2=3.14 $Y2=2.91
r18 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=2.405
+ $X2=3.14 $Y2=2.775
r19 11 12 21.2951 $w=2.28e-07 $l=4.25e-07 $layer=LI1_cond $X=3.14 $Y=1.98
+ $X2=3.14 $Y2=2.405
r20 10 11 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.14 $Y=1.665
+ $X2=3.14 $Y2=1.98
r21 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.665
r22 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=0.925 $X2=3.14
+ $Y2=1.295
r23 7 8 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=0.555 $X2=3.14
+ $Y2=0.925
r24 7 22 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.14 $Y=0.555
+ $X2=3.14 $Y2=0.42
r25 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.835 $X2=3.12 $Y2=2.91
r26 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.835 $X2=3.12 $Y2=1.98
r27 1 22 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.98
+ $Y=0.245 $X2=3.12 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_2%VGND 1 2 9 11 13 16 17 18 27 33
r38 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r39 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r40 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 27 32 4.34925 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.632
+ $Y2=0
r42 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.12
+ $Y2=0
r43 26 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r44 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r45 21 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r46 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 18 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r48 18 22 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.24
+ $Y2=0
r49 16 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.16
+ $Y2=0
r50 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.525
+ $Y2=0
r51 15 29 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=3.12
+ $Y2=0
r52 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.525
+ $Y2=0
r53 11 32 3.0886 $w=2.9e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.632 $Y2=0
r54 11 13 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.39
r55 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0
r56 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0.39
r57 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.245 $X2=3.55 $Y2=0.39
r58 1 9 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.245 $X2=2.525 $Y2=0.39
.ends

