* File: sky130_fd_sc_lp__and2b_2.pxi.spice
* Created: Wed Sep  2 09:31:01 2020
* 
x_PM_SKY130_FD_SC_LP__AND2B_2%A_N N_A_N_M1006_g N_A_N_M1004_g A_N A_N
+ N_A_N_c_61_n N_A_N_c_62_n PM_SKY130_FD_SC_LP__AND2B_2%A_N
x_PM_SKY130_FD_SC_LP__AND2B_2%A_186_239# N_A_186_239#_M1005_d
+ N_A_186_239#_M1003_d N_A_186_239#_M1000_g N_A_186_239#_c_89_n
+ N_A_186_239#_M1002_g N_A_186_239#_M1001_g N_A_186_239#_M1008_g
+ N_A_186_239#_c_91_n N_A_186_239#_c_92_n N_A_186_239#_c_93_n
+ N_A_186_239#_c_102_n N_A_186_239#_c_103_n N_A_186_239#_c_94_n
+ N_A_186_239#_c_95_n N_A_186_239#_c_96_n N_A_186_239#_c_97_n
+ PM_SKY130_FD_SC_LP__AND2B_2%A_186_239#
x_PM_SKY130_FD_SC_LP__AND2B_2%B N_B_M1003_g N_B_M1009_g B B N_B_c_174_n
+ N_B_c_175_n PM_SKY130_FD_SC_LP__AND2B_2%B
x_PM_SKY130_FD_SC_LP__AND2B_2%A_28_367# N_A_28_367#_M1004_s N_A_28_367#_M1006_s
+ N_A_28_367#_M1005_g N_A_28_367#_M1007_g N_A_28_367#_c_213_n
+ N_A_28_367#_c_214_n N_A_28_367#_c_215_n N_A_28_367#_c_216_n
+ N_A_28_367#_c_220_n N_A_28_367#_c_217_n PM_SKY130_FD_SC_LP__AND2B_2%A_28_367#
x_PM_SKY130_FD_SC_LP__AND2B_2%VPWR N_VPWR_M1006_d N_VPWR_M1001_d N_VPWR_M1007_d
+ N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n VPWR
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_269_n N_VPWR_c_278_n
+ N_VPWR_c_279_n N_VPWR_c_280_n PM_SKY130_FD_SC_LP__AND2B_2%VPWR
x_PM_SKY130_FD_SC_LP__AND2B_2%X N_X_M1002_s N_X_M1000_s N_X_c_302_n X X X X X
+ PM_SKY130_FD_SC_LP__AND2B_2%X
x_PM_SKY130_FD_SC_LP__AND2B_2%VGND N_VGND_M1004_d N_VGND_M1008_d N_VGND_c_326_n
+ N_VGND_c_327_n VGND N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n
+ PM_SKY130_FD_SC_LP__AND2B_2%VGND
cc_1 VNB N_A_N_M1006_g 0.00623951f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.045
cc_2 VNB A_N 0.00810002f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_61_n 0.033098f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_4 VNB N_A_N_c_62_n 0.0206187f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.21
cc_5 VNB N_A_186_239#_M1000_g 0.00854382f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_A_186_239#_c_89_n 0.0184547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_186_239#_M1008_g 0.0271515f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.375
cc_8 VNB N_A_186_239#_c_91_n 8.22047e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_186_239#_c_92_n 0.0527582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_186_239#_c_93_n 0.00808088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_186_239#_c_94_n 0.00521995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_186_239#_c_95_n 0.0330429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_186_239#_c_96_n 0.00167923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_186_239#_c_97_n 0.0194624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1003_g 0.00681804f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.045
cc_16 VNB B 0.0111861f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_B_c_174_n 0.0296069f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_18 VNB N_B_c_175_n 0.0167171f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.21
cc_19 VNB N_A_28_367#_M1005_g 0.0147438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_28_367#_M1007_g 0.0175016f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_21 VNB N_A_28_367#_c_213_n 0.0103904f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.54
cc_22 VNB N_A_28_367#_c_214_n 0.0296923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_28_367#_c_215_n 0.0225285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_28_367#_c_216_n 0.0263246f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.665
cc_25 VNB N_A_28_367#_c_217_n 0.0466779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_269_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_302_n 0.00484367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.00509885f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_29 VNB N_VGND_c_326_n 0.0123607f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_30 VNB N_VGND_c_327_n 0.0182193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_328_n 0.0354643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_329_n 0.205758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_330_n 0.0375842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A_N_M1006_g 0.0296729f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.045
cc_35 VPB A_N 0.00567575f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_36 VPB N_A_186_239#_M1000_g 0.0232636f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_37 VPB N_A_186_239#_M1001_g 0.0213337f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.54
cc_38 VPB N_A_186_239#_c_92_n 0.0078604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_186_239#_c_93_n 0.00443634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_186_239#_c_102_n 0.00208455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_186_239#_c_103_n 6.98108e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_186_239#_c_94_n 0.0207772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_B_M1003_g 0.0243661f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.045
cc_44 VPB N_A_28_367#_M1007_g 0.0272785f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.375
cc_45 VPB N_A_28_367#_c_214_n 0.0117787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_28_367#_c_220_n 0.0132504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_270_n 0.0342452f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.375
cc_48 VPB N_VPWR_c_271_n 0.019861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_272_n 0.016802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_273_n 0.0646812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_274_n 0.0212365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_275_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_276_n 0.0155085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_269_n 0.0998106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_278_n 0.00612923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_279_n 0.0102056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_280_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB X 0.00377612f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.375
cc_59 N_A_N_M1006_g N_A_186_239#_M1000_g 0.0159868f $X=0.48 $Y=2.045 $X2=0 $Y2=0
cc_60 N_A_N_c_62_n N_A_186_239#_c_89_n 0.0162792f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_61 A_N N_A_186_239#_c_92_n 0.00517551f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A_N_c_61_n N_A_186_239#_c_92_n 0.0174182f $X=0.525 $Y=1.375 $X2=0 $Y2=0
cc_63 N_A_N_c_62_n N_A_186_239#_c_92_n 6.55063e-19 $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A_N_M1006_g N_A_28_367#_c_214_n 0.00890363f $X=0.48 $Y=2.045 $X2=0 $Y2=0
cc_65 A_N N_A_28_367#_c_214_n 0.0419357f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A_N_c_61_n N_A_28_367#_c_214_n 0.00808178f $X=0.525 $Y=1.375 $X2=0 $Y2=0
cc_67 N_A_N_c_62_n N_A_28_367#_c_214_n 0.00459057f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_68 A_N N_A_28_367#_c_215_n 0.0135954f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_N_c_62_n N_A_28_367#_c_215_n 0.0107043f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_70 A_N N_A_28_367#_c_216_n 0.00438436f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_N_c_61_n N_A_28_367#_c_216_n 0.00384498f $X=0.525 $Y=1.375 $X2=0 $Y2=0
cc_72 N_A_N_c_62_n N_A_28_367#_c_216_n 0.00956965f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_N_M1006_g N_A_28_367#_c_220_n 0.00508365f $X=0.48 $Y=2.045 $X2=0 $Y2=0
cc_74 N_A_N_M1006_g N_VPWR_c_270_n 0.00368396f $X=0.48 $Y=2.045 $X2=0 $Y2=0
cc_75 A_N N_VPWR_c_270_n 0.0262547f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_N_c_61_n N_VPWR_c_270_n 4.09642e-19 $X=0.525 $Y=1.375 $X2=0 $Y2=0
cc_77 N_A_N_c_62_n N_X_c_302_n 0.00141298f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_78 A_N X 0.0458946f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_N_c_62_n X 0.00106591f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A_N_c_62_n N_VGND_c_329_n 0.0044629f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_N_c_62_n N_VGND_c_330_n 0.00292942f $X=0.525 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_186_239#_M1001_g N_B_M1003_g 0.00866908f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_186_239#_c_91_n N_B_M1003_g 6.04156e-19 $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_84 N_A_186_239#_c_92_n N_B_M1003_g 0.0060897f $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_85 N_A_186_239#_c_93_n N_B_M1003_g 0.0148844f $X=2.25 $Y=1.71 $X2=0 $Y2=0
cc_86 N_A_186_239#_c_103_n N_B_M1003_g 0.00101119f $X=2.345 $Y=2.045 $X2=0 $Y2=0
cc_87 N_A_186_239#_M1008_g B 5.70717e-19 $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_88 N_A_186_239#_c_91_n B 0.00719646f $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_89 N_A_186_239#_c_92_n B 4.39421e-19 $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_90 N_A_186_239#_c_93_n B 0.0218791f $X=2.25 $Y=1.71 $X2=0 $Y2=0
cc_91 N_A_186_239#_c_94_n B 0.0217213f $X=2.905 $Y=1.71 $X2=0 $Y2=0
cc_92 N_A_186_239#_c_95_n B 0.0219735f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_93 N_A_186_239#_c_96_n B 0.0162075f $X=2.345 $Y=1.71 $X2=0 $Y2=0
cc_94 N_A_186_239#_c_97_n B 0.00738076f $X=3.032 $Y=0.877 $X2=0 $Y2=0
cc_95 N_A_186_239#_M1008_g N_B_c_174_n 0.00688898f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_96 N_A_186_239#_c_91_n N_B_c_174_n 6.46921e-19 $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_97 N_A_186_239#_c_92_n N_B_c_174_n 0.0122859f $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_98 N_A_186_239#_c_93_n N_B_c_174_n 0.00396368f $X=2.25 $Y=1.71 $X2=0 $Y2=0
cc_99 N_A_186_239#_c_96_n N_B_c_174_n 7.36548e-19 $X=2.345 $Y=1.71 $X2=0 $Y2=0
cc_100 N_A_186_239#_M1008_g N_B_c_175_n 0.0193329f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_101 N_A_186_239#_c_97_n N_B_c_175_n 0.00151061f $X=3.032 $Y=0.877 $X2=0 $Y2=0
cc_102 N_A_186_239#_c_95_n N_A_28_367#_M1005_g 0.0044767f $X=3.032 $Y=1.625
+ $X2=0 $Y2=0
cc_103 N_A_186_239#_c_97_n N_A_28_367#_M1005_g 0.00621676f $X=3.032 $Y=0.877
+ $X2=0 $Y2=0
cc_104 N_A_186_239#_c_103_n N_A_28_367#_M1007_g 0.00101119f $X=2.345 $Y=2.045
+ $X2=0 $Y2=0
cc_105 N_A_186_239#_c_94_n N_A_28_367#_M1007_g 0.0158751f $X=2.905 $Y=1.71 $X2=0
+ $Y2=0
cc_106 N_A_186_239#_c_95_n N_A_28_367#_M1007_g 0.00612008f $X=3.032 $Y=1.625
+ $X2=0 $Y2=0
cc_107 N_A_186_239#_c_95_n N_A_28_367#_c_213_n 0.0010809f $X=3.032 $Y=1.625
+ $X2=0 $Y2=0
cc_108 N_A_186_239#_c_89_n N_A_28_367#_c_215_n 0.0121074f $X=1.18 $Y=1.195 $X2=0
+ $Y2=0
cc_109 N_A_186_239#_M1008_g N_A_28_367#_c_215_n 0.0185176f $X=1.61 $Y=0.665
+ $X2=0 $Y2=0
cc_110 N_A_186_239#_c_91_n N_A_28_367#_c_215_n 0.00368472f $X=1.57 $Y=1.51 $X2=0
+ $Y2=0
cc_111 N_A_186_239#_c_92_n N_A_28_367#_c_215_n 0.00424322f $X=1.57 $Y=1.51 $X2=0
+ $Y2=0
cc_112 N_A_186_239#_c_97_n N_A_28_367#_c_215_n 0.0129811f $X=3.032 $Y=0.877
+ $X2=0 $Y2=0
cc_113 N_A_186_239#_c_89_n N_A_28_367#_c_216_n 9.59264e-19 $X=1.18 $Y=1.195
+ $X2=0 $Y2=0
cc_114 N_A_186_239#_c_97_n N_A_28_367#_c_217_n 0.00109491f $X=3.032 $Y=0.877
+ $X2=0 $Y2=0
cc_115 N_A_186_239#_M1000_g N_VPWR_c_270_n 0.00696463f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_186_239#_M1000_g N_VPWR_c_271_n 7.88315e-19 $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_186_239#_M1001_g N_VPWR_c_271_n 0.0249753f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_186_239#_c_92_n N_VPWR_c_271_n 0.00117518f $X=1.57 $Y=1.51 $X2=0
+ $Y2=0
cc_119 N_A_186_239#_c_93_n N_VPWR_c_271_n 0.0256507f $X=2.25 $Y=1.71 $X2=0 $Y2=0
cc_120 N_A_186_239#_c_102_n N_VPWR_c_271_n 0.0194526f $X=1.735 $Y=1.71 $X2=0
+ $Y2=0
cc_121 N_A_186_239#_c_94_n N_VPWR_c_273_n 0.0247108f $X=2.905 $Y=1.71 $X2=0
+ $Y2=0
cc_122 N_A_186_239#_M1000_g N_VPWR_c_275_n 0.00585385f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_186_239#_M1001_g N_VPWR_c_275_n 0.00486043f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_186_239#_M1000_g N_VPWR_c_269_n 0.0118221f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_186_239#_M1001_g N_VPWR_c_269_n 0.00824727f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_126 N_A_186_239#_c_89_n N_X_c_302_n 0.00811314f $X=1.18 $Y=1.195 $X2=0 $Y2=0
cc_127 N_A_186_239#_M1008_g N_X_c_302_n 0.00651662f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_128 N_A_186_239#_c_91_n N_X_c_302_n 0.00475211f $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A_186_239#_c_92_n N_X_c_302_n 0.00419321f $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A_186_239#_M1000_g X 0.00494518f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_186_239#_c_89_n X 0.00223387f $X=1.18 $Y=1.195 $X2=0 $Y2=0
cc_132 N_A_186_239#_M1008_g X 0.00294768f $X=1.61 $Y=0.665 $X2=0 $Y2=0
cc_133 N_A_186_239#_c_91_n X 0.0204439f $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A_186_239#_c_92_n X 0.0175785f $X=1.57 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A_186_239#_c_102_n X 0.0138212f $X=1.735 $Y=1.71 $X2=0 $Y2=0
cc_136 N_A_186_239#_M1008_g N_VGND_c_326_n 0.00679012f $X=1.61 $Y=0.665 $X2=0
+ $Y2=0
cc_137 N_A_186_239#_c_89_n N_VGND_c_327_n 0.0040165f $X=1.18 $Y=1.195 $X2=0
+ $Y2=0
cc_138 N_A_186_239#_M1008_g N_VGND_c_327_n 0.0040165f $X=1.61 $Y=0.665 $X2=0
+ $Y2=0
cc_139 N_A_186_239#_c_97_n N_VGND_c_328_n 0.00541298f $X=3.032 $Y=0.877 $X2=0
+ $Y2=0
cc_140 N_A_186_239#_c_89_n N_VGND_c_329_n 0.00686329f $X=1.18 $Y=1.195 $X2=0
+ $Y2=0
cc_141 N_A_186_239#_M1008_g N_VGND_c_329_n 0.00686329f $X=1.61 $Y=0.665 $X2=0
+ $Y2=0
cc_142 N_A_186_239#_c_97_n N_VGND_c_329_n 0.00979855f $X=3.032 $Y=0.877 $X2=0
+ $Y2=0
cc_143 N_A_186_239#_c_89_n N_VGND_c_330_n 0.00679012f $X=1.18 $Y=1.195 $X2=0
+ $Y2=0
cc_144 N_B_M1003_g N_A_28_367#_M1007_g 0.0205012f $X=2.13 $Y=2.045 $X2=0 $Y2=0
cc_145 B N_A_28_367#_M1007_g 0.00633695f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_146 B N_A_28_367#_c_213_n 0.0105618f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B_c_174_n N_A_28_367#_c_213_n 0.0310111f $X=2.11 $Y=1.36 $X2=0 $Y2=0
cc_148 B N_A_28_367#_c_215_n 0.0187318f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_149 N_B_c_174_n N_A_28_367#_c_215_n 0.00319182f $X=2.11 $Y=1.36 $X2=0 $Y2=0
cc_150 N_B_c_175_n N_A_28_367#_c_215_n 0.011638f $X=2.11 $Y=1.195 $X2=0 $Y2=0
cc_151 N_B_c_175_n N_A_28_367#_c_217_n 0.0310111f $X=2.11 $Y=1.195 $X2=0 $Y2=0
cc_152 N_B_M1003_g N_VPWR_c_271_n 0.00905665f $X=2.13 $Y=2.045 $X2=0 $Y2=0
cc_153 N_B_M1003_g N_VPWR_c_273_n 5.19665e-19 $X=2.13 $Y=2.045 $X2=0 $Y2=0
cc_154 N_B_c_175_n N_X_c_302_n 0.00111702f $X=2.11 $Y=1.195 $X2=0 $Y2=0
cc_155 B X 0.00427822f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B_c_175_n N_VGND_c_328_n 0.00275208f $X=2.11 $Y=1.195 $X2=0 $Y2=0
cc_157 N_B_c_175_n N_VGND_c_329_n 0.00412665f $X=2.11 $Y=1.195 $X2=0 $Y2=0
cc_158 N_A_28_367#_M1007_g N_VPWR_c_271_n 5.16628e-19 $X=2.56 $Y=2.045 $X2=0
+ $Y2=0
cc_159 N_A_28_367#_M1007_g N_VPWR_c_273_n 0.00908229f $X=2.56 $Y=2.045 $X2=0
+ $Y2=0
cc_160 N_A_28_367#_c_215_n N_X_M1002_s 0.00421127f $X=2.26 $Y=0.62 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_28_367#_c_215_n N_X_c_302_n 0.0245674f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_162 N_A_28_367#_c_215_n N_VGND_M1004_d 0.00951914f $X=2.26 $Y=0.62 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_28_367#_c_215_n N_VGND_M1008_d 0.0134236f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_164 N_A_28_367#_c_215_n N_VGND_c_326_n 0.0329712f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_165 N_A_28_367#_c_217_n N_VGND_c_326_n 0.00118565f $X=2.65 $Y=0.39 $X2=0
+ $Y2=0
cc_166 N_A_28_367#_c_215_n N_VGND_c_327_n 0.0128109f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_167 N_A_28_367#_c_215_n N_VGND_c_328_n 0.0408356f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_168 N_A_28_367#_c_217_n N_VGND_c_328_n 0.00600801f $X=2.65 $Y=0.39 $X2=0
+ $Y2=0
cc_169 N_A_28_367#_c_215_n N_VGND_c_329_n 0.054925f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_170 N_A_28_367#_c_216_n N_VGND_c_329_n 0.0138393f $X=0.305 $Y=0.62 $X2=0
+ $Y2=0
cc_171 N_A_28_367#_c_217_n N_VGND_c_329_n 0.00824115f $X=2.65 $Y=0.39 $X2=0
+ $Y2=0
cc_172 N_A_28_367#_c_215_n N_VGND_c_330_n 0.0284102f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_173 N_A_28_367#_c_216_n N_VGND_c_330_n 0.0106657f $X=0.305 $Y=0.62 $X2=0
+ $Y2=0
cc_174 N_A_28_367#_c_215_n A_455_133# 0.00178136f $X=2.26 $Y=0.62 $X2=-0.19
+ $Y2=-0.245
cc_175 N_VPWR_c_269_n N_X_M1000_s 0.0041489f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_176 N_VPWR_c_275_n X 0.0136943f $X=1.485 $Y=3.33 $X2=0 $Y2=0
cc_177 N_VPWR_c_269_n X 0.00866972f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_178 N_X_M1002_s N_VGND_c_329_n 0.00287061f $X=1.255 $Y=0.245 $X2=0 $Y2=0
