* File: sky130_fd_sc_lp__nand3_1.pex.spice
* Created: Fri Aug 28 10:48:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3_1%C 3 6 8 10 17 19
r28 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.495
+ $X2=0.54 $Y2=1.66
r29 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.495
+ $X2=0.54 $Y2=1.33
r30 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.495 $X2=0.54 $Y2=1.495
r31 10 18 3.98693 $w=5.38e-07 $l=1.8e-07 $layer=LI1_cond $X=0.72 $Y=1.48
+ $X2=0.54 $Y2=1.48
r32 8 18 6.64488 $w=5.38e-07 $l=3e-07 $layer=LI1_cond $X=0.24 $Y=1.48 $X2=0.54
+ $Y2=1.48
r33 6 20 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.63 $Y=2.465
+ $X2=0.63 $Y2=1.66
r34 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.63 $Y=0.8 $X2=0.63
+ $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_1%B 3 6 8 9 10 11 17 19
r36 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.495
+ $X2=1.11 $Y2=1.66
r37 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.495
+ $X2=1.11 $Y2=1.33
r38 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.495 $X2=1.11 $Y2=1.495
r39 11 18 6.21953 $w=3.13e-07 $l=1.7e-07 $layer=LI1_cond $X=1.182 $Y=1.665
+ $X2=1.182 $Y2=1.495
r40 10 18 7.3171 $w=3.13e-07 $l=2e-07 $layer=LI1_cond $X=1.182 $Y=1.295
+ $X2=1.182 $Y2=1.495
r41 9 10 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.182 $Y=0.925
+ $X2=1.182 $Y2=1.295
r42 8 9 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.182 $Y=0.555
+ $X2=1.182 $Y2=0.925
r43 6 20 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=1.06 $Y=2.465
+ $X2=1.06 $Y2=1.66
r44 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.02 $Y=0.8 $X2=1.02
+ $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_1%A 3 6 8 9 10 11 17 19
r31 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.495
+ $X2=1.68 $Y2=1.66
r32 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.495
+ $X2=1.68 $Y2=1.33
r33 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.495 $X2=1.68 $Y2=1.495
r34 11 18 7.68295 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=1.637 $Y=1.665
+ $X2=1.637 $Y2=1.495
r35 10 18 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=1.637 $Y=1.295
+ $X2=1.637 $Y2=1.495
r36 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.637 $Y=0.925
+ $X2=1.637 $Y2=1.295
r37 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.637 $Y=0.555
+ $X2=1.637 $Y2=0.925
r38 6 20 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=1.59 $Y=2.465
+ $X2=1.59 $Y2=1.66
r39 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.59 $Y=0.8 $X2=1.59
+ $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_1%VPWR 1 2 7 9 13 17 19 23 24 30
r29 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 21 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.33 $Y2=3.33
r32 21 23 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 19 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 19 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 19 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 15 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=3.245
+ $X2=1.33 $Y2=3.33
r37 15 17 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=1.33 $Y=3.245
+ $X2=1.33 $Y2=2.4
r38 14 27 3.90694 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r39 13 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=1.33 $Y2=3.33
r40 13 14 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=0.465 $Y2=3.33
r41 9 12 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=0.34 $Y=2.085
+ $X2=0.34 $Y2=2.95
r42 7 27 3.23622 $w=2.5e-07 $l=1.44375e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.232 $Y2=3.33
r43 7 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.34 $Y2=2.95
r44 2 17 300 $w=1.7e-07 $l=6.55286e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.835 $X2=1.33 $Y2=2.4
r45 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=1.835 $X2=0.38 $Y2=2.95
r46 1 9 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=1.835 $X2=0.38 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_1%Y 1 2 3 12 14 15 16 26 33 38
r34 16 26 4.88885 $w=2e-07 $l=3.25e-07 $layer=LI1_cond $X=1.99 $Y=2.02 $X2=1.665
+ $Y2=2.02
r35 16 38 11.5426 $w=9.18e-07 $l=7.9e-07 $layer=LI1_cond $X=1.99 $Y=2.12
+ $X2=1.99 $Y2=2.91
r36 16 26 1.94091 $w=1.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.63 $Y=2.02
+ $X2=1.665 $Y2=2.02
r37 15 16 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=1.63
+ $Y2=2.02
r38 15 27 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=1.2 $Y=2.02
+ $X2=0.995 $Y2=2.02
r39 14 27 4.86411 $w=2e-07 $l=1.8e-07 $layer=LI1_cond $X=0.815 $Y=2.02 $X2=0.995
+ $Y2=2.02
r40 14 33 19.066 $w=5.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.815 $Y=2.12
+ $X2=0.815 $Y2=2.91
r41 10 16 2.22342 $w=5.15e-07 $l=1.78115e-07 $layer=LI1_cond $X=2.125 $Y=1.92
+ $X2=1.99 $Y2=2.02
r42 10 12 42.3068 $w=3.78e-07 $l=1.395e-06 $layer=LI1_cond $X=2.125 $Y=1.92
+ $X2=2.125 $Y2=0.525
r43 3 16 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.835 $X2=1.805 $Y2=2.005
r44 3 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.835 $X2=1.805 $Y2=2.91
r45 2 14 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.835 $X2=0.845 $Y2=2.005
r46 2 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.835 $X2=0.845 $Y2=2.91
r47 1 12 91 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_NDIFF $count=2 $X=1.665
+ $Y=0.38 $X2=2.02 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_1%VGND 1 4 6 8 15 16
r22 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r23 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r24 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r25 12 15 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r26 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r27 10 19 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.29
+ $Y2=0
r28 10 12 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.72
+ $Y2=0
r29 8 16 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r30 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r31 4 19 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.29 $Y2=0
r32 4 6 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.415 $Y2=0.525
r33 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.29
+ $Y=0.38 $X2=0.415 $Y2=0.525
.ends

