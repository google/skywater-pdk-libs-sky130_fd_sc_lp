* File: sky130_fd_sc_lp__nor3_m.pex.spice
* Created: Fri Aug 28 10:56:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3_M%A 2 5 6 8 10 11 13 16 18 19 20 21 27
c37 27 0 4.44504e-20 $X=0.27 $Y=1.02
c38 18 0 1.77859e-19 $X=0.24 $Y=0.925
r39 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.02 $X2=0.27 $Y2=1.02
r40 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r41 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r42 19 28 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.02
r43 18 28 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.02
r44 14 16 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.36 $Y=2.23
+ $X2=0.54 $Y2=2.23
r45 12 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.36
+ $X2=0.27 $Y2=1.02
r46 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.36
+ $X2=0.27 $Y2=1.525
r47 11 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.005
+ $X2=0.27 $Y2=1.02
r48 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.34 $Y=0.855
+ $X2=0.34 $Y2=1.005
r49 6 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.54 $Y=2.305
+ $X2=0.54 $Y2=2.23
r50 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=2.305 $X2=0.54
+ $Y2=2.625
r51 5 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.5 $Y=0.535 $X2=0.5
+ $Y2=0.855
r52 2 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.155
+ $X2=0.36 $Y2=2.23
r53 2 13 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.155
+ $X2=0.36 $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_M%B 3 7 11 12 13 14 15 16 17 24
c44 13 0 6.97414e-20 $X=0.72 $Y=1.295
c45 7 0 1.77859e-19 $X=0.93 $Y=2.625
r46 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.41 $X2=0.84 $Y2=1.41
r47 16 17 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.78 $Y=2.405
+ $X2=0.78 $Y2=2.775
r48 15 16 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.78 $Y=2.035
+ $X2=0.78 $Y2=2.405
r49 14 15 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.78 $Y=1.665
+ $X2=0.78 $Y2=2.035
r50 14 25 10.1336 $w=2.88e-07 $l=2.55e-07 $layer=LI1_cond $X=0.78 $Y=1.665
+ $X2=0.78 $Y2=1.41
r51 13 25 4.57003 $w=2.88e-07 $l=1.15e-07 $layer=LI1_cond $X=0.78 $Y=1.295
+ $X2=0.78 $Y2=1.41
r52 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.84 $Y=1.75
+ $X2=0.84 $Y2=1.41
r53 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.75
+ $X2=0.84 $Y2=1.915
r54 10 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.245
+ $X2=0.84 $Y2=1.41
r55 7 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.93 $Y=2.625
+ $X2=0.93 $Y2=1.915
r56 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.93 $Y=0.535
+ $X2=0.93 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_M%C 3 7 11 12 13 14 15 20
r34 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=1.375 $X2=1.38 $Y2=1.375
r35 14 15 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.29 $Y=1.665
+ $X2=1.29 $Y2=2.035
r36 14 21 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.29 $Y=1.665
+ $X2=1.29 $Y2=1.375
r37 13 21 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=1.29 $Y=1.295 $X2=1.29
+ $Y2=1.375
r38 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.38 $Y=1.715
+ $X2=1.38 $Y2=1.375
r39 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.715
+ $X2=1.38 $Y2=1.88
r40 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.21
+ $X2=1.38 $Y2=1.375
r41 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.36 $Y=0.535
+ $X2=1.36 $Y2=1.21
r42 3 12 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.32 $Y=2.625
+ $X2=1.32 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_M%VPWR 1 4 6 8 15 16
r19 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r20 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r21 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r22 12 15 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r23 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r24 10 19 3.64151 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r25 10 12 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 8 16 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 4 19 3.27368 $w=2.1e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.197 $Y2=3.33
r29 4 6 32.4805 $w=2.08e-07 $l=6.15e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.63
r30 1 6 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.415 $X2=0.29 $Y2=2.63
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_M%Y 1 2 3 10 14 17 21 23 24 29
c38 24 0 4.44504e-20 $X=0.72 $Y=0.925
r39 24 29 9.56757 $w=3.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.715 $Y=0.84
+ $X2=0.715 $Y2=0.6
r40 19 21 5.18301 $w=4.48e-07 $l=1.95e-07 $layer=LI1_cond $X=1.535 $Y=2.62
+ $X2=1.73 $Y2=2.62
r41 17 21 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.73 $Y=2.395
+ $X2=1.73 $Y2=2.62
r42 16 23 3.6114 $w=2.57e-07 $l=1.23386e-07 $layer=LI1_cond $X=1.73 $Y=1.01
+ $X2=1.642 $Y2=0.925
r43 16 17 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=1.73 $Y=1.01
+ $X2=1.73 $Y2=2.395
r44 12 23 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=1.642 $Y=0.84
+ $X2=1.642 $Y2=0.925
r45 12 14 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=1.642 $Y=0.84
+ $X2=1.642 $Y2=0.6
r46 11 24 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.82 $Y=0.925
+ $X2=0.715 $Y2=0.925
r47 10 23 2.87242 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.47 $Y=0.925
+ $X2=1.642 $Y2=0.925
r48 10 11 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.47 $Y=0.925
+ $X2=0.82 $Y2=0.925
r49 3 19 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=2.415 $X2=1.535 $Y2=2.62
r50 2 14 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.325 $X2=1.575 $Y2=0.6
r51 1 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.325 $X2=0.715 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_M%VGND 1 2 7 9 13 16 17 18 25 26
r26 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r27 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r28 23 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r29 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 20 29 3.64449 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r31 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.72
+ $Y2=0
r32 18 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r33 18 23 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r34 16 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.72
+ $Y2=0
r35 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=1.145
+ $Y2=0
r36 15 25 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.68
+ $Y2=0
r37 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.145
+ $Y2=0
r38 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0
r39 11 13 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0.47
r40 7 29 3.2707 $w=2.1e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.195 $Y2=0
r41 7 9 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.285 $Y2=0.47
r42 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.325 $X2=1.145 $Y2=0.47
r43 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.325 $X2=0.285 $Y2=0.47
.ends

