# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a22oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.880000 1.210000 6.580000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.750000 1.425000 8.005000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.775000 1.355000 4.645000 1.525000 ;
        RECT 2.985000 1.210000 4.645000 1.355000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 1.210000 2.245000 1.525000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.705000 3.825000 1.875000 ;
        RECT 0.835000 1.875000 1.165000 2.735000 ;
        RECT 1.695000 1.875000 2.025000 2.735000 ;
        RECT 2.425000 0.595000 2.815000 0.815000 ;
        RECT 2.425000 0.815000 5.845000 1.040000 ;
        RECT 2.425000 1.040000 2.815000 1.145000 ;
        RECT 2.425000 1.145000 2.595000 1.705000 ;
        RECT 2.555000 1.875000 2.885000 2.735000 ;
        RECT 3.495000 1.875000 3.825000 2.735000 ;
        RECT 5.645000 0.695000 5.845000 0.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.160000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 8.350000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.275000  0.315000 0.535000 0.870000 ;
      RECT 0.275000  0.870000 2.245000 1.040000 ;
      RECT 0.405000  1.825000 0.665000 2.905000 ;
      RECT 0.405000  2.905000 4.290000 3.075000 ;
      RECT 0.705000  0.085000 1.035000 0.700000 ;
      RECT 1.205000  0.315000 1.395000 0.870000 ;
      RECT 1.335000  2.045000 1.525000 2.905000 ;
      RECT 1.565000  0.085000 1.895000 0.700000 ;
      RECT 2.065000  0.255000 4.045000 0.425000 ;
      RECT 2.065000  0.425000 2.245000 0.870000 ;
      RECT 2.195000  2.045000 2.385000 2.905000 ;
      RECT 2.995000  0.425000 4.045000 0.635000 ;
      RECT 3.055000  2.045000 3.325000 2.905000 ;
      RECT 3.995000  1.755000 6.045000 1.925000 ;
      RECT 3.995000  1.925000 4.290000 2.905000 ;
      RECT 4.295000  0.275000 6.275000 0.525000 ;
      RECT 4.460000  2.095000 4.790000 3.245000 ;
      RECT 4.960000  1.925000 5.150000 3.075000 ;
      RECT 5.320000  2.095000 5.650000 3.245000 ;
      RECT 5.820000  1.925000 6.045000 1.930000 ;
      RECT 5.820000  1.930000 7.845000 2.100000 ;
      RECT 5.820000  2.100000 6.055000 3.075000 ;
      RECT 6.015000  0.525000 6.275000 0.775000 ;
      RECT 6.015000  0.775000 7.135000 1.040000 ;
      RECT 6.225000  2.270000 6.555000 3.245000 ;
      RECT 6.445000  0.085000 6.775000 0.605000 ;
      RECT 6.725000  2.100000 6.915000 3.075000 ;
      RECT 6.855000  1.040000 7.135000 1.065000 ;
      RECT 6.855000  1.065000 8.065000 1.255000 ;
      RECT 6.945000  0.255000 7.135000 0.775000 ;
      RECT 7.085000  2.270000 7.415000 3.245000 ;
      RECT 7.305000  0.085000 7.635000 0.895000 ;
      RECT 7.585000  2.100000 7.845000 3.075000 ;
      RECT 7.805000  0.255000 8.065000 1.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__a22oi_4
END LIBRARY
