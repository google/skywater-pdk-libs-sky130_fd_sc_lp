* File: sky130_fd_sc_lp__nor4_1.pex.spice
* Created: Wed Sep  2 10:10:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4_1%A 3 7 9 12 13
c23 13 0 5.81704e-20 $X=0.38 $Y=1.51
r24 12 15 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.38 $Y=1.51
+ $X2=0.38 $Y2=1.675
r25 12 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.38 $Y=1.51
+ $X2=0.38 $Y2=1.345
r26 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.38
+ $Y=1.51 $X2=0.38 $Y2=1.51
r27 9 13 4.70075 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.275 $Y=1.665
+ $X2=0.275 $Y2=1.51
r28 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.675
r29 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_1%B 3 7 9 10 11 12 19 23 35
c43 7 0 1.82149e-19 $X=0.955 $Y=2.465
r44 23 35 2.00169 $w=4.17e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.757 $Y=2.082
+ $X2=0.842 $Y2=2.035
r45 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.675
r46 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.345
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.51 $X2=0.925 $Y2=1.51
r48 11 12 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.757 $Y=2.405
+ $X2=0.757 $Y2=2.775
r49 10 35 0.555875 $w=4.17e-07 $l=1.9e-08 $layer=LI1_cond $X=0.842 $Y=2.016
+ $X2=0.842 $Y2=2.035
r50 10 11 10.7798 $w=3.23e-07 $l=3.04e-07 $layer=LI1_cond $X=0.757 $Y=2.101
+ $X2=0.757 $Y2=2.405
r51 10 23 0.673736 $w=3.23e-07 $l=1.9e-08 $layer=LI1_cond $X=0.757 $Y=2.101
+ $X2=0.757 $Y2=2.082
r52 9 10 10.2691 $w=4.17e-07 $l=3.51e-07 $layer=LI1_cond $X=0.842 $Y=1.665
+ $X2=0.842 $Y2=2.016
r53 9 20 4.53477 $w=4.17e-07 $l=1.55e-07 $layer=LI1_cond $X=0.842 $Y=1.665
+ $X2=0.842 $Y2=1.51
r54 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.955 $Y=2.465
+ $X2=0.955 $Y2=1.675
r55 3 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.905 $Y=0.655
+ $X2=0.905 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_1%C 3 7 9 10 11 12 19 20 36
c44 20 0 1.23978e-19 $X=1.465 $Y=1.51
c45 7 0 4.25493e-20 $X=1.555 $Y=0.655
r46 36 37 1.83035 $w=4.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.535 $Y=1.665
+ $X2=1.535 $Y2=1.71
r47 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.51
+ $X2=1.465 $Y2=1.675
r48 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.51
+ $X2=1.465 $Y2=1.345
r49 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.51 $X2=1.465 $Y2=1.51
r50 11 12 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.59 $Y=2.405
+ $X2=1.59 $Y2=2.775
r51 10 11 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.59 $Y=2.035
+ $X2=1.59 $Y2=2.405
r52 9 36 0.50897 $w=4.68e-07 $l=2e-08 $layer=LI1_cond $X=1.535 $Y=1.645
+ $X2=1.535 $Y2=1.665
r53 9 20 3.43554 $w=4.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=1.645
+ $X2=1.535 $Y2=1.51
r54 9 10 9.76375 $w=3.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.59 $Y=1.73
+ $X2=1.59 $Y2=2.035
r55 9 37 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=1.59 $Y=1.73 $X2=1.59
+ $Y2=1.71
r56 7 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.555 $Y=0.655
+ $X2=1.555 $Y2=1.345
r57 3 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.445 $Y=2.465
+ $X2=1.445 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_1%D 3 7 10 11 12 16
c32 11 0 4.25493e-20 $X=2.64 $Y=1.295
r33 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=1.375 $X2=2.365 $Y2=1.375
r34 12 17 7.5103 $w=4.43e-07 $l=2.9e-07 $layer=LI1_cond $X=2.502 $Y=1.665
+ $X2=2.502 $Y2=1.375
r35 11 17 2.07181 $w=4.43e-07 $l=8e-08 $layer=LI1_cond $X=2.502 $Y=1.295
+ $X2=2.502 $Y2=1.375
r36 9 16 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.06 $Y=1.375
+ $X2=2.365 $Y2=1.375
r37 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=1.375
+ $X2=1.985 $Y2=1.375
r38 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.54
+ $X2=1.985 $Y2=1.375
r39 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.985 $Y=1.54
+ $X2=1.985 $Y2=2.465
r40 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.21
+ $X2=1.985 $Y2=1.375
r41 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.985 $Y=1.21
+ $X2=1.985 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_1%VPWR 1 4 6 10 17 18
r27 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r29 15 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 14 17 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 12 21 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r33 12 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 10 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 10 15 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 6 9 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.26 $Y=2.005
+ $X2=0.26 $Y2=2.95
r37 4 21 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r38 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r39 1 9 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r40 1 6 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_1%Y 1 2 3 12 14 15 18 23 25 26 27 41
r55 27 37 4.74535 $w=4.23e-07 $l=1.75e-07 $layer=LI1_cond $X=2.152 $Y=2.775
+ $X2=2.152 $Y2=2.95
r56 26 27 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.152 $Y=2.405
+ $X2=2.152 $Y2=2.775
r57 26 31 7.13159 $w=4.23e-07 $l=2.63e-07 $layer=LI1_cond $X=2.152 $Y=2.405
+ $X2=2.152 $Y2=2.142
r58 25 31 3.44377 $w=4.23e-07 $l=1.27e-07 $layer=LI1_cond $X=2.152 $Y=2.015
+ $X2=2.152 $Y2=2.142
r59 25 41 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=2.152 $Y=2.015
+ $X2=2.152 $Y2=1.93
r60 20 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.235
+ $X2=2.025 $Y2=1.15
r61 20 41 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.025 $Y=1.235
+ $X2=2.025 $Y2=1.93
r62 16 23 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.735 $Y=1.15
+ $X2=2.025 $Y2=1.15
r63 16 18 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=1.735 $Y=1.065
+ $X2=1.735 $Y2=0.42
r64 14 16 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.605 $Y=1.15
+ $X2=1.735 $Y2=1.15
r65 14 15 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.605 $Y=1.15
+ $X2=0.855 $Y2=1.15
r66 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.725 $Y=1.065
+ $X2=0.855 $Y2=1.15
r67 10 12 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=0.725 $Y=1.065
+ $X2=0.725 $Y2=0.42
r68 3 25 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=2.06 $Y=1.835
+ $X2=2.2 $Y2=2.015
r69 3 37 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=1.835 $X2=2.2 $Y2=2.95
r70 2 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.63
+ $Y=0.235 $X2=1.77 $Y2=0.42
r71 1 12 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_1%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r41 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 37 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r45 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.2
+ $Y2=0
r47 34 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.64
+ $Y2=0
r48 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r49 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.23
+ $Y2=0
r51 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.68
+ $Y2=0
r52 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.2
+ $Y2=0
r53 29 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.68
+ $Y2=0
r54 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r55 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r56 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 25 40 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r58 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r59 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.23
+ $Y2=0
r60 24 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r61 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r62 22 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r63 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r64 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.2 $Y=0.085
+ $X2=2.2 $Y2=0.38
r65 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r66 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.38
r67 10 40 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r68 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r69 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.235 $X2=2.2 $Y2=0.38
r70 2 16 91 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.23 $Y2=0.38
r71 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

