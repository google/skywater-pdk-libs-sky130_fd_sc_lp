* File: sky130_fd_sc_lp__o221ai_0.spice
* Created: Fri Aug 28 11:08:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o221ai_0  VNB VPB C1 B1 B2 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_A_110_47#_M1002_d N_C1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_196_47#_M1006_d N_B1_M1006_g N_A_110_47#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_196_47#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1953 AS=0.0588 PD=1.3 PS=0.7 NRD=24.276 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_196_47#_M1004_d N_A1_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1953 PD=0.7 PS=1.3 NRD=0 NRS=24.276 M=1 R=2.8 SA=75002
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_110_47#_M1007_d N_B2_M1007_g N_A_196_47#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_C1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1003 A_214_468# N_B1_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g A_214_468# VPB PHIGHVT L=0.15 W=0.64 AD=0.1248
+ AS=0.0672 PD=1.03 PS=0.85 NRD=18.4589 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 A_394_468# N_A2_M1008_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1248 PD=0.85 PS=1.03 NRD=15.3857 NRS=15.3857 M=1 R=4.26667 SA=75001.5
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_394_468# VPB PHIGHVT L=0.15 W=0.64 AD=0.208
+ AS=0.0672 PD=1.93 PS=0.85 NRD=18.4589 NRS=15.3857 M=1 R=4.26667 SA=75001.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o221ai_0.pxi.spice"
*
.ends
*
*
