* File: sky130_fd_sc_lp__a2111o_4.spice
* Created: Fri Aug 28 09:46:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111o_4.pex.spice"
.subckt sky130_fd_sc_lp__a2111o_4  VNB VPB D1 C1 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_D1_M1004_g N_A_77_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1004_d N_D1_M1022_g N_A_77_47#_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_C1_M1002_g N_A_77_47#_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1002_d N_C1_M1012_g N_A_77_47#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1005 N_A_77_47#_M1012_s N_B1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3717 PD=1.12 PS=1.725 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75002.1
+ A=0.126 P=1.98 MULT=1
MM1014 N_A_77_47#_M1014_d N_B1_M1014_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3717 PD=1.12 PS=1.725 NRD=0 NRS=0 M=1 R=5.6 SA=75003 SB=75001.1
+ A=0.126 P=1.98 MULT=1
MM1003 N_A_77_47#_M1014_d N_A1_M1003_g N_A_813_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1016 N_A_77_47#_M1016_d N_A1_M1016_g N_A_813_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_A_813_47#_M1010_d N_A2_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1021 N_A_813_47#_M1010_d N_A2_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1021_s N_A_77_47#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A_77_47#_M1008_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1008_d N_A_77_47#_M1019_g N_X_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1027 N_VGND_M1027_d N_A_77_47#_M1027_g N_X_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_63_367#_M1006_d N_D1_M1006_g N_A_77_47#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1018 N_A_63_367#_M1018_d N_D1_M1018_g N_A_77_47#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1000 N_A_63_367#_M1018_d N_C1_M1000_g N_A_318_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_A_63_367#_M1013_d N_C1_M1013_g N_A_318_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_A_318_367#_M1009_d N_B1_M1009_g N_A_511_349#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1025 N_A_318_367#_M1009_d N_B1_M1025_g N_A_511_349#_M1025_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.32445 PD=1.54 PS=1.775 NRD=0 NRS=18.7544 M=1 R=8.4
+ SA=75000.6 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1015 N_A_511_349#_M1025_s N_A1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.32445 AS=0.1764 PD=1.775 PS=1.54 NRD=17.9664 NRS=0 M=1 R=8.4
+ SA=75001.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1023 N_A_511_349#_M1023_d N_A1_M1023_g N_VPWR_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_A_511_349#_M1001_d N_A2_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1020 N_A_511_349#_M1001_d N_A2_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1011 N_X_M1011_d N_A_77_47#_M1011_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1017 N_X_M1011_d N_A_77_47#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1024 N_X_M1024_d N_A_77_47#_M1024_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1026 N_X_M1024_d N_A_77_47#_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=16.1579 P=20.99
*
.include "sky130_fd_sc_lp__a2111o_4.pxi.spice"
*
.ends
*
*
