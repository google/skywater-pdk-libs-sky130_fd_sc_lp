* File: sky130_fd_sc_lp__o2bb2a_0.pxi.spice
* Created: Wed Sep  2 10:21:13 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2A_0%A_80_176# N_A_80_176#_M1001_s N_A_80_176#_M1011_d
+ N_A_80_176#_c_96_n N_A_80_176#_M1005_g N_A_80_176#_M1002_g N_A_80_176#_c_98_n
+ N_A_80_176#_c_99_n N_A_80_176#_c_100_n N_A_80_176#_c_101_n N_A_80_176#_c_108_n
+ N_A_80_176#_c_186_p N_A_80_176#_c_109_n N_A_80_176#_c_110_n
+ N_A_80_176#_c_111_n N_A_80_176#_c_112_n N_A_80_176#_c_113_n
+ N_A_80_176#_c_114_n N_A_80_176#_c_102_n N_A_80_176#_c_103_n
+ N_A_80_176#_c_116_n N_A_80_176#_c_117_n N_A_80_176#_c_104_n
+ N_A_80_176#_c_118_n N_A_80_176#_c_105_n PM_SKY130_FD_SC_LP__O2BB2A_0%A_80_176#
x_PM_SKY130_FD_SC_LP__O2BB2A_0%A1_N N_A1_N_M1003_g N_A1_N_M1007_g A1_N A1_N
+ N_A1_N_c_229_n PM_SKY130_FD_SC_LP__O2BB2A_0%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2A_0%A2_N N_A2_N_M1004_g N_A2_N_c_267_n N_A2_N_c_272_n
+ N_A2_N_M1009_g N_A2_N_c_273_n A2_N A2_N N_A2_N_c_269_n N_A2_N_c_270_n
+ PM_SKY130_FD_SC_LP__O2BB2A_0%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2A_0%A_229_483# N_A_229_483#_M1004_d
+ N_A_229_483#_M1007_d N_A_229_483#_c_332_n N_A_229_483#_c_325_n
+ N_A_229_483#_c_326_n N_A_229_483#_c_333_n N_A_229_483#_c_334_n
+ N_A_229_483#_c_327_n N_A_229_483#_M1001_g N_A_229_483#_M1011_g
+ N_A_229_483#_c_336_n N_A_229_483#_c_328_n N_A_229_483#_c_337_n
+ N_A_229_483#_c_338_n N_A_229_483#_c_329_n N_A_229_483#_c_330_n
+ N_A_229_483#_c_331_n PM_SKY130_FD_SC_LP__O2BB2A_0%A_229_483#
x_PM_SKY130_FD_SC_LP__O2BB2A_0%B2 N_B2_M1010_g N_B2_M1008_g N_B2_c_415_n
+ N_B2_c_419_n B2 B2 N_B2_c_417_n PM_SKY130_FD_SC_LP__O2BB2A_0%B2
x_PM_SKY130_FD_SC_LP__O2BB2A_0%B1 N_B1_M1006_g N_B1_M1000_g N_B1_c_458_n
+ N_B1_c_459_n B1 B1 B1 N_B1_c_456_n PM_SKY130_FD_SC_LP__O2BB2A_0%B1
x_PM_SKY130_FD_SC_LP__O2BB2A_0%X N_X_M1002_s N_X_M1005_s N_X_c_488_n X X X X X X
+ N_X_c_487_n X PM_SKY130_FD_SC_LP__O2BB2A_0%X
x_PM_SKY130_FD_SC_LP__O2BB2A_0%VPWR N_VPWR_M1005_d N_VPWR_M1009_d N_VPWR_M1006_d
+ N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n VPWR
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n
+ N_VPWR_c_505_n PM_SKY130_FD_SC_LP__O2BB2A_0%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2A_0%VGND N_VGND_M1002_d N_VGND_M1010_d N_VGND_c_559_n
+ N_VGND_c_560_n VGND N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n
+ N_VGND_c_564_n N_VGND_c_565_n PM_SKY130_FD_SC_LP__O2BB2A_0%VGND
x_PM_SKY130_FD_SC_LP__O2BB2A_0%A_512_47# N_A_512_47#_M1001_d N_A_512_47#_M1000_d
+ N_A_512_47#_c_606_n N_A_512_47#_c_607_n N_A_512_47#_c_608_n
+ N_A_512_47#_c_609_n PM_SKY130_FD_SC_LP__O2BB2A_0%A_512_47#
cc_1 VNB N_A_80_176#_c_96_n 0.0241005f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.37
cc_2 VNB N_A_80_176#_M1005_g 0.00576953f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_3 VNB N_A_80_176#_c_98_n 0.0213087f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.55
cc_4 VNB N_A_80_176#_c_99_n 0.00174117f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.045
cc_5 VNB N_A_80_176#_c_100_n 0.0197466f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.045
cc_6 VNB N_A_80_176#_c_101_n 6.52195e-19 $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.3
cc_7 VNB N_A_80_176#_c_102_n 0.003158f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.445
cc_8 VNB N_A_80_176#_c_103_n 0.0156683f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=2.175
cc_9 VNB N_A_80_176#_c_104_n 0.00180775f $X=-0.19 $Y=-0.245 $X2=2.252 $Y2=0.675
cc_10 VNB N_A_80_176#_c_105_n 0.0208858f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.88
cc_11 VNB N_A1_N_M1003_g 0.0522451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A1_N 0.00659389f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.55
cc_13 VNB N_A2_N_M1004_g 0.0280469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_N_c_267_n 0.0171458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A2_N 8.29463e-19 $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.56
cc_16 VNB N_A2_N_c_269_n 0.0317087f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.55
cc_17 VNB N_A2_N_c_270_n 0.00940639f $X=-0.19 $Y=-0.245 $X2=2.252 $Y2=0.553
cc_18 VNB N_A_229_483#_c_325_n 0.0360514f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_19 VNB N_A_229_483#_c_326_n 0.0117309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_229_483#_c_327_n 0.0188286f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.56
cc_21 VNB N_A_229_483#_c_328_n 0.0171229f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.385
cc_22 VNB N_A_229_483#_c_329_n 0.0112804f $X=-0.19 $Y=-0.245 $X2=2.252 $Y2=0.445
cc_23 VNB N_A_229_483#_c_330_n 0.00738094f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=2.175
cc_24 VNB N_A_229_483#_c_331_n 0.03944f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=2.345
cc_25 VNB N_B2_M1010_g 0.0380349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B2_c_415_n 0.0249666f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_27 VNB B2 0.00642155f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.88
cc_28 VNB N_B2_c_417_n 0.0176224f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.045
cc_29 VNB N_B1_M1000_g 0.069589f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.06
cc_30 VNB B1 0.029059f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.88
cc_31 VNB N_B1_c_456_n 0.0139323f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.045
cc_32 VNB X 0.0474828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_487_n 0.0168605f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=2.26
cc_34 VNB N_VPWR_c_505_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.252 $Y2=0.675
cc_35 VNB N_VGND_c_559_n 0.00533988f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_36 VNB N_VGND_c_560_n 0.00522139f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.56
cc_37 VNB N_VGND_c_561_n 0.0560521f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.045
cc_38 VNB N_VGND_c_562_n 0.017975f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=2.99
cc_39 VNB N_VGND_c_563_n 0.224147f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=2.345
cc_40 VNB N_VGND_c_564_n 0.0249905f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=2.26
cc_41 VNB N_VGND_c_565_n 0.00497572f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.445
cc_42 VNB N_A_512_47#_c_606_n 9.95328e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.55
cc_43 VNB N_A_512_47#_c_607_n 0.0212533f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_44 VNB N_A_512_47#_c_608_n 0.00258687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_512_47#_c_609_n 0.0207448f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.56
cc_46 VPB N_A_80_176#_M1005_g 0.0557586f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_47 VPB N_A_80_176#_c_101_n 0.0046111f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.3
cc_48 VPB N_A_80_176#_c_108_n 0.00630799f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.385
cc_49 VPB N_A_80_176#_c_109_n 6.75941e-19 $X=-0.19 $Y=1.655 $X2=1.09 $Y2=2.905
cc_50 VPB N_A_80_176#_c_110_n 0.0184887f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.99
cc_51 VPB N_A_80_176#_c_111_n 0.00202489f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=2.99
cc_52 VPB N_A_80_176#_c_112_n 0.00244512f $X=-0.19 $Y=1.655 $X2=1.89 $Y2=2.905
cc_53 VPB N_A_80_176#_c_113_n 0.00637188f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=2.26
cc_54 VPB N_A_80_176#_c_114_n 0.00215786f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=2.26
cc_55 VPB N_A_80_176#_c_103_n 0.00858407f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=2.175
cc_56 VPB N_A_80_176#_c_116_n 0.0037321f $X=-0.19 $Y=1.655 $X2=2.575 $Y2=2.26
cc_57 VPB N_A_80_176#_c_117_n 5.5039e-19 $X=-0.19 $Y=1.655 $X2=2.7 $Y2=2.625
cc_58 VPB N_A_80_176#_c_118_n 0.00157448f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=2.26
cc_59 VPB N_A1_N_M1003_g 0.00627446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A1_N_M1007_g 0.028039f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.06
cc_61 VPB A1_N 0.0100813f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.55
cc_62 VPB N_A1_N_c_229_n 0.033141f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.56
cc_63 VPB N_A2_N_c_267_n 0.0246425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A2_N_c_272_n 0.0194287f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.06
cc_65 VPB N_A2_N_c_273_n 0.0219766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_229_483#_c_332_n 0.00726183f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_67 VPB N_A_229_483#_c_333_n 0.0371729f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.88
cc_68 VPB N_A_229_483#_c_334_n 0.00970743f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.56
cc_69 VPB N_A_229_483#_M1011_g 0.0239386f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.045
cc_70 VPB N_A_229_483#_c_336_n 0.00350761f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.3
cc_71 VPB N_A_229_483#_c_337_n 0.0025531f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=2.99
cc_72 VPB N_A_229_483#_c_338_n 0.0101685f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=2.26
cc_73 VPB N_A_229_483#_c_329_n 0.0248586f $X=-0.19 $Y=1.655 $X2=2.252 $Y2=0.445
cc_74 VPB N_B2_M1008_g 0.0417221f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.06
cc_75 VPB N_B2_c_419_n 0.0171647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB B2 0.004821f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.88
cc_77 VPB N_B1_M1006_g 0.027875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_B1_c_458_n 0.0271413f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_79 VPB N_B1_c_459_n 0.0183916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB B1 0.0304874f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.88
cc_81 VPB N_B1_c_456_n 0.00441166f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.045
cc_82 VPB N_X_c_488_n 0.0223211f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.55
cc_83 VPB X 0.037232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB X 0.00634768f $X=-0.19 $Y=1.655 $X2=2.72 $Y2=2.625
cc_85 VPB N_VPWR_c_506_n 0.00575715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_507_n 0.0158288f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.55
cc_87 VPB N_VPWR_c_508_n 0.0144238f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.045
cc_88 VPB N_VPWR_c_509_n 0.0354408f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.045
cc_89 VPB N_VPWR_c_510_n 0.0156862f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.385
cc_90 VPB N_VPWR_c_511_n 0.0325093f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=2.99
cc_91 VPB N_VPWR_c_512_n 0.0276135f $X=-0.19 $Y=1.655 $X2=2.252 $Y2=0.553
cc_92 VPB N_VPWR_c_513_n 0.00502701f $X=-0.19 $Y=1.655 $X2=2.575 $Y2=2.26
cc_93 VPB N_VPWR_c_514_n 0.00497514f $X=-0.19 $Y=1.655 $X2=2.72 $Y2=2.625
cc_94 VPB N_VPWR_c_505_n 0.0882059f $X=-0.19 $Y=1.655 $X2=2.252 $Y2=0.675
cc_95 N_A_80_176#_M1005_g N_A1_N_M1003_g 0.00613484f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_96 N_A_80_176#_c_99_n N_A1_N_M1003_g 0.00246601f $X=0.595 $Y=1.045 $X2=0
+ $Y2=0
cc_97 N_A_80_176#_c_100_n N_A1_N_M1003_g 0.0403484f $X=0.595 $Y=1.045 $X2=0
+ $Y2=0
cc_98 N_A_80_176#_c_101_n N_A1_N_M1003_g 6.86917e-19 $X=0.63 $Y=2.3 $X2=0 $Y2=0
cc_99 N_A_80_176#_c_105_n N_A1_N_M1003_g 0.0121541f $X=0.58 $Y=0.88 $X2=0 $Y2=0
cc_100 N_A_80_176#_M1005_g N_A1_N_M1007_g 0.0143639f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_101 N_A_80_176#_c_101_n N_A1_N_M1007_g 0.00332335f $X=0.63 $Y=2.3 $X2=0 $Y2=0
cc_102 N_A_80_176#_c_108_n N_A1_N_M1007_g 0.008628f $X=1.005 $Y=2.385 $X2=0
+ $Y2=0
cc_103 N_A_80_176#_c_109_n N_A1_N_M1007_g 0.0123674f $X=1.09 $Y=2.905 $X2=0
+ $Y2=0
cc_104 N_A_80_176#_c_111_n N_A1_N_M1007_g 0.00433919f $X=1.175 $Y=2.99 $X2=0
+ $Y2=0
cc_105 N_A_80_176#_M1005_g A1_N 9.73752e-19 $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_106 N_A_80_176#_c_101_n A1_N 0.0453453f $X=0.63 $Y=2.3 $X2=0 $Y2=0
cc_107 N_A_80_176#_c_108_n A1_N 0.0242891f $X=1.005 $Y=2.385 $X2=0 $Y2=0
cc_108 N_A_80_176#_M1005_g N_A1_N_c_229_n 0.0150528f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_109 N_A_80_176#_c_101_n N_A1_N_c_229_n 0.00227831f $X=0.63 $Y=2.3 $X2=0 $Y2=0
cc_110 N_A_80_176#_c_108_n N_A1_N_c_229_n 0.00338248f $X=1.005 $Y=2.385 $X2=0
+ $Y2=0
cc_111 N_A_80_176#_c_102_n N_A2_N_M1004_g 0.00256737f $X=2.27 $Y=0.445 $X2=0
+ $Y2=0
cc_112 N_A_80_176#_c_103_n N_A2_N_c_267_n 4.06443e-19 $X=2.29 $Y=2.175 $X2=0
+ $Y2=0
cc_113 N_A_80_176#_c_108_n N_A2_N_c_272_n 4.05202e-19 $X=1.005 $Y=2.385 $X2=0
+ $Y2=0
cc_114 N_A_80_176#_c_109_n N_A2_N_c_272_n 7.5767e-19 $X=1.09 $Y=2.905 $X2=0
+ $Y2=0
cc_115 N_A_80_176#_c_110_n N_A2_N_c_272_n 0.00982427f $X=1.805 $Y=2.99 $X2=0
+ $Y2=0
cc_116 N_A_80_176#_c_112_n N_A2_N_c_272_n 0.00700223f $X=1.89 $Y=2.905 $X2=0
+ $Y2=0
cc_117 N_A_80_176#_c_114_n N_A2_N_c_273_n 0.00200225f $X=1.975 $Y=2.26 $X2=0
+ $Y2=0
cc_118 N_A_80_176#_c_105_n A2_N 7.15918e-19 $X=0.58 $Y=0.88 $X2=0 $Y2=0
cc_119 N_A_80_176#_c_99_n N_A2_N_c_270_n 0.025033f $X=0.595 $Y=1.045 $X2=0 $Y2=0
cc_120 N_A_80_176#_c_100_n N_A2_N_c_270_n 0.00173875f $X=0.595 $Y=1.045 $X2=0
+ $Y2=0
cc_121 N_A_80_176#_c_103_n N_A_229_483#_c_325_n 0.0140172f $X=2.29 $Y=2.175
+ $X2=0 $Y2=0
cc_122 N_A_80_176#_c_104_n N_A_229_483#_c_325_n 0.00306861f $X=2.252 $Y=0.675
+ $X2=0 $Y2=0
cc_123 N_A_80_176#_c_113_n N_A_229_483#_c_333_n 0.00543979f $X=2.205 $Y=2.26
+ $X2=0 $Y2=0
cc_124 N_A_80_176#_c_103_n N_A_229_483#_c_333_n 0.00961963f $X=2.29 $Y=2.175
+ $X2=0 $Y2=0
cc_125 N_A_80_176#_c_116_n N_A_229_483#_c_333_n 0.00828064f $X=2.575 $Y=2.26
+ $X2=0 $Y2=0
cc_126 N_A_80_176#_c_118_n N_A_229_483#_c_333_n 0.00351786f $X=2.29 $Y=2.26
+ $X2=0 $Y2=0
cc_127 N_A_80_176#_c_113_n N_A_229_483#_c_334_n 0.00708637f $X=2.205 $Y=2.26
+ $X2=0 $Y2=0
cc_128 N_A_80_176#_c_114_n N_A_229_483#_c_334_n 9.69133e-19 $X=1.975 $Y=2.26
+ $X2=0 $Y2=0
cc_129 N_A_80_176#_c_104_n N_A_229_483#_c_327_n 0.00274617f $X=2.252 $Y=0.675
+ $X2=0 $Y2=0
cc_130 N_A_80_176#_c_112_n N_A_229_483#_M1011_g 0.00188505f $X=1.89 $Y=2.905
+ $X2=0 $Y2=0
cc_131 N_A_80_176#_c_116_n N_A_229_483#_M1011_g 0.0122497f $X=2.575 $Y=2.26
+ $X2=0 $Y2=0
cc_132 N_A_80_176#_c_117_n N_A_229_483#_M1011_g 0.00106454f $X=2.7 $Y=2.625
+ $X2=0 $Y2=0
cc_133 N_A_80_176#_c_108_n N_A_229_483#_c_336_n 0.00605043f $X=1.005 $Y=2.385
+ $X2=0 $Y2=0
cc_134 N_A_80_176#_c_112_n N_A_229_483#_c_336_n 0.00425336f $X=1.89 $Y=2.905
+ $X2=0 $Y2=0
cc_135 N_A_80_176#_c_114_n N_A_229_483#_c_336_n 0.0136805f $X=1.975 $Y=2.26
+ $X2=0 $Y2=0
cc_136 N_A_80_176#_c_103_n N_A_229_483#_c_336_n 0.00790546f $X=2.29 $Y=2.175
+ $X2=0 $Y2=0
cc_137 N_A_80_176#_c_103_n N_A_229_483#_c_328_n 0.0495179f $X=2.29 $Y=2.175
+ $X2=0 $Y2=0
cc_138 N_A_80_176#_c_108_n N_A_229_483#_c_337_n 0.00292628f $X=1.005 $Y=2.385
+ $X2=0 $Y2=0
cc_139 N_A_80_176#_c_110_n N_A_229_483#_c_337_n 0.0187021f $X=1.805 $Y=2.99
+ $X2=0 $Y2=0
cc_140 N_A_80_176#_c_112_n N_A_229_483#_c_337_n 0.0241115f $X=1.89 $Y=2.905
+ $X2=0 $Y2=0
cc_141 N_A_80_176#_c_113_n N_A_229_483#_c_338_n 0.00303815f $X=2.205 $Y=2.26
+ $X2=0 $Y2=0
cc_142 N_A_80_176#_c_114_n N_A_229_483#_c_338_n 0.0108937f $X=1.975 $Y=2.26
+ $X2=0 $Y2=0
cc_143 N_A_80_176#_c_103_n N_A_229_483#_c_338_n 0.0252104f $X=2.29 $Y=2.175
+ $X2=0 $Y2=0
cc_144 N_A_80_176#_c_114_n N_A_229_483#_c_329_n 0.00116505f $X=1.975 $Y=2.26
+ $X2=0 $Y2=0
cc_145 N_A_80_176#_c_102_n N_A_229_483#_c_330_n 0.0233014f $X=2.27 $Y=0.445
+ $X2=0 $Y2=0
cc_146 N_A_80_176#_c_103_n N_A_229_483#_c_330_n 0.00306197f $X=2.29 $Y=2.175
+ $X2=0 $Y2=0
cc_147 N_A_80_176#_c_103_n N_A_229_483#_c_331_n 0.014054f $X=2.29 $Y=2.175 $X2=0
+ $Y2=0
cc_148 N_A_80_176#_c_103_n N_B2_M1010_g 0.00536471f $X=2.29 $Y=2.175 $X2=0 $Y2=0
cc_149 N_A_80_176#_c_103_n N_B2_M1008_g 0.00649491f $X=2.29 $Y=2.175 $X2=0 $Y2=0
cc_150 N_A_80_176#_c_116_n N_B2_M1008_g 0.00549002f $X=2.575 $Y=2.26 $X2=0 $Y2=0
cc_151 N_A_80_176#_c_117_n N_B2_M1008_g 0.00839431f $X=2.7 $Y=2.625 $X2=0 $Y2=0
cc_152 N_A_80_176#_c_116_n N_B2_c_419_n 0.00126263f $X=2.575 $Y=2.26 $X2=0 $Y2=0
cc_153 N_A_80_176#_c_103_n B2 0.0544053f $X=2.29 $Y=2.175 $X2=0 $Y2=0
cc_154 N_A_80_176#_c_116_n B2 0.0165989f $X=2.575 $Y=2.26 $X2=0 $Y2=0
cc_155 N_A_80_176#_c_103_n N_B2_c_417_n 0.00193283f $X=2.29 $Y=2.175 $X2=0 $Y2=0
cc_156 N_A_80_176#_c_117_n N_B1_M1006_g 0.00147394f $X=2.7 $Y=2.625 $X2=0 $Y2=0
cc_157 N_A_80_176#_c_116_n N_B1_c_459_n 7.58773e-19 $X=2.575 $Y=2.26 $X2=0 $Y2=0
cc_158 N_A_80_176#_c_116_n B1 0.00192203f $X=2.575 $Y=2.26 $X2=0 $Y2=0
cc_159 N_A_80_176#_c_99_n X 0.0499124f $X=0.595 $Y=1.045 $X2=0 $Y2=0
cc_160 N_A_80_176#_c_100_n X 0.0360585f $X=0.595 $Y=1.045 $X2=0 $Y2=0
cc_161 N_A_80_176#_c_101_n X 0.0452834f $X=0.63 $Y=2.3 $X2=0 $Y2=0
cc_162 N_A_80_176#_c_186_p X 0.00631516f $X=0.715 $Y=2.385 $X2=0 $Y2=0
cc_163 N_A_80_176#_c_105_n X 0.00503573f $X=0.58 $Y=0.88 $X2=0 $Y2=0
cc_164 N_A_80_176#_c_100_n N_X_c_487_n 0.00399648f $X=0.595 $Y=1.045 $X2=0 $Y2=0
cc_165 N_A_80_176#_M1005_g X 6.74683e-19 $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_166 N_A_80_176#_c_186_p X 0.00356269f $X=0.715 $Y=2.385 $X2=0 $Y2=0
cc_167 N_A_80_176#_c_108_n N_VPWR_M1005_d 0.00361947f $X=1.005 $Y=2.385
+ $X2=-0.19 $Y2=-0.245
cc_168 N_A_80_176#_c_186_p N_VPWR_M1005_d 0.0011806f $X=0.715 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_80_176#_c_112_n N_VPWR_M1009_d 0.0115983f $X=1.89 $Y=2.905 $X2=0
+ $Y2=0
cc_170 N_A_80_176#_M1005_g N_VPWR_c_506_n 0.0126684f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_171 N_A_80_176#_c_108_n N_VPWR_c_506_n 0.00945038f $X=1.005 $Y=2.385 $X2=0
+ $Y2=0
cc_172 N_A_80_176#_c_186_p N_VPWR_c_506_n 0.00989174f $X=0.715 $Y=2.385 $X2=0
+ $Y2=0
cc_173 N_A_80_176#_c_109_n N_VPWR_c_506_n 0.0195802f $X=1.09 $Y=2.905 $X2=0
+ $Y2=0
cc_174 N_A_80_176#_c_111_n N_VPWR_c_506_n 0.0146986f $X=1.175 $Y=2.99 $X2=0
+ $Y2=0
cc_175 N_A_80_176#_c_110_n N_VPWR_c_507_n 0.0147863f $X=1.805 $Y=2.99 $X2=0
+ $Y2=0
cc_176 N_A_80_176#_c_112_n N_VPWR_c_507_n 0.0294149f $X=1.89 $Y=2.905 $X2=0
+ $Y2=0
cc_177 N_A_80_176#_c_113_n N_VPWR_c_507_n 0.00484086f $X=2.205 $Y=2.26 $X2=0
+ $Y2=0
cc_178 N_A_80_176#_c_118_n N_VPWR_c_507_n 0.0145425f $X=2.29 $Y=2.26 $X2=0 $Y2=0
cc_179 N_A_80_176#_c_117_n N_VPWR_c_509_n 0.0109327f $X=2.7 $Y=2.625 $X2=0 $Y2=0
cc_180 N_A_80_176#_M1005_g N_VPWR_c_510_n 0.00452967f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_181 N_A_80_176#_c_110_n N_VPWR_c_511_n 0.052712f $X=1.805 $Y=2.99 $X2=0 $Y2=0
cc_182 N_A_80_176#_c_111_n N_VPWR_c_511_n 0.0121867f $X=1.175 $Y=2.99 $X2=0
+ $Y2=0
cc_183 N_A_80_176#_c_117_n N_VPWR_c_512_n 0.00572876f $X=2.7 $Y=2.625 $X2=0
+ $Y2=0
cc_184 N_A_80_176#_M1005_g N_VPWR_c_505_n 0.0088676f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_185 N_A_80_176#_c_108_n N_VPWR_c_505_n 0.00613077f $X=1.005 $Y=2.385 $X2=0
+ $Y2=0
cc_186 N_A_80_176#_c_186_p N_VPWR_c_505_n 5.99092e-19 $X=0.715 $Y=2.385 $X2=0
+ $Y2=0
cc_187 N_A_80_176#_c_110_n N_VPWR_c_505_n 0.0302878f $X=1.805 $Y=2.99 $X2=0
+ $Y2=0
cc_188 N_A_80_176#_c_111_n N_VPWR_c_505_n 0.00660921f $X=1.175 $Y=2.99 $X2=0
+ $Y2=0
cc_189 N_A_80_176#_c_117_n N_VPWR_c_505_n 0.00928473f $X=2.7 $Y=2.625 $X2=0
+ $Y2=0
cc_190 N_A_80_176#_c_99_n N_VGND_c_559_n 0.00197252f $X=0.595 $Y=1.045 $X2=0
+ $Y2=0
cc_191 N_A_80_176#_c_100_n N_VGND_c_559_n 0.00137917f $X=0.595 $Y=1.045 $X2=0
+ $Y2=0
cc_192 N_A_80_176#_c_105_n N_VGND_c_559_n 0.0109289f $X=0.58 $Y=0.88 $X2=0 $Y2=0
cc_193 N_A_80_176#_c_102_n N_VGND_c_561_n 0.0139397f $X=2.27 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A_80_176#_M1001_s N_VGND_c_563_n 0.00259026f $X=2.145 $Y=0.235 $X2=0
+ $Y2=0
cc_195 N_A_80_176#_c_102_n N_VGND_c_563_n 0.0092904f $X=2.27 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_A_80_176#_c_105_n N_VGND_c_563_n 0.00852247f $X=0.58 $Y=0.88 $X2=0
+ $Y2=0
cc_197 N_A_80_176#_c_105_n N_VGND_c_564_n 0.00428763f $X=0.58 $Y=0.88 $X2=0
+ $Y2=0
cc_198 N_A_80_176#_c_104_n N_A_512_47#_c_606_n 0.0228836f $X=2.252 $Y=0.675
+ $X2=0 $Y2=0
cc_199 N_A_80_176#_c_103_n N_A_512_47#_c_608_n 0.0132397f $X=2.29 $Y=2.175 $X2=0
+ $Y2=0
cc_200 N_A1_N_M1003_g N_A2_N_M1004_g 0.0579678f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A1_N_M1003_g N_A2_N_c_267_n 0.0201289f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_202 A1_N N_A2_N_c_267_n 0.00482843f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A1_N_c_229_n N_A2_N_c_267_n 0.0130418f $X=0.98 $Y=1.955 $X2=0 $Y2=0
cc_204 N_A1_N_M1007_g N_A2_N_c_272_n 0.0120225f $X=1.07 $Y=2.625 $X2=0 $Y2=0
cc_205 N_A1_N_M1007_g N_A2_N_c_273_n 0.0130418f $X=1.07 $Y=2.625 $X2=0 $Y2=0
cc_206 N_A1_N_M1003_g A2_N 0.00965228f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A1_N_M1003_g N_A2_N_c_270_n 0.0195311f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_208 A1_N N_A2_N_c_270_n 0.0259696f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A1_N_M1007_g N_A_229_483#_c_336_n 0.00128518f $X=1.07 $Y=2.625 $X2=0
+ $Y2=0
cc_210 A1_N N_A_229_483#_c_336_n 0.0164968f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_211 A1_N N_A_229_483#_c_328_n 0.00132032f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A1_N_M1007_g N_A_229_483#_c_337_n 0.00117927f $X=1.07 $Y=2.625 $X2=0
+ $Y2=0
cc_213 A1_N N_A_229_483#_c_338_n 0.0199777f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A1_N_M1007_g N_VPWR_c_506_n 0.0024872f $X=1.07 $Y=2.625 $X2=0 $Y2=0
cc_215 N_A1_N_M1007_g N_VPWR_c_511_n 9.95699e-19 $X=1.07 $Y=2.625 $X2=0 $Y2=0
cc_216 N_A1_N_M1007_g N_VPWR_c_505_n 3.37918e-19 $X=1.07 $Y=2.625 $X2=0 $Y2=0
cc_217 N_A1_N_M1003_g N_VGND_c_559_n 0.00331718f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_218 N_A1_N_M1003_g N_VGND_c_561_n 0.00462244f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A1_N_M1003_g N_VGND_c_563_n 0.00573903f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A2_N_c_267_n N_A_229_483#_c_332_n 0.00603899f $X=1.46 $Y=2.155 $X2=0
+ $Y2=0
cc_221 N_A2_N_M1004_g N_A_229_483#_c_326_n 0.0049739f $X=1.435 $Y=0.56 $X2=0
+ $Y2=0
cc_222 N_A2_N_c_273_n N_A_229_483#_c_334_n 0.00325283f $X=1.645 $Y=2.23 $X2=0
+ $Y2=0
cc_223 N_A2_N_c_273_n N_A_229_483#_M1011_g 0.00521603f $X=1.645 $Y=2.23 $X2=0
+ $Y2=0
cc_224 N_A2_N_c_267_n N_A_229_483#_c_336_n 0.00544286f $X=1.46 $Y=2.155 $X2=0
+ $Y2=0
cc_225 N_A2_N_c_272_n N_A_229_483#_c_336_n 0.00243681f $X=1.645 $Y=2.305 $X2=0
+ $Y2=0
cc_226 N_A2_N_c_273_n N_A_229_483#_c_336_n 0.00944911f $X=1.645 $Y=2.23 $X2=0
+ $Y2=0
cc_227 N_A2_N_M1004_g N_A_229_483#_c_328_n 0.00237619f $X=1.435 $Y=0.56 $X2=0
+ $Y2=0
cc_228 N_A2_N_c_267_n N_A_229_483#_c_328_n 0.00379665f $X=1.46 $Y=2.155 $X2=0
+ $Y2=0
cc_229 A2_N N_A_229_483#_c_328_n 0.00442864f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_230 N_A2_N_c_269_n N_A_229_483#_c_328_n 0.00234298f $X=1.525 $Y=1.18 $X2=0
+ $Y2=0
cc_231 N_A2_N_c_270_n N_A_229_483#_c_328_n 0.0342211f $X=1.227 $Y=1.12 $X2=0
+ $Y2=0
cc_232 N_A2_N_c_272_n N_A_229_483#_c_337_n 0.00556363f $X=1.645 $Y=2.305 $X2=0
+ $Y2=0
cc_233 N_A2_N_c_273_n N_A_229_483#_c_337_n 0.00455272f $X=1.645 $Y=2.23 $X2=0
+ $Y2=0
cc_234 N_A2_N_c_267_n N_A_229_483#_c_338_n 0.00607839f $X=1.46 $Y=2.155 $X2=0
+ $Y2=0
cc_235 N_A2_N_c_273_n N_A_229_483#_c_338_n 0.00327969f $X=1.645 $Y=2.23 $X2=0
+ $Y2=0
cc_236 N_A2_N_c_269_n N_A_229_483#_c_338_n 0.00298284f $X=1.525 $Y=1.18 $X2=0
+ $Y2=0
cc_237 N_A2_N_c_270_n N_A_229_483#_c_338_n 0.00697105f $X=1.227 $Y=1.12 $X2=0
+ $Y2=0
cc_238 N_A2_N_c_267_n N_A_229_483#_c_329_n 0.0175891f $X=1.46 $Y=2.155 $X2=0
+ $Y2=0
cc_239 N_A2_N_c_269_n N_A_229_483#_c_330_n 0.00329767f $X=1.525 $Y=1.18 $X2=0
+ $Y2=0
cc_240 N_A2_N_c_270_n N_A_229_483#_c_330_n 0.00341302f $X=1.227 $Y=1.12 $X2=0
+ $Y2=0
cc_241 N_A2_N_c_267_n N_A_229_483#_c_331_n 0.00473966f $X=1.46 $Y=2.155 $X2=0
+ $Y2=0
cc_242 N_A2_N_c_269_n N_A_229_483#_c_331_n 0.0129557f $X=1.525 $Y=1.18 $X2=0
+ $Y2=0
cc_243 N_A2_N_c_270_n X 5.35562e-19 $X=1.227 $Y=1.12 $X2=0 $Y2=0
cc_244 N_A2_N_c_272_n N_VPWR_c_507_n 7.34082e-19 $X=1.645 $Y=2.305 $X2=0 $Y2=0
cc_245 N_A2_N_c_272_n N_VPWR_c_511_n 7.17276e-19 $X=1.645 $Y=2.305 $X2=0 $Y2=0
cc_246 N_A2_N_M1004_g N_VGND_c_561_n 0.00478016f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_247 A2_N N_VGND_c_561_n 0.00712146f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_248 N_A2_N_M1004_g N_VGND_c_563_n 0.00969038f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_249 A2_N N_VGND_c_563_n 0.00865835f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_250 N_A2_N_c_270_n N_VGND_c_563_n 0.00316723f $X=1.227 $Y=1.12 $X2=0 $Y2=0
cc_251 A2_N A_224_70# 0.00168395f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_252 N_A_229_483#_c_327_n N_B2_M1010_g 0.0189723f $X=2.485 $Y=0.765 $X2=0
+ $Y2=0
cc_253 N_A_229_483#_c_333_n N_B2_M1008_g 0.0229999f $X=2.41 $Y=2.14 $X2=0 $Y2=0
cc_254 N_A_229_483#_c_329_n N_B2_c_415_n 0.00488278f $X=1.94 $Y=1.75 $X2=0 $Y2=0
cc_255 N_A_229_483#_c_333_n B2 3.84588e-19 $X=2.41 $Y=2.14 $X2=0 $Y2=0
cc_256 N_A_229_483#_c_331_n N_B2_c_417_n 0.00488278f $X=1.942 $Y=1.585 $X2=0
+ $Y2=0
cc_257 N_A_229_483#_c_333_n N_VPWR_c_507_n 0.00140613f $X=2.41 $Y=2.14 $X2=0
+ $Y2=0
cc_258 N_A_229_483#_M1011_g N_VPWR_c_507_n 0.00420885f $X=2.485 $Y=2.625 $X2=0
+ $Y2=0
cc_259 N_A_229_483#_M1011_g N_VPWR_c_512_n 0.00490845f $X=2.485 $Y=2.625 $X2=0
+ $Y2=0
cc_260 N_A_229_483#_M1011_g N_VPWR_c_505_n 0.00506877f $X=2.485 $Y=2.625 $X2=0
+ $Y2=0
cc_261 N_A_229_483#_c_325_n N_VGND_c_561_n 9.32665e-19 $X=2.41 $Y=0.84 $X2=0
+ $Y2=0
cc_262 N_A_229_483#_c_326_n N_VGND_c_561_n 0.00334504f $X=2.11 $Y=0.84 $X2=0
+ $Y2=0
cc_263 N_A_229_483#_c_327_n N_VGND_c_561_n 0.00564615f $X=2.485 $Y=0.765 $X2=0
+ $Y2=0
cc_264 N_A_229_483#_c_330_n N_VGND_c_561_n 0.014764f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_265 N_A_229_483#_c_326_n N_VGND_c_563_n 0.00521322f $X=2.11 $Y=0.84 $X2=0
+ $Y2=0
cc_266 N_A_229_483#_c_327_n N_VGND_c_563_n 0.0118895f $X=2.485 $Y=0.765 $X2=0
+ $Y2=0
cc_267 N_A_229_483#_c_330_n N_VGND_c_563_n 0.0153934f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_268 N_A_229_483#_c_325_n N_A_512_47#_c_606_n 3.34403e-19 $X=2.41 $Y=0.84
+ $X2=0 $Y2=0
cc_269 N_A_229_483#_c_327_n N_A_512_47#_c_606_n 0.00617712f $X=2.485 $Y=0.765
+ $X2=0 $Y2=0
cc_270 N_A_229_483#_c_325_n N_A_512_47#_c_608_n 0.00396239f $X=2.41 $Y=0.84
+ $X2=0 $Y2=0
cc_271 N_B2_M1010_g N_B1_M1000_g 0.0478389f $X=2.915 $Y=0.445 $X2=0 $Y2=0
cc_272 B2 N_B1_M1000_g 4.46599e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_273 N_B2_c_419_n N_B1_c_458_n 0.0287191f $X=2.825 $Y=1.825 $X2=0 $Y2=0
cc_274 N_B2_M1008_g N_B1_c_459_n 0.0287191f $X=2.915 $Y=2.625 $X2=0 $Y2=0
cc_275 N_B2_c_415_n B1 0.00340986f $X=2.825 $Y=1.66 $X2=0 $Y2=0
cc_276 B2 B1 0.046868f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_277 N_B2_c_417_n B1 0.00269945f $X=2.825 $Y=1.32 $X2=0 $Y2=0
cc_278 N_B2_c_415_n N_B1_c_456_n 0.0287191f $X=2.825 $Y=1.66 $X2=0 $Y2=0
cc_279 B2 N_B1_c_456_n 9.70401e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_280 N_B2_M1008_g N_VPWR_c_509_n 0.00177594f $X=2.915 $Y=2.625 $X2=0 $Y2=0
cc_281 N_B2_M1008_g N_VPWR_c_512_n 0.00471331f $X=2.915 $Y=2.625 $X2=0 $Y2=0
cc_282 N_B2_M1008_g N_VPWR_c_505_n 0.00506877f $X=2.915 $Y=2.625 $X2=0 $Y2=0
cc_283 N_B2_M1010_g N_VGND_c_560_n 0.00316145f $X=2.915 $Y=0.445 $X2=0 $Y2=0
cc_284 N_B2_M1010_g N_VGND_c_561_n 0.00585385f $X=2.915 $Y=0.445 $X2=0 $Y2=0
cc_285 N_B2_M1010_g N_VGND_c_563_n 0.00619488f $X=2.915 $Y=0.445 $X2=0 $Y2=0
cc_286 N_B2_M1010_g N_A_512_47#_c_606_n 0.00187663f $X=2.915 $Y=0.445 $X2=0
+ $Y2=0
cc_287 N_B2_M1010_g N_A_512_47#_c_607_n 0.0121455f $X=2.915 $Y=0.445 $X2=0 $Y2=0
cc_288 B2 N_A_512_47#_c_607_n 0.0104103f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_289 B2 N_A_512_47#_c_608_n 0.0224564f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_290 N_B2_c_417_n N_A_512_47#_c_608_n 0.00129195f $X=2.825 $Y=1.32 $X2=0 $Y2=0
cc_291 N_B1_M1006_g N_VPWR_c_509_n 0.0121538f $X=3.275 $Y=2.625 $X2=0 $Y2=0
cc_292 N_B1_c_459_n N_VPWR_c_509_n 0.00114054f $X=3.365 $Y=2.215 $X2=0 $Y2=0
cc_293 B1 N_VPWR_c_509_n 0.0201981f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_294 N_B1_M1006_g N_VPWR_c_512_n 0.00407914f $X=3.275 $Y=2.625 $X2=0 $Y2=0
cc_295 N_B1_M1006_g N_VPWR_c_505_n 0.00425776f $X=3.275 $Y=2.625 $X2=0 $Y2=0
cc_296 N_B1_M1000_g N_VGND_c_560_n 0.00316145f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_297 N_B1_M1000_g N_VGND_c_562_n 0.00585385f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_298 N_B1_M1000_g N_VGND_c_563_n 0.00719175f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_299 N_B1_M1000_g N_A_512_47#_c_607_n 0.0133098f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_300 B1 N_A_512_47#_c_607_n 0.0398182f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_301 N_B1_c_456_n N_A_512_47#_c_607_n 6.00835e-19 $X=3.365 $Y=1.71 $X2=0 $Y2=0
cc_302 N_B1_M1000_g N_A_512_47#_c_609_n 0.00405726f $X=3.345 $Y=0.445 $X2=0
+ $Y2=0
cc_303 N_X_c_488_n N_VPWR_c_506_n 0.0161562f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_304 N_X_c_488_n N_VPWR_c_510_n 0.0173933f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_305 N_X_c_488_n N_VPWR_c_505_n 0.00998238f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_306 N_X_c_487_n N_VGND_c_563_n 0.0144905f $X=0.4 $Y=0.545 $X2=0 $Y2=0
cc_307 N_X_c_487_n N_VGND_c_564_n 0.0148629f $X=0.4 $Y=0.545 $X2=0 $Y2=0
cc_308 N_VGND_c_563_n N_A_512_47#_M1001_d 0.0023104f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_309 N_VGND_c_563_n N_A_512_47#_M1000_d 0.00221783f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_561_n N_A_512_47#_c_606_n 0.0140193f $X=3 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_563_n N_A_512_47#_c_606_n 0.0107884f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_560_n N_A_512_47#_c_607_n 0.0166313f $X=3.13 $Y=0.445 $X2=0
+ $Y2=0
cc_313 N_VGND_c_563_n N_A_512_47#_c_607_n 0.0110733f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_562_n N_A_512_47#_c_609_n 0.0164158f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_563_n N_A_512_47#_c_609_n 0.011248f $X=3.6 $Y=0 $X2=0 $Y2=0
