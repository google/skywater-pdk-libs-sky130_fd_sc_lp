* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4bb_m A B C_N D_N VGND VNB VPB VPWR X
X0 a_27_530# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_196_530# a_336_439# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_336_439# a_27_530# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_336_439# a_196_530# a_419_439# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND B a_336_439# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_336_439# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_336_439# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_419_439# a_27_530# a_491_439# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND D_N a_196_530# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_336_439# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_27_530# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_491_439# B a_593_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR D_N a_196_530# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_593_485# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
