* NGSPICE file created from sky130_fd_sc_lp__o2111a_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2111a_lp A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_232_419# A2 a_134_419# VPB phighvt w=1e+06u l=250000u
+  ad=6.2e+11p pd=5.24e+06u as=2.4e+11p ps=2.48e+06u
M1001 X a_232_419# a_708_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1002 X a_232_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=1.165e+12p ps=8.33e+06u
M1003 a_404_51# C1 a_326_51# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_232_419# D1 a_404_51# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1005 a_326_51# B1 a_29_51# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.835e+11p ps=3.03e+06u
M1006 a_708_47# a_232_419# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.709e+11p ps=2.97e+06u
M1007 a_232_419# C1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR D1 a_232_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B1 a_232_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_29_51# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_134_419# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1 a_29_51# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

