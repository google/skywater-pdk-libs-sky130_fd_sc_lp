* File: sky130_fd_sc_lp__a22oi_1.pxi.spice
* Created: Wed Sep  2 09:23:05 2020
* 
x_PM_SKY130_FD_SC_LP__A22OI_1%B2 N_B2_c_47_n N_B2_M1004_g N_B2_M1002_g B2 B2
+ N_B2_c_50_n PM_SKY130_FD_SC_LP__A22OI_1%B2
x_PM_SKY130_FD_SC_LP__A22OI_1%B1 N_B1_M1007_g N_B1_M1006_g B1 B1 N_B1_c_75_n
+ N_B1_c_76_n PM_SKY130_FD_SC_LP__A22OI_1%B1
x_PM_SKY130_FD_SC_LP__A22OI_1%A1 N_A1_M1005_g N_A1_M1003_g A1 A1 A1 A1
+ N_A1_c_112_n N_A1_c_113_n N_A1_c_114_n A1 PM_SKY130_FD_SC_LP__A22OI_1%A1
x_PM_SKY130_FD_SC_LP__A22OI_1%A2 N_A2_c_158_n N_A2_M1001_g N_A2_M1000_g A2 A2
+ N_A2_c_161_n PM_SKY130_FD_SC_LP__A22OI_1%A2
x_PM_SKY130_FD_SC_LP__A22OI_1%A_65_367# N_A_65_367#_M1002_s N_A_65_367#_M1006_d
+ N_A_65_367#_M1000_d N_A_65_367#_c_193_n N_A_65_367#_c_194_n
+ N_A_65_367#_c_200_n N_A_65_367#_c_213_p N_A_65_367#_c_202_n
+ N_A_65_367#_c_195_n N_A_65_367#_c_196_n N_A_65_367#_c_197_n
+ PM_SKY130_FD_SC_LP__A22OI_1%A_65_367#
x_PM_SKY130_FD_SC_LP__A22OI_1%Y N_Y_M1007_d N_Y_M1002_d N_Y_c_228_n N_Y_c_240_n
+ N_Y_c_235_n N_Y_c_229_n N_Y_c_236_n Y Y Y PM_SKY130_FD_SC_LP__A22OI_1%Y
x_PM_SKY130_FD_SC_LP__A22OI_1%VPWR N_VPWR_M1003_d VPWR N_VPWR_c_275_n
+ N_VPWR_c_276_n N_VPWR_c_274_n N_VPWR_c_278_n PM_SKY130_FD_SC_LP__A22OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A22OI_1%VGND N_VGND_M1004_s N_VGND_M1001_d N_VGND_c_305_n
+ N_VGND_c_306_n N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n N_VGND_c_310_n
+ VGND N_VGND_c_311_n N_VGND_c_312_n PM_SKY130_FD_SC_LP__A22OI_1%VGND
cc_1 VNB N_B2_c_47_n 0.0180716f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.295
cc_2 VNB N_B2_M1002_g 0.00146606f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_3 VNB B2 0.0284509f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B2_c_50_n 0.0486134f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.46
cc_5 VNB N_B1_M1006_g 0.00145774f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_6 VNB B1 0.005002f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_B1_c_75_n 0.032038f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=1.46
cc_8 VNB N_B1_c_76_n 0.017595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_M1003_g 0.00171994f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_10 VNB A1 0.001944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_112_n 0.0306645f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.295
cc_12 VNB N_A1_c_113_n 0.0190041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_114_n 0.00108015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_158_n 0.0208991f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.295
cc_15 VNB N_A2_M1000_g 0.00194731f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_16 VNB A2 0.0368879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_161_n 0.0659525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_228_n 0.00282534f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_Y_c_229_n 0.00224142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_274_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=1.46
cc_21 VNB N_VGND_c_305_n 0.0372931f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_VGND_c_306_n 0.0340604f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=1.46
cc_23 VNB N_VGND_c_307_n 0.0112126f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.46
cc_24 VNB N_VGND_c_308_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_309_n 0.0482447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_310_n 0.00596836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_311_n 0.0142356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_312_n 0.209251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_B2_M1002_g 0.0246393f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_30 VPB B2 0.0145386f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_31 VPB N_B1_M1006_g 0.0205742f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_32 VPB B1 0.00224104f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_33 VPB N_A1_M1003_g 0.0232733f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_34 VPB A1 0.00243051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A2_M1000_g 0.028593f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_36 VPB A2 0.0125463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_65_367#_c_193_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_65_367#_c_194_n 0.0371196f $X=-0.19 $Y=1.655 $X2=0.45 $Y2=1.46
cc_39 VPB N_A_65_367#_c_195_n 0.0148865f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.665
cc_40 VPB N_A_65_367#_c_196_n 0.0230171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_65_367#_c_197_n 0.00717518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_Y_c_228_n 0.00136759f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_43 VPB N_VPWR_c_275_n 0.0416698f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_44 VPB N_VPWR_c_276_n 0.0171493f $X=-0.19 $Y=1.655 $X2=0.45 $Y2=1.46
cc_45 VPB N_VPWR_c_274_n 0.0547623f $X=-0.19 $Y=1.655 $X2=0.45 $Y2=1.46
cc_46 VPB N_VPWR_c_278_n 0.0124205f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 N_B2_M1002_g N_B1_M1006_g 0.0365037f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_48 N_B2_c_47_n B1 4.66746e-19 $X=0.665 $Y=1.295 $X2=0 $Y2=0
cc_49 N_B2_c_50_n N_B1_c_75_n 0.0426606f $X=0.665 $Y=1.46 $X2=0 $Y2=0
cc_50 N_B2_c_47_n N_B1_c_76_n 0.0426606f $X=0.665 $Y=1.295 $X2=0 $Y2=0
cc_51 B2 N_A_65_367#_c_194_n 0.0224262f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_B2_c_50_n N_A_65_367#_c_194_n 0.00144108f $X=0.665 $Y=1.46 $X2=0 $Y2=0
cc_53 N_B2_M1002_g N_A_65_367#_c_200_n 0.0111507f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_54 N_B2_c_47_n N_Y_c_228_n 0.00924987f $X=0.665 $Y=1.295 $X2=0 $Y2=0
cc_55 N_B2_M1002_g N_Y_c_228_n 0.00987152f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_56 B2 N_Y_c_228_n 0.0403735f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_B2_c_50_n N_Y_c_228_n 0.00730885f $X=0.665 $Y=1.46 $X2=0 $Y2=0
cc_58 N_B2_c_47_n N_Y_c_235_n 0.00464098f $X=0.665 $Y=1.295 $X2=0 $Y2=0
cc_59 N_B2_M1002_g N_Y_c_236_n 0.0123534f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_60 N_B2_M1002_g N_VPWR_c_275_n 0.00357877f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_61 N_B2_M1002_g N_VPWR_c_274_n 0.00644799f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_62 N_B2_c_47_n N_VGND_c_305_n 0.00483749f $X=0.665 $Y=1.295 $X2=0 $Y2=0
cc_63 B2 N_VGND_c_305_n 0.022426f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_64 N_B2_c_50_n N_VGND_c_305_n 0.0015759f $X=0.665 $Y=1.46 $X2=0 $Y2=0
cc_65 N_B2_c_47_n N_VGND_c_309_n 0.00482246f $X=0.665 $Y=1.295 $X2=0 $Y2=0
cc_66 N_B2_c_47_n N_VGND_c_312_n 0.00867022f $X=0.665 $Y=1.295 $X2=0 $Y2=0
cc_67 N_B1_M1006_g N_A1_M1003_g 0.0302518f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_68 N_B1_c_76_n A1 5.50431e-19 $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_69 B1 A1 0.0319764f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_70 N_B1_c_75_n A1 3.08006e-19 $X=1.13 $Y=1.46 $X2=0 $Y2=0
cc_71 N_B1_c_75_n N_A1_c_112_n 0.0205893f $X=1.13 $Y=1.46 $X2=0 $Y2=0
cc_72 B1 N_A1_c_113_n 0.00333976f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_73 N_B1_c_76_n N_A1_c_113_n 0.0180895f $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_74 B1 N_A1_c_114_n 0.0103827f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_75 N_B1_c_76_n N_A1_c_114_n 5.87509e-19 $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_76 N_B1_M1006_g N_A_65_367#_c_200_n 0.011368f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_77 N_B1_M1006_g N_Y_c_228_n 0.00404985f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_78 B1 N_Y_c_228_n 0.0402635f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B1_c_76_n N_Y_c_228_n 0.0060627f $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_80 B1 N_Y_c_240_n 0.0235232f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_81 N_B1_c_75_n N_Y_c_240_n 0.00105055f $X=1.13 $Y=1.46 $X2=0 $Y2=0
cc_82 N_B1_c_76_n N_Y_c_240_n 0.0149115f $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_83 N_B1_c_76_n N_Y_c_229_n 0.00729656f $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_84 N_B1_M1006_g N_Y_c_236_n 0.0123441f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_85 N_B1_c_75_n N_Y_c_236_n 0.00175681f $X=1.13 $Y=1.46 $X2=0 $Y2=0
cc_86 N_B1_M1006_g Y 0.0125596f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_87 B1 Y 0.0220648f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B1_c_75_n Y 5.51443e-19 $X=1.13 $Y=1.46 $X2=0 $Y2=0
cc_89 N_B1_M1006_g N_VPWR_c_275_n 0.00357877f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_90 N_B1_M1006_g N_VPWR_c_274_n 0.00553095f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B1_M1006_g N_VPWR_c_278_n 0.00106633f $X=1.095 $Y=2.465 $X2=0 $Y2=0
cc_92 N_B1_c_76_n N_VGND_c_309_n 0.00482246f $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_93 N_B1_c_76_n N_VGND_c_312_n 0.0051802f $X=1.122 $Y=1.295 $X2=0 $Y2=0
cc_94 A1 N_A2_c_158_n 0.00724778f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_95 N_A1_c_113_n N_A2_c_158_n 0.0290128f $X=1.67 $Y=1.295 $X2=-0.19 $Y2=-0.245
cc_96 N_A1_c_114_n N_A2_c_158_n 0.0029989f $X=1.682 $Y=1.342 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A1_M1003_g N_A2_M1000_g 0.02025f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_98 A1 N_A2_M1000_g 2.97473e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A1_M1003_g A2 3.89186e-19 $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_100 A1 A2 0.0359129f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A1_c_112_n A2 0.00122263f $X=1.67 $Y=1.46 $X2=0 $Y2=0
cc_102 N_A1_c_113_n A2 2.34757e-19 $X=1.67 $Y=1.295 $X2=0 $Y2=0
cc_103 N_A1_c_114_n A2 0.0116265f $X=1.682 $Y=1.342 $X2=0 $Y2=0
cc_104 A1 N_A2_c_161_n 8.55195e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A1_c_112_n N_A2_c_161_n 0.0214885f $X=1.67 $Y=1.46 $X2=0 $Y2=0
cc_106 N_A1_M1003_g N_A_65_367#_c_202_n 0.0110757f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A1_c_114_n N_Y_c_228_n 8.01339e-19 $X=1.682 $Y=1.342 $X2=0 $Y2=0
cc_108 A1 N_Y_c_240_n 0.0145292f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_109 A1 N_Y_c_229_n 0.0360309f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_110 N_A1_c_113_n N_Y_c_229_n 0.0022412f $X=1.67 $Y=1.295 $X2=0 $Y2=0
cc_111 N_A1_M1003_g N_Y_c_236_n 7.37186e-19 $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A1_M1003_g Y 0.0143794f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_113 A1 Y 0.0240632f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_114 N_A1_c_112_n Y 8.39197e-19 $X=1.67 $Y=1.46 $X2=0 $Y2=0
cc_115 N_A1_M1003_g N_VPWR_c_275_n 0.00487821f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A1_M1003_g N_VPWR_c_274_n 0.00473514f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A1_M1003_g N_VPWR_c_278_n 0.0136185f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_118 A1 N_VGND_c_306_n 0.0266803f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A1_c_113_n N_VGND_c_306_n 0.0013162f $X=1.67 $Y=1.295 $X2=0 $Y2=0
cc_120 A1 N_VGND_c_309_n 0.00790735f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A1_c_113_n N_VGND_c_309_n 0.00401979f $X=1.67 $Y=1.295 $X2=0 $Y2=0
cc_122 A1 N_VGND_c_312_n 0.00782639f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A1_c_113_n N_VGND_c_312_n 0.00715176f $X=1.67 $Y=1.295 $X2=0 $Y2=0
cc_124 A1 A_331_69# 0.00993848f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_125 N_A1_c_114_n A_331_69# 0.00258727f $X=1.682 $Y=1.342 $X2=-0.19 $Y2=-0.245
cc_126 N_A2_M1000_g N_A_65_367#_c_202_n 0.012257f $X=2.35 $Y=2.465 $X2=0 $Y2=0
cc_127 A2 N_A_65_367#_c_202_n 0.00455279f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A2_c_161_n N_A_65_367#_c_202_n 2.05858e-19 $X=2.55 $Y=1.46 $X2=0 $Y2=0
cc_129 N_A2_M1000_g N_A_65_367#_c_195_n 0.00941554f $X=2.35 $Y=2.465 $X2=0 $Y2=0
cc_130 A2 N_A_65_367#_c_195_n 0.0255384f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A2_c_161_n N_A_65_367#_c_195_n 0.00155535f $X=2.55 $Y=1.46 $X2=0 $Y2=0
cc_132 N_A2_M1000_g N_A_65_367#_c_197_n 5.71016e-19 $X=2.35 $Y=2.465 $X2=0 $Y2=0
cc_133 A2 Y 0.0179252f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A2_c_161_n Y 9.89558e-19 $X=2.55 $Y=1.46 $X2=0 $Y2=0
cc_135 N_A2_M1000_g N_VPWR_c_276_n 0.00487821f $X=2.35 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_M1000_g N_VPWR_c_274_n 0.00556317f $X=2.35 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A2_M1000_g N_VPWR_c_278_n 0.0141009f $X=2.35 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A2_c_158_n N_VGND_c_306_n 0.0163463f $X=2.12 $Y=1.295 $X2=0 $Y2=0
cc_139 A2 N_VGND_c_306_n 0.0225959f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A2_c_161_n N_VGND_c_306_n 0.00175224f $X=2.55 $Y=1.46 $X2=0 $Y2=0
cc_141 N_A2_c_158_n N_VGND_c_309_n 0.00400407f $X=2.12 $Y=1.295 $X2=0 $Y2=0
cc_142 N_A2_c_158_n N_VGND_c_312_n 0.00780677f $X=2.12 $Y=1.295 $X2=0 $Y2=0
cc_143 N_A_65_367#_c_200_n N_Y_M1002_d 0.00332344f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_144 N_A_65_367#_c_200_n N_Y_c_236_n 0.016693f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_145 N_A_65_367#_M1006_d Y 0.00741718f $X=1.17 $Y=1.835 $X2=0 $Y2=0
cc_146 N_A_65_367#_c_213_p Y 0.0182397f $X=1.337 $Y=2.47 $X2=0 $Y2=0
cc_147 N_A_65_367#_c_202_n Y 0.047645f $X=2.415 $Y=2.385 $X2=0 $Y2=0
cc_148 N_A_65_367#_c_202_n N_VPWR_M1003_d 0.0129036f $X=2.415 $Y=2.385 $X2=-0.19
+ $Y2=1.655
cc_149 N_A_65_367#_c_193_n N_VPWR_c_275_n 0.0175634f $X=0.41 $Y=2.905 $X2=0
+ $Y2=0
cc_150 N_A_65_367#_c_200_n N_VPWR_c_275_n 0.0528605f $X=1.215 $Y=2.99 $X2=0
+ $Y2=0
cc_151 N_A_65_367#_c_196_n N_VPWR_c_276_n 0.0178111f $X=2.565 $Y=2.505 $X2=0
+ $Y2=0
cc_152 N_A_65_367#_M1002_s N_VPWR_c_274_n 0.00215162f $X=0.325 $Y=1.835 $X2=0
+ $Y2=0
cc_153 N_A_65_367#_M1006_d N_VPWR_c_274_n 0.0029829f $X=1.17 $Y=1.835 $X2=0
+ $Y2=0
cc_154 N_A_65_367#_M1000_d N_VPWR_c_274_n 0.00244787f $X=2.425 $Y=1.835 $X2=0
+ $Y2=0
cc_155 N_A_65_367#_c_193_n N_VPWR_c_274_n 0.00970886f $X=0.41 $Y=2.905 $X2=0
+ $Y2=0
cc_156 N_A_65_367#_c_200_n N_VPWR_c_274_n 0.033577f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_157 N_A_65_367#_c_202_n N_VPWR_c_274_n 0.00999856f $X=2.415 $Y=2.385 $X2=0
+ $Y2=0
cc_158 N_A_65_367#_c_196_n N_VPWR_c_274_n 0.0100304f $X=2.565 $Y=2.505 $X2=0
+ $Y2=0
cc_159 N_A_65_367#_c_197_n N_VPWR_c_274_n 0.00194326f $X=2.572 $Y=2.385 $X2=0
+ $Y2=0
cc_160 N_A_65_367#_c_202_n N_VPWR_c_278_n 0.0438303f $X=2.415 $Y=2.385 $X2=0
+ $Y2=0
cc_161 Y N_VPWR_M1003_d 0.0194525f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_162 N_Y_M1002_d N_VPWR_c_274_n 0.00225186f $X=0.74 $Y=1.835 $X2=0 $Y2=0
cc_163 N_Y_c_229_n N_VGND_c_305_n 0.00735592f $X=1.33 $Y=0.49 $X2=0 $Y2=0
cc_164 N_Y_c_229_n N_VGND_c_309_n 0.0103515f $X=1.33 $Y=0.49 $X2=0 $Y2=0
cc_165 N_Y_c_240_n N_VGND_c_312_n 0.0101598f $X=1.205 $Y=0.95 $X2=0 $Y2=0
cc_166 N_Y_c_235_n N_VGND_c_312_n 0.00631872f $X=0.875 $Y=0.95 $X2=0 $Y2=0
cc_167 N_Y_c_229_n N_VGND_c_312_n 0.00780843f $X=1.33 $Y=0.49 $X2=0 $Y2=0
cc_168 N_Y_c_228_n A_148_69# 0.00160653f $X=0.79 $Y=1.92 $X2=-0.19 $Y2=-0.245
cc_169 N_Y_c_240_n A_148_69# 0.00100313f $X=1.205 $Y=0.95 $X2=-0.19 $Y2=-0.245
cc_170 N_Y_c_235_n A_148_69# 0.00188384f $X=0.875 $Y=0.95 $X2=-0.19 $Y2=-0.245
