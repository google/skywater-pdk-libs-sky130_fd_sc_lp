* NGSPICE file created from sky130_fd_sc_lp__and4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4b_1 A_N B C D VGND VNB VPB VPWR X
M1000 X a_215_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=8.463e+11p ps=7.17e+06u
M1001 a_300_47# a_27_49# a_215_367# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1002 VPWR B a_215_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1003 a_372_47# B a_300_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_444_47# C a_372_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 VGND A_N a_27_49# VNB nshort w=420000u l=150000u
+  ad=4.977e+11p pd=4.36e+06u as=1.113e+11p ps=1.37e+06u
M1006 X a_215_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1007 VPWR D a_215_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_215_367# a_27_49# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_215_367# C VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A_N a_27_49# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 VGND D a_444_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

