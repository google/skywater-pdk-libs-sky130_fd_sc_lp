* File: sky130_fd_sc_lp__buflp_m.pex.spice
* Created: Fri Aug 28 10:12:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFLP_M%A_90_94# 1 2 9 13 17 21 25 29 33 36 37 38
c60 21 0 1.43438e-19 $X=0.915 $Y=2.66
r61 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.825
+ $Y=1.375 $X2=0.825 $Y2=1.375
r62 31 38 2.70057 $w=3.55e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.09 $Y=1.38
+ $X2=1.985 $Y2=1.295
r63 31 33 59.0051 $w=2.48e-07 $l=1.28e-06 $layer=LI1_cond $X=2.09 $Y=1.38
+ $X2=2.09 $Y2=2.66
r64 27 38 2.70057 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=1.21
+ $X2=1.985 $Y2=1.295
r65 27 29 10.4007 $w=4.58e-07 $l=4e-07 $layer=LI1_cond $X=1.985 $Y=1.21
+ $X2=1.985 $Y2=0.81
r66 26 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=1.295
+ $X2=0.825 $Y2=1.295
r67 25 38 4.08752 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.755 $Y=1.295
+ $X2=1.985 $Y2=1.295
r68 25 26 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.755 $Y=1.295
+ $X2=0.99 $Y2=1.295
r69 19 37 92.2311 $w=2.7e-07 $l=5.94559e-07 $layer=POLY_cond $X=0.915 $Y=1.88
+ $X2=0.72 $Y2=1.375
r70 19 21 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.915 $Y=1.88
+ $X2=0.915 $Y2=2.66
r71 15 37 31.5348 $w=2.7e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.885 $Y=1.21
+ $X2=0.72 $Y2=1.375
r72 15 17 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.885 $Y=1.21
+ $X2=0.885 $Y2=0.81
r73 11 37 92.2311 $w=2.7e-07 $l=5.94559e-07 $layer=POLY_cond $X=0.525 $Y=1.88
+ $X2=0.72 $Y2=1.375
r74 11 13 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.525 $Y=1.88
+ $X2=0.525 $Y2=2.66
r75 7 37 31.5348 $w=2.7e-07 $l=1.95e-07 $layer=POLY_cond $X=0.525 $Y=1.375
+ $X2=0.72 $Y2=1.375
r76 7 9 205.106 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.525 $Y=1.375
+ $X2=0.525 $Y2=0.81
r77 2 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=2.45 $X2=2.05 $Y2=2.66
r78 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.78
+ $Y=0.6 $X2=1.92 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_M%A 3 7 11 15 17 18 19 20 26
c42 17 0 1.43438e-19 $X=1.68 $Y=1.665
r43 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=2.405
+ $X2=1.63 $Y2=2.775
r44 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=2.035
+ $X2=1.63 $Y2=2.405
r45 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=2.035
r46 17 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.715 $X2=1.63 $Y2=1.715
r47 13 26 88.1262 $w=2.84e-07 $l=6.2155e-07 $layer=POLY_cond $X=1.835 $Y=2.22
+ $X2=1.575 $Y2=1.715
r48 13 15 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.835 $Y=2.22
+ $X2=1.835 $Y2=2.66
r49 9 26 30.422 $w=2.84e-07 $l=2.20624e-07 $layer=POLY_cond $X=1.705 $Y=1.55
+ $X2=1.575 $Y2=1.715
r50 9 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.705 $Y=1.55
+ $X2=1.705 $Y2=0.81
r51 5 26 88.1262 $w=2.84e-07 $l=5.66282e-07 $layer=POLY_cond $X=1.445 $Y=2.22
+ $X2=1.575 $Y2=1.715
r52 5 7 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.445 $Y=2.22
+ $X2=1.445 $Y2=2.66
r53 1 26 30.422 $w=2.84e-07 $l=3.32415e-07 $layer=POLY_cond $X=1.315 $Y=1.55
+ $X2=1.575 $Y2=1.715
r54 1 3 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.315 $Y=1.55
+ $X2=1.315 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_M%X 1 2 7 8 9 10 11 12 13
r14 13 37 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.3 $Y=2.775 $X2=0.3
+ $Y2=2.66
r15 12 37 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.3 $Y=2.405
+ $X2=0.3 $Y2=2.66
r16 11 12 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=2.035 $X2=0.3
+ $Y2=2.405
r17 10 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=1.665 $X2=0.3
+ $Y2=2.035
r18 9 10 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=1.295 $X2=0.3
+ $Y2=1.665
r19 8 9 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=0.925 $X2=0.3
+ $Y2=1.295
r20 8 25 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.3 $Y=0.925 $X2=0.3
+ $Y2=0.81
r21 7 25 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.3 $Y=0.555 $X2=0.3
+ $Y2=0.81
r22 2 37 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.45 $X2=0.31 $Y2=2.66
r23 1 25 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.6 $X2=0.31 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_M%VPWR 1 6 8 10 17 18 21
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=3.33
+ $X2=1.13 $Y2=3.33
r28 15 17 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.295 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.13 $Y2=3.33
r31 10 12 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r33 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.72
+ $Y2=3.33
r34 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=3.245 $X2=1.13
+ $Y2=3.33
r36 4 6 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=2.66
r37 1 6 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=2.45 $X2=1.13 $Y2=2.66
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_M%VGND 1 6 8 10 17 18 21
r26 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r28 15 17 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=2.16
+ $Y2=0
r29 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r31 10 12 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.72
+ $Y2=0
r32 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r33 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r34 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r36 4 6 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0.81
r37 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.6 $X2=1.1 $Y2=0.81
.ends

