* File: sky130_fd_sc_lp__or3_lp.pxi.spice
* Created: Wed Sep  2 10:30:49 2020
* 
x_PM_SKY130_FD_SC_LP__OR3_LP%A_108_31# N_A_108_31#_M1010_d N_A_108_31#_M1004_d
+ N_A_108_31#_M1006_d N_A_108_31#_M1008_g N_A_108_31#_c_76_n N_A_108_31#_c_77_n
+ N_A_108_31#_c_91_n N_A_108_31#_M1005_g N_A_108_31#_M1001_g N_A_108_31#_c_79_n
+ N_A_108_31#_c_80_n N_A_108_31#_c_81_n N_A_108_31#_c_82_n N_A_108_31#_c_83_n
+ N_A_108_31#_c_84_n N_A_108_31#_c_85_n N_A_108_31#_c_86_n N_A_108_31#_c_87_n
+ N_A_108_31#_c_88_n N_A_108_31#_c_94_n N_A_108_31#_c_89_n N_A_108_31#_c_90_n
+ PM_SKY130_FD_SC_LP__OR3_LP%A_108_31#
x_PM_SKY130_FD_SC_LP__OR3_LP%A N_A_c_184_n N_A_M1009_g N_A_c_185_n N_A_c_186_n
+ N_A_c_187_n N_A_M1010_g N_A_c_188_n N_A_c_194_n N_A_M1007_g N_A_c_189_n A A A
+ A N_A_c_190_n N_A_c_191_n N_A_c_192_n PM_SKY130_FD_SC_LP__OR3_LP%A
x_PM_SKY130_FD_SC_LP__OR3_LP%B N_B_c_249_n N_B_M1002_g N_B_c_250_n N_B_c_251_n
+ N_B_M1000_g N_B_c_252_n N_B_M1011_g N_B_c_253_n N_B_c_254_n N_B_c_255_n
+ N_B_c_260_n B B B B N_B_c_256_n N_B_c_257_n PM_SKY130_FD_SC_LP__OR3_LP%B
x_PM_SKY130_FD_SC_LP__OR3_LP%C N_C_c_309_n N_C_M1003_g N_C_M1006_g N_C_c_310_n
+ N_C_M1004_g N_C_c_311_n N_C_c_312_n N_C_c_313_n N_C_c_318_n C N_C_c_314_n
+ N_C_c_315_n PM_SKY130_FD_SC_LP__OR3_LP%C
x_PM_SKY130_FD_SC_LP__OR3_LP%X N_X_M1008_s N_X_M1005_s X X X X X X X N_X_c_357_n
+ PM_SKY130_FD_SC_LP__OR3_LP%X
x_PM_SKY130_FD_SC_LP__OR3_LP%VPWR N_VPWR_M1005_d N_VPWR_c_378_n VPWR
+ N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_377_n N_VPWR_c_382_n
+ PM_SKY130_FD_SC_LP__OR3_LP%VPWR
x_PM_SKY130_FD_SC_LP__OR3_LP%VGND N_VGND_M1001_d N_VGND_M1011_d N_VGND_c_409_n
+ N_VGND_c_410_n VGND N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n
+ N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n PM_SKY130_FD_SC_LP__OR3_LP%VGND
cc_1 VNB N_A_108_31#_M1008_g 0.0384442f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.495
cc_2 VNB N_A_108_31#_c_76_n 0.00977956f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.245
cc_3 VNB N_A_108_31#_c_77_n 0.0109496f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.245
cc_4 VNB N_A_108_31#_M1001_g 0.0336192f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.495
cc_5 VNB N_A_108_31#_c_79_n 0.00393417f $X=-0.19 $Y=-0.245 $X2=1.127 $Y2=1.613
cc_6 VNB N_A_108_31#_c_80_n 0.0188054f $X=-0.19 $Y=-0.245 $X2=1.127 $Y2=1.245
cc_7 VNB N_A_108_31#_c_81_n 0.00160059f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.335
cc_8 VNB N_A_108_31#_c_82_n 0.0272582f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.335
cc_9 VNB N_A_108_31#_c_83_n 0.00837335f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=0.95
cc_10 VNB N_A_108_31#_c_84_n 0.00255387f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.95
cc_11 VNB N_A_108_31#_c_85_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.495
cc_12 VNB N_A_108_31#_c_86_n 0.0214043f $X=-0.19 $Y=-0.245 $X2=3.395 $Y2=0.95
cc_13 VNB N_A_108_31#_c_87_n 0.0256923f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.495
cc_14 VNB N_A_108_31#_c_88_n 0.00200962f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.95
cc_15 VNB N_A_108_31#_c_89_n 0.0296144f $X=-0.19 $Y=-0.245 $X2=3.487 $Y2=2.065
cc_16 VNB N_A_108_31#_c_90_n 0.014226f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.95
cc_17 VNB N_A_c_184_n 0.0138865f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.285
cc_18 VNB N_A_c_185_n 0.0100944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_c_186_n 0.00876493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_187_n 0.0137713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_188_n 0.0172809f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.495
cc_22 VNB N_A_c_189_n 0.00437176f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.965
cc_23 VNB N_A_c_190_n 0.0239877f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.495
cc_24 VNB N_A_c_191_n 0.0102402f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.495
cc_25 VNB N_A_c_192_n 0.0193716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_249_n 0.0137713f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.285
cc_27 VNB N_B_c_250_n 0.00901152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_251_n 0.00862406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_c_252_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.495
cc_30 VNB N_B_c_253_n 0.00568287f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.245
cc_31 VNB N_B_c_254_n 0.0183459f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.545
cc_32 VNB N_B_c_255_n 0.0203691f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.545
cc_33 VNB N_B_c_256_n 0.0169853f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.335
cc_34 VNB N_B_c_257_n 0.00163377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C_c_309_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.285
cc_36 VNB N_C_c_310_n 0.0175316f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.17
cc_37 VNB N_C_c_311_n 0.0235553f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.965
cc_38 VNB N_C_c_312_n 0.0193953f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.17
cc_39 VNB N_C_c_313_n 0.0195165f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.495
cc_40 VNB N_C_c_314_n 0.0141684f $X=-0.19 $Y=-0.245 $X2=1.127 $Y2=1.245
cc_41 VNB N_C_c_315_n 0.00428838f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.035
cc_42 VNB X 0.0497339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_357_n 0.0286364f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.495
cc_44 VNB N_VPWR_c_377_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.127 $Y2=1.613
cc_45 VNB N_VGND_c_409_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_410_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_411_n 0.0281509f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.545
cc_48 VNB N_VGND_c_412_n 0.0352526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_413_n 0.0271986f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.335
cc_50 VNB N_VGND_c_414_n 0.243774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_415_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.865
cc_52 VNB N_VGND_c_416_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_A_108_31#_c_91_n 0.0266708f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.965
cc_54 VPB N_A_108_31#_c_79_n 0.0379886f $X=-0.19 $Y=1.655 $X2=1.127 $Y2=1.613
cc_55 VPB N_A_108_31#_c_81_n 0.00274039f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=1.335
cc_56 VPB N_A_108_31#_c_94_n 0.0483921f $X=-0.19 $Y=1.655 $X2=3.415 $Y2=2.23
cc_57 VPB N_A_108_31#_c_89_n 0.0197367f $X=-0.19 $Y=1.655 $X2=3.487 $Y2=2.065
cc_58 VPB N_A_c_188_n 0.0367997f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.495
cc_59 VPB N_A_c_194_n 0.0202769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_c_191_n 0.00666239f $X=-0.19 $Y=1.655 $X2=1.98 $Y2=0.495
cc_61 VPB N_B_M1000_g 0.0253196f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.17
cc_62 VPB N_B_c_255_n 0.00475774f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.545
cc_63 VPB N_B_c_260_n 0.014521f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.17
cc_64 VPB N_B_c_257_n 0.00175682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_C_M1006_g 0.0310133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_C_c_313_n 0.0045586f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.495
cc_67 VPB N_C_c_318_n 0.0140076f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=0.495
cc_68 VPB N_C_c_315_n 0.00308283f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=1.035
cc_69 VPB X 0.0870256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_378_n 0.00731138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_379_n 0.0280556f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.495
cc_72 VPB N_VPWR_c_380_n 0.069426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_377_n 0.084531f $X=-0.19 $Y=1.655 $X2=1.127 $Y2=1.613
cc_74 VPB N_VPWR_c_382_n 0.00548753f $X=-0.19 $Y=1.655 $X2=1.19 $Y2=1.035
cc_75 N_A_108_31#_M1001_g N_A_c_184_n 0.0181569f $X=0.975 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_108_31#_c_85_n N_A_c_184_n 0.00161464f $X=1.98 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A_108_31#_c_83_n N_A_c_185_n 0.0135868f $X=1.815 $Y=0.95 $X2=0 $Y2=0
cc_78 N_A_108_31#_c_80_n N_A_c_186_n 0.00139458f $X=1.127 $Y=1.245 $X2=0 $Y2=0
cc_79 N_A_108_31#_c_83_n N_A_c_186_n 0.00825744f $X=1.815 $Y=0.95 $X2=0 $Y2=0
cc_80 N_A_108_31#_c_84_n N_A_c_186_n 0.00154334f $X=1.355 $Y=0.95 $X2=0 $Y2=0
cc_81 N_A_108_31#_c_85_n N_A_c_187_n 0.00995781f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_82 N_A_108_31#_c_79_n N_A_c_188_n 0.00852381f $X=1.127 $Y=1.613 $X2=0 $Y2=0
cc_83 N_A_108_31#_c_83_n N_A_c_189_n 0.00623175f $X=1.815 $Y=0.95 $X2=0 $Y2=0
cc_84 N_A_108_31#_c_85_n N_A_c_189_n 0.00495788f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_85 N_A_108_31#_c_88_n N_A_c_189_n 9.26094e-19 $X=1.98 $Y=0.95 $X2=0 $Y2=0
cc_86 N_A_108_31#_c_81_n N_A_c_190_n 6.55437e-19 $X=1.19 $Y=1.335 $X2=0 $Y2=0
cc_87 N_A_108_31#_c_82_n N_A_c_190_n 0.00791004f $X=1.19 $Y=1.335 $X2=0 $Y2=0
cc_88 N_A_108_31#_c_88_n N_A_c_190_n 0.00213629f $X=1.98 $Y=0.95 $X2=0 $Y2=0
cc_89 N_A_108_31#_c_91_n N_A_c_191_n 0.00164974f $X=0.945 $Y=1.965 $X2=0 $Y2=0
cc_90 N_A_108_31#_c_79_n N_A_c_191_n 0.00523151f $X=1.127 $Y=1.613 $X2=0 $Y2=0
cc_91 N_A_108_31#_c_80_n N_A_c_191_n 0.00509944f $X=1.127 $Y=1.245 $X2=0 $Y2=0
cc_92 N_A_108_31#_c_81_n N_A_c_191_n 0.0449198f $X=1.19 $Y=1.335 $X2=0 $Y2=0
cc_93 N_A_108_31#_c_83_n N_A_c_191_n 0.0191162f $X=1.815 $Y=0.95 $X2=0 $Y2=0
cc_94 N_A_108_31#_c_86_n N_A_c_191_n 0.0104251f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_95 N_A_108_31#_c_88_n N_A_c_191_n 0.0281935f $X=1.98 $Y=0.95 $X2=0 $Y2=0
cc_96 N_A_108_31#_M1001_g N_A_c_192_n 0.00279516f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_97 N_A_108_31#_c_80_n N_A_c_192_n 0.00791004f $X=1.127 $Y=1.245 $X2=0 $Y2=0
cc_98 N_A_108_31#_c_81_n N_A_c_192_n 0.0032112f $X=1.19 $Y=1.335 $X2=0 $Y2=0
cc_99 N_A_108_31#_c_83_n N_A_c_192_n 0.00499491f $X=1.815 $Y=0.95 $X2=0 $Y2=0
cc_100 N_A_108_31#_c_88_n N_A_c_192_n 0.00264924f $X=1.98 $Y=0.95 $X2=0 $Y2=0
cc_101 N_A_108_31#_c_85_n N_B_c_249_n 0.00995781f $X=1.98 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_108_31#_c_86_n N_B_c_250_n 0.0119384f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_103 N_A_108_31#_c_85_n N_B_c_251_n 0.00495788f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_104 N_A_108_31#_c_86_n N_B_c_251_n 0.00825744f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_105 N_A_108_31#_c_88_n N_B_c_251_n 0.00133508f $X=1.98 $Y=0.95 $X2=0 $Y2=0
cc_106 N_A_108_31#_c_94_n N_B_M1000_g 0.00144468f $X=3.415 $Y=2.23 $X2=0 $Y2=0
cc_107 N_A_108_31#_c_85_n N_B_c_252_n 0.00161464f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_108 N_A_108_31#_c_86_n N_B_c_253_n 0.00899008f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_109 N_A_108_31#_c_86_n N_B_c_254_n 0.00718962f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_110 N_A_108_31#_c_86_n N_B_c_256_n 0.00113819f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_111 N_A_108_31#_c_86_n N_B_c_257_n 0.0245349f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_112 N_A_108_31#_c_94_n N_B_c_257_n 0.0301513f $X=3.415 $Y=2.23 $X2=0 $Y2=0
cc_113 N_A_108_31#_c_87_n N_C_c_309_n 0.00161464f $X=3.56 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_108_31#_c_94_n N_C_M1006_g 0.0265254f $X=3.415 $Y=2.23 $X2=0 $Y2=0
cc_115 N_A_108_31#_c_89_n N_C_M1006_g 0.00418088f $X=3.487 $Y=2.065 $X2=0 $Y2=0
cc_116 N_A_108_31#_c_87_n N_C_c_310_n 0.0110144f $X=3.56 $Y=0.495 $X2=0 $Y2=0
cc_117 N_A_108_31#_c_86_n N_C_c_311_n 0.0278107f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_118 N_A_108_31#_c_87_n N_C_c_311_n 0.00565463f $X=3.56 $Y=0.495 $X2=0 $Y2=0
cc_119 N_A_108_31#_c_90_n N_C_c_311_n 0.00187523f $X=3.56 $Y=0.95 $X2=0 $Y2=0
cc_120 N_A_108_31#_c_86_n N_C_c_312_n 0.0075525f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_121 N_A_108_31#_c_89_n N_C_c_312_n 0.00354853f $X=3.487 $Y=2.065 $X2=0 $Y2=0
cc_122 N_A_108_31#_c_94_n N_C_c_318_n 4.35446e-19 $X=3.415 $Y=2.23 $X2=0 $Y2=0
cc_123 N_A_108_31#_c_86_n N_C_c_314_n 5.68334e-19 $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_124 N_A_108_31#_c_89_n N_C_c_314_n 0.0146902f $X=3.487 $Y=2.065 $X2=0 $Y2=0
cc_125 N_A_108_31#_c_86_n N_C_c_315_n 0.0261167f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_126 N_A_108_31#_c_94_n N_C_c_315_n 0.00603187f $X=3.415 $Y=2.23 $X2=0 $Y2=0
cc_127 N_A_108_31#_c_89_n N_C_c_315_n 0.0447009f $X=3.487 $Y=2.065 $X2=0 $Y2=0
cc_128 N_A_108_31#_M1008_g X 0.0152842f $X=0.615 $Y=0.495 $X2=0 $Y2=0
cc_129 N_A_108_31#_c_76_n X 0.00878913f $X=0.9 $Y=1.245 $X2=0 $Y2=0
cc_130 N_A_108_31#_c_77_n X 0.00913756f $X=0.69 $Y=1.245 $X2=0 $Y2=0
cc_131 N_A_108_31#_c_91_n X 0.0241241f $X=0.945 $Y=1.965 $X2=0 $Y2=0
cc_132 N_A_108_31#_M1001_g X 0.00419244f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_133 N_A_108_31#_c_79_n X 0.00949672f $X=1.127 $Y=1.613 $X2=0 $Y2=0
cc_134 N_A_108_31#_c_81_n X 0.0642112f $X=1.19 $Y=1.335 $X2=0 $Y2=0
cc_135 N_A_108_31#_c_82_n X 0.0149008f $X=1.19 $Y=1.335 $X2=0 $Y2=0
cc_136 N_A_108_31#_c_84_n X 0.0145108f $X=1.355 $Y=0.95 $X2=0 $Y2=0
cc_137 N_A_108_31#_M1008_g N_X_c_357_n 0.0152173f $X=0.615 $Y=0.495 $X2=0 $Y2=0
cc_138 N_A_108_31#_M1001_g N_X_c_357_n 0.00422733f $X=0.975 $Y=0.495 $X2=0 $Y2=0
cc_139 N_A_108_31#_c_91_n N_VPWR_c_378_n 0.0249818f $X=0.945 $Y=1.965 $X2=0
+ $Y2=0
cc_140 N_A_108_31#_c_79_n N_VPWR_c_378_n 0.00220014f $X=1.127 $Y=1.613 $X2=0
+ $Y2=0
cc_141 N_A_108_31#_c_81_n N_VPWR_c_378_n 0.0256417f $X=1.19 $Y=1.335 $X2=0 $Y2=0
cc_142 N_A_108_31#_c_91_n N_VPWR_c_379_n 0.00769046f $X=0.945 $Y=1.965 $X2=0
+ $Y2=0
cc_143 N_A_108_31#_c_94_n N_VPWR_c_380_n 0.0318087f $X=3.415 $Y=2.23 $X2=0 $Y2=0
cc_144 N_A_108_31#_c_91_n N_VPWR_c_377_n 0.0143431f $X=0.945 $Y=1.965 $X2=0
+ $Y2=0
cc_145 N_A_108_31#_c_94_n N_VPWR_c_377_n 0.0181913f $X=3.415 $Y=2.23 $X2=0 $Y2=0
cc_146 N_A_108_31#_M1008_g N_VGND_c_409_n 0.00152856f $X=0.615 $Y=0.495 $X2=0
+ $Y2=0
cc_147 N_A_108_31#_M1001_g N_VGND_c_409_n 0.0100628f $X=0.975 $Y=0.495 $X2=0
+ $Y2=0
cc_148 N_A_108_31#_c_80_n N_VGND_c_409_n 9.53999e-19 $X=1.127 $Y=1.245 $X2=0
+ $Y2=0
cc_149 N_A_108_31#_c_84_n N_VGND_c_409_n 0.0228841f $X=1.355 $Y=0.95 $X2=0 $Y2=0
cc_150 N_A_108_31#_c_85_n N_VGND_c_409_n 0.0140521f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_151 N_A_108_31#_c_85_n N_VGND_c_410_n 0.0140521f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_152 N_A_108_31#_c_86_n N_VGND_c_410_n 0.0207959f $X=3.395 $Y=0.95 $X2=0 $Y2=0
cc_153 N_A_108_31#_c_87_n N_VGND_c_410_n 0.0140521f $X=3.56 $Y=0.495 $X2=0 $Y2=0
cc_154 N_A_108_31#_M1008_g N_VGND_c_411_n 0.00352123f $X=0.615 $Y=0.495 $X2=0
+ $Y2=0
cc_155 N_A_108_31#_M1001_g N_VGND_c_411_n 0.00445056f $X=0.975 $Y=0.495 $X2=0
+ $Y2=0
cc_156 N_A_108_31#_c_85_n N_VGND_c_412_n 0.021949f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_157 N_A_108_31#_c_87_n N_VGND_c_413_n 0.0220321f $X=3.56 $Y=0.495 $X2=0 $Y2=0
cc_158 N_A_108_31#_M1008_g N_VGND_c_414_n 0.00560636f $X=0.615 $Y=0.495 $X2=0
+ $Y2=0
cc_159 N_A_108_31#_M1001_g N_VGND_c_414_n 0.00796275f $X=0.975 $Y=0.495 $X2=0
+ $Y2=0
cc_160 N_A_108_31#_c_84_n N_VGND_c_414_n 0.00116576f $X=1.355 $Y=0.95 $X2=0
+ $Y2=0
cc_161 N_A_108_31#_c_85_n N_VGND_c_414_n 0.0124703f $X=1.98 $Y=0.495 $X2=0 $Y2=0
cc_162 N_A_108_31#_c_87_n N_VGND_c_414_n 0.0125808f $X=3.56 $Y=0.495 $X2=0 $Y2=0
cc_163 N_A_c_187_n N_B_c_249_n 0.00899044f $X=1.765 $Y=0.78 $X2=-0.19 $Y2=-0.245
cc_164 N_A_c_189_n N_B_c_251_n 0.00899044f $X=1.765 $Y=0.855 $X2=0 $Y2=0
cc_165 N_A_c_191_n N_B_c_251_n 9.4238e-19 $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_166 N_A_c_188_n N_B_M1000_g 0.0696247f $X=1.902 $Y=1.673 $X2=0 $Y2=0
cc_167 N_A_c_192_n N_B_c_254_n 0.0057515f $X=1.902 $Y=1.215 $X2=0 $Y2=0
cc_168 N_A_c_188_n N_B_c_255_n 0.0110544f $X=1.902 $Y=1.673 $X2=0 $Y2=0
cc_169 N_A_c_190_n N_B_c_256_n 0.0110544f $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_170 N_A_c_191_n N_B_c_256_n 0.0115969f $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_171 N_A_c_188_n N_B_c_257_n 0.0011414f $X=1.902 $Y=1.673 $X2=0 $Y2=0
cc_172 N_A_c_190_n N_B_c_257_n 6.61375e-19 $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_173 N_A_c_191_n N_B_c_257_n 0.133576f $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_174 N_A_c_191_n N_VPWR_M1005_d 0.0234767f $X=1.855 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_c_194_n N_VPWR_c_378_n 0.00904307f $X=2.09 $Y=2.01 $X2=0 $Y2=0
cc_176 N_A_c_191_n N_VPWR_c_378_n 0.0678142f $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_177 N_A_c_194_n N_VPWR_c_380_n 0.00595064f $X=2.09 $Y=2.01 $X2=0 $Y2=0
cc_178 N_A_c_191_n N_VPWR_c_380_n 0.0202921f $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_179 N_A_c_194_n N_VPWR_c_377_n 0.00855176f $X=2.09 $Y=2.01 $X2=0 $Y2=0
cc_180 N_A_c_191_n N_VPWR_c_377_n 0.0234256f $X=1.855 $Y=1.38 $X2=0 $Y2=0
cc_181 N_A_c_191_n A_443_409# 0.00757755f $X=1.855 $Y=1.38 $X2=-0.19 $Y2=-0.245
cc_182 N_A_c_184_n N_VGND_c_409_n 0.0114545f $X=1.405 $Y=0.78 $X2=0 $Y2=0
cc_183 N_A_c_187_n N_VGND_c_409_n 0.00200313f $X=1.765 $Y=0.78 $X2=0 $Y2=0
cc_184 N_A_c_184_n N_VGND_c_412_n 0.00445056f $X=1.405 $Y=0.78 $X2=0 $Y2=0
cc_185 N_A_c_185_n N_VGND_c_412_n 4.57848e-19 $X=1.69 $Y=0.855 $X2=0 $Y2=0
cc_186 N_A_c_187_n N_VGND_c_412_n 0.00502664f $X=1.765 $Y=0.78 $X2=0 $Y2=0
cc_187 N_A_c_184_n N_VGND_c_414_n 0.00796275f $X=1.405 $Y=0.78 $X2=0 $Y2=0
cc_188 N_A_c_185_n N_VGND_c_414_n 6.33118e-19 $X=1.69 $Y=0.855 $X2=0 $Y2=0
cc_189 N_A_c_187_n N_VGND_c_414_n 0.00942073f $X=1.765 $Y=0.78 $X2=0 $Y2=0
cc_190 N_B_c_252_n N_C_c_309_n 0.00973888f $X=2.555 $Y=0.78 $X2=-0.19 $Y2=-0.245
cc_191 N_B_M1000_g N_C_M1006_g 0.0484879f $X=2.58 $Y=2.545 $X2=0 $Y2=0
cc_192 N_B_c_257_n N_C_M1006_g 0.0115796f $X=2.62 $Y=1.38 $X2=0 $Y2=0
cc_193 N_B_c_253_n N_C_c_311_n 0.00973888f $X=2.542 $Y=0.855 $X2=0 $Y2=0
cc_194 N_B_c_254_n N_C_c_312_n 0.00897589f $X=2.62 $Y=1.215 $X2=0 $Y2=0
cc_195 N_B_c_255_n N_C_c_313_n 0.01184f $X=2.62 $Y=1.72 $X2=0 $Y2=0
cc_196 N_B_c_260_n N_C_c_318_n 0.01184f $X=2.62 $Y=1.885 $X2=0 $Y2=0
cc_197 N_B_c_256_n N_C_c_314_n 0.01184f $X=2.62 $Y=1.38 $X2=0 $Y2=0
cc_198 N_B_c_257_n N_C_c_314_n 8.23261e-19 $X=2.62 $Y=1.38 $X2=0 $Y2=0
cc_199 N_B_c_256_n N_C_c_315_n 0.00410205f $X=2.62 $Y=1.38 $X2=0 $Y2=0
cc_200 N_B_c_257_n N_C_c_315_n 0.0438819f $X=2.62 $Y=1.38 $X2=0 $Y2=0
cc_201 N_B_M1000_g N_VPWR_c_380_n 0.00596257f $X=2.58 $Y=2.545 $X2=0 $Y2=0
cc_202 N_B_c_257_n N_VPWR_c_380_n 0.00914393f $X=2.62 $Y=1.38 $X2=0 $Y2=0
cc_203 N_B_M1000_g N_VPWR_c_377_n 0.00771107f $X=2.58 $Y=2.545 $X2=0 $Y2=0
cc_204 N_B_c_257_n N_VPWR_c_377_n 0.0101955f $X=2.62 $Y=1.38 $X2=0 $Y2=0
cc_205 N_B_c_257_n A_541_409# 0.0116447f $X=2.62 $Y=1.38 $X2=-0.19 $Y2=-0.245
cc_206 N_B_c_249_n N_VGND_c_410_n 0.00200313f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_207 N_B_c_252_n N_VGND_c_410_n 0.0114581f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_208 N_B_c_249_n N_VGND_c_412_n 0.00502664f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_209 N_B_c_250_n N_VGND_c_412_n 4.57848e-19 $X=2.455 $Y=0.855 $X2=0 $Y2=0
cc_210 N_B_c_252_n N_VGND_c_412_n 0.00445056f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_211 N_B_c_249_n N_VGND_c_414_n 0.00942073f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_212 N_B_c_250_n N_VGND_c_414_n 6.33118e-19 $X=2.455 $Y=0.855 $X2=0 $Y2=0
cc_213 N_B_c_252_n N_VGND_c_414_n 0.00796275f $X=2.555 $Y=0.78 $X2=0 $Y2=0
cc_214 N_C_M1006_g N_VPWR_c_380_n 0.0086001f $X=3.15 $Y=2.545 $X2=0 $Y2=0
cc_215 N_C_M1006_g N_VPWR_c_377_n 0.0165732f $X=3.15 $Y=2.545 $X2=0 $Y2=0
cc_216 N_C_c_309_n N_VGND_c_410_n 0.0114736f $X=2.985 $Y=0.78 $X2=0 $Y2=0
cc_217 N_C_c_310_n N_VGND_c_410_n 0.00200313f $X=3.345 $Y=0.78 $X2=0 $Y2=0
cc_218 N_C_c_309_n N_VGND_c_413_n 0.00445056f $X=2.985 $Y=0.78 $X2=0 $Y2=0
cc_219 N_C_c_310_n N_VGND_c_413_n 0.00502664f $X=3.345 $Y=0.78 $X2=0 $Y2=0
cc_220 N_C_c_311_n N_VGND_c_413_n 5.63805e-19 $X=3.345 $Y=0.855 $X2=0 $Y2=0
cc_221 N_C_c_309_n N_VGND_c_414_n 0.00796275f $X=2.985 $Y=0.78 $X2=0 $Y2=0
cc_222 N_C_c_310_n N_VGND_c_414_n 0.0100616f $X=3.345 $Y=0.78 $X2=0 $Y2=0
cc_223 N_C_c_311_n N_VGND_c_414_n 7.67806e-19 $X=3.345 $Y=0.855 $X2=0 $Y2=0
cc_224 X N_VPWR_c_378_n 0.0728647f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_225 X N_VPWR_c_379_n 0.0483277f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_226 X N_VPWR_c_377_n 0.0276711f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_227 N_X_c_357_n A_138_57# 0.00133334f $X=0.485 $Y=0.8 $X2=-0.19 $Y2=-0.245
cc_228 N_X_c_357_n N_VGND_c_409_n 0.00600007f $X=0.485 $Y=0.8 $X2=0 $Y2=0
cc_229 N_X_c_357_n N_VGND_c_411_n 0.0373716f $X=0.485 $Y=0.8 $X2=0 $Y2=0
cc_230 N_X_c_357_n N_VGND_c_414_n 0.0260354f $X=0.485 $Y=0.8 $X2=0 $Y2=0
