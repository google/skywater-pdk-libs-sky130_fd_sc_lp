* File: sky130_fd_sc_lp__a211o_m.pxi.spice
* Created: Wed Sep  2 09:17:51 2020
* 
x_PM_SKY130_FD_SC_LP__A211O_M%A2 N_A2_M1002_g N_A2_M1001_g A2 N_A2_c_65_n
+ N_A2_c_66_n PM_SKY130_FD_SC_LP__A211O_M%A2
x_PM_SKY130_FD_SC_LP__A211O_M%A1 N_A1_c_90_n N_A1_M1009_g N_A1_M1008_g
+ N_A1_c_92_n A1 A1 N_A1_c_94_n PM_SKY130_FD_SC_LP__A211O_M%A1
x_PM_SKY130_FD_SC_LP__A211O_M%A_82_483# N_A_82_483#_M1009_d N_A_82_483#_M1004_d
+ N_A_82_483#_M1005_d N_A_82_483#_c_134_n N_A_82_483#_M1006_g
+ N_A_82_483#_M1007_g N_A_82_483#_c_136_n N_A_82_483#_c_137_n
+ N_A_82_483#_c_138_n N_A_82_483#_c_139_n N_A_82_483#_c_140_n
+ N_A_82_483#_c_141_n N_A_82_483#_c_130_n N_A_82_483#_c_143_n
+ N_A_82_483#_c_131_n N_A_82_483#_c_132_n N_A_82_483#_c_144_n
+ N_A_82_483#_c_133_n N_A_82_483#_c_162_p N_A_82_483#_c_145_n
+ PM_SKY130_FD_SC_LP__A211O_M%A_82_483#
x_PM_SKY130_FD_SC_LP__A211O_M%B1 N_B1_M1000_g N_B1_M1003_g B1 B1 N_B1_c_216_n
+ N_B1_c_217_n PM_SKY130_FD_SC_LP__A211O_M%B1
x_PM_SKY130_FD_SC_LP__A211O_M%C1 N_C1_M1005_g N_C1_M1004_g C1 N_C1_c_253_n
+ PM_SKY130_FD_SC_LP__A211O_M%C1
x_PM_SKY130_FD_SC_LP__A211O_M%X N_X_M1007_s N_X_M1006_s X X X X X X X
+ PM_SKY130_FD_SC_LP__A211O_M%X
x_PM_SKY130_FD_SC_LP__A211O_M%VPWR N_VPWR_M1006_d N_VPWR_M1002_d N_VPWR_c_287_n
+ N_VPWR_c_288_n VPWR N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_291_n
+ N_VPWR_c_286_n N_VPWR_c_293_n N_VPWR_c_294_n PM_SKY130_FD_SC_LP__A211O_M%VPWR
x_PM_SKY130_FD_SC_LP__A211O_M%A_225_389# N_A_225_389#_M1002_s
+ N_A_225_389#_M1008_d N_A_225_389#_c_320_n N_A_225_389#_c_321_n
+ N_A_225_389#_c_322_n N_A_225_389#_c_330_n
+ PM_SKY130_FD_SC_LP__A211O_M%A_225_389#
x_PM_SKY130_FD_SC_LP__A211O_M%VGND N_VGND_M1007_d N_VGND_M1000_d N_VGND_c_342_n
+ N_VGND_c_343_n N_VGND_c_344_n N_VGND_c_358_n N_VGND_c_364_n VGND
+ N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n N_VGND_c_349_n
+ PM_SKY130_FD_SC_LP__A211O_M%VGND
cc_1 VNB N_A2_M1002_g 0.00567005f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=2.155
cc_2 VNB A2 0.0136334f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_3 VNB N_A2_c_65_n 0.0384743f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.42
cc_4 VNB N_A2_c_66_n 0.0172004f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.255
cc_5 VNB N_A1_c_90_n 0.0570366f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.585
cc_6 VNB N_A1_M1009_g 0.0442801f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=1.255
cc_7 VNB N_A1_c_92_n 0.00258887f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.255
cc_8 VNB A1 0.0050897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_c_94_n 0.0498264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_82_483#_M1007_g 0.0508975f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.397
cc_11 VNB N_A_82_483#_c_130_n 0.00261227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_82_483#_c_131_n 0.01461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_82_483#_c_132_n 0.00641614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_82_483#_c_133_n 8.72418e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1000_g 0.0312519f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=2.155
cc_16 VNB B1 0.00567693f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_17 VNB N_B1_c_216_n 0.0367242f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.42
cc_18 VNB N_B1_c_217_n 0.00856828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C1_M1004_g 0.0367181f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=0.935
cc_20 VNB C1 0.00700403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C1_c_253_n 0.0292896f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.397
cc_22 VNB X 0.0584269f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=0.935
cc_23 VNB N_VPWR_c_286_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_342_n 0.0195348f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_25 VNB N_VGND_c_343_n 0.0485431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_344_n 0.021601f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.42
cc_27 VNB N_VGND_c_345_n 0.018844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_346_n 0.0204409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_347_n 0.217343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_348_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_349_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_A2_M1002_g 0.0298815f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=2.155
cc_33 VPB N_A1_M1009_g 0.0225482f $X=-0.19 $Y=1.655 $X2=1.535 $Y2=1.255
cc_34 VPB N_A_82_483#_c_134_n 0.0221634f $X=-0.19 $Y=1.655 $X2=1.43 $Y2=1.42
cc_35 VPB N_A_82_483#_M1007_g 0.0552108f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.397
cc_36 VPB N_A_82_483#_c_136_n 0.0382965f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.397
cc_37 VPB N_A_82_483#_c_137_n 0.010626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_82_483#_c_138_n 0.0628418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_82_483#_c_139_n 0.00961157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_82_483#_c_140_n 0.00856122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_82_483#_c_141_n 0.0177625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_82_483#_c_130_n 0.00219637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_82_483#_c_143_n 0.0132497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_82_483#_c_144_n 0.00271508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_82_483#_c_145_n 0.0444191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B1_M1000_g 0.0226442f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=2.155
cc_47 VPB N_C1_M1005_g 0.0287856f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=2.155
cc_48 VPB C1 0.00770225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_C1_c_253_n 0.0238635f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.397
cc_50 VPB X 0.054868f $X=-0.19 $Y=1.655 $X2=1.535 $Y2=0.935
cc_51 VPB N_VPWR_c_287_n 0.00495479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_288_n 0.0224774f $X=-0.19 $Y=1.655 $X2=1.43 $Y2=1.255
cc_53 VPB N_VPWR_c_289_n 0.0192393f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.397
cc_54 VPB N_VPWR_c_290_n 0.0224788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_291_n 0.0453748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_286_n 0.0928832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_293_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_294_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_225_389#_c_320_n 2.17323e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_225_389#_c_321_n 0.0151373f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.42
cc_61 VPB N_A_225_389#_c_322_n 0.00805936f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.42
cc_62 N_A2_c_66_n N_A1_c_90_n 0.00838916f $X=1.43 $Y=1.255 $X2=-0.19 $Y2=-0.245
cc_63 N_A2_M1002_g N_A1_M1009_g 0.0264083f $X=1.465 $Y=2.155 $X2=0 $Y2=0
cc_64 A2 N_A1_M1009_g 0.00427231f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A2_c_66_n N_A1_M1009_g 0.0599631f $X=1.43 $Y=1.255 $X2=0 $Y2=0
cc_66 N_A2_c_65_n A1 0.00135614f $X=1.415 $Y=1.42 $X2=0 $Y2=0
cc_67 N_A2_c_66_n A1 0.0125602f $X=1.43 $Y=1.255 $X2=0 $Y2=0
cc_68 N_A2_c_65_n N_A_82_483#_M1007_g 0.00818352f $X=1.415 $Y=1.42 $X2=0 $Y2=0
cc_69 N_A2_M1002_g N_A_82_483#_c_136_n 0.00330624f $X=1.465 $Y=2.155 $X2=0 $Y2=0
cc_70 N_A2_M1002_g N_A_82_483#_c_138_n 0.00949186f $X=1.465 $Y=2.155 $X2=0 $Y2=0
cc_71 A2 N_A_82_483#_c_130_n 0.0071005f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_72 A2 N_A_82_483#_c_132_n 0.0102211f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A2_c_66_n N_A_82_483#_c_132_n 0.00138946f $X=1.43 $Y=1.255 $X2=0 $Y2=0
cc_74 A2 N_B1_c_217_n 0.00610667f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A2_c_66_n N_B1_c_217_n 0.00157983f $X=1.43 $Y=1.255 $X2=0 $Y2=0
cc_76 N_A2_M1002_g N_VPWR_c_288_n 0.0121052f $X=1.465 $Y=2.155 $X2=0 $Y2=0
cc_77 N_A2_M1002_g N_A_225_389#_c_320_n 3.52891e-19 $X=1.465 $Y=2.155 $X2=0
+ $Y2=0
cc_78 N_A2_M1002_g N_A_225_389#_c_321_n 0.0153304f $X=1.465 $Y=2.155 $X2=0 $Y2=0
cc_79 A2 N_A_225_389#_c_321_n 0.0313141f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A2_c_65_n N_A_225_389#_c_321_n 0.00305514f $X=1.415 $Y=1.42 $X2=0 $Y2=0
cc_81 A2 N_A_225_389#_c_322_n 3.98847e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A2_c_65_n N_A_225_389#_c_322_n 0.00347104f $X=1.415 $Y=1.42 $X2=0 $Y2=0
cc_83 N_A2_c_66_n N_VGND_c_347_n 7.80882e-19 $X=1.43 $Y=1.255 $X2=0 $Y2=0
cc_84 A1 N_A_82_483#_M1007_g 6.97002e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A1_M1009_g N_A_82_483#_c_138_n 0.00955511f $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_86 N_A1_M1009_g N_A_82_483#_c_130_n 0.00171366f $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_87 N_A1_M1009_g N_A_82_483#_c_143_n 6.2062e-19 $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_88 N_A1_M1009_g N_A_82_483#_c_132_n 0.00988514f $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_89 A1 N_A_82_483#_c_132_n 0.00238324f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A1_M1009_g N_B1_M1000_g 0.0533376f $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_91 N_A1_c_90_n N_B1_c_216_n 0.021337f $X=1.82 $Y=0.26 $X2=0 $Y2=0
cc_92 N_A1_c_90_n N_B1_c_217_n 0.0114925f $X=1.82 $Y=0.26 $X2=0 $Y2=0
cc_93 N_A1_M1009_g N_B1_c_217_n 0.0179782f $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_94 N_A1_c_92_n N_B1_c_217_n 0.00925355f $X=1.2 $Y=0.35 $X2=0 $Y2=0
cc_95 A1 N_B1_c_217_n 0.011122f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_96 N_A1_c_94_n N_B1_c_217_n 8.52245e-19 $X=1.085 $Y=0.26 $X2=0 $Y2=0
cc_97 N_A1_M1009_g N_VPWR_c_288_n 0.00782349f $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_98 N_A1_M1009_g N_A_225_389#_c_321_n 0.017636f $X=1.895 $Y=0.935 $X2=0 $Y2=0
cc_99 N_A1_M1009_g N_A_225_389#_c_330_n 2.03427e-19 $X=1.895 $Y=0.935 $X2=0
+ $Y2=0
cc_100 A1 N_VGND_M1007_d 0.0159441f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_101 N_A1_c_92_n N_VGND_c_342_n 0.012244f $X=1.2 $Y=0.35 $X2=0 $Y2=0
cc_102 A1 N_VGND_c_342_n 0.0139502f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_103 N_A1_c_94_n N_VGND_c_342_n 0.00577906f $X=1.085 $Y=0.26 $X2=0 $Y2=0
cc_104 N_A1_c_92_n N_VGND_c_343_n 0.0210617f $X=1.2 $Y=0.35 $X2=0 $Y2=0
cc_105 N_A1_c_94_n N_VGND_c_343_n 0.0233615f $X=1.085 $Y=0.26 $X2=0 $Y2=0
cc_106 N_A1_c_90_n N_VGND_c_344_n 0.00128822f $X=1.82 $Y=0.26 $X2=0 $Y2=0
cc_107 A1 N_VGND_c_358_n 0.0134137f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A1_c_90_n N_VGND_c_347_n 0.0252807f $X=1.82 $Y=0.26 $X2=0 $Y2=0
cc_109 N_A1_c_92_n N_VGND_c_347_n 0.0119374f $X=1.2 $Y=0.35 $X2=0 $Y2=0
cc_110 N_A1_c_94_n N_VGND_c_347_n 0.00896182f $X=1.085 $Y=0.26 $X2=0 $Y2=0
cc_111 N_A_82_483#_c_141_n N_B1_M1000_g 0.00510879f $X=2.395 $Y=2.9 $X2=0 $Y2=0
cc_112 N_A_82_483#_c_130_n N_B1_M1000_g 0.0126624f $X=2.48 $Y=1.93 $X2=0 $Y2=0
cc_113 N_A_82_483#_c_143_n N_B1_M1000_g 0.00526395f $X=2.48 $Y=2.735 $X2=0 $Y2=0
cc_114 N_A_82_483#_c_132_n N_B1_M1000_g 0.0216333f $X=2.565 $Y=1.25 $X2=0 $Y2=0
cc_115 N_A_82_483#_c_162_p N_B1_M1000_g 0.0058533f $X=2.48 $Y=2.095 $X2=0 $Y2=0
cc_116 N_A_82_483#_c_145_n N_B1_M1000_g 0.00155068f $X=2.11 $Y=2.81 $X2=0 $Y2=0
cc_117 N_A_82_483#_c_132_n B1 0.0152748f $X=2.565 $Y=1.25 $X2=0 $Y2=0
cc_118 N_A_82_483#_c_132_n N_B1_c_216_n 0.0012626f $X=2.565 $Y=1.25 $X2=0 $Y2=0
cc_119 N_A_82_483#_c_132_n N_B1_c_217_n 0.00485002f $X=2.565 $Y=1.25 $X2=0 $Y2=0
cc_120 N_A_82_483#_c_143_n N_C1_M1005_g 0.00334436f $X=2.48 $Y=2.735 $X2=0 $Y2=0
cc_121 N_A_82_483#_c_144_n N_C1_M1005_g 0.0176969f $X=2.9 $Y=2.095 $X2=0 $Y2=0
cc_122 N_A_82_483#_c_130_n N_C1_M1004_g 0.00248117f $X=2.48 $Y=1.93 $X2=0 $Y2=0
cc_123 N_A_82_483#_c_131_n N_C1_M1004_g 0.0158459f $X=2.965 $Y=1.25 $X2=0 $Y2=0
cc_124 N_A_82_483#_c_132_n N_C1_M1004_g 6.373e-19 $X=2.565 $Y=1.25 $X2=0 $Y2=0
cc_125 N_A_82_483#_c_133_n N_C1_M1004_g 7.46117e-19 $X=3.05 $Y=1 $X2=0 $Y2=0
cc_126 N_A_82_483#_c_130_n C1 0.0148336f $X=2.48 $Y=1.93 $X2=0 $Y2=0
cc_127 N_A_82_483#_c_131_n C1 0.0262884f $X=2.965 $Y=1.25 $X2=0 $Y2=0
cc_128 N_A_82_483#_c_144_n C1 0.018015f $X=2.9 $Y=2.095 $X2=0 $Y2=0
cc_129 N_A_82_483#_c_130_n N_C1_c_253_n 0.00777645f $X=2.48 $Y=1.93 $X2=0 $Y2=0
cc_130 N_A_82_483#_c_131_n N_C1_c_253_n 0.00934625f $X=2.965 $Y=1.25 $X2=0 $Y2=0
cc_131 N_A_82_483#_c_144_n N_C1_c_253_n 0.00639258f $X=2.9 $Y=2.095 $X2=0 $Y2=0
cc_132 N_A_82_483#_M1007_g X 0.0556139f $X=0.52 $Y=0.935 $X2=0 $Y2=0
cc_133 N_A_82_483#_c_140_n X 0.0120296f $X=0.502 $Y=2.49 $X2=0 $Y2=0
cc_134 N_A_82_483#_c_134_n N_VPWR_c_287_n 0.00460896f $X=0.485 $Y=2.565 $X2=0
+ $Y2=0
cc_135 N_A_82_483#_c_136_n N_VPWR_c_287_n 0.0058931f $X=0.9 $Y=2.49 $X2=0 $Y2=0
cc_136 N_A_82_483#_c_139_n N_VPWR_c_287_n 0.00263239f $X=1.05 $Y=2.81 $X2=0
+ $Y2=0
cc_137 N_A_82_483#_c_136_n N_VPWR_c_288_n 0.00729552f $X=0.9 $Y=2.49 $X2=0 $Y2=0
cc_138 N_A_82_483#_c_138_n N_VPWR_c_288_n 0.0281647f $X=1.945 $Y=2.81 $X2=0
+ $Y2=0
cc_139 N_A_82_483#_c_141_n N_VPWR_c_288_n 0.0252851f $X=2.395 $Y=2.9 $X2=0 $Y2=0
cc_140 N_A_82_483#_c_143_n N_VPWR_c_288_n 0.0147986f $X=2.48 $Y=2.735 $X2=0
+ $Y2=0
cc_141 N_A_82_483#_c_145_n N_VPWR_c_288_n 0.0045032f $X=2.11 $Y=2.81 $X2=0 $Y2=0
cc_142 N_A_82_483#_c_134_n N_VPWR_c_289_n 0.00585385f $X=0.485 $Y=2.565 $X2=0
+ $Y2=0
cc_143 N_A_82_483#_c_139_n N_VPWR_c_290_n 0.0150888f $X=1.05 $Y=2.81 $X2=0 $Y2=0
cc_144 N_A_82_483#_c_138_n N_VPWR_c_291_n 0.0023335f $X=1.945 $Y=2.81 $X2=0
+ $Y2=0
cc_145 N_A_82_483#_c_141_n N_VPWR_c_291_n 0.0341188f $X=2.395 $Y=2.9 $X2=0 $Y2=0
cc_146 N_A_82_483#_c_145_n N_VPWR_c_291_n 0.0081186f $X=2.11 $Y=2.81 $X2=0 $Y2=0
cc_147 N_A_82_483#_c_134_n N_VPWR_c_286_n 0.0130126f $X=0.485 $Y=2.565 $X2=0
+ $Y2=0
cc_148 N_A_82_483#_c_139_n N_VPWR_c_286_n 0.0190562f $X=1.05 $Y=2.81 $X2=0 $Y2=0
cc_149 N_A_82_483#_c_141_n N_VPWR_c_286_n 0.0204578f $X=2.395 $Y=2.9 $X2=0 $Y2=0
cc_150 N_A_82_483#_c_145_n N_VPWR_c_286_n 0.0104909f $X=2.11 $Y=2.81 $X2=0 $Y2=0
cc_151 N_A_82_483#_M1007_g N_A_225_389#_c_320_n 0.00745488f $X=0.52 $Y=0.935
+ $X2=0 $Y2=0
cc_152 N_A_82_483#_c_138_n N_A_225_389#_c_320_n 0.00528775f $X=1.945 $Y=2.81
+ $X2=0 $Y2=0
cc_153 N_A_82_483#_c_130_n N_A_225_389#_c_321_n 0.0127186f $X=2.48 $Y=1.93 $X2=0
+ $Y2=0
cc_154 N_A_82_483#_c_132_n N_A_225_389#_c_321_n 0.0119699f $X=2.565 $Y=1.25
+ $X2=0 $Y2=0
cc_155 N_A_82_483#_c_162_p N_A_225_389#_c_321_n 4.24085e-19 $X=2.48 $Y=2.095
+ $X2=0 $Y2=0
cc_156 N_A_82_483#_M1007_g N_A_225_389#_c_322_n 0.00470066f $X=0.52 $Y=0.935
+ $X2=0 $Y2=0
cc_157 N_A_82_483#_c_141_n N_A_225_389#_c_330_n 0.00632222f $X=2.395 $Y=2.9
+ $X2=0 $Y2=0
cc_158 N_A_82_483#_c_162_p N_A_225_389#_c_330_n 0.0129564f $X=2.48 $Y=2.095
+ $X2=0 $Y2=0
cc_159 N_A_82_483#_c_145_n N_A_225_389#_c_330_n 0.00341808f $X=2.11 $Y=2.81
+ $X2=0 $Y2=0
cc_160 N_A_82_483#_M1007_g N_VGND_c_342_n 0.00473171f $X=0.52 $Y=0.935 $X2=0
+ $Y2=0
cc_161 N_A_82_483#_M1007_g N_VGND_c_358_n 0.00339328f $X=0.52 $Y=0.935 $X2=0
+ $Y2=0
cc_162 N_A_82_483#_c_131_n N_VGND_c_364_n 0.013552f $X=2.965 $Y=1.25 $X2=0 $Y2=0
cc_163 N_A_82_483#_c_132_n N_VGND_c_364_n 0.00882399f $X=2.565 $Y=1.25 $X2=0
+ $Y2=0
cc_164 N_A_82_483#_M1007_g N_VGND_c_345_n 0.0030451f $X=0.52 $Y=0.935 $X2=0
+ $Y2=0
cc_165 N_A_82_483#_M1007_g N_VGND_c_347_n 0.00371829f $X=0.52 $Y=0.935 $X2=0
+ $Y2=0
cc_166 N_A_82_483#_c_133_n N_VGND_c_347_n 0.00720315f $X=3.05 $Y=1 $X2=0 $Y2=0
cc_167 N_B1_M1000_g N_C1_M1004_g 0.0200447f $X=2.325 $Y=0.935 $X2=0 $Y2=0
cc_168 N_B1_M1000_g N_C1_c_253_n 0.0641478f $X=2.325 $Y=0.935 $X2=0 $Y2=0
cc_169 N_B1_M1000_g N_VPWR_c_288_n 6.89369e-19 $X=2.325 $Y=0.935 $X2=0 $Y2=0
cc_170 N_B1_M1000_g N_A_225_389#_c_321_n 0.00146899f $X=2.325 $Y=0.935 $X2=0
+ $Y2=0
cc_171 B1 N_VGND_c_343_n 0.0231034f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_172 N_B1_c_216_n N_VGND_c_343_n 0.004277f $X=2.345 $Y=0.43 $X2=0 $Y2=0
cc_173 N_B1_c_217_n N_VGND_c_343_n 0.0284309f $X=2.058 $Y=0.452 $X2=0 $Y2=0
cc_174 N_B1_M1000_g N_VGND_c_344_n 0.00309591f $X=2.325 $Y=0.935 $X2=0 $Y2=0
cc_175 B1 N_VGND_c_344_n 0.0269264f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_176 N_B1_c_216_n N_VGND_c_344_n 0.00805121f $X=2.345 $Y=0.43 $X2=0 $Y2=0
cc_177 N_B1_c_216_n N_VGND_c_364_n 0.00205504f $X=2.345 $Y=0.43 $X2=0 $Y2=0
cc_178 B1 N_VGND_c_347_n 0.0139986f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_179 N_B1_c_216_n N_VGND_c_347_n 0.00254324f $X=2.345 $Y=0.43 $X2=0 $Y2=0
cc_180 N_B1_c_217_n N_VGND_c_347_n 0.015864f $X=2.058 $Y=0.452 $X2=0 $Y2=0
cc_181 N_C1_M1005_g N_VPWR_c_286_n 0.00384901f $X=2.685 $Y=2.155 $X2=0 $Y2=0
cc_182 N_C1_M1004_g N_VGND_c_344_n 0.00906248f $X=2.835 $Y=0.935 $X2=0 $Y2=0
cc_183 N_C1_M1004_g N_VGND_c_364_n 0.00459536f $X=2.835 $Y=0.935 $X2=0 $Y2=0
cc_184 N_C1_M1004_g N_VGND_c_346_n 0.0030451f $X=2.835 $Y=0.935 $X2=0 $Y2=0
cc_185 N_C1_M1004_g N_VGND_c_347_n 0.00371829f $X=2.835 $Y=0.935 $X2=0 $Y2=0
cc_186 X N_VPWR_c_289_n 0.0095728f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_187 N_X_M1006_s N_VPWR_c_286_n 0.00334315f $X=0.145 $Y=2.675 $X2=0 $Y2=0
cc_188 X N_VPWR_c_286_n 0.00863123f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_189 X N_VGND_c_342_n 0.0196684f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_190 X N_VGND_c_345_n 0.00698589f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_191 X N_VGND_c_347_n 0.00795962f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_192 N_VPWR_c_288_n N_A_225_389#_c_321_n 0.0207154f $X=1.68 $Y=2.22 $X2=0
+ $Y2=0
