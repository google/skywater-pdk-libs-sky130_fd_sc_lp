* File: sky130_fd_sc_lp__edfxbp_1.pex.spice
* Created: Wed Sep  2 09:51:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%DE 3 7 9 15 17 19 20 22 24 25 26 32 34 44
c61 32 0 6.76474e-20 $X=1.25 $Y=2.9
c62 15 0 2.85507e-19 $X=1.515 $Y=0.475
r63 44 45 2.57123 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=1.25 $Y=2.775 $X2=1.25
+ $Y2=2.735
r64 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=2.9
+ $X2=1.25 $Y2=2.735
r65 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=2.9 $X2=1.25 $Y2=2.9
r66 26 33 3.59702 $w=3.28e-07 $l=1.03e-07 $layer=LI1_cond $X=1.25 $Y=2.797
+ $X2=1.25 $Y2=2.9
r67 26 44 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=1.25 $Y=2.797
+ $X2=1.25 $Y2=2.775
r68 26 45 1.17805 $w=2.23e-07 $l=2.3e-08 $layer=LI1_cond $X=1.197 $Y=2.712
+ $X2=1.197 $Y2=2.735
r69 25 26 15.7244 $w=2.23e-07 $l=3.07e-07 $layer=LI1_cond $X=1.197 $Y=2.405
+ $X2=1.197 $Y2=2.712
r70 24 25 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.197 $Y=2.035
+ $X2=1.197 $Y2=2.405
r71 22 23 61.9393 $w=2.14e-07 $l=2.75e-07 $layer=POLY_cond $X=1.515 $Y=1.88
+ $X2=1.79 $Y2=1.88
r72 21 22 79.9579 $w=2.14e-07 $l=3.55e-07 $layer=POLY_cond $X=1.16 $Y=1.88
+ $X2=1.515 $Y2=1.88
r73 17 23 11.1354 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.79 $Y=2.005
+ $X2=1.79 $Y2=1.88
r74 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.79 $Y=2.005
+ $X2=1.79 $Y2=2.325
r75 13 22 11.1354 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.515 $Y=1.755
+ $X2=1.515 $Y2=1.88
r76 13 15 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=1.515 $Y=1.755
+ $X2=1.515 $Y2=0.475
r77 11 21 11.1354 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.16 $Y=2.005
+ $X2=1.16 $Y2=1.88
r78 11 34 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.16 $Y=2.005
+ $X2=1.16 $Y2=2.735
r79 10 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.6 $Y=1.83
+ $X2=0.525 $Y2=1.83
r80 9 21 21.2592 $w=2.14e-07 $l=9.68246e-08 $layer=POLY_cond $X=1.085 $Y=1.83
+ $X2=1.16 $Y2=1.88
r81 9 10 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.085 $Y=1.83
+ $X2=0.6 $Y2=1.83
r82 5 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.525 $Y=1.905
+ $X2=0.525 $Y2=1.83
r83 5 7 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.525 $Y=1.905
+ $X2=0.525 $Y2=2.725
r84 1 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.525 $Y=1.755
+ $X2=0.525 $Y2=1.83
r85 1 3 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.525 $Y=1.755
+ $X2=0.525 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_120_179# 1 2 9 13 17 21 25 26 28
c63 21 0 1.3912e-19 $X=0.74 $Y=2.55
c64 13 0 1.35708e-19 $X=2.22 $Y=2.325
r65 26 29 15.0104 $w=2.89e-07 $l=9e-08 $layer=POLY_cond $X=2.035 $Y=1.4
+ $X2=1.945 $Y2=1.4
r66 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.035
+ $Y=1.4 $X2=2.035 $Y2=1.4
r67 23 28 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.4
+ $X2=0.74 $Y2=1.4
r68 23 25 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.905 $Y=1.4
+ $X2=2.035 $Y2=1.4
r69 19 28 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.74 $Y=1.565
+ $X2=0.74 $Y2=1.4
r70 19 21 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=0.74 $Y=1.565
+ $X2=0.74 $Y2=2.55
r71 15 28 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.74 $Y=1.235
+ $X2=0.74 $Y2=1.4
r72 15 17 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.74 $Y=1.235
+ $X2=0.74 $Y2=1.105
r73 11 26 30.8547 $w=2.89e-07 $l=2.5446e-07 $layer=POLY_cond $X=2.22 $Y=1.565
+ $X2=2.035 $Y2=1.4
r74 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.22 $Y=1.565
+ $X2=2.22 $Y2=2.325
r75 7 29 18.0918 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=1.235
+ $X2=1.945 $Y2=1.4
r76 7 9 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.945 $Y=1.235
+ $X2=1.945 $Y2=0.475
r77 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=2.405 $X2=0.74 $Y2=2.55
r78 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.895 $X2=0.74 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%D 3 7 9 13
r41 11 13 16.2472 $w=2.67e-07 $l=9e-08 $layer=POLY_cond $X=2.58 $Y=1.345
+ $X2=2.67 $Y2=1.345
r42 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.345 $X2=2.67 $Y2=1.345
r43 5 13 47.839 $w=2.67e-07 $l=3.37565e-07 $layer=POLY_cond $X=2.935 $Y=1.18
+ $X2=2.67 $Y2=1.345
r44 5 7 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.935 $Y=1.18
+ $X2=2.935 $Y2=0.77
r45 1 11 16.2448 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.51
+ $X2=2.58 $Y2=1.345
r46 1 3 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.58 $Y=1.51 $X2=2.58
+ $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_587_350# 1 2 9 11 12 15 19 23 25 26 29 33
+ 40 44 45 49 50 53 54 57 60 67 81
c206 67 0 1.11531e-19 $X=11.73 $Y=1.67
c207 60 0 1.75981e-19 $X=12.24 $Y=2.035
c208 53 0 1.52339e-20 $X=12.095 $Y=2.035
c209 49 0 1.61716e-19 $X=3.655 $Y=1.615
r210 71 81 4.84477 $w=5.54e-07 $l=3.16425e-07 $layer=LI1_cond $X=11.96 $Y=1.76
+ $X2=12.185 $Y2=1.98
r211 71 78 5.94585 $w=5.54e-07 $l=2.7e-07 $layer=LI1_cond $X=11.96 $Y=1.76
+ $X2=11.96 $Y2=1.49
r212 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.73
+ $Y=1.76 $X2=11.73 $Y2=1.76
r213 67 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.73 $Y=1.67
+ $X2=11.73 $Y2=1.76
r214 60 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=2.035
+ $X2=12.24 $Y2=2.035
r215 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r216 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r217 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=2.035
+ $X2=12.24 $Y2=2.035
r218 53 54 10.3341 $w=1.4e-07 $l=8.35e-06 $layer=MET1_cond $X=12.095 $Y=2.035
+ $X2=3.745 $Y2=2.035
r219 52 57 14.5035 $w=1.93e-07 $l=2.55e-07 $layer=LI1_cond $X=3.587 $Y=1.78
+ $X2=3.587 $Y2=2.035
r220 50 65 21.1993 $w=5.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.555 $Y=1.615
+ $X2=3.555 $Y2=1.825
r221 50 64 47.4091 $w=5.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.615
+ $X2=3.555 $Y2=1.45
r222 49 52 7.67512 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=1.615
+ $X2=3.655 $Y2=1.78
r223 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=1.615 $X2=3.655 $Y2=1.615
r224 45 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.85 $Y=1.49
+ $X2=12.85 $Y2=1.655
r225 45 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.85 $Y=1.49
+ $X2=12.85 $Y2=1.325
r226 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.85
+ $Y=1.49 $X2=12.85 $Y2=1.49
r227 42 78 3.76816 $w=3.3e-07 $l=3.95e-07 $layer=LI1_cond $X=12.355 $Y=1.49
+ $X2=11.96 $Y2=1.49
r228 42 44 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=12.355 $Y=1.49
+ $X2=12.85 $Y2=1.49
r229 38 78 5.61216 $w=5.54e-07 $l=1.94808e-07 $layer=LI1_cond $X=12.025 $Y=1.325
+ $X2=11.96 $Y2=1.49
r230 38 40 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=12.025 $Y=1.325
+ $X2=12.025 $Y2=0.98
r231 35 37 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=11.13 $Y=1.67
+ $X2=11.28 $Y2=1.67
r232 33 75 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=12.94 $Y=2.445
+ $X2=12.94 $Y2=1.655
r233 29 74 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=12.83 $Y=0.705
+ $X2=12.83 $Y2=1.325
r234 26 37 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.355 $Y=1.67
+ $X2=11.28 $Y2=1.67
r235 25 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.565 $Y=1.67
+ $X2=11.73 $Y2=1.67
r236 25 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=11.565 $Y=1.67
+ $X2=11.355 $Y2=1.67
r237 21 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.28 $Y=1.745
+ $X2=11.28 $Y2=1.67
r238 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=11.28 $Y=1.745
+ $X2=11.28 $Y2=2.295
r239 17 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.13 $Y=1.595
+ $X2=11.13 $Y2=1.67
r240 17 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=11.13 $Y=1.595
+ $X2=11.13 $Y2=0.915
r241 15 64 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.365 $Y=0.77
+ $X2=3.365 $Y2=1.45
r242 11 65 32.8864 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.29 $Y=1.825
+ $X2=3.555 $Y2=1.825
r243 11 12 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=3.29 $Y=1.825
+ $X2=3.085 $Y2=1.825
r244 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.01 $Y=1.9
+ $X2=3.085 $Y2=1.825
r245 7 9 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.01 $Y=1.9 $X2=3.01
+ $Y2=2.325
r246 2 81 600 $w=1.7e-07 $l=2.20624e-07 $layer=licon1_PDIFF $count=1 $X=12.055
+ $Y=1.815 $X2=12.185 $Y2=1.98
r247 1 40 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=11.89
+ $Y=0.705 $X2=12.025 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_958_290# 1 2 9 13 17 21 26 31 35 36 37 39
+ 40 46 53 54 57 62 63
c145 53 0 1.52339e-20 $X=5.08 $Y=1.615
c146 39 0 1.92769e-19 $X=8.255 $Y=1.665
r147 62 63 3.86001 $w=3.83e-07 $l=8.5e-08 $layer=LI1_cond $X=8.477 $Y=1.47
+ $X2=8.477 $Y2=1.385
r148 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.08
+ $Y=1.615 $X2=5.08 $Y2=1.615
r149 51 53 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.945 $Y=1.615
+ $X2=5.08 $Y2=1.615
r150 49 51 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=4.865 $Y=1.615
+ $X2=4.945 $Y2=1.615
r151 47 65 4.85718 $w=3.83e-07 $l=1.15e-07 $layer=LI1_cond $X=8.477 $Y=1.665
+ $X2=8.477 $Y2=1.78
r152 47 62 5.83705 $w=3.83e-07 $l=1.95e-07 $layer=LI1_cond $X=8.477 $Y=1.665
+ $X2=8.477 $Y2=1.47
r153 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r154 42 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r155 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r156 39 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r157 39 40 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.185 $Y2=1.665
r158 36 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.785 $Y=1.41
+ $X2=9.785 $Y2=1.575
r159 36 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.785 $Y=1.41
+ $X2=9.785 $Y2=1.245
r160 35 37 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=9.785 $Y=1.4
+ $X2=9.62 $Y2=1.4
r161 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.785
+ $Y=1.41 $X2=9.785 $Y2=1.41
r162 33 63 21.0151 $w=2.53e-07 $l=4.65e-07 $layer=LI1_cond $X=8.412 $Y=0.92
+ $X2=8.412 $Y2=1.385
r163 31 33 8.65746 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=8.375 $Y=0.69
+ $X2=8.375 $Y2=0.92
r164 29 62 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=8.67 $Y=1.47
+ $X2=8.477 $Y2=1.47
r165 29 37 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=8.67 $Y=1.47
+ $X2=9.62 $Y2=1.47
r166 26 65 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=8.545 $Y=2.145
+ $X2=8.545 $Y2=1.78
r167 21 57 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=9.855 $Y=0.705
+ $X2=9.855 $Y2=1.245
r168 17 58 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.78 $Y=2.15
+ $X2=9.78 $Y2=1.575
r169 11 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.945 $Y=1.45
+ $X2=4.945 $Y2=1.615
r170 11 13 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=4.945 $Y=1.45
+ $X2=4.945 $Y2=0.665
r171 7 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.865 $Y=1.78
+ $X2=4.865 $Y2=1.615
r172 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.865 $Y=1.78
+ $X2=4.865 $Y2=2.19
r173 2 26 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=8.365
+ $Y=1.98 $X2=8.505 $Y2=2.145
r174 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.235
+ $Y=0.48 $X2=8.375 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_1067_65# 1 2 9 12 15 19 23 27 29 37 39 40
+ 41 43 44 45 47 48 49 51 52 53 56 57 62 64 68
c197 53 0 1.8865e-19 $X=9.12 $Y=1.82
c198 27 0 9.64333e-20 $X=5.56 $Y=1.135
r199 60 62 7.19862 $w=5.38e-07 $l=3.25e-07 $layer=LI1_cond $X=6.25 $Y=0.535
+ $X2=6.575 $Y2=0.535
r200 57 70 17.7061 $w=2.45e-07 $l=9e-08 $layer=POLY_cond $X=10.355 $Y=1.51
+ $X2=10.265 $Y2=1.51
r201 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.355
+ $Y=1.51 $X2=10.355 $Y2=1.51
r202 54 56 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=10.355 $Y=1.735
+ $X2=10.355 $Y2=1.51
r203 52 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.19 $Y=1.82
+ $X2=10.355 $Y2=1.735
r204 52 53 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=10.19 $Y=1.82
+ $X2=9.12 $Y2=1.82
r205 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.035 $Y=1.905
+ $X2=9.12 $Y2=1.82
r206 50 51 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.035 $Y=1.905
+ $X2=9.035 $Y2=2.515
r207 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.95 $Y=2.6
+ $X2=9.035 $Y2=2.515
r208 48 49 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.95 $Y=2.6
+ $X2=8.24 $Y2=2.6
r209 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.155 $Y=2.515
+ $X2=8.24 $Y2=2.6
r210 46 47 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.155 $Y=2.13
+ $X2=8.155 $Y2=2.515
r211 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.07 $Y=2.045
+ $X2=8.155 $Y2=2.13
r212 44 45 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.07 $Y=2.045
+ $X2=7.54 $Y2=2.045
r213 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.455 $Y=2.13
+ $X2=7.54 $Y2=2.045
r214 42 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.455 $Y=2.13
+ $X2=7.455 $Y2=2.82
r215 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.37 $Y=2.905
+ $X2=7.455 $Y2=2.82
r216 40 41 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.37 $Y=2.905
+ $X2=6.66 $Y2=2.905
r217 39 64 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=6.575 $Y=1.555
+ $X2=6.535 $Y2=1.72
r218 38 62 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=6.575 $Y=0.805
+ $X2=6.575 $Y2=0.535
r219 38 39 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.575 $Y=0.805
+ $X2=6.575 $Y2=1.555
r220 35 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.535 $Y=2.82
+ $X2=6.66 $Y2=2.905
r221 35 37 37.3392 $w=2.48e-07 $l=8.1e-07 $layer=LI1_cond $X=6.535 $Y=2.82
+ $X2=6.535 $Y2=2.01
r222 34 64 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=1.885
+ $X2=6.535 $Y2=1.72
r223 34 37 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=1.885
+ $X2=6.535 $Y2=2.01
r224 32 68 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.685 $Y=1.72
+ $X2=5.825 $Y2=1.72
r225 32 65 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.685 $Y=1.72
+ $X2=5.56 $Y2=1.72
r226 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.685
+ $Y=1.72 $X2=5.685 $Y2=1.72
r227 29 64 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=1.72
+ $X2=6.535 $Y2=1.72
r228 29 31 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=6.41 $Y=1.72
+ $X2=5.685 $Y2=1.72
r229 25 27 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.41 $Y=1.135
+ $X2=5.56 $Y2=1.135
r230 21 57 75.7429 $w=2.45e-07 $l=4.60163e-07 $layer=POLY_cond $X=10.74 $Y=1.675
+ $X2=10.355 $Y2=1.51
r231 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.74 $Y=1.675
+ $X2=10.74 $Y2=2.465
r232 17 70 14.2527 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.265 $Y=1.345
+ $X2=10.265 $Y2=1.51
r233 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=10.265 $Y=1.345
+ $X2=10.265 $Y2=0.705
r234 13 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.885
+ $X2=5.825 $Y2=1.72
r235 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.825 $Y=1.885
+ $X2=5.825 $Y2=2.495
r236 12 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=1.555
+ $X2=5.56 $Y2=1.72
r237 11 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.56 $Y=1.21
+ $X2=5.56 $Y2=1.135
r238 11 12 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=5.56 $Y=1.21
+ $X2=5.56 $Y2=1.555
r239 7 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.41 $Y=1.06
+ $X2=5.41 $Y2=1.135
r240 7 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.41 $Y=1.06
+ $X2=5.41 $Y2=0.665
r241 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.435
+ $Y=1.865 $X2=6.575 $Y2=2.01
r242 1 60 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=6.11
+ $Y=0.235 $X2=6.25 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_902_396# 1 2 7 9 12 16 20 24 26 28 33
c72 26 0 9.64333e-20 $X=6.135 $Y=1.15
r73 27 33 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=6.135 $Y=1.15
+ $X2=6.36 $Y2=1.15
r74 27 30 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.135 $Y=1.15
+ $X2=6.035 $Y2=1.15
r75 26 28 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.135 $Y=1.15
+ $X2=5.97 $Y2=1.15
r76 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.135
+ $Y=1.15 $X2=6.135 $Y2=1.15
r77 23 24 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=1.16
+ $X2=4.73 $Y2=1.16
r78 23 28 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=4.895 $Y=1.16
+ $X2=5.97 $Y2=1.16
r79 18 24 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.65 $Y=1.245
+ $X2=4.73 $Y2=1.16
r80 18 20 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=4.65 $Y=1.245
+ $X2=4.65 $Y2=2.16
r81 14 24 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=1.075
+ $X2=4.73 $Y2=1.16
r82 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.73 $Y=1.075
+ $X2=4.73 $Y2=0.665
r83 10 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.36 $Y=1.315
+ $X2=6.36 $Y2=1.15
r84 10 12 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=6.36 $Y=1.315
+ $X2=6.36 $Y2=2.285
r85 7 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.035 $Y=0.985
+ $X2=6.035 $Y2=1.15
r86 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.035 $Y=0.985
+ $X2=6.035 $Y2=0.555
r87 2 20 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=4.51 $Y=1.98
+ $X2=4.65 $Y2=2.16
r88 1 16 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.55
+ $Y=0.455 $X2=4.73 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%CLK 1 5 9 12 15 17 18 20
c54 20 0 7.72461e-20 $X=7.005 $Y=1.175
c55 18 0 6.21449e-20 $X=6.96 $Y=1.295
c56 15 0 8.80718e-20 $X=7.46 $Y=1.745
r57 20 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.005 $Y=1.175
+ $X2=7.005 $Y2=1.265
r58 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.005
+ $Y=1.265 $X2=7.005 $Y2=1.265
r59 13 15 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=7.32 $Y=1.745
+ $X2=7.46 $Y2=1.745
r60 12 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.46 $Y=1.67
+ $X2=7.46 $Y2=1.745
r61 11 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.46 $Y=1.25
+ $X2=7.46 $Y2=1.175
r62 11 12 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=7.46 $Y=1.25
+ $X2=7.46 $Y2=1.67
r63 7 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.46 $Y=1.1 $X2=7.46
+ $Y2=1.175
r64 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.46 $Y=1.1 $X2=7.46
+ $Y2=0.69
r65 3 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.32 $Y=1.82 $X2=7.32
+ $Y2=1.745
r66 3 5 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.32 $Y=1.82 $X2=7.32
+ $Y2=2.3
r67 2 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.17 $Y=1.175
+ $X2=7.005 $Y2=1.175
r68 1 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.385 $Y=1.175
+ $X2=7.46 $Y2=1.175
r69 1 2 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=7.385 $Y=1.175
+ $X2=7.17 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_872_324# 1 2 10 13 15 16 21 26 27 29 31
+ 34 37 38 39 41 44 47 49 50 56 59 61 63 64
c173 64 0 6.21449e-20 $X=7.94 $Y=1.265
c174 61 0 2.02548e-19 $X=7.435 $Y=1.185
c175 49 0 8.80718e-20 $X=7.435 $Y=1.61
c176 38 0 1.8865e-19 $X=8.07 $Y=1.65
c177 37 0 1.61716e-19 $X=4.455 $Y=1.77
c178 29 0 9.76166e-20 $X=9.25 $Y=1.725
r179 64 66 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=8.005 $Y=1.265
+ $X2=8.005 $Y2=1.1
r180 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.94
+ $Y=1.265 $X2=7.94 $Y2=1.265
r181 51 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.52 $Y=1.185
+ $X2=7.435 $Y2=1.185
r182 50 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.775 $Y=1.185
+ $X2=7.94 $Y2=1.185
r183 50 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.775 $Y=1.185
+ $X2=7.52 $Y2=1.185
r184 49 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=1.61
+ $X2=7.435 $Y2=1.695
r185 48 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=1.27
+ $X2=7.435 $Y2=1.185
r186 48 49 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.435 $Y=1.27
+ $X2=7.435 $Y2=1.61
r187 47 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=1.1
+ $X2=7.435 $Y2=1.185
r188 46 59 12.6565 $w=2.94e-07 $l=3.88555e-07 $layer=LI1_cond $X=7.435 $Y=0.92
+ $X2=7.13 $Y2=0.73
r189 46 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.435 $Y=0.92
+ $X2=7.435 $Y2=1.1
r190 42 56 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.065 $Y=1.695
+ $X2=7.435 $Y2=1.695
r191 42 44 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=7.065 $Y=1.78
+ $X2=7.065 $Y2=2.125
r192 38 40 45.1092 $w=5.9e-07 $l=1.2e-07 $layer=POLY_cond $X=8.07 $Y=1.65
+ $X2=8.07 $Y2=1.77
r193 38 39 9.54275 $w=5.9e-07 $l=7.5e-08 $layer=POLY_cond $X=8.07 $Y=1.65
+ $X2=8.07 $Y2=1.575
r194 36 37 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=4.455 $Y=1.62
+ $X2=4.455 $Y2=1.77
r195 32 41 20.4101 $w=1.5e-07 $l=8.7892e-08 $layer=POLY_cond $X=9.305 $Y=1.575
+ $X2=9.277 $Y2=1.65
r196 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.305 $Y=1.575
+ $X2=9.305 $Y2=0.915
r197 29 41 20.4101 $w=1.5e-07 $l=8.74643e-08 $layer=POLY_cond $X=9.25 $Y=1.725
+ $X2=9.277 $Y2=1.65
r198 29 31 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.25 $Y=1.725
+ $X2=9.25 $Y2=2.465
r199 28 38 35.6395 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=8.365 $Y=1.65
+ $X2=8.07 $Y2=1.65
r200 27 41 5.30422 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=9.175 $Y=1.65
+ $X2=9.277 $Y2=1.65
r201 27 28 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.175 $Y=1.65
+ $X2=8.365 $Y2=1.65
r202 26 40 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.29 $Y=2.3
+ $X2=8.29 $Y2=1.77
r203 24 26 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=8.29 $Y=3.075
+ $X2=8.29 $Y2=2.3
r204 21 66 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.16 $Y=0.69
+ $X2=8.16 $Y2=1.1
r205 17 64 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=8.005 $Y=1.33
+ $X2=8.005 $Y2=1.265
r206 17 39 29.6212 $w=4.6e-07 $l=2.45e-07 $layer=POLY_cond $X=8.005 $Y=1.33
+ $X2=8.005 $Y2=1.575
r207 15 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.215 $Y=3.15
+ $X2=8.29 $Y2=3.075
r208 15 16 1899.8 $w=1.5e-07 $l=3.705e-06 $layer=POLY_cond $X=8.215 $Y=3.15
+ $X2=4.51 $Y2=3.15
r209 13 36 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=4.475 $Y=0.665
+ $X2=4.475 $Y2=1.62
r210 10 37 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.435 $Y=2.19
+ $X2=4.435 $Y2=1.77
r211 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.435 $Y=3.075
+ $X2=4.51 $Y2=3.15
r212 8 10 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=4.435 $Y=3.075
+ $X2=4.435 $Y2=2.19
r213 2 44 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=6.975
+ $Y=1.98 $X2=7.105 $Y2=2.125
r214 1 59 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.985
+ $Y=0.48 $X2=7.13 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_1865_367# 1 2 8 9 10 11 13 16 18 20 23 26
+ 28 31 32 39 40 42 45 46 47 51 54 58 59 60 64 65 72
c182 46 0 1.75981e-19 $X=13.54 $Y=2.43
c183 18 0 1.44709e-19 $X=13.915 $Y=1.185
r184 71 72 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=13.915 $Y=1.35
+ $X2=13.92 $Y2=1.35
r185 64 65 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=11.8 $Y=0.49
+ $X2=11.97 $Y2=0.49
r186 60 62 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.305 $Y=2.52
+ $X2=11.305 $Y2=2.79
r187 58 59 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=10.94 $Y=0.49
+ $X2=11.11 $Y2=0.49
r188 54 56 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=9.635 $Y=0.49
+ $X2=9.635 $Y2=0.63
r189 52 71 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=13.705 $Y=1.35
+ $X2=13.915 $Y2=1.35
r190 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.705
+ $Y=1.35 $X2=13.705 $Y2=1.35
r191 49 51 35.2825 $w=3.23e-07 $l=9.95e-07 $layer=LI1_cond $X=13.702 $Y=2.345
+ $X2=13.702 $Y2=1.35
r192 48 51 22.517 $w=3.23e-07 $l=6.35e-07 $layer=LI1_cond $X=13.702 $Y=0.715
+ $X2=13.702 $Y2=1.35
r193 46 49 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=13.54 $Y=2.43
+ $X2=13.702 $Y2=2.345
r194 46 47 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=13.54 $Y=2.43
+ $X2=12.38 $Y2=2.43
r195 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.295 $Y=2.515
+ $X2=12.38 $Y2=2.43
r196 44 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.295 $Y=2.515
+ $X2=12.295 $Y2=2.705
r197 42 48 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=13.54 $Y=0.63
+ $X2=13.702 $Y2=0.715
r198 42 65 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=13.54 $Y=0.63
+ $X2=11.97 $Y2=0.63
r199 41 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.39 $Y=2.79
+ $X2=11.305 $Y2=2.79
r200 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.21 $Y=2.79
+ $X2=12.295 $Y2=2.705
r201 40 41 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=12.21 $Y=2.79
+ $X2=11.39 $Y2=2.79
r202 39 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.65 $Y=0.43
+ $X2=11.65 $Y2=0.595
r203 38 64 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=11.65 $Y=0.43
+ $X2=11.8 $Y2=0.43
r204 38 59 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=11.65 $Y=0.43
+ $X2=11.11 $Y2=0.43
r205 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.65
+ $Y=0.43 $X2=11.65 $Y2=0.43
r206 34 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.8 $Y=0.63
+ $X2=9.635 $Y2=0.63
r207 34 58 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=9.8 $Y=0.63
+ $X2=10.94 $Y2=0.63
r208 31 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=2.52
+ $X2=11.305 $Y2=2.52
r209 31 32 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=11.22 $Y=2.52
+ $X2=9.63 $Y2=2.52
r210 28 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.465 $Y=2.435
+ $X2=9.63 $Y2=2.52
r211 28 30 1.84848 $w=3.3e-07 $l=5e-08 $layer=LI1_cond $X=9.465 $Y=2.435
+ $X2=9.465 $Y2=2.385
r212 25 26 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=12.24 $Y=1.31
+ $X2=12.4 $Y2=1.31
r213 21 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.92 $Y=1.515
+ $X2=13.92 $Y2=1.35
r214 21 23 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=13.92 $Y=1.515
+ $X2=13.92 $Y2=2.465
r215 18 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.915 $Y=1.185
+ $X2=13.915 $Y2=1.35
r216 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.915 $Y=1.185
+ $X2=13.915 $Y2=0.655
r217 14 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.4 $Y=1.385
+ $X2=12.4 $Y2=1.31
r218 14 16 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=12.4 $Y=1.385
+ $X2=12.4 $Y2=2.135
r219 11 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.24 $Y=1.235
+ $X2=12.24 $Y2=1.31
r220 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.24 $Y=1.235
+ $X2=12.24 $Y2=0.915
r221 9 25 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.165 $Y=1.31
+ $X2=12.24 $Y2=1.31
r222 9 10 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=12.165 $Y=1.31
+ $X2=11.815 $Y2=1.31
r223 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.74 $Y=1.235
+ $X2=11.815 $Y2=1.31
r224 8 68 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=11.74 $Y=1.235
+ $X2=11.74 $Y2=0.595
r225 2 30 600 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=1 $X=9.325
+ $Y=1.835 $X2=9.465 $Y2=2.385
r226 1 54 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=9.38
+ $Y=0.705 $X2=9.635 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48
+ 51 52 54 55 57 58 59 68 85 92 99 100 106 109 112
c140 100 0 6.76474e-20 $X=14.16 $Y=3.33
c141 32 0 1.92769e-19 $X=6.145 $Y=2.395
r142 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r143 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r144 106 107 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r145 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 100 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r147 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r148 97 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.87 $Y=3.33
+ $X2=13.705 $Y2=3.33
r149 97 99 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.87 $Y=3.33
+ $X2=14.16 $Y2=3.33
r150 96 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r151 96 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r152 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r153 93 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.89 $Y=3.33
+ $X2=12.725 $Y2=3.33
r154 93 95 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=12.89 $Y=3.33
+ $X2=13.2 $Y2=3.33
r155 92 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.705 $Y2=3.33
r156 92 95 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.2 $Y2=3.33
r157 91 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r158 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r159 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r160 87 90 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r161 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r162 85 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.56 $Y=3.33
+ $X2=12.725 $Y2=3.33
r163 85 90 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.56 $Y=3.33
+ $X2=12.24 $Y2=3.33
r164 84 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r165 83 84 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r166 81 84 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.8 $Y2=3.33
r167 80 83 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.8 $Y2=3.33
r168 80 81 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r169 78 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r170 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r171 75 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r172 74 77 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r173 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r174 72 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.23 $Y=3.33
+ $X2=6.105 $Y2=3.33
r175 72 74 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.23 $Y=3.33
+ $X2=6.48 $Y2=3.33
r176 71 107 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=6 $Y2=3.33
r177 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r178 68 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=6.105 $Y2=3.33
r179 68 70 249.219 $w=1.68e-07 $l=3.82e-06 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 67 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r181 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r182 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r183 64 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r184 63 66 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r185 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r186 61 103 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r187 61 63 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.72 $Y2=3.33
r188 59 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r189 59 75 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 57 83 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=10.87 $Y=3.33
+ $X2=10.8 $Y2=3.33
r191 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.87 $Y=3.33
+ $X2=10.955 $Y2=3.33
r192 56 87 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=11.28 $Y2=3.33
r193 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=10.955 $Y2=3.33
r194 54 77 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.72 $Y=3.33
+ $X2=7.44 $Y2=3.33
r195 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.72 $Y=3.33
+ $X2=7.805 $Y2=3.33
r196 53 80 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=7.89 $Y=3.33 $X2=7.92
+ $Y2=3.33
r197 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=3.33
+ $X2=7.805 $Y2=3.33
r198 51 66 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r199 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=2.005 $Y2=3.33
r200 50 70 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.09 $Y=3.33 $X2=2.16
+ $Y2=3.33
r201 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=3.33
+ $X2=2.005 $Y2=3.33
r202 46 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=3.33
r203 46 48 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=2.905
r204 42 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.725 $Y=3.245
+ $X2=12.725 $Y2=3.33
r205 42 44 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.725 $Y=3.245
+ $X2=12.725 $Y2=2.895
r206 38 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.955 $Y=3.245
+ $X2=10.955 $Y2=3.33
r207 38 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.955 $Y=3.245
+ $X2=10.955 $Y2=2.95
r208 34 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.805 $Y=3.245
+ $X2=7.805 $Y2=3.33
r209 34 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.805 $Y=3.245
+ $X2=7.805 $Y2=2.475
r210 30 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.105 $Y=3.245
+ $X2=6.105 $Y2=3.33
r211 30 32 39.1831 $w=2.48e-07 $l=8.5e-07 $layer=LI1_cond $X=6.105 $Y=3.245
+ $X2=6.105 $Y2=2.395
r212 26 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=3.245
+ $X2=2.005 $Y2=3.33
r213 26 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.005 $Y=3.245
+ $X2=2.005 $Y2=2.325
r214 22 103 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.197 $Y2=3.33
r215 22 24 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.55
r216 7 48 600 $w=1.7e-07 $l=1.13785e-06 $layer=licon1_PDIFF $count=1 $X=13.565
+ $Y=1.835 $X2=13.705 $Y2=2.905
r217 6 44 600 $w=1.7e-07 $l=1.1985e-06 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.815 $X2=12.725 $Y2=2.895
r218 5 40 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.815
+ $Y=1.835 $X2=10.955 $Y2=2.95
r219 4 36 600 $w=1.7e-07 $l=6.69309e-07 $layer=licon1_PDIFF $count=1 $X=7.395
+ $Y=1.98 $X2=7.805 $Y2=2.475
r220 3 32 600 $w=1.7e-07 $l=2.94915e-07 $layer=licon1_PDIFF $count=1 $X=5.9
+ $Y=2.285 $X2=6.145 $Y2=2.395
r221 2 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=2.115 $X2=2.005 $Y2=2.325
r222 1 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.405 $X2=0.31 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_286_423# 1 2 9 11 12 14 15 16 19
c49 9 0 1.3912e-19 $X=1.575 $Y=2.325
r50 17 19 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.185 $Y=2.735
+ $X2=3.185 $Y2=2.325
r51 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.06 $Y=2.82
+ $X2=3.185 $Y2=2.735
r52 15 16 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.06 $Y=2.82
+ $X2=2.44 $Y2=2.82
r53 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.355 $Y=2.735
+ $X2=2.44 $Y2=2.82
r54 13 14 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.355 $Y=1.915
+ $X2=2.355 $Y2=2.735
r55 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.27 $Y=1.83
+ $X2=2.355 $Y2=1.915
r56 11 12 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.27 $Y=1.83
+ $X2=1.74 $Y2=1.83
r57 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.615 $Y=1.915
+ $X2=1.74 $Y2=1.83
r58 7 9 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.615 $Y=1.915
+ $X2=1.615 $Y2=2.325
r59 2 19 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=2.115 $X2=3.225 $Y2=2.325
r60 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=2.115 $X2=1.575 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_531_423# 1 2 3 4 15 17 18 19 20 21 25 28
+ 29 30 33 38
c91 18 0 1.35708e-19 $X=2.88 $Y=1.83
r92 36 37 17.4286 $w=2.66e-07 $l=3.8e-07 $layer=LI1_cond $X=3.15 $Y=0.805
+ $X2=3.15 $Y2=1.185
r93 31 33 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.08 $Y=2.545
+ $X2=5.08 $Y2=2.19
r94 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.915 $Y=2.63
+ $X2=5.08 $Y2=2.545
r95 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.915 $Y=2.63
+ $X2=4.385 $Y2=2.63
r96 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.3 $Y=2.545
+ $X2=4.385 $Y2=2.63
r97 27 38 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.3 $Y=1.27
+ $X2=4.22 $Y2=1.185
r98 27 28 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=4.3 $Y=1.27
+ $X2=4.3 $Y2=2.545
r99 23 38 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.22 $Y=1.1 $X2=4.22
+ $Y2=1.185
r100 23 25 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.22 $Y=1.1
+ $X2=4.22 $Y2=0.665
r101 22 37 3.35683 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=1.185
+ $X2=3.15 $Y2=1.185
r102 21 38 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=1.185
+ $X2=4.22 $Y2=1.185
r103 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.055 $Y=1.185
+ $X2=3.315 $Y2=1.185
r104 19 37 5.48216 $w=2.66e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.225 $Y=1.27
+ $X2=3.15 $Y2=1.185
r105 19 20 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.225 $Y=1.27
+ $X2=3.225 $Y2=1.745
r106 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.14 $Y=1.83
+ $X2=3.225 $Y2=1.745
r107 17 18 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.14 $Y=1.83
+ $X2=2.88 $Y2=1.83
r108 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.755 $Y=1.915
+ $X2=2.88 $Y2=1.83
r109 13 15 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=2.755 $Y=1.915
+ $X2=2.755 $Y2=2.325
r110 4 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.94
+ $Y=1.98 $X2=5.08 $Y2=2.19
r111 3 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.655
+ $Y=2.115 $X2=2.795 $Y2=2.325
r112 2 25 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.455 $X2=4.22 $Y2=0.665
r113 1 36 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.56 $X2=3.15 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_761_396# 1 2 9 11 12 15
r33 13 15 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.61 $Y=2.895 $X2=5.61
+ $Y2=2.495
r34 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.445 $Y=2.98
+ $X2=5.61 $Y2=2.895
r35 11 12 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=5.445 $Y=2.98
+ $X2=4.035 $Y2=2.98
r36 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.95 $Y=2.895
+ $X2=4.035 $Y2=2.98
r37 7 9 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.95 $Y=2.895
+ $X2=3.95 $Y2=2.19
r38 2 15 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=5.48
+ $Y=2.285 $X2=5.61 $Y2=2.495
r39 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=1.98 $X2=3.95 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_1781_367# 1 2 12 13
r23 12 13 7.74904 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=10.525 $Y=2.925
+ $X2=10.36 $Y2=2.925
r24 9 13 73.4773 $w=1.98e-07 $l=1.325e-06 $layer=LI1_cond $X=9.035 $Y=2.965
+ $X2=10.36 $Y2=2.965
r25 2 12 600 $w=1.7e-07 $l=1.1131e-06 $layer=licon1_PDIFF $count=1 $X=10.395
+ $Y=1.835 $X2=10.525 $Y2=2.885
r26 1 9 600 $w=1.7e-07 $l=1.17821e-06 $layer=licon1_PDIFF $count=1 $X=8.905
+ $Y=1.835 $X2=9.035 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_1971_388# 1 2 7 11
c28 7 0 2.09147e-19 $X=11.57 $Y=2.17
r29 11 14 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=11.695 $Y=2.17
+ $X2=11.695 $Y2=2.305
r30 7 11 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.57 $Y=2.17
+ $X2=11.695 $Y2=2.17
r31 7 9 102.754 $w=1.68e-07 $l=1.575e-06 $layer=LI1_cond $X=11.57 $Y=2.17
+ $X2=9.995 $Y2=2.17
r32 2 14 600 $w=1.7e-07 $l=3.94968e-07 $layer=licon1_PDIFF $count=1 $X=11.355
+ $Y=2.085 $X2=11.655 $Y2=2.305
r33 1 9 600 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=1 $X=9.855
+ $Y=1.94 $X2=9.995 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%Q_N 1 2 7 12 13 14 18
c27 12 0 1.44709e-19 $X=13.275 $Y=1.835
r28 14 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.275 $Y=2 $X2=13.19
+ $Y2=2
r29 14 18 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=13.152 $Y=2
+ $X2=13.19 $Y2=2
r30 13 14 15.0865 $w=3.28e-07 $l=4.32e-07 $layer=LI1_cond $X=12.72 $Y=2
+ $X2=13.152 $Y2=2
r31 12 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.275 $Y=1.835
+ $X2=13.275 $Y2=2
r32 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.275 $Y=1.145
+ $X2=13.275 $Y2=1.835
r33 7 11 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.19 $Y=1.02
+ $X2=13.275 $Y2=1.145
r34 7 9 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=13.19 $Y=1.02
+ $X2=13.045 $Y2=1.02
r35 2 14 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=13.015
+ $Y=1.815 $X2=13.155 $Y2=2
r36 1 9 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=12.905
+ $Y=0.285 $X2=13.045 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%Q 1 2 9 11 12 13 14 15 24 37
r13 22 37 0.542326 $w=2.53e-07 $l=1.2e-08 $layer=LI1_cond $X=14.172 $Y=2.023
+ $X2=14.172 $Y2=2.035
r14 15 39 3.57031 $w=2.53e-07 $l=7.9e-08 $layer=LI1_cond $X=14.172 $Y=2.071
+ $X2=14.172 $Y2=2.15
r15 15 37 1.62698 $w=2.53e-07 $l=3.6e-08 $layer=LI1_cond $X=14.172 $Y=2.071
+ $X2=14.172 $Y2=2.035
r16 15 22 1.94334 $w=2.53e-07 $l=4.3e-08 $layer=LI1_cond $X=14.172 $Y=1.98
+ $X2=14.172 $Y2=2.023
r17 14 15 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=14.172 $Y=1.665
+ $X2=14.172 $Y2=1.98
r18 13 14 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=14.172 $Y=1.295
+ $X2=14.172 $Y2=1.665
r19 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=14.172 $Y=0.925
+ $X2=14.172 $Y2=1.295
r20 11 12 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=14.172 $Y=0.555
+ $X2=14.172 $Y2=0.925
r21 11 24 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=14.172 $Y=0.555
+ $X2=14.172 $Y2=0.43
r22 9 39 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=14.175 $Y=2.44
+ $X2=14.175 $Y2=2.15
r23 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.995
+ $Y=1.835 $X2=14.135 $Y2=1.98
r24 2 9 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=13.995
+ $Y=1.835 $X2=14.135 $Y2=2.44
r25 1 24 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=13.99
+ $Y=0.235 $X2=14.13 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%VGND 1 2 3 4 5 6 7 22 24 28 32 36 38 39 45
+ 46 52 53 59 61 66 71 96 97 103 106 109
r125 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r126 106 107 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r127 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r128 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r129 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r130 94 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r131 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r132 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r133 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r134 88 91 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=12.24 $Y2=0
r135 87 90 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=10.8 $Y=0
+ $X2=12.24 $Y2=0
r136 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r137 85 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r138 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r139 82 85 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r140 82 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r141 81 84 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.32
+ $Y2=0
r142 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r143 79 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.03 $Y=0
+ $X2=7.865 $Y2=0
r144 79 81 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=8.4
+ $Y2=0
r145 78 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r146 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r147 75 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r148 74 77 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.44
+ $Y2=0
r149 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r150 72 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.79 $Y=0
+ $X2=5.625 $Y2=0
r151 72 74 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.79 $Y=0 $X2=6
+ $Y2=0
r152 71 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.7 $Y=0 $X2=7.865
+ $Y2=0
r153 71 77 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.7 $Y=0 $X2=7.44
+ $Y2=0
r154 70 107 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=5.52 $Y2=0
r155 70 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r156 69 70 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r157 67 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=0
+ $X2=1.69 $Y2=0
r158 67 69 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=2.16
+ $Y2=0
r159 66 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=0
+ $X2=5.625 $Y2=0
r160 66 69 215.294 $w=1.68e-07 $l=3.3e-06 $layer=LI1_cond $X=5.46 $Y=0 $X2=2.16
+ $Y2=0
r161 65 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r162 65 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r163 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r164 62 100 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r165 62 64 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=1.2
+ $Y2=0
r166 61 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.565 $Y=0
+ $X2=1.69 $Y2=0
r167 61 64 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.2
+ $Y2=0
r168 59 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=7.44
+ $Y2=0
r169 59 75 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=6
+ $Y2=0
r170 55 96 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=13.75 $Y=0
+ $X2=14.16 $Y2=0
r171 53 93 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=13.42 $Y=0 $X2=13.2
+ $Y2=0
r172 52 57 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=13.585 $Y=0
+ $X2=13.585 $Y2=0.28
r173 52 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.585 $Y=0
+ $X2=13.75 $Y2=0
r174 52 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.585 $Y=0
+ $X2=13.42 $Y2=0
r175 48 93 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=12.7 $Y=0 $X2=13.2
+ $Y2=0
r176 46 90 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=12.37 $Y=0
+ $X2=12.24 $Y2=0
r177 45 50 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=12.535 $Y=0
+ $X2=12.535 $Y2=0.28
r178 45 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.535 $Y=0
+ $X2=12.7 $Y2=0
r179 45 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.535 $Y=0
+ $X2=12.37 $Y2=0
r180 41 87 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=10.76 $Y=0 $X2=10.8
+ $Y2=0
r181 39 84 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=10.43 $Y=0
+ $X2=10.32 $Y2=0
r182 38 43 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.595 $Y2=0.28
r183 38 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.76 $Y2=0
r184 38 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.43 $Y2=0
r185 34 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=0.085
+ $X2=7.865 $Y2=0
r186 34 36 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=7.865 $Y=0.085
+ $X2=7.865 $Y2=0.69
r187 30 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=0.085
+ $X2=5.625 $Y2=0
r188 30 32 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=5.625 $Y=0.085
+ $X2=5.625 $Y2=0.665
r189 26 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0
r190 26 28 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0.475
r191 22 100 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.197 $Y2=0
r192 22 24 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=1.105
r193 7 57 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=13.45
+ $Y=0.135 $X2=13.585 $Y2=0.28
r194 6 50 182 $w=1.7e-07 $l=5.23569e-07 $layer=licon1_NDIFF $count=1 $X=12.315
+ $Y=0.705 $X2=12.535 $Y2=0.28
r195 5 43 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=10.34
+ $Y=0.285 $X2=10.595 $Y2=0.28
r196 4 36 182 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_NDIFF $count=1 $X=7.535
+ $Y=0.48 $X2=7.865 $Y2=0.69
r197 3 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.485
+ $Y=0.455 $X2=5.625 $Y2=0.665
r198 2 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.265 $X2=1.73 $Y2=0.475
r199 1 24 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.895 $X2=0.31 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_231_53# 1 2 9 12 13 15 16 18
c36 16 0 1.63805e-19 $X=2.165 $Y=0.942
r37 18 20 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=2.68 $Y=0.805
+ $X2=2.68 $Y2=0.915
r38 15 16 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.995 $Y=0.942
+ $X2=2.165 $Y2=0.942
r39 13 20 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=0.915
+ $X2=2.68 $Y2=0.915
r40 13 16 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.555 $Y=0.915
+ $X2=2.165 $Y2=0.915
r41 12 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.385 $Y=0.97
+ $X2=1.995 $Y2=0.97
r42 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.26 $Y=0.885
+ $X2=1.385 $Y2=0.97
r43 7 9 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.26 $Y=0.885 $X2=1.26
+ $Y2=0.485
r44 2 18 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.56 $X2=2.72 $Y2=0.805
r45 1 9 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.265 $X2=1.3 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_404_53# 1 2 7 11 13
c21 13 0 1.21702e-19 $X=2.16 $Y=0.35
r22 13 16 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=0.35
+ $X2=2.16 $Y2=0.455
r23 9 11 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.66 $Y=0.435
+ $X2=3.66 $Y2=0.73
r24 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0.35
+ $X2=2.16 $Y2=0.35
r25 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=3.66 $Y2=0.435
r26 7 8 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=2.325 $Y2=0.35
r27 2 11 182 $w=1.7e-07 $l=2.92916e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.56 $X2=3.66 $Y2=0.73
r28 1 16 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.265 $X2=2.16 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__EDFXBP_1%A_1789_141# 1 2 12 14 15
r35 14 15 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.455 $Y=0.96
+ $X2=11.29 $Y2=0.96
r36 12 15 132.765 $w=1.68e-07 $l=2.035e-06 $layer=LI1_cond $X=9.255 $Y=0.98
+ $X2=11.29 $Y2=0.98
r37 10 12 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.09 $Y=0.915
+ $X2=9.255 $Y2=0.915
r38 2 14 182 $w=1.7e-07 $l=3.58852e-07 $layer=licon1_NDIFF $count=1 $X=11.205
+ $Y=0.705 $X2=11.455 $Y2=0.96
r39 1 10 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.945
+ $Y=0.705 $X2=9.09 $Y2=0.915
.ends

