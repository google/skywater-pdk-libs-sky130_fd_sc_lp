* File: sky130_fd_sc_lp__nand2_2.pex.spice
* Created: Wed Sep  2 10:02:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_2%B 3 7 11 15 17 18 26
c40 11 0 8.47484e-20 $X=0.905 $Y=0.745
r41 24 26 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.635 $Y=1.51
+ $X2=0.905 $Y2=1.51
r42 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=1.51 $X2=0.635 $Y2=1.51
r43 21 24 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.475 $Y=1.51
+ $X2=0.635 $Y2=1.51
r44 18 25 2.92411 $w=3.33e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.582
+ $X2=0.635 $Y2=1.582
r45 17 25 13.5885 $w=3.33e-07 $l=3.95e-07 $layer=LI1_cond $X=0.24 $Y=1.582
+ $X2=0.635 $Y2=1.582
r46 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=1.51
r47 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=2.465
r48 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=1.51
r49 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.905 $Y=1.345 $X2=0.905
+ $Y2=0.745
r50 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=1.51
r51 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=2.465
r52 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=1.51
r53 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.475 $Y=1.345 $X2=0.475
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_2%A 3 7 11 15 17 18 26
r47 24 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.55 $Y=1.51
+ $X2=1.765 $Y2=1.51
r48 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.51 $X2=1.55 $Y2=1.51
r49 21 24 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.55 $Y2=1.51
r50 18 25 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=1.68 $Y=1.582
+ $X2=1.55 $Y2=1.582
r51 17 25 12.0404 $w=3.33e-07 $l=3.5e-07 $layer=LI1_cond $X=1.2 $Y=1.582
+ $X2=1.55 $Y2=1.582
r52 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.675
+ $X2=1.765 $Y2=1.51
r53 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.765 $Y=1.675
+ $X2=1.765 $Y2=2.465
r54 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.51
r55 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.765 $Y=1.345 $X2=1.765
+ $Y2=0.745
r56 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.675
+ $X2=1.335 $Y2=1.51
r57 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.335 $Y=1.675
+ $X2=1.335 $Y2=2.465
r58 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.345
+ $X2=1.335 $Y2=1.51
r59 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.335 $Y=1.345 $X2=1.335
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_2%VPWR 1 2 3 10 12 18 20 22 24 26 31 40 44
r38 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.12 $Y2=3.33
r43 32 34 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 31 43 4.49945 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.107 $Y2=3.33
r45 31 34 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 27 37 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r49 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.12 $Y2=3.33
r51 26 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 24 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 20 43 3.26672 $w=3.3e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=2.107 $Y2=3.33
r56 20 22 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=1.98 $Y2=2.4
r57 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=3.33
r58 16 18 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=2.4
r59 12 15 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=0.26 $Y=2.09
+ $X2=0.26 $Y2=2.95
r60 10 37 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r61 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r62 3 22 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.4
r63 2 18 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.4
r64 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r65 1 12 400 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.09
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_2%Y 1 2 3 10 12 14 18 22 24 26 27 31 34
c43 27 0 8.47484e-20 $X=1.715 $Y=1.16
r44 33 34 9.47977 $w=3.08e-07 $l=2.55e-07 $layer=LI1_cond $X=2.155 $Y=1.92
+ $X2=2.155 $Y2=1.665
r45 32 34 15.6137 $w=3.08e-07 $l=4.2e-07 $layer=LI1_cond $X=2.155 $Y=1.245
+ $X2=2.155 $Y2=1.665
r46 26 32 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2 $Y=1.16
+ $X2=2.155 $Y2=1.245
r47 26 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2 $Y=1.16 $X2=1.715
+ $Y2=1.16
r48 25 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.645 $Y=2.005
+ $X2=1.55 $Y2=2.005
r49 24 33 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2 $Y=2.005
+ $X2=2.155 $Y2=1.92
r50 24 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2 $Y=2.005
+ $X2=1.645 $Y2=2.005
r51 20 31 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=2.09
+ $X2=1.55 $Y2=2.005
r52 20 22 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=1.55 $Y=2.09 $X2=1.55
+ $Y2=2.91
r53 16 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.55 $Y=1.075
+ $X2=1.715 $Y2=1.16
r54 16 18 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.55 $Y=1.075
+ $X2=1.55 $Y2=0.69
r55 15 29 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.785 $Y=2.005
+ $X2=0.69 $Y2=2.005
r56 14 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.455 $Y=2.005
+ $X2=1.55 $Y2=2.005
r57 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.455 $Y=2.005
+ $X2=0.785 $Y2=2.005
r58 10 29 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.09 $X2=0.69
+ $Y2=2.005
r59 10 12 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=0.69 $Y=2.09 $X2=0.69
+ $Y2=2.91
r60 3 31 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.085
r61 3 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.91
r62 2 29 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.085
r63 2 12 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.91
r64 1 18 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.325 $X2=1.55 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_2%A_27_65# 1 2 3 12 14 15 20 21 24
r34 22 24 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.06 $Y=0.435
+ $X2=2.06 $Y2=0.47
r35 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.895 $Y=0.35
+ $X2=2.06 $Y2=0.435
r36 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=0.35
+ $X2=1.205 $Y2=0.35
r37 17 19 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.12 $Y=1.075
+ $X2=1.12 $Y2=0.47
r38 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.435
+ $X2=1.205 $Y2=0.35
r39 16 19 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.12 $Y=0.435
+ $X2=1.12 $Y2=0.47
r40 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=1.12 $Y2=1.075
r41 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=0.355 $Y2=1.16
r42 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.355 $Y2=1.16
r43 10 12 26.8165 $w=2.58e-07 $l=6.05e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.225 $Y2=0.47
r44 3 24 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.325 $X2=2.06 $Y2=0.47
r45 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.325 $X2=1.12 $Y2=0.47
r46 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.325 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_2%VGND 1 6 8 10 20 21 24
r26 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r27 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r28 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r29 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r30 15 17 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r31 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r32 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r34 10 12 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r35 8 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r36 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r37 8 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r39 4 6 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.45
r40 1 6 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.325 $X2=0.69 $Y2=0.45
.ends

