* File: sky130_fd_sc_lp__o311a_m.pxi.spice
* Created: Wed Sep  2 10:23:26 2020
* 
x_PM_SKY130_FD_SC_LP__O311A_M%A1 N_A1_c_85_n N_A1_M1004_g N_A1_M1003_g
+ N_A1_c_86_n N_A1_c_87_n N_A1_c_88_n A1 A1 A1 N_A1_c_90_n N_A1_c_91_n
+ PM_SKY130_FD_SC_LP__O311A_M%A1
x_PM_SKY130_FD_SC_LP__O311A_M%A2 N_A2_M1000_g N_A2_M1008_g N_A2_c_130_n
+ N_A2_c_134_n A2 A2 A2 A2 N_A2_c_132_n PM_SKY130_FD_SC_LP__O311A_M%A2
x_PM_SKY130_FD_SC_LP__O311A_M%A_93_153# N_A_93_153#_M1001_d N_A_93_153#_M1005_d
+ N_A_93_153#_M1006_d N_A_93_153#_M1009_g N_A_93_153#_c_177_n
+ N_A_93_153#_c_178_n N_A_93_153#_c_172_n N_A_93_153#_M1011_g
+ N_A_93_153#_c_173_n N_A_93_153#_c_179_n N_A_93_153#_c_180_n
+ N_A_93_153#_c_181_n N_A_93_153#_c_182_n N_A_93_153#_c_174_n
+ N_A_93_153#_c_184_n N_A_93_153#_c_185_n N_A_93_153#_c_186_n
+ N_A_93_153#_c_175_n PM_SKY130_FD_SC_LP__O311A_M%A_93_153#
x_PM_SKY130_FD_SC_LP__O311A_M%A3 N_A3_M1010_g N_A3_M1005_g N_A3_c_259_n
+ N_A3_c_260_n A3 N_A3_c_261_n N_A3_c_270_n PM_SKY130_FD_SC_LP__O311A_M%A3
x_PM_SKY130_FD_SC_LP__O311A_M%B1 N_B1_M1007_g N_B1_M1002_g N_B1_c_299_n
+ N_B1_c_300_n B1 B1 N_B1_c_302_n PM_SKY130_FD_SC_LP__O311A_M%B1
x_PM_SKY130_FD_SC_LP__O311A_M%C1 N_C1_M1006_g N_C1_M1001_g N_C1_c_347_n
+ N_C1_c_348_n N_C1_c_340_n N_C1_c_341_n N_C1_c_342_n N_C1_c_343_n C1 C1 C1 C1
+ C1 N_C1_c_345_n PM_SKY130_FD_SC_LP__O311A_M%C1
x_PM_SKY130_FD_SC_LP__O311A_M%X N_X_M1011_s N_X_M1009_s N_X_c_384_n N_X_c_382_n
+ X N_X_c_383_n PM_SKY130_FD_SC_LP__O311A_M%X
x_PM_SKY130_FD_SC_LP__O311A_M%VPWR N_VPWR_M1009_d N_VPWR_M1002_d N_VPWR_c_395_n
+ N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n VPWR N_VPWR_c_399_n
+ N_VPWR_c_400_n N_VPWR_c_394_n N_VPWR_c_402_n PM_SKY130_FD_SC_LP__O311A_M%VPWR
x_PM_SKY130_FD_SC_LP__O311A_M%VGND N_VGND_M1011_d N_VGND_M1008_d N_VGND_c_432_n
+ N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n
+ VGND N_VGND_c_438_n N_VGND_c_439_n PM_SKY130_FD_SC_LP__O311A_M%VGND
x_PM_SKY130_FD_SC_LP__O311A_M%A_250_47# N_A_250_47#_M1003_d N_A_250_47#_M1010_d
+ N_A_250_47#_c_484_n N_A_250_47#_c_485_n N_A_250_47#_c_486_n
+ N_A_250_47#_c_487_n PM_SKY130_FD_SC_LP__O311A_M%A_250_47#
cc_1 VNB N_A1_c_85_n 0.0207087f $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.648
cc_2 VNB N_A1_c_86_n 4.61658e-19 $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.825
cc_3 VNB N_A1_c_87_n 0.016567f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.765
cc_4 VNB N_A1_c_88_n 0.011794f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.915
cc_5 VNB A1 0.00949929f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_A1_c_90_n 0.0174962f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.32
cc_7 VNB N_A1_c_91_n 0.0140651f $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.155
cc_8 VNB N_A2_M1008_g 0.036142f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.195
cc_9 VNB N_A2_c_130_n 0.0206593f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.445
cc_10 VNB A2 0.0047141f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.765
cc_11 VNB N_A2_c_132_n 0.0152781f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.32
cc_12 VNB N_A_93_153#_M1009_g 0.0405774f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.765
cc_13 VNB N_A_93_153#_c_172_n 0.0198002f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_14 VNB N_A_93_153#_c_173_n 0.0230527f $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.32
cc_15 VNB N_A_93_153#_c_174_n 0.0194525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_93_153#_c_175_n 0.00889548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_M1010_g 0.0289451f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=0.915
cc_18 VNB N_A3_c_259_n 0.0230706f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.445
cc_19 VNB N_A3_c_260_n 0.0105938f $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.825
cc_20 VNB N_A3_c_261_n 0.0162642f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_21 VNB N_B1_M1007_g 0.0203367f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=0.915
cc_22 VNB N_B1_M1002_g 0.0113666f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.195
cc_23 VNB N_B1_c_299_n 0.0267952f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.445
cc_24 VNB N_B1_c_300_n 0.0183353f $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.825
cc_25 VNB B1 0.00309577f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.765
cc_26 VNB N_B1_c_302_n 0.0185745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_M1001_g 0.0259894f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.195
cc_28 VNB N_C1_c_340_n 0.038267f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.445
cc_29 VNB N_C1_c_341_n 0.00922157f $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.825
cc_30 VNB N_C1_c_342_n 0.00865485f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.915
cc_31 VNB N_C1_c_343_n 0.0250694f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB C1 0.00902883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_C1_c_345_n 0.0380985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_382_n 0.0485966f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.445
cc_35 VNB N_X_c_383_n 0.025359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_394_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_432_n 0.00439692f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.765
cc_38 VNB N_VGND_c_433_n 0.00439692f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.765
cc_39 VNB N_VGND_c_434_n 0.0254545f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_40 VNB N_VGND_c_435_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_41 VNB N_VGND_c_436_n 0.0181538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_437_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_438_n 0.0582479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_439_n 0.216947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_250_47#_c_484_n 0.00134021f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.765
cc_46 VNB N_A_250_47#_c_485_n 0.0159695f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.445
cc_47 VNB N_A_250_47#_c_486_n 0.00816928f $X=-0.19 $Y=-0.245 $X2=1.032 $Y2=1.825
cc_48 VNB N_A_250_47#_c_487_n 0.00135575f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_49 VPB N_A1_M1004_g 0.0201727f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.195
cc_50 VPB N_A1_c_86_n 0.0170631f $X=-0.19 $Y=1.655 $X2=1.032 $Y2=1.825
cc_51 VPB A1 0.0106612f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_52 VPB N_A2_M1000_g 0.0183135f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=0.915
cc_53 VPB N_A2_c_134_n 0.0153433f $X=-0.19 $Y=1.655 $X2=1.032 $Y2=1.825
cc_54 VPB A2 0.0050833f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=0.765
cc_55 VPB N_A_93_153#_M1009_g 0.0666029f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=0.765
cc_56 VPB N_A_93_153#_c_177_n 0.116916f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=0.915
cc_57 VPB N_A_93_153#_c_178_n 0.0151908f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_58 VPB N_A_93_153#_c_179_n 0.0159813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_93_153#_c_180_n 0.0205491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_93_153#_c_181_n 0.00595212f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.295
cc_61 VPB N_A_93_153#_c_182_n 8.99879e-19 $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.665
cc_62 VPB N_A_93_153#_c_174_n 0.00110107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_93_153#_c_184_n 0.00571625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_93_153#_c_185_n 0.0484718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_93_153#_c_186_n 7.66045e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A3_M1005_g 0.0296283f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.195
cc_67 VPB N_A3_c_260_n 0.0062455f $X=-0.19 $Y=1.655 $X2=1.032 $Y2=1.825
cc_68 VPB N_B1_M1002_g 0.0312685f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.195
cc_69 VPB N_C1_M1006_g 0.0225214f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=0.915
cc_70 VPB N_C1_c_347_n 0.0381041f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.765
cc_71 VPB N_C1_c_348_n 0.0121157f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.445
cc_72 VPB N_C1_c_342_n 0.00217846f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=0.915
cc_73 VPB C1 0.0418955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_X_c_384_n 0.01667f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.445
cc_75 VPB N_X_c_382_n 0.0150781f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.445
cc_76 VPB N_VPWR_c_395_n 0.0221855f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.765
cc_77 VPB N_VPWR_c_396_n 0.0376404f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=0.765
cc_78 VPB N_VPWR_c_397_n 0.0530312f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_79 VPB N_VPWR_c_398_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_80 VPB N_VPWR_c_399_n 0.0206615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_400_n 0.0322151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_394_n 0.0953775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_402_n 0.00583335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 N_A1_M1004_g N_A2_M1000_g 0.0211272f $X=1.135 $Y=2.195 $X2=0 $Y2=0
cc_85 N_A1_c_87_n N_A2_M1008_g 0.0201838f $X=1.155 $Y=0.765 $X2=0 $Y2=0
cc_86 A1 N_A2_M1008_g 0.00131349f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A1_c_91_n N_A2_M1008_g 0.00944226f $X=1.032 $Y=1.155 $X2=0 $Y2=0
cc_88 N_A1_c_85_n N_A2_c_130_n 0.0211272f $X=1.032 $Y=1.648 $X2=0 $Y2=0
cc_89 N_A1_c_86_n N_A2_c_134_n 0.0211272f $X=1.032 $Y=1.825 $X2=0 $Y2=0
cc_90 A1 A2 0.0257053f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_91 N_A1_c_90_n A2 0.00512836f $X=1.02 $Y=1.32 $X2=0 $Y2=0
cc_92 A1 N_A2_c_132_n 0.00207835f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A1_c_90_n N_A2_c_132_n 0.0211272f $X=1.02 $Y=1.32 $X2=0 $Y2=0
cc_94 N_A1_M1004_g N_A_93_153#_M1009_g 0.0135543f $X=1.135 $Y=2.195 $X2=0 $Y2=0
cc_95 A1 N_A_93_153#_M1009_g 0.00894002f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A1_c_90_n N_A_93_153#_M1009_g 0.0328755f $X=1.02 $Y=1.32 $X2=0 $Y2=0
cc_97 N_A1_c_91_n N_A_93_153#_M1009_g 0.00303797f $X=1.032 $Y=1.155 $X2=0 $Y2=0
cc_98 N_A1_M1004_g N_A_93_153#_c_177_n 0.00545354f $X=1.135 $Y=2.195 $X2=0 $Y2=0
cc_99 N_A1_c_87_n N_A_93_153#_c_172_n 0.0148797f $X=1.155 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A1_c_88_n N_A_93_153#_c_173_n 0.00853762f $X=1.155 $Y=0.915 $X2=0 $Y2=0
cc_101 A1 N_A_93_153#_c_173_n 0.0127004f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 A1 N_X_c_382_n 0.0525244f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A1_M1004_g N_VPWR_c_395_n 0.00557486f $X=1.135 $Y=2.195 $X2=0 $Y2=0
cc_104 N_A1_c_86_n N_VPWR_c_395_n 4.62461e-19 $X=1.032 $Y=1.825 $X2=0 $Y2=0
cc_105 A1 N_VPWR_c_395_n 0.0148499f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_106 N_A1_M1004_g N_VPWR_c_394_n 8.51218e-19 $X=1.135 $Y=2.195 $X2=0 $Y2=0
cc_107 N_A1_c_87_n N_VGND_c_432_n 0.00156327f $X=1.155 $Y=0.765 $X2=0 $Y2=0
cc_108 A1 N_VGND_c_432_n 0.0103694f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_109 N_A1_c_90_n N_VGND_c_432_n 7.50744e-19 $X=1.02 $Y=1.32 $X2=0 $Y2=0
cc_110 N_A1_c_87_n N_VGND_c_436_n 0.00585385f $X=1.155 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A1_c_88_n N_VGND_c_436_n 6.8925e-19 $X=1.155 $Y=0.915 $X2=0 $Y2=0
cc_112 N_A1_c_87_n N_VGND_c_439_n 0.0106127f $X=1.155 $Y=0.765 $X2=0 $Y2=0
cc_113 N_A1_c_88_n N_VGND_c_439_n 9.8095e-19 $X=1.155 $Y=0.915 $X2=0 $Y2=0
cc_114 A1 N_VGND_c_439_n 0.00965934f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_115 N_A1_c_87_n N_A_250_47#_c_484_n 0.00170671f $X=1.155 $Y=0.765 $X2=0 $Y2=0
cc_116 N_A1_c_87_n N_A_250_47#_c_486_n 0.00423251f $X=1.155 $Y=0.765 $X2=0 $Y2=0
cc_117 A1 N_A_250_47#_c_486_n 0.0045521f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_118 N_A2_M1000_g N_A_93_153#_c_177_n 0.00506318f $X=1.495 $Y=2.195 $X2=0
+ $Y2=0
cc_119 A2 N_A_93_153#_c_177_n 0.00620473f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_120 A2 N_A_93_153#_c_179_n 0.0150504f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_121 A2 N_A_93_153#_c_181_n 0.0084375f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A2_M1008_g N_A3_M1010_g 0.0336068f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A2_M1000_g N_A3_M1005_g 0.0185022f $X=1.495 $Y=2.195 $X2=0 $Y2=0
cc_124 N_A2_c_130_n N_A3_c_259_n 0.0137835f $X=1.585 $Y=1.66 $X2=0 $Y2=0
cc_125 N_A2_c_134_n N_A3_c_260_n 0.0137835f $X=1.585 $Y=1.825 $X2=0 $Y2=0
cc_126 A2 N_A3_c_261_n 0.0126456f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A2_c_132_n N_A3_c_261_n 0.0137835f $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_128 N_A2_M1008_g N_A3_c_270_n 4.98669e-19 $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_129 A2 N_A3_c_270_n 0.0301073f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_132_n N_A3_c_270_n 5.24566e-19 $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_131 A2 N_VPWR_c_395_n 0.00988924f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A2_M1000_g N_VPWR_c_394_n 8.51218e-19 $X=1.495 $Y=2.195 $X2=0 $Y2=0
cc_133 A2 N_VPWR_c_394_n 0.00910345f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 A2 A_314_397# 0.00533621f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_135 N_A2_M1008_g N_VGND_c_433_n 0.00156327f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A2_M1008_g N_VGND_c_436_n 0.00437852f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A2_M1008_g N_VGND_c_439_n 0.00604796f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A2_M1008_g N_A_250_47#_c_484_n 9.4709e-19 $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A2_M1008_g N_A_250_47#_c_485_n 0.0122928f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_140 A2 N_A_250_47#_c_485_n 0.0147462f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A2_c_132_n N_A_250_47#_c_485_n 8.41944e-19 $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_142 N_A2_c_132_n N_A_250_47#_c_486_n 0.00319817f $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_143 N_A_93_153#_c_177_n N_A3_M1005_g 0.00234561f $X=2.025 $Y=3.03 $X2=0 $Y2=0
cc_144 N_A_93_153#_c_179_n N_A3_M1005_g 0.00327966f $X=2.25 $Y=2.13 $X2=0 $Y2=0
cc_145 N_A_93_153#_c_181_n N_A3_M1005_g 0.00238561f $X=2.355 $Y=1.85 $X2=0 $Y2=0
cc_146 N_A_93_153#_c_184_n N_A3_M1005_g 5.45931e-19 $X=2.19 $Y=2.94 $X2=0 $Y2=0
cc_147 N_A_93_153#_c_185_n N_A3_M1005_g 0.00535823f $X=2.19 $Y=2.94 $X2=0 $Y2=0
cc_148 N_A_93_153#_c_181_n N_A3_c_260_n 0.0042802f $X=2.355 $Y=1.85 $X2=0 $Y2=0
cc_149 N_A_93_153#_c_181_n N_A3_c_270_n 0.0120415f $X=2.355 $Y=1.85 $X2=0 $Y2=0
cc_150 N_A_93_153#_c_174_n N_B1_M1007_g 8.82604e-19 $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_93_153#_c_175_n N_B1_M1007_g 0.00101523f $X=3.33 $Y=0.51 $X2=0 $Y2=0
cc_152 N_A_93_153#_c_179_n N_B1_M1002_g 0.00800308f $X=2.25 $Y=2.13 $X2=0 $Y2=0
cc_153 N_A_93_153#_c_180_n N_B1_M1002_g 0.0171998f $X=3.115 $Y=1.85 $X2=0 $Y2=0
cc_154 N_A_93_153#_c_174_n N_B1_M1002_g 0.00614379f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_93_153#_c_174_n N_B1_c_299_n 0.00547185f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_93_153#_c_180_n N_B1_c_300_n 0.00351131f $X=3.115 $Y=1.85 $X2=0 $Y2=0
cc_157 N_A_93_153#_c_180_n B1 0.00968604f $X=3.115 $Y=1.85 $X2=0 $Y2=0
cc_158 N_A_93_153#_c_174_n B1 0.0255335f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_93_153#_c_174_n N_B1_c_302_n 6.17235e-19 $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_93_153#_c_180_n N_C1_M1006_g 0.00985216f $X=3.115 $Y=1.85 $X2=0 $Y2=0
cc_161 N_A_93_153#_c_182_n N_C1_M1006_g 0.00196872f $X=3.22 $Y=2.11 $X2=0 $Y2=0
cc_162 N_A_93_153#_c_174_n N_C1_M1001_g 0.0078528f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_93_153#_c_175_n N_C1_M1001_g 0.00562804f $X=3.33 $Y=0.51 $X2=0 $Y2=0
cc_164 N_A_93_153#_c_180_n N_C1_c_347_n 0.00202586f $X=3.115 $Y=1.85 $X2=0 $Y2=0
cc_165 N_A_93_153#_c_174_n N_C1_c_347_n 0.00632001f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_93_153#_c_186_n N_C1_c_347_n 0.00784395f $X=3.21 $Y=1.85 $X2=0 $Y2=0
cc_167 N_A_93_153#_c_180_n N_C1_c_348_n 0.00790877f $X=3.115 $Y=1.85 $X2=0 $Y2=0
cc_168 N_A_93_153#_c_174_n N_C1_c_340_n 0.00825463f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_93_153#_c_175_n N_C1_c_340_n 0.00709503f $X=3.33 $Y=0.51 $X2=0 $Y2=0
cc_170 N_A_93_153#_c_174_n N_C1_c_341_n 0.00365314f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_93_153#_c_182_n C1 0.0246682f $X=3.22 $Y=2.11 $X2=0 $Y2=0
cc_172 N_A_93_153#_c_174_n C1 0.0631787f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A_93_153#_c_186_n C1 0.0131818f $X=3.21 $Y=1.85 $X2=0 $Y2=0
cc_174 N_A_93_153#_c_175_n C1 5.60103e-19 $X=3.33 $Y=0.51 $X2=0 $Y2=0
cc_175 N_A_93_153#_c_174_n N_C1_c_345_n 0.00752707f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A_93_153#_M1009_g N_X_c_384_n 7.93141e-19 $X=0.54 $Y=2.195 $X2=0 $Y2=0
cc_177 N_A_93_153#_c_172_n N_X_c_382_n 0.00297004f $X=0.745 $Y=0.765 $X2=0 $Y2=0
cc_178 N_A_93_153#_c_173_n N_X_c_382_n 0.02994f $X=0.745 $Y=0.84 $X2=0 $Y2=0
cc_179 N_A_93_153#_c_173_n N_X_c_383_n 0.00793786f $X=0.745 $Y=0.84 $X2=0 $Y2=0
cc_180 N_A_93_153#_M1009_g N_VPWR_c_395_n 0.0397693f $X=0.54 $Y=2.195 $X2=0
+ $Y2=0
cc_181 N_A_93_153#_c_177_n N_VPWR_c_395_n 0.0244106f $X=2.025 $Y=3.03 $X2=0
+ $Y2=0
cc_182 N_A_93_153#_c_178_n N_VPWR_c_395_n 0.00656411f $X=0.615 $Y=3.03 $X2=0
+ $Y2=0
cc_183 N_A_93_153#_c_179_n N_VPWR_c_396_n 0.028417f $X=2.25 $Y=2.13 $X2=0 $Y2=0
cc_184 N_A_93_153#_c_180_n N_VPWR_c_396_n 0.0146902f $X=3.115 $Y=1.85 $X2=0
+ $Y2=0
cc_185 N_A_93_153#_c_184_n N_VPWR_c_396_n 0.00785069f $X=2.19 $Y=2.94 $X2=0
+ $Y2=0
cc_186 N_A_93_153#_c_185_n N_VPWR_c_396_n 0.00533051f $X=2.19 $Y=2.94 $X2=0
+ $Y2=0
cc_187 N_A_93_153#_c_177_n N_VPWR_c_397_n 0.0374824f $X=2.025 $Y=3.03 $X2=0
+ $Y2=0
cc_188 N_A_93_153#_c_184_n N_VPWR_c_397_n 0.0152941f $X=2.19 $Y=2.94 $X2=0 $Y2=0
cc_189 N_A_93_153#_c_178_n N_VPWR_c_399_n 0.00393414f $X=0.615 $Y=3.03 $X2=0
+ $Y2=0
cc_190 N_A_93_153#_c_177_n N_VPWR_c_394_n 0.047087f $X=2.025 $Y=3.03 $X2=0 $Y2=0
cc_191 N_A_93_153#_c_178_n N_VPWR_c_394_n 0.00783176f $X=0.615 $Y=3.03 $X2=0
+ $Y2=0
cc_192 N_A_93_153#_c_184_n N_VPWR_c_394_n 0.0104794f $X=2.19 $Y=2.94 $X2=0 $Y2=0
cc_193 N_A_93_153#_c_185_n N_VPWR_c_394_n 0.00782252f $X=2.19 $Y=2.94 $X2=0
+ $Y2=0
cc_194 N_A_93_153#_c_172_n N_VGND_c_432_n 0.00288714f $X=0.745 $Y=0.765 $X2=0
+ $Y2=0
cc_195 N_A_93_153#_c_172_n N_VGND_c_434_n 0.00585385f $X=0.745 $Y=0.765 $X2=0
+ $Y2=0
cc_196 N_A_93_153#_c_173_n N_VGND_c_434_n 6.59122e-19 $X=0.745 $Y=0.84 $X2=0
+ $Y2=0
cc_197 N_A_93_153#_c_175_n N_VGND_c_438_n 0.0109093f $X=3.33 $Y=0.51 $X2=0 $Y2=0
cc_198 N_A_93_153#_M1001_d N_VGND_c_439_n 0.00236056f $X=3.19 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_A_93_153#_c_172_n N_VGND_c_439_n 0.00749616f $X=0.745 $Y=0.765 $X2=0
+ $Y2=0
cc_200 N_A_93_153#_c_173_n N_VGND_c_439_n 7.45101e-19 $X=0.745 $Y=0.84 $X2=0
+ $Y2=0
cc_201 N_A_93_153#_c_175_n N_VGND_c_439_n 0.0120475f $X=3.33 $Y=0.51 $X2=0 $Y2=0
cc_202 N_A3_M1010_g N_B1_M1007_g 0.0203727f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_203 N_A3_M1005_g N_B1_M1002_g 0.0173544f $X=2.035 $Y=2.195 $X2=0 $Y2=0
cc_204 N_A3_c_260_n N_B1_M1002_g 0.0142171f $X=2.125 $Y=1.665 $X2=0 $Y2=0
cc_205 N_A3_c_261_n N_B1_c_299_n 0.0142171f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A3_c_270_n N_B1_c_299_n 0.00220614f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A3_c_259_n N_B1_c_300_n 0.0142171f $X=2.125 $Y=1.5 $X2=0 $Y2=0
cc_208 N_A3_M1010_g B1 6.11235e-19 $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A3_c_261_n B1 0.00175571f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A3_c_270_n B1 0.0196812f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A3_M1005_g N_VPWR_c_394_n 3.66166e-19 $X=2.035 $Y=2.195 $X2=0 $Y2=0
cc_212 N_A3_M1010_g N_VGND_c_433_n 0.00288714f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A3_M1010_g N_VGND_c_438_n 0.00437852f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A3_M1010_g N_VGND_c_439_n 0.00630876f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A3_M1010_g N_A_250_47#_c_485_n 0.0121375f $X=2.035 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A3_c_261_n N_A_250_47#_c_485_n 0.00523522f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A3_c_270_n N_A_250_47#_c_485_n 0.0250028f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A3_M1010_g N_A_250_47#_c_487_n 0.00103339f $X=2.035 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_B1_M1007_g N_C1_M1001_g 0.0234307f $X=2.575 $Y=0.445 $X2=0 $Y2=0
cc_220 B1 N_C1_M1001_g 6.87366e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_221 N_B1_c_302_n N_C1_M1001_g 0.00630511f $X=2.665 $Y=0.96 $X2=0 $Y2=0
cc_222 N_B1_M1002_g N_C1_c_348_n 0.0217326f $X=2.575 $Y=2.195 $X2=0 $Y2=0
cc_223 N_B1_c_299_n N_C1_c_341_n 0.00630511f $X=2.665 $Y=1.3 $X2=0 $Y2=0
cc_224 N_B1_c_300_n N_C1_c_343_n 0.00266238f $X=2.665 $Y=1.465 $X2=0 $Y2=0
cc_225 N_B1_c_299_n N_C1_c_345_n 0.00266238f $X=2.665 $Y=1.3 $X2=0 $Y2=0
cc_226 N_B1_M1002_g N_VPWR_c_396_n 0.00127738f $X=2.575 $Y=2.195 $X2=0 $Y2=0
cc_227 N_B1_M1002_g N_VPWR_c_394_n 0.00393927f $X=2.575 $Y=2.195 $X2=0 $Y2=0
cc_228 N_B1_M1007_g N_VGND_c_438_n 0.00585385f $X=2.575 $Y=0.445 $X2=0 $Y2=0
cc_229 N_B1_M1007_g N_VGND_c_439_n 0.00869802f $X=2.575 $Y=0.445 $X2=0 $Y2=0
cc_230 B1 N_VGND_c_439_n 0.0067861f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_231 N_B1_c_302_n N_VGND_c_439_n 0.00210244f $X=2.665 $Y=0.96 $X2=0 $Y2=0
cc_232 N_B1_M1007_g N_A_250_47#_c_485_n 0.00294484f $X=2.575 $Y=0.445 $X2=0
+ $Y2=0
cc_233 B1 N_A_250_47#_c_485_n 0.006715f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_234 N_B1_M1007_g N_A_250_47#_c_487_n 0.00849146f $X=2.575 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_C1_M1006_g N_VPWR_c_396_n 0.00225549f $X=3.005 $Y=2.195 $X2=0 $Y2=0
cc_236 C1 N_VPWR_c_396_n 0.0048366f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_237 N_C1_M1006_g N_VPWR_c_394_n 0.00393927f $X=3.005 $Y=2.195 $X2=0 $Y2=0
cc_238 C1 N_VPWR_c_394_n 0.00780715f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_239 N_C1_M1001_g N_VGND_c_438_n 0.00512735f $X=3.115 $Y=0.445 $X2=0 $Y2=0
cc_240 N_C1_M1001_g N_VGND_c_439_n 0.0104507f $X=3.115 $Y=0.445 $X2=0 $Y2=0
cc_241 N_C1_c_340_n N_VGND_c_439_n 0.00128969f $X=3.405 $Y=0.915 $X2=0 $Y2=0
cc_242 C1 N_VGND_c_439_n 0.00672977f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_243 N_X_c_383_n N_VGND_c_434_n 0.0213142f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_244 N_X_M1011_s N_VGND_c_439_n 0.00242809f $X=0.405 $Y=0.235 $X2=0 $Y2=0
cc_245 N_X_c_383_n N_VGND_c_439_n 0.0175272f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_246 N_VGND_c_439_n N_A_250_47#_M1003_d 0.00373063f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_247 N_VGND_c_439_n N_A_250_47#_M1010_d 0.00914164f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_436_n N_A_250_47#_c_484_n 0.008231f $X=1.715 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_439_n N_A_250_47#_c_484_n 0.00765087f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_c_433_n N_A_250_47#_c_485_n 0.0139569f $X=1.82 $Y=0.38 $X2=0 $Y2=0
cc_251 N_VGND_c_436_n N_A_250_47#_c_485_n 0.00305343f $X=1.715 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_438_n N_A_250_47#_c_485_n 0.00305343f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_439_n N_A_250_47#_c_485_n 0.0109462f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_438_n N_A_250_47#_c_487_n 0.00778424f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_439_n N_A_250_47#_c_487_n 0.00691521f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_439_n A_530_47# 0.0120089f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
