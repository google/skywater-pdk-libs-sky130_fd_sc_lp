* File: sky130_fd_sc_lp__a211oi_lp.pex.spice
* Created: Fri Aug 28 09:48:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211OI_LP%C1 1 3 7 10 12 14 16 17 18 19 20 21 22 23
+ 30 32
r49 30 32 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.345
+ $X2=0.72 $Y2=1.18
r50 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=2.405
+ $X2=0.74 $Y2=2.775
r51 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=2.035
+ $X2=0.74 $Y2=2.405
r52 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.665
+ $X2=0.74 $Y2=2.035
r53 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.295
+ $X2=0.74 $Y2=1.665
r54 19 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.74
+ $Y=1.345 $X2=0.74 $Y2=1.345
r55 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.97 $Y=0.78 $X2=0.97
+ $Y2=0.495
r56 13 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.685 $Y=0.855
+ $X2=0.61 $Y2=0.855
r57 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.895 $Y=0.855
+ $X2=0.97 $Y2=0.78
r58 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.895 $Y=0.855
+ $X2=0.685 $Y2=0.855
r59 10 18 172.675 $w=2.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.78 $Y=2.545
+ $X2=0.78 $Y2=1.85
r60 7 18 34.9505 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=1.85
r61 6 30 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=0.72 $Y=1.365 $X2=0.72
+ $Y2=1.345
r62 6 7 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=0.72 $Y=1.365 $X2=0.72
+ $Y2=1.665
r63 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.61 $Y=0.93 $X2=0.61
+ $Y2=0.855
r64 4 32 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.61 $Y=0.93 $X2=0.61
+ $Y2=1.18
r65 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.61 $Y=0.78 $X2=0.61
+ $Y2=0.855
r66 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.61 $Y=0.78 $X2=0.61
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_LP%B1 3 5 7 10 12 14 16 17 18 19 20 22 29
r55 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.31
+ $Y=1.335 $X2=1.31 $Y2=1.335
r56 22 30 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.505
+ $X2=1.31 $Y2=1.505
r57 20 30 1.96371 $w=6.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=1.505
+ $X2=1.31 $Y2=1.505
r58 17 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.31 $Y=1.675
+ $X2=1.31 $Y2=1.335
r59 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.675
+ $X2=1.31 $Y2=1.84
r60 16 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.17
+ $X2=1.31 $Y2=1.335
r61 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.76 $Y=0.78 $X2=1.76
+ $Y2=0.495
r62 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.475 $Y=0.855
+ $X2=1.4 $Y2=0.855
r63 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.685 $Y=0.855
+ $X2=1.76 $Y2=0.78
r64 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.685 $Y=0.855
+ $X2=1.475 $Y2=0.855
r65 8 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.4 $Y=0.93 $X2=1.4
+ $Y2=0.855
r66 8 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.4 $Y=0.93 $X2=1.4
+ $Y2=1.17
r67 5 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.4 $Y=0.78 $X2=1.4
+ $Y2=0.855
r68 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.4 $Y=0.78 $X2=1.4
+ $Y2=0.495
r69 3 18 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.27 $Y=2.545
+ $X2=1.27 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_LP%A1 3 7 9 10 14
r37 14 17 63.9614 $w=5.9e-07 $l=5.05e-07 $layer=POLY_cond $X=2.01 $Y=1.335
+ $X2=2.01 $Y2=1.84
r38 14 16 49.19 $w=5.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.335
+ $X2=2.01 $Y2=1.17
r39 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=1.295
+ $X2=2.14 $Y2=1.665
r40 9 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.14
+ $Y=1.335 $X2=2.14 $Y2=1.335
r41 7 16 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.19 $Y=0.495
+ $X2=2.19 $Y2=1.17
r42 3 17 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.84 $Y=2.545
+ $X2=1.84 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_LP%A2 3 7 11 12 13 15 22
r30 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.71
+ $Y=1.275 $X2=2.71 $Y2=1.275
r31 15 23 7.31929 $w=6.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.12 $Y=1.445
+ $X2=2.71 $Y2=1.445
r32 13 23 1.24963 $w=6.68e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=1.445 $X2=2.71
+ $Y2=1.445
r33 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.71 $Y=1.615
+ $X2=2.71 $Y2=1.275
r34 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.615
+ $X2=2.71 $Y2=1.78
r35 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.11
+ $X2=2.71 $Y2=1.275
r36 7 12 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.67 $Y=2.545
+ $X2=2.67 $Y2=1.78
r37 3 10 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.62 $Y=0.495
+ $X2=2.62 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_LP%Y 1 2 3 10 14 16 17 18 19 20 21 22 33
r43 22 52 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=2.775
+ $X2=0.26 $Y2=2.9
r44 21 22 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r45 21 46 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.19
r46 20 46 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.26 $Y=2.035
+ $X2=0.26 $Y2=2.19
r47 19 20 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r48 18 19 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r49 17 31 2.71818 $w=3.52e-07 $l=8.5e-08 $layer=LI1_cond $X=0.342 $Y=0.905
+ $X2=0.342 $Y2=0.82
r50 17 37 2.71818 $w=3.52e-07 $l=1.19143e-07 $layer=LI1_cond $X=0.342 $Y=0.905
+ $X2=0.26 $Y2=0.99
r51 17 18 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=1 $X2=0.26
+ $Y2=1.295
r52 17 37 0.426831 $w=2.68e-07 $l=1e-08 $layer=LI1_cond $X=0.26 $Y=1 $X2=0.26
+ $Y2=0.99
r53 16 31 7.02063 $w=4.33e-07 $l=2.65e-07 $layer=LI1_cond $X=0.342 $Y=0.555
+ $X2=0.342 $Y2=0.82
r54 16 33 1.58958 $w=4.33e-07 $l=6e-08 $layer=LI1_cond $X=0.342 $Y=0.555
+ $X2=0.342 $Y2=0.495
r55 12 14 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.975 $Y=0.82
+ $X2=1.975 $Y2=0.495
r56 11 17 4.06059 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.56 $Y=0.905
+ $X2=0.342 $Y2=0.905
r57 10 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.81 $Y=0.905
+ $X2=1.975 $Y2=0.82
r58 10 11 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.81 $Y=0.905
+ $X2=0.56 $Y2=0.905
r59 3 52 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.045 $X2=0.31 $Y2=2.9
r60 3 46 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.045 $X2=0.31 $Y2=2.19
r61 2 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.835
+ $Y=0.285 $X2=1.975 $Y2=0.495
r62 1 33 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.25
+ $Y=0.285 $X2=0.395 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_LP%A_279_409# 1 2 11 13 14 19
r27 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.935 $Y=2.19
+ $X2=2.935 $Y2=2.9
r28 13 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.77 $Y=2.105
+ $X2=2.935 $Y2=2.19
r29 13 14 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.77 $Y=2.105
+ $X2=1.74 $Y2=2.105
r30 9 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.575 $Y=2.19
+ $X2=1.74 $Y2=2.105
r31 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.575 $Y=2.19
+ $X2=1.575 $Y2=2.9
r32 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=2.045 $X2=2.935 $Y2=2.9
r33 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=2.045 $X2=2.935 $Y2=2.19
r34 1 11 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=2.045 $X2=1.575 $Y2=2.9
r35 1 9 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=2.045 $X2=1.575 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_LP%VPWR 1 6 8 10 20 21 24
r29 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=3.33
+ $X2=2.105 $Y2=3.33
r33 18 20 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.27 $Y=3.33
+ $X2=3.12 $Y2=3.33
r34 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.105 $Y2=3.33
r37 10 16 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=3.245
+ $X2=2.105 $Y2=3.33
r42 4 6 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.105 $Y=3.245
+ $X2=2.105 $Y2=2.535
r43 1 6 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=2.045 $X2=2.105 $Y2=2.535
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_LP%VGND 1 2 9 13 16 17 18 20 33 34 37
r41 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r44 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r45 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r46 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.185
+ $Y2=0
r47 25 27 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.68
+ $Y2=0
r48 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r49 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.185
+ $Y2=0
r51 20 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.72
+ $Y2=0
r52 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r53 18 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 18 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 16 30 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.64
+ $Y2=0
r56 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.835
+ $Y2=0
r57 15 33 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.12
+ $Y2=0
r58 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=0 $X2=2.835
+ $Y2=0
r59 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.835 $Y=0.085
+ $X2=2.835 $Y2=0
r60 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.835 $Y=0.085
+ $X2=2.835 $Y2=0.495
r61 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r62 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.45
r63 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.285 $X2=2.835 $Y2=0.495
r64 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.285 $X2=1.185 $Y2=0.45
.ends

