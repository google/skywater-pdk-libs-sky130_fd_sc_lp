* File: sky130_fd_sc_lp__o21bai_2.pex.spice
* Created: Fri Aug 28 11:06:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BAI_2%B1_N 2 5 6 7 10 12 13 17 19
c29 2 0 5.82284e-20 $X=0.362 $Y=1.36
r30 17 19 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.005
+ $X2=0.362 $Y2=0.84
r31 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.34
+ $Y=1.005 $X2=0.34 $Y2=1.005
r32 13 18 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.005
r33 12 18 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.005
r34 8 10 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.84 $Y=1.51 $X2=0.84
+ $Y2=2.045
r35 6 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.765 $Y=1.435
+ $X2=0.84 $Y2=1.51
r36 6 7 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.765 $Y=1.435
+ $X2=0.55 $Y2=1.435
r37 5 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.52
+ $X2=0.475 $Y2=0.84
r38 2 7 33.9315 $w=1.5e-07 $l=2.2236e-07 $layer=POLY_cond $X=0.362 $Y=1.36
+ $X2=0.55 $Y2=1.435
r39 1 17 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.362 $Y=1.027
+ $X2=0.362 $Y2=1.005
r40 1 2 49.3865 $w=3.75e-07 $l=3.33e-07 $layer=POLY_cond $X=0.362 $Y=1.027
+ $X2=0.362 $Y2=1.36
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%A_100_367# 1 2 7 9 12 14 16 18 21 23 26 32
+ 36 37 39 43
c69 39 0 5.82284e-20 $X=0.725 $Y=1.48
r70 42 43 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.505 $Y=1.44
+ $X2=1.58 $Y2=1.44
r71 36 37 11.8331 $w=3.33e-07 $l=2.9e-07 $layer=LI1_cond $X=0.627 $Y=2.045
+ $X2=0.627 $Y2=1.755
r72 33 42 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.29 $Y=1.44
+ $X2=1.505 $Y2=1.44
r73 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.29
+ $Y=1.44 $X2=1.29 $Y2=1.44
r74 30 39 1.04409 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=0.855 $Y=1.48
+ $X2=0.725 $Y2=1.48
r75 30 32 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=0.855 $Y=1.48
+ $X2=1.29 $Y2=1.48
r76 28 39 5.53409 $w=2.3e-07 $l=1.39194e-07 $layer=LI1_cond $X=0.695 $Y=1.605
+ $X2=0.725 $Y2=1.48
r77 28 37 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=0.695 $Y=1.605
+ $X2=0.695 $Y2=1.755
r78 24 39 5.53409 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.725 $Y=1.355
+ $X2=0.725 $Y2=1.48
r79 24 26 37.0112 $w=2.58e-07 $l=8.35e-07 $layer=LI1_cond $X=0.725 $Y=1.355
+ $X2=0.725 $Y2=0.52
r80 19 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.425
+ $X2=1.935 $Y2=1.35
r81 19 21 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.935 $Y=1.425
+ $X2=1.935 $Y2=2.465
r82 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.275
+ $X2=1.935 $Y2=1.35
r83 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.935 $Y=1.275
+ $X2=1.935 $Y2=0.745
r84 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.935 $Y2=1.35
r85 14 43 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.58 $Y2=1.35
r86 10 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.605
+ $X2=1.505 $Y2=1.44
r87 10 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.505 $Y=1.605
+ $X2=1.505 $Y2=2.465
r88 7 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.275
+ $X2=1.505 $Y2=1.44
r89 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.505 $Y=1.275
+ $X2=1.505 $Y2=0.745
r90 2 36 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.5
+ $Y=1.835 $X2=0.625 $Y2=2.045
r91 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.31 $X2=0.69 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%A1 3 7 11 15 18 19 21 22 24 26 27 35 36 45
c83 18 0 5.32484e-20 $X=3.605 $Y=1.92
c84 7 0 8.53043e-20 $X=2.445 $Y=2.465
r85 43 52 6.90441 $w=2e-07 $l=2.83e-07 $layer=LI1_cond $X=2.58 $Y=2.02 $X2=2.297
+ $Y2=2.02
r86 43 45 3.32727 $w=1.98e-07 $l=6e-08 $layer=LI1_cond $X=2.58 $Y=2.02 $X2=2.64
+ $Y2=2.02
r87 36 52 10.7965 $w=5.63e-07 $l=5.1e-07 $layer=LI1_cond $X=2.297 $Y=1.51
+ $X2=2.297 $Y2=2.02
r88 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.51
+ $X2=2.415 $Y2=1.675
r89 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.51
+ $X2=2.415 $Y2=1.345
r90 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.51 $X2=2.415 $Y2=1.51
r91 26 27 14.7198 $w=3.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.12 $Y=2.02
+ $X2=3.515 $Y2=2.02
r92 24 52 0.317543 $w=5.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.297 $Y=2.035
+ $X2=2.297 $Y2=2.02
r93 24 26 25.9527 $w=1.98e-07 $l=4.68e-07 $layer=LI1_cond $X=2.652 $Y=2.02
+ $X2=3.12 $Y2=2.02
r94 24 45 0.665455 $w=1.98e-07 $l=1.2e-08 $layer=LI1_cond $X=2.652 $Y=2.02
+ $X2=2.64 $Y2=2.02
r95 22 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.51
+ $X2=3.825 $Y2=1.675
r96 22 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.51
+ $X2=3.825 $Y2=1.345
r97 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.51 $X2=3.825 $Y2=1.51
r98 19 21 6.80989 $w=2.18e-07 $l=1.3e-07 $layer=LI1_cond $X=3.695 $Y=1.535
+ $X2=3.825 $Y2=1.535
r99 18 27 3.60057 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=3.605 $Y=1.92 $X2=3.605
+ $Y2=2.02
r100 17 19 6.90553 $w=2.2e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.605 $Y=1.645
+ $X2=3.695 $Y2=1.535
r101 17 18 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.605 $Y=1.645
+ $X2=3.605 $Y2=1.92
r102 15 41 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.735 $Y=2.465
+ $X2=3.735 $Y2=1.675
r103 11 40 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.735 $Y=0.745
+ $X2=3.735 $Y2=1.345
r104 7 38 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.445 $Y=2.465
+ $X2=2.445 $Y2=1.675
r105 3 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.365 $Y=0.745
+ $X2=2.365 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%A2 3 7 11 15 17 24
c52 17 0 8.53043e-20 $X=3.12 $Y=1.665
r53 22 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.965 $Y=1.51
+ $X2=3.305 $Y2=1.51
r54 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.51 $X2=2.965 $Y2=1.51
r55 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.875 $Y=1.51
+ $X2=2.965 $Y2=1.51
r56 17 23 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=3.12 $Y=1.587
+ $X2=2.965 $Y2=1.587
r57 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.675
+ $X2=3.305 $Y2=1.51
r58 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.305 $Y=1.675
+ $X2=3.305 $Y2=2.465
r59 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.345
+ $X2=3.305 $Y2=1.51
r60 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.305 $Y=1.345 $X2=3.305
+ $Y2=0.745
r61 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.675
+ $X2=2.875 $Y2=1.51
r62 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.875 $Y=1.675
+ $X2=2.875 $Y2=2.465
r63 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.345
+ $X2=2.875 $Y2=1.51
r64 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.875 $Y=1.345 $X2=2.875
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%VPWR 1 2 3 12 18 20 22 26 28 33 38 47 50 54
r52 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r57 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 39 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 39 41 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 38 53 3.91666 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=4.092 $Y2=3.33
r62 38 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 34 47 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.195 $Y2=3.33
r66 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 33 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.16 $Y2=3.33
r68 33 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 28 47 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.195 $Y2=3.33
r72 28 30 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 26 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 26 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 22 25 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=3.99 $Y=1.98
+ $X2=3.99 $Y2=2.95
r77 20 53 3.2265 $w=2.5e-07 $l=1.38109e-07 $layer=LI1_cond $X=3.99 $Y=3.245
+ $X2=4.092 $Y2=3.33
r78 20 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.99 $Y=3.245
+ $X2=3.99 $Y2=2.95
r79 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=3.33
r80 16 18 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=2.915
r81 12 15 11.5708 $w=4.58e-07 $l=4.45e-07 $layer=LI1_cond $X=1.195 $Y=1.98
+ $X2=1.195 $Y2=2.425
r82 10 47 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=3.33
r83 10 15 21.3214 $w=4.58e-07 $l=8.2e-07 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=2.425
r84 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.835 $X2=3.95 $Y2=2.95
r85 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.835 $X2=3.95 $Y2=1.98
r86 2 18 600 $w=1.7e-07 $l=1.15256e-06 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.16 $Y2=2.915
r87 1 15 300 $w=1.7e-07 $l=7.54553e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=1.835 $X2=1.29 $Y2=2.425
r88 1 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.915
+ $Y=1.835 $X2=1.055 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%Y 1 2 3 12 16 22 24 25 26 27 28
r42 28 31 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=2.455
+ $X2=1.72 $Y2=2.29
r43 27 31 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=1.72 $Y=1.98
+ $X2=1.72 $Y2=2.29
r44 25 27 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=1.72 $Y=1.94 $X2=1.72
+ $Y2=1.98
r45 25 26 5.95733 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.72 $Y=1.94
+ $X2=1.72 $Y2=1.815
r46 24 26 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=1.735 $Y=1.145
+ $X2=1.735 $Y2=1.815
r47 20 28 0.225187 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.845 $Y=2.455
+ $X2=1.72 $Y2=2.455
r48 20 22 43.4785 $w=3.28e-07 $l=1.245e-06 $layer=LI1_cond $X=1.845 $Y=2.455
+ $X2=3.09 $Y2=2.455
r49 14 28 6.67463 $w=2.4e-07 $l=1.69926e-07 $layer=LI1_cond $X=1.71 $Y=2.62
+ $X2=1.72 $Y2=2.455
r50 14 16 14.5308 $w=2.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.71 $Y=2.62
+ $X2=1.71 $Y2=2.91
r51 10 24 6.50529 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=0.98
+ $X2=1.72 $Y2=1.145
r52 10 12 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.72 $Y=0.98 $X2=1.72
+ $Y2=0.68
r53 3 22 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=1.835 $X2=3.09 $Y2=2.455
r54 2 28 600 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.835 $X2=1.72 $Y2=2.445
r55 2 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.835 $X2=1.72 $Y2=1.98
r56 2 16 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.835 $X2=1.72 $Y2=2.91
r57 1 12 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=1.58
+ $Y=0.325 $X2=1.72 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%A_504_367# 1 2 7 13
r20 11 13 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=3.52 $Y=2.8
+ $X2=3.52 $Y2=2.375
r21 7 11 6.89002 $w=2.75e-07 $l=2.23226e-07 $layer=LI1_cond $X=3.355 $Y=2.937
+ $X2=3.52 $Y2=2.8
r22 7 9 29.1254 $w=2.73e-07 $l=6.95e-07 $layer=LI1_cond $X=3.355 $Y=2.937
+ $X2=2.66 $Y2=2.937
r23 2 13 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=3.38
+ $Y=1.835 $X2=3.52 $Y2=2.375
r24 1 9 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=1.835 $X2=2.66 $Y2=2.915
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%VGND 1 2 3 10 12 16 20 22 24 32 39 40 46 49
r52 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r53 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r56 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.52
+ $Y2=0
r58 37 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=4.08
+ $Y2=0
r59 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r60 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r61 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r62 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.765 $Y=0 $X2=2.6
+ $Y2=0
r63 33 35 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.765 $Y=0 $X2=3.12
+ $Y2=0
r64 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.52
+ $Y2=0
r65 32 35 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.12
+ $Y2=0
r66 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r67 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r68 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 25 43 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r70 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r71 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=0 $X2=2.6
+ $Y2=0
r72 24 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=0 $X2=2.16
+ $Y2=0
r73 22 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r74 22 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.72
+ $Y2=0
r75 22 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r76 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.52 $Y2=0
r77 18 20 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.52 $Y2=0.45
r78 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=0.085 $X2=2.6
+ $Y2=0
r79 14 16 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.6 $Y=0.085
+ $X2=2.6 $Y2=0.45
r80 10 43 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r81 10 12 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.535
r82 3 20 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.38
+ $Y=0.325 $X2=3.52 $Y2=0.45
r83 2 16 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=2.44
+ $Y=0.325 $X2=2.6 $Y2=0.45
r84 1 12 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.31 $X2=0.26 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_2%A_233_65# 1 2 3 4 15 17 18 23 24 27 29 33
+ 35
r62 31 33 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=3.995 $Y=1.085
+ $X2=3.995 $Y2=0.47
r63 30 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.185 $Y=1.17
+ $X2=3.06 $Y2=1.17
r64 29 31 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.855 $Y=1.17
+ $X2=3.995 $Y2=1.085
r65 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.855 $Y=1.17
+ $X2=3.185 $Y2=1.17
r66 25 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=1.085
+ $X2=3.06 $Y2=1.17
r67 25 27 28.3501 $w=2.48e-07 $l=6.15e-07 $layer=LI1_cond $X=3.06 $Y=1.085
+ $X2=3.06 $Y2=0.47
r68 23 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.935 $Y=1.17
+ $X2=3.06 $Y2=1.17
r69 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.935 $Y=1.17
+ $X2=2.265 $Y2=1.17
r70 20 24 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.165 $Y=1.085
+ $X2=2.265 $Y2=1.17
r71 20 22 34.1045 $w=1.98e-07 $l=6.15e-07 $layer=LI1_cond $X=2.165 $Y=1.085
+ $X2=2.165 $Y2=0.47
r72 19 22 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=2.165 $Y=0.425
+ $X2=2.165 $Y2=0.47
r73 17 19 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.065 $Y=0.34
+ $X2=2.165 $Y2=0.425
r74 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.065 $Y=0.34
+ $X2=1.375 $Y2=0.34
r75 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.25 $Y=0.425
+ $X2=1.375 $Y2=0.34
r76 13 15 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=1.25 $Y=0.425
+ $X2=1.25 $Y2=0.47
r77 4 33 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=3.81
+ $Y=0.325 $X2=3.97 $Y2=0.47
r78 3 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.95
+ $Y=0.325 $X2=3.09 $Y2=0.47
r79 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.325 $X2=2.15 $Y2=0.47
r80 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.165
+ $Y=0.325 $X2=1.29 $Y2=0.47
.ends

