# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o41ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o41ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.210000 10.475000 1.525000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.745000 1.345000 8.435000 1.525000 ;
        RECT 6.745000 1.525000 7.335000 1.750000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845000 1.345000 6.575000 1.750000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 1.355000 4.255000 1.525000 ;
        RECT 2.985000 1.525000 3.685000 1.760000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.375000 2.815000 1.760000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.881600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.930000 4.350000 2.100000 ;
        RECT 0.990000 2.100000 1.180000 3.075000 ;
        RECT 1.385000 0.595000 1.610000 1.015000 ;
        RECT 1.385000 1.015000 4.675000 1.185000 ;
        RECT 1.860000 2.100000 2.040000 3.075000 ;
        RECT 2.280000 0.595000 2.470000 1.015000 ;
        RECT 3.160000 2.100000 3.490000 2.725000 ;
        RECT 4.020000 1.705000 4.675000 1.875000 ;
        RECT 4.020000 1.875000 4.350000 1.930000 ;
        RECT 4.020000 2.100000 4.350000 2.725000 ;
        RECT 4.425000 1.185000 4.675000 1.705000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.490000  1.930000  0.820000 3.245000 ;
      RECT  0.920000  0.255000  2.970000 0.425000 ;
      RECT  0.920000  0.425000  1.215000 1.095000 ;
      RECT  1.350000  2.270000  1.680000 3.245000 ;
      RECT  1.780000  0.425000  2.110000 0.845000 ;
      RECT  2.210000  2.270000  2.540000 3.245000 ;
      RECT  2.640000  0.425000  2.970000 0.675000 ;
      RECT  2.640000  0.675000  5.015000 0.845000 ;
      RECT  2.730000  2.270000  2.990000 2.895000 ;
      RECT  2.730000  2.895000  4.710000 3.075000 ;
      RECT  3.150000  0.085000  3.480000 0.505000 ;
      RECT  3.660000  0.255000  3.990000 0.675000 ;
      RECT  3.660000  2.270000  3.850000 2.895000 ;
      RECT  4.170000  0.085000  4.500000 0.505000 ;
      RECT  4.520000  2.045000  6.500000 2.225000 ;
      RECT  4.520000  2.225000  4.710000 2.895000 ;
      RECT  4.680000  0.255000  5.015000 0.675000 ;
      RECT  4.845000  0.845000  5.015000 1.005000 ;
      RECT  4.845000  1.005000 10.390000 1.040000 ;
      RECT  4.845000  1.040000  8.585000 1.175000 ;
      RECT  4.845000  1.920000  6.500000 2.045000 ;
      RECT  4.880000  2.395000  5.210000 2.855000 ;
      RECT  4.880000  2.855000  8.310000 3.075000 ;
      RECT  5.185000  0.085000  5.515000 0.835000 ;
      RECT  5.380000  2.225000  5.570000 2.685000 ;
      RECT  5.690000  0.255000  5.880000 1.005000 ;
      RECT  5.740000  2.395000  6.070000 2.855000 ;
      RECT  6.050000  0.085000  6.380000 0.835000 ;
      RECT  6.240000  2.225000  6.500000 2.685000 ;
      RECT  6.550000  0.255000  6.740000 1.005000 ;
      RECT  6.690000  1.920000  7.880000 2.100000 ;
      RECT  6.690000  2.100000  6.950000 2.685000 ;
      RECT  6.910000  0.085000  7.240000 0.835000 ;
      RECT  7.120000  2.270000  7.450000 2.735000 ;
      RECT  7.120000  2.735000  8.310000 2.855000 ;
      RECT  7.410000  0.255000  7.670000 1.005000 ;
      RECT  7.620000  1.695000 10.460000 1.875000 ;
      RECT  7.620000  1.875000  7.880000 1.920000 ;
      RECT  7.620000  2.100000  7.880000 2.490000 ;
      RECT  7.840000  0.085000  8.170000 0.835000 ;
      RECT  8.050000  2.045000  8.310000 2.735000 ;
      RECT  8.340000  0.255000  8.625000 0.870000 ;
      RECT  8.340000  0.870000 10.390000 1.005000 ;
      RECT  8.480000  1.875000  8.670000 3.075000 ;
      RECT  8.795000  0.085000  9.070000 0.700000 ;
      RECT  8.840000  2.045000  9.170000 3.245000 ;
      RECT  9.240000  0.255000  9.490000 0.870000 ;
      RECT  9.340000  1.875000  9.530000 3.075000 ;
      RECT  9.660000  0.085000  9.940000 0.700000 ;
      RECT  9.700000  2.045000 10.030000 3.245000 ;
      RECT 10.110000  0.255000 10.390000 0.870000 ;
      RECT 10.200000  1.875000 10.460000 3.075000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__o41ai_4
END LIBRARY
