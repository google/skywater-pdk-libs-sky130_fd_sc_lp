* File: sky130_fd_sc_lp__a32o_0.pxi.spice
* Created: Fri Aug 28 10:00:47 2020
* 
x_PM_SKY130_FD_SC_LP__A32O_0%A_80_21# N_A_80_21#_M1007_d N_A_80_21#_M1001_d
+ N_A_80_21#_M1005_g N_A_80_21#_M1009_g N_A_80_21#_c_79_n N_A_80_21#_c_88_n
+ N_A_80_21#_c_80_n N_A_80_21#_c_81_n N_A_80_21#_c_82_n N_A_80_21#_c_83_n
+ N_A_80_21#_c_113_p N_A_80_21#_c_84_n N_A_80_21#_c_125_p N_A_80_21#_c_85_n
+ N_A_80_21#_c_90_n PM_SKY130_FD_SC_LP__A32O_0%A_80_21#
x_PM_SKY130_FD_SC_LP__A32O_0%A3 N_A3_c_177_n N_A3_M1006_g N_A3_M1004_g
+ N_A3_c_180_n A3 A3 N_A3_c_182_n N_A3_c_200_n PM_SKY130_FD_SC_LP__A32O_0%A3
x_PM_SKY130_FD_SC_LP__A32O_0%A2 N_A2_M1000_g N_A2_M1003_g N_A2_c_229_n
+ N_A2_c_230_n A2 N_A2_c_231_n N_A2_c_232_n PM_SKY130_FD_SC_LP__A32O_0%A2
x_PM_SKY130_FD_SC_LP__A32O_0%A1 N_A1_M1007_g N_A1_M1011_g N_A1_c_282_n
+ N_A1_c_283_n A1 A1 N_A1_c_285_n PM_SKY130_FD_SC_LP__A32O_0%A1
x_PM_SKY130_FD_SC_LP__A32O_0%B1 N_B1_M1010_g N_B1_M1001_g N_B1_c_323_n
+ N_B1_c_324_n B1 B1 N_B1_c_326_n PM_SKY130_FD_SC_LP__A32O_0%B1
x_PM_SKY130_FD_SC_LP__A32O_0%B2 N_B2_c_361_n N_B2_M1008_g N_B2_M1002_g
+ N_B2_c_363_n B2 B2 B2 N_B2_c_365_n PM_SKY130_FD_SC_LP__A32O_0%B2
x_PM_SKY130_FD_SC_LP__A32O_0%X N_X_M1005_s N_X_M1009_s X X X X X X X N_X_c_397_n
+ X N_X_c_399_n PM_SKY130_FD_SC_LP__A32O_0%X
x_PM_SKY130_FD_SC_LP__A32O_0%VPWR N_VPWR_M1009_d N_VPWR_M1003_d N_VPWR_c_414_n
+ N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n VPWR N_VPWR_c_418_n
+ N_VPWR_c_419_n N_VPWR_c_413_n N_VPWR_c_421_n PM_SKY130_FD_SC_LP__A32O_0%VPWR
x_PM_SKY130_FD_SC_LP__A32O_0%A_269_429# N_A_269_429#_M1006_d
+ N_A_269_429#_M1011_d N_A_269_429#_M1008_d N_A_269_429#_c_454_n
+ N_A_269_429#_c_455_n N_A_269_429#_c_456_n N_A_269_429#_c_457_n
+ N_A_269_429#_c_458_n N_A_269_429#_c_459_n N_A_269_429#_c_460_n
+ PM_SKY130_FD_SC_LP__A32O_0%A_269_429#
x_PM_SKY130_FD_SC_LP__A32O_0%VGND N_VGND_M1005_d N_VGND_M1002_d N_VGND_c_498_n
+ N_VGND_c_499_n VGND N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ N_VGND_c_503_n PM_SKY130_FD_SC_LP__A32O_0%VGND
cc_1 VNB N_A_80_21#_M1005_g 0.0508614f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_80_21#_c_79_n 0.015303f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.845
cc_3 VNB N_A_80_21#_c_80_n 0.00400194f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.45
cc_4 VNB N_A_80_21#_c_81_n 0.0195569f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.45
cc_5 VNB N_A_80_21#_c_82_n 0.0232395f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.76
cc_6 VNB N_A_80_21#_c_83_n 0.00190857f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.76
cc_7 VNB N_A_80_21#_c_84_n 0.00295776f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=0.445
cc_8 VNB N_A_80_21#_c_85_n 0.0122225f $X=-0.19 $Y=-0.245 $X2=3.037 $Y2=1.785
cc_9 VNB N_A3_c_177_n 0.0208983f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.145
cc_10 VNB N_A3_M1006_g 0.00226735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_M1004_g 0.0281203f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_12 VNB N_A3_c_180_n 0.0235099f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.462
cc_13 VNB A3 9.8895e-19 $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.995
cc_14 VNB N_A3_c_182_n 0.0240474f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.845
cc_15 VNB N_A2_M1000_g 0.0286921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_229_n 0.0209127f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.462
cc_17 VNB N_A2_c_230_n 0.00907649f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.845
cc_18 VNB N_A2_c_231_n 0.0151177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_232_n 0.00444844f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.845
cc_20 VNB N_A1_M1007_g 0.0216368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_M1011_g 0.00816805f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.285
cc_22 VNB N_A1_c_282_n 0.0208947f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.462
cc_23 VNB N_A1_c_283_n 0.0153831f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.845
cc_24 VNB A1 0.0101603f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.995
cc_25 VNB N_A1_c_285_n 0.0158444f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.995
cc_26 VNB N_B1_M1010_g 0.0224914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_M1001_g 0.0090804f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.285
cc_28 VNB N_B1_c_323_n 0.0225239f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.462
cc_29 VNB N_B1_c_324_n 0.0164289f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.845
cc_30 VNB B1 0.0105768f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.995
cc_31 VNB N_B1_c_326_n 0.0151969f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.995
cc_32 VNB N_B2_c_361_n 0.0221374f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=0.235
cc_33 VNB N_B2_M1002_g 0.0325755f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.285
cc_34 VNB N_B2_c_363_n 0.0321505f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.465
cc_35 VNB B2 0.0373643f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.845
cc_36 VNB N_B2_c_365_n 0.0287002f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.76
cc_37 VNB X 0.0534056f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.285
cc_38 VNB N_X_c_397_n 0.0129546f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=0.61
cc_39 VNB N_VPWR_c_413_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=2.27
cc_40 VNB N_VGND_c_498_n 0.0122476f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.285
cc_41 VNB N_VGND_c_499_n 0.0192289f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_42 VNB N_VGND_c_500_n 0.0518269f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.995
cc_43 VNB N_VGND_c_501_n 0.0151978f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=0.445
cc_44 VNB N_VGND_c_502_n 0.0137467f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=2.27
cc_45 VNB N_VGND_c_503_n 0.208255f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=1.785
cc_46 VPB N_A_80_21#_M1009_g 0.0207482f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.465
cc_47 VPB N_A_80_21#_c_79_n 0.0161944f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.845
cc_48 VPB N_A_80_21#_c_88_n 0.0330914f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.995
cc_49 VPB N_A_80_21#_c_85_n 0.00216222f $X=-0.19 $Y=1.655 $X2=3.037 $Y2=1.785
cc_50 VPB N_A_80_21#_c_90_n 0.00519098f $X=-0.19 $Y=1.655 $X2=3.037 $Y2=1.955
cc_51 VPB N_A3_M1006_g 0.0381593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB A3 0.00517849f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.995
cc_53 VPB N_A2_M1003_g 0.0372701f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.285
cc_54 VPB N_A2_c_230_n 0.00674491f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.845
cc_55 VPB N_A2_c_232_n 7.98174e-19 $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.845
cc_56 VPB N_A1_M1011_g 0.0370037f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.285
cc_57 VPB N_B1_M1001_g 0.0362532f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.285
cc_58 VPB N_B2_c_361_n 0.0346852f $X=-0.19 $Y=1.655 $X2=2.275 $Y2=0.235
cc_59 VPB N_B2_M1008_g 0.0296736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB B2 0.0141072f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.845
cc_61 VPB X 0.024818f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.285
cc_62 VPB N_X_c_399_n 0.0593182f $X=-0.19 $Y=1.655 $X2=3.037 $Y2=1.955
cc_63 VPB N_VPWR_c_414_n 0.0187723f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_64 VPB N_VPWR_c_415_n 0.0123137f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.995
cc_65 VPB N_VPWR_c_416_n 0.0268012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_417_n 0.00535984f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.845
cc_67 VPB N_VPWR_c_418_n 0.0191784f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.76
cc_68 VPB N_VPWR_c_419_n 0.0431088f $X=-0.19 $Y=1.655 $X2=2.985 $Y2=1.955
cc_69 VPB N_VPWR_c_413_n 0.0838826f $X=-0.19 $Y=1.655 $X2=2.985 $Y2=2.27
cc_70 VPB N_VPWR_c_421_n 0.00632158f $X=-0.19 $Y=1.655 $X2=3.17 $Y2=0.61
cc_71 VPB N_A_269_429#_c_454_n 0.00657963f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.845
cc_72 VPB N_A_269_429#_c_455_n 0.0194059f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.465
cc_73 VPB N_A_269_429#_c_456_n 0.00935967f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.465
cc_74 VPB N_A_269_429#_c_457_n 0.0018231f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.845
cc_75 VPB N_A_269_429#_c_458_n 0.02034f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.45
cc_76 VPB N_A_269_429#_c_459_n 0.00352015f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.45
cc_77 VPB N_A_269_429#_c_460_n 0.0338423f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.76
cc_78 N_A_80_21#_c_80_n N_A3_c_177_n 9.69718e-19 $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_81_n N_A3_c_177_n 0.00996263f $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_79_n N_A3_M1006_g 0.00541352f $X=0.657 $Y=1.845 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_88_n N_A3_M1006_g 0.0191485f $X=0.657 $Y=1.995 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_80_n N_A3_M1006_g 6.7053e-19 $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_83 N_A_80_21#_M1005_g N_A3_M1004_g 0.00616886f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_80_n N_A3_M1004_g 0.0015996f $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_82_n N_A3_M1004_g 0.0135205f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_84_n N_A3_M1004_g 0.00540729f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_79_n N_A3_c_180_n 0.00996263f $X=0.657 $Y=1.845 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_79_n A3 0.0022238f $X=0.657 $Y=1.845 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_80_n A3 0.0203488f $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_90 N_A_80_21#_M1005_g N_A3_c_182_n 0.00875552f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_80_n N_A3_c_182_n 0.00409386f $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_82_n N_A3_c_182_n 0.00743976f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_93 N_A_80_21#_M1005_g N_A3_c_200_n 2.58994e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_80_n N_A3_c_200_n 0.0347552f $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_81_n N_A3_c_200_n 9.41415e-19 $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_82_n N_A3_c_200_n 0.030142f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_82_n N_A2_M1000_g 3.04808e-19 $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_84_n N_A2_M1000_g 0.0173012f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_82_n N_A2_c_231_n 2.59669e-19 $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_113_p N_A2_c_231_n 0.0018885f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_84_n N_A2_c_231_n 0.00276163f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_82_n N_A2_c_232_n 0.00625348f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_84_n N_A2_c_232_n 0.0214428f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_113_p N_A1_M1007_g 0.0116485f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_84_n N_A1_M1007_g 0.00279606f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_90_n N_A1_M1011_g 7.45437e-19 $X=3.037 $Y=1.955 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_113_p A1 0.0240205f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_84_n A1 0.00533757f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_113_p N_A1_c_285_n 0.00383504f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_113_p N_B1_M1010_g 0.0180668f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_85_n N_B1_M1010_g 0.00342368f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_125_p N_B1_M1001_g 0.0103348f $X=2.985 $Y=2.27 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_85_n N_B1_M1001_g 0.00670863f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_90_n N_B1_M1001_g 0.00488833f $X=3.037 $Y=1.955 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_90_n N_B1_c_324_n 0.00398454f $X=3.037 $Y=1.955 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_113_p B1 0.0253192f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_85_n B1 0.0555174f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_90_n B1 0.00566449f $X=3.037 $Y=1.955 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_113_p N_B1_c_326_n 0.00382778f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_85_n N_B1_c_326_n 0.00671634f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_85_n N_B2_c_361_n 0.0040358f $X=3.037 $Y=1.785 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_80_21#_c_90_n N_B2_c_361_n 0.00591762f $X=3.037 $Y=1.955 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_80_21#_c_125_p N_B2_M1008_g 0.0162559f $X=2.985 $Y=2.27 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_90_n N_B2_M1008_g 0.00890089f $X=3.037 $Y=1.955 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_113_p N_B2_M1002_g 0.00956751f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_85_n N_B2_M1002_g 0.0119297f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_85_n N_B2_c_363_n 0.00447877f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_85_n B2 0.0797417f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_85_n N_B2_c_365_n 0.0039597f $X=3.037 $Y=1.785 $X2=0 $Y2=0
cc_130 N_A_80_21#_M1005_g X 0.0358513f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_80_21#_M1009_g X 0.00351437f $X=0.84 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_80_n X 0.0840532f $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_83_n X 0.0139714f $X=0.755 $Y=0.76 $X2=0 $Y2=0
cc_134 N_A_80_21#_M1009_g N_X_c_399_n 0.00364023f $X=0.84 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_88_n N_X_c_399_n 0.0124202f $X=0.657 $Y=1.995 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_80_n N_X_c_399_n 0.0221091f $X=0.59 $Y=1.45 $X2=0 $Y2=0
cc_137 N_A_80_21#_M1009_g N_VPWR_c_414_n 0.00120184f $X=0.84 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_A_80_21#_M1009_g N_VPWR_c_416_n 0.00460069f $X=0.84 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_M1009_g N_VPWR_c_413_n 0.00492109f $X=0.84 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_c_90_n N_A_269_429#_c_455_n 0.0144432f $X=3.037 $Y=1.955 $X2=0
+ $Y2=0
cc_141 N_A_80_21#_c_125_p N_A_269_429#_c_457_n 0.0302852f $X=2.985 $Y=2.27 $X2=0
+ $Y2=0
cc_142 N_A_80_21#_c_125_p N_A_269_429#_c_458_n 0.0205458f $X=2.985 $Y=2.27 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_c_125_p N_A_269_429#_c_460_n 0.0232845f $X=2.985 $Y=2.27 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_c_113_p N_VGND_c_499_n 0.0266531f $X=3.085 $Y=0.445 $X2=0
+ $Y2=0
cc_145 N_A_80_21#_c_82_n N_VGND_c_500_n 0.00554648f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_113_p N_VGND_c_500_n 0.071924f $X=3.085 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_84_n N_VGND_c_500_n 0.0121945f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_80_21#_M1005_g N_VGND_c_501_n 0.00466457f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_149 N_A_80_21#_c_83_n N_VGND_c_501_n 3.18906e-19 $X=0.755 $Y=0.76 $X2=0 $Y2=0
cc_150 N_A_80_21#_M1005_g N_VGND_c_502_n 0.00958841f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_151 N_A_80_21#_c_82_n N_VGND_c_502_n 0.0358737f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_152 N_A_80_21#_c_83_n N_VGND_c_502_n 0.0171546f $X=0.755 $Y=0.76 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_84_n N_VGND_c_502_n 0.0104834f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_154 N_A_80_21#_M1007_d N_VGND_c_503_n 0.00316088f $X=2.275 $Y=0.235 $X2=0
+ $Y2=0
cc_155 N_A_80_21#_M1005_g N_VGND_c_503_n 0.00848288f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_156 N_A_80_21#_c_82_n N_VGND_c_503_n 0.0109888f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_157 N_A_80_21#_c_83_n N_VGND_c_503_n 0.00156811f $X=0.755 $Y=0.76 $X2=0 $Y2=0
cc_158 N_A_80_21#_c_113_p N_VGND_c_503_n 0.0513675f $X=3.085 $Y=0.445 $X2=0
+ $Y2=0
cc_159 N_A_80_21#_c_84_n N_VGND_c_503_n 0.00896865f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_80_21#_c_84_n A_275_47# 0.00461957f $X=1.85 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_80_21#_c_113_p A_363_47# 0.00753381f $X=3.085 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_80_21#_c_113_p A_563_47# 0.0084488f $X=3.085 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_80_21#_c_85_n A_563_47# 5.5126e-19 $X=3.037 $Y=1.785 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A3_M1004_g N_A2_M1000_g 0.0391232f $X=1.3 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A3_M1006_g N_A2_M1003_g 0.0163736f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_166 A3 N_A2_M1003_g 0.00181896f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A3_c_177_n N_A2_c_229_n 0.0124058f $X=1.17 $Y=1.4 $X2=0 $Y2=0
cc_168 N_A3_M1006_g N_A2_c_230_n 0.00436066f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A3_c_180_n N_A2_c_230_n 0.0124058f $X=1.17 $Y=1.605 $X2=0 $Y2=0
cc_170 A3 N_A2_c_230_n 2.88706e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A3_c_182_n N_A2_c_231_n 0.0124058f $X=1.13 $Y=1.1 $X2=0 $Y2=0
cc_172 N_A3_c_200_n N_A2_c_231_n 5.59836e-19 $X=1.13 $Y=1.1 $X2=0 $Y2=0
cc_173 N_A3_M1006_g N_A2_c_232_n 2.63865e-19 $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_174 A3 N_A2_c_232_n 0.0109178f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A3_c_182_n N_A2_c_232_n 0.003579f $X=1.13 $Y=1.1 $X2=0 $Y2=0
cc_176 N_A3_c_200_n N_A2_c_232_n 0.0430735f $X=1.13 $Y=1.1 $X2=0 $Y2=0
cc_177 N_A3_M1006_g N_VPWR_c_414_n 0.0102013f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A3_c_180_n N_VPWR_c_414_n 0.00105351f $X=1.17 $Y=1.605 $X2=0 $Y2=0
cc_179 A3 N_VPWR_c_414_n 0.0163082f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A3_M1006_g N_VPWR_c_415_n 4.58776e-19 $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A3_M1006_g N_VPWR_c_418_n 0.00428369f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A3_M1006_g N_VPWR_c_413_n 0.00462582f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A3_M1006_g N_A_269_429#_c_454_n 0.00294979f $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A3_M1006_g N_A_269_429#_c_456_n 0.00510928f $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A3_M1004_g N_VGND_c_500_n 0.00358332f $X=1.3 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A3_M1004_g N_VGND_c_502_n 0.010295f $X=1.3 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A3_M1004_g N_VGND_c_503_n 0.00431053f $X=1.3 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A2_M1000_g N_A1_M1007_g 0.0357011f $X=1.74 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A2_M1003_g N_A1_M1011_g 0.026273f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A2_c_229_n N_A1_M1011_g 0.00710144f $X=1.75 $Y=1.52 $X2=0 $Y2=0
cc_191 N_A2_c_232_n N_A1_M1011_g 9.22229e-19 $X=1.75 $Y=1.18 $X2=0 $Y2=0
cc_192 N_A2_c_231_n N_A1_c_282_n 0.0153117f $X=1.75 $Y=1.18 $X2=0 $Y2=0
cc_193 N_A2_c_232_n N_A1_c_282_n 4.52426e-19 $X=1.75 $Y=1.18 $X2=0 $Y2=0
cc_194 N_A2_c_229_n N_A1_c_283_n 0.0153117f $X=1.75 $Y=1.52 $X2=0 $Y2=0
cc_195 N_A2_M1000_g A1 0.00415834f $X=1.74 $Y=0.445 $X2=0 $Y2=0
cc_196 N_A2_c_231_n A1 0.00319995f $X=1.75 $Y=1.18 $X2=0 $Y2=0
cc_197 N_A2_c_232_n A1 0.0394742f $X=1.75 $Y=1.18 $X2=0 $Y2=0
cc_198 N_A2_M1003_g N_VPWR_c_414_n 4.81366e-19 $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A2_M1003_g N_VPWR_c_415_n 0.00903649f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A2_M1003_g N_VPWR_c_418_n 0.00443704f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A2_M1003_g N_VPWR_c_413_n 0.00478986f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A2_M1003_g N_A_269_429#_c_454_n 0.0019806f $X=1.795 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_A2_M1003_g N_A_269_429#_c_455_n 0.0158891f $X=1.795 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A2_c_230_n N_A_269_429#_c_455_n 0.00248229f $X=1.75 $Y=1.685 $X2=0
+ $Y2=0
cc_205 N_A2_c_232_n N_A_269_429#_c_455_n 0.0112663f $X=1.75 $Y=1.18 $X2=0 $Y2=0
cc_206 N_A2_c_230_n N_A_269_429#_c_456_n 0.00294791f $X=1.75 $Y=1.685 $X2=0
+ $Y2=0
cc_207 N_A2_c_232_n N_A_269_429#_c_456_n 0.0151547f $X=1.75 $Y=1.18 $X2=0 $Y2=0
cc_208 N_A2_M1003_g N_A_269_429#_c_457_n 6.00829e-19 $X=1.795 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_A2_M1000_g N_VGND_c_500_n 0.00362854f $X=1.74 $Y=0.445 $X2=0 $Y2=0
cc_210 N_A2_M1000_g N_VGND_c_502_n 0.00151897f $X=1.74 $Y=0.445 $X2=0 $Y2=0
cc_211 N_A2_M1000_g N_VGND_c_503_n 0.00558459f $X=1.74 $Y=0.445 $X2=0 $Y2=0
cc_212 N_A1_M1007_g N_B1_M1010_g 0.0178629f $X=2.2 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A1_M1011_g N_B1_M1001_g 0.0306498f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A1_c_282_n N_B1_c_323_n 0.0137828f $X=2.29 $Y=1.345 $X2=0 $Y2=0
cc_215 N_A1_c_283_n N_B1_c_324_n 0.0137828f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_216 A1 B1 0.0587775f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_217 N_A1_c_285_n B1 0.00448642f $X=2.29 $Y=1.005 $X2=0 $Y2=0
cc_218 A1 N_B1_c_326_n 5.83031e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_219 N_A1_c_285_n N_B1_c_326_n 0.0137828f $X=2.29 $Y=1.005 $X2=0 $Y2=0
cc_220 N_A1_M1011_g N_VPWR_c_415_n 0.00430572f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A1_M1011_g N_VPWR_c_419_n 0.00380959f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A1_M1011_g N_VPWR_c_413_n 0.00393687f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A1_M1011_g N_A_269_429#_c_455_n 0.0155194f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A1_c_283_n N_A_269_429#_c_455_n 0.0030797f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_225 A1 N_A_269_429#_c_455_n 0.016231f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_226 N_A1_M1011_g N_A_269_429#_c_457_n 0.0129564f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A1_M1011_g N_A_269_429#_c_459_n 9.82662e-19 $X=2.32 $Y=2.465 $X2=0
+ $Y2=0
cc_228 N_A1_M1007_g N_VGND_c_500_n 0.00363059f $X=2.2 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A1_M1007_g N_VGND_c_503_n 0.00581984f $X=2.2 $Y=0.445 $X2=0 $Y2=0
cc_230 N_B1_M1001_g N_B2_c_361_n 0.0251518f $X=2.77 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_231 N_B1_c_324_n N_B2_c_361_n 0.00356221f $X=2.83 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_232 N_B1_M1010_g N_B2_M1002_g 0.0216316f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_233 B1 N_B2_M1002_g 4.06374e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_234 N_B1_c_326_n N_B2_M1002_g 0.00816758f $X=2.83 $Y=1.005 $X2=0 $Y2=0
cc_235 N_B1_c_323_n N_B2_c_363_n 0.00816758f $X=2.83 $Y=1.345 $X2=0 $Y2=0
cc_236 N_B1_c_323_n N_B2_c_365_n 0.00356221f $X=2.83 $Y=1.345 $X2=0 $Y2=0
cc_237 N_B1_M1001_g N_VPWR_c_419_n 6.46133e-19 $X=2.77 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_M1001_g N_A_269_429#_c_455_n 0.00144788f $X=2.77 $Y=2.465 $X2=0
+ $Y2=0
cc_239 B1 N_A_269_429#_c_455_n 0.00583079f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_240 N_B1_M1001_g N_A_269_429#_c_457_n 0.00244297f $X=2.77 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_B1_M1001_g N_A_269_429#_c_458_n 0.00922642f $X=2.77 $Y=2.465 $X2=0
+ $Y2=0
cc_242 N_B1_M1010_g N_VGND_c_500_n 0.00363059f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_243 N_B1_M1010_g N_VGND_c_503_n 0.00600426f $X=2.74 $Y=0.445 $X2=0 $Y2=0
cc_244 N_B2_M1008_g N_VPWR_c_419_n 6.46133e-19 $X=3.2 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B2_M1008_g N_A_269_429#_c_458_n 0.00938123f $X=3.2 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B2_c_361_n N_A_269_429#_c_460_n 0.00791268f $X=3.2 $Y=1.9 $X2=0 $Y2=0
cc_247 N_B2_M1008_g N_A_269_429#_c_460_n 0.0036673f $X=3.2 $Y=2.465 $X2=0 $Y2=0
cc_248 B2 N_A_269_429#_c_460_n 0.0109535f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_249 N_B2_M1002_g N_VGND_c_499_n 0.00643628f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_250 N_B2_c_363_n N_VGND_c_499_n 0.00128212f $X=3.57 $Y=1.105 $X2=0 $Y2=0
cc_251 B2 N_VGND_c_499_n 0.0222009f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_252 N_B2_M1002_g N_VGND_c_500_n 0.00511208f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_253 N_B2_M1002_g N_VGND_c_503_n 0.0104194f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_254 B2 N_VGND_c_503_n 0.00431497f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_255 N_X_c_399_n N_VPWR_c_414_n 0.0145975f $X=0.625 $Y=2.29 $X2=0 $Y2=0
cc_256 N_X_c_399_n N_VPWR_c_416_n 0.025232f $X=0.625 $Y=2.29 $X2=0 $Y2=0
cc_257 N_X_c_399_n N_VPWR_c_413_n 0.0239906f $X=0.625 $Y=2.29 $X2=0 $Y2=0
cc_258 N_X_c_397_n N_VGND_c_501_n 0.0184996f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_259 N_X_M1005_s N_VGND_c_503_n 0.00371702f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_260 N_X_c_397_n N_VGND_c_503_n 0.0104061f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_261 N_VPWR_c_414_n N_A_269_429#_c_454_n 0.0264547f $X=1.055 $Y=2.29 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_415_n N_A_269_429#_c_454_n 0.0233002f $X=2.03 $Y=2.29 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_418_n N_A_269_429#_c_454_n 0.00825385f $X=1.865 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_413_n N_A_269_429#_c_454_n 0.0104525f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_c_415_n N_A_269_429#_c_455_n 0.0242265f $X=2.03 $Y=2.29 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_415_n N_A_269_429#_c_457_n 0.0298138f $X=2.03 $Y=2.29 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_419_n N_A_269_429#_c_458_n 0.0594494f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_c_413_n N_A_269_429#_c_458_n 0.0358658f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_c_415_n N_A_269_429#_c_459_n 0.0149473f $X=2.03 $Y=2.29 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_419_n N_A_269_429#_c_459_n 0.019216f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_271 N_VPWR_c_413_n N_A_269_429#_c_459_n 0.0110276f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VGND_c_503_n A_275_47# 0.00324374f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_273 N_VGND_c_503_n A_363_47# 0.00249632f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_274 N_VGND_c_503_n A_563_47# 0.00316062f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
