/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_LP__BUSHOLD0_1_V
`define SKY130_FD_SC_LP__BUSHOLD0_1_V

/**
 * bushold0: Bus signal holder (back-to-back inverter) with
 *           noninverting reset (gates internal node weak driver).
 *
 * Verilog wrapper for bushold0 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_lp__bushold0.v"

`ifdef USE_POWER_PINS
/*********************************************************/

`celldefine
module sky130_fd_sc_lp__bushold0_1 (
    X    ,
    RESET,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    inout X    ;
    input RESET;
    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_lp__bushold0 base (
        .X(X),
        .RESET(RESET),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/
`else // If not USE_POWER_PINS
/*********************************************************/

`celldefine
module sky130_fd_sc_lp__bushold0_1 (
    X    ,
    RESET,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    inout X    ;
    input RESET;
    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;

    // Voltage supply signals
    supply1 VPWR;
    supply0 VGND;
    supply1 VPB ;
    supply0 VNB ;

    sky130_fd_sc_lp__bushold0 base (
        .X(X),
        .RESET(RESET)
    );

endmodule
`endcelldefine

/*********************************************************/
`endif // USE_POWER_PINS

`default_nettype wire
`endif  // SKY130_FD_SC_LP__BUSHOLD0_1_V
