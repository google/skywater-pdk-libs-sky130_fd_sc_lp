* File: sky130_fd_sc_lp__a221o_m.pex.spice
* Created: Fri Aug 28 09:52:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221O_M%A_33_153# 1 2 3 12 14 17 21 25 27 31 34 35
+ 39 42 43 44 48 50 55
c112 50 0 2.87424e-20 $X=3.08 $Y=0.51
c113 39 0 1.83705e-19 $X=3.1 $Y=2.13
c114 31 0 1.46329e-19 $X=1.705 $Y=0.51
r115 52 53 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.75
+ $X2=3.08 $Y2=0.835
r116 50 52 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.08 $Y=0.51
+ $X2=3.08 $Y2=0.75
r117 44 46 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.07 $Y=1.48 $X2=1.07
+ $Y2=1.78
r118 43 56 79.6082 $w=6.1e-07 $l=5.05e-07 $layer=POLY_cond $X=0.47 $Y=1.86
+ $X2=0.47 $Y2=2.365
r119 43 55 49.7869 $w=6.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.86
+ $X2=0.47 $Y2=1.695
r120 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.86 $X2=0.61 $Y2=1.86
r121 39 53 59.6965 $w=2.48e-07 $l=1.295e-06 $layer=LI1_cond $X=3.12 $Y=2.13
+ $X2=3.12 $Y2=0.835
r122 36 48 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.81 $Y=0.75
+ $X2=1.715 $Y2=0.75
r123 35 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.75
+ $X2=3.08 $Y2=0.75
r124 35 36 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.915 $Y=0.75
+ $X2=1.81 $Y2=0.75
r125 33 48 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.705 $Y=0.835
+ $X2=1.715 $Y2=0.75
r126 33 34 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.705 $Y=0.835
+ $X2=1.705 $Y2=1.395
r127 29 48 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=0.665
+ $X2=1.715 $Y2=0.75
r128 29 31 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.715 $Y=0.665
+ $X2=1.715 $Y2=0.51
r129 28 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=1.48
+ $X2=1.07 $Y2=1.48
r130 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=1.48
+ $X2=1.705 $Y2=1.395
r131 27 28 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.62 $Y=1.48
+ $X2=1.155 $Y2=1.48
r132 26 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.78
+ $X2=0.61 $Y2=1.78
r133 25 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=1.78
+ $X2=1.07 $Y2=1.78
r134 25 26 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.985 $Y=1.78
+ $X2=0.695 $Y2=1.78
r135 19 21 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=0.24 $Y=0.84
+ $X2=0.475 $Y2=0.84
r136 17 56 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.66 $Y=2.885
+ $X2=0.66 $Y2=2.365
r137 12 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=0.765
+ $X2=0.475 $Y2=0.84
r138 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.765
+ $X2=0.475 $Y2=0.445
r139 10 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.24 $Y=0.915
+ $X2=0.24 $Y2=0.84
r140 10 55 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.24 $Y=0.915
+ $X2=0.24 $Y2=1.695
r141 3 39 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.985 $X2=3.1 $Y2=2.13
r142 2 50 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.51
r143 1 31 182 $w=1.7e-07 $l=4.83322e-07 $layer=licon1_NDIFF $count=1 $X=1.34
+ $Y=0.235 $X2=1.705 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%A2 3 7 9 10 16
c48 7 0 1.17366e-19 $X=1.09 $Y=2.885
r49 14 16 32.4255 $w=2.75e-07 $l=1.85e-07 $layer=POLY_cond $X=0.72 $Y=1.32
+ $X2=0.905 $Y2=1.32
r50 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.32 $X2=0.72 $Y2=1.32
r51 9 10 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=0.925 $X2=0.72
+ $Y2=1.295
r52 5 16 32.4255 $w=2.75e-07 $l=2.5446e-07 $layer=POLY_cond $X=1.09 $Y=1.485
+ $X2=0.905 $Y2=1.32
r53 5 7 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=1.09 $Y=1.485 $X2=1.09
+ $Y2=2.885
r54 1 16 16.9318 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.155
+ $X2=0.905 $Y2=1.32
r55 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.905 $Y=1.155
+ $X2=0.905 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%A1 1 3 6 8 9 17
c46 6 0 1.47633e-19 $X=1.52 $Y=2.885
r47 15 17 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=0.93
+ $X2=1.52 $Y2=0.93
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.355
+ $Y=0.93 $X2=1.355 $Y2=0.93
r49 12 15 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.265 $Y=0.93
+ $X2=1.355 $Y2=0.93
r50 9 16 0.177299 $w=3.23e-07 $l=5e-09 $layer=LI1_cond $X=1.277 $Y=0.925
+ $X2=1.277 $Y2=0.93
r51 8 9 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.277 $Y=0.555
+ $X2=1.277 $Y2=0.925
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.095
+ $X2=1.52 $Y2=0.93
r53 4 6 917.851 $w=1.5e-07 $l=1.79e-06 $layer=POLY_cond $X=1.52 $Y=1.095
+ $X2=1.52 $Y2=2.885
r54 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=0.765
+ $X2=1.265 $Y2=0.93
r55 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.265 $Y=0.765
+ $X2=1.265 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%B1 3 7 9 12
c39 9 0 1.47633e-19 $X=2.16 $Y=1.295
r40 12 15 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.032 $Y=1.32
+ $X2=2.032 $Y2=1.485
r41 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.032 $Y=1.32
+ $X2=2.032 $Y2=1.155
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.32 $X2=2.055 $Y2=1.32
r43 9 13 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=1.32
+ $X2=2.055 $Y2=1.32
r44 7 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.025 $Y=2.195
+ $X2=2.025 $Y2=1.485
r45 3 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.92 $Y=0.445
+ $X2=1.92 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%B2 1 3 6 14 16 17 18 21 23
c49 17 0 1.63183e-19 $X=2.48 $Y=1.845
c50 14 0 2.87424e-20 $X=2.505 $Y=0.84
c51 6 0 2.05222e-20 $X=2.455 $Y=2.195
r52 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.595 $Y=1.32
+ $X2=2.595 $Y2=1.485
r53 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.595 $Y=1.32
+ $X2=2.595 $Y2=1.155
r54 18 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.595
+ $Y=1.32 $X2=2.595 $Y2=1.32
r55 16 17 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.48 $Y=1.695 $X2=2.48
+ $Y2=1.845
r56 16 24 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.505 $Y=1.695
+ $X2=2.505 $Y2=1.485
r57 12 14 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.28 $Y=0.84
+ $X2=2.505 $Y2=0.84
r58 8 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=0.915
+ $X2=2.505 $Y2=0.84
r59 8 23 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.505 $Y=0.915
+ $X2=2.505 $Y2=1.155
r60 6 17 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.455 $Y=2.195
+ $X2=2.455 $Y2=1.845
r61 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=0.765
+ $X2=2.28 $Y2=0.84
r62 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.28 $Y=0.765 $X2=2.28
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%C1 1 3 7 9 12 16 18 19 26
r39 23 26 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.785 $Y=2.91
+ $X2=2.885 $Y2=2.91
r40 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=2.91 $X2=2.785 $Y2=2.91
r41 19 24 10.0278 $w=3.83e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=2.882
+ $X2=2.785 $Y2=2.882
r42 18 24 4.34037 $w=3.83e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=2.882
+ $X2=2.785 $Y2=2.882
r43 14 16 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.885 $Y=1.8
+ $X2=3.075 $Y2=1.8
r44 10 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.865 $Y=0.84
+ $X2=3.075 $Y2=0.84
r45 9 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.075 $Y=1.725
+ $X2=3.075 $Y2=1.8
r46 8 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.075 $Y=0.915
+ $X2=3.075 $Y2=0.84
r47 8 9 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.075 $Y=0.915
+ $X2=3.075 $Y2=1.725
r48 5 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=2.745
+ $X2=2.885 $Y2=2.91
r49 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.885 $Y=2.745
+ $X2=2.885 $Y2=2.195
r50 4 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=1.875
+ $X2=2.885 $Y2=1.8
r51 4 7 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.885 $Y=1.875
+ $X2=2.885 $Y2=2.195
r52 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=0.765
+ $X2=2.865 $Y2=0.84
r53 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.865 $Y=0.765
+ $X2=2.865 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%X 1 2 7 8 9 10 11 12 13 41
r25 39 41 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.25 $Y=2.82
+ $X2=0.445 $Y2=2.82
r26 21 39 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.25 $Y=2.655
+ $X2=0.25 $Y2=2.82
r27 13 39 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=2.82 $X2=0.25
+ $Y2=2.82
r28 12 21 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=0.25 $Y=2.405
+ $X2=0.25 $Y2=2.655
r29 11 12 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.035
+ $X2=0.25 $Y2=2.405
r30 10 11 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=2.035
r31 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r32 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=0.925 $X2=0.25
+ $Y2=1.295
r33 7 8 24.2249 $w=1.88e-07 $l=4.15e-07 $layer=LI1_cond $X=0.25 $Y=0.51 $X2=0.25
+ $Y2=0.925
r34 2 41 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.32
+ $Y=2.675 $X2=0.445 $Y2=2.82
r35 1 7 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%VPWR 1 2 9 13 16 17 18 24 33 34 37
r35 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r38 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=3.33
+ $X2=1.735 $Y2=3.33
r40 28 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.9 $Y=3.33 $X2=2.16
+ $Y2=3.33
r41 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.735 $Y2=3.33
r43 24 26 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 18 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 16 21 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=3.33 $X2=0.72
+ $Y2=3.33
r50 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.77 $Y=3.33
+ $X2=0.875 $Y2=3.33
r51 15 26 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.875 $Y2=3.33
r53 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=3.245
+ $X2=1.735 $Y2=3.33
r54 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.735 $Y=3.245
+ $X2=1.735 $Y2=2.95
r55 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r56 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.95
r57 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.675 $X2=1.735 $Y2=2.95
r58 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=2.675 $X2=0.875 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%A_233_535# 1 2 9 11 12 15
c23 9 0 2.86637e-19 $X=1.305 $Y=2.82
r24 13 15 12.4113 $w=2.08e-07 $l=2.35e-07 $layer=LI1_cond $X=2.24 $Y=2.495
+ $X2=2.24 $Y2=2.26
r25 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.135 $Y=2.58
+ $X2=2.24 $Y2=2.495
r26 11 12 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.135 $Y=2.58
+ $X2=1.39 $Y2=2.58
r27 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.295 $Y=2.665
+ $X2=1.39 $Y2=2.58
r28 7 9 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.295 $Y=2.665
+ $X2=1.295 $Y2=2.82
r29 2 15 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.985 $X2=2.24 $Y2=2.26
r30 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=2.675 $X2=1.305 $Y2=2.82
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%A_337_397# 1 2 9 11 12 15
r27 13 15 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.67 $Y=1.915
+ $X2=2.67 $Y2=2.13
r28 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.565 $Y=1.83
+ $X2=2.67 $Y2=1.915
r29 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.565 $Y=1.83
+ $X2=1.915 $Y2=1.83
r30 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.81 $Y=1.915
+ $X2=1.915 $Y2=1.83
r31 7 9 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.81 $Y=1.915 $X2=1.81
+ $Y2=2.13
r32 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.985 $X2=2.67 $Y2=2.13
r33 1 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.985 $X2=1.81 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_M%VGND 1 2 9 13 16 17 18 20 33 34 37
r54 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r56 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r57 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r58 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r59 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r60 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r62 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r63 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r64 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r66 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r67 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r68 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r69 16 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.16
+ $Y2=0
r70 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.495
+ $Y2=0
r71 15 33 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.66 $Y=0 $X2=3.12
+ $Y2=0
r72 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.66 $Y=0 $X2=2.495
+ $Y2=0
r73 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=0.085
+ $X2=2.495 $Y2=0
r74 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.495 $Y=0.085
+ $X2=2.495 $Y2=0.38
r75 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r76 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r77 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.495 $Y2=0.38
r78 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

