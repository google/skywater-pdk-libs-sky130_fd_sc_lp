* File: sky130_fd_sc_lp__clkinv_8.spice
* Created: Wed Sep  2 09:40:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkinv_8.pex.spice"
.subckt sky130_fd_sc_lp__clkinv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.2 A=0.063
+ P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002.8 A=0.063
+ P=1.14 MULT=1
MM1004 N_VGND_M1002_d N_A_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.3 A=0.063
+ P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75001.9 A=0.063
+ P=1.14 MULT=1
MM1009 N_VGND_M1006_d N_A_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75001.5 A=0.063
+ P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75001.1 A=0.063
+ P=1.14 MULT=1
MM1013 N_VGND_M1011_d N_A_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1005_d N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1008_d N_A_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1012_d N_A_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1015_d N_A_M1015_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1015_d N_A_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1017_d N_A_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__clkinv_8.pxi.spice"
*
.ends
*
*
