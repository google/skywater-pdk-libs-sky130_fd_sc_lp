* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand2b_1 A_N B VGND VNB VPB VPWR Y
M1000 VGND A_N a_40_367# VNB nshort w=420000u l=150000u
+  ad=2.562e+11p pd=2.4e+06u as=1.113e+11p ps=1.37e+06u
M1001 Y a_40_367# a_269_47# VNB nshort w=840000u l=150000u
+  ad=2.856e+11p pd=2.36e+06u as=1.764e+11p ps=2.1e+06u
M1002 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=7.14e+11p ps=6.32e+06u
M1003 a_269_47# B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A_N a_40_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VPWR a_40_367# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
