* File: sky130_fd_sc_lp__or3b_m.pxi.spice
* Created: Wed Sep  2 10:31:34 2020
* 
x_PM_SKY130_FD_SC_LP__OR3B_M%C_N N_C_N_c_80_n N_C_N_M1000_g N_C_N_M1005_g
+ N_C_N_c_82_n N_C_N_c_83_n N_C_N_c_88_n C_N C_N C_N C_N C_N N_C_N_c_85_n
+ PM_SKY130_FD_SC_LP__OR3B_M%C_N
x_PM_SKY130_FD_SC_LP__OR3B_M%A_112_55# N_A_112_55#_M1000_d N_A_112_55#_M1005_d
+ N_A_112_55#_c_116_n N_A_112_55#_c_117_n N_A_112_55#_c_118_n
+ N_A_112_55#_c_119_n N_A_112_55#_M1004_g N_A_112_55#_c_121_n
+ N_A_112_55#_M1008_g N_A_112_55#_c_122_n N_A_112_55#_c_123_n
+ N_A_112_55#_c_124_n N_A_112_55#_c_125_n N_A_112_55#_c_126_n
+ N_A_112_55#_c_130_n N_A_112_55#_c_131_n PM_SKY130_FD_SC_LP__OR3B_M%A_112_55#
x_PM_SKY130_FD_SC_LP__OR3B_M%B N_B_M1003_g N_B_M1002_g N_B_c_175_n N_B_c_180_n B
+ B N_B_c_177_n PM_SKY130_FD_SC_LP__OR3B_M%B
x_PM_SKY130_FD_SC_LP__OR3B_M%A N_A_M1007_g N_A_M1009_g A A A N_A_c_212_n
+ N_A_c_213_n PM_SKY130_FD_SC_LP__OR3B_M%A
x_PM_SKY130_FD_SC_LP__OR3B_M%A_212_418# N_A_212_418#_M1008_s
+ N_A_212_418#_M1002_d N_A_212_418#_M1004_s N_A_212_418#_M1001_g
+ N_A_212_418#_M1006_g N_A_212_418#_c_243_n N_A_212_418#_c_244_n
+ N_A_212_418#_c_245_n N_A_212_418#_c_246_n N_A_212_418#_c_258_n
+ N_A_212_418#_c_259_n N_A_212_418#_c_247_n N_A_212_418#_c_248_n
+ N_A_212_418#_c_249_n N_A_212_418#_c_250_n N_A_212_418#_c_251_n
+ N_A_212_418#_c_252_n N_A_212_418#_c_253_n N_A_212_418#_c_254_n
+ N_A_212_418#_c_255_n PM_SKY130_FD_SC_LP__OR3B_M%A_212_418#
x_PM_SKY130_FD_SC_LP__OR3B_M%VPWR N_VPWR_M1005_s N_VPWR_M1009_d N_VPWR_c_328_n
+ N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_344_n N_VPWR_c_331_n N_VPWR_c_332_n
+ VPWR N_VPWR_c_333_n N_VPWR_c_327_n PM_SKY130_FD_SC_LP__OR3B_M%VPWR
x_PM_SKY130_FD_SC_LP__OR3B_M%X N_X_M1001_d N_X_M1006_d X X X X X X X N_X_c_366_n
+ X PM_SKY130_FD_SC_LP__OR3B_M%X
x_PM_SKY130_FD_SC_LP__OR3B_M%VGND N_VGND_M1000_s N_VGND_M1008_d N_VGND_M1007_d
+ N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n
+ N_VGND_c_386_n VGND N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n
+ N_VGND_c_390_n PM_SKY130_FD_SC_LP__OR3B_M%VGND
cc_1 VNB N_C_N_c_80_n 0.0089214f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.14
cc_2 VNB N_C_N_M1000_g 0.0279762f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.485
cc_3 VNB N_C_N_c_82_n 0.0349411f $X=-0.19 $Y=-0.245 $X2=0.332 $Y2=0.99
cc_4 VNB N_C_N_c_83_n 0.0236153f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_5 VNB C_N 0.00722069f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_C_N_c_85_n 0.0381401f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_A_112_55#_c_116_n 0.0148937f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.885
cc_8 VNB N_A_112_55#_c_117_n 0.0330738f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.885
cc_9 VNB N_A_112_55#_c_118_n 0.0110125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_112_55#_c_119_n 0.0248141f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_11 VNB N_A_112_55#_M1004_g 0.0130713f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_12 VNB N_A_112_55#_c_121_n 0.0194921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_112_55#_c_122_n 0.0121271f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_A_112_55#_c_123_n 0.010886f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_15 VNB N_A_112_55#_c_124_n 0.00175081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_112_55#_c_125_n 0.00314808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_112_55#_c_126_n 0.0181041f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_18 VNB N_B_M1002_g 0.0397239f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.29
cc_19 VNB N_B_c_175_n 0.02037f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_20 VNB B 0.00492219f $X=-0.19 $Y=-0.245 $X2=0.332 $Y2=0.99
cc_21 VNB N_B_c_177_n 0.0189317f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.215
cc_22 VNB N_A_M1007_g 0.0595293f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.84
cc_23 VNB N_A_212_418#_M1006_g 0.0111309f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_24 VNB N_A_212_418#_c_243_n 0.0199613f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.215
cc_25 VNB N_A_212_418#_c_244_n 0.0231252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_212_418#_c_245_n 0.0181522f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_27 VNB N_A_212_418#_c_246_n 0.0103079f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_A_212_418#_c_247_n 0.00227233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_212_418#_c_248_n 0.00980478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_212_418#_c_249_n 0.00902549f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_31 VNB N_A_212_418#_c_250_n 0.00186787f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_32 VNB N_A_212_418#_c_251_n 0.00358309f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_33 VNB N_A_212_418#_c_252_n 0.00191403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_212_418#_c_253_n 7.39423e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_212_418#_c_254_n 0.0162882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_212_418#_c_255_n 0.0012964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_327_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_38 VNB X 0.0646428f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.29
cc_39 VNB N_VGND_c_381_n 0.0114773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_382_n 0.00685879f $X=-0.19 $Y=-0.245 $X2=0.332 $Y2=0.84
cc_41 VNB N_VGND_c_383_n 0.00454526f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.215
cc_42 VNB N_VGND_c_384_n 0.00454526f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_43 VNB N_VGND_c_385_n 0.0190583f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_44 VNB N_VGND_c_386_n 0.00401194f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_45 VNB N_VGND_c_387_n 0.0348217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_388_n 0.0218749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_389_n 0.203509f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_48 VNB N_VGND_c_390_n 0.00401194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VPB N_C_N_c_80_n 0.0311274f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.14
cc_50 VPB N_C_N_M1005_g 0.0430703f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.885
cc_51 VPB N_C_N_c_88_n 0.0240241f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.215
cc_52 VPB C_N 0.0329613f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_53 VPB N_A_112_55#_M1004_g 0.0349293f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_54 VPB N_A_112_55#_c_124_n 5.34031e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_112_55#_c_126_n 0.0277708f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_56 VPB N_A_112_55#_c_130_n 0.0192296f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_57 VPB N_A_112_55#_c_131_n 0.00595322f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_58 VPB N_B_M1003_g 0.0233139f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.84
cc_59 VPB N_B_c_175_n 5.57233e-19 $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_60 VPB N_B_c_180_n 0.0152787f $X=-0.19 $Y=1.655 $X2=0.332 $Y2=0.84
cc_61 VPB B 0.00167341f $X=-0.19 $Y=1.655 $X2=0.332 $Y2=0.99
cc_62 VPB N_A_M1007_g 0.033037f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.84
cc_63 VPB N_A_c_212_n 0.042888f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_64 VPB N_A_c_213_n 0.0324212f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_65 VPB N_A_212_418#_M1006_g 0.0359485f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_66 VPB N_A_212_418#_c_246_n 0.00408061f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_67 VPB N_A_212_418#_c_258_n 0.0146034f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_68 VPB N_A_212_418#_c_259_n 0.0089521f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_69 VPB N_A_212_418#_c_252_n 0.00259989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_328_n 0.0110915f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.29
cc_71 VPB N_VPWR_c_329_n 0.00484226f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.885
cc_72 VPB N_VPWR_c_330_n 0.0255447f $X=-0.19 $Y=1.655 $X2=0.332 $Y2=0.84
cc_73 VPB N_VPWR_c_331_n 0.0575352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_332_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_75 VPB N_VPWR_c_333_n 0.0214303f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_76 VPB N_VPWR_c_327_n 0.0823103f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_77 VPB X 0.0246939f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.29
cc_78 VPB X 0.00536733f $X=-0.19 $Y=1.655 $X2=0.332 $Y2=0.84
cc_79 VPB N_X_c_366_n 0.0283187f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_80 N_C_N_c_82_n N_A_112_55#_c_116_n 0.00422685f $X=0.332 $Y=0.99 $X2=0 $Y2=0
cc_81 N_C_N_c_85_n N_A_112_55#_c_116_n 0.00519952f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_82 N_C_N_M1000_g N_A_112_55#_c_118_n 0.00422685f $X=0.485 $Y=0.485 $X2=0
+ $Y2=0
cc_83 C_N N_A_112_55#_c_122_n 6.67444e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_C_N_c_85_n N_A_112_55#_c_122_n 0.0170497f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_85 N_C_N_M1000_g N_A_112_55#_c_123_n 0.00633408f $X=0.485 $Y=0.485 $X2=0
+ $Y2=0
cc_86 C_N N_A_112_55#_c_123_n 0.0959007f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_87 N_C_N_c_85_n N_A_112_55#_c_123_n 0.00384495f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_88 N_C_N_c_83_n N_A_112_55#_c_125_n 0.00384495f $X=0.27 $Y=1.51 $X2=0 $Y2=0
cc_89 N_C_N_c_83_n N_A_112_55#_c_126_n 0.0170497f $X=0.27 $Y=1.51 $X2=0 $Y2=0
cc_90 N_C_N_c_88_n N_A_112_55#_c_130_n 0.0162282f $X=0.485 $Y=2.215 $X2=0 $Y2=0
cc_91 N_C_N_c_80_n N_A_112_55#_c_131_n 0.00384495f $X=0.36 $Y=2.14 $X2=0 $Y2=0
cc_92 N_C_N_M1000_g N_A_212_418#_c_253_n 0.00107555f $X=0.485 $Y=0.485 $X2=0
+ $Y2=0
cc_93 N_C_N_M1005_g N_VPWR_c_329_n 0.00442088f $X=0.485 $Y=2.885 $X2=0 $Y2=0
cc_94 N_C_N_c_88_n N_VPWR_c_329_n 3.39155e-19 $X=0.485 $Y=2.215 $X2=0 $Y2=0
cc_95 C_N N_VPWR_c_329_n 0.0104807f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_96 N_C_N_M1005_g N_VPWR_c_331_n 0.00585385f $X=0.485 $Y=2.885 $X2=0 $Y2=0
cc_97 N_C_N_M1005_g N_VPWR_c_327_n 0.0130948f $X=0.485 $Y=2.885 $X2=0 $Y2=0
cc_98 C_N N_VPWR_c_327_n 0.00131218f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_99 N_C_N_M1000_g N_VGND_c_382_n 0.00468315f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_100 N_C_N_c_82_n N_VGND_c_382_n 0.00138828f $X=0.332 $Y=0.99 $X2=0 $Y2=0
cc_101 C_N N_VGND_c_382_n 0.0111969f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_102 N_C_N_M1000_g N_VGND_c_387_n 0.00545548f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_103 N_C_N_M1000_g N_VGND_c_389_n 0.0120886f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_104 N_C_N_c_82_n N_VGND_c_389_n 0.00221078f $X=0.332 $Y=0.99 $X2=0 $Y2=0
cc_105 C_N N_VGND_c_389_n 0.00110271f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_106 N_A_112_55#_c_121_n N_B_M1002_g 0.0214476f $X=1.46 $Y=0.77 $X2=0 $Y2=0
cc_107 N_A_112_55#_M1004_g N_B_c_180_n 0.0430988f $X=1.42 $Y=2.3 $X2=0 $Y2=0
cc_108 N_A_112_55#_c_119_n B 0.00400714f $X=1.345 $Y=1.305 $X2=0 $Y2=0
cc_109 N_A_112_55#_c_119_n N_B_c_177_n 0.0430988f $X=1.345 $Y=1.305 $X2=0 $Y2=0
cc_110 N_A_112_55#_M1004_g N_A_c_213_n 0.00514348f $X=1.42 $Y=2.3 $X2=0 $Y2=0
cc_111 N_A_112_55#_c_130_n N_A_c_213_n 0.0172341f $X=0.7 $Y=2.82 $X2=0 $Y2=0
cc_112 N_A_112_55#_c_116_n N_A_212_418#_c_246_n 0.00275765f $X=0.93 $Y=1.23
+ $X2=0 $Y2=0
cc_113 N_A_112_55#_c_117_n N_A_212_418#_c_246_n 0.0135252f $X=1.385 $Y=0.845
+ $X2=0 $Y2=0
cc_114 N_A_112_55#_c_119_n N_A_212_418#_c_246_n 0.0103097f $X=1.345 $Y=1.305
+ $X2=0 $Y2=0
cc_115 N_A_112_55#_M1004_g N_A_212_418#_c_246_n 0.0162797f $X=1.42 $Y=2.3 $X2=0
+ $Y2=0
cc_116 N_A_112_55#_c_123_n N_A_212_418#_c_246_n 0.0236591f $X=0.7 $Y=0.55 $X2=0
+ $Y2=0
cc_117 N_A_112_55#_c_125_n N_A_212_418#_c_246_n 0.0365252f $X=0.84 $Y=1.395
+ $X2=0 $Y2=0
cc_118 N_A_112_55#_c_126_n N_A_212_418#_c_246_n 0.00407346f $X=0.84 $Y=1.395
+ $X2=0 $Y2=0
cc_119 N_A_112_55#_c_130_n N_A_212_418#_c_246_n 0.0100854f $X=0.7 $Y=2.82 $X2=0
+ $Y2=0
cc_120 N_A_112_55#_M1004_g N_A_212_418#_c_259_n 0.0117862f $X=1.42 $Y=2.3 $X2=0
+ $Y2=0
cc_121 N_A_112_55#_c_130_n N_A_212_418#_c_259_n 0.0152527f $X=0.7 $Y=2.82 $X2=0
+ $Y2=0
cc_122 N_A_112_55#_c_117_n N_A_212_418#_c_253_n 0.00158117f $X=1.385 $Y=0.845
+ $X2=0 $Y2=0
cc_123 N_A_112_55#_c_121_n N_A_212_418#_c_253_n 0.00311102f $X=1.46 $Y=0.77
+ $X2=0 $Y2=0
cc_124 N_A_112_55#_c_123_n N_A_212_418#_c_253_n 0.0134648f $X=0.7 $Y=0.55 $X2=0
+ $Y2=0
cc_125 N_A_112_55#_c_130_n N_VPWR_c_331_n 0.00877924f $X=0.7 $Y=2.82 $X2=0 $Y2=0
cc_126 N_A_112_55#_M1005_d N_VPWR_c_327_n 0.0042053f $X=0.56 $Y=2.675 $X2=0
+ $Y2=0
cc_127 N_A_112_55#_c_130_n N_VPWR_c_327_n 0.00770513f $X=0.7 $Y=2.82 $X2=0 $Y2=0
cc_128 N_A_112_55#_c_121_n N_VGND_c_383_n 0.00284272f $X=1.46 $Y=0.77 $X2=0
+ $Y2=0
cc_129 N_A_112_55#_c_117_n N_VGND_c_387_n 9.55955e-19 $X=1.385 $Y=0.845 $X2=0
+ $Y2=0
cc_130 N_A_112_55#_c_118_n N_VGND_c_387_n 0.00509037f $X=1.005 $Y=0.845 $X2=0
+ $Y2=0
cc_131 N_A_112_55#_c_121_n N_VGND_c_387_n 0.0058025f $X=1.46 $Y=0.77 $X2=0 $Y2=0
cc_132 N_A_112_55#_c_123_n N_VGND_c_387_n 0.0075246f $X=0.7 $Y=0.55 $X2=0 $Y2=0
cc_133 N_A_112_55#_c_118_n N_VGND_c_389_n 0.00763919f $X=1.005 $Y=0.845 $X2=0
+ $Y2=0
cc_134 N_A_112_55#_c_121_n N_VGND_c_389_n 0.0120492f $X=1.46 $Y=0.77 $X2=0 $Y2=0
cc_135 N_A_112_55#_c_123_n N_VGND_c_389_n 0.00751788f $X=0.7 $Y=0.55 $X2=0 $Y2=0
cc_136 N_B_M1003_g N_A_M1007_g 0.0261114f $X=1.78 $Y=2.3 $X2=0 $Y2=0
cc_137 N_B_M1002_g N_A_M1007_g 0.0317119f $X=1.89 $Y=0.45 $X2=0 $Y2=0
cc_138 B N_A_M1007_g 0.00205514f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_139 N_B_c_177_n N_A_M1007_g 0.0416221f $X=1.87 $Y=1.325 $X2=0 $Y2=0
cc_140 N_B_M1003_g N_A_c_213_n 0.00565832f $X=1.78 $Y=2.3 $X2=0 $Y2=0
cc_141 N_B_M1002_g N_A_212_418#_c_246_n 0.00621165f $X=1.89 $Y=0.45 $X2=0 $Y2=0
cc_142 N_B_c_180_n N_A_212_418#_c_246_n 9.05089e-19 $X=1.87 $Y=1.83 $X2=0 $Y2=0
cc_143 B N_A_212_418#_c_246_n 0.0318941f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_B_c_177_n N_A_212_418#_c_246_n 0.00209001f $X=1.87 $Y=1.325 $X2=0 $Y2=0
cc_145 N_B_M1003_g N_A_212_418#_c_258_n 0.0117159f $X=1.78 $Y=2.3 $X2=0 $Y2=0
cc_146 N_B_c_180_n N_A_212_418#_c_258_n 0.00515738f $X=1.87 $Y=1.83 $X2=0 $Y2=0
cc_147 B N_A_212_418#_c_258_n 0.0245115f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 B N_A_212_418#_c_259_n 0.00885311f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_149 N_B_M1002_g N_A_212_418#_c_247_n 0.00156803f $X=1.89 $Y=0.45 $X2=0 $Y2=0
cc_150 N_B_M1002_g N_A_212_418#_c_249_n 0.00287294f $X=1.89 $Y=0.45 $X2=0 $Y2=0
cc_151 B N_A_212_418#_c_249_n 0.00210796f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B_c_177_n N_A_212_418#_c_249_n 9.50511e-19 $X=1.87 $Y=1.325 $X2=0 $Y2=0
cc_153 B N_A_212_418#_c_251_n 0.0174819f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_B_M1003_g N_VPWR_c_344_n 8.77009e-19 $X=1.78 $Y=2.3 $X2=0 $Y2=0
cc_155 N_B_M1002_g N_VGND_c_383_n 0.00154346f $X=1.89 $Y=0.45 $X2=0 $Y2=0
cc_156 B N_VGND_c_383_n 0.00545902f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_157 N_B_c_177_n N_VGND_c_383_n 0.00137474f $X=1.87 $Y=1.325 $X2=0 $Y2=0
cc_158 N_B_M1002_g N_VGND_c_385_n 0.0058025f $X=1.89 $Y=0.45 $X2=0 $Y2=0
cc_159 N_B_M1002_g N_VGND_c_389_n 0.0107259f $X=1.89 $Y=0.45 $X2=0 $Y2=0
cc_160 N_A_M1007_g N_A_212_418#_M1006_g 0.0297496f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_161 N_A_M1007_g N_A_212_418#_c_243_n 0.0148859f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_162 N_A_M1007_g N_A_212_418#_c_258_n 0.0178606f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_163 N_A_c_212_n N_A_212_418#_c_258_n 0.00229431f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_164 N_A_c_213_n N_A_212_418#_c_258_n 0.0177235f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_165 N_A_c_213_n N_A_212_418#_c_259_n 0.0256842f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_166 N_A_M1007_g N_A_212_418#_c_247_n 0.00288865f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_167 N_A_M1007_g N_A_212_418#_c_248_n 0.0154054f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_168 N_A_M1007_g N_A_212_418#_c_251_n 0.0145707f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_169 N_A_M1007_g N_A_212_418#_c_254_n 0.0405345f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_170 N_A_M1007_g N_VPWR_c_330_n 0.00428126f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_171 N_A_c_212_n N_VPWR_c_330_n 0.00808304f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_172 N_A_c_213_n N_VPWR_c_330_n 0.0245778f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_173 N_A_M1007_g N_VPWR_c_344_n 0.00507333f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_174 N_A_c_212_n N_VPWR_c_331_n 0.00815497f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_175 N_A_c_213_n N_VPWR_c_331_n 0.0556879f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_176 N_A_c_212_n N_VPWR_c_327_n 0.0106807f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_177 N_A_c_213_n N_VPWR_c_327_n 0.0447256f $X=2.26 $Y=2.835 $X2=0 $Y2=0
cc_178 N_A_M1007_g N_VGND_c_384_n 0.00154346f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_179 N_A_M1007_g N_VGND_c_385_n 0.0058025f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_180 N_A_M1007_g N_VGND_c_389_n 0.00614687f $X=2.32 $Y=0.45 $X2=0 $Y2=0
cc_181 N_A_212_418#_c_258_n N_VPWR_M1009_d 0.00233158f $X=2.575 $Y=2.015 $X2=0
+ $Y2=0
cc_182 N_A_212_418#_M1006_g N_VPWR_c_330_n 0.00116737f $X=2.795 $Y=2.3 $X2=0
+ $Y2=0
cc_183 N_A_212_418#_c_258_n N_VPWR_c_344_n 0.017236f $X=2.575 $Y=2.015 $X2=0
+ $Y2=0
cc_184 N_A_212_418#_M1006_g N_VPWR_c_333_n 0.00325938f $X=2.795 $Y=2.3 $X2=0
+ $Y2=0
cc_185 N_A_212_418#_M1006_g N_VPWR_c_327_n 0.00418739f $X=2.795 $Y=2.3 $X2=0
+ $Y2=0
cc_186 N_A_212_418#_c_259_n A_299_418# 0.00143222f $X=1.7 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_212_418#_c_258_n A_371_418# 0.00510366f $X=2.575 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_212_418#_M1006_g X 0.0163771f $X=2.795 $Y=2.3 $X2=0 $Y2=0
cc_189 N_A_212_418#_c_243_n X 0.00540106f $X=2.77 $Y=0.775 $X2=0 $Y2=0
cc_190 N_A_212_418#_c_258_n X 0.00907059f $X=2.575 $Y=2.015 $X2=0 $Y2=0
cc_191 N_A_212_418#_c_250_n X 0.0129659f $X=2.715 $Y=0.945 $X2=0 $Y2=0
cc_192 N_A_212_418#_c_251_n X 0.0354397f $X=2.715 $Y=1.305 $X2=0 $Y2=0
cc_193 N_A_212_418#_c_252_n X 0.0232649f $X=2.66 $Y=1.93 $X2=0 $Y2=0
cc_194 N_A_212_418#_c_254_n X 0.0191893f $X=2.77 $Y=0.94 $X2=0 $Y2=0
cc_195 N_A_212_418#_M1006_g N_X_c_366_n 0.00300841f $X=2.795 $Y=2.3 $X2=0 $Y2=0
cc_196 N_A_212_418#_c_243_n N_VGND_c_384_n 0.00284272f $X=2.77 $Y=0.775 $X2=0
+ $Y2=0
cc_197 N_A_212_418#_c_248_n N_VGND_c_384_n 0.00833303f $X=2.575 $Y=0.86 $X2=0
+ $Y2=0
cc_198 N_A_212_418#_c_250_n N_VGND_c_384_n 0.00357657f $X=2.715 $Y=0.945 $X2=0
+ $Y2=0
cc_199 N_A_212_418#_c_247_n N_VGND_c_385_n 0.00748063f $X=2.105 $Y=0.535 $X2=0
+ $Y2=0
cc_200 N_A_212_418#_c_253_n N_VGND_c_387_n 0.0085197f $X=1.245 $Y=0.515 $X2=0
+ $Y2=0
cc_201 N_A_212_418#_c_243_n N_VGND_c_388_n 0.0058025f $X=2.77 $Y=0.775 $X2=0
+ $Y2=0
cc_202 N_A_212_418#_c_254_n N_VGND_c_388_n 5.91418e-19 $X=2.77 $Y=0.94 $X2=0
+ $Y2=0
cc_203 N_A_212_418#_M1008_s N_VGND_c_389_n 0.00288564f $X=1.12 $Y=0.24 $X2=0
+ $Y2=0
cc_204 N_A_212_418#_M1002_d N_VGND_c_389_n 0.00379116f $X=1.965 $Y=0.24 $X2=0
+ $Y2=0
cc_205 N_A_212_418#_c_243_n N_VGND_c_389_n 0.00710949f $X=2.77 $Y=0.775 $X2=0
+ $Y2=0
cc_206 N_A_212_418#_c_247_n N_VGND_c_389_n 0.00754439f $X=2.105 $Y=0.535 $X2=0
+ $Y2=0
cc_207 N_A_212_418#_c_248_n N_VGND_c_389_n 0.00747856f $X=2.575 $Y=0.86 $X2=0
+ $Y2=0
cc_208 N_A_212_418#_c_250_n N_VGND_c_389_n 0.00775001f $X=2.715 $Y=0.945 $X2=0
+ $Y2=0
cc_209 N_A_212_418#_c_253_n N_VGND_c_389_n 0.00764888f $X=1.245 $Y=0.515 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_330_n N_X_c_366_n 0.0224421f $X=2.615 $Y=3.245 $X2=0 $Y2=0
cc_211 N_VPWR_c_333_n N_X_c_366_n 0.00832801f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_327_n N_X_c_366_n 0.00949235f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_213 X N_VGND_c_388_n 0.0210075f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_214 N_X_M1001_d N_VGND_c_389_n 0.00236247f $X=2.825 $Y=0.24 $X2=0 $Y2=0
cc_215 X N_VGND_c_389_n 0.0130934f $X=3.035 $Y=0.47 $X2=0 $Y2=0
