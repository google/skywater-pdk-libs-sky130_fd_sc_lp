* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2oi_0 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 Y a_110_47# a_420_387# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_420_387# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND A1_N a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR B1 a_420_387# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_481_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_110_47# Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y B2 a_481_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_110_427# A2_N a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_110_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR A1_N a_110_427# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
