* NGSPICE file created from sky130_fd_sc_lp__sdlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 VGND a_737_329# a_721_133# VNB nshort w=420000u l=150000u
+  ad=9.706e+11p pd=9.31e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_623_133# a_334_69# a_154_69# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.809e+11p ps=3.18e+06u
M1002 a_1231_367# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.656e+12p ps=1.346e+07u
M1003 VGND CLK a_254_357# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 a_334_69# a_254_357# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1005 GCLK a_1231_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1006 a_721_133# a_334_69# a_623_133# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.428e+11p ps=1.52e+06u
M1007 VPWR CLK a_254_357# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1008 VPWR a_737_329# a_1231_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_737_329# a_736_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 GCLK a_1231_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1011 a_154_69# SCE VGND VNB nshort w=420000u l=150000u
+  ad=2.457e+11p pd=2.85e+06u as=0p ps=0u
M1012 a_1194_52# CLK VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 a_1231_367# a_737_329# a_1194_52# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1014 a_737_329# a_623_133# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1015 a_154_69# GATE a_110_468# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1016 a_334_69# a_254_357# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1017 a_736_463# a_254_357# a_623_133# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND GATE a_154_69# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_623_133# a_254_357# a_154_69# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_110_468# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_737_329# a_623_133# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
.ends

