* File: sky130_fd_sc_lp__clkinvlp_16.pex.spice
* Created: Wed Sep  2 09:41:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINVLP_16%A 3 7 11 15 19 23 27 31 35 39 43 47 51
+ 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131 135 139
+ 141 143 145 172 206 211 224 230 237 238
c382 224 0 1.8905e-19 $X=5.04 $Y=1.295
c383 143 0 5.28023e-20 $X=8.475 $Y=2.48
c384 139 0 4.8318e-20 $X=7.945 $Y=0.61
c385 111 0 1.9352e-19 $X=6.365 $Y=0.61
c386 87 0 6.16522e-20 $X=5.215 $Y=0.61
c387 59 0 1.07873e-19 $X=3.635 $Y=0.61
c388 31 0 5.41591e-20 $X=2.055 $Y=0.61
r389 237 238 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=1.295
+ $X2=8.4 $Y2=1.295
r390 231 238 1.23188 $w=2.3e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=1.295
+ $X2=8.4 $Y2=1.295
r391 230 231 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.295
+ $X2=6.48 $Y2=1.295
r392 225 231 0.92391 $w=2.3e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=1.295
+ $X2=6.48 $Y2=1.295
r393 224 225 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r394 215 221 0.92391 $w=2.3e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=1.295
+ $X2=3.6 $Y2=1.295
r395 212 215 0.61594 $w=2.3e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=1.295
+ $X2=2.16 $Y2=1.295
r396 211 215 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.295
r397 211 212 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=1.295
+ $X2=1.2 $Y2=1.295
r398 207 212 0.61594 $w=2.3e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=1.295
+ $X2=1.2 $Y2=1.295
r399 206 207 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.295
r400 203 237 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.55
+ $Y=1.4 $X2=8.55 $Y2=1.4
r401 199 237 15.8648 $w=3.83e-07 $l=5.3e-07 $layer=LI1_cond $X=7.87 $Y=1.372
+ $X2=8.4 $Y2=1.372
r402 198 199 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.87
+ $Y=1.4 $X2=7.87 $Y2=1.4
r403 196 198 41.6273 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=7.585 $Y=1.407
+ $X2=7.87 $Y2=1.407
r404 190 192 37.9758 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=6.535 $Y=1.407
+ $X2=6.795 $Y2=1.407
r405 190 230 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.535
+ $Y=1.4 $X2=6.535 $Y2=1.4
r406 188 190 24.8303 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=6.365 $Y=1.407
+ $X2=6.535 $Y2=1.407
r407 182 224 1.73225 $w=7.23e-07 $l=1.05e-07 $layer=LI1_cond $X=5.017 $Y=1.4
+ $X2=5.017 $Y2=1.295
r408 181 182 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.215
+ $Y=1.4 $X2=5.215 $Y2=1.4
r409 179 181 62.8061 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.785 $Y=1.407
+ $X2=5.215 $Y2=1.407
r410 172 221 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=1.295
+ $X2=3.6 $Y2=1.295
r411 171 173 28.4818 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.44 $Y=1.407
+ $X2=3.635 $Y2=1.407
r412 171 172 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.4 $X2=3.44 $Y2=1.4
r413 169 171 34.3242 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.205 $Y=1.407
+ $X2=3.44 $Y2=1.407
r414 161 163 8.76364 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.995 $Y=1.407
+ $X2=2.055 $Y2=1.407
r415 159 161 54.0424 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.625 $Y=1.407
+ $X2=1.995 $Y2=1.407
r416 157 211 1.07647 $w=1.188e-06 $l=1.05e-07 $layer=LI1_cond $X=1.67 $Y=1.4
+ $X2=1.67 $Y2=1.295
r417 157 161 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.995
+ $Y=1.4 $X2=1.995 $Y2=1.4
r418 156 157 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.315
+ $Y=1.4 $X2=1.315 $Y2=1.4
r419 154 156 7.30303 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.265 $Y=1.407
+ $X2=1.315 $Y2=1.407
r420 151 152 45.2788 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.525 $Y=1.407
+ $X2=0.835 $Y2=1.407
r421 150 151 7.30303 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.407
+ $X2=0.525 $Y2=1.407
r422 148 150 22.6394 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.32 $Y=1.407
+ $X2=0.475 $Y2=1.407
r423 148 206 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.415 $X2=0.32 $Y2=1.415
r424 145 225 0.468371 $w=2.3e-07 $l=7.3e-07 $layer=MET1_cond $X=4.31 $Y=1.295
+ $X2=5.04 $Y2=1.295
r425 145 221 0.455539 $w=2.3e-07 $l=7.1e-07 $layer=MET1_cond $X=4.31 $Y=1.295
+ $X2=3.6 $Y2=1.295
r426 141 203 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.475 $Y=1.407
+ $X2=8.55 $Y2=1.407
r427 141 143 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=8.475 $Y=1.565
+ $X2=8.475 $Y2=2.48
r428 137 139 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=7.945 $Y=1.235
+ $X2=7.945 $Y2=0.61
r429 133 141 77.4121 $w=3.3e-07 $l=5.3e-07 $layer=POLY_cond $X=7.945 $Y=1.407
+ $X2=8.475 $Y2=1.407
r430 133 198 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.945 $Y=1.407
+ $X2=7.87 $Y2=1.407
r431 133 137 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=7.945 $Y=1.407
+ $X2=7.945 $Y2=1.235
r432 133 135 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=7.945 $Y=1.565
+ $X2=7.945 $Y2=2.48
r433 129 196 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=7.585 $Y=1.235
+ $X2=7.585 $Y2=1.407
r434 129 131 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=7.585 $Y=1.235
+ $X2=7.585 $Y2=0.61
r435 125 196 24.8303 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=7.415 $Y=1.407
+ $X2=7.585 $Y2=1.407
r436 125 194 37.9758 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=7.415 $Y=1.407
+ $X2=7.155 $Y2=1.407
r437 125 127 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=7.415 $Y=1.565
+ $X2=7.415 $Y2=2.48
r438 121 194 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=7.155 $Y=1.235
+ $X2=7.155 $Y2=1.407
r439 121 123 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=7.155 $Y=1.235
+ $X2=7.155 $Y2=0.61
r440 117 194 39.4364 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.885 $Y=1.407
+ $X2=7.155 $Y2=1.407
r441 117 192 13.1455 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.885 $Y=1.407
+ $X2=6.795 $Y2=1.407
r442 117 119 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=6.885 $Y=1.565
+ $X2=6.885 $Y2=2.48
r443 113 192 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=6.795 $Y=1.235
+ $X2=6.795 $Y2=1.407
r444 113 115 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=6.795 $Y=1.235
+ $X2=6.795 $Y2=0.61
r445 109 188 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=6.365 $Y=1.235
+ $X2=6.365 $Y2=1.407
r446 109 111 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=6.365 $Y=1.235
+ $X2=6.365 $Y2=0.61
r447 105 188 1.46061 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.355 $Y=1.407
+ $X2=6.365 $Y2=1.407
r448 105 186 51.1212 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=6.355 $Y=1.407
+ $X2=6.005 $Y2=1.407
r449 105 107 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=6.355 $Y=1.565
+ $X2=6.355 $Y2=2.48
r450 101 186 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=6.005 $Y=1.235
+ $X2=6.005 $Y2=1.407
r451 101 103 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=6.005 $Y=1.235
+ $X2=6.005 $Y2=0.61
r452 97 186 26.2909 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.825 $Y=1.407
+ $X2=6.005 $Y2=1.407
r453 97 184 36.5152 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.825 $Y=1.407
+ $X2=5.575 $Y2=1.407
r454 97 99 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=5.825 $Y=1.565
+ $X2=5.825 $Y2=2.48
r455 93 184 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=5.575 $Y=1.235
+ $X2=5.575 $Y2=1.407
r456 93 95 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=5.575 $Y=1.235
+ $X2=5.575 $Y2=0.61
r457 89 184 40.897 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=5.295 $Y=1.407
+ $X2=5.575 $Y2=1.407
r458 89 181 11.6848 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.295 $Y=1.407
+ $X2=5.215 $Y2=1.407
r459 89 91 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=5.295 $Y=1.565
+ $X2=5.295 $Y2=2.48
r460 85 181 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=5.215 $Y=1.235
+ $X2=5.215 $Y2=1.407
r461 85 87 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=5.215 $Y=1.235
+ $X2=5.215 $Y2=0.61
r462 81 179 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=4.785 $Y=1.235
+ $X2=4.785 $Y2=1.407
r463 81 83 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=4.785 $Y=1.235
+ $X2=4.785 $Y2=0.61
r464 77 179 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.765 $Y=1.407
+ $X2=4.785 $Y2=1.407
r465 77 177 49.6606 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.765 $Y=1.407
+ $X2=4.425 $Y2=1.407
r466 77 79 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=4.765 $Y=1.565
+ $X2=4.765 $Y2=2.48
r467 73 177 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=4.425 $Y=1.235
+ $X2=4.425 $Y2=1.407
r468 73 75 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=4.425 $Y=1.235
+ $X2=4.425 $Y2=0.61
r469 69 177 27.7515 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.235 $Y=1.407
+ $X2=4.425 $Y2=1.407
r470 69 175 35.0545 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.235 $Y=1.407
+ $X2=3.995 $Y2=1.407
r471 69 71 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=4.235 $Y=1.565
+ $X2=4.235 $Y2=2.48
r472 65 175 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=3.995 $Y=1.235
+ $X2=3.995 $Y2=1.407
r473 65 67 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=3.995 $Y=1.235
+ $X2=3.995 $Y2=0.61
r474 61 175 42.3576 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=3.705 $Y=1.407
+ $X2=3.995 $Y2=1.407
r475 61 173 10.2242 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.705 $Y=1.407
+ $X2=3.635 $Y2=1.407
r476 61 63 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.705 $Y=1.565
+ $X2=3.705 $Y2=2.48
r477 57 173 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=3.635 $Y=1.235
+ $X2=3.635 $Y2=1.407
r478 57 59 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=3.635 $Y=1.235
+ $X2=3.635 $Y2=0.61
r479 53 169 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=3.205 $Y=1.235
+ $X2=3.205 $Y2=1.407
r480 53 55 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=3.205 $Y=1.235
+ $X2=3.205 $Y2=0.61
r481 49 169 4.38182 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.175 $Y=1.407
+ $X2=3.205 $Y2=1.407
r482 49 167 48.2 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.175 $Y=1.407
+ $X2=2.845 $Y2=1.407
r483 49 51 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.175 $Y=1.565
+ $X2=3.175 $Y2=2.48
r484 45 167 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.845 $Y=1.235
+ $X2=2.845 $Y2=1.407
r485 45 47 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.845 $Y=1.235
+ $X2=2.845 $Y2=0.61
r486 41 167 29.2121 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.645 $Y=1.407
+ $X2=2.845 $Y2=1.407
r487 41 165 33.5939 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.645 $Y=1.407
+ $X2=2.415 $Y2=1.407
r488 41 43 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.645 $Y=1.565
+ $X2=2.645 $Y2=2.48
r489 37 165 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.415 $Y=1.235
+ $X2=2.415 $Y2=1.407
r490 37 39 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.415 $Y=1.235
+ $X2=2.415 $Y2=0.61
r491 33 165 43.8182 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.115 $Y=1.407
+ $X2=2.415 $Y2=1.407
r492 33 163 8.76364 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.115 $Y=1.407
+ $X2=2.055 $Y2=1.407
r493 33 35 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.115 $Y=1.565
+ $X2=2.115 $Y2=2.48
r494 29 163 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.055 $Y=1.235
+ $X2=2.055 $Y2=1.407
r495 29 31 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.055 $Y=1.235
+ $X2=2.055 $Y2=0.61
r496 25 159 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=1.407
r497 25 27 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=0.61
r498 21 159 5.84242 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.585 $Y=1.407
+ $X2=1.625 $Y2=1.407
r499 21 156 39.4364 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.585 $Y=1.407
+ $X2=1.315 $Y2=1.407
r500 21 23 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=1.585 $Y=1.565
+ $X2=1.585 $Y2=2.48
r501 17 154 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=1.407
r502 17 19 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=0.61
r503 13 154 30.6727 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.055 $Y=1.407
+ $X2=1.265 $Y2=1.407
r504 13 152 32.1333 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.055 $Y=1.407
+ $X2=0.835 $Y2=1.407
r505 13 15 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=2.48
r506 9 152 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=1.407
r507 9 11 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=0.61
r508 5 151 9.34494 $w=2.5e-07 $l=1.73e-07 $layer=POLY_cond $X=0.525 $Y=1.58
+ $X2=0.525 $Y2=1.407
r509 5 7 223.608 $w=2.5e-07 $l=9e-07 $layer=POLY_cond $X=0.525 $Y=1.58 $X2=0.525
+ $Y2=2.48
r510 1 150 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=1.407
r511 1 3 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_16%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 44 50
+ 56 62 66 70 76 80 82 87 88 90 91 93 94 95 104 108 117 125 128 131 134 138 146
c161 56 0 1.8905e-19 $X=4.5 $Y=2.125
r162 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r163 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r164 132 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r165 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r166 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r167 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r169 120 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r170 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r171 117 137 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.847 $Y2=3.33
r172 117 119 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.4 $Y2=3.33
r173 116 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r174 116 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r175 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r176 113 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=6.62 $Y2=3.33
r177 113 115 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=7.44 $Y2=3.33
r178 112 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r179 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r180 109 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=4.5 $Y2=3.33
r181 109 111 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=5.04 $Y2=3.33
r182 108 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.56 $Y2=3.33
r183 108 111 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.04 $Y2=3.33
r184 107 146 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.32 $Y2=3.33
r185 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r186 104 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.5 $Y2=3.33
r187 104 106 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.08 $Y2=3.33
r188 103 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r190 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r191 100 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r192 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r193 97 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.32 $Y2=3.33
r194 97 99 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r195 95 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r196 95 146 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.32 $Y2=3.33
r197 95 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r198 93 115 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.44 $Y2=3.33
r199 93 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.68 $Y2=3.33
r200 92 119 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.845 $Y=3.33
+ $X2=8.4 $Y2=3.33
r201 92 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.845 $Y=3.33
+ $X2=7.68 $Y2=3.33
r202 90 102 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r203 90 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.44 $Y2=3.33
r204 89 106 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.08 $Y2=3.33
r205 89 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.44 $Y2=3.33
r206 87 99 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.16 $Y2=3.33
r207 87 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.38 $Y2=3.33
r208 86 102 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=3.12 $Y2=3.33
r209 86 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.38 $Y2=3.33
r210 82 85 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.74 $Y=2.125
+ $X2=8.74 $Y2=2.835
r211 80 137 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=8.74 $Y=3.245
+ $X2=8.847 $Y2=3.33
r212 80 85 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=8.74 $Y=3.245
+ $X2=8.74 $Y2=2.835
r213 76 79 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.68 $Y=2.125
+ $X2=7.68 $Y2=2.835
r214 74 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.68 $Y=3.245
+ $X2=7.68 $Y2=3.33
r215 74 79 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.68 $Y=3.245
+ $X2=7.68 $Y2=2.835
r216 70 73 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.62 $Y=2.125
+ $X2=6.62 $Y2=2.835
r217 68 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.62 $Y=3.245
+ $X2=6.62 $Y2=3.33
r218 68 73 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.62 $Y=3.245
+ $X2=6.62 $Y2=2.835
r219 67 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=3.33
+ $X2=5.56 $Y2=3.33
r220 66 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=6.62 $Y2=3.33
r221 66 67 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=5.725 $Y2=3.33
r222 62 65 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=5.56 $Y=2.125
+ $X2=5.56 $Y2=2.835
r223 60 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=3.245
+ $X2=5.56 $Y2=3.33
r224 60 65 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.56 $Y=3.245
+ $X2=5.56 $Y2=2.835
r225 56 59 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.5 $Y=2.125 $X2=4.5
+ $Y2=2.835
r226 54 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=3.245
+ $X2=4.5 $Y2=3.33
r227 54 59 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.5 $Y=3.245
+ $X2=4.5 $Y2=2.835
r228 50 53 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.44 $Y=2.125
+ $X2=3.44 $Y2=2.835
r229 48 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=3.33
r230 48 53 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.835
r231 44 47 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.38 $Y=2.125
+ $X2=2.38 $Y2=2.835
r232 42 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r233 42 47 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.835
r234 38 41 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.32 $Y=2.125
+ $X2=1.32 $Y2=2.835
r235 36 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=3.33
r236 36 41 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=2.835
r237 35 122 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r238 34 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.32 $Y2=3.33
r239 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.425 $Y2=3.33
r240 30 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.26 $Y=2.125
+ $X2=0.26 $Y2=2.835
r241 28 122 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r242 28 33 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.835
r243 9 85 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.6
+ $Y=1.98 $X2=8.74 $Y2=2.835
r244 9 82 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.6
+ $Y=1.98 $X2=8.74 $Y2=2.125
r245 8 79 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.98 $X2=7.68 $Y2=2.835
r246 8 76 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.98 $X2=7.68 $Y2=2.125
r247 7 73 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.98 $X2=6.62 $Y2=2.835
r248 7 70 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.98 $X2=6.62 $Y2=2.125
r249 6 65 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.98 $X2=5.56 $Y2=2.835
r250 6 62 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.98 $X2=5.56 $Y2=2.125
r251 5 59 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=1.98 $X2=4.5 $Y2=2.835
r252 5 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=1.98 $X2=4.5 $Y2=2.125
r253 4 53 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.98 $X2=3.44 $Y2=2.835
r254 4 50 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.98 $X2=3.44 $Y2=2.125
r255 3 47 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.98 $X2=2.38 $Y2=2.835
r256 3 44 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.98 $X2=2.38 $Y2=2.125
r257 2 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.98 $X2=1.32 $Y2=2.835
r258 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.98 $X2=1.32 $Y2=2.125
r259 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.98 $X2=0.26 $Y2=2.835
r260 1 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.98 $X2=0.26 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 40 44 50
+ 54 60 66 70 71 74 77 78 80 83 88 90 93 100 108 115 122 130 137 138 145 147
c244 138 0 5.28023e-20 $X=8.21 $Y=2.035
c245 88 0 4.8318e-20 $X=7.37 $Y=1.38
c246 83 0 2.55172e-19 $X=6.042 $Y=1.38
c247 80 0 1.07873e-19 $X=4.127 $Y=1.565
c248 74 0 5.41591e-20 $X=2.91 $Y=1.38
r249 145 147 5.53173 $w=3.58e-07 $l=1.6e-07 $layer=LI1_cond $X=6.075 $Y=2.035
+ $X2=6.075 $Y2=1.875
r250 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=2.035 $X2=6
+ $Y2=2.035
r251 137 142 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=8.21 $Y=2.035
+ $X2=8.21 $Y2=2.835
r252 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.21 $Y=2.035
+ $X2=8.21 $Y2=2.035
r253 131 138 0.680101 $w=2.3e-07 $l=1.06e-06 $layer=MET1_cond $X=7.15 $Y=2.035
+ $X2=8.21 $Y2=2.035
r254 131 146 0.737845 $w=2.3e-07 $l=1.15e-06 $layer=MET1_cond $X=7.15 $Y=2.035
+ $X2=6 $Y2=2.035
r255 130 134 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=7.15 $Y=2.035
+ $X2=7.15 $Y2=2.835
r256 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.15 $Y=2.035
+ $X2=7.15 $Y2=2.035
r257 123 146 0.61594 $w=2.3e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=2.035
+ $X2=6 $Y2=2.035
r258 122 127 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=5.03 $Y=2.035
+ $X2=5.03 $Y2=2.835
r259 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r260 115 119 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=3.97 $Y=2.035
+ $X2=3.97 $Y2=2.835
r261 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.97 $Y=2.035
+ $X2=3.97 $Y2=2.035
r262 109 116 0.680101 $w=2.3e-07 $l=1.06e-06 $layer=MET1_cond $X=2.91 $Y=2.035
+ $X2=3.97 $Y2=2.035
r263 108 112 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=2.91 $Y=2.035
+ $X2=2.91 $Y2=2.835
r264 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.91 $Y=2.035
+ $X2=2.91 $Y2=2.035
r265 101 109 0.680101 $w=2.3e-07 $l=1.06e-06 $layer=MET1_cond $X=1.85 $Y=2.035
+ $X2=2.91 $Y2=2.035
r266 100 105 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=1.85 $Y=2.035
+ $X2=1.85 $Y2=2.835
r267 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.85 $Y=2.035
+ $X2=1.85 $Y2=2.035
r268 94 101 0.725013 $w=2.3e-07 $l=1.13e-06 $layer=MET1_cond $X=0.72 $Y=2.035
+ $X2=1.85 $Y2=2.035
r269 93 97 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=0.79 $Y=2.035 $X2=0.79
+ $Y2=2.835
r270 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.035
r271 90 123 0.368923 $w=2.3e-07 $l=5.75e-07 $layer=MET1_cond $X=4.465 $Y=2.035
+ $X2=5.04 $Y2=2.035
r272 90 116 0.317594 $w=2.3e-07 $l=4.95e-07 $layer=MET1_cond $X=4.465 $Y=2.035
+ $X2=3.97 $Y2=2.035
r273 86 130 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=7.15 $Y=1.565
+ $X2=7.15 $Y2=2.035
r274 85 88 6.85236 $w=3.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.15 $Y=1.38
+ $X2=7.37 $Y2=1.38
r275 85 86 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=7.15 $Y=1.38
+ $X2=7.15 $Y2=1.565
r276 81 83 7.84907 $w=3.68e-07 $l=2.52e-07 $layer=LI1_cond $X=5.79 $Y=1.38
+ $X2=6.042 $Y2=1.38
r277 79 80 13.5466 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.127 $Y=1.195
+ $X2=4.127 $Y2=1.565
r278 78 80 10.8465 $w=2.53e-07 $l=2.4e-07 $layer=LI1_cond $X=4.007 $Y=1.805
+ $X2=4.007 $Y2=1.565
r279 77 115 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.97 $Y=1.97
+ $X2=3.97 $Y2=2.035
r280 77 78 6.3875 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=1.97
+ $X2=3.97 $Y2=1.805
r281 75 108 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.91 $Y=1.565
+ $X2=2.91 $Y2=2.035
r282 74 75 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=2.91 $Y=1.38
+ $X2=2.91 $Y2=1.565
r283 72 74 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.63 $Y=1.38
+ $X2=2.91 $Y2=1.38
r284 70 93 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.79 $Y=1.9
+ $X2=0.79 $Y2=2.035
r285 70 71 6.05995 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=1.9
+ $X2=0.79 $Y2=1.735
r286 64 88 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=7.37 $Y=1.195
+ $X2=7.37 $Y2=1.38
r287 64 66 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=7.37 $Y=1.195
+ $X2=7.37 $Y2=0.61
r288 60 62 22.7287 $w=3.58e-07 $l=7.1e-07 $layer=LI1_cond $X=6.075 $Y=2.125
+ $X2=6.075 $Y2=2.835
r289 58 145 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=6.075 $Y=2.055
+ $X2=6.075 $Y2=2.035
r290 58 60 2.24086 $w=3.58e-07 $l=7e-08 $layer=LI1_cond $X=6.075 $Y=2.055
+ $X2=6.075 $Y2=2.125
r291 56 83 2.08285 $w=2.95e-07 $l=1.85e-07 $layer=LI1_cond $X=6.042 $Y=1.565
+ $X2=6.042 $Y2=1.38
r292 56 147 12.1104 $w=2.93e-07 $l=3.1e-07 $layer=LI1_cond $X=6.042 $Y=1.565
+ $X2=6.042 $Y2=1.875
r293 52 81 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=5.79 $Y=1.195
+ $X2=5.79 $Y2=1.38
r294 52 54 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=5.79 $Y=1.195
+ $X2=5.79 $Y2=0.61
r295 50 79 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=4.21 $Y=0.61
+ $X2=4.21 $Y2=1.195
r296 42 72 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=2.63 $Y=1.195
+ $X2=2.63 $Y2=1.38
r297 42 44 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.63 $Y=1.195
+ $X2=2.63 $Y2=0.61
r298 40 69 13.6575 $w=5.03e-07 $l=5.36936e-07 $layer=LI1_cond $X=0.765 $Y=1.01
+ $X2=0.92 $Y2=0.545
r299 40 71 29.84 $w=2.78e-07 $l=7.25e-07 $layer=LI1_cond $X=0.765 $Y=1.01
+ $X2=0.765 $Y2=1.735
r300 13 142 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.98 $X2=8.21 $Y2=2.835
r301 13 137 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=1.98 $X2=8.21 $Y2=2.125
r302 12 134 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.01
+ $Y=1.98 $X2=7.15 $Y2=2.835
r303 12 130 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.01
+ $Y=1.98 $X2=7.15 $Y2=2.125
r304 11 62 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=5.95
+ $Y=1.98 $X2=6.09 $Y2=2.835
r305 11 60 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.95
+ $Y=1.98 $X2=6.09 $Y2=2.125
r306 10 127 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.98 $X2=5.03 $Y2=2.835
r307 10 122 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.98 $X2=5.03 $Y2=2.125
r308 9 119 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.98 $X2=3.97 $Y2=2.835
r309 9 115 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.98 $X2=3.97 $Y2=2.125
r310 8 112 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.98 $X2=2.91 $Y2=2.835
r311 8 108 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.98 $X2=2.91 $Y2=2.125
r312 7 105 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.98 $X2=1.85 $Y2=2.835
r313 7 100 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.98 $X2=1.85 $Y2=2.125
r314 6 97 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.98 $X2=0.79 $Y2=2.835
r315 6 93 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.98 $X2=0.79 $Y2=2.125
r316 5 66 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=7.23
+ $Y=0.335 $X2=7.37 $Y2=0.61
r317 4 54 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.65
+ $Y=0.335 $X2=5.79 $Y2=0.61
r318 3 50 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.07
+ $Y=0.335 $X2=4.21 $Y2=0.61
r319 2 44 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.335 $X2=2.63 $Y2=0.61
r320 1 69 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.335 $X2=1.05 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_16%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44
+ 45 47 48 49 51 63 70 83 84 90 93 96 106
r117 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r118 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r119 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r120 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r121 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r122 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r123 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r124 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r125 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r126 77 80 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r127 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r128 75 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.745 $Y=0 $X2=6.58
+ $Y2=0
r129 75 77 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.96 $Y2=0
r130 74 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r131 74 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r132 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r133 71 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r134 71 73 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r135 70 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=0 $X2=6.58
+ $Y2=0
r136 70 73 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=6.415 $Y=0
+ $X2=5.52 $Y2=0
r137 66 106 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.32
+ $Y2=0
r138 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r139 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r140 63 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r141 63 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.56 $Y2=0
r142 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r143 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r144 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r145 59 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r146 58 61 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r147 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r148 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.84
+ $Y2=0
r149 56 58 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.16 $Y2=0
r150 55 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r151 55 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r152 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r153 52 87 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r154 52 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r155 51 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.84
+ $Y2=0
r156 51 54 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.675 $Y=0
+ $X2=0.72 $Y2=0
r157 49 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r158 49 106 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.32 $Y2=0
r159 49 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r160 47 80 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.995 $Y=0 $X2=7.92
+ $Y2=0
r161 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=8.16
+ $Y2=0
r162 46 83 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.88 $Y2=0
r163 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.325 $Y=0 $X2=8.16
+ $Y2=0
r164 44 61 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0
+ $X2=3.12 $Y2=0
r165 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r166 43 65 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.6
+ $Y2=0
r167 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r168 39 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.16 $Y=0.085
+ $X2=8.16 $Y2=0
r169 39 41 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=8.16 $Y=0.085
+ $X2=8.16 $Y2=0.61
r170 35 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0
r171 35 37 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0.61
r172 31 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r173 31 33 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.61
r174 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r175 27 29 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.61
r176 23 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r177 23 25 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.61
r178 19 87 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r179 19 21 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.61
r180 6 41 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=8.02
+ $Y=0.335 $X2=8.16 $Y2=0.61
r181 5 37 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=6.44
+ $Y=0.335 $X2=6.58 $Y2=0.61
r182 4 33 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.335 $X2=5 $Y2=0.61
r183 3 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.335 $X2=3.42 $Y2=0.61
r184 2 25 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.335 $X2=1.84 $Y2=0.61
r185 1 21 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.335 $X2=0.26 $Y2=0.61
.ends

