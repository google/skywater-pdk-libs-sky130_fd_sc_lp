# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxtp_lp2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dlxtp_lp2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 0.905000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.460000 0.440000 8.050000 2.925000 ;
        RECT 7.720000 0.395000 8.050000 0.440000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.175000 1.380000 1.845000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.265000 0.445000 0.725000 ;
      RECT 0.115000  0.725000 0.285000 2.025000 ;
      RECT 0.115000  2.025000 0.445000 2.455000 ;
      RECT 0.115000  2.455000 1.325000 2.585000 ;
      RECT 0.115000  2.585000 3.650000 2.625000 ;
      RECT 0.115000  2.625000 0.445000 3.065000 ;
      RECT 0.645000  2.805000 0.975000 3.245000 ;
      RECT 0.905000  0.085000 1.235000 0.725000 ;
      RECT 1.155000  2.625000 3.650000 2.755000 ;
      RECT 1.175000  2.025000 2.025000 2.275000 ;
      RECT 1.695000  0.265000 2.025000 2.025000 ;
      RECT 2.240000  0.265000 2.585000 0.915000 ;
      RECT 2.240000  0.915000 4.880000 1.085000 ;
      RECT 2.240000  1.085000 2.570000 2.405000 ;
      RECT 2.750000  1.265000 4.400000 1.435000 ;
      RECT 2.750000  1.435000 3.080000 1.935000 ;
      RECT 2.850000  2.935000 3.180000 3.245000 ;
      RECT 3.045000  0.085000 3.375000 0.675000 ;
      RECT 3.320000  1.615000 3.650000 2.585000 ;
      RECT 3.710000  0.765000 4.880000 0.915000 ;
      RECT 3.945000  0.295000 5.230000 0.585000 ;
      RECT 4.070000  1.435000 4.400000 1.665000 ;
      RECT 4.305000  2.075000 5.230000 2.245000 ;
      RECT 4.305000  2.245000 4.635000 3.065000 ;
      RECT 4.610000  1.085000 4.880000 1.895000 ;
      RECT 5.060000  0.585000 5.230000 0.855000 ;
      RECT 5.060000  0.855000 6.215000 1.025000 ;
      RECT 5.060000  1.025000 5.230000 2.075000 ;
      RECT 5.410000  0.085000 5.740000 0.675000 ;
      RECT 5.410000  1.205000 5.675000 1.705000 ;
      RECT 5.410000  1.705000 6.565000 1.875000 ;
      RECT 5.410000  2.075000 5.740000 3.245000 ;
      RECT 5.885000  1.025000 6.215000 1.525000 ;
      RECT 6.140000  2.075000 6.565000 3.065000 ;
      RECT 6.370000  0.265000 6.700000 0.675000 ;
      RECT 6.395000  0.675000 6.700000 1.035000 ;
      RECT 6.395000  1.035000 6.965000 1.705000 ;
      RECT 6.395000  1.875000 6.565000 2.075000 ;
      RECT 6.930000  0.085000 7.260000 0.855000 ;
      RECT 6.930000  1.885000 7.260000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__dlxtp_lp2
END LIBRARY
