* File: sky130_fd_sc_lp__a221o_m.pxi.spice
* Created: Wed Sep  2 09:21:36 2020
* 
x_PM_SKY130_FD_SC_LP__A221O_M%A_33_153# N_A_33_153#_M1008_d N_A_33_153#_M1011_d
+ N_A_33_153#_M1009_d N_A_33_153#_c_79_n N_A_33_153#_M1004_g N_A_33_153#_M1002_g
+ N_A_33_153#_c_80_n N_A_33_153#_c_90_n N_A_33_153#_c_81_n N_A_33_153#_c_117_p
+ N_A_33_153#_c_82_n N_A_33_153#_c_83_n N_A_33_153#_c_84_n N_A_33_153#_c_92_n
+ N_A_33_153#_c_93_n N_A_33_153#_c_85_n N_A_33_153#_c_86_n N_A_33_153#_c_87_n
+ N_A_33_153#_c_88_n PM_SKY130_FD_SC_LP__A221O_M%A_33_153#
x_PM_SKY130_FD_SC_LP__A221O_M%A2 N_A2_M1007_g N_A2_M1010_g A2 A2 N_A2_c_194_n
+ PM_SKY130_FD_SC_LP__A221O_M%A2
x_PM_SKY130_FD_SC_LP__A221O_M%A1 N_A1_c_239_n N_A1_M1008_g N_A1_M1000_g A1 A1
+ N_A1_c_242_n PM_SKY130_FD_SC_LP__A221O_M%A1
x_PM_SKY130_FD_SC_LP__A221O_M%B1 N_B1_M1005_g N_B1_M1006_g B1 N_B1_c_288_n
+ PM_SKY130_FD_SC_LP__A221O_M%B1
x_PM_SKY130_FD_SC_LP__A221O_M%B2 N_B2_c_324_n N_B2_M1003_g N_B2_M1001_g
+ N_B2_c_325_n N_B2_c_326_n N_B2_c_332_n B2 N_B2_c_328_n N_B2_c_329_n
+ PM_SKY130_FD_SC_LP__A221O_M%B2
x_PM_SKY130_FD_SC_LP__A221O_M%C1 N_C1_c_373_n N_C1_M1011_g N_C1_M1009_g
+ N_C1_c_374_n N_C1_c_375_n N_C1_c_378_n C1 C1 N_C1_c_380_n
+ PM_SKY130_FD_SC_LP__A221O_M%C1
x_PM_SKY130_FD_SC_LP__A221O_M%X N_X_M1004_s N_X_M1002_s X X X X X X X
+ N_X_c_414_n PM_SKY130_FD_SC_LP__A221O_M%X
x_PM_SKY130_FD_SC_LP__A221O_M%VPWR N_VPWR_M1002_d N_VPWR_M1000_d N_VPWR_c_438_n
+ N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n VPWR N_VPWR_c_442_n
+ N_VPWR_c_443_n N_VPWR_c_437_n N_VPWR_c_445_n PM_SKY130_FD_SC_LP__A221O_M%VPWR
x_PM_SKY130_FD_SC_LP__A221O_M%A_233_535# N_A_233_535#_M1010_d
+ N_A_233_535#_M1006_d N_A_233_535#_c_476_n N_A_233_535#_c_472_n
+ N_A_233_535#_c_473_n N_A_233_535#_c_474_n
+ PM_SKY130_FD_SC_LP__A221O_M%A_233_535#
x_PM_SKY130_FD_SC_LP__A221O_M%A_337_397# N_A_337_397#_M1006_s
+ N_A_337_397#_M1001_d N_A_337_397#_c_495_n N_A_337_397#_c_496_n
+ N_A_337_397#_c_497_n N_A_337_397#_c_498_n
+ PM_SKY130_FD_SC_LP__A221O_M%A_337_397#
x_PM_SKY130_FD_SC_LP__A221O_M%VGND N_VGND_M1004_d N_VGND_M1003_d N_VGND_c_522_n
+ N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n VGND N_VGND_c_526_n
+ N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n PM_SKY130_FD_SC_LP__A221O_M%VGND
cc_1 VNB N_A_33_153#_c_79_n 0.0192606f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_2 VNB N_A_33_153#_c_80_n 0.0319856f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_3 VNB N_A_33_153#_c_81_n 0.0193364f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.48
cc_4 VNB N_A_33_153#_c_82_n 0.0101614f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.395
cc_5 VNB N_A_33_153#_c_83_n 0.0130002f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=0.75
cc_6 VNB N_A_33_153#_c_84_n 0.0373854f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=2.13
cc_7 VNB N_A_33_153#_c_85_n 0.00237091f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.48
cc_8 VNB N_A_33_153#_c_86_n 0.00210752f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.75
cc_9 VNB N_A_33_153#_c_87_n 0.0166521f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.51
cc_10 VNB N_A_33_153#_c_88_n 0.0426912f $X=-0.19 $Y=-0.245 $X2=0.47 $Y2=1.695
cc_11 VNB N_A2_M1007_g 0.0373876f $X=-0.19 $Y=-0.245 $X2=2.96 $Y2=1.985
cc_12 VNB N_A2_M1010_g 0.00974066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A2 0.0090795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_194_n 0.0570985f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.885
cc_15 VNB N_A1_c_239_n 0.016341f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.235
cc_16 VNB N_A1_M1000_g 0.0297364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A1 0.00808717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_242_n 0.0394344f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.885
cc_19 VNB N_B1_M1005_g 0.0371047f $X=-0.19 $Y=-0.245 $X2=2.96 $Y2=1.985
cc_20 VNB N_B1_M1006_g 0.00990908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB B1 0.00306009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_288_n 0.034585f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_23 VNB N_B2_c_324_n 0.0157999f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.235
cc_24 VNB N_B2_c_325_n 0.0270519f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_25 VNB N_B2_c_326_n 0.010326f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.885
cc_26 VNB B2 0.00256734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B2_c_328_n 0.0298736f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_28 VNB N_B2_c_329_n 0.0155313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C1_c_373_n 0.0209741f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.235
cc_30 VNB N_C1_c_374_n 0.0422065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C1_c_375_n 0.0289772f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_32 VNB X 0.042507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_437_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.395
cc_34 VNB N_VGND_c_522_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_523_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_36 VNB N_VGND_c_524_n 0.0391189f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.885
cc_37 VNB N_VGND_c_525_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.885
cc_38 VNB N_VGND_c_526_n 0.0163199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_527_n 0.0210426f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=0.835
cc_40 VNB N_VGND_c_528_n 0.190785f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.395
cc_41 VNB N_VGND_c_529_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=0.835
cc_42 VPB N_A_33_153#_M1002_g 0.0313352f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.885
cc_43 VPB N_A_33_153#_c_90_n 0.00950519f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.78
cc_44 VPB N_A_33_153#_c_84_n 0.0255469f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=2.13
cc_45 VPB N_A_33_153#_c_92_n 0.00421235f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.86
cc_46 VPB N_A_33_153#_c_93_n 0.102127f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.86
cc_47 VPB N_A_33_153#_c_85_n 0.00213358f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.48
cc_48 VPB N_A_33_153#_c_88_n 0.00173387f $X=-0.19 $Y=1.655 $X2=0.47 $Y2=1.695
cc_49 VPB N_A2_M1010_g 0.0642455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A1_M1000_g 0.0701669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B1_M1006_g 0.0280439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_B2_M1001_g 0.0199932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B2_c_326_n 0.00247588f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.885
cc_54 VPB N_B2_c_332_n 0.0119057f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.885
cc_55 VPB N_C1_M1009_g 0.0352824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_C1_c_374_n 0.00306762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_C1_c_378_n 0.0283266f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.885
cc_58 VPB C1 0.0374604f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=0.84
cc_59 VPB N_C1_c_380_n 0.0446672f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.78
cc_60 VPB X 0.0395852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_X_c_414_n 0.0188832f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.78
cc_62 VPB N_VPWR_c_438_n 0.00432637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_439_n 0.00789712f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_64 VPB N_VPWR_c_440_n 0.0235313f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.885
cc_65 VPB N_VPWR_c_441_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.885
cc_66 VPB N_VPWR_c_442_n 0.0154194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_443_n 0.0404331f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=0.835
cc_68 VPB N_VPWR_c_437_n 0.0664491f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=1.395
cc_69 VPB N_VPWR_c_445_n 0.00510247f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=0.835
cc_70 VPB N_A_233_535#_c_472_n 0.0207741f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.695
cc_71 VPB N_A_233_535#_c_473_n 0.00957895f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_72 VPB N_A_233_535#_c_474_n 0.00184352f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.365
cc_73 VPB N_A_337_397#_c_495_n 0.00139403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_337_397#_c_496_n 0.014756f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.695
cc_75 VPB N_A_337_397#_c_497_n 0.00586694f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_76 VPB N_A_337_397#_c_498_n 0.00103653f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.365
cc_77 N_A_33_153#_c_79_n N_A2_M1007_g 0.0201937f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_78 N_A_33_153#_c_88_n N_A2_M1007_g 0.00238033f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_79 N_A_33_153#_M1002_g N_A2_M1010_g 0.0238008f $X=0.66 $Y=2.885 $X2=0 $Y2=0
cc_80 N_A_33_153#_c_90_n N_A2_M1010_g 4.00469e-19 $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_81 N_A_33_153#_c_81_n N_A2_M1010_g 0.00167166f $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_82 N_A_33_153#_c_92_n N_A2_M1010_g 0.00273792f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_83 N_A_33_153#_c_93_n N_A2_M1010_g 0.0392983f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_84 N_A_33_153#_c_85_n N_A2_M1010_g 0.0189694f $X=1.07 $Y=1.48 $X2=0 $Y2=0
cc_85 N_A_33_153#_c_88_n N_A2_M1010_g 0.00115135f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_86 N_A_33_153#_c_80_n A2 6.8402e-19 $X=0.475 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A_33_153#_c_90_n A2 0.0070566f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_88 N_A_33_153#_c_92_n A2 0.00418826f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_89 N_A_33_153#_c_93_n A2 3.93723e-19 $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_90 N_A_33_153#_c_85_n A2 0.00582693f $X=1.07 $Y=1.48 $X2=0 $Y2=0
cc_91 N_A_33_153#_c_88_n A2 9.12968e-19 $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_92 N_A_33_153#_c_90_n N_A2_c_194_n 0.00735965f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_93 N_A_33_153#_c_81_n N_A2_c_194_n 0.00179395f $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_94 N_A_33_153#_c_92_n N_A2_c_194_n 6.47257e-19 $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_95 N_A_33_153#_c_93_n N_A2_c_194_n 0.0142818f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_96 N_A_33_153#_c_85_n N_A2_c_194_n 0.00938108f $X=1.07 $Y=1.48 $X2=0 $Y2=0
cc_97 N_A_33_153#_c_88_n N_A2_c_194_n 0.0179931f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_98 N_A_33_153#_c_117_p N_A1_c_239_n 0.00312784f $X=1.705 $Y=0.51 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_33_153#_c_86_n N_A1_c_239_n 3.68224e-19 $X=1.715 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_33_153#_c_81_n N_A1_M1000_g 0.0188418f $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_101 N_A_33_153#_c_85_n N_A1_M1000_g 0.00168292f $X=1.07 $Y=1.48 $X2=0 $Y2=0
cc_102 N_A_33_153#_M1008_d A1 0.00237889f $X=1.34 $Y=0.235 $X2=0 $Y2=0
cc_103 N_A_33_153#_c_81_n A1 0.0148315f $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_104 N_A_33_153#_c_117_p A1 0.0143718f $X=1.705 $Y=0.51 $X2=0 $Y2=0
cc_105 N_A_33_153#_c_82_n A1 0.0186556f $X=1.705 $Y=1.395 $X2=0 $Y2=0
cc_106 N_A_33_153#_c_85_n A1 0.00214118f $X=1.07 $Y=1.48 $X2=0 $Y2=0
cc_107 N_A_33_153#_c_86_n A1 0.0141319f $X=1.715 $Y=0.75 $X2=0 $Y2=0
cc_108 N_A_33_153#_c_81_n N_A1_c_242_n 0.00174306f $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_109 N_A_33_153#_c_82_n N_A1_c_242_n 0.00941744f $X=1.705 $Y=1.395 $X2=0 $Y2=0
cc_110 N_A_33_153#_c_86_n N_A1_c_242_n 6.60269e-19 $X=1.715 $Y=0.75 $X2=0 $Y2=0
cc_111 N_A_33_153#_c_117_p N_B1_M1005_g 2.36833e-19 $X=1.705 $Y=0.51 $X2=0 $Y2=0
cc_112 N_A_33_153#_c_82_n N_B1_M1005_g 0.00932327f $X=1.705 $Y=1.395 $X2=0 $Y2=0
cc_113 N_A_33_153#_c_83_n N_B1_M1005_g 0.0151836f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_114 N_A_33_153#_c_81_n N_B1_M1006_g 0.00223406f $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_115 N_A_33_153#_c_81_n B1 0.00709266f $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_116 N_A_33_153#_c_82_n B1 0.0170107f $X=1.705 $Y=1.395 $X2=0 $Y2=0
cc_117 N_A_33_153#_c_83_n B1 0.0127503f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_118 N_A_33_153#_c_81_n N_B1_c_288_n 7.99853e-19 $X=1.62 $Y=1.48 $X2=0 $Y2=0
cc_119 N_A_33_153#_c_83_n N_B1_c_288_n 0.00463618f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_120 N_A_33_153#_c_83_n N_B2_c_324_n 0.00714485f $X=2.915 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_33_153#_c_87_n N_B2_c_324_n 6.42446e-19 $X=3.08 $Y=0.51 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_33_153#_c_83_n N_B2_c_325_n 0.0178779f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_123 N_A_33_153#_c_84_n N_B2_c_325_n 3.72317e-19 $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_124 N_A_33_153#_c_84_n N_B2_c_326_n 0.00515217f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_125 N_A_33_153#_c_83_n B2 0.012657f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_126 N_A_33_153#_c_84_n B2 0.0117755f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_127 N_A_33_153#_c_83_n N_B2_c_328_n 0.00370862f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_128 N_A_33_153#_c_84_n N_B2_c_328_n 0.0035129f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_129 N_A_33_153#_c_84_n N_B2_c_329_n 0.00512563f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_130 N_A_33_153#_c_83_n N_C1_c_373_n 0.00601136f $X=2.915 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_33_153#_c_87_n N_C1_c_373_n 0.00776354f $X=3.08 $Y=0.51 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_33_153#_c_84_n N_C1_M1009_g 0.00256993f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_133 N_A_33_153#_c_84_n N_C1_c_374_n 0.0268226f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_134 N_A_33_153#_c_83_n N_C1_c_375_n 0.00634747f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_135 N_A_33_153#_c_84_n N_C1_c_375_n 0.00369048f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_136 N_A_33_153#_c_87_n N_C1_c_375_n 0.0105901f $X=3.08 $Y=0.51 $X2=0 $Y2=0
cc_137 N_A_33_153#_c_84_n N_C1_c_378_n 0.0095267f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_138 N_A_33_153#_c_84_n C1 0.00950954f $X=3.1 $Y=2.13 $X2=0 $Y2=0
cc_139 N_A_33_153#_c_79_n X 0.00428617f $X=0.475 $Y=0.765 $X2=0 $Y2=0
cc_140 N_A_33_153#_M1002_g X 0.00931507f $X=0.66 $Y=2.885 $X2=0 $Y2=0
cc_141 N_A_33_153#_c_80_n X 0.0113996f $X=0.475 $Y=0.84 $X2=0 $Y2=0
cc_142 N_A_33_153#_c_92_n X 0.0446903f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_143 N_A_33_153#_c_93_n X 0.0341779f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_144 N_A_33_153#_c_85_n X 0.00635638f $X=1.07 $Y=1.48 $X2=0 $Y2=0
cc_145 N_A_33_153#_c_88_n X 0.0253171f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_146 N_A_33_153#_M1002_g N_X_c_414_n 5.68606e-19 $X=0.66 $Y=2.885 $X2=0 $Y2=0
cc_147 N_A_33_153#_c_92_n N_X_c_414_n 0.00134781f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_148 N_A_33_153#_c_93_n N_X_c_414_n 0.00781211f $X=0.61 $Y=1.86 $X2=0 $Y2=0
cc_149 N_A_33_153#_M1002_g N_VPWR_c_438_n 0.00288714f $X=0.66 $Y=2.885 $X2=0
+ $Y2=0
cc_150 N_A_33_153#_M1002_g N_VPWR_c_440_n 0.00585385f $X=0.66 $Y=2.885 $X2=0
+ $Y2=0
cc_151 N_A_33_153#_M1002_g N_VPWR_c_437_n 0.0118727f $X=0.66 $Y=2.885 $X2=0
+ $Y2=0
cc_152 N_A_33_153#_c_84_n N_A_337_397#_c_496_n 0.0117604f $X=3.1 $Y=2.13 $X2=0
+ $Y2=0
cc_153 N_A_33_153#_c_81_n N_A_337_397#_c_497_n 0.00752735f $X=1.62 $Y=1.48 $X2=0
+ $Y2=0
cc_154 N_A_33_153#_c_85_n N_A_337_397#_c_497_n 0.00399561f $X=1.07 $Y=1.48 $X2=0
+ $Y2=0
cc_155 N_A_33_153#_c_84_n N_A_337_397#_c_498_n 0.00450152f $X=3.1 $Y=2.13 $X2=0
+ $Y2=0
cc_156 N_A_33_153#_c_79_n N_VGND_c_522_n 0.0119058f $X=0.475 $Y=0.765 $X2=0
+ $Y2=0
cc_157 N_A_33_153#_c_83_n N_VGND_c_523_n 0.0218188f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_158 N_A_33_153#_c_87_n N_VGND_c_523_n 0.00455041f $X=3.08 $Y=0.51 $X2=0 $Y2=0
cc_159 N_A_33_153#_c_117_p N_VGND_c_524_n 0.00789274f $X=1.705 $Y=0.51 $X2=0
+ $Y2=0
cc_160 N_A_33_153#_c_83_n N_VGND_c_524_n 0.00837164f $X=2.915 $Y=0.75 $X2=0
+ $Y2=0
cc_161 N_A_33_153#_c_79_n N_VGND_c_526_n 0.00486043f $X=0.475 $Y=0.765 $X2=0
+ $Y2=0
cc_162 N_A_33_153#_c_80_n N_VGND_c_526_n 0.00129882f $X=0.475 $Y=0.84 $X2=0
+ $Y2=0
cc_163 N_A_33_153#_c_83_n N_VGND_c_527_n 0.00412321f $X=2.915 $Y=0.75 $X2=0
+ $Y2=0
cc_164 N_A_33_153#_c_87_n N_VGND_c_527_n 0.010639f $X=3.08 $Y=0.51 $X2=0 $Y2=0
cc_165 N_A_33_153#_M1008_d N_VGND_c_528_n 0.00717444f $X=1.34 $Y=0.235 $X2=0
+ $Y2=0
cc_166 N_A_33_153#_M1011_d N_VGND_c_528_n 0.00235821f $X=2.94 $Y=0.235 $X2=0
+ $Y2=0
cc_167 N_A_33_153#_c_79_n N_VGND_c_528_n 0.0093594f $X=0.475 $Y=0.765 $X2=0
+ $Y2=0
cc_168 N_A_33_153#_c_80_n N_VGND_c_528_n 0.00119216f $X=0.475 $Y=0.84 $X2=0
+ $Y2=0
cc_169 N_A_33_153#_c_117_p N_VGND_c_528_n 0.00695668f $X=1.705 $Y=0.51 $X2=0
+ $Y2=0
cc_170 N_A_33_153#_c_83_n N_VGND_c_528_n 0.0211166f $X=2.915 $Y=0.75 $X2=0 $Y2=0
cc_171 N_A_33_153#_c_87_n N_VGND_c_528_n 0.011528f $X=3.08 $Y=0.51 $X2=0 $Y2=0
cc_172 N_A2_M1007_g N_A1_c_239_n 0.0599225f $X=0.905 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A2_M1007_g N_A1_M1000_g 0.00581076f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_174 A2 N_A1_M1000_g 9.45479e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_175 N_A2_c_194_n N_A1_M1000_g 0.0707665f $X=0.905 $Y=1.32 $X2=0 $Y2=0
cc_176 N_A2_M1007_g A1 0.0104022f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_177 A2 A1 0.0132816f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_178 N_A2_c_194_n A1 0.00132825f $X=0.905 $Y=1.32 $X2=0 $Y2=0
cc_179 N_A2_M1007_g X 3.47729e-19 $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A2_M1010_g X 8.92979e-19 $X=1.09 $Y=2.885 $X2=0 $Y2=0
cc_181 A2 X 0.0322201f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_182 N_A2_c_194_n X 0.0022841f $X=0.905 $Y=1.32 $X2=0 $Y2=0
cc_183 N_A2_M1010_g N_VPWR_c_438_n 0.00148932f $X=1.09 $Y=2.885 $X2=0 $Y2=0
cc_184 N_A2_M1010_g N_VPWR_c_439_n 7.58747e-19 $X=1.09 $Y=2.885 $X2=0 $Y2=0
cc_185 N_A2_M1010_g N_VPWR_c_442_n 0.00585385f $X=1.09 $Y=2.885 $X2=0 $Y2=0
cc_186 N_A2_M1010_g N_VPWR_c_437_n 0.0107511f $X=1.09 $Y=2.885 $X2=0 $Y2=0
cc_187 N_A2_M1010_g N_A_233_535#_c_473_n 0.00537389f $X=1.09 $Y=2.885 $X2=0
+ $Y2=0
cc_188 N_A2_M1007_g N_VGND_c_522_n 0.010197f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_189 A2 N_VGND_c_522_n 0.00706417f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_190 N_A2_c_194_n N_VGND_c_522_n 0.00198887f $X=0.905 $Y=1.32 $X2=0 $Y2=0
cc_191 N_A2_M1007_g N_VGND_c_524_n 0.00486043f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A2_M1007_g N_VGND_c_528_n 0.00818711f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_193 A2 N_VGND_c_528_n 9.09151e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_194 N_A1_c_239_n N_B1_M1005_g 0.0107736f $X=1.265 $Y=0.765 $X2=0 $Y2=0
cc_195 A1 N_B1_M1005_g 7.15839e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_196 N_A1_c_242_n N_B1_M1005_g 0.0162059f $X=1.52 $Y=0.93 $X2=0 $Y2=0
cc_197 N_A1_M1000_g N_B1_M1006_g 0.0281989f $X=1.52 $Y=2.885 $X2=0 $Y2=0
cc_198 N_A1_M1000_g N_B1_c_288_n 0.0162059f $X=1.52 $Y=2.885 $X2=0 $Y2=0
cc_199 N_A1_M1000_g N_VPWR_c_439_n 0.0086261f $X=1.52 $Y=2.885 $X2=0 $Y2=0
cc_200 N_A1_M1000_g N_VPWR_c_442_n 0.0035715f $X=1.52 $Y=2.885 $X2=0 $Y2=0
cc_201 N_A1_M1000_g N_VPWR_c_437_n 0.00428043f $X=1.52 $Y=2.885 $X2=0 $Y2=0
cc_202 N_A1_M1000_g N_A_233_535#_c_476_n 2.03427e-19 $X=1.52 $Y=2.885 $X2=0
+ $Y2=0
cc_203 N_A1_M1000_g N_A_233_535#_c_472_n 0.0175512f $X=1.52 $Y=2.885 $X2=0 $Y2=0
cc_204 N_A1_M1000_g N_A_337_397#_c_495_n 0.00912319f $X=1.52 $Y=2.885 $X2=0
+ $Y2=0
cc_205 N_A1_M1000_g N_A_337_397#_c_497_n 0.00322362f $X=1.52 $Y=2.885 $X2=0
+ $Y2=0
cc_206 N_A1_c_239_n N_VGND_c_522_n 0.00232421f $X=1.265 $Y=0.765 $X2=0 $Y2=0
cc_207 A1 N_VGND_c_522_n 8.39633e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_208 N_A1_c_239_n N_VGND_c_524_n 0.00398598f $X=1.265 $Y=0.765 $X2=0 $Y2=0
cc_209 A1 N_VGND_c_524_n 0.00755004f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_210 N_A1_c_242_n N_VGND_c_524_n 0.00335219f $X=1.52 $Y=0.93 $X2=0 $Y2=0
cc_211 N_A1_c_239_n N_VGND_c_528_n 0.00600116f $X=1.265 $Y=0.765 $X2=0 $Y2=0
cc_212 A1 N_VGND_c_528_n 0.0102437f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_213 N_A1_c_242_n N_VGND_c_528_n 0.00415065f $X=1.52 $Y=0.93 $X2=0 $Y2=0
cc_214 A1 A_196_47# 0.00248426f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_215 N_B1_M1005_g N_B2_c_324_n 0.0512219f $X=1.92 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_216 B1 N_B2_c_325_n 7.26181e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_217 N_B1_c_288_n N_B2_c_325_n 8.38584e-19 $X=2.055 $Y=1.32 $X2=0 $Y2=0
cc_218 N_B1_M1006_g N_B2_c_326_n 0.00883253f $X=2.025 $Y=2.195 $X2=0 $Y2=0
cc_219 N_B1_M1006_g N_B2_c_332_n 0.0212173f $X=2.025 $Y=2.195 $X2=0 $Y2=0
cc_220 B1 B2 0.0142588f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_221 N_B1_c_288_n B2 2.30229e-19 $X=2.055 $Y=1.32 $X2=0 $Y2=0
cc_222 B1 N_B2_c_328_n 0.00361248f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_223 N_B1_c_288_n N_B2_c_328_n 0.0211399f $X=2.055 $Y=1.32 $X2=0 $Y2=0
cc_224 N_B1_M1005_g N_B2_c_329_n 0.00705744f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B1_M1006_g N_A_233_535#_c_472_n 0.00802595f $X=2.025 $Y=2.195 $X2=0
+ $Y2=0
cc_226 N_B1_M1006_g N_A_233_535#_c_474_n 0.00225151f $X=2.025 $Y=2.195 $X2=0
+ $Y2=0
cc_227 N_B1_M1006_g N_A_337_397#_c_495_n 0.00101696f $X=2.025 $Y=2.195 $X2=0
+ $Y2=0
cc_228 N_B1_M1006_g N_A_337_397#_c_496_n 0.0133367f $X=2.025 $Y=2.195 $X2=0
+ $Y2=0
cc_229 B1 N_A_337_397#_c_496_n 0.0146523f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_230 N_B1_c_288_n N_A_337_397#_c_496_n 0.00383326f $X=2.055 $Y=1.32 $X2=0
+ $Y2=0
cc_231 N_B1_c_288_n N_A_337_397#_c_497_n 0.00298504f $X=2.055 $Y=1.32 $X2=0
+ $Y2=0
cc_232 N_B1_M1005_g N_VGND_c_523_n 0.00207709f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_233 N_B1_M1005_g N_VGND_c_524_n 0.00429465f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_234 N_B1_M1005_g N_VGND_c_528_n 0.00643997f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_235 N_B2_c_324_n N_C1_c_373_n 0.012457f $X=2.28 $Y=0.765 $X2=-0.19 $Y2=-0.245
cc_236 N_B2_c_326_n N_C1_c_374_n 0.00364831f $X=2.48 $Y=1.695 $X2=0 $Y2=0
cc_237 B2 N_C1_c_374_n 2.47792e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_238 N_B2_c_328_n N_C1_c_374_n 0.0178489f $X=2.595 $Y=1.32 $X2=0 $Y2=0
cc_239 N_B2_c_329_n N_C1_c_374_n 0.00364831f $X=2.595 $Y=1.155 $X2=0 $Y2=0
cc_240 N_B2_c_325_n N_C1_c_375_n 0.010244f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_241 N_B2_M1001_g N_C1_c_378_n 0.0149601f $X=2.455 $Y=2.195 $X2=0 $Y2=0
cc_242 N_B2_c_332_n N_C1_c_378_n 0.00671262f $X=2.48 $Y=1.845 $X2=0 $Y2=0
cc_243 N_B2_M1001_g N_VPWR_c_437_n 0.00393928f $X=2.455 $Y=2.195 $X2=0 $Y2=0
cc_244 N_B2_M1001_g N_A_233_535#_c_472_n 0.00129737f $X=2.455 $Y=2.195 $X2=0
+ $Y2=0
cc_245 N_B2_M1001_g N_A_233_535#_c_474_n 0.00225151f $X=2.455 $Y=2.195 $X2=0
+ $Y2=0
cc_246 N_B2_M1001_g N_A_337_397#_c_496_n 0.00878543f $X=2.455 $Y=2.195 $X2=0
+ $Y2=0
cc_247 N_B2_c_332_n N_A_337_397#_c_496_n 0.00940151f $X=2.48 $Y=1.845 $X2=0
+ $Y2=0
cc_248 B2 N_A_337_397#_c_496_n 0.0145365f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_249 N_B2_c_328_n N_A_337_397#_c_496_n 0.00412243f $X=2.595 $Y=1.32 $X2=0
+ $Y2=0
cc_250 N_B2_M1001_g N_A_337_397#_c_498_n 9.4709e-19 $X=2.455 $Y=2.195 $X2=0
+ $Y2=0
cc_251 N_B2_c_324_n N_VGND_c_523_n 0.00964222f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_252 N_B2_c_325_n N_VGND_c_523_n 0.00121104f $X=2.505 $Y=0.84 $X2=0 $Y2=0
cc_253 N_B2_c_324_n N_VGND_c_524_n 0.0035715f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_254 N_B2_c_324_n N_VGND_c_528_n 0.0040852f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_255 C1 N_VPWR_c_439_n 0.00785184f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_256 C1 N_VPWR_c_443_n 0.0432658f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_257 N_C1_c_380_n N_VPWR_c_443_n 0.00805502f $X=2.885 $Y=2.91 $X2=0 $Y2=0
cc_258 C1 N_VPWR_c_437_n 0.0246955f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_259 N_C1_c_380_n N_VPWR_c_437_n 0.0114868f $X=2.885 $Y=2.91 $X2=0 $Y2=0
cc_260 N_C1_M1009_g N_A_233_535#_c_472_n 0.00399585f $X=2.885 $Y=2.195 $X2=0
+ $Y2=0
cc_261 N_C1_c_378_n N_A_337_397#_c_496_n 0.00164109f $X=3.075 $Y=1.8 $X2=0 $Y2=0
cc_262 N_C1_M1009_g N_A_337_397#_c_498_n 5.6852e-19 $X=2.885 $Y=2.195 $X2=0
+ $Y2=0
cc_263 C1 N_A_337_397#_c_498_n 0.00883186f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_264 N_C1_c_380_n N_A_337_397#_c_498_n 8.73645e-19 $X=2.885 $Y=2.91 $X2=0
+ $Y2=0
cc_265 N_C1_c_373_n N_VGND_c_523_n 0.00779467f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_266 N_C1_c_373_n N_VGND_c_527_n 0.00423721f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_267 N_C1_c_375_n N_VGND_c_527_n 5.35341e-19 $X=3.075 $Y=0.84 $X2=0 $Y2=0
cc_268 N_C1_c_373_n N_VGND_c_528_n 0.00740085f $X=2.865 $Y=0.765 $X2=0 $Y2=0
cc_269 N_X_c_414_n N_VPWR_c_440_n 0.0163326f $X=0.445 $Y=2.82 $X2=0 $Y2=0
cc_270 N_X_M1002_s N_VPWR_c_437_n 0.00344799f $X=0.32 $Y=2.675 $X2=0 $Y2=0
cc_271 N_X_c_414_n N_VPWR_c_437_n 0.0142805f $X=0.445 $Y=2.82 $X2=0 $Y2=0
cc_272 N_X_c_414_n N_A_233_535#_c_476_n 2.66198e-19 $X=0.445 $Y=2.82 $X2=0 $Y2=0
cc_273 N_X_c_414_n N_A_233_535#_c_473_n 3.09595e-19 $X=0.445 $Y=2.82 $X2=0 $Y2=0
cc_274 X N_VGND_c_526_n 0.00831216f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_275 N_X_M1004_s N_VGND_c_528_n 0.0036043f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_276 X N_VGND_c_528_n 0.0069578f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_277 N_VPWR_c_437_n N_A_233_535#_M1010_d 0.00377398f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_278 N_VPWR_c_442_n N_A_233_535#_c_476_n 0.00770662f $X=1.57 $Y=3.33 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_437_n N_A_233_535#_c_476_n 0.00688329f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_439_n N_A_233_535#_c_472_n 0.0218865f $X=1.735 $Y=2.95 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_442_n N_A_233_535#_c_472_n 0.00283061f $X=1.57 $Y=3.33 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_443_n N_A_233_535#_c_472_n 0.00795485f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_437_n N_A_233_535#_c_472_n 0.0186195f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_284 N_A_233_535#_c_472_n N_A_337_397#_c_495_n 0.0142166f $X=2.135 $Y=2.58
+ $X2=0 $Y2=0
cc_285 N_A_233_535#_c_472_n N_A_337_397#_c_496_n 0.0059116f $X=2.135 $Y=2.58
+ $X2=0 $Y2=0
cc_286 N_A_233_535#_c_474_n N_A_337_397#_c_496_n 0.0145058f $X=2.24 $Y=2.26
+ $X2=0 $Y2=0
cc_287 N_VGND_c_528_n A_196_47# 0.00652402f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_288 N_VGND_c_528_n A_399_47# 0.00253354f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
