# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__inv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  5.040000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.170000 1.920000 0.465000 3.245000 ;
        RECT 1.065000 1.920000 1.325000 3.245000 ;
        RECT 1.925000 1.920000 2.185000 3.245000 ;
        RECT 2.785000 1.920000 3.045000 3.245000 ;
        RECT 3.645000 1.920000 3.905000 3.245000 ;
        RECT 4.505000 1.920000 4.765000 3.245000 ;
        RECT 5.365000 1.920000 5.625000 3.245000 ;
        RECT 6.225000 1.920000 6.485000 3.245000 ;
        RECT 7.085000 1.920000 7.380000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.050000 1.550000 6.500000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.704000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.620000 1.920000 6.930000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.085000 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.170000  0.085000 0.465000 1.005000 ;
      RECT 0.635000  0.305000 0.895000 3.050000 ;
      RECT 1.065000  0.085000 1.325000 1.005000 ;
      RECT 1.065000  1.335000 1.325000 1.750000 ;
      RECT 1.495000  0.305000 1.755000 3.050000 ;
      RECT 1.925000  0.085000 2.185000 1.005000 ;
      RECT 1.925000  1.335000 2.185000 1.750000 ;
      RECT 2.355000  0.305000 2.615000 3.050000 ;
      RECT 2.785000  0.085000 3.045000 1.005000 ;
      RECT 2.785000  1.335000 3.045000 1.750000 ;
      RECT 3.215000  0.305000 3.475000 3.050000 ;
      RECT 3.645000  0.085000 3.905000 1.005000 ;
      RECT 3.645000  1.335000 3.905000 1.750000 ;
      RECT 4.075000  0.305000 4.335000 3.050000 ;
      RECT 4.505000  0.085000 4.765000 1.005000 ;
      RECT 4.505000  1.335000 4.765000 1.750000 ;
      RECT 4.935000  0.305000 5.195000 3.050000 ;
      RECT 5.365000  0.085000 5.625000 1.005000 ;
      RECT 5.365000  1.335000 5.625000 1.750000 ;
      RECT 5.795000  0.305000 6.055000 3.050000 ;
      RECT 6.225000  0.085000 6.485000 1.005000 ;
      RECT 6.225000  1.335000 6.485000 1.750000 ;
      RECT 6.655000  0.305000 6.915000 3.050000 ;
      RECT 7.085000  0.085000 7.380000 1.005000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.680000  1.950000 0.850000 2.120000 ;
      RECT 1.110000  1.580000 1.280000 1.750000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.540000  1.950000 1.710000 2.120000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.970000  1.580000 2.140000 1.750000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.400000  1.950000 2.570000 2.120000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.830000  1.580000 3.000000 1.750000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.260000  1.950000 3.430000 2.120000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.690000  1.580000 3.860000 1.750000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 4.120000  1.950000 4.290000 2.120000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.550000  1.580000 4.720000 1.750000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.980000  1.950000 5.150000 2.120000 ;
      RECT 5.410000  1.580000 5.580000 1.750000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.840000  1.950000 6.010000 2.120000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 6.270000  1.580000 6.440000 1.750000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.700000  1.950000 6.870000 2.120000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
  END
END sky130_fd_sc_lp__inv_16
END LIBRARY
