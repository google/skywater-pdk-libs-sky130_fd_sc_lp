* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__clkbuf_16 A VGND VNB VPB VPWR X
X0 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_116_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A a_116_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_116_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND A a_116_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR A a_116_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VPWR A a_116_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_116_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_116_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VPWR a_116_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 X a_116_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 X a_116_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 VGND a_116_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
