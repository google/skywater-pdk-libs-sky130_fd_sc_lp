* File: sky130_fd_sc_lp__dlrbn_lp.pxi.spice
* Created: Wed Sep  2 09:46:22 2020
* 
x_PM_SKY130_FD_SC_LP__DLRBN_LP%D N_D_M1015_g N_D_M1013_g N_D_M1002_g N_D_c_190_n
+ N_D_c_191_n D D N_D_c_192_n N_D_c_193_n PM_SKY130_FD_SC_LP__DLRBN_LP%D
x_PM_SKY130_FD_SC_LP__DLRBN_LP%GATE_N N_GATE_N_M1003_g N_GATE_N_M1018_g
+ N_GATE_N_M1019_g N_GATE_N_c_236_n N_GATE_N_c_237_n GATE_N GATE_N
+ N_GATE_N_c_238_n N_GATE_N_c_239_n PM_SKY130_FD_SC_LP__DLRBN_LP%GATE_N
x_PM_SKY130_FD_SC_LP__DLRBN_LP%A_252_396# N_A_252_396#_M1019_d
+ N_A_252_396#_M1003_d N_A_252_396#_c_301_n N_A_252_396#_c_302_n
+ N_A_252_396#_c_303_n N_A_252_396#_M1017_g N_A_252_396#_M1021_g
+ N_A_252_396#_c_288_n N_A_252_396#_M1007_g N_A_252_396#_M1012_g
+ N_A_252_396#_c_291_n N_A_252_396#_c_305_n N_A_252_396#_M1009_g
+ N_A_252_396#_c_292_n N_A_252_396#_c_293_n N_A_252_396#_c_306_n
+ N_A_252_396#_c_294_n N_A_252_396#_c_308_n N_A_252_396#_c_309_n
+ N_A_252_396#_c_295_n N_A_252_396#_c_296_n N_A_252_396#_c_311_n
+ N_A_252_396#_c_312_n N_A_252_396#_c_297_n N_A_252_396#_c_298_n
+ N_A_252_396#_c_299_n N_A_252_396#_c_300_n
+ PM_SKY130_FD_SC_LP__DLRBN_LP%A_252_396#
x_PM_SKY130_FD_SC_LP__DLRBN_LP%A_27_68# N_A_27_68#_M1015_s N_A_27_68#_M1013_s
+ N_A_27_68#_M1020_g N_A_27_68#_c_439_n N_A_27_68#_c_440_n N_A_27_68#_c_441_n
+ N_A_27_68#_M1011_g N_A_27_68#_c_448_n N_A_27_68#_c_449_n N_A_27_68#_c_461_n
+ N_A_27_68#_c_463_n N_A_27_68#_c_450_n N_A_27_68#_c_451_n N_A_27_68#_c_497_n
+ N_A_27_68#_c_452_n N_A_27_68#_c_453_n N_A_27_68#_c_442_n N_A_27_68#_c_443_n
+ N_A_27_68#_c_444_n N_A_27_68#_c_456_n N_A_27_68#_c_445_n N_A_27_68#_c_458_n
+ N_A_27_68#_c_446_n PM_SKY130_FD_SC_LP__DLRBN_LP%A_27_68#
x_PM_SKY130_FD_SC_LP__DLRBN_LP%A_451_419# N_A_451_419#_M1021_s
+ N_A_451_419#_M1017_s N_A_451_419#_M1000_g N_A_451_419#_M1022_g
+ N_A_451_419#_c_564_n N_A_451_419#_c_577_n N_A_451_419#_c_578_n
+ N_A_451_419#_c_565_n N_A_451_419#_c_566_n N_A_451_419#_c_567_n
+ N_A_451_419#_c_568_n N_A_451_419#_c_569_n N_A_451_419#_c_570_n
+ N_A_451_419#_c_580_n N_A_451_419#_c_571_n N_A_451_419#_c_572_n
+ N_A_451_419#_c_573_n N_A_451_419#_c_574_n
+ PM_SKY130_FD_SC_LP__DLRBN_LP%A_451_419#
x_PM_SKY130_FD_SC_LP__DLRBN_LP%A_952_305# N_A_952_305#_M1024_s
+ N_A_952_305#_M1005_d N_A_952_305#_M1026_g N_A_952_305#_M1029_g
+ N_A_952_305#_c_700_n N_A_952_305#_M1014_g N_A_952_305#_c_701_n
+ N_A_952_305#_M1008_g N_A_952_305#_M1001_g N_A_952_305#_c_703_n
+ N_A_952_305#_M1004_g N_A_952_305#_M1027_g N_A_952_305#_M1006_g
+ N_A_952_305#_c_707_n N_A_952_305#_c_708_n N_A_952_305#_c_720_n
+ N_A_952_305#_c_777_p N_A_952_305#_c_744_p N_A_952_305#_c_709_n
+ N_A_952_305#_c_710_n N_A_952_305#_c_711_n N_A_952_305#_c_712_n
+ N_A_952_305#_c_713_n N_A_952_305#_c_714_n N_A_952_305#_c_715_n
+ N_A_952_305#_c_716_n PM_SKY130_FD_SC_LP__DLRBN_LP%A_952_305#
x_PM_SKY130_FD_SC_LP__DLRBN_LP%A_796_419# N_A_796_419#_M1012_d
+ N_A_796_419#_M1000_d N_A_796_419#_M1005_g N_A_796_419#_c_862_n
+ N_A_796_419#_M1024_g N_A_796_419#_c_876_n N_A_796_419#_c_871_n
+ N_A_796_419#_c_872_n N_A_796_419#_c_863_n N_A_796_419#_c_873_n
+ N_A_796_419#_c_864_n N_A_796_419#_c_865_n N_A_796_419#_c_866_n
+ N_A_796_419#_c_867_n N_A_796_419#_c_868_n N_A_796_419#_c_869_n
+ PM_SKY130_FD_SC_LP__DLRBN_LP%A_796_419#
x_PM_SKY130_FD_SC_LP__DLRBN_LP%RESET_B N_RESET_B_M1028_g N_RESET_B_M1010_g
+ RESET_B RESET_B N_RESET_B_c_973_n N_RESET_B_c_974_n
+ PM_SKY130_FD_SC_LP__DLRBN_LP%RESET_B
x_PM_SKY130_FD_SC_LP__DLRBN_LP%A_1617_76# N_A_1617_76#_M1004_s
+ N_A_1617_76#_M1027_s N_A_1617_76#_M1023_g N_A_1617_76#_M1016_g
+ N_A_1617_76#_M1025_g N_A_1617_76#_c_1015_n N_A_1617_76#_c_1016_n
+ N_A_1617_76#_c_1017_n N_A_1617_76#_c_1018_n N_A_1617_76#_c_1019_n
+ N_A_1617_76#_c_1020_n N_A_1617_76#_c_1021_n N_A_1617_76#_c_1022_n
+ N_A_1617_76#_c_1023_n PM_SKY130_FD_SC_LP__DLRBN_LP%A_1617_76#
x_PM_SKY130_FD_SC_LP__DLRBN_LP%VPWR N_VPWR_M1013_d N_VPWR_M1017_d N_VPWR_M1026_d
+ N_VPWR_M1028_d N_VPWR_M1027_d N_VPWR_c_1080_n N_VPWR_c_1081_n N_VPWR_c_1082_n
+ N_VPWR_c_1083_n N_VPWR_c_1084_n VPWR N_VPWR_c_1085_n N_VPWR_c_1086_n
+ N_VPWR_c_1087_n N_VPWR_c_1088_n N_VPWR_c_1089_n N_VPWR_c_1079_n
+ N_VPWR_c_1091_n N_VPWR_c_1092_n N_VPWR_c_1093_n N_VPWR_c_1094_n
+ N_VPWR_c_1095_n PM_SKY130_FD_SC_LP__DLRBN_LP%VPWR
x_PM_SKY130_FD_SC_LP__DLRBN_LP%Q N_Q_M1008_d N_Q_M1001_d N_Q_c_1181_n
+ N_Q_c_1182_n Q Q Q Q Q PM_SKY130_FD_SC_LP__DLRBN_LP%Q
x_PM_SKY130_FD_SC_LP__DLRBN_LP%Q_N N_Q_N_M1025_d N_Q_N_M1016_d N_Q_N_c_1209_n
+ Q_N Q_N Q_N N_Q_N_c_1212_n N_Q_N_c_1210_n PM_SKY130_FD_SC_LP__DLRBN_LP%Q_N
x_PM_SKY130_FD_SC_LP__DLRBN_LP%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_M1029_d
+ N_VGND_M1010_d N_VGND_M1006_d N_VGND_c_1232_n N_VGND_c_1233_n N_VGND_c_1234_n
+ N_VGND_c_1235_n N_VGND_c_1236_n N_VGND_c_1237_n VGND N_VGND_c_1238_n
+ N_VGND_c_1239_n N_VGND_c_1240_n N_VGND_c_1241_n N_VGND_c_1242_n
+ N_VGND_c_1243_n N_VGND_c_1244_n N_VGND_c_1245_n N_VGND_c_1246_n
+ N_VGND_c_1247_n N_VGND_c_1248_n PM_SKY130_FD_SC_LP__DLRBN_LP%VGND
cc_1 VNB N_D_M1015_g 0.0327748f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.55
cc_2 VNB N_D_M1002_g 0.0263836f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.55
cc_3 VNB N_D_c_190_n 0.0225774f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.24
cc_4 VNB N_D_c_191_n 0.00510434f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.76
cc_5 VNB N_D_c_192_n 0.0264349f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.255
cc_6 VNB N_D_c_193_n 0.00424976f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.255
cc_7 VNB N_GATE_N_M1003_g 0.00174718f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.55
cc_8 VNB N_GATE_N_M1018_g 0.0201686f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.48
cc_9 VNB N_GATE_N_M1019_g 0.0242712f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.55
cc_10 VNB N_GATE_N_c_236_n 0.0264059f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.24
cc_11 VNB N_GATE_N_c_237_n 0.0275909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_GATE_N_c_238_n 0.0276074f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.295
cc_13 VNB N_GATE_N_c_239_n 0.00685502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_252_396#_M1021_g 0.0236418f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.09
cc_15 VNB N_A_252_396#_c_288_n 0.00629424f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.76
cc_16 VNB N_A_252_396#_M1007_g 0.0213175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_252_396#_M1012_g 0.0226041f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.255
cc_18 VNB N_A_252_396#_c_291_n 0.0216673f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.295
cc_19 VNB N_A_252_396#_c_292_n 0.0292109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_252_396#_c_293_n 0.019506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_252_396#_c_294_n 0.0111577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_252_396#_c_295_n 0.0173039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_252_396#_c_296_n 0.0185803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_252_396#_c_297_n 0.0015711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_252_396#_c_298_n 0.0307941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_252_396#_c_299_n 0.00495302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_252_396#_c_300_n 0.0378262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_68#_c_439_n 0.022027f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.24
cc_29 VNB N_A_27_68#_c_440_n 0.00963373f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.09
cc_30 VNB N_A_27_68#_c_441_n 0.0162651f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.24
cc_31 VNB N_A_27_68#_c_442_n 0.00108032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_68#_c_443_n 0.00852979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_68#_c_444_n 0.0270872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_68#_c_445_n 0.0415592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_68#_c_446_n 0.0466695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_451_419#_M1022_g 0.0286554f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.24
cc_37 VNB N_A_451_419#_c_564_n 0.0212764f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.585
cc_38 VNB N_A_451_419#_c_565_n 0.00453274f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.255
cc_39 VNB N_A_451_419#_c_566_n 0.0144723f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.255
cc_40 VNB N_A_451_419#_c_567_n 0.00329503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_451_419#_c_568_n 0.014608f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.295
cc_42 VNB N_A_451_419#_c_569_n 0.00255857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_451_419#_c_570_n 0.0122615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_451_419#_c_571_n 0.00873275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_451_419#_c_572_n 0.0217466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_451_419#_c_573_n 0.00344066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_451_419#_c_574_n 0.0342421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_952_305#_M1029_g 0.0614304f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.24
cc_49 VNB N_A_952_305#_c_700_n 0.0156466f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.24
cc_50 VNB N_A_952_305#_c_701_n 0.0186123f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_51 VNB N_A_952_305#_M1001_g 0.00245261f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.255
cc_52 VNB N_A_952_305#_c_703_n 0.0430236f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.255
cc_53 VNB N_A_952_305#_M1004_g 0.0412967f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.665
cc_54 VNB N_A_952_305#_M1027_g 0.0155544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_952_305#_M1006_g 0.0321101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_952_305#_c_707_n 0.0168085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_952_305#_c_708_n 0.00181198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_952_305#_c_709_n 9.97909e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_952_305#_c_710_n 0.00593009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_952_305#_c_711_n 0.00728432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_952_305#_c_712_n 0.0256529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_952_305#_c_713_n 0.0140978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_952_305#_c_714_n 0.0103112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_952_305#_c_715_n 0.0228474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_952_305#_c_716_n 0.0603297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_796_419#_c_862_n 0.0136353f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.24
cc_67 VNB N_A_796_419#_c_863_n 0.0134543f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.255
cc_68 VNB N_A_796_419#_c_864_n 0.00918331f $X=-0.19 $Y=-0.245 $X2=0.637
+ $Y2=1.295
cc_69 VNB N_A_796_419#_c_865_n 0.00355608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_796_419#_c_866_n 0.0109602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_796_419#_c_867_n 0.00435324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_796_419#_c_868_n 0.0611428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_796_419#_c_869_n 0.0541145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_RESET_B_M1010_g 0.0343342f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.48
cc_75 VNB N_RESET_B_c_973_n 0.00233667f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.76
cc_76 VNB N_RESET_B_c_974_n 0.0167278f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_77 VNB N_A_1617_76#_M1023_g 0.0193316f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.09
cc_78 VNB N_A_1617_76#_M1025_g 0.0253324f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.76
cc_79 VNB N_A_1617_76#_c_1015_n 0.021457f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.255
cc_80 VNB N_A_1617_76#_c_1016_n 0.0121906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1617_76#_c_1017_n 0.00220477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1617_76#_c_1018_n 0.00390811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1617_76#_c_1019_n 0.0172769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1617_76#_c_1020_n 0.0181067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1617_76#_c_1021_n 0.00728657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1617_76#_c_1022_n 0.00144692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1617_76#_c_1023_n 0.0286062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VPWR_c_1079_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_Q_c_1181_n 0.00990997f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.09
cc_90 VNB N_Q_c_1182_n 0.0117837f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.24
cc_91 VNB Q 0.00316993f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.09
cc_92 VNB N_Q_N_c_1209_n 0.0255865f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.55
cc_93 VNB N_Q_N_c_1210_n 0.0402092f $X=-0.19 $Y=-0.245 $X2=0.637 $Y2=1.665
cc_94 VNB N_VGND_c_1232_n 0.00874652f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_95 VNB N_VGND_c_1233_n 0.0498566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1234_n 0.00584537f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.255
cc_97 VNB N_VGND_c_1235_n 0.00931215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1236_n 0.0294546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1237_n 0.00714724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1238_n 0.0276622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1239_n 0.0558072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1240_n 0.0296297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1241_n 0.0531988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1242_n 0.0281784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1243_n 0.574183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1244_n 0.00567616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1245_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1246_n 0.00631189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1247_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1248_n 0.00616439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VPB N_D_M1013_g 0.035779f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.48
cc_112 VPB N_D_c_191_n 0.0104703f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.76
cc_113 VPB N_D_c_193_n 0.00314739f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.255
cc_114 VPB N_GATE_N_M1003_g 0.0411957f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.55
cc_115 VPB N_GATE_N_c_239_n 0.00351153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_252_396#_c_301_n 0.0339811f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.48
cc_117 VPB N_A_252_396#_c_302_n 0.0192157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_252_396#_c_303_n 0.0242663f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.09
cc_119 VPB N_A_252_396#_c_288_n 0.0105671f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.76
cc_120 VPB N_A_252_396#_c_305_n 0.0294557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_252_396#_c_306_n 0.00918958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_252_396#_c_294_n 0.00361674f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_252_396#_c_308_n 0.0116164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_252_396#_c_309_n 0.0142262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_252_396#_c_295_n 0.00537892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_252_396#_c_311_n 0.00700891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_252_396#_c_312_n 0.0570783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_27_68#_M1020_g 0.025561f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.09
cc_129 VPB N_A_27_68#_c_448_n 0.00932077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_27_68#_c_449_n 0.0218177f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.255
cc_131 VPB N_A_27_68#_c_450_n 0.0240189f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_27_68#_c_451_n 9.26011e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_27_68#_c_452_n 0.00488334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_27_68#_c_453_n 4.309e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_27_68#_c_442_n 0.001519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_27_68#_c_443_n 0.0229362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_27_68#_c_456_n 0.015815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_27_68#_c_445_n 0.0147035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_27_68#_c_458_n 0.00758388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_451_419#_M1000_g 0.0371888f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.09
cc_141 VPB N_A_451_419#_c_564_n 0.00111416f $X=-0.19 $Y=1.655 $X2=0.595
+ $Y2=1.585
cc_142 VPB N_A_451_419#_c_577_n 0.010451f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_143 VPB N_A_451_419#_c_578_n 0.00776781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_451_419#_c_565_n 8.14307e-19 $X=-0.19 $Y=1.655 $X2=0.605
+ $Y2=1.255
cc_145 VPB N_A_451_419#_c_580_n 0.00689333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_451_419#_c_571_n 0.00433789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_451_419#_c_572_n 0.00825912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_952_305#_M1026_g 0.0328108f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.09
cc_149 VPB N_A_952_305#_M1001_g 0.0570086f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.255
cc_150 VPB N_A_952_305#_M1027_g 0.031868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_952_305#_c_720_n 0.00901773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_952_305#_c_709_n 0.0100814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_952_305#_c_710_n 0.00270582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_952_305#_c_715_n 0.0277804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_796_419#_M1005_g 0.0300962f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.09
cc_156 VPB N_A_796_419#_c_871_n 0.0109933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_796_419#_c_872_n 0.0036128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_796_419#_c_873_n 0.00196714f $X=-0.19 $Y=1.655 $X2=0.637
+ $Y2=1.255
cc_159 VPB N_A_796_419#_c_865_n 0.00414265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_796_419#_c_866_n 0.0165024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_M1028_g 0.0298341f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.55
cc_162 VPB N_RESET_B_c_973_n 0.00151586f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.76
cc_163 VPB N_RESET_B_c_974_n 0.0429796f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_164 VPB N_A_1617_76#_M1016_g 0.033609f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.24
cc_165 VPB N_A_1617_76#_c_1016_n 0.00347372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_1617_76#_c_1018_n 0.0186203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_1617_76#_c_1022_n 7.54819e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1080_n 0.00344978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1081_n 0.00240024f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.255
cc_170 VPB N_VPWR_c_1082_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1083_n 0.00696923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1084_n 0.0226092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1085_n 0.0477173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1086_n 0.0495506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1087_n 0.0513003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1088_n 0.0351395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1089_n 0.0269338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1079_n 0.081426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1091_n 0.0267049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1092_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1093_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1094_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1095_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB Q 0.0163455f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.09
cc_185 VPB Q_N 0.043146f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.09
cc_186 VPB N_Q_N_c_1212_n 0.0241524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_Q_N_c_1210_n 0.0098162f $X=-0.19 $Y=1.655 $X2=0.637 $Y2=1.665
cc_188 N_D_M1013_g N_GATE_N_M1003_g 0.0481777f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_189 N_D_c_191_n N_GATE_N_M1003_g 0.00740834f $X=0.595 $Y=1.76 $X2=0 $Y2=0
cc_190 N_D_M1002_g N_GATE_N_M1018_g 0.0172222f $X=0.855 $Y=0.55 $X2=0 $Y2=0
cc_191 N_D_c_192_n N_GATE_N_c_236_n 0.00740834f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_192 N_D_c_193_n N_GATE_N_c_236_n 0.00218125f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_193 N_D_M1002_g N_GATE_N_c_237_n 0.00728901f $X=0.855 $Y=0.55 $X2=0 $Y2=0
cc_194 N_D_c_190_n N_GATE_N_c_238_n 0.00728901f $X=0.675 $Y=1.24 $X2=0 $Y2=0
cc_195 N_D_c_192_n N_GATE_N_c_238_n 0.00666611f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_196 N_D_c_193_n N_GATE_N_c_238_n 8.42766e-19 $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_197 N_D_M1002_g N_GATE_N_c_239_n 0.00438409f $X=0.855 $Y=0.55 $X2=0 $Y2=0
cc_198 N_D_c_192_n N_GATE_N_c_239_n 0.00117005f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_199 N_D_c_193_n N_GATE_N_c_239_n 0.043276f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_200 N_D_M1013_g N_A_252_396#_c_309_n 0.0010579f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_201 N_D_M1013_g N_A_27_68#_c_448_n 0.00458765f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_202 N_D_M1013_g N_A_27_68#_c_449_n 0.00874038f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_203 N_D_M1013_g N_A_27_68#_c_461_n 0.0163275f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_204 N_D_c_193_n N_A_27_68#_c_461_n 0.00857499f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_205 N_D_M1013_g N_A_27_68#_c_463_n 5.84508e-19 $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_206 N_D_M1015_g N_A_27_68#_c_444_n 0.0101793f $X=0.495 $Y=0.55 $X2=0 $Y2=0
cc_207 N_D_M1002_g N_A_27_68#_c_444_n 0.00125133f $X=0.855 $Y=0.55 $X2=0 $Y2=0
cc_208 N_D_M1013_g N_A_27_68#_c_456_n 0.00506206f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_209 N_D_c_191_n N_A_27_68#_c_456_n 0.00127074f $X=0.595 $Y=1.76 $X2=0 $Y2=0
cc_210 N_D_c_193_n N_A_27_68#_c_456_n 0.005453f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_211 N_D_M1015_g N_A_27_68#_c_445_n 0.0246835f $X=0.495 $Y=0.55 $X2=0 $Y2=0
cc_212 N_D_M1013_g N_A_27_68#_c_445_n 0.00459653f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_213 N_D_c_193_n N_A_27_68#_c_445_n 0.0503719f $X=0.605 $Y=1.255 $X2=0 $Y2=0
cc_214 N_D_M1013_g N_A_27_68#_c_458_n 3.84191e-19 $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_215 N_D_M1013_g N_VPWR_c_1080_n 0.0112691f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_216 N_D_M1013_g N_VPWR_c_1079_n 0.00688048f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_217 N_D_M1013_g N_VPWR_c_1091_n 0.00687065f $X=0.605 $Y=2.48 $X2=0 $Y2=0
cc_218 N_D_M1015_g N_VGND_c_1232_n 0.00192363f $X=0.495 $Y=0.55 $X2=0 $Y2=0
cc_219 N_D_M1002_g N_VGND_c_1232_n 0.0131321f $X=0.855 $Y=0.55 $X2=0 $Y2=0
cc_220 N_D_M1015_g N_VGND_c_1238_n 0.00457319f $X=0.495 $Y=0.55 $X2=0 $Y2=0
cc_221 N_D_M1002_g N_VGND_c_1238_n 0.0040395f $X=0.855 $Y=0.55 $X2=0 $Y2=0
cc_222 N_D_M1015_g N_VGND_c_1243_n 0.00895391f $X=0.495 $Y=0.55 $X2=0 $Y2=0
cc_223 N_D_M1002_g N_VGND_c_1243_n 0.00772493f $X=0.855 $Y=0.55 $X2=0 $Y2=0
cc_224 N_GATE_N_M1003_g N_A_252_396#_c_302_n 0.014168f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_225 N_GATE_N_M1019_g N_A_252_396#_c_292_n 0.00121063f $X=1.645 $Y=0.55 $X2=0
+ $Y2=0
cc_226 N_GATE_N_M1003_g N_A_252_396#_c_309_n 0.00643729f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_227 N_GATE_N_c_236_n N_A_252_396#_c_309_n 0.00118564f $X=1.255 $Y=1.63 $X2=0
+ $Y2=0
cc_228 N_GATE_N_c_239_n N_A_252_396#_c_309_n 0.0217744f $X=1.335 $Y=1.125 $X2=0
+ $Y2=0
cc_229 N_GATE_N_M1003_g N_A_252_396#_c_295_n 0.00485081f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_230 N_GATE_N_M1018_g N_A_252_396#_c_295_n 0.00215465f $X=1.285 $Y=0.55 $X2=0
+ $Y2=0
cc_231 N_GATE_N_M1019_g N_A_252_396#_c_295_n 0.0150526f $X=1.645 $Y=0.55 $X2=0
+ $Y2=0
cc_232 N_GATE_N_c_237_n N_A_252_396#_c_295_n 0.00560285f $X=1.645 $Y=1.035 $X2=0
+ $Y2=0
cc_233 N_GATE_N_c_238_n N_A_252_396#_c_295_n 0.0118479f $X=1.335 $Y=1.125 $X2=0
+ $Y2=0
cc_234 N_GATE_N_c_239_n N_A_252_396#_c_295_n 0.0585837f $X=1.335 $Y=1.125 $X2=0
+ $Y2=0
cc_235 N_GATE_N_M1003_g N_A_252_396#_c_311_n 0.00362226f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_236 N_GATE_N_c_237_n N_A_252_396#_c_298_n 0.00121063f $X=1.645 $Y=1.035 $X2=0
+ $Y2=0
cc_237 N_GATE_N_M1003_g N_A_27_68#_c_449_n 6.28179e-19 $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_238 N_GATE_N_M1003_g N_A_27_68#_c_461_n 0.0196757f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_239 N_GATE_N_c_239_n N_A_27_68#_c_461_n 0.00397107f $X=1.335 $Y=1.125 $X2=0
+ $Y2=0
cc_240 N_GATE_N_M1003_g N_A_27_68#_c_463_n 0.0114944f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_241 N_GATE_N_M1003_g N_A_27_68#_c_451_n 0.00755618f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_242 N_GATE_N_M1003_g N_A_27_68#_c_456_n 0.00183997f $X=1.135 $Y=2.48 $X2=0
+ $Y2=0
cc_243 N_GATE_N_M1019_g N_A_451_419#_c_564_n 0.00115627f $X=1.645 $Y=0.55 $X2=0
+ $Y2=0
cc_244 N_GATE_N_M1019_g N_A_451_419#_c_570_n 0.0023132f $X=1.645 $Y=0.55 $X2=0
+ $Y2=0
cc_245 N_GATE_N_M1003_g N_VPWR_c_1080_n 0.00923464f $X=1.135 $Y=2.48 $X2=0 $Y2=0
cc_246 N_GATE_N_M1003_g N_VPWR_c_1085_n 0.00659216f $X=1.135 $Y=2.48 $X2=0 $Y2=0
cc_247 N_GATE_N_M1003_g N_VPWR_c_1079_n 0.0068215f $X=1.135 $Y=2.48 $X2=0 $Y2=0
cc_248 N_GATE_N_M1018_g N_VGND_c_1232_n 0.0123258f $X=1.285 $Y=0.55 $X2=0 $Y2=0
cc_249 N_GATE_N_M1019_g N_VGND_c_1232_n 0.00192363f $X=1.645 $Y=0.55 $X2=0 $Y2=0
cc_250 N_GATE_N_c_236_n N_VGND_c_1232_n 0.00237457f $X=1.255 $Y=1.63 $X2=0 $Y2=0
cc_251 N_GATE_N_c_237_n N_VGND_c_1232_n 3.10581e-19 $X=1.645 $Y=1.035 $X2=0
+ $Y2=0
cc_252 N_GATE_N_c_239_n N_VGND_c_1232_n 0.0129101f $X=1.335 $Y=1.125 $X2=0 $Y2=0
cc_253 N_GATE_N_M1018_g N_VGND_c_1233_n 0.0040395f $X=1.285 $Y=0.55 $X2=0 $Y2=0
cc_254 N_GATE_N_M1019_g N_VGND_c_1233_n 0.00457319f $X=1.645 $Y=0.55 $X2=0 $Y2=0
cc_255 N_GATE_N_M1018_g N_VGND_c_1243_n 0.00772493f $X=1.285 $Y=0.55 $X2=0 $Y2=0
cc_256 N_GATE_N_M1019_g N_VGND_c_1243_n 0.00904779f $X=1.645 $Y=0.55 $X2=0 $Y2=0
cc_257 N_A_252_396#_c_306_n N_A_27_68#_M1020_g 0.0219891f $X=2.665 $Y=1.945
+ $X2=0 $Y2=0
cc_258 N_A_252_396#_c_296_n N_A_27_68#_c_439_n 0.0135657f $X=4.03 $Y=0.94 $X2=0
+ $Y2=0
cc_259 N_A_252_396#_c_300_n N_A_27_68#_c_439_n 0.0217199f $X=4.195 $Y=1.02 $X2=0
+ $Y2=0
cc_260 N_A_252_396#_M1007_g N_A_27_68#_c_440_n 0.00810819f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_261 N_A_252_396#_c_296_n N_A_27_68#_c_440_n 0.00294904f $X=4.03 $Y=0.94 $X2=0
+ $Y2=0
cc_262 N_A_252_396#_M1007_g N_A_27_68#_c_441_n 0.00702535f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_263 N_A_252_396#_M1012_g N_A_27_68#_c_441_n 0.0217199f $X=4.105 $Y=0.445
+ $X2=0 $Y2=0
cc_264 N_A_252_396#_M1003_d N_A_27_68#_c_461_n 0.00278736f $X=1.26 $Y=1.98 $X2=0
+ $Y2=0
cc_265 N_A_252_396#_c_309_n N_A_27_68#_c_461_n 0.00727153f $X=1.695 $Y=2.085
+ $X2=0 $Y2=0
cc_266 N_A_252_396#_c_311_n N_A_27_68#_c_461_n 0.00943257f $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_267 N_A_252_396#_c_312_n N_A_27_68#_c_461_n 8.26094e-19 $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_268 N_A_252_396#_M1003_d N_A_27_68#_c_463_n 0.0108565f $X=1.26 $Y=1.98 $X2=0
+ $Y2=0
cc_269 N_A_252_396#_c_311_n N_A_27_68#_c_463_n 0.00347514f $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_270 N_A_252_396#_c_312_n N_A_27_68#_c_463_n 2.58224e-19 $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_271 N_A_252_396#_M1003_d N_A_27_68#_c_450_n 0.0063409f $X=1.26 $Y=1.98 $X2=0
+ $Y2=0
cc_272 N_A_252_396#_c_303_n N_A_27_68#_c_450_n 0.0171246f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_273 N_A_252_396#_c_311_n N_A_27_68#_c_450_n 0.0137582f $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_274 N_A_252_396#_c_312_n N_A_27_68#_c_450_n 0.00415059f $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_275 N_A_252_396#_c_303_n N_A_27_68#_c_497_n 0.0239661f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_276 N_A_252_396#_c_303_n N_A_27_68#_c_453_n 0.00813192f $X=2.665 $Y=2.02
+ $X2=0 $Y2=0
cc_277 N_A_252_396#_c_306_n N_A_27_68#_c_442_n 0.00261321f $X=2.665 $Y=1.945
+ $X2=0 $Y2=0
cc_278 N_A_252_396#_c_288_n N_A_27_68#_c_443_n 0.00955809f $X=2.715 $Y=1.87
+ $X2=0 $Y2=0
cc_279 N_A_252_396#_c_292_n N_A_27_68#_c_446_n 0.00810819f $X=2.995 $Y=0.93
+ $X2=0 $Y2=0
cc_280 N_A_252_396#_c_296_n N_A_27_68#_c_446_n 0.00872696f $X=4.03 $Y=0.94 $X2=0
+ $Y2=0
cc_281 N_A_252_396#_c_297_n N_A_27_68#_c_446_n 0.00117811f $X=2.595 $Y=1.02
+ $X2=0 $Y2=0
cc_282 N_A_252_396#_c_298_n N_A_27_68#_c_446_n 0.0119789f $X=2.595 $Y=1.02 $X2=0
+ $Y2=0
cc_283 N_A_252_396#_c_299_n N_A_27_68#_c_446_n 9.0165e-19 $X=4.195 $Y=0.94 $X2=0
+ $Y2=0
cc_284 N_A_252_396#_c_300_n N_A_27_68#_c_446_n 0.00589881f $X=4.195 $Y=1.02
+ $X2=0 $Y2=0
cc_285 N_A_252_396#_c_305_n N_A_451_419#_M1000_g 0.0286238f $X=4.395 $Y=2.01
+ $X2=0 $Y2=0
cc_286 N_A_252_396#_c_308_n N_A_451_419#_M1000_g 0.0050503f $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_287 N_A_252_396#_M1012_g N_A_451_419#_M1022_g 0.0146609f $X=4.105 $Y=0.445
+ $X2=0 $Y2=0
cc_288 N_A_252_396#_c_299_n N_A_451_419#_M1022_g 0.0014395f $X=4.195 $Y=0.94
+ $X2=0 $Y2=0
cc_289 N_A_252_396#_c_300_n N_A_451_419#_M1022_g 0.0097061f $X=4.195 $Y=1.02
+ $X2=0 $Y2=0
cc_290 N_A_252_396#_M1021_g N_A_451_419#_c_564_n 0.00567024f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_291 N_A_252_396#_c_288_n N_A_451_419#_c_564_n 0.00170613f $X=2.715 $Y=1.87
+ $X2=0 $Y2=0
cc_292 N_A_252_396#_c_292_n N_A_451_419#_c_564_n 0.0134812f $X=2.995 $Y=0.93
+ $X2=0 $Y2=0
cc_293 N_A_252_396#_c_295_n N_A_451_419#_c_564_n 0.0770425f $X=1.86 $Y=0.55
+ $X2=0 $Y2=0
cc_294 N_A_252_396#_c_297_n N_A_451_419#_c_564_n 0.0475656f $X=2.595 $Y=1.02
+ $X2=0 $Y2=0
cc_295 N_A_252_396#_c_301_n N_A_451_419#_c_577_n 0.0188424f $X=2.54 $Y=1.945
+ $X2=0 $Y2=0
cc_296 N_A_252_396#_c_303_n N_A_451_419#_c_577_n 0.00448325f $X=2.665 $Y=2.02
+ $X2=0 $Y2=0
cc_297 N_A_252_396#_c_295_n N_A_451_419#_c_577_n 0.00594398f $X=1.86 $Y=0.55
+ $X2=0 $Y2=0
cc_298 N_A_252_396#_c_311_n N_A_451_419#_c_577_n 0.051268f $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_299 N_A_252_396#_c_312_n N_A_451_419#_c_577_n 0.00636351f $X=1.865 $Y=2.125
+ $X2=0 $Y2=0
cc_300 N_A_252_396#_c_301_n N_A_451_419#_c_578_n 0.00283071f $X=2.54 $Y=1.945
+ $X2=0 $Y2=0
cc_301 N_A_252_396#_c_288_n N_A_451_419#_c_578_n 0.0108564f $X=2.715 $Y=1.87
+ $X2=0 $Y2=0
cc_302 N_A_252_396#_c_293_n N_A_451_419#_c_578_n 7.14025e-19 $X=2.61 $Y=1.525
+ $X2=0 $Y2=0
cc_303 N_A_252_396#_c_306_n N_A_451_419#_c_578_n 0.0082979f $X=2.665 $Y=1.945
+ $X2=0 $Y2=0
cc_304 N_A_252_396#_c_297_n N_A_451_419#_c_578_n 0.0149283f $X=2.595 $Y=1.02
+ $X2=0 $Y2=0
cc_305 N_A_252_396#_c_293_n N_A_451_419#_c_565_n 0.00366786f $X=2.61 $Y=1.525
+ $X2=0 $Y2=0
cc_306 N_A_252_396#_c_297_n N_A_451_419#_c_565_n 0.00689674f $X=2.595 $Y=1.02
+ $X2=0 $Y2=0
cc_307 N_A_252_396#_c_296_n N_A_451_419#_c_566_n 0.037492f $X=4.03 $Y=0.94 $X2=0
+ $Y2=0
cc_308 N_A_252_396#_c_292_n N_A_451_419#_c_567_n 0.00120761f $X=2.995 $Y=0.93
+ $X2=0 $Y2=0
cc_309 N_A_252_396#_c_296_n N_A_451_419#_c_567_n 0.0115201f $X=4.03 $Y=0.94
+ $X2=0 $Y2=0
cc_310 N_A_252_396#_c_297_n N_A_451_419#_c_567_n 0.0132448f $X=2.595 $Y=1.02
+ $X2=0 $Y2=0
cc_311 N_A_252_396#_c_298_n N_A_451_419#_c_567_n 0.00202826f $X=2.595 $Y=1.02
+ $X2=0 $Y2=0
cc_312 N_A_252_396#_c_291_n N_A_451_419#_c_568_n 0.00752306f $X=4.315 $Y=1.525
+ $X2=0 $Y2=0
cc_313 N_A_252_396#_c_305_n N_A_451_419#_c_568_n 3.86518e-19 $X=4.395 $Y=2.01
+ $X2=0 $Y2=0
cc_314 N_A_252_396#_c_294_n N_A_451_419#_c_568_n 0.0103644f $X=4.445 $Y=1.6
+ $X2=0 $Y2=0
cc_315 N_A_252_396#_c_299_n N_A_451_419#_c_568_n 0.0186556f $X=4.195 $Y=0.94
+ $X2=0 $Y2=0
cc_316 N_A_252_396#_c_300_n N_A_451_419#_c_568_n 0.00135872f $X=4.195 $Y=1.02
+ $X2=0 $Y2=0
cc_317 N_A_252_396#_c_291_n N_A_451_419#_c_569_n 0.00455784f $X=4.315 $Y=1.525
+ $X2=0 $Y2=0
cc_318 N_A_252_396#_M1021_g N_A_451_419#_c_570_n 0.00769509f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_319 N_A_252_396#_M1007_g N_A_451_419#_c_570_n 0.00110975f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_320 N_A_252_396#_c_292_n N_A_451_419#_c_570_n 0.00337384f $X=2.995 $Y=0.93
+ $X2=0 $Y2=0
cc_321 N_A_252_396#_c_295_n N_A_451_419#_c_570_n 0.028143f $X=1.86 $Y=0.55 $X2=0
+ $Y2=0
cc_322 N_A_252_396#_c_297_n N_A_451_419#_c_570_n 0.0070399f $X=2.595 $Y=1.02
+ $X2=0 $Y2=0
cc_323 N_A_252_396#_c_301_n N_A_451_419#_c_580_n 0.0068694f $X=2.54 $Y=1.945
+ $X2=0 $Y2=0
cc_324 N_A_252_396#_c_293_n N_A_451_419#_c_580_n 0.00162168f $X=2.61 $Y=1.525
+ $X2=0 $Y2=0
cc_325 N_A_252_396#_c_295_n N_A_451_419#_c_580_n 0.0141938f $X=1.86 $Y=0.55
+ $X2=0 $Y2=0
cc_326 N_A_252_396#_c_291_n N_A_451_419#_c_571_n 0.00553492f $X=4.315 $Y=1.525
+ $X2=0 $Y2=0
cc_327 N_A_252_396#_c_294_n N_A_451_419#_c_571_n 5.63343e-19 $X=4.445 $Y=1.6
+ $X2=0 $Y2=0
cc_328 N_A_252_396#_c_308_n N_A_451_419#_c_571_n 4.77012e-19 $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_329 N_A_252_396#_c_296_n N_A_451_419#_c_571_n 0.0184764f $X=4.03 $Y=0.94
+ $X2=0 $Y2=0
cc_330 N_A_252_396#_c_291_n N_A_451_419#_c_572_n 0.0159456f $X=4.315 $Y=1.525
+ $X2=0 $Y2=0
cc_331 N_A_252_396#_c_308_n N_A_451_419#_c_572_n 0.00259054f $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_332 N_A_252_396#_c_296_n N_A_451_419#_c_572_n 0.00155643f $X=4.03 $Y=0.94
+ $X2=0 $Y2=0
cc_333 N_A_252_396#_c_299_n N_A_451_419#_c_573_n 0.0131032f $X=4.195 $Y=0.94
+ $X2=0 $Y2=0
cc_334 N_A_252_396#_c_300_n N_A_451_419#_c_573_n 0.00150212f $X=4.195 $Y=1.02
+ $X2=0 $Y2=0
cc_335 N_A_252_396#_c_300_n N_A_451_419#_c_574_n 0.0156433f $X=4.195 $Y=1.02
+ $X2=0 $Y2=0
cc_336 N_A_252_396#_c_308_n N_A_952_305#_M1026_g 0.0488001f $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_337 N_A_252_396#_c_294_n N_A_952_305#_c_710_n 0.0011747f $X=4.445 $Y=1.6
+ $X2=0 $Y2=0
cc_338 N_A_252_396#_c_294_n N_A_952_305#_c_715_n 0.0488001f $X=4.445 $Y=1.6
+ $X2=0 $Y2=0
cc_339 N_A_252_396#_c_305_n N_A_796_419#_c_876_n 0.0203859f $X=4.395 $Y=2.01
+ $X2=0 $Y2=0
cc_340 N_A_252_396#_c_305_n N_A_796_419#_c_871_n 0.0196763f $X=4.395 $Y=2.01
+ $X2=0 $Y2=0
cc_341 N_A_252_396#_c_294_n N_A_796_419#_c_871_n 2.48776e-19 $X=4.445 $Y=1.6
+ $X2=0 $Y2=0
cc_342 N_A_252_396#_c_305_n N_A_796_419#_c_872_n 0.00145441f $X=4.395 $Y=2.01
+ $X2=0 $Y2=0
cc_343 N_A_252_396#_c_294_n N_A_796_419#_c_872_n 8.26447e-19 $X=4.445 $Y=1.6
+ $X2=0 $Y2=0
cc_344 N_A_252_396#_M1012_g N_A_796_419#_c_864_n 0.0139825f $X=4.105 $Y=0.445
+ $X2=0 $Y2=0
cc_345 N_A_252_396#_c_299_n N_A_796_419#_c_864_n 0.00485793f $X=4.195 $Y=0.94
+ $X2=0 $Y2=0
cc_346 N_A_252_396#_c_300_n N_A_796_419#_c_864_n 0.00158217f $X=4.195 $Y=1.02
+ $X2=0 $Y2=0
cc_347 N_A_252_396#_c_303_n N_VPWR_c_1081_n 0.00507552f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_348 N_A_252_396#_c_305_n N_VPWR_c_1082_n 0.00397509f $X=4.395 $Y=2.01 $X2=0
+ $Y2=0
cc_349 N_A_252_396#_c_303_n N_VPWR_c_1085_n 0.00599768f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_350 N_A_252_396#_c_305_n N_VPWR_c_1086_n 0.00939541f $X=4.395 $Y=2.01 $X2=0
+ $Y2=0
cc_351 N_A_252_396#_c_303_n N_VPWR_c_1079_n 0.00973979f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_352 N_A_252_396#_c_305_n N_VPWR_c_1079_n 0.0161763f $X=4.395 $Y=2.01 $X2=0
+ $Y2=0
cc_353 N_A_252_396#_c_295_n N_VGND_c_1232_n 0.0151574f $X=1.86 $Y=0.55 $X2=0
+ $Y2=0
cc_354 N_A_252_396#_M1021_g N_VGND_c_1233_n 0.00547815f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_355 N_A_252_396#_M1007_g N_VGND_c_1233_n 0.00486043f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_356 N_A_252_396#_c_295_n N_VGND_c_1233_n 0.013514f $X=1.86 $Y=0.55 $X2=0
+ $Y2=0
cc_357 N_A_252_396#_M1021_g N_VGND_c_1234_n 0.00240189f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_252_396#_M1007_g N_VGND_c_1234_n 0.0134651f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_359 N_A_252_396#_c_296_n N_VGND_c_1234_n 0.0255241f $X=4.03 $Y=0.94 $X2=0
+ $Y2=0
cc_360 N_A_252_396#_M1012_g N_VGND_c_1239_n 0.00585385f $X=4.105 $Y=0.445 $X2=0
+ $Y2=0
cc_361 N_A_252_396#_M1021_g N_VGND_c_1243_n 0.00756669f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_362 N_A_252_396#_M1007_g N_VGND_c_1243_n 0.00443987f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_363 N_A_252_396#_M1012_g N_VGND_c_1243_n 0.00682102f $X=4.105 $Y=0.445 $X2=0
+ $Y2=0
cc_364 N_A_252_396#_c_292_n N_VGND_c_1243_n 6.06194e-19 $X=2.995 $Y=0.93 $X2=0
+ $Y2=0
cc_365 N_A_252_396#_c_295_n N_VGND_c_1243_n 0.00995894f $X=1.86 $Y=0.55 $X2=0
+ $Y2=0
cc_366 N_A_252_396#_c_296_n N_VGND_c_1243_n 0.0316578f $X=4.03 $Y=0.94 $X2=0
+ $Y2=0
cc_367 N_A_252_396#_c_297_n N_VGND_c_1243_n 0.00356796f $X=2.595 $Y=1.02 $X2=0
+ $Y2=0
cc_368 N_A_252_396#_c_299_n N_VGND_c_1243_n 0.00814301f $X=4.195 $Y=0.94 $X2=0
+ $Y2=0
cc_369 N_A_27_68#_c_450_n N_A_451_419#_M1017_s 0.00564752f $X=2.665 $Y=2.98
+ $X2=0 $Y2=0
cc_370 N_A_27_68#_c_452_n N_A_451_419#_M1000_g 6.80311e-19 $X=3.225 $Y=2.14
+ $X2=0 $Y2=0
cc_371 N_A_27_68#_c_442_n N_A_451_419#_M1000_g 0.00198073f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_372 N_A_27_68#_c_443_n N_A_451_419#_M1000_g 0.0821494f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_373 N_A_27_68#_c_450_n N_A_451_419#_c_577_n 0.0247944f $X=2.665 $Y=2.98 $X2=0
+ $Y2=0
cc_374 N_A_27_68#_c_453_n N_A_451_419#_c_577_n 0.00841003f $X=2.835 $Y=2.14
+ $X2=0 $Y2=0
cc_375 N_A_27_68#_c_443_n N_A_451_419#_c_577_n 2.28825e-19 $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_376 N_A_27_68#_c_452_n N_A_451_419#_c_578_n 0.0164153f $X=3.225 $Y=2.14 $X2=0
+ $Y2=0
cc_377 N_A_27_68#_c_453_n N_A_451_419#_c_578_n 0.0127426f $X=2.835 $Y=2.14 $X2=0
+ $Y2=0
cc_378 N_A_27_68#_c_442_n N_A_451_419#_c_578_n 0.0135289f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_379 N_A_27_68#_c_443_n N_A_451_419#_c_578_n 0.00157856f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_380 N_A_27_68#_c_442_n N_A_451_419#_c_565_n 0.00704355f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_381 N_A_27_68#_c_443_n N_A_451_419#_c_565_n 8.24224e-19 $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_382 N_A_27_68#_c_446_n N_A_451_419#_c_565_n 0.00188238f $X=3.325 $Y=1.605
+ $X2=0 $Y2=0
cc_383 N_A_27_68#_c_439_n N_A_451_419#_c_566_n 0.00106725f $X=3.64 $Y=0.805
+ $X2=0 $Y2=0
cc_384 N_A_27_68#_c_452_n N_A_451_419#_c_566_n 0.00538303f $X=3.225 $Y=2.14
+ $X2=0 $Y2=0
cc_385 N_A_27_68#_c_442_n N_A_451_419#_c_566_n 0.0194099f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_386 N_A_27_68#_c_443_n N_A_451_419#_c_566_n 0.00254894f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_387 N_A_27_68#_c_446_n N_A_451_419#_c_566_n 0.0132717f $X=3.325 $Y=1.605
+ $X2=0 $Y2=0
cc_388 N_A_27_68#_c_439_n N_A_451_419#_c_571_n 4.10172e-19 $X=3.64 $Y=0.805
+ $X2=0 $Y2=0
cc_389 N_A_27_68#_c_442_n N_A_451_419#_c_571_n 0.0108501f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_390 N_A_27_68#_c_443_n N_A_451_419#_c_571_n 8.58022e-19 $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_391 N_A_27_68#_c_446_n N_A_451_419#_c_571_n 0.00202608f $X=3.325 $Y=1.605
+ $X2=0 $Y2=0
cc_392 N_A_27_68#_c_439_n N_A_451_419#_c_572_n 0.00149818f $X=3.64 $Y=0.805
+ $X2=0 $Y2=0
cc_393 N_A_27_68#_c_443_n N_A_451_419#_c_572_n 0.00940465f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_394 N_A_27_68#_c_446_n N_A_451_419#_c_572_n 0.0090275f $X=3.325 $Y=1.605
+ $X2=0 $Y2=0
cc_395 N_A_27_68#_M1020_g N_A_796_419#_c_876_n 0.00358544f $X=3.365 $Y=2.595
+ $X2=0 $Y2=0
cc_396 N_A_27_68#_c_452_n N_A_796_419#_c_876_n 6.73957e-19 $X=3.225 $Y=2.14
+ $X2=0 $Y2=0
cc_397 N_A_27_68#_c_452_n N_A_796_419#_c_872_n 0.00547397f $X=3.225 $Y=2.14
+ $X2=0 $Y2=0
cc_398 N_A_27_68#_c_442_n N_A_796_419#_c_872_n 6.63768e-19 $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_399 N_A_27_68#_c_461_n N_VPWR_M1013_d 0.00725427f $X=1.215 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_400 N_A_27_68#_c_452_n N_VPWR_M1017_d 0.00889375f $X=3.225 $Y=2.14 $X2=0
+ $Y2=0
cc_401 N_A_27_68#_c_449_n N_VPWR_c_1080_n 0.0174373f $X=0.34 $Y=2.835 $X2=0
+ $Y2=0
cc_402 N_A_27_68#_c_461_n N_VPWR_c_1080_n 0.0157965f $X=1.215 $Y=2.475 $X2=0
+ $Y2=0
cc_403 N_A_27_68#_c_463_n N_VPWR_c_1080_n 0.0105407f $X=1.3 $Y=2.895 $X2=0 $Y2=0
cc_404 N_A_27_68#_c_451_n N_VPWR_c_1080_n 0.0129587f $X=1.385 $Y=2.98 $X2=0
+ $Y2=0
cc_405 N_A_27_68#_M1020_g N_VPWR_c_1081_n 0.0185889f $X=3.365 $Y=2.595 $X2=0
+ $Y2=0
cc_406 N_A_27_68#_c_452_n N_VPWR_c_1081_n 0.0149038f $X=3.225 $Y=2.14 $X2=0
+ $Y2=0
cc_407 N_A_27_68#_c_450_n N_VPWR_c_1085_n 0.0849142f $X=2.665 $Y=2.98 $X2=0
+ $Y2=0
cc_408 N_A_27_68#_c_451_n N_VPWR_c_1085_n 0.0113001f $X=1.385 $Y=2.98 $X2=0
+ $Y2=0
cc_409 N_A_27_68#_M1020_g N_VPWR_c_1086_n 0.008763f $X=3.365 $Y=2.595 $X2=0
+ $Y2=0
cc_410 N_A_27_68#_M1020_g N_VPWR_c_1079_n 0.0144563f $X=3.365 $Y=2.595 $X2=0
+ $Y2=0
cc_411 N_A_27_68#_c_449_n N_VPWR_c_1079_n 0.0153197f $X=0.34 $Y=2.835 $X2=0
+ $Y2=0
cc_412 N_A_27_68#_c_461_n N_VPWR_c_1079_n 0.0124161f $X=1.215 $Y=2.475 $X2=0
+ $Y2=0
cc_413 N_A_27_68#_c_450_n N_VPWR_c_1079_n 0.0532597f $X=2.665 $Y=2.98 $X2=0
+ $Y2=0
cc_414 N_A_27_68#_c_451_n N_VPWR_c_1079_n 0.00636923f $X=1.385 $Y=2.98 $X2=0
+ $Y2=0
cc_415 N_A_27_68#_c_449_n N_VPWR_c_1091_n 0.0199586f $X=0.34 $Y=2.835 $X2=0
+ $Y2=0
cc_416 N_A_27_68#_c_444_n N_VGND_c_1232_n 0.0154769f $X=0.28 $Y=0.55 $X2=0 $Y2=0
cc_417 N_A_27_68#_c_440_n N_VGND_c_1234_n 0.00201563f $X=3.46 $Y=0.805 $X2=0
+ $Y2=0
cc_418 N_A_27_68#_c_441_n N_VGND_c_1234_n 0.0123433f $X=3.715 $Y=0.73 $X2=0
+ $Y2=0
cc_419 N_A_27_68#_c_444_n N_VGND_c_1238_n 0.0175663f $X=0.28 $Y=0.55 $X2=0 $Y2=0
cc_420 N_A_27_68#_c_440_n N_VGND_c_1239_n 0.00465854f $X=3.46 $Y=0.805 $X2=0
+ $Y2=0
cc_421 N_A_27_68#_c_441_n N_VGND_c_1239_n 0.00585385f $X=3.715 $Y=0.73 $X2=0
+ $Y2=0
cc_422 N_A_27_68#_c_440_n N_VGND_c_1243_n 0.00623841f $X=3.46 $Y=0.805 $X2=0
+ $Y2=0
cc_423 N_A_27_68#_c_441_n N_VGND_c_1243_n 0.00710641f $X=3.715 $Y=0.73 $X2=0
+ $Y2=0
cc_424 N_A_27_68#_c_444_n N_VGND_c_1243_n 0.0130705f $X=0.28 $Y=0.55 $X2=0 $Y2=0
cc_425 N_A_451_419#_M1022_g N_A_952_305#_M1029_g 0.0272389f $X=4.675 $Y=0.445
+ $X2=0 $Y2=0
cc_426 N_A_451_419#_c_568_n N_A_952_305#_M1029_g 7.0348e-19 $X=4.6 $Y=1.51 $X2=0
+ $Y2=0
cc_427 N_A_451_419#_c_569_n N_A_952_305#_M1029_g 8.2093e-19 $X=4.685 $Y=1.425
+ $X2=0 $Y2=0
cc_428 N_A_451_419#_c_573_n N_A_952_305#_M1029_g 4.09151e-19 $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_429 N_A_451_419#_c_574_n N_A_952_305#_M1029_g 0.020616f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_430 N_A_451_419#_c_573_n N_A_952_305#_c_708_n 0.019019f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_431 N_A_451_419#_c_574_n N_A_952_305#_c_708_n 0.00155751f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_432 N_A_451_419#_c_568_n N_A_952_305#_c_710_n 0.00500321f $X=4.6 $Y=1.51
+ $X2=0 $Y2=0
cc_433 N_A_451_419#_c_568_n N_A_952_305#_c_711_n 0.00504036f $X=4.6 $Y=1.51
+ $X2=0 $Y2=0
cc_434 N_A_451_419#_c_569_n N_A_952_305#_c_711_n 0.00628872f $X=4.685 $Y=1.425
+ $X2=0 $Y2=0
cc_435 N_A_451_419#_c_573_n N_A_952_305#_c_711_n 0.00538911f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_436 N_A_451_419#_c_574_n N_A_952_305#_c_711_n 4.21682e-19 $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_437 N_A_451_419#_c_568_n N_A_952_305#_c_715_n 0.00223279f $X=4.6 $Y=1.51
+ $X2=0 $Y2=0
cc_438 N_A_451_419#_c_573_n N_A_952_305#_c_715_n 0.00120658f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_439 N_A_451_419#_c_574_n N_A_952_305#_c_715_n 0.00962379f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_440 N_A_451_419#_M1000_g N_A_796_419#_c_876_n 0.0196421f $X=3.855 $Y=2.595
+ $X2=0 $Y2=0
cc_441 N_A_451_419#_c_568_n N_A_796_419#_c_871_n 0.017454f $X=4.6 $Y=1.51 $X2=0
+ $Y2=0
cc_442 N_A_451_419#_M1000_g N_A_796_419#_c_872_n 0.00407559f $X=3.855 $Y=2.595
+ $X2=0 $Y2=0
cc_443 N_A_451_419#_c_568_n N_A_796_419#_c_872_n 0.0112252f $X=4.6 $Y=1.51 $X2=0
+ $Y2=0
cc_444 N_A_451_419#_c_571_n N_A_796_419#_c_872_n 0.00372187f $X=3.855 $Y=1.51
+ $X2=0 $Y2=0
cc_445 N_A_451_419#_c_572_n N_A_796_419#_c_872_n 3.72389e-19 $X=3.865 $Y=1.59
+ $X2=0 $Y2=0
cc_446 N_A_451_419#_M1022_g N_A_796_419#_c_863_n 0.00454824f $X=4.675 $Y=0.445
+ $X2=0 $Y2=0
cc_447 N_A_451_419#_c_573_n N_A_796_419#_c_863_n 0.0158849f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_448 N_A_451_419#_c_574_n N_A_796_419#_c_863_n 0.00124625f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_449 N_A_451_419#_M1022_g N_A_796_419#_c_864_n 0.0143689f $X=4.675 $Y=0.445
+ $X2=0 $Y2=0
cc_450 N_A_451_419#_c_568_n N_A_796_419#_c_864_n 0.00192133f $X=4.6 $Y=1.51
+ $X2=0 $Y2=0
cc_451 N_A_451_419#_c_573_n N_A_796_419#_c_864_n 0.0085796f $X=4.765 $Y=1.12
+ $X2=0 $Y2=0
cc_452 N_A_451_419#_M1000_g N_VPWR_c_1081_n 0.00388058f $X=3.855 $Y=2.595 $X2=0
+ $Y2=0
cc_453 N_A_451_419#_M1000_g N_VPWR_c_1086_n 0.00954582f $X=3.855 $Y=2.595 $X2=0
+ $Y2=0
cc_454 N_A_451_419#_M1017_s N_VPWR_c_1079_n 0.00233022f $X=2.255 $Y=2.095 $X2=0
+ $Y2=0
cc_455 N_A_451_419#_M1000_g N_VPWR_c_1079_n 0.0165468f $X=3.855 $Y=2.595 $X2=0
+ $Y2=0
cc_456 N_A_451_419#_c_570_n N_VGND_c_1233_n 0.026255f $X=2.42 $Y=0.47 $X2=0
+ $Y2=0
cc_457 N_A_451_419#_c_570_n N_VGND_c_1234_n 0.0139887f $X=2.42 $Y=0.47 $X2=0
+ $Y2=0
cc_458 N_A_451_419#_M1022_g N_VGND_c_1239_n 0.00375982f $X=4.675 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_A_451_419#_M1021_s N_VGND_c_1243_n 0.00233022f $X=2.275 $Y=0.235 $X2=0
+ $Y2=0
cc_460 N_A_451_419#_M1022_g N_VGND_c_1243_n 0.00620332f $X=4.675 $Y=0.445 $X2=0
+ $Y2=0
cc_461 N_A_451_419#_c_570_n N_VGND_c_1243_n 0.0166743f $X=2.42 $Y=0.47 $X2=0
+ $Y2=0
cc_462 N_A_952_305#_M1026_g N_A_796_419#_M1005_g 0.0161037f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_463 N_A_952_305#_c_720_n N_A_796_419#_M1005_g 0.0205565f $X=5.99 $Y=2.24
+ $X2=0 $Y2=0
cc_464 N_A_952_305#_c_744_p N_A_796_419#_M1005_g 0.00803707f $X=6.155 $Y=2.785
+ $X2=0 $Y2=0
cc_465 N_A_952_305#_c_712_n N_A_796_419#_c_862_n 0.00752537f $X=6.095 $Y=1.04
+ $X2=0 $Y2=0
cc_466 N_A_952_305#_c_713_n N_A_796_419#_c_862_n 0.00792203f $X=6.845 $Y=1.44
+ $X2=0 $Y2=0
cc_467 N_A_952_305#_M1026_g N_A_796_419#_c_876_n 0.00371531f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_468 N_A_952_305#_M1026_g N_A_796_419#_c_871_n 0.028309f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_469 N_A_952_305#_c_720_n N_A_796_419#_c_871_n 0.00990958f $X=5.99 $Y=2.24
+ $X2=0 $Y2=0
cc_470 N_A_952_305#_c_710_n N_A_796_419#_c_871_n 0.0242646f $X=5.13 $Y=1.69
+ $X2=0 $Y2=0
cc_471 N_A_952_305#_c_715_n N_A_796_419#_c_871_n 0.00292987f $X=5.215 $Y=1.69
+ $X2=0 $Y2=0
cc_472 N_A_952_305#_M1029_g N_A_796_419#_c_863_n 0.013037f $X=5.215 $Y=0.445
+ $X2=0 $Y2=0
cc_473 N_A_952_305#_c_708_n N_A_796_419#_c_863_n 0.0125335f $X=5.295 $Y=1.08
+ $X2=0 $Y2=0
cc_474 N_A_952_305#_c_712_n N_A_796_419#_c_863_n 0.0407129f $X=6.095 $Y=1.04
+ $X2=0 $Y2=0
cc_475 N_A_952_305#_M1026_g N_A_796_419#_c_873_n 0.00235648f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_476 N_A_952_305#_M1029_g N_A_796_419#_c_864_n 0.00154872f $X=5.215 $Y=0.445
+ $X2=0 $Y2=0
cc_477 N_A_952_305#_M1026_g N_A_796_419#_c_865_n 7.61128e-19 $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_478 N_A_952_305#_c_720_n N_A_796_419#_c_865_n 0.00506068f $X=5.99 $Y=2.24
+ $X2=0 $Y2=0
cc_479 N_A_952_305#_c_710_n N_A_796_419#_c_865_n 0.0224186f $X=5.13 $Y=1.69
+ $X2=0 $Y2=0
cc_480 N_A_952_305#_c_712_n N_A_796_419#_c_865_n 0.0181148f $X=6.095 $Y=1.04
+ $X2=0 $Y2=0
cc_481 N_A_952_305#_c_715_n N_A_796_419#_c_865_n 0.00201464f $X=5.215 $Y=1.69
+ $X2=0 $Y2=0
cc_482 N_A_952_305#_M1026_g N_A_796_419#_c_866_n 6.72839e-19 $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_483 N_A_952_305#_c_720_n N_A_796_419#_c_866_n 0.00104429f $X=5.99 $Y=2.24
+ $X2=0 $Y2=0
cc_484 N_A_952_305#_c_710_n N_A_796_419#_c_866_n 2.99648e-19 $X=5.13 $Y=1.69
+ $X2=0 $Y2=0
cc_485 N_A_952_305#_c_712_n N_A_796_419#_c_866_n 0.00398877f $X=6.095 $Y=1.04
+ $X2=0 $Y2=0
cc_486 N_A_952_305#_c_715_n N_A_796_419#_c_866_n 0.0158582f $X=5.215 $Y=1.69
+ $X2=0 $Y2=0
cc_487 N_A_952_305#_M1024_s N_A_796_419#_c_867_n 0.00248891f $X=5.955 $Y=0.765
+ $X2=0 $Y2=0
cc_488 N_A_952_305#_M1029_g N_A_796_419#_c_867_n 9.14714e-19 $X=5.215 $Y=0.445
+ $X2=0 $Y2=0
cc_489 N_A_952_305#_c_712_n N_A_796_419#_c_867_n 0.0253293f $X=6.095 $Y=1.04
+ $X2=0 $Y2=0
cc_490 N_A_952_305#_M1029_g N_A_796_419#_c_868_n 0.0311791f $X=5.215 $Y=0.445
+ $X2=0 $Y2=0
cc_491 N_A_952_305#_c_712_n N_A_796_419#_c_868_n 9.47502e-19 $X=6.095 $Y=1.04
+ $X2=0 $Y2=0
cc_492 N_A_952_305#_c_710_n N_A_796_419#_c_869_n 2.15142e-19 $X=5.13 $Y=1.69
+ $X2=0 $Y2=0
cc_493 N_A_952_305#_c_711_n N_A_796_419#_c_869_n 0.00515145f $X=5.13 $Y=1.525
+ $X2=0 $Y2=0
cc_494 N_A_952_305#_c_712_n N_A_796_419#_c_869_n 0.0204785f $X=6.095 $Y=1.04
+ $X2=0 $Y2=0
cc_495 N_A_952_305#_c_715_n N_A_796_419#_c_869_n 0.00135098f $X=5.215 $Y=1.69
+ $X2=0 $Y2=0
cc_496 N_A_952_305#_c_720_n N_RESET_B_M1028_g 0.0193574f $X=5.99 $Y=2.24 $X2=0
+ $Y2=0
cc_497 N_A_952_305#_c_777_p N_RESET_B_M1028_g 0.0198884f $X=6.845 $Y=2.785 $X2=0
+ $Y2=0
cc_498 N_A_952_305#_c_744_p N_RESET_B_M1028_g 0.00937074f $X=6.155 $Y=2.785
+ $X2=0 $Y2=0
cc_499 N_A_952_305#_c_709_n N_RESET_B_M1028_g 0.00698955f $X=6.93 $Y=2.7 $X2=0
+ $Y2=0
cc_500 N_A_952_305#_c_700_n N_RESET_B_M1010_g 0.0152567f $X=7.1 $Y=1.295 $X2=0
+ $Y2=0
cc_501 N_A_952_305#_c_712_n N_RESET_B_M1010_g 0.00140579f $X=6.095 $Y=1.04 $X2=0
+ $Y2=0
cc_502 N_A_952_305#_c_713_n N_RESET_B_M1010_g 0.0167205f $X=6.845 $Y=1.44 $X2=0
+ $Y2=0
cc_503 N_A_952_305#_c_714_n N_RESET_B_M1010_g 0.0050844f $X=7.165 $Y=1.46 $X2=0
+ $Y2=0
cc_504 N_A_952_305#_c_716_n N_RESET_B_M1010_g 0.0158987f $X=7.75 $Y=1.46 $X2=0
+ $Y2=0
cc_505 N_A_952_305#_c_720_n N_RESET_B_c_973_n 0.0318988f $X=5.99 $Y=2.24 $X2=0
+ $Y2=0
cc_506 N_A_952_305#_c_777_p N_RESET_B_c_973_n 0.020152f $X=6.845 $Y=2.785 $X2=0
+ $Y2=0
cc_507 N_A_952_305#_c_709_n N_RESET_B_c_973_n 0.0656264f $X=6.93 $Y=2.7 $X2=0
+ $Y2=0
cc_508 N_A_952_305#_c_713_n N_RESET_B_c_973_n 0.0248367f $X=6.845 $Y=1.44 $X2=0
+ $Y2=0
cc_509 N_A_952_305#_c_714_n N_RESET_B_c_973_n 0.00149249f $X=7.165 $Y=1.46 $X2=0
+ $Y2=0
cc_510 N_A_952_305#_c_709_n N_RESET_B_c_974_n 0.00862438f $X=6.93 $Y=2.7 $X2=0
+ $Y2=0
cc_511 N_A_952_305#_c_712_n N_RESET_B_c_974_n 0.00511633f $X=6.095 $Y=1.04 $X2=0
+ $Y2=0
cc_512 N_A_952_305#_c_713_n N_RESET_B_c_974_n 0.00328942f $X=6.845 $Y=1.44 $X2=0
+ $Y2=0
cc_513 N_A_952_305#_M1006_g N_A_1617_76#_M1023_g 0.0210576f $X=8.8 $Y=0.59 $X2=0
+ $Y2=0
cc_514 N_A_952_305#_c_707_n N_A_1617_76#_c_1015_n 0.0210576f $X=8.8 $Y=1.37
+ $X2=0 $Y2=0
cc_515 N_A_952_305#_M1027_g N_A_1617_76#_c_1016_n 0.0210576f $X=8.75 $Y=2.37
+ $X2=0 $Y2=0
cc_516 N_A_952_305#_M1004_g N_A_1617_76#_c_1017_n 0.00610891f $X=8.44 $Y=0.59
+ $X2=0 $Y2=0
cc_517 N_A_952_305#_c_703_n N_A_1617_76#_c_1018_n 0.00812265f $X=8.365 $Y=1.37
+ $X2=0 $Y2=0
cc_518 N_A_952_305#_M1004_g N_A_1617_76#_c_1018_n 0.00446336f $X=8.44 $Y=0.59
+ $X2=0 $Y2=0
cc_519 N_A_952_305#_M1027_g N_A_1617_76#_c_1018_n 0.035433f $X=8.75 $Y=2.37
+ $X2=0 $Y2=0
cc_520 N_A_952_305#_M1006_g N_A_1617_76#_c_1018_n 0.00142801f $X=8.8 $Y=0.59
+ $X2=0 $Y2=0
cc_521 N_A_952_305#_c_707_n N_A_1617_76#_c_1018_n 0.0114797f $X=8.8 $Y=1.37
+ $X2=0 $Y2=0
cc_522 N_A_952_305#_c_716_n N_A_1617_76#_c_1018_n 0.00444532f $X=7.75 $Y=1.46
+ $X2=0 $Y2=0
cc_523 N_A_952_305#_M1006_g N_A_1617_76#_c_1019_n 0.0183825f $X=8.8 $Y=0.59
+ $X2=0 $Y2=0
cc_524 N_A_952_305#_c_701_n N_A_1617_76#_c_1020_n 0.00301769f $X=7.46 $Y=1.295
+ $X2=0 $Y2=0
cc_525 N_A_952_305#_c_703_n N_A_1617_76#_c_1020_n 0.00489384f $X=8.365 $Y=1.37
+ $X2=0 $Y2=0
cc_526 N_A_952_305#_M1004_g N_A_1617_76#_c_1020_n 0.00948225f $X=8.44 $Y=0.59
+ $X2=0 $Y2=0
cc_527 N_A_952_305#_M1006_g N_A_1617_76#_c_1020_n 0.00221647f $X=8.8 $Y=0.59
+ $X2=0 $Y2=0
cc_528 N_A_952_305#_M1004_g N_A_1617_76#_c_1021_n 0.0125397f $X=8.44 $Y=0.59
+ $X2=0 $Y2=0
cc_529 N_A_952_305#_M1006_g N_A_1617_76#_c_1022_n 0.00213442f $X=8.8 $Y=0.59
+ $X2=0 $Y2=0
cc_530 N_A_952_305#_c_777_p N_VPWR_M1028_d 0.0232819f $X=6.845 $Y=2.785 $X2=0
+ $Y2=0
cc_531 N_A_952_305#_c_709_n N_VPWR_M1028_d 0.0181798f $X=6.93 $Y=2.7 $X2=0 $Y2=0
cc_532 N_A_952_305#_M1026_g N_VPWR_c_1082_n 0.019954f $X=4.885 $Y=2.595 $X2=0
+ $Y2=0
cc_533 N_A_952_305#_c_720_n N_VPWR_c_1082_n 0.0103902f $X=5.99 $Y=2.24 $X2=0
+ $Y2=0
cc_534 N_A_952_305#_c_744_p N_VPWR_c_1082_n 0.0123852f $X=6.155 $Y=2.785 $X2=0
+ $Y2=0
cc_535 N_A_952_305#_M1001_g N_VPWR_c_1083_n 0.0252947f $X=7.625 $Y=2.595 $X2=0
+ $Y2=0
cc_536 N_A_952_305#_c_777_p N_VPWR_c_1083_n 0.0138719f $X=6.845 $Y=2.785 $X2=0
+ $Y2=0
cc_537 N_A_952_305#_c_709_n N_VPWR_c_1083_n 0.0458f $X=6.93 $Y=2.7 $X2=0 $Y2=0
cc_538 N_A_952_305#_c_714_n N_VPWR_c_1083_n 0.00550891f $X=7.165 $Y=1.46 $X2=0
+ $Y2=0
cc_539 N_A_952_305#_c_716_n N_VPWR_c_1083_n 0.00903609f $X=7.75 $Y=1.46 $X2=0
+ $Y2=0
cc_540 N_A_952_305#_M1027_g N_VPWR_c_1084_n 0.0266261f $X=8.75 $Y=2.37 $X2=0
+ $Y2=0
cc_541 N_A_952_305#_M1026_g N_VPWR_c_1086_n 0.008763f $X=4.885 $Y=2.595 $X2=0
+ $Y2=0
cc_542 N_A_952_305#_c_777_p N_VPWR_c_1087_n 0.0227869f $X=6.845 $Y=2.785 $X2=0
+ $Y2=0
cc_543 N_A_952_305#_c_744_p N_VPWR_c_1087_n 0.0179231f $X=6.155 $Y=2.785 $X2=0
+ $Y2=0
cc_544 N_A_952_305#_M1001_g N_VPWR_c_1088_n 0.00810115f $X=7.625 $Y=2.595 $X2=0
+ $Y2=0
cc_545 N_A_952_305#_M1027_g N_VPWR_c_1088_n 0.00747382f $X=8.75 $Y=2.37 $X2=0
+ $Y2=0
cc_546 N_A_952_305#_M1005_d N_VPWR_c_1079_n 0.00223819f $X=5.85 $Y=2.095 $X2=0
+ $Y2=0
cc_547 N_A_952_305#_M1026_g N_VPWR_c_1079_n 0.0144563f $X=4.885 $Y=2.595 $X2=0
+ $Y2=0
cc_548 N_A_952_305#_M1001_g N_VPWR_c_1079_n 0.0141561f $X=7.625 $Y=2.595 $X2=0
+ $Y2=0
cc_549 N_A_952_305#_M1027_g N_VPWR_c_1079_n 0.00779694f $X=8.75 $Y=2.37 $X2=0
+ $Y2=0
cc_550 N_A_952_305#_c_777_p N_VPWR_c_1079_n 0.0272561f $X=6.845 $Y=2.785 $X2=0
+ $Y2=0
cc_551 N_A_952_305#_c_744_p N_VPWR_c_1079_n 0.0123929f $X=6.155 $Y=2.785 $X2=0
+ $Y2=0
cc_552 N_A_952_305#_c_700_n N_Q_c_1181_n 0.00154458f $X=7.1 $Y=1.295 $X2=0 $Y2=0
cc_553 N_A_952_305#_c_701_n N_Q_c_1181_n 0.00843873f $X=7.46 $Y=1.295 $X2=0
+ $Y2=0
cc_554 N_A_952_305#_M1004_g N_Q_c_1181_n 0.0021139f $X=8.44 $Y=0.59 $X2=0 $Y2=0
cc_555 N_A_952_305#_c_701_n N_Q_c_1182_n 0.00221594f $X=7.46 $Y=1.295 $X2=0
+ $Y2=0
cc_556 N_A_952_305#_M1004_g N_Q_c_1182_n 6.28884e-19 $X=8.44 $Y=0.59 $X2=0 $Y2=0
cc_557 N_A_952_305#_c_716_n N_Q_c_1182_n 0.00401765f $X=7.75 $Y=1.46 $X2=0 $Y2=0
cc_558 N_A_952_305#_c_701_n Q 0.00273191f $X=7.46 $Y=1.295 $X2=0 $Y2=0
cc_559 N_A_952_305#_M1001_g Q 0.0546456f $X=7.625 $Y=2.595 $X2=0 $Y2=0
cc_560 N_A_952_305#_c_703_n Q 0.0174068f $X=8.365 $Y=1.37 $X2=0 $Y2=0
cc_561 N_A_952_305#_M1027_g Q 0.00567446f $X=8.75 $Y=2.37 $X2=0 $Y2=0
cc_562 N_A_952_305#_c_714_n Q 0.0156997f $X=7.165 $Y=1.46 $X2=0 $Y2=0
cc_563 N_A_952_305#_c_716_n Q 0.0131727f $X=7.75 $Y=1.46 $X2=0 $Y2=0
cc_564 N_A_952_305#_M1027_g N_Q_N_c_1212_n 2.74877e-19 $X=8.75 $Y=2.37 $X2=0
+ $Y2=0
cc_565 N_A_952_305#_M1029_g N_VGND_c_1235_n 0.00689783f $X=5.215 $Y=0.445 $X2=0
+ $Y2=0
cc_566 N_A_952_305#_c_700_n N_VGND_c_1236_n 0.0096192f $X=7.1 $Y=1.295 $X2=0
+ $Y2=0
cc_567 N_A_952_305#_c_701_n N_VGND_c_1236_n 0.00144992f $X=7.46 $Y=1.295 $X2=0
+ $Y2=0
cc_568 N_A_952_305#_c_712_n N_VGND_c_1236_n 0.00382056f $X=6.095 $Y=1.04 $X2=0
+ $Y2=0
cc_569 N_A_952_305#_c_713_n N_VGND_c_1236_n 0.0215957f $X=6.845 $Y=1.44 $X2=0
+ $Y2=0
cc_570 N_A_952_305#_M1004_g N_VGND_c_1237_n 0.00179299f $X=8.44 $Y=0.59 $X2=0
+ $Y2=0
cc_571 N_A_952_305#_M1006_g N_VGND_c_1237_n 0.0120741f $X=8.8 $Y=0.59 $X2=0
+ $Y2=0
cc_572 N_A_952_305#_M1029_g N_VGND_c_1239_n 0.00420601f $X=5.215 $Y=0.445 $X2=0
+ $Y2=0
cc_573 N_A_952_305#_c_700_n N_VGND_c_1241_n 0.00289826f $X=7.1 $Y=1.295 $X2=0
+ $Y2=0
cc_574 N_A_952_305#_c_701_n N_VGND_c_1241_n 0.00337154f $X=7.46 $Y=1.295 $X2=0
+ $Y2=0
cc_575 N_A_952_305#_M1004_g N_VGND_c_1241_n 0.00527781f $X=8.44 $Y=0.59 $X2=0
+ $Y2=0
cc_576 N_A_952_305#_M1006_g N_VGND_c_1241_n 0.0047441f $X=8.8 $Y=0.59 $X2=0
+ $Y2=0
cc_577 N_A_952_305#_M1029_g N_VGND_c_1243_n 0.00752048f $X=5.215 $Y=0.445 $X2=0
+ $Y2=0
cc_578 N_A_952_305#_c_700_n N_VGND_c_1243_n 0.00363223f $X=7.1 $Y=1.295 $X2=0
+ $Y2=0
cc_579 N_A_952_305#_c_701_n N_VGND_c_1243_n 0.00432409f $X=7.46 $Y=1.295 $X2=0
+ $Y2=0
cc_580 N_A_952_305#_M1004_g N_VGND_c_1243_n 0.00542671f $X=8.44 $Y=0.59 $X2=0
+ $Y2=0
cc_581 N_A_952_305#_M1006_g N_VGND_c_1243_n 0.00455844f $X=8.8 $Y=0.59 $X2=0
+ $Y2=0
cc_582 N_A_796_419#_c_871_n N_RESET_B_M1028_g 2.148e-19 $X=5.475 $Y=2.12 $X2=0
+ $Y2=0
cc_583 N_A_796_419#_c_866_n N_RESET_B_M1010_g 6.18407e-19 $X=5.725 $Y=1.73 $X2=0
+ $Y2=0
cc_584 N_A_796_419#_c_868_n N_RESET_B_M1010_g 0.0408593f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_585 N_A_796_419#_c_869_n N_RESET_B_M1010_g 0.00393524f $X=5.725 $Y=1.565
+ $X2=0 $Y2=0
cc_586 N_A_796_419#_M1005_g N_RESET_B_c_973_n 9.43546e-19 $X=5.725 $Y=2.595
+ $X2=0 $Y2=0
cc_587 N_A_796_419#_c_865_n N_RESET_B_c_973_n 0.0101473f $X=5.725 $Y=1.73 $X2=0
+ $Y2=0
cc_588 N_A_796_419#_c_866_n N_RESET_B_c_973_n 2.76197e-19 $X=5.725 $Y=1.73 $X2=0
+ $Y2=0
cc_589 N_A_796_419#_M1005_g N_RESET_B_c_974_n 0.0280157f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_590 N_A_796_419#_c_862_n N_RESET_B_c_974_n 0.00658209f $X=6.31 $Y=0.655 $X2=0
+ $Y2=0
cc_591 N_A_796_419#_c_873_n N_RESET_B_c_974_n 6.4147e-19 $X=5.56 $Y=2.035 $X2=0
+ $Y2=0
cc_592 N_A_796_419#_c_865_n N_RESET_B_c_974_n 0.001332f $X=5.725 $Y=1.73 $X2=0
+ $Y2=0
cc_593 N_A_796_419#_c_866_n N_RESET_B_c_974_n 0.0162323f $X=5.725 $Y=1.73 $X2=0
+ $Y2=0
cc_594 N_A_796_419#_c_871_n N_VPWR_M1026_d 0.012933f $X=5.475 $Y=2.12 $X2=0
+ $Y2=0
cc_595 N_A_796_419#_M1005_g N_VPWR_c_1082_n 0.0103029f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_596 N_A_796_419#_c_871_n N_VPWR_c_1082_n 0.0209601f $X=5.475 $Y=2.12 $X2=0
+ $Y2=0
cc_597 N_A_796_419#_c_876_n N_VPWR_c_1086_n 0.0178162f $X=4.13 $Y=2.24 $X2=0
+ $Y2=0
cc_598 N_A_796_419#_M1005_g N_VPWR_c_1087_n 0.00938036f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_599 N_A_796_419#_M1000_d N_VPWR_c_1079_n 0.0023187f $X=3.98 $Y=2.095 $X2=0
+ $Y2=0
cc_600 N_A_796_419#_M1005_g N_VPWR_c_1079_n 0.0168486f $X=5.725 $Y=2.595 $X2=0
+ $Y2=0
cc_601 N_A_796_419#_c_876_n N_VPWR_c_1079_n 0.0123708f $X=4.13 $Y=2.24 $X2=0
+ $Y2=0
cc_602 N_A_796_419#_c_871_n A_904_419# 0.0048076f $X=5.475 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_603 N_A_796_419#_c_863_n N_VGND_M1029_d 0.00336501f $X=5.855 $Y=0.69 $X2=0
+ $Y2=0
cc_604 N_A_796_419#_c_863_n N_VGND_c_1235_n 0.0235175f $X=5.855 $Y=0.69 $X2=0
+ $Y2=0
cc_605 N_A_796_419#_c_867_n N_VGND_c_1235_n 0.00758005f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_606 N_A_796_419#_c_868_n N_VGND_c_1235_n 0.00113758f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_607 N_A_796_419#_c_867_n N_VGND_c_1236_n 0.0147375f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_608 N_A_796_419#_c_868_n N_VGND_c_1236_n 0.00822975f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_609 N_A_796_419#_c_863_n N_VGND_c_1239_n 0.0102604f $X=5.855 $Y=0.69 $X2=0
+ $Y2=0
cc_610 N_A_796_419#_c_864_n N_VGND_c_1239_n 0.0246051f $X=4.46 $Y=0.47 $X2=0
+ $Y2=0
cc_611 N_A_796_419#_c_863_n N_VGND_c_1240_n 0.00325096f $X=5.855 $Y=0.69 $X2=0
+ $Y2=0
cc_612 N_A_796_419#_c_867_n N_VGND_c_1240_n 0.0148168f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_613 N_A_796_419#_c_868_n N_VGND_c_1240_n 0.0107095f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_614 N_A_796_419#_M1012_d N_VGND_c_1243_n 0.00417932f $X=4.18 $Y=0.235 $X2=0
+ $Y2=0
cc_615 N_A_796_419#_c_863_n N_VGND_c_1243_n 0.0243775f $X=5.855 $Y=0.69 $X2=0
+ $Y2=0
cc_616 N_A_796_419#_c_864_n N_VGND_c_1243_n 0.0153758f $X=4.46 $Y=0.47 $X2=0
+ $Y2=0
cc_617 N_A_796_419#_c_867_n N_VGND_c_1243_n 0.011889f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_618 N_A_796_419#_c_868_n N_VGND_c_1243_n 0.0106168f $X=6.02 $Y=0.49 $X2=0
+ $Y2=0
cc_619 N_A_796_419#_c_863_n A_950_47# 0.00471833f $X=5.855 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_620 N_RESET_B_c_973_n N_VPWR_M1028_d 0.00960281f $X=6.5 $Y=1.77 $X2=0 $Y2=0
cc_621 N_RESET_B_M1028_g N_VPWR_c_1087_n 0.00655523f $X=6.255 $Y=2.595 $X2=0
+ $Y2=0
cc_622 N_RESET_B_M1028_g N_VPWR_c_1079_n 0.00960922f $X=6.255 $Y=2.595 $X2=0
+ $Y2=0
cc_623 N_RESET_B_M1010_g N_VGND_c_1236_n 0.00987521f $X=6.67 $Y=0.975 $X2=0
+ $Y2=0
cc_624 N_RESET_B_M1010_g N_VGND_c_1240_n 0.00289826f $X=6.67 $Y=0.975 $X2=0
+ $Y2=0
cc_625 N_RESET_B_M1010_g N_VGND_c_1243_n 0.00363223f $X=6.67 $Y=0.975 $X2=0
+ $Y2=0
cc_626 N_A_1617_76#_M1016_g N_VPWR_c_1084_n 0.0257226f $X=9.28 $Y=2.37 $X2=0
+ $Y2=0
cc_627 N_A_1617_76#_c_1018_n N_VPWR_c_1084_n 0.0697491f $X=8.485 $Y=2.015 $X2=0
+ $Y2=0
cc_628 N_A_1617_76#_c_1022_n N_VPWR_c_1084_n 0.00185662f $X=9.32 $Y=1.165 $X2=0
+ $Y2=0
cc_629 N_A_1617_76#_c_1018_n N_VPWR_c_1088_n 0.0134413f $X=8.485 $Y=2.015 $X2=0
+ $Y2=0
cc_630 N_A_1617_76#_M1016_g N_VPWR_c_1089_n 0.00747382f $X=9.28 $Y=2.37 $X2=0
+ $Y2=0
cc_631 N_A_1617_76#_M1016_g N_VPWR_c_1079_n 0.00779694f $X=9.28 $Y=2.37 $X2=0
+ $Y2=0
cc_632 N_A_1617_76#_c_1018_n N_VPWR_c_1079_n 0.0143765f $X=8.485 $Y=2.015 $X2=0
+ $Y2=0
cc_633 N_A_1617_76#_c_1017_n N_Q_c_1181_n 0.00851846f $X=8.32 $Y=1 $X2=0 $Y2=0
cc_634 N_A_1617_76#_c_1018_n N_Q_c_1181_n 4.57377e-19 $X=8.485 $Y=2.015 $X2=0
+ $Y2=0
cc_635 N_A_1617_76#_c_1020_n N_Q_c_1181_n 0.00594923f $X=8.225 $Y=0.59 $X2=0
+ $Y2=0
cc_636 N_A_1617_76#_c_1021_n N_Q_c_1181_n 0.00899597f $X=8.442 $Y=1.085 $X2=0
+ $Y2=0
cc_637 N_A_1617_76#_c_1018_n N_Q_c_1182_n 0.138549f $X=8.485 $Y=2.015 $X2=0
+ $Y2=0
cc_638 N_A_1617_76#_M1023_g N_Q_N_c_1209_n 0.00125204f $X=9.23 $Y=0.59 $X2=0
+ $Y2=0
cc_639 N_A_1617_76#_M1025_g N_Q_N_c_1209_n 0.0100697f $X=9.59 $Y=0.59 $X2=0
+ $Y2=0
cc_640 N_A_1617_76#_M1016_g Q_N 0.0134647f $X=9.28 $Y=2.37 $X2=0 $Y2=0
cc_641 N_A_1617_76#_M1016_g N_Q_N_c_1212_n 0.00584696f $X=9.28 $Y=2.37 $X2=0
+ $Y2=0
cc_642 N_A_1617_76#_c_1015_n N_Q_N_c_1212_n 0.00505259f $X=9.59 $Y=1.075 $X2=0
+ $Y2=0
cc_643 N_A_1617_76#_c_1016_n N_Q_N_c_1212_n 6.13565e-19 $X=9.32 $Y=1.67 $X2=0
+ $Y2=0
cc_644 N_A_1617_76#_c_1022_n N_Q_N_c_1212_n 0.00867382f $X=9.32 $Y=1.165 $X2=0
+ $Y2=0
cc_645 N_A_1617_76#_M1016_g N_Q_N_c_1210_n 0.00370596f $X=9.28 $Y=2.37 $X2=0
+ $Y2=0
cc_646 N_A_1617_76#_M1025_g N_Q_N_c_1210_n 0.00869848f $X=9.59 $Y=0.59 $X2=0
+ $Y2=0
cc_647 N_A_1617_76#_c_1022_n N_Q_N_c_1210_n 0.0321883f $X=9.32 $Y=1.165 $X2=0
+ $Y2=0
cc_648 N_A_1617_76#_c_1023_n N_Q_N_c_1210_n 0.0102238f $X=9.32 $Y=1.165 $X2=0
+ $Y2=0
cc_649 N_A_1617_76#_M1023_g N_VGND_c_1237_n 0.0121945f $X=9.23 $Y=0.59 $X2=0
+ $Y2=0
cc_650 N_A_1617_76#_M1025_g N_VGND_c_1237_n 0.00180376f $X=9.59 $Y=0.59 $X2=0
+ $Y2=0
cc_651 N_A_1617_76#_c_1019_n N_VGND_c_1237_n 0.024419f $X=9.155 $Y=1.085 $X2=0
+ $Y2=0
cc_652 N_A_1617_76#_c_1020_n N_VGND_c_1237_n 0.0158869f $X=8.225 $Y=0.59 $X2=0
+ $Y2=0
cc_653 N_A_1617_76#_c_1022_n N_VGND_c_1237_n 0.00193744f $X=9.32 $Y=1.165 $X2=0
+ $Y2=0
cc_654 N_A_1617_76#_c_1020_n N_VGND_c_1241_n 0.0143928f $X=8.225 $Y=0.59 $X2=0
+ $Y2=0
cc_655 N_A_1617_76#_M1023_g N_VGND_c_1242_n 0.0047441f $X=9.23 $Y=0.59 $X2=0
+ $Y2=0
cc_656 N_A_1617_76#_M1025_g N_VGND_c_1242_n 0.00544382f $X=9.59 $Y=0.59 $X2=0
+ $Y2=0
cc_657 N_A_1617_76#_M1023_g N_VGND_c_1243_n 0.00455844f $X=9.23 $Y=0.59 $X2=0
+ $Y2=0
cc_658 N_A_1617_76#_M1025_g N_VGND_c_1243_n 0.00542671f $X=9.59 $Y=0.59 $X2=0
+ $Y2=0
cc_659 N_A_1617_76#_c_1020_n N_VGND_c_1243_n 0.0124752f $X=8.225 $Y=0.59 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_1079_n A_698_419# 0.010279f $X=9.84 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_661 N_VPWR_c_1079_n A_904_419# 0.010279f $X=9.84 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_662 N_VPWR_c_1079_n N_Q_M1001_d 0.0023218f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_663 N_VPWR_c_1083_n Q 0.0712868f $X=7.36 $Y=2.24 $X2=0 $Y2=0
cc_664 N_VPWR_c_1088_n Q 0.0210372f $X=8.85 $Y=3.33 $X2=0 $Y2=0
cc_665 N_VPWR_c_1079_n Q 0.0131898f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_666 N_VPWR_c_1089_n Q_N 0.0191637f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_667 N_VPWR_c_1079_n Q_N 0.0204781f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_668 N_VPWR_c_1084_n N_Q_N_c_1212_n 0.071673f $X=9.015 $Y=2.015 $X2=0 $Y2=0
cc_669 N_Q_c_1181_n N_VGND_c_1236_n 0.0111268f $X=7.675 $Y=0.975 $X2=0 $Y2=0
cc_670 N_Q_c_1181_n N_VGND_c_1241_n 0.00579094f $X=7.675 $Y=0.975 $X2=0 $Y2=0
cc_671 N_Q_c_1181_n N_VGND_c_1243_n 0.0100214f $X=7.675 $Y=0.975 $X2=0 $Y2=0
cc_672 N_Q_N_c_1209_n N_VGND_c_1237_n 0.0153904f $X=9.805 $Y=0.59 $X2=0 $Y2=0
cc_673 N_Q_N_c_1209_n N_VGND_c_1242_n 0.013815f $X=9.805 $Y=0.59 $X2=0 $Y2=0
cc_674 N_Q_N_c_1209_n N_VGND_c_1243_n 0.0119446f $X=9.805 $Y=0.59 $X2=0 $Y2=0
cc_675 N_VGND_c_1243_n A_542_47# 0.00312872f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_676 N_VGND_c_1243_n A_758_47# 0.00357568f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_677 N_VGND_c_1243_n A_950_47# 0.00437871f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
