* File: sky130_fd_sc_lp__o311a_1.pex.spice
* Created: Fri Aug 28 11:13:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311A_1%A_80_21# 1 2 3 12 16 20 23 24 27 31 34 35 37
+ 41 43 52
r91 43 45 20.1147 $w=5.43e-07 $l=6.35e-07 $layer=LI1_cond $X=3.347 $Y=0.38
+ $X2=3.347 $Y2=1.015
r92 37 39 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.515 $Y=1.98
+ $X2=3.515 $Y2=2.91
r93 35 46 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.515 $Y=1.79
+ $X2=3.16 $Y2=1.79
r94 35 37 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.515 $Y=1.875
+ $X2=3.515 $Y2=1.98
r95 34 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=1.705
+ $X2=3.16 $Y2=1.79
r96 34 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.16 $Y=1.705
+ $X2=3.16 $Y2=1.015
r97 32 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=1.79
+ $X2=2.425 $Y2=1.79
r98 31 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=1.79
+ $X2=3.16 $Y2=1.79
r99 31 32 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.075 $Y=1.79
+ $X2=2.59 $Y2=1.79
r100 27 29 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=2.425 $Y=1.98
+ $X2=2.425 $Y2=2.91
r101 25 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=1.875
+ $X2=2.425 $Y2=1.79
r102 25 27 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.425 $Y=1.875
+ $X2=2.425 $Y2=1.98
r103 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=1.79
+ $X2=2.425 $Y2=1.79
r104 23 24 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=2.26 $Y=1.79
+ $X2=0.795 $Y2=1.79
r105 21 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.63 $Y=1.51 $X2=0.72
+ $Y2=1.51
r106 21 49 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.63 $Y=1.51
+ $X2=0.475 $Y2=1.51
r107 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.51 $X2=0.63 $Y2=1.51
r108 18 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.665 $Y=1.705
+ $X2=0.795 $Y2=1.79
r109 18 20 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=0.665 $Y=1.705
+ $X2=0.665 $Y2=1.51
r110 14 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.675
+ $X2=0.72 $Y2=1.51
r111 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.72 $Y=1.675
+ $X2=0.72 $Y2=2.465
r112 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=1.51
r113 10 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=0.655
r114 3 39 400 $w=1.7e-07 $l=1.15688e-06 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.835 $X2=3.485 $Y2=2.91
r115 3 37 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.835 $X2=3.485 $Y2=1.98
r116 2 29 400 $w=1.7e-07 $l=1.16614e-06 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.835 $X2=2.425 $Y2=2.91
r117 2 27 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.835 $X2=2.425 $Y2=1.98
r118 1 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.315
+ $Y=0.235 $X2=3.455 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%A1 3 6 8 9 10 15 17
r40 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.35
+ $X2=1.17 $Y2=1.515
r41 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.35
+ $X2=1.17 $Y2=1.185
r42 10 26 5.51891 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=1.215 $Y=1.295
+ $X2=1.215 $Y2=1.185
r43 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.35 $X2=1.17 $Y2=1.35
r44 9 26 14.4182 $w=1.98e-07 $l=2.6e-07 $layer=LI1_cond $X=1.185 $Y=0.925
+ $X2=1.185 $Y2=1.185
r45 8 9 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.185 $Y=0.555
+ $X2=1.185 $Y2=0.925
r46 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.26 $Y=2.465
+ $X2=1.26 $Y2=1.515
r47 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.26 $Y=0.655
+ $X2=1.26 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%A2 3 7 8 11 13
r30 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.35
+ $X2=1.71 $Y2=1.515
r31 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.35
+ $X2=1.71 $Y2=1.185
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.35 $X2=1.71 $Y2=1.35
r33 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.755 $Y=0.655
+ $X2=1.755 $Y2=1.185
r34 3 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.705 $Y=2.465
+ $X2=1.705 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%A3 3 7 8 11 12 13
r30 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.35
+ $X2=2.25 $Y2=1.515
r31 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.35
+ $X2=2.25 $Y2=1.185
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.35 $X2=2.25 $Y2=1.35
r33 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.35 $X2=2.25
+ $Y2=1.35
r34 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.34 $Y=0.655
+ $X2=2.34 $Y2=1.185
r35 3 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.16 $Y=2.465
+ $X2=2.16 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%B1 3 7 8 11 12 13
r30 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.35
+ $X2=2.79 $Y2=1.515
r31 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.35
+ $X2=2.79 $Y2=1.185
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.35 $X2=2.79 $Y2=1.35
r33 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=1.35 $X2=2.79
+ $Y2=1.35
r34 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.88 $Y=0.655
+ $X2=2.88 $Y2=1.185
r35 3 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.7 $Y=2.465 $X2=2.7
+ $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%C1 1 3 6 8 13
r25 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.51
+ $Y=1.36 $X2=3.51 $Y2=1.36
r26 10 13 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.24 $Y=1.36
+ $X2=3.51 $Y2=1.36
r27 8 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.6 $Y=1.36 $X2=3.51
+ $Y2=1.36
r28 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.525
+ $X2=3.24 $Y2=1.36
r29 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.24 $Y=1.525 $X2=3.24
+ $Y2=2.465
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.195
+ $X2=3.24 $Y2=1.36
r31 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.24 $Y=1.195 $X2=3.24
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%X 1 2 7 8 9 10 11 12 13 25 37 40
r20 38 40 1.5185 $w=5.73e-07 $l=7.3e-08 $layer=LI1_cond $X=0.382 $Y=2.332
+ $X2=0.382 $Y2=2.405
r21 37 48 0.426831 $w=2.68e-07 $l=1e-08 $layer=LI1_cond $X=0.23 $Y=2.035
+ $X2=0.23 $Y2=2.045
r22 13 45 3.64024 $w=5.73e-07 $l=1.75e-07 $layer=LI1_cond $X=0.382 $Y=2.775
+ $X2=0.382 $Y2=2.95
r23 12 38 0.124808 $w=5.73e-07 $l=6e-09 $layer=LI1_cond $X=0.382 $Y=2.326
+ $X2=0.382 $Y2=2.332
r24 12 50 4.07707 $w=5.73e-07 $l=1.96e-07 $layer=LI1_cond $X=0.382 $Y=2.326
+ $X2=0.382 $Y2=2.13
r25 12 13 7.5717 $w=5.73e-07 $l=3.64e-07 $layer=LI1_cond $X=0.382 $Y=2.411
+ $X2=0.382 $Y2=2.775
r26 12 40 0.124808 $w=5.73e-07 $l=6e-09 $layer=LI1_cond $X=0.382 $Y=2.411
+ $X2=0.382 $Y2=2.405
r27 11 50 0.998465 $w=5.73e-07 $l=4.8e-08 $layer=LI1_cond $X=0.382 $Y=2.082
+ $X2=0.382 $Y2=2.13
r28 11 48 4.15721 $w=5.73e-07 $l=3.7e-08 $layer=LI1_cond $X=0.382 $Y=2.082
+ $X2=0.382 $Y2=2.045
r29 11 37 1.62196 $w=2.68e-07 $l=3.8e-08 $layer=LI1_cond $X=0.23 $Y=1.997
+ $X2=0.23 $Y2=2.035
r30 10 11 14.1708 $w=2.68e-07 $l=3.32e-07 $layer=LI1_cond $X=0.23 $Y=1.665
+ $X2=0.23 $Y2=1.997
r31 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.665
r32 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.925 $X2=0.23
+ $Y2=1.295
r33 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.555 $X2=0.23
+ $Y2=0.925
r34 7 25 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.23 $Y=0.555
+ $X2=0.23 $Y2=0.42
r35 2 50 400 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=1.835 $X2=0.505 $Y2=2.13
r36 2 45 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=1.835 $X2=0.505 $Y2=2.95
r37 1 25 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%VPWR 1 2 9 15 20 21 23 24 25 38 39
r41 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 29 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 25 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 25 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 23 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=3.33 $X2=2.64
+ $Y2=3.33
r51 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=3.33
+ $X2=2.965 $Y2=3.33
r52 22 38 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.13 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=3.33
+ $X2=2.965 $Y2=3.33
r54 20 28 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=1.005 $Y2=3.33
r56 19 32 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.17 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=3.33
+ $X2=1.005 $Y2=3.33
r58 15 18 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=2.965 $Y=2.13
+ $X2=2.965 $Y2=2.95
r59 13 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=3.245
+ $X2=2.965 $Y2=3.33
r60 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.965 $Y=3.245
+ $X2=2.965 $Y2=2.95
r61 9 12 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.005 $Y=2.13
+ $X2=1.005 $Y2=2.95
r62 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.005 $Y=3.245
+ $X2=1.005 $Y2=3.33
r63 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.005 $Y=3.245
+ $X2=1.005 $Y2=2.95
r64 2 18 400 $w=1.7e-07 $l=1.20626e-06 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.965 $Y2=2.95
r65 2 15 400 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.965 $Y2=2.13
r66 1 12 400 $w=1.7e-07 $l=1.21547e-06 $layer=licon1_PDIFF $count=1 $X=0.795
+ $Y=1.835 $X2=1.005 $Y2=2.95
r67 1 9 400 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_PDIFF $count=1 $X=0.795
+ $Y=1.835 $X2=1.005 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r49 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r50 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 30 37 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r52 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r53 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.05
+ $Y2=0
r54 27 29 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=2.215 $Y=0 $X2=3.6
+ $Y2=0
r55 26 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r56 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r58 23 25 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.68
+ $Y2=0
r59 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.05
+ $Y2=0
r60 22 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=1.68
+ $Y2=0
r61 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r64 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r65 15 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r66 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r67 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0
r68 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0.55
r69 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r70 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.38
r71 2 13 182 $w=1.7e-07 $l=4.10518e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.235 $X2=2.05 $Y2=0.55
r72 1 9 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_1%A_267_47# 1 2 9 11 12 13 15
r23 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0.845
+ $X2=2.615 $Y2=0.93
r24 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.615 $Y=0.845
+ $X2=2.615 $Y2=0.38
r25 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0.93
+ $X2=2.615 $Y2=0.93
r26 11 12 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.45 $Y=0.93
+ $X2=1.675 $Y2=0.93
r27 7 12 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.565 $Y=0.845
+ $X2=1.675 $Y2=0.93
r28 7 9 22.2631 $w=2.18e-07 $l=4.25e-07 $layer=LI1_cond $X=1.565 $Y=0.845
+ $X2=1.565 $Y2=0.42
r29 2 18 182 $w=1.7e-07 $l=7.88686e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.615 $Y2=0.93
r30 2 15 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.615 $Y2=0.38
r31 1 9 91 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=2 $X=1.335
+ $Y=0.235 $X2=1.54 $Y2=0.42
.ends

