* File: sky130_fd_sc_lp__o41a_m.pex.spice
* Created: Wed Sep  2 10:27:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41A_M%A_80_21# 1 2 9 11 14 16 20 21 22 23 24 25 28
+ 32 35
c74 22 0 5.36468e-20 $X=1.105 $Y=0.81
c75 21 0 1.12474e-19 $X=0.63 $Y=0.93
r76 30 32 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=1.32 $Y=2.615
+ $X2=1.32 $Y2=2.82
r77 26 28 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=1.21 $Y=0.725
+ $X2=1.21 $Y2=0.53
r78 24 30 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.225 $Y=2.53
+ $X2=1.32 $Y2=2.615
r79 24 25 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.225 $Y=2.53
+ $X2=0.715 $Y2=2.53
r80 22 26 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.105 $Y=0.81
+ $X2=1.21 $Y2=0.725
r81 22 23 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.105 $Y=0.81
+ $X2=0.715 $Y2=0.81
r82 21 35 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=0.93
+ $X2=0.597 $Y2=0.765
r83 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=0.93 $X2=0.63 $Y2=0.93
r84 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=2.445
+ $X2=0.715 $Y2=2.53
r85 18 20 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=0.63 $Y=2.445
+ $X2=0.63 $Y2=0.93
r86 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=0.895
+ $X2=0.715 $Y2=0.81
r87 17 20 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.63 $Y=0.895
+ $X2=0.63 $Y2=0.93
r88 14 16 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=0.67 $Y=2.885
+ $X2=0.67 $Y2=1.435
r89 11 16 43.6889 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.597 $Y=1.238
+ $X2=0.597 $Y2=1.435
r90 10 21 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.597 $Y=0.962
+ $X2=0.597 $Y2=0.93
r91 10 11 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.597 $Y=0.962
+ $X2=0.597 $Y2=1.238
r92 9 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.765
r93 2 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.19
+ $Y=2.675 $X2=1.33 $Y2=2.82
r94 1 28 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.255 $X2=1.21 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%B1 3 9 12 13 14 17 19 20 21 26
c53 19 0 1.38473e-19 $X=1.2 $Y=1.295
r54 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.12
+ $Y=1.84 $X2=1.12 $Y2=1.84
r55 21 27 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.12 $Y=2.035
+ $X2=1.12 $Y2=1.84
r56 20 27 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.84
r57 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=1.295
+ $X2=1.12 $Y2=1.665
r58 15 17 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.21 $Y=0.895
+ $X2=1.425 $Y2=0.895
r59 13 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.12 $Y=2.18
+ $X2=1.12 $Y2=1.84
r60 13 14 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=2.18
+ $X2=1.12 $Y2=2.345
r61 12 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.675
+ $X2=1.12 $Y2=1.84
r62 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=0.82
+ $X2=1.425 $Y2=0.895
r63 7 9 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=1.425 $Y=0.82
+ $X2=1.425 $Y2=0.465
r64 5 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.21 $Y=0.97 $X2=1.21
+ $Y2=0.895
r65 5 12 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.21 $Y=0.97 $X2=1.21
+ $Y2=1.675
r66 3 14 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.115 $Y=2.885
+ $X2=1.115 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%A4 2 5 11 12 13 14 15 16 17 18 19 26 28
c55 14 0 8.00614e-20 $X=1.82 $Y=0.935
r56 26 28 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.677 $Y=1.375
+ $X2=1.677 $Y2=1.21
r57 18 19 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.405
+ $X2=1.68 $Y2=2.775
r58 17 18 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.405
r59 16 17 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=2.035
r60 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.665
r61 15 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.375 $X2=1.68 $Y2=1.375
r62 14 28 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.785 $Y=0.935
+ $X2=1.785 $Y2=1.21
r63 13 14 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.82 $Y=0.785
+ $X2=1.82 $Y2=0.935
r64 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.855 $Y=0.465
+ $X2=1.855 $Y2=0.785
r65 5 12 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.57 $Y=2.885
+ $X2=1.57 $Y2=1.88
r66 2 12 49.3547 $w=3.65e-07 $l=1.82e-07 $layer=POLY_cond $X=1.677 $Y=1.698
+ $X2=1.677 $Y2=1.88
r67 1 26 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=1.677 $Y=1.392
+ $X2=1.677 $Y2=1.375
r68 1 2 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=1.677 $Y=1.392
+ $X2=1.677 $Y2=1.698
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%A3 3 7 11 12 13 14 15 16 22
r43 15 16 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.197 $Y=2.035
+ $X2=2.197 $Y2=2.405
r44 14 15 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.197 $Y=1.665
+ $X2=2.197 $Y2=2.035
r45 13 14 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.197 $Y=1.295
+ $X2=2.197 $Y2=1.665
r46 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.235
+ $Y=1.31 $X2=2.235 $Y2=1.31
r47 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.235 $Y=1.65
+ $X2=2.235 $Y2=1.31
r48 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.65
+ $X2=2.235 $Y2=1.815
r49 10 22 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.145
+ $X2=2.235 $Y2=1.31
r50 7 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.285 $Y=0.465
+ $X2=2.285 $Y2=1.145
r51 3 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.145 $Y=2.885
+ $X2=2.145 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%A2 3 7 9 11 14 15 16 17 23
c47 9 0 1.08688e-19 $X=2.505 $Y=2.13
r48 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.805
+ $Y=1.67 $X2=2.805 $Y2=1.67
r49 16 17 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.722 $Y=2.035
+ $X2=2.722 $Y2=2.405
r50 16 24 12.5565 $w=3.33e-07 $l=3.65e-07 $layer=LI1_cond $X=2.722 $Y=2.035
+ $X2=2.722 $Y2=1.67
r51 15 24 0.172006 $w=3.33e-07 $l=5e-09 $layer=LI1_cond $X=2.722 $Y=1.665
+ $X2=2.722 $Y2=1.67
r52 14 15 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.722 $Y=1.295
+ $X2=2.722 $Y2=1.665
r53 13 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.505
+ $X2=2.805 $Y2=1.67
r54 11 23 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=2.805 $Y=2.055
+ $X2=2.805 $Y2=1.67
r55 9 11 103.286 $w=1.4e-07 $l=3e-07 $layer=POLY_cond $X=2.505 $Y=2.13 $X2=2.805
+ $Y2=2.13
r56 7 13 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.715 $Y=0.465
+ $X2=2.715 $Y2=1.505
r57 1 9 1.15097 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=2.205
+ $X2=2.505 $Y2=2.13
r58 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.505 $Y=2.205
+ $X2=2.505 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%A1 1 3 4 5 8 14 17 18 19 20 21 22 28
c40 19 0 2.87744e-20 $X=3.6 $Y=1.295
r41 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.455
+ $Y=1.835 $X2=3.455 $Y2=1.835
r42 21 22 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.527 $Y=2.035
+ $X2=3.527 $Y2=2.405
r43 21 29 7.3171 $w=3.13e-07 $l=2e-07 $layer=LI1_cond $X=3.527 $Y=2.035
+ $X2=3.527 $Y2=1.835
r44 20 29 6.21953 $w=3.13e-07 $l=1.7e-07 $layer=LI1_cond $X=3.527 $Y=1.665
+ $X2=3.527 $Y2=1.835
r45 19 20 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.527 $Y=1.295
+ $X2=3.527 $Y2=1.665
r46 18 28 101.42 $w=3.3e-07 $l=5.8e-07 $layer=POLY_cond $X=3.455 $Y=2.415
+ $X2=3.455 $Y2=1.835
r47 17 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.455 $Y=1.67
+ $X2=3.455 $Y2=1.835
r48 12 14 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.145 $Y=1.19
+ $X2=3.365 $Y2=1.19
r49 10 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=1.265
+ $X2=3.365 $Y2=1.19
r50 10 17 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.365 $Y=1.265
+ $X2=3.365 $Y2=1.67
r51 6 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.145 $Y=1.115
+ $X2=3.145 $Y2=1.19
r52 6 8 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.145 $Y=1.115
+ $X2=3.145 $Y2=0.465
r53 4 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.29 $Y=2.49
+ $X2=3.455 $Y2=2.415
r54 4 5 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.29 $Y=2.49 $X2=2.94
+ $Y2=2.49
r55 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.865 $Y=2.565
+ $X2=2.94 $Y2=2.49
r56 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.865 $Y=2.565
+ $X2=2.865 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%X 1 2 7 8 9 10 11 20 32 37
r16 35 37 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=0.26 $Y=2.9
+ $X2=0.455 $Y2=2.9
r17 18 35 0.716491 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=0.26 $Y=2.795
+ $X2=0.26 $Y2=2.9
r18 18 32 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=0.26 $Y=2.795 $X2=0.26
+ $Y2=2.775
r19 11 35 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=2.9 $X2=0.26
+ $Y2=2.9
r20 11 32 1.74286 $w=2.08e-07 $l=3.3e-08 $layer=LI1_cond $X=0.26 $Y=2.742
+ $X2=0.26 $Y2=2.775
r21 10 11 17.7983 $w=2.08e-07 $l=3.37e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.742
r22 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.035
+ $X2=0.26 $Y2=2.405
r23 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665 $X2=0.26
+ $Y2=2.035
r24 7 8 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295 $X2=0.26
+ $Y2=1.665
r25 7 20 41.4589 $w=2.08e-07 $l=7.85e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=0.51
r26 2 37 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=2.675 $X2=0.455 $Y2=2.9
r27 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%VPWR 1 2 9 13 16 17 18 24 33 34 37
c48 13 0 7.99132e-20 $X=3.08 $Y=2.95
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 34 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 31 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.08 $Y2=3.33
r53 31 33 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.08 $Y2=3.33
r59 24 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 18 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 16 21 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.8 $Y=3.33 $X2=0.72
+ $Y2=3.33
r65 16 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=3.33 $X2=0.895
+ $Y2=3.33
r66 15 26 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.2
+ $Y2=3.33
r67 15 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.895 $Y2=3.33
r68 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=3.33
r69 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.95
r70 7 17 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=3.33
r71 7 9 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=2.97
r72 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=2.675 $X2=3.08 $Y2=2.95
r73 1 9 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=0.745
+ $Y=2.675 $X2=0.885 $Y2=2.97
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%VGND 1 2 3 12 16 20 23 24 26 27 28 30 43 44
+ 47
c57 44 0 2.64147e-20 $X=3.6 $Y=0
c58 30 0 1.12474e-19 $X=0.585 $Y=0
r59 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r60 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r62 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 38 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r64 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r65 35 47 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.69
+ $Y2=0
r66 35 37 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.68
+ $Y2=0
r67 33 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r68 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r69 30 47 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.69
+ $Y2=0
r70 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r71 28 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r72 28 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r73 26 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.64
+ $Y2=0
r74 26 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.93
+ $Y2=0
r75 25 43 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=3.6
+ $Y2=0
r76 25 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=2.93
+ $Y2=0
r77 23 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=1.68
+ $Y2=0
r78 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=2.07
+ $Y2=0
r79 22 40 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.64
+ $Y2=0
r80 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.07
+ $Y2=0
r81 18 27 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=0.085
+ $X2=2.93 $Y2=0
r82 18 20 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=2.93 $Y=0.085
+ $X2=2.93 $Y2=0.4
r83 14 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0
r84 14 16 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0.4
r85 10 47 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r86 10 12 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r87 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.255 $X2=2.93 $Y2=0.4
r88 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.255 $X2=2.07 $Y2=0.4
r89 1 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_M%A_300_51# 1 2 3 12 14 15 18 20 24 26
r47 22 24 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=3.36 $Y=0.745
+ $X2=3.36 $Y2=0.53
r48 21 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.605 $Y=0.83
+ $X2=2.5 $Y2=0.83
r49 20 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.255 $Y=0.83
+ $X2=3.36 $Y2=0.745
r50 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.255 $Y=0.83
+ $X2=2.605 $Y2=0.83
r51 16 26 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=0.745 $X2=2.5
+ $Y2=0.83
r52 16 18 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.5 $Y=0.745 $X2=2.5
+ $Y2=0.53
r53 14 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.395 $Y=0.83
+ $X2=2.5 $Y2=0.83
r54 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.395 $Y=0.83
+ $X2=1.745 $Y2=0.83
r55 10 15 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.64 $Y=0.745
+ $X2=1.745 $Y2=0.83
r56 10 12 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.64 $Y=0.745
+ $X2=1.64 $Y2=0.53
r57 3 24 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.255 $X2=3.36 $Y2=0.53
r58 2 18 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.255 $X2=2.5 $Y2=0.53
r59 1 12 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.255 $X2=1.64 $Y2=0.53
.ends

