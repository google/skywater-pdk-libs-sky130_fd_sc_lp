* File: sky130_fd_sc_lp__dfrbp_2.pxi.spice
* Created: Wed Sep  2 09:43:21 2020
* 
x_PM_SKY130_FD_SC_LP__DFRBP_2%CLK N_CLK_M1033_g N_CLK_c_246_n N_CLK_M1005_g CLK
+ CLK PM_SKY130_FD_SC_LP__DFRBP_2%CLK
x_PM_SKY130_FD_SC_LP__DFRBP_2%D N_D_M1027_g N_D_M1008_g N_D_c_280_n N_D_c_281_n
+ N_D_c_286_n D D N_D_c_283_n PM_SKY130_FD_SC_LP__DFRBP_2%D
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_196_79# N_A_196_79#_M1006_d N_A_196_79#_M1020_d
+ N_A_196_79#_M1019_g N_A_196_79#_c_331_n N_A_196_79#_M1002_g
+ N_A_196_79#_c_332_n N_A_196_79#_M1013_g N_A_196_79#_c_333_n
+ N_A_196_79#_M1031_g N_A_196_79#_c_350_n N_A_196_79#_c_351_n
+ N_A_196_79#_c_334_n N_A_196_79#_c_335_n N_A_196_79#_c_336_n
+ N_A_196_79#_c_337_n N_A_196_79#_c_338_n N_A_196_79#_c_339_n
+ N_A_196_79#_c_340_n N_A_196_79#_c_341_n N_A_196_79#_c_354_n
+ N_A_196_79#_c_342_n N_A_196_79#_c_343_n N_A_196_79#_c_344_n
+ N_A_196_79#_c_345_n N_A_196_79#_c_346_n PM_SKY130_FD_SC_LP__DFRBP_2%A_196_79#
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_811_341# N_A_811_341#_M1007_d
+ N_A_811_341#_M1025_d N_A_811_341#_M1034_g N_A_811_341#_c_519_n
+ N_A_811_341#_M1000_g N_A_811_341#_c_520_n N_A_811_341#_c_521_n
+ N_A_811_341#_c_522_n N_A_811_341#_c_523_n N_A_811_341#_c_530_n
+ N_A_811_341#_c_531_n N_A_811_341#_c_524_n N_A_811_341#_c_533_n
+ N_A_811_341#_c_525_n N_A_811_341#_c_561_p
+ PM_SKY130_FD_SC_LP__DFRBP_2%A_811_341#
x_PM_SKY130_FD_SC_LP__DFRBP_2%RESET_B N_RESET_B_M1016_g N_RESET_B_M1001_g
+ N_RESET_B_c_631_n N_RESET_B_c_632_n N_RESET_B_M1032_g N_RESET_B_M1012_g
+ N_RESET_B_M1003_g N_RESET_B_M1011_g N_RESET_B_c_635_n N_RESET_B_c_644_n
+ N_RESET_B_c_636_n N_RESET_B_c_645_n N_RESET_B_c_646_n N_RESET_B_c_647_n
+ N_RESET_B_c_648_n N_RESET_B_c_649_n RESET_B N_RESET_B_c_637_n
+ N_RESET_B_c_638_n N_RESET_B_c_653_n N_RESET_B_c_639_n N_RESET_B_c_655_n
+ N_RESET_B_c_656_n PM_SKY130_FD_SC_LP__DFRBP_2%RESET_B
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_637_191# N_A_637_191#_M1028_d
+ N_A_637_191#_M1019_d N_A_637_191#_M1012_d N_A_637_191#_c_824_n
+ N_A_637_191#_M1007_g N_A_637_191#_M1025_g N_A_637_191#_c_825_n
+ N_A_637_191#_c_830_n N_A_637_191#_c_831_n N_A_637_191#_c_846_n
+ N_A_637_191#_c_848_n N_A_637_191#_c_826_n N_A_637_191#_c_827_n
+ PM_SKY130_FD_SC_LP__DFRBP_2%A_637_191#
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_27_79# N_A_27_79#_M1033_s N_A_27_79#_M1005_s
+ N_A_27_79#_M1006_g N_A_27_79#_M1020_g N_A_27_79#_c_929_n N_A_27_79#_c_930_n
+ N_A_27_79#_c_941_n N_A_27_79#_c_942_n N_A_27_79#_c_931_n N_A_27_79#_c_944_n
+ N_A_27_79#_c_932_n N_A_27_79#_c_933_n N_A_27_79#_M1028_g N_A_27_79#_c_946_n
+ N_A_27_79#_M1035_g N_A_27_79#_c_948_n N_A_27_79#_M1024_g N_A_27_79#_M1015_g
+ N_A_27_79#_c_950_n N_A_27_79#_c_951_n N_A_27_79#_c_952_n N_A_27_79#_c_953_n
+ N_A_27_79#_c_935_n N_A_27_79#_c_954_n N_A_27_79#_c_955_n N_A_27_79#_c_936_n
+ N_A_27_79#_c_937_n N_A_27_79#_c_938_n N_A_27_79#_c_939_n
+ PM_SKY130_FD_SC_LP__DFRBP_2%A_27_79#
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_1444_320# N_A_1444_320#_M1029_d
+ N_A_1444_320#_M1011_d N_A_1444_320#_M1036_g N_A_1444_320#_M1037_g
+ N_A_1444_320#_c_1097_n N_A_1444_320#_c_1098_n N_A_1444_320#_c_1099_n
+ N_A_1444_320#_c_1100_n N_A_1444_320#_c_1093_n N_A_1444_320#_c_1101_n
+ N_A_1444_320#_c_1094_n N_A_1444_320#_c_1103_n N_A_1444_320#_c_1104_n
+ N_A_1444_320#_c_1105_n PM_SKY130_FD_SC_LP__DFRBP_2%A_1444_320#
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_1272_128# N_A_1272_128#_M1013_d
+ N_A_1272_128#_M1024_d N_A_1272_128#_c_1182_n N_A_1272_128#_M1029_g
+ N_A_1272_128#_M1017_g N_A_1272_128#_c_1183_n N_A_1272_128#_c_1184_n
+ N_A_1272_128#_M1009_g N_A_1272_128#_M1010_g N_A_1272_128#_c_1186_n
+ N_A_1272_128#_M1023_g N_A_1272_128#_M1022_g N_A_1272_128#_c_1188_n
+ N_A_1272_128#_c_1189_n N_A_1272_128#_M1014_g N_A_1272_128#_M1004_g
+ N_A_1272_128#_c_1192_n N_A_1272_128#_c_1193_n N_A_1272_128#_c_1194_n
+ N_A_1272_128#_c_1195_n N_A_1272_128#_c_1210_n N_A_1272_128#_c_1211_n
+ N_A_1272_128#_c_1196_n N_A_1272_128#_c_1197_n N_A_1272_128#_c_1198_n
+ N_A_1272_128#_c_1199_n PM_SKY130_FD_SC_LP__DFRBP_2%A_1272_128#
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_2028_367# N_A_2028_367#_M1004_s
+ N_A_2028_367#_M1014_s N_A_2028_367#_M1021_g N_A_2028_367#_M1018_g
+ N_A_2028_367#_c_1347_n N_A_2028_367#_M1030_g N_A_2028_367#_M1026_g
+ N_A_2028_367#_c_1350_n N_A_2028_367#_c_1351_n N_A_2028_367#_c_1352_n
+ N_A_2028_367#_c_1353_n N_A_2028_367#_c_1354_n N_A_2028_367#_c_1355_n
+ N_A_2028_367#_c_1356_n PM_SKY130_FD_SC_LP__DFRBP_2%A_2028_367#
x_PM_SKY130_FD_SC_LP__DFRBP_2%VPWR N_VPWR_M1005_d N_VPWR_M1016_d N_VPWR_M1000_d
+ N_VPWR_M1025_s N_VPWR_M1036_d N_VPWR_M1017_d N_VPWR_M1023_d N_VPWR_M1014_d
+ N_VPWR_M1026_d N_VPWR_c_1414_n N_VPWR_c_1415_n N_VPWR_c_1416_n N_VPWR_c_1417_n
+ N_VPWR_c_1418_n N_VPWR_c_1419_n N_VPWR_c_1420_n N_VPWR_c_1421_n
+ N_VPWR_c_1422_n N_VPWR_c_1423_n N_VPWR_c_1424_n N_VPWR_c_1425_n VPWR
+ N_VPWR_c_1426_n N_VPWR_c_1427_n N_VPWR_c_1428_n N_VPWR_c_1429_n
+ N_VPWR_c_1430_n N_VPWR_c_1431_n N_VPWR_c_1432_n N_VPWR_c_1433_n
+ N_VPWR_c_1434_n N_VPWR_c_1435_n N_VPWR_c_1436_n N_VPWR_c_1437_n
+ N_VPWR_c_1438_n N_VPWR_c_1439_n N_VPWR_c_1440_n N_VPWR_c_1413_n
+ PM_SKY130_FD_SC_LP__DFRBP_2%VPWR
x_PM_SKY130_FD_SC_LP__DFRBP_2%A_308_463# N_A_308_463#_M1027_d
+ N_A_308_463#_M1016_s N_A_308_463#_M1008_d N_A_308_463#_M1019_s
+ N_A_308_463#_c_1573_n N_A_308_463#_c_1568_n N_A_308_463#_c_1570_n
+ N_A_308_463#_c_1571_n PM_SKY130_FD_SC_LP__DFRBP_2%A_308_463#
x_PM_SKY130_FD_SC_LP__DFRBP_2%Q_N N_Q_N_M1010_d N_Q_N_M1009_s Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1638_p Q_N PM_SKY130_FD_SC_LP__DFRBP_2%Q_N
x_PM_SKY130_FD_SC_LP__DFRBP_2%Q N_Q_M1021_d N_Q_M1018_s Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DFRBP_2%Q
x_PM_SKY130_FD_SC_LP__DFRBP_2%VGND N_VGND_M1033_d N_VGND_M1001_s N_VGND_M1032_d
+ N_VGND_M1037_d N_VGND_M1010_s N_VGND_M1022_s N_VGND_M1004_d N_VGND_M1030_s
+ N_VGND_c_1658_n N_VGND_c_1659_n N_VGND_c_1660_n N_VGND_c_1661_n
+ N_VGND_c_1662_n N_VGND_c_1663_n N_VGND_c_1664_n N_VGND_c_1665_n
+ N_VGND_c_1666_n N_VGND_c_1667_n N_VGND_c_1668_n VGND N_VGND_c_1669_n
+ N_VGND_c_1670_n N_VGND_c_1671_n N_VGND_c_1672_n N_VGND_c_1673_n
+ N_VGND_c_1674_n N_VGND_c_1675_n N_VGND_c_1676_n N_VGND_c_1677_n
+ N_VGND_c_1678_n N_VGND_c_1679_n N_VGND_c_1680_n N_VGND_c_1681_n
+ N_VGND_c_1682_n PM_SKY130_FD_SC_LP__DFRBP_2%VGND
cc_1 VNB N_CLK_M1033_g 0.0449989f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.605
cc_2 VNB N_CLK_c_246_n 0.026977f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.97
cc_3 VNB CLK 0.00427655f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_D_c_280_n 0.0153758f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_D_c_281_n 0.00470711f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_6 VNB D 0.00123743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_D_c_283_n 0.0165182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_196_79#_c_331_n 0.0146213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_196_79#_c_332_n 0.0190363f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.805
cc_10 VNB N_A_196_79#_c_333_n 0.0227536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_196_79#_c_334_n 0.01263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_196_79#_c_335_n 0.0105577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_196_79#_c_336_n 0.0248022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_196_79#_c_337_n 0.00954372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_196_79#_c_338_n 0.0363288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_196_79#_c_339_n 0.0072662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_196_79#_c_340_n 0.00100954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_196_79#_c_341_n 0.0160226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_196_79#_c_342_n 0.00409486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_196_79#_c_343_n 0.00236147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_196_79#_c_344_n 0.00105935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_196_79#_c_345_n 0.038855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_196_79#_c_346_n 0.0297902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_811_341#_M1034_g 0.0221174f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_25 VNB N_A_811_341#_c_519_n 0.00911289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_811_341#_c_520_n 2.66712e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_811_341#_c_521_n 0.0154978f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.035
cc_28 VNB N_A_811_341#_c_522_n 0.00125933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_811_341#_c_523_n 0.00222243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_811_341#_c_524_n 0.00696357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_811_341#_c_525_n 0.00221877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_RESET_B_M1001_g 0.0279316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_c_631_n 0.135141f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_RESET_B_c_632_n 0.00871646f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_35 VNB N_RESET_B_M1032_g 0.0297865f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.805
cc_36 VNB N_RESET_B_M1003_g 0.0295296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_RESET_B_c_635_n 0.0285628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_RESET_B_c_636_n 0.00867826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_c_637_n 0.00610935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_c_638_n 0.00615306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_RESET_B_c_639_n 0.00913631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_637_191#_c_824_n 0.0193257f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_43 VNB N_A_637_191#_c_825_n 0.00283785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_637_191#_c_826_n 0.004564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_637_191#_c_827_n 0.0400756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_79#_M1006_g 0.0153952f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_47 VNB N_A_27_79#_c_929_n 0.436891f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.805
cc_48 VNB N_A_27_79#_c_930_n 0.0125015f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.665
cc_49 VNB N_A_27_79#_c_931_n 0.0250505f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.035
cc_50 VNB N_A_27_79#_c_932_n 0.00824733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_27_79#_c_933_n 0.0239387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_79#_M1015_g 0.0418487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_27_79#_c_935_n 0.020003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_27_79#_c_936_n 0.00453417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_79#_c_937_n 0.0399207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_27_79#_c_938_n 0.0165056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_79#_c_939_n 0.0199478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1444_320#_M1037_g 0.0332213f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.805
cc_59 VNB N_A_1444_320#_c_1093_n 0.010102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1444_320#_c_1094_n 0.00503684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1272_128#_c_1182_n 0.0190463f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.68
cc_62 VNB N_A_1272_128#_c_1183_n 0.0147703f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.805
cc_63 VNB N_A_1272_128#_c_1184_n 0.0332711f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.805
cc_64 VNB N_A_1272_128#_M1010_g 0.0258364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1272_128#_c_1186_n 0.00516739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1272_128#_M1022_g 0.0281977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1272_128#_c_1188_n 0.0382019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1272_128#_c_1189_n 0.0196586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1272_128#_M1014_g 0.00882207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1272_128#_M1004_g 0.0229598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1272_128#_c_1192_n 0.00538399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1272_128#_c_1193_n 0.00268506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1272_128#_c_1194_n 0.0161994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1272_128#_c_1195_n 0.00480528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1272_128#_c_1196_n 0.00204963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1272_128#_c_1197_n 0.0339392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1272_128#_c_1198_n 0.00261607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1272_128#_c_1199_n 0.0017303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_2028_367#_M1018_g 0.00166771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_2028_367#_c_1347_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.805
cc_81 VNB N_A_2028_367#_M1030_g 0.0350845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2028_367#_M1026_g 0.00232429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2028_367#_c_1350_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2028_367#_c_1351_n 0.0101699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2028_367#_c_1352_n 2.45317e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2028_367#_c_1353_n 0.00696185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2028_367#_c_1354_n 0.0315211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2028_367#_c_1355_n 0.00226177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2028_367#_c_1356_n 0.0176749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VPWR_c_1413_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_308_463#_c_1568_n 0.00264963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB Q_N 0.00254628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB Q 0.00817696f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.68
cc_94 VNB N_VGND_c_1658_n 0.010397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1659_n 0.0154299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1660_n 0.0199285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1661_n 0.020095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1662_n 0.0157783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1663_n 0.0151473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1664_n 0.00894546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1665_n 0.0118625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1666_n 0.0486161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1667_n 0.0544705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1668_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1669_n 0.0183946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1670_n 0.0197005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1671_n 0.0902275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1672_n 0.0311219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1673_n 0.0131373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1674_n 0.0197233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1675_n 0.0157992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1676_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1677_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1678_n 0.00436638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1679_n 0.00524804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1680_n 0.00524804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1681_n 0.00644923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1682_n 0.605539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VPB N_CLK_c_246_n 0.0295591f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.97
cc_120 VPB N_CLK_M1005_g 0.0353151f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.68
cc_121 VPB CLK 0.00659054f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_122 VPB N_D_M1008_g 0.0203453f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.68
cc_123 VPB N_D_c_281_n 0.0190045f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_124 VPB N_D_c_286_n 0.0157172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB D 0.00738864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_196_79#_M1019_g 0.0316109f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_127 VPB N_A_196_79#_c_333_n 0.00985235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_196_79#_M1031_g 0.0506738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_196_79#_c_350_n 0.00975005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_196_79#_c_351_n 0.0103072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_196_79#_c_340_n 0.00116442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_196_79#_c_341_n 0.00482124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_196_79#_c_354_n 0.00664861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_196_79#_c_344_n 0.00292906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_196_79#_c_345_n 0.0218117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_196_79#_c_346_n 0.00936221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_811_341#_c_519_n 0.0258294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_811_341#_M1000_g 0.0285501f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.805
cc_139 VPB N_A_811_341#_c_520_n 3.5247e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_811_341#_c_523_n 0.00471895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_811_341#_c_530_n 0.00458022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_811_341#_c_531_n 0.00370116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_811_341#_c_524_n 0.00529145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_811_341#_c_533_n 0.00155678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_RESET_B_M1016_g 0.0221154f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.605
cc_146 VPB N_RESET_B_M1012_g 0.0264161f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.805
cc_147 VPB N_RESET_B_M1003_g 0.0269703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_RESET_B_M1011_g 0.0253564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_RESET_B_c_644_n 0.0172544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_645_n 0.0256272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_646_n 0.00442505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_647_n 0.0287003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_648_n 0.00395121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_RESET_B_c_649_n 0.00593005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB RESET_B 0.00129998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_RESET_B_c_637_n 0.0210637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_638_n 0.00429526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_653_n 0.0378735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_c_639_n 0.0043119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_655_n 0.0417697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_c_656_n 0.00366977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_637_191#_M1025_g 0.023071f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.805
cc_163 VPB N_A_637_191#_c_825_n 0.00931749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_637_191#_c_830_n 0.00776232f $X=-0.19 $Y=1.655 $X2=0.715
+ $Y2=1.805
cc_165 VPB N_A_637_191#_c_831_n 0.0018946f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.035
cc_166 VPB N_A_637_191#_c_826_n 0.00151023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_637_191#_c_827_n 0.0104976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_27_79#_M1020_g 0.00916224f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.805
cc_169 VPB N_A_27_79#_c_941_n 0.136091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_27_79#_c_942_n 0.0107679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_27_79#_c_931_n 0.0274575f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.035
cc_172 VPB N_A_27_79#_c_944_n 0.0644572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_27_79#_c_932_n 0.0032926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_27_79#_c_946_n 0.0528886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_27_79#_M1035_g 0.0346455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_27_79#_c_948_n 0.190742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_27_79#_M1024_g 0.0230034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_27_79#_c_950_n 0.0251614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_27_79#_c_951_n 0.0155812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_27_79#_c_952_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_27_79#_c_953_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_27_79#_c_954_n 0.0061967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_27_79#_c_955_n 0.0231767f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_27_79#_c_939_n 0.0345055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1444_320#_M1036_g 0.02434f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_186 VPB N_A_1444_320#_M1037_g 0.00855851f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.805
cc_187 VPB N_A_1444_320#_c_1097_n 0.02131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1444_320#_c_1098_n 0.0163792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1444_320#_c_1099_n 0.0106559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1444_320#_c_1100_n 0.00661469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1444_320#_c_1101_n 0.0042747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_1444_320#_c_1094_n 9.85704e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_1444_320#_c_1103_n 0.00511252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_1444_320#_c_1104_n 0.0142737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1444_320#_c_1105_n 0.00188063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1272_128#_M1017_g 0.0637553f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_1272_128#_c_1183_n 0.00685636f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.805
cc_198 VPB N_A_1272_128#_c_1184_n 0.00792678f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.805
cc_199 VPB N_A_1272_128#_M1009_g 0.0174365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1272_128#_c_1186_n 0.00369644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1272_128#_M1023_g 0.018988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1272_128#_c_1188_n 0.0131365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1272_128#_M1014_g 0.026691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1272_128#_c_1192_n 9.76387e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1272_128#_c_1193_n 9.76387e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1272_128#_c_1210_n 0.00351642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1272_128#_c_1211_n 0.00694105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1272_128#_c_1198_n 0.0073371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_2028_367#_M1018_g 0.0236461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_2028_367#_M1026_g 0.0272176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_2028_367#_c_1352_n 0.0136775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1414_n 0.00375836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1415_n 0.0110762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1416_n 0.0139596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1417_n 0.0191964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1418_n 0.0139738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1419_n 0.0118281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1420_n 0.0390346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1421_n 0.0306981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1422_n 0.0118367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1423_n 0.0586484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1424_n 0.0175562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1425_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1426_n 0.0170443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1427_n 0.0294397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1428_n 0.0560743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1429_n 0.0182786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1430_n 0.0475998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1431_n 0.0193013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1432_n 0.0230073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1433_n 0.0177272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1434_n 0.0048079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1435_n 0.00463502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1436_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1437_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1438_n 0.0130537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1439_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1440_n 0.00680245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1413_n 0.11107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_308_463#_c_1568_n 0.00201962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_308_463#_c_1570_n 0.0016432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_308_463#_c_1571_n 0.0123439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB Q_N 0.00307485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB Q 0.00347098f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.68
cc_245 CLK N_A_196_79#_c_341_n 0.0222884f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_246 CLK N_A_196_79#_c_354_n 0.012378f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_247 N_CLK_M1033_g N_A_27_79#_M1006_g 0.0105017f $X=0.475 $Y=0.605 $X2=0 $Y2=0
cc_248 N_CLK_M1033_g N_A_27_79#_c_931_n 0.00221527f $X=0.475 $Y=0.605 $X2=0
+ $Y2=0
cc_249 N_CLK_c_246_n N_A_27_79#_c_931_n 0.0261731f $X=0.5 $Y=1.97 $X2=0 $Y2=0
cc_250 N_CLK_M1005_g N_A_27_79#_c_931_n 0.00316724f $X=0.5 $Y=2.68 $X2=0 $Y2=0
cc_251 CLK N_A_27_79#_c_931_n 0.00593747f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_252 N_CLK_M1005_g N_A_27_79#_c_950_n 0.0158428f $X=0.5 $Y=2.68 $X2=0 $Y2=0
cc_253 CLK N_A_27_79#_c_950_n 0.00308799f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_254 N_CLK_M1033_g N_A_27_79#_c_935_n 0.00538039f $X=0.475 $Y=0.605 $X2=0
+ $Y2=0
cc_255 N_CLK_M1005_g N_A_27_79#_c_954_n 0.00100612f $X=0.5 $Y=2.68 $X2=0 $Y2=0
cc_256 N_CLK_M1033_g N_A_27_79#_c_936_n 0.0210006f $X=0.475 $Y=0.605 $X2=0 $Y2=0
cc_257 N_CLK_c_246_n N_A_27_79#_c_936_n 0.00185523f $X=0.5 $Y=1.97 $X2=0 $Y2=0
cc_258 CLK N_A_27_79#_c_936_n 0.0253827f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_259 N_CLK_M1033_g N_A_27_79#_c_937_n 0.0185774f $X=0.475 $Y=0.605 $X2=0 $Y2=0
cc_260 N_CLK_c_246_n N_A_27_79#_c_937_n 4.20175e-19 $X=0.5 $Y=1.97 $X2=0 $Y2=0
cc_261 CLK N_A_27_79#_c_937_n 0.00272099f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_262 N_CLK_M1033_g N_A_27_79#_c_938_n 0.00649739f $X=0.475 $Y=0.605 $X2=0
+ $Y2=0
cc_263 N_CLK_M1033_g N_A_27_79#_c_939_n 0.0107719f $X=0.475 $Y=0.605 $X2=0 $Y2=0
cc_264 N_CLK_c_246_n N_A_27_79#_c_939_n 0.0218482f $X=0.5 $Y=1.97 $X2=0 $Y2=0
cc_265 CLK N_A_27_79#_c_939_n 0.0521297f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_266 N_CLK_c_246_n N_VPWR_c_1414_n 0.00113385f $X=0.5 $Y=1.97 $X2=0 $Y2=0
cc_267 N_CLK_M1005_g N_VPWR_c_1414_n 0.0137033f $X=0.5 $Y=2.68 $X2=0 $Y2=0
cc_268 CLK N_VPWR_c_1414_n 0.0303715f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_269 N_CLK_M1005_g N_VPWR_c_1426_n 0.00411131f $X=0.5 $Y=2.68 $X2=0 $Y2=0
cc_270 N_CLK_M1005_g N_VPWR_c_1413_n 0.00817336f $X=0.5 $Y=2.68 $X2=0 $Y2=0
cc_271 N_CLK_M1033_g N_VGND_c_1658_n 0.00349517f $X=0.475 $Y=0.605 $X2=0 $Y2=0
cc_272 N_CLK_M1033_g N_VGND_c_1669_n 0.00559701f $X=0.475 $Y=0.605 $X2=0 $Y2=0
cc_273 N_CLK_M1033_g N_VGND_c_1682_n 0.00537853f $X=0.475 $Y=0.605 $X2=0 $Y2=0
cc_274 D N_A_196_79#_c_335_n 0.00106645f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_275 N_D_c_280_n N_A_196_79#_c_336_n 0.00169995f $X=2.51 $Y=1.485 $X2=0 $Y2=0
cc_276 D N_A_196_79#_c_336_n 0.0117669f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_277 N_D_c_283_n N_A_196_79#_c_336_n 0.00139454f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_278 D N_A_196_79#_c_341_n 0.00682544f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_279 N_D_c_280_n N_A_196_79#_c_342_n 0.00355938f $X=2.51 $Y=1.485 $X2=0 $Y2=0
cc_280 D N_A_196_79#_c_342_n 0.013152f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_281 N_D_M1008_g N_RESET_B_M1016_g 0.0185316f $X=2.45 $Y=2.525 $X2=0 $Y2=0
cc_282 N_D_c_280_n N_RESET_B_M1001_g 0.0253896f $X=2.51 $Y=1.485 $X2=0 $Y2=0
cc_283 D N_RESET_B_M1001_g 0.0100879f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_284 N_D_c_280_n N_RESET_B_c_631_n 0.00881753f $X=2.51 $Y=1.485 $X2=0 $Y2=0
cc_285 D N_RESET_B_c_635_n 0.00625935f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_286 N_D_c_283_n N_RESET_B_c_635_n 0.0253896f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_287 N_D_c_281_n N_RESET_B_c_644_n 0.00742007f $X=2.51 $Y=1.99 $X2=0 $Y2=0
cc_288 N_D_c_281_n N_RESET_B_c_645_n 0.00145948f $X=2.51 $Y=1.99 $X2=0 $Y2=0
cc_289 N_D_c_286_n N_RESET_B_c_645_n 8.64093e-19 $X=2.51 $Y=2.155 $X2=0 $Y2=0
cc_290 D N_RESET_B_c_645_n 0.0473699f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_291 D N_RESET_B_c_646_n 6.3482e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_292 D N_RESET_B_c_637_n 0.00455607f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_293 N_D_c_283_n N_RESET_B_c_637_n 0.00742007f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_294 D N_RESET_B_c_638_n 0.0548266f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_295 N_D_c_283_n N_RESET_B_c_638_n 5.26329e-19 $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_296 N_D_M1008_g N_A_27_79#_c_941_n 0.0100449f $X=2.45 $Y=2.525 $X2=0 $Y2=0
cc_297 N_D_M1008_g N_A_27_79#_c_944_n 0.0164796f $X=2.45 $Y=2.525 $X2=0 $Y2=0
cc_298 N_D_c_286_n N_A_27_79#_c_944_n 0.0118377f $X=2.51 $Y=2.155 $X2=0 $Y2=0
cc_299 N_D_c_281_n N_A_27_79#_c_932_n 0.00486698f $X=2.51 $Y=1.99 $X2=0 $Y2=0
cc_300 N_D_c_280_n N_A_27_79#_c_933_n 0.00896418f $X=2.51 $Y=1.485 $X2=0 $Y2=0
cc_301 D N_A_27_79#_c_933_n 3.64068e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_302 N_D_c_283_n N_A_27_79#_c_933_n 0.00486698f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_303 N_D_c_281_n N_A_27_79#_c_951_n 0.0118377f $X=2.51 $Y=1.99 $X2=0 $Y2=0
cc_304 D N_A_27_79#_c_951_n 4.61148e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_305 N_D_M1008_g N_VPWR_c_1415_n 0.00430022f $X=2.45 $Y=2.525 $X2=0 $Y2=0
cc_306 N_D_M1008_g N_VPWR_c_1413_n 9.39239e-19 $X=2.45 $Y=2.525 $X2=0 $Y2=0
cc_307 D N_A_308_463#_M1027_d 0.00287204f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_308 N_D_M1008_g N_A_308_463#_c_1573_n 0.00847642f $X=2.45 $Y=2.525 $X2=0
+ $Y2=0
cc_309 D N_A_308_463#_c_1573_n 0.0343273f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_310 N_D_c_280_n N_A_308_463#_c_1568_n 0.00477394f $X=2.51 $Y=1.485 $X2=0
+ $Y2=0
cc_311 D N_A_308_463#_c_1568_n 0.0715318f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_312 N_D_c_283_n N_A_308_463#_c_1568_n 0.00399394f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_313 N_D_M1008_g N_A_308_463#_c_1571_n 0.00371719f $X=2.45 $Y=2.525 $X2=0
+ $Y2=0
cc_314 N_D_c_286_n N_A_308_463#_c_1571_n 0.00239771f $X=2.51 $Y=2.155 $X2=0
+ $Y2=0
cc_315 D N_A_308_463#_c_1571_n 0.00866914f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_316 D A_427_191# 0.00100186f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_317 N_A_196_79#_c_339_n N_A_811_341#_M1007_d 0.00860509f $X=6.29 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_318 N_A_196_79#_c_331_n N_A_811_341#_M1034_g 0.0381068f $X=3.845 $Y=1.45
+ $X2=0 $Y2=0
cc_319 N_A_196_79#_c_338_n N_A_811_341#_M1034_g 0.00255041f $X=4.56 $Y=0.715
+ $X2=0 $Y2=0
cc_320 N_A_196_79#_c_345_n N_A_811_341#_M1034_g 0.00559644f $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_321 N_A_196_79#_M1019_g N_A_811_341#_c_519_n 7.76632e-19 $X=3.46 $Y=2.525
+ $X2=0 $Y2=0
cc_322 N_A_196_79#_c_345_n N_A_811_341#_c_519_n 0.0089709f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_323 N_A_196_79#_M1019_g N_A_811_341#_M1000_g 0.00278369f $X=3.46 $Y=2.525
+ $X2=0 $Y2=0
cc_324 N_A_196_79#_c_331_n N_A_811_341#_c_522_n 2.60124e-19 $X=3.845 $Y=1.45
+ $X2=0 $Y2=0
cc_325 N_A_196_79#_c_345_n N_A_811_341#_c_522_n 3.12549e-19 $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_326 N_A_196_79#_c_346_n N_A_811_341#_c_524_n 0.00288694f $X=6.55 $Y=1.555
+ $X2=0 $Y2=0
cc_327 N_A_196_79#_c_332_n N_A_811_341#_c_525_n 0.00288694f $X=6.285 $Y=1.39
+ $X2=0 $Y2=0
cc_328 N_A_196_79#_c_339_n N_A_811_341#_c_525_n 0.0212846f $X=6.29 $Y=0.805
+ $X2=0 $Y2=0
cc_329 N_A_196_79#_c_340_n N_A_811_341#_c_525_n 0.0480309f $X=6.385 $Y=1.555
+ $X2=0 $Y2=0
cc_330 N_A_196_79#_c_350_n N_RESET_B_M1016_g 0.00268993f $X=1.145 $Y=2.515 $X2=0
+ $Y2=0
cc_331 N_A_196_79#_c_351_n N_RESET_B_M1016_g 0.00320043f $X=1.295 $Y=2.305 $X2=0
+ $Y2=0
cc_332 N_A_196_79#_c_334_n N_RESET_B_M1001_g 0.00282489f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_333 N_A_196_79#_c_335_n N_RESET_B_M1001_g 0.011107f $X=2.075 $Y=0.955 $X2=0
+ $Y2=0
cc_334 N_A_196_79#_c_336_n N_RESET_B_M1001_g 8.12301e-19 $X=3.205 $Y=0.715 $X2=0
+ $Y2=0
cc_335 N_A_196_79#_c_341_n N_RESET_B_M1001_g 0.00741517f $X=1.312 $Y=1.935 $X2=0
+ $Y2=0
cc_336 N_A_196_79#_c_342_n N_RESET_B_M1001_g 0.0132086f $X=2.195 $Y=0.715 $X2=0
+ $Y2=0
cc_337 N_A_196_79#_c_331_n N_RESET_B_c_631_n 0.00881437f $X=3.845 $Y=1.45 $X2=0
+ $Y2=0
cc_338 N_A_196_79#_c_336_n N_RESET_B_c_631_n 0.0201374f $X=3.205 $Y=0.715 $X2=0
+ $Y2=0
cc_339 N_A_196_79#_c_338_n N_RESET_B_c_631_n 0.0264802f $X=4.56 $Y=0.715 $X2=0
+ $Y2=0
cc_340 N_A_196_79#_c_342_n N_RESET_B_c_631_n 0.00267555f $X=2.195 $Y=0.715 $X2=0
+ $Y2=0
cc_341 N_A_196_79#_c_343_n N_RESET_B_c_631_n 0.0053441f $X=3.29 $Y=0.715 $X2=0
+ $Y2=0
cc_342 N_A_196_79#_c_338_n N_RESET_B_M1032_g 0.0173357f $X=4.56 $Y=0.715 $X2=0
+ $Y2=0
cc_343 N_A_196_79#_c_339_n N_RESET_B_M1032_g 0.00167209f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_344 N_A_196_79#_c_335_n N_RESET_B_c_635_n 0.00350047f $X=2.075 $Y=0.955 $X2=0
+ $Y2=0
cc_345 N_A_196_79#_c_341_n N_RESET_B_c_635_n 0.00110712f $X=1.312 $Y=1.935 $X2=0
+ $Y2=0
cc_346 N_A_196_79#_M1019_g N_RESET_B_c_645_n 0.0107955f $X=3.46 $Y=2.525 $X2=0
+ $Y2=0
cc_347 N_A_196_79#_c_344_n N_RESET_B_c_645_n 0.0171139f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_348 N_A_196_79#_c_345_n N_RESET_B_c_645_n 0.00709661f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_349 N_A_196_79#_c_341_n N_RESET_B_c_646_n 0.00766499f $X=1.312 $Y=1.935 $X2=0
+ $Y2=0
cc_350 N_A_196_79#_M1031_g N_RESET_B_c_647_n 0.0102691f $X=6.935 $Y=2.69 $X2=0
+ $Y2=0
cc_351 N_A_196_79#_c_340_n N_RESET_B_c_647_n 0.00749067f $X=6.385 $Y=1.555 $X2=0
+ $Y2=0
cc_352 N_A_196_79#_c_346_n N_RESET_B_c_647_n 0.00599408f $X=6.55 $Y=1.555 $X2=0
+ $Y2=0
cc_353 N_A_196_79#_c_354_n N_RESET_B_c_637_n 0.00110712f $X=1.312 $Y=2.155 $X2=0
+ $Y2=0
cc_354 N_A_196_79#_c_335_n N_RESET_B_c_638_n 0.0134823f $X=2.075 $Y=0.955 $X2=0
+ $Y2=0
cc_355 N_A_196_79#_c_341_n N_RESET_B_c_638_n 0.0528734f $X=1.312 $Y=1.935 $X2=0
+ $Y2=0
cc_356 N_A_196_79#_c_337_n N_A_637_191#_M1028_d 0.00729588f $X=3.29 $Y=1.615
+ $X2=-0.19 $Y2=-0.245
cc_357 N_A_196_79#_c_332_n N_A_637_191#_c_824_n 0.0213037f $X=6.285 $Y=1.39
+ $X2=0 $Y2=0
cc_358 N_A_196_79#_c_339_n N_A_637_191#_c_824_n 0.0175928f $X=6.29 $Y=0.805
+ $X2=0 $Y2=0
cc_359 N_A_196_79#_c_340_n N_A_637_191#_c_824_n 6.74483e-19 $X=6.385 $Y=1.555
+ $X2=0 $Y2=0
cc_360 N_A_196_79#_M1019_g N_A_637_191#_c_825_n 0.00460853f $X=3.46 $Y=2.525
+ $X2=0 $Y2=0
cc_361 N_A_196_79#_c_331_n N_A_637_191#_c_825_n 0.00389476f $X=3.845 $Y=1.45
+ $X2=0 $Y2=0
cc_362 N_A_196_79#_c_337_n N_A_637_191#_c_825_n 0.0113315f $X=3.29 $Y=1.615
+ $X2=0 $Y2=0
cc_363 N_A_196_79#_c_344_n N_A_637_191#_c_825_n 0.0252326f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_364 N_A_196_79#_c_345_n N_A_637_191#_c_825_n 0.0104038f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_365 N_A_196_79#_M1019_g N_A_637_191#_c_831_n 2.37983e-19 $X=3.46 $Y=2.525
+ $X2=0 $Y2=0
cc_366 N_A_196_79#_c_344_n N_A_637_191#_c_831_n 0.00109494f $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_367 N_A_196_79#_c_345_n N_A_637_191#_c_831_n 0.00486918f $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_368 N_A_196_79#_c_338_n N_A_637_191#_c_846_n 0.0284286f $X=4.56 $Y=0.715
+ $X2=0 $Y2=0
cc_369 N_A_196_79#_c_339_n N_A_637_191#_c_846_n 0.0621646f $X=6.29 $Y=0.805
+ $X2=0 $Y2=0
cc_370 N_A_196_79#_c_331_n N_A_637_191#_c_848_n 0.00992945f $X=3.845 $Y=1.45
+ $X2=0 $Y2=0
cc_371 N_A_196_79#_c_337_n N_A_637_191#_c_848_n 0.0267332f $X=3.29 $Y=1.615
+ $X2=0 $Y2=0
cc_372 N_A_196_79#_c_338_n N_A_637_191#_c_848_n 0.0467716f $X=4.56 $Y=0.715
+ $X2=0 $Y2=0
cc_373 N_A_196_79#_c_344_n N_A_637_191#_c_848_n 0.00388181f $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_374 N_A_196_79#_c_345_n N_A_637_191#_c_848_n 0.00687444f $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_375 N_A_196_79#_c_339_n N_A_637_191#_c_827_n 7.37384e-19 $X=6.29 $Y=0.805
+ $X2=0 $Y2=0
cc_376 N_A_196_79#_c_346_n N_A_637_191#_c_827_n 0.00867074f $X=6.55 $Y=1.555
+ $X2=0 $Y2=0
cc_377 N_A_196_79#_c_334_n N_A_27_79#_M1006_g 0.00518808f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_378 N_A_196_79#_c_350_n N_A_27_79#_M1020_g 4.50163e-19 $X=1.145 $Y=2.515
+ $X2=0 $Y2=0
cc_379 N_A_196_79#_c_351_n N_A_27_79#_M1020_g 0.00235767f $X=1.295 $Y=2.305
+ $X2=0 $Y2=0
cc_380 N_A_196_79#_c_332_n N_A_27_79#_c_929_n 0.007882f $X=6.285 $Y=1.39 $X2=0
+ $Y2=0
cc_381 N_A_196_79#_c_334_n N_A_27_79#_c_929_n 0.00693171f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_382 N_A_196_79#_c_335_n N_A_27_79#_c_929_n 0.0064402f $X=2.075 $Y=0.955 $X2=0
+ $Y2=0
cc_383 N_A_196_79#_c_338_n N_A_27_79#_c_929_n 0.00368313f $X=4.56 $Y=0.715 $X2=0
+ $Y2=0
cc_384 N_A_196_79#_c_339_n N_A_27_79#_c_929_n 0.0187555f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_385 N_A_196_79#_c_342_n N_A_27_79#_c_929_n 9.31264e-19 $X=2.195 $Y=0.715
+ $X2=0 $Y2=0
cc_386 N_A_196_79#_c_350_n N_A_27_79#_c_941_n 0.00685929f $X=1.145 $Y=2.515
+ $X2=0 $Y2=0
cc_387 N_A_196_79#_c_354_n N_A_27_79#_c_931_n 0.00312265f $X=1.312 $Y=2.155
+ $X2=0 $Y2=0
cc_388 N_A_196_79#_M1019_g N_A_27_79#_c_944_n 0.0253619f $X=3.46 $Y=2.525 $X2=0
+ $Y2=0
cc_389 N_A_196_79#_c_345_n N_A_27_79#_c_944_n 3.1318e-19 $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_390 N_A_196_79#_c_337_n N_A_27_79#_c_932_n 5.71391e-19 $X=3.29 $Y=1.615 $X2=0
+ $Y2=0
cc_391 N_A_196_79#_c_344_n N_A_27_79#_c_932_n 0.00227118f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_392 N_A_196_79#_c_345_n N_A_27_79#_c_932_n 0.0204458f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_393 N_A_196_79#_c_331_n N_A_27_79#_c_933_n 0.00512483f $X=3.845 $Y=1.45 $X2=0
+ $Y2=0
cc_394 N_A_196_79#_c_336_n N_A_27_79#_c_933_n 0.00384262f $X=3.205 $Y=0.715
+ $X2=0 $Y2=0
cc_395 N_A_196_79#_c_337_n N_A_27_79#_c_933_n 0.00894805f $X=3.29 $Y=1.615 $X2=0
+ $Y2=0
cc_396 N_A_196_79#_c_345_n N_A_27_79#_c_933_n 0.00232889f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_397 N_A_196_79#_M1019_g N_A_27_79#_c_946_n 0.0104164f $X=3.46 $Y=2.525 $X2=0
+ $Y2=0
cc_398 N_A_196_79#_M1019_g N_A_27_79#_M1035_g 0.0132354f $X=3.46 $Y=2.525 $X2=0
+ $Y2=0
cc_399 N_A_196_79#_c_345_n N_A_27_79#_M1035_g 0.00142998f $X=3.54 $Y=1.78 $X2=0
+ $Y2=0
cc_400 N_A_196_79#_M1031_g N_A_27_79#_M1024_g 0.0205389f $X=6.935 $Y=2.69 $X2=0
+ $Y2=0
cc_401 N_A_196_79#_c_340_n N_A_27_79#_M1024_g 0.00102182f $X=6.385 $Y=1.555
+ $X2=0 $Y2=0
cc_402 N_A_196_79#_c_346_n N_A_27_79#_M1024_g 0.0101866f $X=6.55 $Y=1.555 $X2=0
+ $Y2=0
cc_403 N_A_196_79#_c_332_n N_A_27_79#_M1015_g 0.00953452f $X=6.285 $Y=1.39 $X2=0
+ $Y2=0
cc_404 N_A_196_79#_c_333_n N_A_27_79#_M1015_g 0.00114049f $X=6.86 $Y=1.645 $X2=0
+ $Y2=0
cc_405 N_A_196_79#_c_351_n N_A_27_79#_c_950_n 0.00926193f $X=1.295 $Y=2.305
+ $X2=0 $Y2=0
cc_406 N_A_196_79#_c_334_n N_A_27_79#_c_936_n 0.0125385f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_407 N_A_196_79#_c_341_n N_A_27_79#_c_936_n 0.0164032f $X=1.312 $Y=1.935 $X2=0
+ $Y2=0
cc_408 N_A_196_79#_c_334_n N_A_27_79#_c_937_n 0.00789011f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_409 N_A_196_79#_c_341_n N_A_27_79#_c_937_n 0.0195166f $X=1.312 $Y=1.935 $X2=0
+ $Y2=0
cc_410 N_A_196_79#_c_333_n N_A_1444_320#_M1037_g 0.00136835f $X=6.86 $Y=1.645
+ $X2=0 $Y2=0
cc_411 N_A_196_79#_M1031_g N_A_1444_320#_c_1098_n 0.0435595f $X=6.935 $Y=2.69
+ $X2=0 $Y2=0
cc_412 N_A_196_79#_c_333_n N_A_1444_320#_c_1103_n 7.38872e-19 $X=6.86 $Y=1.645
+ $X2=0 $Y2=0
cc_413 N_A_196_79#_M1031_g N_A_1444_320#_c_1103_n 0.00178548f $X=6.935 $Y=2.69
+ $X2=0 $Y2=0
cc_414 N_A_196_79#_c_333_n N_A_1444_320#_c_1104_n 0.0435595f $X=6.86 $Y=1.645
+ $X2=0 $Y2=0
cc_415 N_A_196_79#_c_339_n N_A_1272_128#_M1013_d 0.00253806f $X=6.29 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_416 N_A_196_79#_c_340_n N_A_1272_128#_M1013_d 0.00378572f $X=6.385 $Y=1.555
+ $X2=-0.19 $Y2=-0.245
cc_417 N_A_196_79#_c_346_n N_A_1272_128#_c_1210_n 0.00327665f $X=6.55 $Y=1.555
+ $X2=0 $Y2=0
cc_418 N_A_196_79#_c_332_n N_A_1272_128#_c_1196_n 0.00365381f $X=6.285 $Y=1.39
+ $X2=0 $Y2=0
cc_419 N_A_196_79#_c_339_n N_A_1272_128#_c_1196_n 0.0139838f $X=6.29 $Y=0.805
+ $X2=0 $Y2=0
cc_420 N_A_196_79#_c_340_n N_A_1272_128#_c_1196_n 0.0257706f $X=6.385 $Y=1.555
+ $X2=0 $Y2=0
cc_421 N_A_196_79#_c_333_n N_A_1272_128#_c_1197_n 0.00644827f $X=6.86 $Y=1.645
+ $X2=0 $Y2=0
cc_422 N_A_196_79#_c_333_n N_A_1272_128#_c_1198_n 0.0165099f $X=6.86 $Y=1.645
+ $X2=0 $Y2=0
cc_423 N_A_196_79#_M1031_g N_A_1272_128#_c_1198_n 0.0183166f $X=6.935 $Y=2.69
+ $X2=0 $Y2=0
cc_424 N_A_196_79#_c_340_n N_A_1272_128#_c_1198_n 0.0204881f $X=6.385 $Y=1.555
+ $X2=0 $Y2=0
cc_425 N_A_196_79#_c_346_n N_A_1272_128#_c_1198_n 0.00348284f $X=6.55 $Y=1.555
+ $X2=0 $Y2=0
cc_426 N_A_196_79#_c_332_n N_A_1272_128#_c_1199_n 9.1124e-19 $X=6.285 $Y=1.39
+ $X2=0 $Y2=0
cc_427 N_A_196_79#_c_340_n N_A_1272_128#_c_1199_n 0.0158319f $X=6.385 $Y=1.555
+ $X2=0 $Y2=0
cc_428 N_A_196_79#_c_346_n N_A_1272_128#_c_1199_n 0.00103307f $X=6.55 $Y=1.555
+ $X2=0 $Y2=0
cc_429 N_A_196_79#_c_350_n N_VPWR_c_1414_n 0.0203021f $X=1.145 $Y=2.515 $X2=0
+ $Y2=0
cc_430 N_A_196_79#_c_351_n N_VPWR_c_1414_n 0.00722421f $X=1.295 $Y=2.305 $X2=0
+ $Y2=0
cc_431 N_A_196_79#_c_350_n N_VPWR_c_1415_n 0.00973716f $X=1.145 $Y=2.515 $X2=0
+ $Y2=0
cc_432 N_A_196_79#_M1031_g N_VPWR_c_1418_n 0.00165226f $X=6.935 $Y=2.69 $X2=0
+ $Y2=0
cc_433 N_A_196_79#_c_350_n N_VPWR_c_1427_n 0.0174327f $X=1.145 $Y=2.515 $X2=0
+ $Y2=0
cc_434 N_A_196_79#_M1031_g N_VPWR_c_1430_n 0.00534427f $X=6.935 $Y=2.69 $X2=0
+ $Y2=0
cc_435 N_A_196_79#_M1019_g N_VPWR_c_1413_n 9.39239e-19 $X=3.46 $Y=2.525 $X2=0
+ $Y2=0
cc_436 N_A_196_79#_M1031_g N_VPWR_c_1413_n 0.00526787f $X=6.935 $Y=2.69 $X2=0
+ $Y2=0
cc_437 N_A_196_79#_c_350_n N_VPWR_c_1413_n 0.011091f $X=1.145 $Y=2.515 $X2=0
+ $Y2=0
cc_438 N_A_196_79#_M1019_g N_A_308_463#_c_1568_n 0.00139453f $X=3.46 $Y=2.525
+ $X2=0 $Y2=0
cc_439 N_A_196_79#_c_336_n N_A_308_463#_c_1568_n 0.0152777f $X=3.205 $Y=0.715
+ $X2=0 $Y2=0
cc_440 N_A_196_79#_c_337_n N_A_308_463#_c_1568_n 0.0322257f $X=3.29 $Y=1.615
+ $X2=0 $Y2=0
cc_441 N_A_196_79#_c_344_n N_A_308_463#_c_1568_n 0.0258122f $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_442 N_A_196_79#_c_345_n N_A_308_463#_c_1568_n 2.47453e-19 $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_443 N_A_196_79#_c_350_n N_A_308_463#_c_1570_n 0.0184871f $X=1.145 $Y=2.515
+ $X2=0 $Y2=0
cc_444 N_A_196_79#_c_351_n N_A_308_463#_c_1570_n 0.0138514f $X=1.295 $Y=2.305
+ $X2=0 $Y2=0
cc_445 N_A_196_79#_M1019_g N_A_308_463#_c_1571_n 0.00243201f $X=3.46 $Y=2.525
+ $X2=0 $Y2=0
cc_446 N_A_196_79#_c_344_n N_A_308_463#_c_1571_n 0.00441604f $X=3.54 $Y=1.78
+ $X2=0 $Y2=0
cc_447 N_A_196_79#_c_335_n N_VGND_M1001_s 0.00968368f $X=2.075 $Y=0.955 $X2=0
+ $Y2=0
cc_448 N_A_196_79#_c_339_n N_VGND_M1032_d 0.0141895f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_449 N_A_196_79#_c_334_n N_VGND_c_1659_n 0.0259141f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_450 N_A_196_79#_c_335_n N_VGND_c_1659_n 0.0268035f $X=2.075 $Y=0.955 $X2=0
+ $Y2=0
cc_451 N_A_196_79#_c_342_n N_VGND_c_1659_n 0.00541398f $X=2.195 $Y=0.715 $X2=0
+ $Y2=0
cc_452 N_A_196_79#_c_339_n N_VGND_c_1660_n 0.025714f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_453 N_A_196_79#_c_339_n N_VGND_c_1667_n 0.0113618f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_454 N_A_196_79#_c_334_n N_VGND_c_1670_n 0.0140761f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_455 N_A_196_79#_c_336_n N_VGND_c_1671_n 0.0162925f $X=3.205 $Y=0.715 $X2=0
+ $Y2=0
cc_456 N_A_196_79#_c_338_n N_VGND_c_1671_n 0.0254515f $X=4.56 $Y=0.715 $X2=0
+ $Y2=0
cc_457 N_A_196_79#_c_339_n N_VGND_c_1671_n 0.00719708f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_458 N_A_196_79#_c_342_n N_VGND_c_1671_n 0.00454428f $X=2.195 $Y=0.715 $X2=0
+ $Y2=0
cc_459 N_A_196_79#_c_343_n N_VGND_c_1671_n 0.00345508f $X=3.29 $Y=0.715 $X2=0
+ $Y2=0
cc_460 N_A_196_79#_c_332_n N_VGND_c_1682_n 9.54497e-19 $X=6.285 $Y=1.39 $X2=0
+ $Y2=0
cc_461 N_A_196_79#_c_334_n N_VGND_c_1682_n 0.0127335f $X=1.325 $Y=1.04 $X2=0
+ $Y2=0
cc_462 N_A_196_79#_c_336_n N_VGND_c_1682_n 0.0220207f $X=3.205 $Y=0.715 $X2=0
+ $Y2=0
cc_463 N_A_196_79#_c_338_n N_VGND_c_1682_n 0.0345366f $X=4.56 $Y=0.715 $X2=0
+ $Y2=0
cc_464 N_A_196_79#_c_339_n N_VGND_c_1682_n 0.0325179f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_465 N_A_196_79#_c_342_n N_VGND_c_1682_n 0.00607984f $X=2.195 $Y=0.715 $X2=0
+ $Y2=0
cc_466 N_A_196_79#_c_343_n N_VGND_c_1682_n 0.00450883f $X=3.29 $Y=0.715 $X2=0
+ $Y2=0
cc_467 N_A_196_79#_c_342_n A_427_191# 0.00104609f $X=2.195 $Y=0.715 $X2=-0.19
+ $Y2=-0.245
cc_468 N_A_811_341#_M1034_g N_RESET_B_c_631_n 0.00881753f $X=4.23 $Y=1.165 $X2=0
+ $Y2=0
cc_469 N_A_811_341#_M1034_g N_RESET_B_M1032_g 0.0344425f $X=4.23 $Y=1.165 $X2=0
+ $Y2=0
cc_470 N_A_811_341#_c_521_n N_RESET_B_M1032_g 0.00247026f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_471 N_A_811_341#_M1000_g N_RESET_B_M1012_g 0.0212261f $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_472 N_A_811_341#_c_521_n N_RESET_B_c_636_n 0.00655257f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_473 N_A_811_341#_c_519_n N_RESET_B_c_645_n 0.00549094f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_474 N_A_811_341#_M1000_g N_RESET_B_c_645_n 0.00301677f $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_475 N_A_811_341#_c_520_n N_RESET_B_c_645_n 0.01185f $X=4.22 $Y=1.82 $X2=0
+ $Y2=0
cc_476 N_A_811_341#_c_521_n N_RESET_B_c_645_n 0.00384677f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_477 N_A_811_341#_M1025_d N_RESET_B_c_647_n 0.0132501f $X=5.825 $Y=1.895 $X2=0
+ $Y2=0
cc_478 N_A_811_341#_c_521_n N_RESET_B_c_647_n 0.00724899f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_479 N_A_811_341#_c_530_n N_RESET_B_c_647_n 0.0361186f $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_480 N_A_811_341#_c_531_n N_RESET_B_c_647_n 0.0144162f $X=5.26 $Y=1.985 $X2=0
+ $Y2=0
cc_481 N_A_811_341#_c_533_n N_RESET_B_c_647_n 0.013839f $X=6.06 $Y=2.745 $X2=0
+ $Y2=0
cc_482 N_A_811_341#_c_561_p N_RESET_B_c_647_n 0.0156787f $X=6.06 $Y=2.065 $X2=0
+ $Y2=0
cc_483 N_A_811_341#_c_519_n N_RESET_B_c_648_n 7.7286e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_484 N_A_811_341#_M1000_g N_RESET_B_c_648_n 7.54641e-19 $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_485 N_A_811_341#_c_520_n N_RESET_B_c_648_n 0.00136259f $X=4.22 $Y=1.82 $X2=0
+ $Y2=0
cc_486 N_A_811_341#_c_521_n N_RESET_B_c_648_n 0.00412915f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_487 N_A_811_341#_c_531_n N_RESET_B_c_648_n 2.35195e-19 $X=5.26 $Y=1.985 $X2=0
+ $Y2=0
cc_488 N_A_811_341#_c_519_n N_RESET_B_c_649_n 0.00135286f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_489 N_A_811_341#_M1000_g N_RESET_B_c_649_n 9.86771e-19 $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_490 N_A_811_341#_c_520_n N_RESET_B_c_649_n 0.0164096f $X=4.22 $Y=1.82 $X2=0
+ $Y2=0
cc_491 N_A_811_341#_c_521_n N_RESET_B_c_649_n 0.0293134f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_492 N_A_811_341#_c_523_n N_RESET_B_c_649_n 0.00843238f $X=5.175 $Y=1.9 $X2=0
+ $Y2=0
cc_493 N_A_811_341#_c_531_n N_RESET_B_c_649_n 0.0127868f $X=5.26 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_A_811_341#_M1000_g N_RESET_B_c_653_n 0.00582569f $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_495 N_A_811_341#_c_520_n N_RESET_B_c_653_n 2.42948e-19 $X=4.22 $Y=1.82 $X2=0
+ $Y2=0
cc_496 N_A_811_341#_c_521_n N_RESET_B_c_653_n 0.00360183f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_497 N_A_811_341#_c_523_n N_RESET_B_c_653_n 0.00135298f $X=5.175 $Y=1.9 $X2=0
+ $Y2=0
cc_498 N_A_811_341#_c_531_n N_RESET_B_c_653_n 0.00191056f $X=5.26 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A_811_341#_M1034_g N_RESET_B_c_639_n 0.00359153f $X=4.23 $Y=1.165 $X2=0
+ $Y2=0
cc_500 N_A_811_341#_c_519_n N_RESET_B_c_639_n 0.0179185f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_501 N_A_811_341#_c_520_n N_RESET_B_c_639_n 0.0010074f $X=4.22 $Y=1.82 $X2=0
+ $Y2=0
cc_502 N_A_811_341#_c_521_n N_RESET_B_c_639_n 0.00423447f $X=5.09 $Y=1.525 $X2=0
+ $Y2=0
cc_503 N_A_811_341#_c_523_n N_RESET_B_c_639_n 0.00418579f $X=5.175 $Y=1.9 $X2=0
+ $Y2=0
cc_504 N_A_811_341#_c_524_n N_A_637_191#_c_824_n 6.27467e-19 $X=6.035 $Y=1.9
+ $X2=0 $Y2=0
cc_505 N_A_811_341#_c_525_n N_A_637_191#_c_824_n 0.00421799f $X=5.955 $Y=1.155
+ $X2=0 $Y2=0
cc_506 N_A_811_341#_c_523_n N_A_637_191#_M1025_g 0.00380112f $X=5.175 $Y=1.9
+ $X2=0 $Y2=0
cc_507 N_A_811_341#_c_530_n N_A_637_191#_M1025_g 0.0176376f $X=5.95 $Y=1.985
+ $X2=0 $Y2=0
cc_508 N_A_811_341#_c_533_n N_A_637_191#_M1025_g 0.0101559f $X=6.06 $Y=2.745
+ $X2=0 $Y2=0
cc_509 N_A_811_341#_M1034_g N_A_637_191#_c_825_n 0.00212077f $X=4.23 $Y=1.165
+ $X2=0 $Y2=0
cc_510 N_A_811_341#_c_519_n N_A_637_191#_c_825_n 0.00268928f $X=4.25 $Y=1.985
+ $X2=0 $Y2=0
cc_511 N_A_811_341#_M1000_g N_A_637_191#_c_825_n 0.00323797f $X=4.25 $Y=2.525
+ $X2=0 $Y2=0
cc_512 N_A_811_341#_c_520_n N_A_637_191#_c_825_n 0.029906f $X=4.22 $Y=1.82 $X2=0
+ $Y2=0
cc_513 N_A_811_341#_c_522_n N_A_637_191#_c_825_n 0.0143537f $X=4.305 $Y=1.525
+ $X2=0 $Y2=0
cc_514 N_A_811_341#_c_519_n N_A_637_191#_c_830_n 0.00393537f $X=4.25 $Y=1.985
+ $X2=0 $Y2=0
cc_515 N_A_811_341#_M1000_g N_A_637_191#_c_830_n 0.0113848f $X=4.25 $Y=2.525
+ $X2=0 $Y2=0
cc_516 N_A_811_341#_c_520_n N_A_637_191#_c_830_n 0.00614672f $X=4.22 $Y=1.82
+ $X2=0 $Y2=0
cc_517 N_A_811_341#_c_531_n N_A_637_191#_c_830_n 0.00127506f $X=5.26 $Y=1.985
+ $X2=0 $Y2=0
cc_518 N_A_811_341#_M1034_g N_A_637_191#_c_846_n 0.00539263f $X=4.23 $Y=1.165
+ $X2=0 $Y2=0
cc_519 N_A_811_341#_c_521_n N_A_637_191#_c_846_n 0.0628915f $X=5.09 $Y=1.525
+ $X2=0 $Y2=0
cc_520 N_A_811_341#_c_522_n N_A_637_191#_c_846_n 0.00505695f $X=4.305 $Y=1.525
+ $X2=0 $Y2=0
cc_521 N_A_811_341#_c_530_n N_A_637_191#_c_846_n 0.00479835f $X=5.95 $Y=1.985
+ $X2=0 $Y2=0
cc_522 N_A_811_341#_M1034_g N_A_637_191#_c_848_n 0.00835823f $X=4.23 $Y=1.165
+ $X2=0 $Y2=0
cc_523 N_A_811_341#_c_519_n N_A_637_191#_c_848_n 0.00192612f $X=4.25 $Y=1.985
+ $X2=0 $Y2=0
cc_524 N_A_811_341#_c_522_n N_A_637_191#_c_848_n 0.00688432f $X=4.305 $Y=1.525
+ $X2=0 $Y2=0
cc_525 N_A_811_341#_c_521_n N_A_637_191#_c_826_n 0.0138148f $X=5.09 $Y=1.525
+ $X2=0 $Y2=0
cc_526 N_A_811_341#_c_523_n N_A_637_191#_c_826_n 0.00789367f $X=5.175 $Y=1.9
+ $X2=0 $Y2=0
cc_527 N_A_811_341#_c_530_n N_A_637_191#_c_826_n 0.0127445f $X=5.95 $Y=1.985
+ $X2=0 $Y2=0
cc_528 N_A_811_341#_c_524_n N_A_637_191#_c_826_n 0.0178408f $X=6.035 $Y=1.9
+ $X2=0 $Y2=0
cc_529 N_A_811_341#_c_525_n N_A_637_191#_c_826_n 0.00374369f $X=5.955 $Y=1.155
+ $X2=0 $Y2=0
cc_530 N_A_811_341#_c_521_n N_A_637_191#_c_827_n 0.00216925f $X=5.09 $Y=1.525
+ $X2=0 $Y2=0
cc_531 N_A_811_341#_c_523_n N_A_637_191#_c_827_n 0.00128747f $X=5.175 $Y=1.9
+ $X2=0 $Y2=0
cc_532 N_A_811_341#_c_530_n N_A_637_191#_c_827_n 0.00321696f $X=5.95 $Y=1.985
+ $X2=0 $Y2=0
cc_533 N_A_811_341#_c_524_n N_A_637_191#_c_827_n 0.00992828f $X=6.035 $Y=1.9
+ $X2=0 $Y2=0
cc_534 N_A_811_341#_c_525_n N_A_637_191#_c_827_n 3.54818e-19 $X=5.955 $Y=1.155
+ $X2=0 $Y2=0
cc_535 N_A_811_341#_M1000_g N_A_27_79#_M1035_g 0.0415361f $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_536 N_A_811_341#_M1000_g N_A_27_79#_c_948_n 0.0100709f $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_537 N_A_811_341#_c_533_n N_A_27_79#_c_948_n 0.00483184f $X=6.06 $Y=2.745
+ $X2=0 $Y2=0
cc_538 N_A_811_341#_c_533_n N_A_27_79#_M1024_g 0.00888318f $X=6.06 $Y=2.745
+ $X2=0 $Y2=0
cc_539 N_A_811_341#_c_561_p N_A_27_79#_M1024_g 0.00143143f $X=6.06 $Y=2.065
+ $X2=0 $Y2=0
cc_540 N_A_811_341#_c_533_n N_A_1272_128#_c_1210_n 0.0186837f $X=6.06 $Y=2.745
+ $X2=0 $Y2=0
cc_541 N_A_811_341#_c_561_p N_A_1272_128#_c_1210_n 9.06256e-19 $X=6.06 $Y=2.065
+ $X2=0 $Y2=0
cc_542 N_A_811_341#_c_524_n N_A_1272_128#_c_1198_n 0.0063049f $X=6.035 $Y=1.9
+ $X2=0 $Y2=0
cc_543 N_A_811_341#_c_561_p N_A_1272_128#_c_1198_n 0.00429906f $X=6.06 $Y=2.065
+ $X2=0 $Y2=0
cc_544 N_A_811_341#_c_530_n N_VPWR_M1025_s 0.00366342f $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_545 N_A_811_341#_M1000_g N_VPWR_c_1416_n 0.00429952f $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_546 N_A_811_341#_c_530_n N_VPWR_c_1417_n 0.0200875f $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_547 N_A_811_341#_c_533_n N_VPWR_c_1417_n 0.0376436f $X=6.06 $Y=2.745 $X2=0
+ $Y2=0
cc_548 N_A_811_341#_c_533_n N_VPWR_c_1430_n 0.00739966f $X=6.06 $Y=2.745 $X2=0
+ $Y2=0
cc_549 N_A_811_341#_M1000_g N_VPWR_c_1413_n 9.39239e-19 $X=4.25 $Y=2.525 $X2=0
+ $Y2=0
cc_550 N_A_811_341#_c_533_n N_VPWR_c_1413_n 0.00667223f $X=6.06 $Y=2.745 $X2=0
+ $Y2=0
cc_551 N_RESET_B_c_647_n N_A_637_191#_M1025_g 0.0061151f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_552 N_RESET_B_c_653_n N_A_637_191#_M1025_g 0.00405126f $X=4.825 $Y=1.955
+ $X2=0 $Y2=0
cc_553 N_RESET_B_c_645_n N_A_637_191#_c_825_n 0.0203507f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_648_n N_A_637_191#_c_825_n 0.00148346f $X=4.705 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_649_n N_A_637_191#_c_825_n 0.00197853f $X=4.56 $Y=2.035 $X2=0
+ $Y2=0
cc_556 N_RESET_B_M1012_g N_A_637_191#_c_830_n 0.0143386f $X=4.8 $Y=2.525 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_645_n N_A_637_191#_c_830_n 0.0152059f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_647_n N_A_637_191#_c_830_n 0.0102274f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_648_n N_A_637_191#_c_830_n 0.00941699f $X=4.705 $Y=2.035
+ $X2=0 $Y2=0
cc_560 N_RESET_B_c_649_n N_A_637_191#_c_830_n 0.027894f $X=4.56 $Y=2.035 $X2=0
+ $Y2=0
cc_561 N_RESET_B_c_653_n N_A_637_191#_c_830_n 0.00392088f $X=4.825 $Y=1.955
+ $X2=0 $Y2=0
cc_562 N_RESET_B_c_645_n N_A_637_191#_c_831_n 0.0109728f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_563 N_RESET_B_M1032_g N_A_637_191#_c_846_n 0.0140326f $X=4.655 $Y=1.165 $X2=0
+ $Y2=0
cc_564 N_RESET_B_M1032_g N_A_637_191#_c_848_n 4.85016e-19 $X=4.655 $Y=1.165
+ $X2=0 $Y2=0
cc_565 N_RESET_B_c_647_n N_A_637_191#_c_826_n 0.00128557f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_566 N_RESET_B_M1032_g N_A_637_191#_c_827_n 0.00143425f $X=4.655 $Y=1.165
+ $X2=0 $Y2=0
cc_567 N_RESET_B_c_636_n N_A_637_191#_c_827_n 0.0036356f $X=4.677 $Y=1.56 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_632_n N_A_27_79#_c_929_n 0.161595f $X=2.135 $Y=0.54 $X2=0
+ $Y2=0
cc_569 N_RESET_B_M1016_g N_A_27_79#_c_941_n 0.0100449f $X=1.88 $Y=2.525 $X2=0
+ $Y2=0
cc_570 N_RESET_B_c_635_n N_A_27_79#_c_931_n 0.00627607f $X=2.06 $Y=1.56 $X2=0
+ $Y2=0
cc_571 N_RESET_B_c_645_n N_A_27_79#_c_944_n 0.00105595f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_572 N_RESET_B_c_631_n N_A_27_79#_c_933_n 0.00881596f $X=4.58 $Y=0.54 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_645_n N_A_27_79#_c_933_n 4.76806e-19 $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_574 N_RESET_B_M1012_g N_A_27_79#_c_948_n 0.0100824f $X=4.8 $Y=2.525 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_647_n N_A_27_79#_M1024_g 0.0101661f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_576 N_RESET_B_M1016_g N_A_27_79#_c_950_n 0.00143956f $X=1.88 $Y=2.525 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_637_n N_A_27_79#_c_950_n 0.00627607f $X=1.795 $Y=1.65 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_645_n N_A_27_79#_c_951_n 0.00393457f $X=4.415 $Y=2.035 $X2=0
+ $Y2=0
cc_579 N_RESET_B_M1011_g N_A_1444_320#_M1036_g 0.00631849f $X=8.11 $Y=2.69 $X2=0
+ $Y2=0
cc_580 N_RESET_B_c_655_n N_A_1444_320#_M1036_g 3.3445e-19 $X=8.11 $Y=2.115 $X2=0
+ $Y2=0
cc_581 N_RESET_B_M1003_g N_A_1444_320#_M1037_g 0.03361f $X=7.835 $Y=0.85 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_647_n N_A_1444_320#_c_1097_n 0.00137917f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_655_n N_A_1444_320#_c_1097_n 0.0216196f $X=8.11 $Y=2.115
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_656_n N_A_1444_320#_c_1097_n 0.00109517f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_585 N_RESET_B_M1003_g N_A_1444_320#_c_1099_n 0.0114281f $X=7.835 $Y=0.85
+ $X2=0 $Y2=0
cc_586 N_RESET_B_c_647_n N_A_1444_320#_c_1099_n 0.0095383f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_587 RESET_B N_A_1444_320#_c_1099_n 0.00799866f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_588 N_RESET_B_c_655_n N_A_1444_320#_c_1099_n 0.00557608f $X=8.11 $Y=2.115
+ $X2=0 $Y2=0
cc_589 N_RESET_B_c_656_n N_A_1444_320#_c_1099_n 0.0178895f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_590 N_RESET_B_M1003_g N_A_1444_320#_c_1100_n 0.00179055f $X=7.835 $Y=0.85
+ $X2=0 $Y2=0
cc_591 RESET_B N_A_1444_320#_c_1100_n 0.00683437f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_592 N_RESET_B_c_655_n N_A_1444_320#_c_1100_n 0.00828798f $X=8.11 $Y=2.115
+ $X2=0 $Y2=0
cc_593 N_RESET_B_c_656_n N_A_1444_320#_c_1100_n 0.0230474f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_594 N_RESET_B_M1003_g N_A_1444_320#_c_1093_n 7.93776e-19 $X=7.835 $Y=0.85
+ $X2=0 $Y2=0
cc_595 N_RESET_B_M1003_g N_A_1444_320#_c_1103_n 0.00182999f $X=7.835 $Y=0.85
+ $X2=0 $Y2=0
cc_596 N_RESET_B_c_647_n N_A_1444_320#_c_1103_n 0.0238107f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_597 RESET_B N_A_1444_320#_c_1103_n 0.00125932f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_598 N_RESET_B_c_656_n N_A_1444_320#_c_1103_n 0.0180739f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_599 N_RESET_B_M1003_g N_A_1444_320#_c_1104_n 0.0216196f $X=7.835 $Y=0.85
+ $X2=0 $Y2=0
cc_600 N_RESET_B_c_647_n N_A_1272_128#_M1024_d 0.00125515f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_601 N_RESET_B_M1003_g N_A_1272_128#_c_1182_n 0.05024f $X=7.835 $Y=0.85 $X2=0
+ $Y2=0
cc_602 N_RESET_B_M1003_g N_A_1272_128#_M1017_g 0.0082055f $X=7.835 $Y=0.85 $X2=0
+ $Y2=0
cc_603 N_RESET_B_c_655_n N_A_1272_128#_M1017_g 0.028768f $X=8.11 $Y=2.115 $X2=0
+ $Y2=0
cc_604 N_RESET_B_c_656_n N_A_1272_128#_M1017_g 3.07357e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_605 N_RESET_B_M1003_g N_A_1272_128#_c_1184_n 0.00764743f $X=7.835 $Y=0.85
+ $X2=0 $Y2=0
cc_606 N_RESET_B_c_655_n N_A_1272_128#_c_1184_n 8.2446e-19 $X=8.11 $Y=2.115
+ $X2=0 $Y2=0
cc_607 N_RESET_B_c_647_n N_A_1272_128#_c_1210_n 0.0243493f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_RESET_B_M1003_g N_A_1272_128#_c_1197_n 0.015056f $X=7.835 $Y=0.85 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_647_n N_A_1272_128#_c_1197_n 0.0129844f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_RESET_B_c_647_n N_A_1272_128#_c_1198_n 0.00985101f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_611 N_RESET_B_c_647_n N_VPWR_M1025_s 0.00202f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_612 N_RESET_B_M1016_g N_VPWR_c_1415_n 0.00254223f $X=1.88 $Y=2.525 $X2=0
+ $Y2=0
cc_613 N_RESET_B_M1012_g N_VPWR_c_1416_n 0.00429952f $X=4.8 $Y=2.525 $X2=0 $Y2=0
cc_614 N_RESET_B_M1012_g N_VPWR_c_1417_n 0.00600604f $X=4.8 $Y=2.525 $X2=0 $Y2=0
cc_615 N_RESET_B_c_647_n N_VPWR_c_1417_n 0.00882035f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_616 N_RESET_B_M1011_g N_VPWR_c_1418_n 0.00303577f $X=8.11 $Y=2.69 $X2=0 $Y2=0
cc_617 N_RESET_B_c_647_n N_VPWR_c_1418_n 0.0100416f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_618 RESET_B N_VPWR_c_1418_n 0.00160242f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_619 N_RESET_B_c_655_n N_VPWR_c_1418_n 0.00181082f $X=8.11 $Y=2.115 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_656_n N_VPWR_c_1418_n 0.0133104f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_621 N_RESET_B_M1011_g N_VPWR_c_1431_n 0.00534427f $X=8.11 $Y=2.69 $X2=0 $Y2=0
cc_622 N_RESET_B_M1016_g N_VPWR_c_1413_n 9.39239e-19 $X=1.88 $Y=2.525 $X2=0
+ $Y2=0
cc_623 N_RESET_B_M1012_g N_VPWR_c_1413_n 9.39239e-19 $X=4.8 $Y=2.525 $X2=0 $Y2=0
cc_624 N_RESET_B_M1011_g N_VPWR_c_1413_n 0.00526787f $X=8.11 $Y=2.69 $X2=0 $Y2=0
cc_625 N_RESET_B_M1016_g N_A_308_463#_c_1573_n 0.00868565f $X=1.88 $Y=2.525
+ $X2=0 $Y2=0
cc_626 N_RESET_B_c_635_n N_A_308_463#_c_1573_n 0.00200701f $X=2.06 $Y=1.56 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_645_n N_A_308_463#_c_1573_n 0.0106423f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_628 N_RESET_B_c_646_n N_A_308_463#_c_1573_n 5.50958e-19 $X=1.825 $Y=2.035
+ $X2=0 $Y2=0
cc_629 N_RESET_B_c_638_n N_A_308_463#_c_1573_n 0.00822764f $X=1.795 $Y=1.65
+ $X2=0 $Y2=0
cc_630 N_RESET_B_c_645_n N_A_308_463#_c_1568_n 0.0325106f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_631 N_RESET_B_c_644_n N_A_308_463#_c_1570_n 8.85503e-19 $X=1.795 $Y=2.155
+ $X2=0 $Y2=0
cc_632 N_RESET_B_c_646_n N_A_308_463#_c_1570_n 0.00313019f $X=1.825 $Y=2.035
+ $X2=0 $Y2=0
cc_633 N_RESET_B_c_638_n N_A_308_463#_c_1570_n 0.0126646f $X=1.795 $Y=1.65 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_645_n N_A_308_463#_c_1571_n 0.0230897f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_635 N_RESET_B_c_632_n N_VGND_c_1659_n 0.00945428f $X=2.135 $Y=0.54 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_631_n N_VGND_c_1660_n 0.00262778f $X=4.58 $Y=0.54 $X2=0 $Y2=0
cc_637 N_RESET_B_M1003_g N_VGND_c_1661_n 0.0111122f $X=7.835 $Y=0.85 $X2=0 $Y2=0
cc_638 N_RESET_B_M1003_g N_VGND_c_1672_n 0.00338717f $X=7.835 $Y=0.85 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_632_n N_VGND_c_1682_n 0.0150436f $X=2.135 $Y=0.54 $X2=0 $Y2=0
cc_640 N_RESET_B_M1003_g N_VGND_c_1682_n 0.00390857f $X=7.835 $Y=0.85 $X2=0
+ $Y2=0
cc_641 N_A_637_191#_c_824_n N_A_27_79#_c_929_n 0.00788265f $X=5.74 $Y=1.39 $X2=0
+ $Y2=0
cc_642 N_A_637_191#_c_831_n N_A_27_79#_c_946_n 0.00335258f $X=3.985 $Y=2.385
+ $X2=0 $Y2=0
cc_643 N_A_637_191#_c_825_n N_A_27_79#_M1035_g 0.00656721f $X=3.88 $Y=2.3 $X2=0
+ $Y2=0
cc_644 N_A_637_191#_c_831_n N_A_27_79#_M1035_g 0.0115272f $X=3.985 $Y=2.385
+ $X2=0 $Y2=0
cc_645 N_A_637_191#_M1025_g N_A_27_79#_c_948_n 0.0103107f $X=5.75 $Y=2.315 $X2=0
+ $Y2=0
cc_646 N_A_637_191#_c_830_n N_A_27_79#_c_948_n 0.00817682f $X=4.87 $Y=2.385
+ $X2=0 $Y2=0
cc_647 N_A_637_191#_M1025_g N_A_27_79#_M1024_g 0.0146248f $X=5.75 $Y=2.315 $X2=0
+ $Y2=0
cc_648 N_A_637_191#_c_830_n N_VPWR_M1000_d 0.00315285f $X=4.87 $Y=2.385 $X2=0
+ $Y2=0
cc_649 N_A_637_191#_c_830_n N_VPWR_c_1416_n 0.0207781f $X=4.87 $Y=2.385 $X2=0
+ $Y2=0
cc_650 N_A_637_191#_M1025_g N_VPWR_c_1417_n 0.0141302f $X=5.75 $Y=2.315 $X2=0
+ $Y2=0
cc_651 N_A_637_191#_c_830_n N_VPWR_c_1417_n 0.0260566f $X=4.87 $Y=2.385 $X2=0
+ $Y2=0
cc_652 N_A_637_191#_c_831_n N_VPWR_c_1428_n 0.00775274f $X=3.985 $Y=2.385 $X2=0
+ $Y2=0
cc_653 N_A_637_191#_c_830_n N_VPWR_c_1429_n 0.00441176f $X=4.87 $Y=2.385 $X2=0
+ $Y2=0
cc_654 N_A_637_191#_M1025_g N_VPWR_c_1413_n 7.88961e-19 $X=5.75 $Y=2.315 $X2=0
+ $Y2=0
cc_655 N_A_637_191#_c_830_n N_VPWR_c_1413_n 0.0233341f $X=4.87 $Y=2.385 $X2=0
+ $Y2=0
cc_656 N_A_637_191#_c_831_n N_VPWR_c_1413_n 0.0118236f $X=3.985 $Y=2.385 $X2=0
+ $Y2=0
cc_657 N_A_637_191#_c_825_n N_A_308_463#_c_1571_n 0.00589641f $X=3.88 $Y=2.3
+ $X2=0 $Y2=0
cc_658 N_A_637_191#_c_831_n N_A_308_463#_c_1571_n 6.73614e-19 $X=3.985 $Y=2.385
+ $X2=0 $Y2=0
cc_659 N_A_637_191#_c_830_n A_793_463# 0.00124295f $X=4.87 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_660 N_A_637_191#_c_846_n N_VGND_M1032_d 0.0234753f $X=5.43 $Y=1.16 $X2=0
+ $Y2=0
cc_661 N_A_637_191#_c_826_n N_VGND_M1032_d 7.34787e-19 $X=5.525 $Y=1.555 $X2=0
+ $Y2=0
cc_662 N_A_637_191#_c_824_n N_VGND_c_1660_n 0.00161872f $X=5.74 $Y=1.39 $X2=0
+ $Y2=0
cc_663 N_A_637_191#_c_824_n N_VGND_c_1682_n 9.54497e-19 $X=5.74 $Y=1.39 $X2=0
+ $Y2=0
cc_664 N_A_637_191#_c_848_n A_784_191# 0.00493373f $X=4.235 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_665 N_A_637_191#_c_846_n A_861_191# 0.00358338f $X=5.43 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_666 N_A_27_79#_M1015_g N_A_1444_320#_M1037_g 0.040708f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_667 N_A_27_79#_M1024_g N_A_1272_128#_c_1210_n 0.00142005f $X=6.41 $Y=2.48
+ $X2=0 $Y2=0
cc_668 N_A_27_79#_c_929_n N_A_1272_128#_c_1196_n 0.00385409f $X=6.97 $Y=0.18
+ $X2=0 $Y2=0
cc_669 N_A_27_79#_M1015_g N_A_1272_128#_c_1196_n 0.0100435f $X=7.045 $Y=0.85
+ $X2=0 $Y2=0
cc_670 N_A_27_79#_M1015_g N_A_1272_128#_c_1197_n 0.0063885f $X=7.045 $Y=0.85
+ $X2=0 $Y2=0
cc_671 N_A_27_79#_M1024_g N_A_1272_128#_c_1198_n 9.60337e-19 $X=6.41 $Y=2.48
+ $X2=0 $Y2=0
cc_672 N_A_27_79#_M1020_g N_VPWR_c_1414_n 0.0109938f $X=0.93 $Y=2.68 $X2=0 $Y2=0
cc_673 N_A_27_79#_c_942_n N_VPWR_c_1414_n 0.0071807f $X=1.005 $Y=3.15 $X2=0
+ $Y2=0
cc_674 N_A_27_79#_c_954_n N_VPWR_c_1414_n 0.0274284f $X=0.25 $Y=2.465 $X2=0
+ $Y2=0
cc_675 N_A_27_79#_c_941_n N_VPWR_c_1415_n 0.0264276f $X=2.885 $Y=3.15 $X2=0
+ $Y2=0
cc_676 N_A_27_79#_c_944_n N_VPWR_c_1415_n 0.00557219f $X=2.96 $Y=3.075 $X2=0
+ $Y2=0
cc_677 N_A_27_79#_M1035_g N_VPWR_c_1416_n 0.0063441f $X=3.89 $Y=2.525 $X2=0
+ $Y2=0
cc_678 N_A_27_79#_c_948_n N_VPWR_c_1416_n 0.0254009f $X=6.335 $Y=3.15 $X2=0
+ $Y2=0
cc_679 N_A_27_79#_c_948_n N_VPWR_c_1417_n 0.025796f $X=6.335 $Y=3.15 $X2=0 $Y2=0
cc_680 N_A_27_79#_M1024_g N_VPWR_c_1417_n 0.00384505f $X=6.41 $Y=2.48 $X2=0
+ $Y2=0
cc_681 N_A_27_79#_c_955_n N_VPWR_c_1426_n 0.0137038f $X=0.285 $Y=2.515 $X2=0
+ $Y2=0
cc_682 N_A_27_79#_c_942_n N_VPWR_c_1427_n 0.0329955f $X=1.005 $Y=3.15 $X2=0
+ $Y2=0
cc_683 N_A_27_79#_c_941_n N_VPWR_c_1428_n 0.0597153f $X=2.885 $Y=3.15 $X2=0
+ $Y2=0
cc_684 N_A_27_79#_c_948_n N_VPWR_c_1429_n 0.0212709f $X=6.335 $Y=3.15 $X2=0
+ $Y2=0
cc_685 N_A_27_79#_c_948_n N_VPWR_c_1430_n 0.0257875f $X=6.335 $Y=3.15 $X2=0
+ $Y2=0
cc_686 N_A_27_79#_c_941_n N_VPWR_c_1413_n 0.046746f $X=2.885 $Y=3.15 $X2=0 $Y2=0
cc_687 N_A_27_79#_c_942_n N_VPWR_c_1413_n 0.00749832f $X=1.005 $Y=3.15 $X2=0
+ $Y2=0
cc_688 N_A_27_79#_c_946_n N_VPWR_c_1413_n 0.0222444f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_689 N_A_27_79#_c_948_n N_VPWR_c_1413_n 0.0742071f $X=6.335 $Y=3.15 $X2=0
+ $Y2=0
cc_690 N_A_27_79#_c_952_n N_VPWR_c_1413_n 0.00421372f $X=2.96 $Y=3.15 $X2=0
+ $Y2=0
cc_691 N_A_27_79#_c_953_n N_VPWR_c_1413_n 0.00421372f $X=3.89 $Y=3.15 $X2=0
+ $Y2=0
cc_692 N_A_27_79#_c_955_n N_VPWR_c_1413_n 0.00975186f $X=0.285 $Y=2.515 $X2=0
+ $Y2=0
cc_693 N_A_27_79#_c_941_n N_A_308_463#_c_1573_n 0.00199547f $X=2.885 $Y=3.15
+ $X2=0 $Y2=0
cc_694 N_A_27_79#_c_944_n N_A_308_463#_c_1568_n 0.00589298f $X=2.96 $Y=3.075
+ $X2=0 $Y2=0
cc_695 N_A_27_79#_c_932_n N_A_308_463#_c_1568_n 0.00459821f $X=3.09 $Y=1.785
+ $X2=0 $Y2=0
cc_696 N_A_27_79#_c_933_n N_A_308_463#_c_1568_n 0.00362455f $X=3.11 $Y=1.45
+ $X2=0 $Y2=0
cc_697 N_A_27_79#_c_951_n N_A_308_463#_c_1568_n 0.00709685f $X=3.09 $Y=1.86
+ $X2=0 $Y2=0
cc_698 N_A_27_79#_c_941_n N_A_308_463#_c_1570_n 0.003815f $X=2.885 $Y=3.15 $X2=0
+ $Y2=0
cc_699 N_A_27_79#_c_941_n N_A_308_463#_c_1571_n 0.00442011f $X=2.885 $Y=3.15
+ $X2=0 $Y2=0
cc_700 N_A_27_79#_c_944_n N_A_308_463#_c_1571_n 0.0257295f $X=2.96 $Y=3.075
+ $X2=0 $Y2=0
cc_701 N_A_27_79#_c_946_n N_A_308_463#_c_1571_n 0.00447307f $X=3.815 $Y=3.15
+ $X2=0 $Y2=0
cc_702 N_A_27_79#_c_951_n N_A_308_463#_c_1571_n 0.00611822f $X=3.09 $Y=1.86
+ $X2=0 $Y2=0
cc_703 N_A_27_79#_c_930_n N_VGND_c_1658_n 0.0103152f $X=0.98 $Y=0.18 $X2=0 $Y2=0
cc_704 N_A_27_79#_c_936_n N_VGND_c_1658_n 0.0180563f $X=0.95 $Y=1.09 $X2=0 $Y2=0
cc_705 N_A_27_79#_M1006_g N_VGND_c_1659_n 0.00368838f $X=0.905 $Y=0.605 $X2=0
+ $Y2=0
cc_706 N_A_27_79#_c_929_n N_VGND_c_1659_n 0.0254714f $X=6.97 $Y=0.18 $X2=0 $Y2=0
cc_707 N_A_27_79#_c_929_n N_VGND_c_1660_n 0.0248335f $X=6.97 $Y=0.18 $X2=0 $Y2=0
cc_708 N_A_27_79#_c_929_n N_VGND_c_1661_n 0.0115518f $X=6.97 $Y=0.18 $X2=0 $Y2=0
cc_709 N_A_27_79#_M1015_g N_VGND_c_1661_n 0.00173779f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_710 N_A_27_79#_c_929_n N_VGND_c_1667_n 0.0444293f $X=6.97 $Y=0.18 $X2=0 $Y2=0
cc_711 N_A_27_79#_c_935_n N_VGND_c_1669_n 0.00836745f $X=0.26 $Y=0.59 $X2=0
+ $Y2=0
cc_712 N_A_27_79#_c_930_n N_VGND_c_1670_n 0.0217311f $X=0.98 $Y=0.18 $X2=0 $Y2=0
cc_713 N_A_27_79#_c_929_n N_VGND_c_1671_n 0.0842794f $X=6.97 $Y=0.18 $X2=0 $Y2=0
cc_714 N_A_27_79#_c_929_n N_VGND_c_1682_n 0.17041f $X=6.97 $Y=0.18 $X2=0 $Y2=0
cc_715 N_A_27_79#_c_930_n N_VGND_c_1682_n 0.0113334f $X=0.98 $Y=0.18 $X2=0 $Y2=0
cc_716 N_A_27_79#_c_935_n N_VGND_c_1682_n 0.00979051f $X=0.26 $Y=0.59 $X2=0
+ $Y2=0
cc_717 N_A_1444_320#_c_1093_n N_A_1272_128#_c_1182_n 0.00518837f $X=8.745
+ $Y=0.945 $X2=0 $Y2=0
cc_718 N_A_1444_320#_c_1094_n N_A_1272_128#_c_1182_n 0.00261146f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_719 N_A_1444_320#_c_1100_n N_A_1272_128#_M1017_g 0.0209504f $X=8.325 $Y=2.69
+ $X2=0 $Y2=0
cc_720 N_A_1444_320#_c_1101_n N_A_1272_128#_M1017_g 0.0121089f $X=8.745 $Y=1.685
+ $X2=0 $Y2=0
cc_721 N_A_1444_320#_c_1094_n N_A_1272_128#_M1017_g 0.00247268f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_722 N_A_1444_320#_c_1105_n N_A_1272_128#_M1017_g 0.00432208f $X=8.355 $Y=1.69
+ $X2=0 $Y2=0
cc_723 N_A_1444_320#_c_1093_n N_A_1272_128#_c_1183_n 0.00319647f $X=8.745
+ $Y=0.945 $X2=0 $Y2=0
cc_724 N_A_1444_320#_c_1101_n N_A_1272_128#_c_1183_n 9.93321e-19 $X=8.745
+ $Y=1.685 $X2=0 $Y2=0
cc_725 N_A_1444_320#_c_1094_n N_A_1272_128#_c_1183_n 0.0162673f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_726 N_A_1444_320#_c_1099_n N_A_1272_128#_c_1184_n 3.81724e-19 $X=8.22 $Y=1.69
+ $X2=0 $Y2=0
cc_727 N_A_1444_320#_c_1093_n N_A_1272_128#_c_1184_n 0.0093527f $X=8.745
+ $Y=0.945 $X2=0 $Y2=0
cc_728 N_A_1444_320#_c_1094_n N_A_1272_128#_c_1184_n 0.00303117f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_729 N_A_1444_320#_c_1105_n N_A_1272_128#_c_1184_n 0.00607159f $X=8.355
+ $Y=1.69 $X2=0 $Y2=0
cc_730 N_A_1444_320#_c_1100_n N_A_1272_128#_M1009_g 4.83721e-19 $X=8.325 $Y=2.69
+ $X2=0 $Y2=0
cc_731 N_A_1444_320#_c_1101_n N_A_1272_128#_M1009_g 0.0052769f $X=8.745 $Y=1.685
+ $X2=0 $Y2=0
cc_732 N_A_1444_320#_c_1094_n N_A_1272_128#_M1009_g 0.00218965f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_733 N_A_1444_320#_c_1094_n N_A_1272_128#_M1010_g 0.00392194f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_734 N_A_1444_320#_c_1094_n N_A_1272_128#_c_1192_n 0.00335286f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_735 N_A_1444_320#_M1037_g N_A_1272_128#_c_1196_n 0.00203381f $X=7.405 $Y=0.85
+ $X2=0 $Y2=0
cc_736 N_A_1444_320#_M1037_g N_A_1272_128#_c_1197_n 0.0173892f $X=7.405 $Y=0.85
+ $X2=0 $Y2=0
cc_737 N_A_1444_320#_c_1099_n N_A_1272_128#_c_1197_n 0.0485743f $X=8.22 $Y=1.69
+ $X2=0 $Y2=0
cc_738 N_A_1444_320#_c_1093_n N_A_1272_128#_c_1197_n 0.0237006f $X=8.745
+ $Y=0.945 $X2=0 $Y2=0
cc_739 N_A_1444_320#_c_1101_n N_A_1272_128#_c_1197_n 0.00509352f $X=8.745
+ $Y=1.685 $X2=0 $Y2=0
cc_740 N_A_1444_320#_c_1094_n N_A_1272_128#_c_1197_n 0.014602f $X=8.885 $Y=1.6
+ $X2=0 $Y2=0
cc_741 N_A_1444_320#_c_1103_n N_A_1272_128#_c_1197_n 0.0252419f $X=7.385
+ $Y=1.765 $X2=0 $Y2=0
cc_742 N_A_1444_320#_c_1104_n N_A_1272_128#_c_1197_n 0.00126277f $X=7.385
+ $Y=1.765 $X2=0 $Y2=0
cc_743 N_A_1444_320#_c_1105_n N_A_1272_128#_c_1197_n 0.0218861f $X=8.355 $Y=1.69
+ $X2=0 $Y2=0
cc_744 N_A_1444_320#_M1037_g N_A_1272_128#_c_1198_n 0.00361072f $X=7.405 $Y=0.85
+ $X2=0 $Y2=0
cc_745 N_A_1444_320#_c_1103_n N_A_1272_128#_c_1198_n 0.0261814f $X=7.385
+ $Y=1.765 $X2=0 $Y2=0
cc_746 N_A_1444_320#_c_1101_n N_VPWR_M1017_d 0.00235715f $X=8.745 $Y=1.685 $X2=0
+ $Y2=0
cc_747 N_A_1444_320#_M1036_g N_VPWR_c_1418_n 0.0124921f $X=7.295 $Y=2.69 $X2=0
+ $Y2=0
cc_748 N_A_1444_320#_c_1098_n N_VPWR_c_1418_n 0.00112295f $X=7.385 $Y=2.27 $X2=0
+ $Y2=0
cc_749 N_A_1444_320#_c_1103_n N_VPWR_c_1418_n 0.00998092f $X=7.385 $Y=1.765
+ $X2=0 $Y2=0
cc_750 N_A_1444_320#_c_1100_n N_VPWR_c_1419_n 0.0638102f $X=8.325 $Y=2.69 $X2=0
+ $Y2=0
cc_751 N_A_1444_320#_c_1101_n N_VPWR_c_1419_n 0.0238243f $X=8.745 $Y=1.685 $X2=0
+ $Y2=0
cc_752 N_A_1444_320#_M1036_g N_VPWR_c_1430_n 0.00444095f $X=7.295 $Y=2.69 $X2=0
+ $Y2=0
cc_753 N_A_1444_320#_c_1100_n N_VPWR_c_1431_n 0.00656052f $X=8.325 $Y=2.69 $X2=0
+ $Y2=0
cc_754 N_A_1444_320#_M1036_g N_VPWR_c_1413_n 0.00442501f $X=7.295 $Y=2.69 $X2=0
+ $Y2=0
cc_755 N_A_1444_320#_c_1100_n N_VPWR_c_1413_n 0.00908564f $X=8.325 $Y=2.69 $X2=0
+ $Y2=0
cc_756 N_A_1444_320#_c_1101_n Q_N 0.00873276f $X=8.745 $Y=1.685 $X2=0 $Y2=0
cc_757 N_A_1444_320#_c_1094_n Q_N 0.0391181f $X=8.885 $Y=1.6 $X2=0 $Y2=0
cc_758 N_A_1444_320#_c_1093_n N_VGND_M1010_s 0.00507763f $X=8.745 $Y=0.945 $X2=0
+ $Y2=0
cc_759 N_A_1444_320#_c_1094_n N_VGND_M1010_s 2.18744e-19 $X=8.885 $Y=1.6 $X2=0
+ $Y2=0
cc_760 N_A_1444_320#_M1037_g N_VGND_c_1661_n 0.011788f $X=7.405 $Y=0.85 $X2=0
+ $Y2=0
cc_761 N_A_1444_320#_c_1093_n N_VGND_c_1661_n 0.00688436f $X=8.745 $Y=0.945
+ $X2=0 $Y2=0
cc_762 N_A_1444_320#_c_1093_n N_VGND_c_1662_n 0.021825f $X=8.745 $Y=0.945 $X2=0
+ $Y2=0
cc_763 N_A_1444_320#_M1037_g N_VGND_c_1667_n 0.00338717f $X=7.405 $Y=0.85 $X2=0
+ $Y2=0
cc_764 N_A_1444_320#_M1037_g N_VGND_c_1682_n 0.00390857f $X=7.405 $Y=0.85 $X2=0
+ $Y2=0
cc_765 N_A_1444_320#_c_1093_n N_VGND_c_1682_n 0.0198821f $X=8.745 $Y=0.945 $X2=0
+ $Y2=0
cc_766 N_A_1272_128#_M1014_g N_A_2028_367#_M1018_g 0.0127981f $X=10.48 $Y=2.155
+ $X2=0 $Y2=0
cc_767 N_A_1272_128#_M1022_g N_A_2028_367#_c_1351_n 0.00470548f $X=9.575 $Y=0.67
+ $X2=0 $Y2=0
cc_768 N_A_1272_128#_c_1189_n N_A_2028_367#_c_1351_n 0.010439f $X=10.45 $Y=1.35
+ $X2=0 $Y2=0
cc_769 N_A_1272_128#_M1004_g N_A_2028_367#_c_1351_n 0.00890635f $X=10.54
+ $Y=0.555 $X2=0 $Y2=0
cc_770 N_A_1272_128#_c_1194_n N_A_2028_367#_c_1351_n 0.00775873f $X=10.54
+ $Y=0.98 $X2=0 $Y2=0
cc_771 N_A_1272_128#_M1014_g N_A_2028_367#_c_1352_n 0.0156826f $X=10.48 $Y=2.155
+ $X2=0 $Y2=0
cc_772 N_A_1272_128#_c_1189_n N_A_2028_367#_c_1353_n 0.00233283f $X=10.45
+ $Y=1.35 $X2=0 $Y2=0
cc_773 N_A_1272_128#_M1014_g N_A_2028_367#_c_1353_n 0.00489928f $X=10.48
+ $Y=2.155 $X2=0 $Y2=0
cc_774 N_A_1272_128#_c_1194_n N_A_2028_367#_c_1353_n 0.00316245f $X=10.54
+ $Y=0.98 $X2=0 $Y2=0
cc_775 N_A_1272_128#_c_1195_n N_A_2028_367#_c_1353_n 0.0024322f $X=10.465
+ $Y=1.425 $X2=0 $Y2=0
cc_776 N_A_1272_128#_c_1189_n N_A_2028_367#_c_1354_n 0.00299317f $X=10.45
+ $Y=1.35 $X2=0 $Y2=0
cc_777 N_A_1272_128#_c_1195_n N_A_2028_367#_c_1354_n 0.0178725f $X=10.465
+ $Y=1.425 $X2=0 $Y2=0
cc_778 N_A_1272_128#_M1023_g N_A_2028_367#_c_1355_n 0.00197723f $X=9.495 $Y=2.27
+ $X2=0 $Y2=0
cc_779 N_A_1272_128#_M1022_g N_A_2028_367#_c_1355_n 9.85611e-19 $X=9.575 $Y=0.67
+ $X2=0 $Y2=0
cc_780 N_A_1272_128#_c_1188_n N_A_2028_367#_c_1355_n 0.0165991f $X=10.375
+ $Y=1.425 $X2=0 $Y2=0
cc_781 N_A_1272_128#_c_1189_n N_A_2028_367#_c_1355_n 0.00162718f $X=10.45
+ $Y=1.35 $X2=0 $Y2=0
cc_782 N_A_1272_128#_M1014_g N_A_2028_367#_c_1355_n 0.00656374f $X=10.48
+ $Y=2.155 $X2=0 $Y2=0
cc_783 N_A_1272_128#_c_1195_n N_A_2028_367#_c_1355_n 0.00162434f $X=10.465
+ $Y=1.425 $X2=0 $Y2=0
cc_784 N_A_1272_128#_c_1189_n N_A_2028_367#_c_1356_n 0.00368094f $X=10.45
+ $Y=1.35 $X2=0 $Y2=0
cc_785 N_A_1272_128#_M1004_g N_A_2028_367#_c_1356_n 0.0152494f $X=10.54 $Y=0.555
+ $X2=0 $Y2=0
cc_786 N_A_1272_128#_c_1211_n N_VPWR_c_1418_n 0.00698907f $X=6.625 $Y=2.205
+ $X2=0 $Y2=0
cc_787 N_A_1272_128#_M1017_g N_VPWR_c_1419_n 0.0107062f $X=8.54 $Y=2.69 $X2=0
+ $Y2=0
cc_788 N_A_1272_128#_c_1183_n N_VPWR_c_1419_n 7.69258e-19 $X=8.99 $Y=1.425 $X2=0
+ $Y2=0
cc_789 N_A_1272_128#_M1009_g N_VPWR_c_1419_n 0.0146528f $X=9.065 $Y=2.27 $X2=0
+ $Y2=0
cc_790 N_A_1272_128#_M1023_g N_VPWR_c_1419_n 7.22232e-19 $X=9.495 $Y=2.27 $X2=0
+ $Y2=0
cc_791 N_A_1272_128#_M1023_g N_VPWR_c_1420_n 0.00761725f $X=9.495 $Y=2.27 $X2=0
+ $Y2=0
cc_792 N_A_1272_128#_c_1188_n N_VPWR_c_1420_n 0.00631861f $X=10.375 $Y=1.425
+ $X2=0 $Y2=0
cc_793 N_A_1272_128#_M1014_g N_VPWR_c_1420_n 0.00499281f $X=10.48 $Y=2.155 $X2=0
+ $Y2=0
cc_794 N_A_1272_128#_M1014_g N_VPWR_c_1421_n 0.00573215f $X=10.48 $Y=2.155 $X2=0
+ $Y2=0
cc_795 N_A_1272_128#_M1009_g N_VPWR_c_1424_n 0.00444095f $X=9.065 $Y=2.27 $X2=0
+ $Y2=0
cc_796 N_A_1272_128#_M1023_g N_VPWR_c_1424_n 0.00500904f $X=9.495 $Y=2.27 $X2=0
+ $Y2=0
cc_797 N_A_1272_128#_c_1211_n N_VPWR_c_1430_n 0.0112394f $X=6.625 $Y=2.205 $X2=0
+ $Y2=0
cc_798 N_A_1272_128#_M1017_g N_VPWR_c_1431_n 0.00511894f $X=8.54 $Y=2.69 $X2=0
+ $Y2=0
cc_799 N_A_1272_128#_M1014_g N_VPWR_c_1432_n 0.00312414f $X=10.48 $Y=2.155 $X2=0
+ $Y2=0
cc_800 N_A_1272_128#_M1017_g N_VPWR_c_1413_n 0.00526787f $X=8.54 $Y=2.69 $X2=0
+ $Y2=0
cc_801 N_A_1272_128#_M1009_g N_VPWR_c_1413_n 0.00442501f $X=9.065 $Y=2.27 $X2=0
+ $Y2=0
cc_802 N_A_1272_128#_M1023_g N_VPWR_c_1413_n 0.00526787f $X=9.495 $Y=2.27 $X2=0
+ $Y2=0
cc_803 N_A_1272_128#_M1014_g N_VPWR_c_1413_n 0.00410284f $X=10.48 $Y=2.155 $X2=0
+ $Y2=0
cc_804 N_A_1272_128#_c_1211_n N_VPWR_c_1413_n 0.0112734f $X=6.625 $Y=2.205 $X2=0
+ $Y2=0
cc_805 N_A_1272_128#_M1009_g Q_N 0.00195544f $X=9.065 $Y=2.27 $X2=0 $Y2=0
cc_806 N_A_1272_128#_M1010_g Q_N 0.00861353f $X=9.145 $Y=0.67 $X2=0 $Y2=0
cc_807 N_A_1272_128#_c_1186_n Q_N 0.00778231f $X=9.42 $Y=1.425 $X2=0 $Y2=0
cc_808 N_A_1272_128#_M1023_g Q_N 0.021036f $X=9.495 $Y=2.27 $X2=0 $Y2=0
cc_809 N_A_1272_128#_M1022_g Q_N 0.0042171f $X=9.575 $Y=0.67 $X2=0 $Y2=0
cc_810 N_A_1272_128#_c_1192_n Q_N 0.00243059f $X=9.105 $Y=1.425 $X2=0 $Y2=0
cc_811 N_A_1272_128#_c_1193_n Q_N 0.00489593f $X=9.535 $Y=1.425 $X2=0 $Y2=0
cc_812 N_A_1272_128#_c_1182_n N_VGND_c_1661_n 0.00208759f $X=8.195 $Y=1.17 $X2=0
+ $Y2=0
cc_813 N_A_1272_128#_c_1196_n N_VGND_c_1661_n 0.010409f $X=6.735 $Y=0.905 $X2=0
+ $Y2=0
cc_814 N_A_1272_128#_c_1197_n N_VGND_c_1661_n 0.0177658f $X=8.4 $Y=1.335 $X2=0
+ $Y2=0
cc_815 N_A_1272_128#_c_1182_n N_VGND_c_1662_n 0.00369302f $X=8.195 $Y=1.17 $X2=0
+ $Y2=0
cc_816 N_A_1272_128#_c_1183_n N_VGND_c_1662_n 7.17904e-19 $X=8.99 $Y=1.425 $X2=0
+ $Y2=0
cc_817 N_A_1272_128#_M1010_g N_VGND_c_1662_n 0.0115853f $X=9.145 $Y=0.67 $X2=0
+ $Y2=0
cc_818 N_A_1272_128#_M1022_g N_VGND_c_1662_n 5.38127e-19 $X=9.575 $Y=0.67 $X2=0
+ $Y2=0
cc_819 N_A_1272_128#_M1010_g N_VGND_c_1663_n 6.77346e-19 $X=9.145 $Y=0.67 $X2=0
+ $Y2=0
cc_820 N_A_1272_128#_M1022_g N_VGND_c_1663_n 0.0177674f $X=9.575 $Y=0.67 $X2=0
+ $Y2=0
cc_821 N_A_1272_128#_c_1188_n N_VGND_c_1663_n 0.00609477f $X=10.375 $Y=1.425
+ $X2=0 $Y2=0
cc_822 N_A_1272_128#_M1004_g N_VGND_c_1663_n 0.00482158f $X=10.54 $Y=0.555 $X2=0
+ $Y2=0
cc_823 N_A_1272_128#_c_1194_n N_VGND_c_1663_n 8.71609e-19 $X=10.54 $Y=0.98 $X2=0
+ $Y2=0
cc_824 N_A_1272_128#_c_1189_n N_VGND_c_1664_n 5.76908e-19 $X=10.45 $Y=1.35 $X2=0
+ $Y2=0
cc_825 N_A_1272_128#_M1004_g N_VGND_c_1664_n 0.00669066f $X=10.54 $Y=0.555 $X2=0
+ $Y2=0
cc_826 N_A_1272_128#_c_1196_n N_VGND_c_1667_n 0.00404505f $X=6.735 $Y=0.905
+ $X2=0 $Y2=0
cc_827 N_A_1272_128#_c_1182_n N_VGND_c_1672_n 0.00407505f $X=8.195 $Y=1.17 $X2=0
+ $Y2=0
cc_828 N_A_1272_128#_M1010_g N_VGND_c_1673_n 0.00473366f $X=9.145 $Y=0.67 $X2=0
+ $Y2=0
cc_829 N_A_1272_128#_M1022_g N_VGND_c_1673_n 0.00473366f $X=9.575 $Y=0.67 $X2=0
+ $Y2=0
cc_830 N_A_1272_128#_M1004_g N_VGND_c_1674_n 0.0045478f $X=10.54 $Y=0.555 $X2=0
+ $Y2=0
cc_831 N_A_1272_128#_c_1182_n N_VGND_c_1682_n 0.00465306f $X=8.195 $Y=1.17 $X2=0
+ $Y2=0
cc_832 N_A_1272_128#_M1010_g N_VGND_c_1682_n 0.00755886f $X=9.145 $Y=0.67 $X2=0
+ $Y2=0
cc_833 N_A_1272_128#_M1022_g N_VGND_c_1682_n 0.00827881f $X=9.575 $Y=0.67 $X2=0
+ $Y2=0
cc_834 N_A_1272_128#_M1004_g N_VGND_c_1682_n 0.00895354f $X=10.54 $Y=0.555 $X2=0
+ $Y2=0
cc_835 N_A_1272_128#_c_1196_n N_VGND_c_1682_n 0.00525146f $X=6.735 $Y=0.905
+ $X2=0 $Y2=0
cc_836 N_A_2028_367#_c_1352_n N_VPWR_c_1420_n 0.0532557f $X=10.265 $Y=1.98 $X2=0
+ $Y2=0
cc_837 N_A_2028_367#_c_1355_n N_VPWR_c_1420_n 3.31042e-19 $X=10.307 $Y=1.46
+ $X2=0 $Y2=0
cc_838 N_A_2028_367#_M1018_g N_VPWR_c_1421_n 0.00810646f $X=11.065 $Y=2.465
+ $X2=0 $Y2=0
cc_839 N_A_2028_367#_c_1352_n N_VPWR_c_1421_n 0.0260164f $X=10.265 $Y=1.98 $X2=0
+ $Y2=0
cc_840 N_A_2028_367#_c_1353_n N_VPWR_c_1421_n 0.0280703f $X=10.93 $Y=1.46 $X2=0
+ $Y2=0
cc_841 N_A_2028_367#_c_1354_n N_VPWR_c_1421_n 0.00435887f $X=10.93 $Y=1.46 $X2=0
+ $Y2=0
cc_842 N_A_2028_367#_M1026_g N_VPWR_c_1423_n 0.00776549f $X=11.495 $Y=2.465
+ $X2=0 $Y2=0
cc_843 N_A_2028_367#_M1018_g N_VPWR_c_1433_n 0.00585385f $X=11.065 $Y=2.465
+ $X2=0 $Y2=0
cc_844 N_A_2028_367#_M1026_g N_VPWR_c_1433_n 0.00585385f $X=11.495 $Y=2.465
+ $X2=0 $Y2=0
cc_845 N_A_2028_367#_M1018_g N_VPWR_c_1413_n 0.0118904f $X=11.065 $Y=2.465 $X2=0
+ $Y2=0
cc_846 N_A_2028_367#_M1026_g N_VPWR_c_1413_n 0.0114822f $X=11.495 $Y=2.465 $X2=0
+ $Y2=0
cc_847 N_A_2028_367#_c_1352_n N_VPWR_c_1413_n 0.0118013f $X=10.265 $Y=1.98 $X2=0
+ $Y2=0
cc_848 N_A_2028_367#_c_1351_n Q_N 0.00576235f $X=10.325 $Y=0.55 $X2=0 $Y2=0
cc_849 N_A_2028_367#_c_1355_n Q_N 0.00904289f $X=10.307 $Y=1.46 $X2=0 $Y2=0
cc_850 N_A_2028_367#_M1018_g Q 0.00564634f $X=11.065 $Y=2.465 $X2=0 $Y2=0
cc_851 N_A_2028_367#_c_1347_n Q 0.0159372f $X=11.42 $Y=1.55 $X2=0 $Y2=0
cc_852 N_A_2028_367#_M1030_g Q 0.00811794f $X=11.495 $Y=0.765 $X2=0 $Y2=0
cc_853 N_A_2028_367#_M1026_g Q 0.00590937f $X=11.495 $Y=2.465 $X2=0 $Y2=0
cc_854 N_A_2028_367#_c_1353_n Q 0.0261708f $X=10.93 $Y=1.46 $X2=0 $Y2=0
cc_855 N_A_2028_367#_c_1356_n Q 0.0050075f $X=10.952 $Y=1.295 $X2=0 $Y2=0
cc_856 N_A_2028_367#_c_1351_n N_VGND_c_1663_n 0.0608331f $X=10.325 $Y=0.55 $X2=0
+ $Y2=0
cc_857 N_A_2028_367#_M1030_g N_VGND_c_1664_n 5.9294e-19 $X=11.495 $Y=0.765 $X2=0
+ $Y2=0
cc_858 N_A_2028_367#_c_1351_n N_VGND_c_1664_n 0.0432248f $X=10.325 $Y=0.55 $X2=0
+ $Y2=0
cc_859 N_A_2028_367#_c_1353_n N_VGND_c_1664_n 0.0270253f $X=10.93 $Y=1.46 $X2=0
+ $Y2=0
cc_860 N_A_2028_367#_c_1354_n N_VGND_c_1664_n 0.00506784f $X=10.93 $Y=1.46 $X2=0
+ $Y2=0
cc_861 N_A_2028_367#_c_1356_n N_VGND_c_1664_n 0.0187402f $X=10.952 $Y=1.295
+ $X2=0 $Y2=0
cc_862 N_A_2028_367#_M1030_g N_VGND_c_1666_n 0.00737423f $X=11.495 $Y=0.765
+ $X2=0 $Y2=0
cc_863 N_A_2028_367#_c_1351_n N_VGND_c_1674_n 0.0127991f $X=10.325 $Y=0.55 $X2=0
+ $Y2=0
cc_864 N_A_2028_367#_M1030_g N_VGND_c_1675_n 0.00482246f $X=11.495 $Y=0.765
+ $X2=0 $Y2=0
cc_865 N_A_2028_367#_c_1356_n N_VGND_c_1675_n 0.00400407f $X=10.952 $Y=1.295
+ $X2=0 $Y2=0
cc_866 N_A_2028_367#_M1030_g N_VGND_c_1682_n 0.00964708f $X=11.495 $Y=0.765
+ $X2=0 $Y2=0
cc_867 N_A_2028_367#_c_1351_n N_VGND_c_1682_n 0.01299f $X=10.325 $Y=0.55 $X2=0
+ $Y2=0
cc_868 N_A_2028_367#_c_1356_n N_VGND_c_1682_n 0.00774504f $X=10.952 $Y=1.295
+ $X2=0 $Y2=0
cc_869 N_VPWR_M1016_d N_A_308_463#_c_1573_n 0.00624472f $X=1.955 $Y=2.315 $X2=0
+ $Y2=0
cc_870 N_VPWR_c_1415_n N_A_308_463#_c_1573_n 0.0235704f $X=2.165 $Y=2.75 $X2=0
+ $Y2=0
cc_871 N_VPWR_c_1413_n N_A_308_463#_c_1573_n 0.0143212f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_872 N_VPWR_c_1427_n N_A_308_463#_c_1570_n 0.00401414f $X=1.99 $Y=3.33 $X2=0
+ $Y2=0
cc_873 N_VPWR_c_1413_n N_A_308_463#_c_1570_n 0.00526109f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_874 N_VPWR_c_1428_n N_A_308_463#_c_1571_n 0.0159855f $X=4.36 $Y=3.33 $X2=0
+ $Y2=0
cc_875 N_VPWR_c_1413_n N_A_308_463#_c_1571_n 0.0214334f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_876 N_VPWR_c_1419_n Q_N 0.0358568f $X=8.85 $Y=2.025 $X2=0 $Y2=0
cc_877 N_VPWR_c_1420_n Q_N 0.0485453f $X=9.71 $Y=1.785 $X2=0 $Y2=0
cc_878 N_VPWR_c_1424_n Q_N 0.00917475f $X=9.625 $Y=3.33 $X2=0 $Y2=0
cc_879 N_VPWR_c_1413_n Q_N 0.00914479f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_880 N_VPWR_c_1413_n N_Q_M1018_s 0.0041489f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_881 N_VPWR_c_1421_n Q 0.00125019f $X=10.695 $Y=1.98 $X2=0 $Y2=0
cc_882 N_VPWR_c_1423_n Q 0.0015231f $X=11.71 $Y=1.98 $X2=0 $Y2=0
cc_883 N_VPWR_c_1433_n Q 0.0136943f $X=11.58 $Y=3.33 $X2=0 $Y2=0
cc_884 N_VPWR_c_1413_n Q 0.00866972f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_885 N_VPWR_c_1420_n N_VGND_c_1663_n 0.010631f $X=9.71 $Y=1.785 $X2=0 $Y2=0
cc_886 N_VPWR_c_1423_n N_VGND_c_1666_n 0.0112202f $X=11.71 $Y=1.98 $X2=0 $Y2=0
cc_887 Q_N N_VGND_c_1663_n 0.0328441f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_888 N_Q_N_c_1638_p N_VGND_c_1673_n 0.0124525f $X=9.36 $Y=0.42 $X2=0 $Y2=0
cc_889 Q_N N_VGND_c_1682_n 0.00254576f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_890 N_Q_N_c_1638_p N_VGND_c_1682_n 0.00730901f $X=9.36 $Y=0.42 $X2=0 $Y2=0
cc_891 Q N_VGND_c_1664_n 0.0303292f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_892 Q N_VGND_c_1666_n 0.00224457f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_893 Q N_VGND_c_1675_n 0.0105866f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_894 Q N_VGND_c_1682_n 0.00830966f $X=11.195 $Y=0.47 $X2=0 $Y2=0
