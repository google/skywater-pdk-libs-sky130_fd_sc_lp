* File: sky130_fd_sc_lp__and2_m.spice
* Created: Fri Aug 28 10:04:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and2_m.pex.spice"
.subckt sky130_fd_sc_lp__and2_m  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_117_141# N_A_M1004_g N_A_34_141#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g A_117_141# VNB NSHORT L=0.15 W=0.42 AD=0.08925
+ AS=0.0441 PD=0.845 PS=0.63 NRD=41.424 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_34_141#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.08925 PD=1.37 PS=0.845 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_34_141#_M1003_d N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1512 PD=0.7 PS=1.56 NRD=0 NRS=44.5417 M=1 R=2.8 SA=75000.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_A_34_141#_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_34_141#_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__and2_m.pxi.spice"
*
.ends
*
*
