* File: sky130_fd_sc_lp__dfsbp_1.pex.spice
* Created: Fri Aug 28 10:22:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFSBP_1%CLK 2 5 8 10 11 12 13 14 21 23 38
r34 38 39 1.79674 $w=3.83e-07 $l=5.5e-08 $layer=LI1_cond $X=0.277 $Y=2.035
+ $X2=0.277 $Y2=2.09
r35 21 23 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.387 $Y=1.475
+ $X2=0.387 $Y2=1.31
r36 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.475 $X2=0.385 $Y2=1.475
r37 13 38 0.449004 $w=3.83e-07 $l=1.5e-08 $layer=LI1_cond $X=0.277 $Y=2.02
+ $X2=0.277 $Y2=2.035
r38 13 24 3.6519 $w=3.83e-07 $l=1.22e-07 $layer=LI1_cond $X=0.277 $Y=2.02
+ $X2=0.277 $Y2=1.898
r39 13 14 10.0212 $w=3.43e-07 $l=3e-07 $layer=LI1_cond $X=0.257 $Y=2.105
+ $X2=0.257 $Y2=2.405
r40 13 39 0.501062 $w=3.43e-07 $l=1.5e-08 $layer=LI1_cond $X=0.257 $Y=2.105
+ $X2=0.257 $Y2=2.09
r41 12 24 6.97452 $w=3.83e-07 $l=2.33e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.898
r42 12 22 5.68738 $w=3.83e-07 $l=1.9e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.475
r43 11 22 5.38805 $w=3.83e-07 $l=1.8e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.475
r44 8 10 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.48 $Y=2.6 $X2=0.48
+ $Y2=1.98
r45 5 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.48 $Y=0.99 $X2=0.48
+ $Y2=1.31
r46 2 10 46.5995 $w=3.35e-07 $l=1.67e-07 $layer=POLY_cond $X=0.387 $Y=1.813
+ $X2=0.387 $Y2=1.98
r47 1 21 0.344503 $w=3.35e-07 $l=2e-09 $layer=POLY_cond $X=0.387 $Y=1.477
+ $X2=0.387 $Y2=1.475
r48 1 2 57.8765 $w=3.35e-07 $l=3.36e-07 $layer=POLY_cond $X=0.387 $Y=1.477
+ $X2=0.387 $Y2=1.813
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_111_156# 1 2 7 9 11 12 14 17 19 20 23 27
+ 31 35 38 39 42 45 48 51 52 53 55 58 59 61 64 65 66 68 69 70 71 74 77 78 79 82
+ 83 85 88
c265 88 0 1.50513e-19 $X=6.67 $Y=1.5
c266 77 0 1.81645e-19 $X=1.15 $Y=2.94
c267 71 0 2.18694e-19 $X=6.635 $Y=1.505
c268 69 0 1.79345e-19 $X=6.27 $Y=1.33
c269 59 0 1.80116e-19 $X=3.495 $Y=1.66
c270 52 0 4.25888e-20 $X=3.325 $Y=0.385
c271 38 0 5.22705e-20 $X=6.67 $Y=1.84
c272 31 0 4.22624e-20 $X=6.76 $Y=2.665
c273 27 0 1.77516e-19 $X=6.58 $Y=0.965
c274 23 0 2.19324e-19 $X=3.36 $Y=2.875
r275 83 95 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.72 $Y=1.29
+ $X2=1.585 $Y2=1.29
r276 82 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.29 $X2=1.72 $Y2=1.29
r277 79 82 10.8065 $w=1.93e-07 $l=1.9e-07 $layer=LI1_cond $X=1.732 $Y=1.1
+ $X2=1.732 $Y2=1.29
r278 77 93 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.15 $Y=2.94
+ $X2=1.15 $Y2=3.15
r279 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=2.94 $X2=1.15 $Y2=2.94
r280 74 76 9.66615 $w=6.5e-07 $l=6.03838e-07 $layer=LI1_cond $X=0.957 $Y=2.425
+ $X2=1.15 $Y2=2.94
r281 71 88 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.67
+ $Y=1.5 $X2=6.67 $Y2=1.5
r282 69 71 21.1264 $w=2.17e-07 $l=3.86846e-07 $layer=LI1_cond $X=6.27 $Y=1.33
+ $X2=6.635 $Y2=1.375
r283 69 70 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=6.27 $Y=1.33
+ $X2=4.985 $Y2=1.33
r284 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.9 $Y=1.245
+ $X2=4.985 $Y2=1.33
r285 67 68 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.9 $Y=0.775
+ $X2=4.9 $Y2=1.245
r286 65 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=0.69
+ $X2=4.9 $Y2=0.775
r287 65 66 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.815 $Y=0.69
+ $X2=4.265 $Y2=0.69
r288 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.18 $Y=0.775
+ $X2=4.265 $Y2=0.69
r289 63 64 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.18 $Y=0.775
+ $X2=4.18 $Y2=1.075
r290 62 85 1.79375 $w=1.7e-07 $l=3.29773e-07 $layer=LI1_cond $X=3.615 $Y=1.16
+ $X2=3.325 $Y2=1.075
r291 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.095 $Y=1.16
+ $X2=4.18 $Y2=1.075
r292 61 62 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.095 $Y=1.16
+ $X2=3.615 $Y2=1.16
r293 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.495
+ $Y=1.66 $X2=3.495 $Y2=1.66
r294 56 85 4.65272 $w=1.92e-07 $l=2.53109e-07 $layer=LI1_cond $X=3.507 $Y=1.245
+ $X2=3.325 $Y2=1.075
r295 56 58 22.2448 $w=2.13e-07 $l=4.15e-07 $layer=LI1_cond $X=3.507 $Y=1.245
+ $X2=3.507 $Y2=1.66
r296 55 85 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.075
+ $X2=3.325 $Y2=1.075
r297 54 55 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.41 $Y=0.47
+ $X2=3.41 $Y2=1.075
r298 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.325 $Y=0.385
+ $X2=3.41 $Y2=0.47
r299 52 53 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.325 $Y=0.385
+ $X2=2.315 $Y2=0.385
r300 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.23 $Y=0.47
+ $X2=2.315 $Y2=0.385
r301 50 51 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.23 $Y=0.47
+ $X2=2.23 $Y2=1.015
r302 49 79 1.54022 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.83 $Y=1.1
+ $X2=1.732 $Y2=1.1
r303 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.145 $Y=1.1
+ $X2=2.23 $Y2=1.015
r304 48 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.145 $Y=1.1
+ $X2=1.83 $Y2=1.1
r305 47 78 2.45049 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.9 $Y=1.37 $X2=0.77
+ $Y2=1.37
r306 47 82 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.9 $Y=1.37
+ $X2=1.635 $Y2=1.37
r307 45 74 9.49849 $w=6.5e-07 $l=2.87913e-07 $layer=LI1_cond $X=0.74 $Y=2.26
+ $X2=0.957 $Y2=2.425
r308 44 78 3.98977 $w=2.3e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.74 $Y=1.455
+ $X2=0.77 $Y2=1.37
r309 44 45 44.6409 $w=1.98e-07 $l=8.05e-07 $layer=LI1_cond $X=0.74 $Y=1.455
+ $X2=0.74 $Y2=2.26
r310 40 78 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=1.285
+ $X2=0.77 $Y2=1.37
r311 40 42 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.77 $Y=1.285
+ $X2=0.77 $Y2=0.995
r312 38 88 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.67 $Y=1.84
+ $X2=6.67 $Y2=1.5
r313 38 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.67 $Y=1.84
+ $X2=6.67 $Y2=2.005
r314 37 88 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.67 $Y=1.335
+ $X2=6.67 $Y2=1.5
r315 34 59 35.3689 $w=4.45e-07 $l=2.83e-07 $layer=POLY_cond $X=3.437 $Y=1.943
+ $X2=3.437 $Y2=1.66
r316 34 35 45.5004 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=3.437 $Y=1.943
+ $X2=3.437 $Y2=2.165
r317 33 59 6.87381 $w=4.45e-07 $l=5.5e-08 $layer=POLY_cond $X=3.437 $Y=1.605
+ $X2=3.437 $Y2=1.66
r318 31 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.76 $Y=2.665
+ $X2=6.76 $Y2=2.005
r319 27 37 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.58 $Y=0.965
+ $X2=6.58 $Y2=1.335
r320 23 35 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.36 $Y=2.875
+ $X2=3.36 $Y2=2.165
r321 19 33 131.942 $w=8.2e-08 $l=2.56776e-07 $layer=POLY_cond $X=3.215 $Y=1.53
+ $X2=3.437 $Y2=1.605
r322 19 20 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.215 $Y=1.53
+ $X2=2.9 $Y2=1.53
r323 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.825 $Y=1.455
+ $X2=2.9 $Y2=1.53
r324 15 17 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.825 $Y=1.455
+ $X2=2.825 $Y2=0.805
r325 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.815 $Y=3.075
+ $X2=1.815 $Y2=2.645
r326 9 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.125
+ $X2=1.585 $Y2=1.29
r327 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.585 $Y=1.125
+ $X2=1.585 $Y2=0.805
r328 8 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.315 $Y=3.15
+ $X2=1.15 $Y2=3.15
r329 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.74 $Y=3.15
+ $X2=1.815 $Y2=3.075
r330 7 8 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.74 $Y=3.15
+ $X2=1.315 $Y2=3.15
r331 2 74 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=2.28 $X2=0.695 $Y2=2.425
r332 1 42 182 $w=1.7e-07 $l=2.91419e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.78 $X2=0.735 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%D 3 7 9 10 11 17 19 22 23
c57 17 0 6.00859e-20 $X=2.26 $Y=1.44
r58 23 34 4.23719 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=2.34
+ $X2=2.275 $Y2=2.175
r59 22 25 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=2.472 $Y=2.34
+ $X2=2.472 $Y2=2.505
r60 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.465
+ $Y=2.34 $X2=2.465 $Y2=2.34
r61 16 19 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.26 $Y=1.44
+ $X2=2.395 $Y2=1.44
r62 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.44 $X2=2.26 $Y2=1.44
r63 11 23 1.41355 $w=5.48e-07 $l=6.5e-08 $layer=LI1_cond $X=2.275 $Y=2.405
+ $X2=2.275 $Y2=2.34
r64 10 34 3.79628 $w=4.23e-07 $l=1.4e-07 $layer=LI1_cond $X=2.212 $Y=2.035
+ $X2=2.212 $Y2=2.175
r65 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.212 $Y=1.665
+ $X2=2.212 $Y2=2.035
r66 9 17 6.10117 $w=4.23e-07 $l=2.25e-07 $layer=LI1_cond $X=2.212 $Y=1.665
+ $X2=2.212 $Y2=1.44
r67 7 25 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.5 $Y=2.875 $X2=2.5
+ $Y2=2.505
r68 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.275
+ $X2=2.395 $Y2=1.44
r69 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.395 $Y=1.275 $X2=2.395
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_708_93# 1 2 7 9 10 12 13 14 15 16 21 24 27
+ 30 32 34 38 40 43 45
c103 40 0 5.27659e-20 $X=4.365 $Y=2.34
c104 7 0 4.25888e-20 $X=3.615 $Y=1.135
r105 43 45 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.13 $Y=1.665
+ $X2=4.13 $Y2=2.175
r106 38 46 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.22 $Y=2.34
+ $X2=4.22 $Y2=2.48
r107 38 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.22 $Y=2.34
+ $X2=4.22 $Y2=2.175
r108 37 40 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.22 $Y=2.34
+ $X2=4.365 $Y2=2.34
r109 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=2.34 $X2=4.22 $Y2=2.34
r110 32 34 35.2717 $w=3.28e-07 $l=1.01e-06 $layer=LI1_cond $X=4.45 $Y=2.85
+ $X2=5.46 $Y2=2.85
r111 28 30 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.54 $Y=1.415
+ $X2=4.54 $Y2=1.12
r112 27 32 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.365 $Y=2.685
+ $X2=4.45 $Y2=2.85
r113 26 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=2.505
+ $X2=4.365 $Y2=2.34
r114 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.365 $Y=2.505
+ $X2=4.365 $Y2=2.685
r115 24 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.065 $Y=1.5
+ $X2=4.065 $Y2=1.665
r116 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.065
+ $Y=1.5 $X2=4.065 $Y2=1.5
r117 21 28 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.445 $Y=1.5
+ $X2=4.54 $Y2=1.415
r118 21 23 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.445 $Y=1.5
+ $X2=4.065 $Y2=1.5
r119 17 24 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.065 $Y=1.285
+ $X2=4.065 $Y2=1.5
r120 15 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.055 $Y=2.48
+ $X2=4.22 $Y2=2.48
r121 15 16 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=4.055 $Y=2.48
+ $X2=3.795 $Y2=2.48
r122 13 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.9 $Y=1.21
+ $X2=4.065 $Y2=1.285
r123 13 14 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.9 $Y=1.21
+ $X2=3.69 $Y2=1.21
r124 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.72 $Y=2.555
+ $X2=3.795 $Y2=2.48
r125 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.72 $Y=2.555
+ $X2=3.72 $Y2=2.875
r126 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.615 $Y=1.135
+ $X2=3.69 $Y2=1.21
r127 7 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.615 $Y=1.135
+ $X2=3.615 $Y2=0.805
r128 2 34 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=5.32
+ $Y=2.665 $X2=5.46 $Y2=2.85
r129 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.845 $X2=4.53 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_580_119# 1 2 9 11 12 13 15 18 20 21 26 30
+ 33 36 39 41 44 45 46 47 49 50 56 57 60 61 64 65 68
c173 68 0 5.8525e-20 $X=6.13 $Y=2.015
c174 65 0 5.22705e-20 $X=5.845 $Y=1.805
c175 56 0 4.22624e-20 $X=6.13 $Y=1.85
c176 49 0 5.27152e-20 $X=4.76 $Y=2
c177 39 0 2.29862e-19 $X=3.145 $Y=2.885
c178 36 0 6.00859e-20 $X=3.145 $Y=2.485
c179 21 0 1.81116e-19 $X=5.705 $Y=1.55
c180 20 0 1.11656e-19 $X=5.965 $Y=1.55
c181 11 0 7.94915e-20 $X=5.17 $Y=2.48
r182 64 65 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.675 $Y=1.805
+ $X2=5.845 $Y2=1.805
r183 62 63 8.64167 $w=2.4e-07 $l=1.7e-07 $layer=LI1_cond $X=4.83 $Y=1.68
+ $X2=4.83 $Y2=1.85
r184 59 60 9.41323 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=3.087 $Y=1.415
+ $X2=3.087 $Y2=1.585
r185 57 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=1.85
+ $X2=6.13 $Y2=2.015
r186 56 65 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.13 $Y=1.85
+ $X2=5.845 $Y2=1.85
r187 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.13
+ $Y=1.85 $X2=6.13 $Y2=1.85
r188 53 62 2.75731 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.985 $Y=1.68
+ $X2=4.83 $Y2=1.68
r189 53 64 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.985 $Y=1.68
+ $X2=5.675 $Y2=1.68
r190 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.76 $Y=2
+ $X2=4.76 $Y2=2
r191 47 63 3.99923 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=1.935
+ $X2=4.83 $Y2=1.85
r192 47 49 2.41641 $w=3.08e-07 $l=6.5e-08 $layer=LI1_cond $X=4.83 $Y=1.935
+ $X2=4.83 $Y2=2
r193 45 63 2.75731 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.675 $Y=1.85
+ $X2=4.83 $Y2=1.85
r194 45 46 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.675 $Y=1.85
+ $X2=3.955 $Y2=1.85
r195 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.87 $Y=1.935
+ $X2=3.955 $Y2=1.85
r196 43 44 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.87 $Y=1.935
+ $X2=3.87 $Y2=2.485
r197 42 61 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.31 $Y=2.57
+ $X2=3.185 $Y2=2.57
r198 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.785 $Y=2.57
+ $X2=3.87 $Y2=2.485
r199 41 42 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.785 $Y=2.57
+ $X2=3.31 $Y2=2.57
r200 37 61 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=2.655
+ $X2=3.185 $Y2=2.57
r201 37 39 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=3.185 $Y=2.655
+ $X2=3.185 $Y2=2.885
r202 36 61 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.145 $Y=2.485
+ $X2=3.185 $Y2=2.57
r203 36 60 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=3.145 $Y=2.485
+ $X2=3.145 $Y2=1.585
r204 33 59 31.9524 $w=2.08e-07 $l=6.05e-07 $layer=LI1_cond $X=3.05 $Y=0.81
+ $X2=3.05 $Y2=1.415
r205 30 50 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=4.76 $Y=2.405
+ $X2=4.76 $Y2=2
r206 29 50 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.76 $Y=1.835
+ $X2=4.76 $Y2=2
r207 26 68 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=6.22 $Y=2.665
+ $X2=6.22 $Y2=2.015
r208 22 57 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=6.13 $Y=1.625
+ $X2=6.13 $Y2=1.85
r209 20 22 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.965 $Y=1.55
+ $X2=6.13 $Y2=1.625
r210 20 21 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.965 $Y=1.55
+ $X2=5.705 $Y2=1.55
r211 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.63 $Y=1.475
+ $X2=5.705 $Y2=1.55
r212 16 18 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.63 $Y=1.475
+ $X2=5.63 $Y2=0.945
r213 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.245 $Y=2.555
+ $X2=5.245 $Y2=2.875
r214 12 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.925 $Y=2.48
+ $X2=4.76 $Y2=2.405
r215 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.17 $Y=2.48
+ $X2=5.245 $Y2=2.555
r216 11 12 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=5.17 $Y=2.48
+ $X2=4.925 $Y2=2.48
r217 9 29 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.745 $Y=1.055
+ $X2=4.745 $Y2=1.835
r218 2 39 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=2.665 $X2=3.145 $Y2=2.885
r219 1 33 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.9
+ $Y=0.595 $X2=3.04 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%SET_B 3 6 9 13 17 21 24 25 26 28 29 31 35 36
+ 41 42 50
c127 41 0 2.60608e-19 $X=6.33 $Y=2.367
c128 36 0 1.79345e-19 $X=5.33 $Y=2.03
c129 35 0 5.8525e-20 $X=5.33 $Y=2.03
c130 17 0 1.283e-20 $X=8.57 $Y=0.565
c131 9 0 5.27152e-20 $X=5.675 $Y=2.875
r132 41 42 15.5227 $w=2.43e-07 $l=3.3e-07 $layer=LI1_cond $X=6.33 $Y=2.367 $X2=6
+ $Y2=2.367
r133 39 42 23.7544 $w=2.43e-07 $l=5.05e-07 $layer=LI1_cond $X=5.495 $Y=2.367
+ $X2=6 $Y2=2.367
r134 38 39 2.50173 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=5.33 $Y=2.367
+ $X2=5.495 $Y2=2.367
r135 36 44 17.2829 $w=2.51e-07 $l=9e-08 $layer=POLY_cond $X=5.33 $Y=2.03
+ $X2=5.24 $Y2=2.03
r136 35 38 11.7689 $w=3.28e-07 $l=3.37e-07 $layer=LI1_cond $X=5.33 $Y=2.03
+ $X2=5.33 $Y2=2.367
r137 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=2.03 $X2=5.33 $Y2=2.03
r138 32 50 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=8.27 $Y=1.88 $X2=8.57
+ $Y2=1.88
r139 32 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.27 $Y=1.88 $X2=8.18
+ $Y2=1.88
r140 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.27
+ $Y=1.88 $X2=8.27 $Y2=1.88
r141 29 31 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=7.68 $Y=1.88
+ $X2=8.27 $Y2=1.88
r142 27 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.595 $Y=2.045
+ $X2=7.68 $Y2=1.88
r143 27 28 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.595 $Y=2.045
+ $X2=7.595 $Y2=2.845
r144 25 28 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.51 $Y=2.96
+ $X2=7.595 $Y2=2.845
r145 25 26 50.6073 $w=2.28e-07 $l=1.01e-06 $layer=LI1_cond $X=7.51 $Y=2.96
+ $X2=6.5 $Y2=2.96
r146 24 26 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.415 $Y=2.845
+ $X2=6.5 $Y2=2.96
r147 23 41 7.11011 $w=2.45e-07 $l=1.5995e-07 $layer=LI1_cond $X=6.415 $Y=2.49
+ $X2=6.33 $Y2=2.367
r148 23 24 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.415 $Y=2.49
+ $X2=6.415 $Y2=2.845
r149 19 21 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.105 $Y=1.52
+ $X2=5.24 $Y2=1.52
r150 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.57 $Y=1.715
+ $X2=8.57 $Y2=1.88
r151 15 17 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=8.57 $Y=1.715
+ $X2=8.57 $Y2=0.565
r152 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.18 $Y=2.045
+ $X2=8.18 $Y2=1.88
r153 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.18 $Y=2.045
+ $X2=8.18 $Y2=2.455
r154 7 36 66.251 $w=2.51e-07 $l=4.19464e-07 $layer=POLY_cond $X=5.675 $Y=2.195
+ $X2=5.33 $Y2=2.03
r155 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.675 $Y=2.195
+ $X2=5.675 $Y2=2.875
r156 6 44 14.812 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.865
+ $X2=5.24 $Y2=2.03
r157 5 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.24 $Y=1.595
+ $X2=5.24 $Y2=1.52
r158 5 6 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.24 $Y=1.595
+ $X2=5.24 $Y2=1.865
r159 1 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.105 $Y=1.445
+ $X2=5.105 $Y2=1.52
r160 1 3 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=5.105 $Y=1.445
+ $X2=5.105 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_161_21# 1 2 8 9 11 15 19 21 26 29 31 34 36
+ 41 48 52 54 61
c145 41 0 1.81645e-19 $X=1.485 $Y=1.952
c146 34 0 8.90566e-20 $X=7.285 $Y=1.36
c147 29 0 4.55038e-20 $X=7.285 $Y=2.455
c148 26 0 8.41339e-20 $X=7.125 $Y=0.855
c149 15 0 1.71596e-19 $X=2.93 $Y=2.875
r150 50 52 15.6403 $w=2.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.625 $Y=2.09
+ $X2=1.625 $Y2=2.47
r151 46 48 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=1.335 $Y=0.515
+ $X2=1.335 $Y2=0.78
r152 44 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.98
+ $X2=1.35 $Y2=1.98
r153 44 58 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.185 $Y=1.98
+ $X2=1.06 $Y2=1.98
r154 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.185
+ $Y=1.98 $X2=1.185 $Y2=1.98
r155 41 50 6.81721 $w=2.75e-07 $l=1.97282e-07 $layer=LI1_cond $X=1.485 $Y=1.952
+ $X2=1.625 $Y2=2.09
r156 41 43 12.5721 $w=2.73e-07 $l=3e-07 $layer=LI1_cond $X=1.485 $Y=1.952
+ $X2=1.185 $Y2=1.952
r157 39 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=0.35
+ $X2=0.97 $Y2=0.515
r158 39 54 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.97 $Y=0.35
+ $X2=0.97 $Y2=0.18
r159 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=0.35 $X2=0.97 $Y2=0.35
r160 36 46 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=1.205 $Y=0.39
+ $X2=1.335 $Y2=0.515
r161 36 38 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=1.205 $Y=0.39
+ $X2=0.97 $Y2=0.39
r162 32 34 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.125 $Y=1.36
+ $X2=7.285 $Y2=1.36
r163 27 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.285 $Y=1.435
+ $X2=7.285 $Y2=1.36
r164 27 29 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=7.285 $Y=1.435
+ $X2=7.285 $Y2=2.455
r165 24 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.125 $Y=1.285
+ $X2=7.125 $Y2=1.36
r166 24 26 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.125 $Y=1.285
+ $X2=7.125 $Y2=0.855
r167 23 26 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.125 $Y=0.255
+ $X2=7.125 $Y2=0.855
r168 22 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.33 $Y=0.18
+ $X2=3.255 $Y2=0.18
r169 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.05 $Y=0.18
+ $X2=7.125 $Y2=0.255
r170 21 22 1907.49 $w=1.5e-07 $l=3.72e-06 $layer=POLY_cond $X=7.05 $Y=0.18
+ $X2=3.33 $Y2=0.18
r171 17 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=0.255
+ $X2=3.255 $Y2=0.18
r172 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.255 $Y=0.255
+ $X2=3.255 $Y2=0.805
r173 13 15 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.93 $Y=1.965
+ $X2=2.93 $Y2=2.875
r174 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.855 $Y=1.89
+ $X2=2.93 $Y2=1.965
r175 11 61 771.713 $w=1.5e-07 $l=1.505e-06 $layer=POLY_cond $X=2.855 $Y=1.89
+ $X2=1.35 $Y2=1.89
r176 10 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=0.18
+ $X2=0.97 $Y2=0.18
r177 9 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=0.18
+ $X2=3.255 $Y2=0.18
r178 9 10 1048.61 $w=1.5e-07 $l=2.045e-06 $layer=POLY_cond $X=3.18 $Y=0.18
+ $X2=1.135 $Y2=0.18
r179 8 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.815
+ $X2=1.06 $Y2=1.98
r180 8 57 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=1.06 $Y=1.815
+ $X2=1.06 $Y2=0.515
r181 2 52 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.475
+ $Y=2.325 $X2=1.6 $Y2=2.47
r182 1 48 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.245
+ $Y=0.595 $X2=1.37 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_1535_177# 1 2 10 11 12 13 15 16 23 24 28
+ 33 38
r74 30 33 8.13695 $w=3.28e-07 $l=2.33e-07 $layer=LI1_cond $X=9.002 $Y=2.365
+ $X2=9.235 $Y2=2.365
r75 26 28 5.85988 $w=2.93e-07 $l=1.5e-07 $layer=LI1_cond $X=9.287 $Y=0.955
+ $X2=9.287 $Y2=0.805
r76 24 42 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.97 $Y=2.9 $X2=8.97
+ $Y2=3.11
r77 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.97
+ $Y=2.9 $X2=8.97 $Y2=2.9
r78 21 30 2.26808 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=9.002 $Y=2.53
+ $X2=9.002 $Y2=2.365
r79 21 23 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=9.002 $Y=2.53
+ $X2=9.002 $Y2=2.9
r80 19 38 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=7.97 $Y=1.05
+ $X2=8.21 $Y2=1.05
r81 19 35 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=7.97 $Y=1.05
+ $X2=7.75 $Y2=1.05
r82 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.05 $X2=7.97 $Y2=1.05
r83 16 26 7.24045 $w=1.9e-07 $l=1.88611e-07 $layer=LI1_cond $X=9.14 $Y=1.05
+ $X2=9.287 $Y2=0.955
r84 16 18 68.2967 $w=1.88e-07 $l=1.17e-06 $layer=LI1_cond $X=9.14 $Y=1.05
+ $X2=7.97 $Y2=1.05
r85 13 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.21 $Y=0.885
+ $X2=8.21 $Y2=1.05
r86 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.21 $Y=0.885
+ $X2=8.21 $Y2=0.565
r87 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.805 $Y=3.11
+ $X2=8.97 $Y2=3.11
r88 11 12 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=8.805 $Y=3.11
+ $X2=7.825 $Y2=3.11
r89 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.75 $Y=3.035
+ $X2=7.825 $Y2=3.11
r90 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.75 $Y=3.035
+ $X2=7.75 $Y2=2.455
r91 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.75 $Y=1.215
+ $X2=7.75 $Y2=1.05
r92 7 10 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=7.75 $Y=1.215
+ $X2=7.75 $Y2=2.455
r93 2 33 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=9.11
+ $Y=2.155 $X2=9.235 $Y2=2.365
r94 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.18
+ $Y=0.595 $X2=9.305 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_1331_151# 1 2 3 10 12 13 15 16 18 20 22 23
+ 25 28 30 32 33 36 38 41 44 45 49 52 53 54 56 60 63 64 66 70 72 74 75 79 86
c179 74 0 1.18176e-19 $X=9.43 $Y=1.48
c180 66 0 1.77516e-19 $X=7.037 $Y=1.4
r181 80 86 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=11.87 $Y=1.395
+ $X2=12.005 $Y2=1.395
r182 80 83 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=11.87 $Y=1.395
+ $X2=11.82 $Y2=1.395
r183 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.87
+ $Y=1.395 $X2=11.87 $Y2=1.395
r184 76 79 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=11.665 $Y=1.395
+ $X2=11.87 $Y2=1.395
r185 74 75 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.43
+ $Y=1.48 $X2=9.43 $Y2=1.48
r186 68 70 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=8.395 $Y=2.39
+ $X2=8.62 $Y2=2.39
r187 63 64 9.50131 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=6.975 $Y=2.51
+ $X2=6.975 $Y2=2.285
r188 58 60 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=6.865 $Y=1.06
+ $X2=7.02 $Y2=1.06
r189 55 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.665 $Y=1.56
+ $X2=11.665 $Y2=1.395
r190 55 56 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=11.665 $Y=1.56
+ $X2=11.665 $Y2=2.395
r191 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.58 $Y=2.48
+ $X2=11.665 $Y2=2.395
r192 53 54 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=11.58 $Y=2.48
+ $X2=10.87 $Y2=2.48
r193 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.785 $Y=2.395
+ $X2=10.87 $Y2=2.48
r194 51 52 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=10.785 $Y=1.495
+ $X2=10.785 $Y2=2.395
r195 50 74 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=9.595 $Y=1.41
+ $X2=9.43 $Y2=1.405
r196 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.7 $Y=1.41
+ $X2=10.785 $Y2=1.495
r197 49 50 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=10.7 $Y=1.41
+ $X2=9.595 $Y2=1.41
r198 46 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.705 $Y=1.4
+ $X2=8.62 $Y2=1.4
r199 45 74 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=9.265 $Y=1.4
+ $X2=9.43 $Y2=1.405
r200 45 46 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.265 $Y=1.4
+ $X2=8.705 $Y2=1.4
r201 44 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=2.225
+ $X2=8.62 $Y2=2.39
r202 43 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.62 $Y=1.485
+ $X2=8.62 $Y2=1.4
r203 43 44 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=8.62 $Y=1.485
+ $X2=8.62 $Y2=2.225
r204 42 66 1.69765 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=7.14 $Y=1.4
+ $X2=7.037 $Y2=1.4
r205 41 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.535 $Y=1.4
+ $X2=8.62 $Y2=1.4
r206 41 42 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.535 $Y=1.4
+ $X2=7.14 $Y2=1.4
r207 39 66 4.7579 $w=1.87e-07 $l=8.5e-08 $layer=LI1_cond $X=7.037 $Y=1.485
+ $X2=7.037 $Y2=1.4
r208 39 64 43.2816 $w=2.03e-07 $l=8e-07 $layer=LI1_cond $X=7.037 $Y=1.485
+ $X2=7.037 $Y2=2.285
r209 38 66 4.7579 $w=1.87e-07 $l=9.31128e-08 $layer=LI1_cond $X=7.02 $Y=1.315
+ $X2=7.037 $Y2=1.4
r210 37 60 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.02 $Y=1.165
+ $X2=7.02 $Y2=1.06
r211 37 38 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.02 $Y=1.165
+ $X2=7.02 $Y2=1.315
r212 35 75 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=9.43 $Y=1.895
+ $X2=9.43 $Y2=1.48
r213 35 36 13.5877 $w=2.4e-07 $l=1.65e-07 $layer=POLY_cond $X=9.43 $Y=1.895
+ $X2=9.265 $Y2=1.895
r214 33 75 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=9.43 $Y=1.44 $X2=9.43
+ $Y2=1.48
r215 30 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.005 $Y=1.23
+ $X2=12.005 $Y2=1.395
r216 30 32 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=12.005 $Y=1.23
+ $X2=12.005 $Y2=0.7
r217 26 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.82 $Y=1.56
+ $X2=11.82 $Y2=1.395
r218 26 28 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=11.82 $Y=1.56
+ $X2=11.82 $Y2=2.465
r219 23 25 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.995 $Y=2.045
+ $X2=9.995 $Y2=2.475
r220 20 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.95 $Y=1.125
+ $X2=9.95 $Y2=0.805
r221 19 36 12.1617 $w=1.5e-07 $l=3.65582e-07 $layer=POLY_cond $X=9.595 $Y=1.97
+ $X2=9.265 $Y2=1.895
r222 18 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.92 $Y=1.97
+ $X2=9.995 $Y2=2.045
r223 18 19 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=9.92 $Y=1.97
+ $X2=9.595 $Y2=1.97
r224 17 33 38.4264 $w=3.3e-07 $l=3.11769e-07 $layer=POLY_cond $X=9.595 $Y=1.2
+ $X2=9.43 $Y2=1.44
r225 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.875 $Y=1.2
+ $X2=9.95 $Y2=1.125
r226 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.875 $Y=1.2
+ $X2=9.595 $Y2=1.2
r227 13 17 21.9219 $w=2.44e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.52 $Y=1.125
+ $X2=9.595 $Y2=1.2
r228 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.52 $Y=1.125
+ $X2=9.52 $Y2=0.805
r229 10 36 13.5877 $w=2.4e-07 $l=2.48948e-07 $layer=POLY_cond $X=9.45 $Y=2.045
+ $X2=9.265 $Y2=1.895
r230 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.45 $Y=2.045
+ $X2=9.45 $Y2=2.365
r231 3 68 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=2.245 $X2=8.395 $Y2=2.39
r232 2 63 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=6.835
+ $Y=2.245 $X2=6.975 $Y2=2.51
r233 1 58 182 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.755 $X2=6.865 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_2005_119# 1 2 7 11 15 17 22 23 27 29 31 41
r63 38 41 10.9545 $w=3.3e-07 $l=1.00623e-07 $layer=POLY_cond $X=10.565 $Y=1.485
+ $X2=10.505 $Y2=1.56
r64 32 41 40.4161 $w=3.22e-07 $l=2.7e-07 $layer=POLY_cond $X=10.505 $Y=1.83
+ $X2=10.505 $Y2=1.56
r65 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.445
+ $Y=1.83 $X2=10.445 $Y2=1.83
r66 29 31 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=10.405 $Y=1.985
+ $X2=10.405 $Y2=1.83
r67 25 29 13.5701 $w=1.68e-07 $l=2.08e-07 $layer=LI1_cond $X=10.197 $Y=2.07
+ $X2=10.405 $Y2=2.07
r68 25 27 5.86331 $w=2.83e-07 $l=1.45e-07 $layer=LI1_cond $X=10.197 $Y=2.155
+ $X2=10.197 $Y2=2.3
r69 23 38 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=10.565 $Y=1.07
+ $X2=10.565 $Y2=1.485
r70 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.565
+ $Y=1.07 $X2=10.565 $Y2=1.07
r71 19 22 9.28993 $w=5.13e-07 $l=4e-07 $layer=LI1_cond $X=10.165 $Y=0.897
+ $X2=10.565 $Y2=0.897
r72 13 17 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.42 $Y=1.485
+ $X2=11.405 $Y2=1.56
r73 13 15 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=11.42 $Y=1.485
+ $X2=11.42 $Y2=0.7
r74 9 17 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.39 $Y=1.635
+ $X2=11.405 $Y2=1.56
r75 9 11 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=11.39 $Y=1.635
+ $X2=11.39 $Y2=2.465
r76 8 41 20.6399 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=10.73 $Y=1.56
+ $X2=10.505 $Y2=1.56
r77 7 17 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.315 $Y=1.56
+ $X2=11.405 $Y2=1.56
r78 7 8 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=11.315 $Y=1.56
+ $X2=10.73 $Y2=1.56
r79 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=10.07
+ $Y=2.155 $X2=10.21 $Y2=2.3
r80 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.025
+ $Y=0.595 $X2=10.165 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48
+ 51 52 53 55 63 71 76 81 94 95 101 104 107 110 113
r147 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r148 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r149 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r150 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r151 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r154 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r155 92 114 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=9.84 $Y2=3.33
r156 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r157 89 113 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=9.885 $Y=3.33
+ $X2=9.727 $Y2=3.33
r158 89 91 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=9.885 $Y=3.33
+ $X2=11.28 $Y2=3.33
r159 88 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r160 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r162 85 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r163 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33 $X2=9.36
+ $Y2=3.33
r164 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r165 82 110 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=8.09 $Y=3.33
+ $X2=7.97 $Y2=3.33
r166 82 84 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.09 $Y=3.33
+ $X2=8.4 $Y2=3.33
r167 81 113 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=9.57 $Y=3.33
+ $X2=9.727 $Y2=3.33
r168 81 87 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.57 $Y=3.33
+ $X2=9.36 $Y2=3.33
r169 80 111 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r170 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r171 77 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.15 $Y=3.33
+ $X2=5.985 $Y2=3.33
r172 77 79 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.15 $Y=3.33
+ $X2=6.48 $Y2=3.33
r173 76 110 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.85 $Y=3.33
+ $X2=7.97 $Y2=3.33
r174 76 79 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=7.85 $Y=3.33
+ $X2=6.48 $Y2=3.33
r175 75 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r176 75 105 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.08 $Y2=3.33
r177 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r178 72 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=3.33
+ $X2=3.935 $Y2=3.33
r179 72 74 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=4.1 $Y=3.33
+ $X2=5.52 $Y2=3.33
r180 71 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=3.33
+ $X2=5.985 $Y2=3.33
r181 71 74 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.82 $Y=3.33 $X2=5.52
+ $Y2=3.33
r182 70 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r183 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r184 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r185 67 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r186 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r187 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r188 64 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.165 $Y2=3.33
r189 64 66 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.64 $Y2=3.33
r190 63 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.77 $Y=3.33
+ $X2=3.935 $Y2=3.33
r191 63 69 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.77 $Y=3.33
+ $X2=3.6 $Y2=3.33
r192 62 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r193 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r194 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r195 59 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r196 58 61 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r197 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r198 56 98 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.215 $Y2=3.33
r199 56 58 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.72 $Y2=3.33
r200 55 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=3.33
+ $X2=2.165 $Y2=3.33
r201 55 61 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r202 53 80 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r203 53 108 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6 $Y2=3.33
r204 51 91 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=11.44 $Y=3.33
+ $X2=11.28 $Y2=3.33
r205 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.44 $Y=3.33
+ $X2=11.605 $Y2=3.33
r206 50 94 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=11.77 $Y=3.33
+ $X2=12.24 $Y2=3.33
r207 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.77 $Y=3.33
+ $X2=11.605 $Y2=3.33
r208 46 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.605 $Y=3.245
+ $X2=11.605 $Y2=3.33
r209 46 48 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=11.605 $Y=3.245
+ $X2=11.605 $Y2=2.9
r210 42 113 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=9.727 $Y=3.245
+ $X2=9.727 $Y2=3.33
r211 42 44 33.8416 $w=3.13e-07 $l=9.25e-07 $layer=LI1_cond $X=9.727 $Y=3.245
+ $X2=9.727 $Y2=2.32
r212 38 110 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=3.33
r213 38 40 38.4148 $w=2.38e-07 $l=8e-07 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=2.445
r214 34 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=3.33
r215 34 36 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=2.825
r216 30 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=3.245
+ $X2=3.935 $Y2=3.33
r217 30 32 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.935 $Y=3.245
+ $X2=3.935 $Y2=2.93
r218 26 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=3.33
r219 26 28 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=2.84
r220 22 98 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=3.245
+ $X2=0.215 $Y2=3.33
r221 22 24 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.265 $Y=3.245
+ $X2=0.265 $Y2=2.775
r222 7 48 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=11.465
+ $Y=1.835 $X2=11.605 $Y2=2.9
r223 6 44 300 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=2 $X=9.525
+ $Y=2.155 $X2=9.665 $Y2=2.32
r224 5 40 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=7.825
+ $Y=2.245 $X2=7.965 $Y2=2.445
r225 4 36 600 $w=1.7e-07 $l=3.04672e-07 $layer=licon1_PDIFF $count=1 $X=5.75
+ $Y=2.665 $X2=5.985 $Y2=2.825
r226 3 32 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=2.665 $X2=3.935 $Y2=2.93
r227 2 28 600 $w=1.7e-07 $l=6.37848e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=2.325 $X2=2.165 $Y2=2.84
r228 1 24 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=2.28 $X2=0.265 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_494_119# 1 2 8 10 12 18 22
c39 10 0 3.46675e-19 $X=2.805 $Y=2.72
r40 20 22 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.69 $Y=1.85
+ $X2=2.805 $Y2=1.85
r41 16 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.715 $Y=2.885
+ $X2=2.805 $Y2=2.885
r42 12 14 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=0.81
+ $X2=2.63 $Y2=0.975
r43 10 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=2.72
+ $X2=2.805 $Y2=2.885
r44 9 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=1.935
+ $X2=2.805 $Y2=1.85
r45 9 10 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.805 $Y=1.935
+ $X2=2.805 $Y2=2.72
r46 8 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=1.765
+ $X2=2.69 $Y2=1.85
r47 8 14 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.69 $Y=1.765
+ $X2=2.69 $Y2=0.975
r48 2 16 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.665 $X2=2.715 $Y2=2.885
r49 1 12 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.595 $X2=2.61 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%Q 1 2 7 8 9 10 11
r21 11 30 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=11.225 $Y=2.035
+ $X2=11.225 $Y2=2.06
r22 10 11 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.225 $Y=1.665
+ $X2=11.225 $Y2=2.035
r23 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.225 $Y=1.295
+ $X2=11.225 $Y2=1.665
r24 8 9 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.225 $Y=0.925
+ $X2=11.225 $Y2=1.295
r25 7 8 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.225 $Y=0.555
+ $X2=11.225 $Y2=0.925
r26 2 30 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=11.05
+ $Y=1.835 $X2=11.175 $Y2=2.06
r27 1 7 91 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_NDIFF $count=2 $X=11.08
+ $Y=0.28 $X2=11.205 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%Q_N 1 2 7 8 9 10 11 12 13 25 35 38 40
r18 38 40 1.44581 $w=4.53e-07 $l=5.5e-08 $layer=LI1_cond $X=12.167 $Y=1.98
+ $X2=12.167 $Y2=2.035
r19 36 38 0.341737 $w=4.53e-07 $l=1.3e-08 $layer=LI1_cond $X=12.167 $Y=1.967
+ $X2=12.167 $Y2=1.98
r20 35 50 3.20123 $w=2.68e-07 $l=7.5e-08 $layer=LI1_cond $X=12.26 $Y=1.665
+ $X2=12.26 $Y2=1.74
r21 13 47 3.5488 $w=4.53e-07 $l=1.35e-07 $layer=LI1_cond $X=12.167 $Y=2.775
+ $X2=12.167 $Y2=2.91
r22 12 13 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=12.167 $Y=2.405
+ $X2=12.167 $Y2=2.775
r23 11 36 0.236587 $w=4.53e-07 $l=9e-09 $layer=LI1_cond $X=12.167 $Y=1.958
+ $X2=12.167 $Y2=1.967
r24 11 12 9.51605 $w=4.53e-07 $l=3.62e-07 $layer=LI1_cond $X=12.167 $Y=2.043
+ $X2=12.167 $Y2=2.405
r25 11 40 0.210299 $w=4.53e-07 $l=8e-09 $layer=LI1_cond $X=12.167 $Y=2.043
+ $X2=12.167 $Y2=2.035
r26 10 11 5.59922 $w=4.53e-07 $l=2.13e-07 $layer=LI1_cond $X=12.167 $Y=1.745
+ $X2=12.167 $Y2=1.958
r27 10 50 2.09279 $w=4.53e-07 $l=5e-09 $layer=LI1_cond $X=12.167 $Y=1.745
+ $X2=12.167 $Y2=1.74
r28 10 35 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=12.26 $Y=1.66
+ $X2=12.26 $Y2=1.665
r29 9 10 15.5793 $w=2.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.26 $Y=1.295
+ $X2=12.26 $Y2=1.66
r30 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.26 $Y=0.925
+ $X2=12.26 $Y2=1.295
r31 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.26 $Y=0.555
+ $X2=12.26 $Y2=0.925
r32 7 25 5.5488 $w=2.68e-07 $l=1.3e-07 $layer=LI1_cond $X=12.26 $Y=0.555
+ $X2=12.26 $Y2=0.425
r33 2 47 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.895
+ $Y=1.835 $X2=12.035 $Y2=2.91
r34 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.895
+ $Y=1.835 $X2=12.035 $Y2=1.98
r35 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.08
+ $Y=0.28 $X2=12.22 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48
+ 51 52 54 55 57 58 59 61 85 89 96 97 103 106 109
r130 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r131 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r132 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r133 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r134 97 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r135 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r136 94 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.91 $Y=0
+ $X2=11.745 $Y2=0
r137 94 96 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=11.91 $Y=0
+ $X2=12.24 $Y2=0
r138 93 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r139 93 107 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=9.84 $Y2=0
r140 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r141 90 106 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.865 $Y=0
+ $X2=9.735 $Y2=0
r142 90 92 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=9.865 $Y=0
+ $X2=11.28 $Y2=0
r143 89 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.58 $Y=0
+ $X2=11.745 $Y2=0
r144 89 92 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=11.58 $Y=0 $X2=11.28
+ $Y2=0
r145 88 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r146 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r147 85 106 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.605 $Y=0
+ $X2=9.735 $Y2=0
r148 85 87 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.605 $Y=0 $X2=9.36
+ $Y2=0
r149 84 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r150 83 84 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r151 80 83 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=8.4
+ $Y2=0
r152 80 81 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r153 78 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r154 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r155 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r156 74 77 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r157 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r158 72 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r159 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r160 69 72 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r161 69 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r162 68 71 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r163 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r164 66 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.81 $Y2=0
r165 66 68 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=2.16 $Y2=0
r166 65 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r167 65 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r168 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r169 62 100 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0
+ $X2=0.215 $Y2=0
r170 62 64 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r171 61 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0
+ $X2=1.81 $Y2=0
r172 61 64 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.645 $Y=0
+ $X2=0.72 $Y2=0
r173 59 84 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=6.24 $Y=0 $X2=8.4
+ $Y2=0
r174 59 81 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=0 $X2=5.52
+ $Y2=0
r175 57 83 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.62 $Y=0 $X2=8.4
+ $Y2=0
r176 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=0 $X2=8.785
+ $Y2=0
r177 56 87 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.95 $Y=0 $X2=9.36
+ $Y2=0
r178 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.95 $Y=0 $X2=8.785
+ $Y2=0
r179 55 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.52
+ $Y2=0
r180 54 77 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.25 $Y=0 $X2=5.04
+ $Y2=0
r181 54 55 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.25 $Y=0 $X2=5.385
+ $Y2=0
r182 51 71 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.725 $Y=0 $X2=3.6
+ $Y2=0
r183 51 52 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.725 $Y=0 $X2=3.825
+ $Y2=0
r184 50 74 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.925 $Y=0
+ $X2=4.08 $Y2=0
r185 50 52 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.825
+ $Y2=0
r186 46 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.745 $Y=0.085
+ $X2=11.745 $Y2=0
r187 46 48 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.745 $Y=0.085
+ $X2=11.745 $Y2=0.425
r188 42 106 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.735 $Y=0.085
+ $X2=9.735 $Y2=0
r189 42 44 31.9138 $w=2.58e-07 $l=7.2e-07 $layer=LI1_cond $X=9.735 $Y=0.085
+ $X2=9.735 $Y2=0.805
r190 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0
r191 38 40 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0.565
r192 34 55 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=0.085
+ $X2=5.385 $Y2=0
r193 34 36 35.2135 $w=2.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.385 $Y=0.085
+ $X2=5.385 $Y2=0.91
r194 30 52 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=0.085
+ $X2=3.825 $Y2=0
r195 30 32 36.3227 $w=1.98e-07 $l=6.55e-07 $layer=LI1_cond $X=3.825 $Y=0.085
+ $X2=3.825 $Y2=0.74
r196 26 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0
r197 26 28 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.735
r198 22 100 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.215 $Y2=0
r199 22 24 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.935
r200 7 48 91 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=2 $X=11.495
+ $Y=0.28 $X2=11.745 $Y2=0.425
r201 6 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.595
+ $Y=0.595 $X2=9.735 $Y2=0.805
r202 5 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.645
+ $Y=0.355 $X2=8.785 $Y2=0.565
r203 4 36 182 $w=1.7e-07 $l=2.65518e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.845 $X2=5.415 $Y2=0.91
r204 3 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.69
+ $Y=0.595 $X2=3.83 $Y2=0.74
r205 2 28 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.595 $X2=1.81 $Y2=0.735
r206 1 24 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.78 $X2=0.265 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_1141_125# 1 2 9 11 13
r24 11 13 89.0354 $w=1.78e-07 $l=1.445e-06 $layer=LI1_cond $X=6.01 $Y=0.355
+ $X2=7.455 $Y2=0.355
r25 7 11 7.17723 $w=1.8e-07 $l=1.74284e-07 $layer=LI1_cond $X=5.875 $Y=0.445
+ $X2=6.01 $Y2=0.355
r26 7 9 19.8476 $w=2.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.875 $Y=0.445
+ $X2=5.875 $Y2=0.91
r27 2 13 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.535 $X2=7.455 $Y2=0.35
r28 1 9 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.625 $X2=5.845 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_1%A_1248_151# 1 2 7 9 15
c30 9 0 1.11656e-19 $X=6.365 $Y=0.7
c31 7 0 1.50513e-19 $X=7.83 $Y=0.7
r32 15 17 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.965 $Y=0.565
+ $X2=7.965 $Y2=0.7
r33 9 12 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=6.365 $Y=0.7
+ $X2=6.365 $Y2=0.96
r34 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.53 $Y=0.7 $X2=6.365
+ $Y2=0.7
r35 7 17 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.83 $Y=0.7 $X2=7.965
+ $Y2=0.7
r36 7 8 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=7.83 $Y=0.7 $X2=6.53
+ $Y2=0.7
r37 2 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=7.87
+ $Y=0.355 $X2=7.995 $Y2=0.565
r38 1 12 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=6.24
+ $Y=0.755 $X2=6.365 $Y2=0.96
.ends

