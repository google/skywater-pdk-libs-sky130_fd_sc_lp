* File: sky130_fd_sc_lp__o31ai_m.pxi.spice
* Created: Fri Aug 28 11:16:53 2020
* 
x_PM_SKY130_FD_SC_LP__O31AI_M%A1 N_A1_c_64_n N_A1_M1007_g N_A1_c_65_n
+ N_A1_M1002_g N_A1_c_60_n N_A1_c_61_n N_A1_c_66_n N_A1_c_67_n A1 A1 A1 A1
+ N_A1_c_63_n PM_SKY130_FD_SC_LP__O31AI_M%A1
x_PM_SKY130_FD_SC_LP__O31AI_M%A2 N_A2_M1005_g N_A2_M1000_g N_A2_c_102_n
+ N_A2_c_103_n A2 A2 A2 N_A2_c_100_n PM_SKY130_FD_SC_LP__O31AI_M%A2
x_PM_SKY130_FD_SC_LP__O31AI_M%A3 N_A3_M1003_g N_A3_M1001_g N_A3_c_145_n
+ N_A3_c_149_n A3 A3 N_A3_c_151_n PM_SKY130_FD_SC_LP__O31AI_M%A3
x_PM_SKY130_FD_SC_LP__O31AI_M%B1 N_B1_M1004_g N_B1_c_194_n N_B1_M1006_g
+ N_B1_c_189_n N_B1_c_190_n N_B1_c_195_n N_B1_c_196_n N_B1_c_191_n B1 B1
+ N_B1_c_193_n PM_SKY130_FD_SC_LP__O31AI_M%B1
x_PM_SKY130_FD_SC_LP__O31AI_M%VPWR N_VPWR_M1002_s N_VPWR_M1006_d N_VPWR_c_232_n
+ N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n VPWR
+ N_VPWR_c_237_n N_VPWR_c_231_n PM_SKY130_FD_SC_LP__O31AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O31AI_M%Y N_Y_M1004_d N_Y_M1001_d N_Y_c_268_n N_Y_c_267_n
+ Y PM_SKY130_FD_SC_LP__O31AI_M%Y
x_PM_SKY130_FD_SC_LP__O31AI_M%VGND N_VGND_M1007_s N_VGND_M1005_d N_VGND_c_299_n
+ N_VGND_c_300_n N_VGND_c_301_n VGND N_VGND_c_302_n N_VGND_c_303_n
+ N_VGND_c_304_n N_VGND_c_305_n PM_SKY130_FD_SC_LP__O31AI_M%VGND
x_PM_SKY130_FD_SC_LP__O31AI_M%A_126_129# N_A_126_129#_M1007_d
+ N_A_126_129#_M1003_d N_A_126_129#_c_327_n N_A_126_129#_c_328_n
+ N_A_126_129#_c_329_n N_A_126_129#_c_330_n
+ PM_SKY130_FD_SC_LP__O31AI_M%A_126_129#
cc_1 VNB N_A1_c_60_n 0.0209549f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.175
cc_2 VNB N_A1_c_61_n 0.0258694f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.325
cc_3 VNB A1 0.0242032f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_63_n 0.0278466f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.34
cc_5 VNB N_A2_M1005_g 0.0357598f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.175
cc_6 VNB A2 0.00360548f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_7 VNB N_A2_c_100_n 0.0126602f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_8 VNB N_A3_M1003_g 0.0367685f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.175
cc_9 VNB N_A3_c_145_n 0.0197307f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.325
cc_10 VNB A3 0.00181747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_M1004_g 0.0119526f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.855
cc_12 VNB N_B1_c_189_n 0.0232145f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.885
cc_13 VNB N_B1_c_190_n 0.0100598f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.325
cc_14 VNB N_B1_c_191_n 0.0187047f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_15 VNB B1 0.0249636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_193_n 0.0468659f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_VPWR_c_231_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.665
cc_18 VNB N_Y_c_267_n 0.0358824f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.325
cc_19 VNB N_VGND_c_299_n 0.0137364f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.885
cc_20 VNB N_VGND_c_300_n 0.0270131f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.325
cc_21 VNB N_VGND_c_301_n 0.0159532f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_22 VNB N_VGND_c_302_n 0.0206207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_303_n 0.0318693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_304_n 0.176361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_305_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_126_129#_c_327_n 9.46579e-19 $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.325
cc_27 VNB N_A_126_129#_c_328_n 0.0103888f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.325
cc_28 VNB N_A_126_129#_c_329_n 0.00786248f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.68
cc_29 VNB N_A_126_129#_c_330_n 0.00249597f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.49
cc_30 VPB N_A1_c_64_n 0.0367588f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.415
cc_31 VPB N_A1_c_65_n 0.0207587f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.565
cc_32 VPB N_A1_c_66_n 0.0186543f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.845
cc_33 VPB N_A1_c_67_n 0.0318954f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.49
cc_34 VPB A1 0.0362996f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_35 VPB N_A1_c_63_n 0.00196603f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.34
cc_36 VPB N_A2_M1000_g 0.0310246f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.885
cc_37 VPB N_A2_c_102_n 0.0220978f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.325
cc_38 VPB N_A2_c_103_n 0.017776f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.68
cc_39 VPB A2 0.0143813f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.845
cc_40 VPB N_A2_c_100_n 0.00288579f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_41 VPB N_A3_M1001_g 0.0362959f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.885
cc_42 VPB N_A3_c_145_n 0.00348819f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.325
cc_43 VPB N_A3_c_149_n 0.0244832f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.49
cc_44 VPB A3 0.00175777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A3_c_151_n 0.0315044f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_46 VPB N_B1_c_194_n 0.0213538f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.855
cc_47 VPB N_B1_c_195_n 0.0237852f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.175
cc_48 VPB N_B1_c_196_n 0.00994894f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.325
cc_49 VPB N_B1_c_191_n 0.0428638f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.845
cc_50 VPB N_VPWR_c_232_n 0.01277f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.325
cc_51 VPB N_VPWR_c_233_n 0.0131778f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.325
cc_52 VPB N_VPWR_c_234_n 0.00495479f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.845
cc_53 VPB N_VPWR_c_235_n 0.0121672f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.49
cc_54 VPB N_VPWR_c_236_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_237_n 0.037847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_231_n 0.0496523f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.665
cc_57 VPB N_Y_c_268_n 0.0113196f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.885
cc_58 VPB N_Y_c_267_n 0.0354271f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.325
cc_59 VPB Y 0.00410841f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.845
cc_60 N_A1_c_60_n N_A2_M1005_g 0.0203928f $X=0.425 $Y=1.175 $X2=0 $Y2=0
cc_61 A1 N_A2_M1005_g 0.00132697f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A1_c_63_n N_A2_M1005_g 0.00782722f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_63 N_A1_c_64_n N_A2_M1000_g 0.00479041f $X=0.475 $Y=2.415 $X2=0 $Y2=0
cc_64 N_A1_c_67_n N_A2_M1000_g 0.0528124f $X=0.695 $Y=2.49 $X2=0 $Y2=0
cc_65 A1 N_A2_M1000_g 2.64504e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A1_c_66_n N_A2_c_102_n 0.011018f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_67 N_A1_c_64_n N_A2_c_103_n 0.011018f $X=0.475 $Y=2.415 $X2=0 $Y2=0
cc_68 N_A1_c_64_n A2 0.00167127f $X=0.475 $Y=2.415 $X2=0 $Y2=0
cc_69 N_A1_c_67_n A2 7.60954e-19 $X=0.695 $Y=2.49 $X2=0 $Y2=0
cc_70 A1 A2 0.0367916f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A1_c_63_n A2 0.00213891f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_72 A1 N_A2_c_100_n 0.00229979f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A1_c_63_n N_A2_c_100_n 0.011018f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_74 N_A1_c_65_n N_VPWR_c_232_n 0.0112929f $X=0.695 $Y=2.565 $X2=0 $Y2=0
cc_75 N_A1_c_67_n N_VPWR_c_232_n 0.00650864f $X=0.695 $Y=2.49 $X2=0 $Y2=0
cc_76 A1 N_VPWR_c_232_n 0.00700086f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A1_c_65_n N_VPWR_c_237_n 0.00486043f $X=0.695 $Y=2.565 $X2=0 $Y2=0
cc_78 N_A1_c_65_n N_VPWR_c_231_n 0.00818711f $X=0.695 $Y=2.565 $X2=0 $Y2=0
cc_79 A1 N_VPWR_c_231_n 0.00709409f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A1_c_60_n N_VGND_c_300_n 0.0037597f $X=0.425 $Y=1.175 $X2=0 $Y2=0
cc_81 N_A1_c_61_n N_VGND_c_300_n 0.00150576f $X=0.425 $Y=1.325 $X2=0 $Y2=0
cc_82 A1 N_VGND_c_300_n 0.0141001f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A1_c_60_n N_VGND_c_302_n 0.00404937f $X=0.425 $Y=1.175 $X2=0 $Y2=0
cc_84 N_A1_c_60_n N_VGND_c_304_n 0.0046394f $X=0.425 $Y=1.175 $X2=0 $Y2=0
cc_85 N_A1_c_60_n N_A_126_129#_c_327_n 0.00123209f $X=0.425 $Y=1.175 $X2=0 $Y2=0
cc_86 N_A1_c_60_n N_A_126_129#_c_329_n 0.00305231f $X=0.425 $Y=1.175 $X2=0 $Y2=0
cc_87 A1 N_A_126_129#_c_329_n 0.00833984f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A2_M1005_g N_A3_M1003_g 0.0309958f $X=0.985 $Y=0.855 $X2=0 $Y2=0
cc_89 N_A2_M1000_g N_A3_M1001_g 0.03628f $X=1.055 $Y=2.885 $X2=0 $Y2=0
cc_90 A2 N_A3_c_145_n 0.00151295f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A2_c_100_n N_A3_c_145_n 0.00955213f $X=0.965 $Y=1.7 $X2=0 $Y2=0
cc_92 N_A2_c_103_n N_A3_c_149_n 0.03628f $X=0.965 $Y=2.205 $X2=0 $Y2=0
cc_93 A2 N_A3_c_149_n 0.0082743f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_94 A2 A3 0.0329214f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A2_c_100_n A3 4.99685e-19 $X=0.965 $Y=1.7 $X2=0 $Y2=0
cc_96 A2 N_A3_c_151_n 0.00364649f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A2_c_100_n N_A3_c_151_n 0.0186467f $X=0.965 $Y=1.7 $X2=0 $Y2=0
cc_98 N_A2_M1000_g N_VPWR_c_232_n 0.00238543f $X=1.055 $Y=2.885 $X2=0 $Y2=0
cc_99 N_A2_M1000_g N_VPWR_c_237_n 0.00585385f $X=1.055 $Y=2.885 $X2=0 $Y2=0
cc_100 N_A2_M1000_g N_VPWR_c_231_n 0.00619515f $X=1.055 $Y=2.885 $X2=0 $Y2=0
cc_101 A2 N_VPWR_c_231_n 0.0147347f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_102 A2 Y 0.00325204f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A2_M1005_g N_VGND_c_301_n 0.00175675f $X=0.985 $Y=0.855 $X2=0 $Y2=0
cc_104 N_A2_M1005_g N_VGND_c_302_n 0.00404937f $X=0.985 $Y=0.855 $X2=0 $Y2=0
cc_105 N_A2_M1005_g N_VGND_c_304_n 0.0046394f $X=0.985 $Y=0.855 $X2=0 $Y2=0
cc_106 N_A2_M1005_g N_A_126_129#_c_327_n 6.39777e-19 $X=0.985 $Y=0.855 $X2=0
+ $Y2=0
cc_107 N_A2_M1005_g N_A_126_129#_c_328_n 0.0148083f $X=0.985 $Y=0.855 $X2=0
+ $Y2=0
cc_108 A2 N_A_126_129#_c_328_n 0.0242269f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A2_c_100_n N_A_126_129#_c_328_n 8.46827e-19 $X=0.965 $Y=1.7 $X2=0 $Y2=0
cc_110 N_A2_c_100_n N_A_126_129#_c_329_n 0.0031789f $X=0.965 $Y=1.7 $X2=0 $Y2=0
cc_111 N_A2_M1005_g N_A_126_129#_c_330_n 5.89464e-19 $X=0.985 $Y=0.855 $X2=0
+ $Y2=0
cc_112 N_A3_c_145_n N_B1_c_190_n 0.00606969f $X=1.592 $Y=1.685 $X2=0 $Y2=0
cc_113 N_A3_M1001_g N_B1_c_196_n 0.0188786f $X=1.415 $Y=2.885 $X2=0 $Y2=0
cc_114 N_A3_c_149_n N_B1_c_196_n 0.00569692f $X=1.592 $Y=2.205 $X2=0 $Y2=0
cc_115 N_A3_M1003_g N_B1_c_191_n 0.00167374f $X=1.415 $Y=0.855 $X2=0 $Y2=0
cc_116 N_A3_M1001_g N_B1_c_191_n 0.00167374f $X=1.415 $Y=2.885 $X2=0 $Y2=0
cc_117 N_A3_c_145_n N_B1_c_191_n 0.0358662f $X=1.592 $Y=1.685 $X2=0 $Y2=0
cc_118 A3 N_B1_c_191_n 6.34285e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_119 N_A3_M1003_g B1 0.00119574f $X=1.415 $Y=0.855 $X2=0 $Y2=0
cc_120 N_A3_M1003_g N_B1_c_193_n 0.0209039f $X=1.415 $Y=0.855 $X2=0 $Y2=0
cc_121 N_A3_M1001_g N_VPWR_c_237_n 0.00585385f $X=1.415 $Y=2.885 $X2=0 $Y2=0
cc_122 N_A3_M1001_g N_VPWR_c_231_n 0.0108402f $X=1.415 $Y=2.885 $X2=0 $Y2=0
cc_123 N_A3_c_149_n N_Y_c_268_n 7.26846e-19 $X=1.592 $Y=2.205 $X2=0 $Y2=0
cc_124 N_A3_M1003_g N_Y_c_267_n 0.00481025f $X=1.415 $Y=0.855 $X2=0 $Y2=0
cc_125 N_A3_M1001_g N_Y_c_267_n 0.00465611f $X=1.415 $Y=2.885 $X2=0 $Y2=0
cc_126 N_A3_c_145_n N_Y_c_267_n 0.00499578f $X=1.592 $Y=1.685 $X2=0 $Y2=0
cc_127 A3 N_Y_c_267_n 0.043153f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A3_M1001_g Y 0.00580523f $X=1.415 $Y=2.885 $X2=0 $Y2=0
cc_129 N_A3_c_149_n Y 0.00313638f $X=1.592 $Y=2.205 $X2=0 $Y2=0
cc_130 A3 Y 0.0117696f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A3_M1003_g N_VGND_c_301_n 0.00125029f $X=1.415 $Y=0.855 $X2=0 $Y2=0
cc_132 N_A3_M1003_g N_VGND_c_303_n 0.00404937f $X=1.415 $Y=0.855 $X2=0 $Y2=0
cc_133 N_A3_M1003_g N_VGND_c_304_n 0.0046394f $X=1.415 $Y=0.855 $X2=0 $Y2=0
cc_134 N_A3_M1003_g N_A_126_129#_c_328_n 0.0151418f $X=1.415 $Y=0.855 $X2=0
+ $Y2=0
cc_135 N_A3_M1003_g N_A_126_129#_c_330_n 0.0095446f $X=1.415 $Y=0.855 $X2=0
+ $Y2=0
cc_136 N_A3_c_145_n N_A_126_129#_c_330_n 0.00604019f $X=1.592 $Y=1.685 $X2=0
+ $Y2=0
cc_137 A3 N_A_126_129#_c_330_n 0.0108317f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_138 N_B1_c_195_n N_VPWR_c_233_n 2.28363e-19 $X=2.085 $Y=2.49 $X2=0 $Y2=0
cc_139 N_B1_c_194_n N_VPWR_c_234_n 0.00460896f $X=1.845 $Y=2.565 $X2=0 $Y2=0
cc_140 N_B1_c_195_n N_VPWR_c_234_n 0.0014062f $X=2.085 $Y=2.49 $X2=0 $Y2=0
cc_141 N_B1_c_194_n N_VPWR_c_237_n 0.00437852f $X=1.845 $Y=2.565 $X2=0 $Y2=0
cc_142 N_B1_c_194_n N_VPWR_c_231_n 0.00702259f $X=1.845 $Y=2.565 $X2=0 $Y2=0
cc_143 N_B1_c_194_n N_Y_c_268_n 0.00544972f $X=1.845 $Y=2.565 $X2=0 $Y2=0
cc_144 N_B1_c_195_n N_Y_c_268_n 0.0123568f $X=2.085 $Y=2.49 $X2=0 $Y2=0
cc_145 N_B1_c_196_n N_Y_c_268_n 0.00653471f $X=1.92 $Y=2.49 $X2=0 $Y2=0
cc_146 N_B1_M1004_g N_Y_c_267_n 0.00686527f $X=1.845 $Y=0.855 $X2=0 $Y2=0
cc_147 N_B1_c_189_n N_Y_c_267_n 0.0156536f $X=2.085 $Y=1.25 $X2=0 $Y2=0
cc_148 N_B1_c_195_n N_Y_c_267_n 0.00369412f $X=2.085 $Y=2.49 $X2=0 $Y2=0
cc_149 N_B1_c_191_n N_Y_c_267_n 0.0386708f $X=2.16 $Y=2.415 $X2=0 $Y2=0
cc_150 B1 N_Y_c_267_n 0.0203829f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_151 N_B1_c_193_n N_Y_c_267_n 4.83328e-19 $X=1.935 $Y=0.37 $X2=0 $Y2=0
cc_152 N_B1_c_194_n Y 0.0017667f $X=1.845 $Y=2.565 $X2=0 $Y2=0
cc_153 B1 N_VGND_c_301_n 0.0196812f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_154 N_B1_c_193_n N_VGND_c_301_n 0.00285822f $X=1.935 $Y=0.37 $X2=0 $Y2=0
cc_155 B1 N_VGND_c_303_n 0.036111f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_156 N_B1_c_193_n N_VGND_c_303_n 0.00634371f $X=1.935 $Y=0.37 $X2=0 $Y2=0
cc_157 B1 N_VGND_c_304_n 0.0229022f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_158 N_B1_c_193_n N_VGND_c_304_n 0.00905322f $X=1.935 $Y=0.37 $X2=0 $Y2=0
cc_159 N_B1_M1004_g N_A_126_129#_c_330_n 0.00531986f $X=1.845 $Y=0.855 $X2=0
+ $Y2=0
cc_160 N_B1_c_190_n N_A_126_129#_c_330_n 0.00347911f $X=1.92 $Y=1.25 $X2=0 $Y2=0
cc_161 B1 N_A_126_129#_c_330_n 0.0124558f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_162 N_VPWR_c_231_n A_154_535# 0.00620535f $X=2.16 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_163 N_VPWR_c_231_n A_226_535# 0.00465602f $X=2.16 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_164 N_VPWR_c_231_n N_Y_M1001_d 0.00352441f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_c_233_n N_Y_c_268_n 0.00237396f $X=2.06 $Y=3.245 $X2=0 $Y2=0
cc_166 N_VPWR_c_234_n N_Y_c_268_n 0.0157159f $X=2.06 $Y=2.95 $X2=0 $Y2=0
cc_167 N_VPWR_c_237_n N_Y_c_268_n 0.00259728f $X=1.955 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_231_n N_Y_c_268_n 0.00919155f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_169 N_VPWR_c_237_n Y 0.0104096f $X=1.955 $Y=3.33 $X2=0 $Y2=0
cc_170 N_VPWR_c_231_n Y 0.00898566f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_171 N_Y_c_267_n N_VGND_c_304_n 0.00290388f $X=2.14 $Y=0.92 $X2=0 $Y2=0
cc_172 N_Y_c_267_n N_A_126_129#_c_330_n 0.0243909f $X=2.14 $Y=0.92 $X2=0 $Y2=0
cc_173 N_VGND_c_304_n N_A_126_129#_c_327_n 0.00844339f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_174 N_VGND_c_301_n N_A_126_129#_c_328_n 0.0139641f $X=1.2 $Y=0.77 $X2=0 $Y2=0
cc_175 N_VGND_c_304_n N_A_126_129#_c_330_n 0.0051571f $X=2.16 $Y=0 $X2=0 $Y2=0
