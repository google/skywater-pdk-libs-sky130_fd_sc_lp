# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux4_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__mux4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685000 1.570000 7.620000 1.855000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.785000 1.345000 6.165000 2.120000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.685000 1.570000 5.615000 1.905000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425000 1.145000 4.165000 2.265000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.790000 1.325000 8.120000 1.905000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065000 1.285000 2.325000 2.120000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 0.255000 3.255000 2.265000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.095000  0.670000 0.385000 2.815000 ;
      RECT 0.095000  2.815000 1.635000 2.985000 ;
      RECT 0.555000  0.325000 1.635000 0.495000 ;
      RECT 0.555000  0.495000 0.775000 2.635000 ;
      RECT 0.955000  0.665000 1.285000 0.895000 ;
      RECT 0.955000  0.895000 1.125000 1.995000 ;
      RECT 0.955000  1.995000 1.295000 2.575000 ;
      RECT 1.295000  1.065000 2.155000 1.115000 ;
      RECT 1.295000  1.115000 1.895000 1.825000 ;
      RECT 1.465000  0.495000 1.635000 0.525000 ;
      RECT 1.465000  0.525000 2.855000 0.695000 ;
      RECT 1.465000  2.435000 4.750000 2.605000 ;
      RECT 1.465000  2.605000 1.635000 2.815000 ;
      RECT 1.565000  1.825000 1.895000 2.265000 ;
      RECT 1.725000  0.865000 2.155000 1.065000 ;
      RECT 2.485000  0.085000 2.815000 0.355000 ;
      RECT 2.525000  2.785000 2.855000 3.245000 ;
      RECT 2.605000  0.695000 2.855000 1.515000 ;
      RECT 3.385000  2.785000 3.715000 3.245000 ;
      RECT 3.425000  0.085000 4.015000 0.975000 ;
      RECT 4.345000  0.565000 4.790000 0.825000 ;
      RECT 4.345000  0.825000 4.515000 2.075000 ;
      RECT 4.345000  2.075000 4.750000 2.435000 ;
      RECT 4.420000  2.605000 4.750000 2.745000 ;
      RECT 4.695000  0.995000 6.155000 1.165000 ;
      RECT 4.695000  1.165000 5.025000 1.400000 ;
      RECT 5.210000  2.075000 5.540000 2.290000 ;
      RECT 5.210000  2.290000 5.990000 3.245000 ;
      RECT 5.485000  0.085000 5.815000 0.825000 ;
      RECT 5.985000  0.265000 7.130000 0.435000 ;
      RECT 5.985000  0.435000 6.155000 0.995000 ;
      RECT 6.335000  0.605000 6.780000 0.815000 ;
      RECT 6.335000  0.815000 6.515000 2.075000 ;
      RECT 6.335000  2.075000 6.830000 2.745000 ;
      RECT 6.685000  0.985000 8.470000 1.155000 ;
      RECT 6.685000  1.155000 7.130000 1.400000 ;
      RECT 6.960000  0.435000 7.130000 0.985000 ;
      RECT 7.350000  0.085000 7.680000 0.815000 ;
      RECT 7.485000  2.085000 7.815000 3.245000 ;
      RECT 7.850000  0.640000 8.110000 0.985000 ;
      RECT 7.985000  2.075000 8.470000 2.745000 ;
      RECT 8.300000  1.155000 8.470000 2.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  2.320000 1.285000 2.490000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  2.320000 6.565000 2.490000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
    LAYER met1 ;
      RECT 1.055000 2.290000 1.345000 2.335000 ;
      RECT 1.055000 2.335000 6.625000 2.475000 ;
      RECT 1.055000 2.475000 1.345000 2.520000 ;
      RECT 6.335000 2.290000 6.625000 2.335000 ;
      RECT 6.335000 2.475000 6.625000 2.520000 ;
  END
END sky130_fd_sc_lp__mux4_2
