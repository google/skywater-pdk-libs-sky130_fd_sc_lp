* File: sky130_fd_sc_lp__nand4_lp.spice
* Created: Wed Sep  2 10:05:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4_lp.pex.spice"
.subckt sky130_fd_sc_lp__nand4_lp  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1002 A_132_47# N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1006 A_210_47# N_C_M1006_g A_132_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1003 A_324_47# N_B_M1003_g A_210_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0882 PD=0.84 PS=0.84 NRD=44.28 NRS=44.28 M=1 R=2.8 SA=75001.2 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g A_324_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0882 PD=1.41 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75001.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_D_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_Y_M1005_d VPB PHIGHVT L=0.25 W=1 AD=0.145
+ AS=0.14 PD=1.29 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.145 PD=1.28 PS=1.29 NRD=0 NRS=1.9503 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_Y_M1007_d VPB PHIGHVT L=0.25 W=1 AD=0.35
+ AS=0.14 PD=2.7 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
c_27 VNB 0 1.38359e-19 $X=0 $Y=0
c_48 VPB 0 1.89209e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nand4_lp.pxi.spice"
*
.ends
*
*
