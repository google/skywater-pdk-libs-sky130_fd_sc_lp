* File: sky130_fd_sc_lp__a221o_m.spice
* Created: Fri Aug 28 09:52:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221o_m.pex.spice"
.subckt sky130_fd_sc_lp__a221o_m  VNB VPB A2 A1 B1 B2 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_33_153#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1007 A_196_47# N_A2_M1007_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_33_153#_M1008_d N_A1_M1008_g A_196_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.10605 AS=0.0441 PD=0.925 PS=0.63 NRD=64.284 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1005 A_399_47# N_B1_M1005_g N_A_33_153#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.10605 PD=0.63 PS=0.925 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B2_M1003_g A_399_47# VNB NSHORT L=0.15 W=0.42 AD=0.09135
+ AS=0.0441 PD=0.855 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_33_153#_M1011_d N_C1_M1011_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.09135 PD=1.37 PS=0.855 NRD=0 NRS=44.28 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_33_153#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_233_535#_M1010_d N_A2_M1010_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_233_535#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_233_535#_M1006_d N_B1_M1006_g N_A_337_397#_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_A_337_397#_M1001_d N_B2_M1001_g N_A_233_535#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_33_153#_M1009_d N_C1_M1009_g N_A_337_397#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_42 VNB 0 1.46329e-19 $X=0 $Y=0
c_78 VPB 0 1.69271e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a221o_m.pxi.spice"
*
.ends
*
*
