* File: sky130_fd_sc_lp__o2bb2ai_lp.pex.spice
* Created: Fri Aug 28 11:13:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%A1_N 3 7 9 10 14
r31 14 17 67.1496 $w=5.05e-07 $l=5.05e-07 $layer=POLY_cond $X=0.472 $Y=1.39
+ $X2=0.472 $Y2=1.895
r32 14 16 46.6818 $w=5.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.472 $Y=1.39
+ $X2=0.472 $Y2=1.225
r33 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.39 $X2=0.385 $Y2=1.39
r34 10 15 8.68279 $w=3.63e-07 $l=2.75e-07 $layer=LI1_cond $X=0.307 $Y=1.665
+ $X2=0.307 $Y2=1.39
r35 9 15 2.99951 $w=3.63e-07 $l=9.5e-08 $layer=LI1_cond $X=0.307 $Y=1.295
+ $X2=0.307 $Y2=1.39
r36 7 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.6 $Y=2.595 $X2=0.6
+ $Y2=1.895
r37 3 16 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.495 $Y=0.495
+ $X2=0.495 $Y2=1.225
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%A2_N 3 5 7 11 13 16
r52 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=1.07 $X2=1.13 $Y2=1.07
r53 13 17 1.24963 $w=6.68e-07 $l=7e-08 $layer=LI1_cond $X=1.2 $Y=1.24 $X2=1.13
+ $Y2=1.24
r54 12 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.13 $Y=1.41
+ $X2=1.13 $Y2=1.07
r55 11 16 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.13 $Y=0.985
+ $X2=1.13 $Y2=1.07
r56 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.052 $Y=0.835
+ $X2=1.052 $Y2=0.985
r57 5 12 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.575
+ $X2=1.13 $Y2=1.41
r58 5 7 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.13 $Y=1.575
+ $X2=1.13 $Y2=2.595
r59 3 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.885 $Y=0.495
+ $X2=0.885 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%A_145_419# 1 2 9 12 13 15 18 20 21 24 26
+ 31 33 41
c80 13 0 1.28636e-19 $X=1.925 $Y=0.91
r81 40 41 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.795 $Y=1.77
+ $X2=1.845 $Y2=1.77
r82 34 40 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.67 $Y=1.77
+ $X2=1.795 $Y2=1.77
r83 33 36 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.63 $Y=1.77 $X2=1.63
+ $Y2=1.85
r84 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.77 $X2=1.67 $Y2=1.77
r85 27 31 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.03 $Y=1.85 $X2=0.85
+ $Y2=1.85
r86 26 36 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.505 $Y=1.85
+ $X2=1.63 $Y2=1.85
r87 26 27 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.505 $Y=1.85
+ $X2=1.03 $Y2=1.85
r88 22 31 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=1.935
+ $X2=0.85 $Y2=1.85
r89 22 24 9.76375 $w=3.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.85 $Y=1.935
+ $X2=0.85 $Y2=2.24
r90 21 31 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.755 $Y=1.765
+ $X2=0.85 $Y2=1.85
r91 20 30 12.7545 $w=3.3e-07 $l=4.45393e-07 $layer=LI1_cond $X=0.755 $Y=0.725
+ $X2=1.1 $Y2=0.495
r92 20 21 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=0.755 $Y=0.725
+ $X2=0.755 $Y2=1.765
r93 16 18 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=1.845 $Y=0.985
+ $X2=1.925 $Y2=0.985
r94 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=0.91
+ $X2=1.925 $Y2=0.985
r95 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.925 $Y=0.91
+ $X2=1.925 $Y2=0.625
r96 12 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.605
+ $X2=1.845 $Y2=1.77
r97 11 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.06
+ $X2=1.845 $Y2=0.985
r98 11 12 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.845 $Y=1.06
+ $X2=1.845 $Y2=1.605
r99 7 40 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.935
+ $X2=1.795 $Y2=1.77
r100 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.795 $Y=1.935
+ $X2=1.795 $Y2=2.595
r101 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.725
+ $Y=2.095 $X2=0.865 $Y2=2.24
r102 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.285 $X2=1.1 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%B2 3 7 9 10 14
c38 3 0 2.28059e-20 $X=2.325 $Y=2.595
r39 14 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.56
+ $X2=2.365 $Y2=1.725
r40 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.56
+ $X2=2.365 $Y2=1.395
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=1.56 $X2=2.365 $Y2=1.56
r42 10 15 2.73018 $w=4.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.495 $Y=1.665
+ $X2=2.495 $Y2=1.56
r43 9 15 6.89045 $w=4.58e-07 $l=2.65e-07 $layer=LI1_cond $X=2.495 $Y=1.295
+ $X2=2.495 $Y2=1.56
r44 7 16 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.355 $Y=0.625
+ $X2=2.355 $Y2=1.395
r45 3 17 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.325 $Y=2.595
+ $X2=2.325 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%B1 1 3 6 10 11 12 16
c28 11 0 2.28059e-20 $X=3.12 $Y=1.295
r29 16 19 36.9161 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.942 $Y=1.56
+ $X2=2.942 $Y2=1.725
r30 16 18 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.942 $Y=1.56
+ $X2=2.942 $Y2=1.395
r31 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=1.56 $X2=2.98 $Y2=1.56
r32 12 17 3.31525 $w=3.63e-07 $l=1.05e-07 $layer=LI1_cond $X=3.077 $Y=1.665
+ $X2=3.077 $Y2=1.56
r33 11 17 8.36705 $w=3.63e-07 $l=2.65e-07 $layer=LI1_cond $X=3.077 $Y=1.295
+ $X2=3.077 $Y2=1.56
r34 10 19 79.5785 $w=2e-07 $l=2.4e-07 $layer=POLY_cond $X=2.84 $Y=1.965 $X2=2.84
+ $Y2=1.725
r35 6 18 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.815 $Y=0.625
+ $X2=2.815 $Y2=1.395
r36 1 10 33.72 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.815 $Y=2.09
+ $X2=2.815 $Y2=1.965
r37 1 3 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.815 $Y=2.09
+ $X2=2.815 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%VPWR 1 2 3 10 12 18 20 22 27 28 29 35 47
r44 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r49 35 46 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r50 35 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 34 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 31 43 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.245 $Y2=3.33
r54 31 33 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.49 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 29 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 29 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 29 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 27 33 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.23 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=3.33
+ $X2=1.395 $Y2=3.33
r60 26 37 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.395 $Y2=3.33
r62 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.08 $Y=2.24 $X2=3.08
+ $Y2=2.95
r63 20 46 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r64 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.95
r65 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=3.245
+ $X2=1.395 $Y2=3.33
r66 16 18 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=1.395 $Y=3.245
+ $X2=1.395 $Y2=2.28
r67 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.325 $Y=2.24
+ $X2=0.325 $Y2=2.95
r68 10 43 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.325 $Y=3.245
+ $X2=0.245 $Y2=3.33
r69 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.325 $Y=3.245
+ $X2=0.325 $Y2=2.95
r70 3 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=2.095 $X2=3.08 $Y2=2.95
r71 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=2.095 $X2=3.08 $Y2=2.24
r72 2 18 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=1.255
+ $Y=2.095 $X2=1.395 $Y2=2.28
r73 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=2.095 $X2=0.325 $Y2=2.95
r74 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=2.095 $X2=0.325 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%Y 1 2 9 16 18 19 20
r41 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=0.555
+ $X2=1.71 $Y2=0.925
r42 14 20 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.71 $Y=1.255
+ $X2=1.71 $Y2=0.925
r43 14 16 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.71 $Y=1.34 $X2=2.01
+ $Y2=1.34
r44 11 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=1.425
+ $X2=2.01 $Y2=1.34
r45 11 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.01 $Y=1.425
+ $X2=2.01 $Y2=2.115
r46 9 18 7.72582 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=2.28
+ $X2=2.06 $Y2=2.115
r47 2 9 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=2.095 $X2=2.06 $Y2=2.28
r48 1 19 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.415 $X2=1.71 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%VGND 1 2 7 9 13 15 17 27 28 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r40 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.57
+ $Y2=0
r42 25 27 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=3.12
+ $Y2=0
r43 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r44 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r45 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r46 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r47 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 18 31 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r49 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r50 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.57
+ $Y2=0
r51 17 23 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.16
+ $Y2=0
r52 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r53 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r54 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0
r55 11 13 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0.56
r56 7 31 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r57 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.495
r58 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.415 $X2=2.57 $Y2=0.56
r59 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_LP%A_400_83# 1 2 9 11 12 15
c22 9 0 2.63001e-19 $X=2.14 $Y=0.625
r23 13 15 9.05491 $w=2.78e-07 $l=2.2e-07 $layer=LI1_cond $X=3.055 $Y=0.845
+ $X2=3.055 $Y2=0.625
r24 11 13 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.915 $Y=0.93
+ $X2=3.055 $Y2=0.845
r25 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.915 $Y=0.93
+ $X2=2.225 $Y2=0.93
r26 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=0.845
+ $X2=2.225 $Y2=0.93
r27 7 9 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.14 $Y=0.845 $X2=2.14
+ $Y2=0.625
r28 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.415 $X2=3.03 $Y2=0.625
r29 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.415
+ $X2=2.14 $Y2=0.625
.ends

