* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or3b_m A B C_N VGND VNB VPB VPWR X
X0 a_371_418# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_212_418# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR C_N a_112_55# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_212_418# a_112_55# a_299_418# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND C_N a_112_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_212_418# a_112_55# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_299_418# B a_371_418# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND B a_212_418# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_212_418# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_212_418# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
