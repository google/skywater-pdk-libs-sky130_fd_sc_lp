* File: sky130_fd_sc_lp__o31ai_lp.pxi.spice
* Created: Fri Aug 28 11:16:45 2020
* 
x_PM_SKY130_FD_SC_LP__O31AI_LP%A1 N_A1_c_56_n N_A1_M1003_g N_A1_c_57_n
+ N_A1_M1000_g N_A1_c_58_n A1 A1 N_A1_c_59_n N_A1_c_60_n N_A1_c_61_n
+ PM_SKY130_FD_SC_LP__O31AI_LP%A1
x_PM_SKY130_FD_SC_LP__O31AI_LP%A2 N_A2_M1006_g N_A2_M1001_g N_A2_c_94_n
+ N_A2_c_99_n A2 A2 A2 A2 N_A2_c_95_n N_A2_c_96_n
+ PM_SKY130_FD_SC_LP__O31AI_LP%A2
x_PM_SKY130_FD_SC_LP__O31AI_LP%A3 N_A3_M1004_g N_A3_M1002_g N_A3_c_143_n
+ N_A3_c_148_n A3 N_A3_c_144_n N_A3_c_145_n PM_SKY130_FD_SC_LP__O31AI_LP%A3
x_PM_SKY130_FD_SC_LP__O31AI_LP%B1 N_B1_M1005_g N_B1_M1007_g N_B1_c_184_n
+ N_B1_c_189_n B1 N_B1_c_185_n N_B1_c_186_n PM_SKY130_FD_SC_LP__O31AI_LP%B1
x_PM_SKY130_FD_SC_LP__O31AI_LP%VPWR N_VPWR_M1003_s N_VPWR_M1005_d N_VPWR_c_220_n
+ N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_223_n VPWR N_VPWR_c_224_n
+ N_VPWR_c_219_n PM_SKY130_FD_SC_LP__O31AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O31AI_LP%Y N_Y_M1007_d N_Y_M1004_d N_Y_c_261_n N_Y_c_257_n
+ N_Y_c_258_n Y Y Y N_Y_c_275_n N_Y_c_260_n PM_SKY130_FD_SC_LP__O31AI_LP%Y
x_PM_SKY130_FD_SC_LP__O31AI_LP%VGND N_VGND_M1000_s N_VGND_M1001_d N_VGND_c_293_n
+ N_VGND_c_294_n N_VGND_c_295_n N_VGND_c_296_n N_VGND_c_297_n VGND
+ N_VGND_c_298_n N_VGND_c_299_n PM_SKY130_FD_SC_LP__O31AI_LP%VGND
x_PM_SKY130_FD_SC_LP__O31AI_LP%A_161_57# N_A_161_57#_M1000_d N_A_161_57#_M1002_d
+ N_A_161_57#_c_326_n N_A_161_57#_c_327_n N_A_161_57#_c_328_n
+ N_A_161_57#_c_329_n PM_SKY130_FD_SC_LP__O31AI_LP%A_161_57#
cc_1 VNB N_A1_c_56_n 0.0321528f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.598
cc_2 VNB N_A1_c_57_n 0.0180612f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.78
cc_3 VNB N_A1_c_58_n 0.0323395f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.855
cc_4 VNB N_A1_c_59_n 0.0231942f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_5 VNB N_A1_c_60_n 0.0289938f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_6 VNB N_A1_c_61_n 0.0158341f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.11
cc_7 VNB N_A2_M1001_g 0.0442255f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_8 VNB N_A2_c_94_n 0.0153076f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.495
cc_9 VNB N_A2_c_95_n 0.0163843f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_10 VNB N_A2_c_96_n 0.00487884f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.11
cc_11 VNB N_A3_M1002_g 0.0397086f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_12 VNB N_A3_c_143_n 0.018654f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.495
cc_13 VNB N_A3_c_144_n 0.0168076f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_A3_c_145_n 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_B1_M1007_g 0.0425181f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_16 VNB N_B1_c_184_n 0.018764f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.495
cc_17 VNB N_B1_c_185_n 0.0168363f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_B1_c_186_n 0.00696084f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_VPWR_c_219_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_257_n 0.0458341f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.855
cc_21 VNB N_Y_c_258_n 0.0327835f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_VGND_c_293_n 0.017161f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_23 VNB N_VGND_c_294_n 0.028311f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.78
cc_24 VNB N_VGND_c_295_n 0.00712794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_296_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_VGND_c_297_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_27 VNB N_VGND_c_298_n 0.035112f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_28 VNB N_VGND_c_299_n 0.191111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_161_57#_c_326_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.78
cc_30 VNB N_A_161_57#_c_327_n 0.0249195f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.495
cc_31 VNB N_A_161_57#_c_328_n 0.00836148f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.855
cc_32 VNB N_A_161_57#_c_329_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A1_c_56_n 0.0345284f $X=-0.19 $Y=1.655 $X2=0.402 $Y2=1.598
cc_34 VPB N_A1_M1003_g 0.0343426f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.595
cc_35 VPB N_A1_c_60_n 0.0085352f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_36 VPB N_A2_M1006_g 0.0248978f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.93
cc_37 VPB N_A2_c_94_n 0.00779048f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.495
cc_38 VPB N_A2_c_99_n 0.0129824f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.855
cc_39 VPB N_A2_c_96_n 0.0035599f $X=-0.19 $Y=1.655 $X2=0.402 $Y2=1.11
cc_40 VPB N_A3_M1004_g 0.0292328f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.93
cc_41 VPB N_A3_c_143_n 0.00522878f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.495
cc_42 VPB N_A3_c_148_n 0.0139133f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.855
cc_43 VPB N_A3_c_145_n 7.54819e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_44 VPB N_B1_M1005_g 0.031908f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.93
cc_45 VPB N_B1_c_184_n 0.0052596f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.495
cc_46 VPB N_B1_c_189_n 0.0139824f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.855
cc_47 VPB N_B1_c_186_n 0.00287156f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_48 VPB N_VPWR_c_220_n 0.0113538f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.595
cc_49 VPB N_VPWR_c_221_n 0.0441418f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.78
cc_50 VPB N_VPWR_c_222_n 0.0156047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_223_n 0.0177824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_224_n 0.0490575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_219_n 0.0479482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_Y_c_257_n 0.0426619f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.855
cc_55 VPB N_Y_c_260_n 0.00977147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 N_A1_M1003_g N_A2_M1006_g 0.0395702f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_57 N_A1_c_57_n N_A2_M1001_g 0.0177653f $X=0.73 $Y=0.78 $X2=0 $Y2=0
cc_58 N_A1_c_60_n N_A2_M1001_g 7.77674e-19 $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_59 N_A1_c_61_n N_A2_M1001_g 0.0080462f $X=0.402 $Y=1.11 $X2=0 $Y2=0
cc_60 N_A1_c_56_n N_A2_c_94_n 0.00881488f $X=0.402 $Y=1.598 $X2=0 $Y2=0
cc_61 N_A1_c_56_n N_A2_c_99_n 0.0395702f $X=0.402 $Y=1.598 $X2=0 $Y2=0
cc_62 N_A1_c_59_n N_A2_c_95_n 0.00881488f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_63 N_A1_c_60_n N_A2_c_95_n 0.00198874f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_64 N_A1_c_56_n N_A2_c_96_n 0.0052472f $X=0.402 $Y=1.598 $X2=0 $Y2=0
cc_65 N_A1_c_59_n N_A2_c_96_n 0.0021714f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_66 N_A1_c_60_n N_A2_c_96_n 0.0210479f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_67 N_A1_c_56_n N_VPWR_c_221_n 0.00157747f $X=0.402 $Y=1.598 $X2=0 $Y2=0
cc_68 N_A1_M1003_g N_VPWR_c_221_n 0.0260828f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_69 N_A1_c_60_n N_VPWR_c_221_n 0.019625f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_70 N_A1_M1003_g N_VPWR_c_224_n 0.008763f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_71 N_A1_M1003_g N_VPWR_c_219_n 0.0144563f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_72 N_A1_c_57_n N_VGND_c_294_n 0.0128977f $X=0.73 $Y=0.78 $X2=0 $Y2=0
cc_73 N_A1_c_58_n N_VGND_c_294_n 0.00665822f $X=0.73 $Y=0.855 $X2=0 $Y2=0
cc_74 N_A1_c_59_n N_VGND_c_294_n 0.00115583f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_75 N_A1_c_60_n N_VGND_c_294_n 0.0133998f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_76 N_A1_c_57_n N_VGND_c_296_n 0.00502664f $X=0.73 $Y=0.78 $X2=0 $Y2=0
cc_77 N_A1_c_58_n N_VGND_c_296_n 8.33978e-19 $X=0.73 $Y=0.855 $X2=0 $Y2=0
cc_78 N_A1_c_57_n N_VGND_c_299_n 0.0101981f $X=0.73 $Y=0.78 $X2=0 $Y2=0
cc_79 N_A1_c_58_n N_VGND_c_299_n 0.00118182f $X=0.73 $Y=0.855 $X2=0 $Y2=0
cc_80 N_A1_c_57_n N_A_161_57#_c_326_n 0.00900602f $X=0.73 $Y=0.78 $X2=0 $Y2=0
cc_81 N_A1_c_58_n N_A_161_57#_c_326_n 0.00542796f $X=0.73 $Y=0.855 $X2=0 $Y2=0
cc_82 N_A1_c_58_n N_A_161_57#_c_328_n 0.00380327f $X=0.73 $Y=0.855 $X2=0 $Y2=0
cc_83 N_A1_c_61_n N_A_161_57#_c_328_n 0.00330698f $X=0.402 $Y=1.11 $X2=0 $Y2=0
cc_84 N_A2_M1006_g N_A3_M1004_g 0.0482007f $X=1.05 $Y=2.595 $X2=0 $Y2=0
cc_85 N_A2_M1001_g N_A3_M1002_g 0.0250107f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_86 N_A2_c_94_n N_A3_c_143_n 0.0117303f $X=1.09 $Y=1.77 $X2=0 $Y2=0
cc_87 N_A2_c_99_n N_A3_c_148_n 0.0117303f $X=1.09 $Y=1.935 $X2=0 $Y2=0
cc_88 N_A2_M1001_g N_A3_c_144_n 0.00203617f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A2_c_95_n N_A3_c_144_n 0.0117303f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_90 N_A2_c_96_n N_A3_c_144_n 0.0147058f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_91 N_A2_M1001_g N_A3_c_145_n 2.52145e-19 $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_92 N_A2_c_95_n N_A3_c_145_n 7.11149e-19 $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_93 N_A2_c_96_n N_A3_c_145_n 0.0483352f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_94 N_A2_M1006_g N_VPWR_c_221_n 0.00382854f $X=1.05 $Y=2.595 $X2=0 $Y2=0
cc_95 N_A2_c_96_n N_VPWR_c_221_n 0.027363f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_96 N_A2_M1006_g N_VPWR_c_224_n 0.00656883f $X=1.05 $Y=2.595 $X2=0 $Y2=0
cc_97 N_A2_c_96_n N_VPWR_c_224_n 0.0110411f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_98 N_A2_M1006_g N_VPWR_c_219_n 0.00824494f $X=1.05 $Y=2.595 $X2=0 $Y2=0
cc_99 N_A2_c_96_n N_VPWR_c_219_n 0.0122875f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_100 N_A2_c_96_n A_235_419# 0.00912939f $X=1.09 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_101 N_A2_M1006_g N_Y_c_261_n 9.77151e-19 $X=1.05 $Y=2.595 $X2=0 $Y2=0
cc_102 N_A2_M1006_g N_Y_c_260_n 7.68855e-19 $X=1.05 $Y=2.595 $X2=0 $Y2=0
cc_103 N_A2_c_96_n N_Y_c_260_n 0.0490535f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_104 N_A2_M1001_g N_VGND_c_295_n 0.00541719f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_105 N_A2_M1001_g N_VGND_c_296_n 0.00502664f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_106 N_A2_M1001_g N_VGND_c_299_n 0.00968694f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_107 N_A2_M1001_g N_A_161_57#_c_326_n 0.0110106f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_108 N_A2_M1001_g N_A_161_57#_c_327_n 0.0121208f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_109 N_A2_c_96_n N_A_161_57#_c_327_n 0.0131837f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_110 N_A2_M1001_g N_A_161_57#_c_328_n 0.00313634f $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_111 N_A2_c_95_n N_A_161_57#_c_328_n 0.00120613f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_112 N_A2_c_96_n N_A_161_57#_c_328_n 0.0133857f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_113 N_A2_M1001_g N_A_161_57#_c_329_n 8.96792e-19 $X=1.16 $Y=0.495 $X2=0 $Y2=0
cc_114 N_A3_M1004_g N_B1_M1005_g 0.0247502f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_115 N_A3_M1002_g N_B1_M1007_g 0.0321124f $X=1.75 $Y=0.495 $X2=0 $Y2=0
cc_116 N_A3_c_143_n N_B1_c_184_n 0.01184f $X=1.66 $Y=1.73 $X2=0 $Y2=0
cc_117 N_A3_c_148_n N_B1_c_189_n 0.01184f $X=1.66 $Y=1.895 $X2=0 $Y2=0
cc_118 N_A3_c_144_n N_B1_c_185_n 0.01184f $X=1.66 $Y=1.39 $X2=0 $Y2=0
cc_119 N_A3_c_145_n N_B1_c_185_n 8.23261e-19 $X=1.66 $Y=1.39 $X2=0 $Y2=0
cc_120 N_A3_c_144_n N_B1_c_186_n 0.00410205f $X=1.66 $Y=1.39 $X2=0 $Y2=0
cc_121 N_A3_c_145_n N_B1_c_186_n 0.0438819f $X=1.66 $Y=1.39 $X2=0 $Y2=0
cc_122 N_A3_M1004_g N_VPWR_c_223_n 9.89243e-19 $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_123 N_A3_M1004_g N_VPWR_c_224_n 0.00706392f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_124 N_A3_M1004_g N_VPWR_c_219_n 0.0107145f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_125 N_A3_M1004_g N_Y_c_261_n 0.018774f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_126 N_A3_M1004_g N_Y_c_260_n 0.0150235f $X=1.62 $Y=2.595 $X2=0 $Y2=0
cc_127 N_A3_c_148_n N_Y_c_260_n 6.13398e-19 $X=1.66 $Y=1.895 $X2=0 $Y2=0
cc_128 N_A3_c_145_n N_Y_c_260_n 0.0211858f $X=1.66 $Y=1.39 $X2=0 $Y2=0
cc_129 N_A3_M1002_g N_VGND_c_295_n 0.00541719f $X=1.75 $Y=0.495 $X2=0 $Y2=0
cc_130 N_A3_M1002_g N_VGND_c_298_n 0.00502664f $X=1.75 $Y=0.495 $X2=0 $Y2=0
cc_131 N_A3_M1002_g N_VGND_c_299_n 0.00968694f $X=1.75 $Y=0.495 $X2=0 $Y2=0
cc_132 N_A3_M1002_g N_A_161_57#_c_326_n 8.96792e-19 $X=1.75 $Y=0.495 $X2=0 $Y2=0
cc_133 N_A3_M1002_g N_A_161_57#_c_327_n 0.014665f $X=1.75 $Y=0.495 $X2=0 $Y2=0
cc_134 N_A3_c_144_n N_A_161_57#_c_327_n 0.00122995f $X=1.66 $Y=1.39 $X2=0 $Y2=0
cc_135 N_A3_c_145_n N_A_161_57#_c_327_n 0.0246663f $X=1.66 $Y=1.39 $X2=0 $Y2=0
cc_136 N_A3_M1002_g N_A_161_57#_c_329_n 0.0109989f $X=1.75 $Y=0.495 $X2=0 $Y2=0
cc_137 N_B1_M1005_g N_VPWR_c_223_n 0.0124068f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_138 N_B1_M1005_g N_VPWR_c_224_n 0.008763f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_139 N_B1_M1005_g N_VPWR_c_219_n 0.00776649f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_140 N_B1_M1005_g N_Y_c_257_n 0.0105891f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_141 N_B1_M1007_g N_Y_c_257_n 0.0109907f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_142 N_B1_c_185_n N_Y_c_257_n 0.0147882f $X=2.23 $Y=1.39 $X2=0 $Y2=0
cc_143 N_B1_c_186_n N_Y_c_257_n 0.0464518f $X=2.23 $Y=1.39 $X2=0 $Y2=0
cc_144 N_B1_M1007_g N_Y_c_258_n 0.00891389f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_145 N_B1_c_185_n N_Y_c_258_n 5.2181e-19 $X=2.23 $Y=1.39 $X2=0 $Y2=0
cc_146 N_B1_c_186_n N_Y_c_258_n 0.00320476f $X=2.23 $Y=1.39 $X2=0 $Y2=0
cc_147 N_B1_M1005_g N_Y_c_275_n 0.0220219f $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_148 N_B1_c_189_n N_Y_c_275_n 2.87537e-19 $X=2.23 $Y=1.895 $X2=0 $Y2=0
cc_149 N_B1_c_186_n N_Y_c_275_n 0.0123265f $X=2.23 $Y=1.39 $X2=0 $Y2=0
cc_150 N_B1_M1005_g N_Y_c_260_n 3.10204e-19 $X=2.19 $Y=2.595 $X2=0 $Y2=0
cc_151 N_B1_M1007_g N_VGND_c_298_n 0.00502664f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_152 N_B1_M1007_g N_VGND_c_299_n 0.0103089f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_153 N_B1_M1007_g N_A_161_57#_c_327_n 0.00540618f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_154 N_B1_c_185_n N_A_161_57#_c_327_n 3.10581e-19 $X=2.23 $Y=1.39 $X2=0 $Y2=0
cc_155 N_B1_c_186_n N_A_161_57#_c_327_n 0.00713614f $X=2.23 $Y=1.39 $X2=0 $Y2=0
cc_156 N_B1_M1007_g N_A_161_57#_c_329_n 0.0104064f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_157 N_VPWR_c_219_n A_137_419# 0.010279f $X=2.64 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_158 N_VPWR_c_219_n A_235_419# 0.00902063f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_159 N_VPWR_c_219_n N_Y_M1004_d 0.00263863f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_224_n N_Y_c_261_n 0.0283111f $X=2.29 $Y=3.33 $X2=0 $Y2=0
cc_161 N_VPWR_c_219_n N_Y_c_261_n 0.0177915f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VPWR_M1005_d N_Y_c_257_n 0.00304367f $X=2.315 $Y=2.095 $X2=0 $Y2=0
cc_163 N_VPWR_c_223_n N_Y_c_257_n 0.00287998f $X=2.455 $Y=2.905 $X2=0 $Y2=0
cc_164 N_VPWR_c_219_n N_Y_c_257_n 0.00561607f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_M1005_d N_Y_c_275_n 0.0112253f $X=2.315 $Y=2.095 $X2=0 $Y2=0
cc_166 N_VPWR_c_223_n N_Y_c_275_n 0.0182202f $X=2.455 $Y=2.905 $X2=0 $Y2=0
cc_167 N_VPWR_c_219_n N_Y_c_275_n 0.00810308f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_168 N_Y_c_258_n N_VGND_c_298_n 0.0289609f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_169 N_Y_c_258_n N_VGND_c_299_n 0.0170302f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_170 N_Y_c_257_n N_A_161_57#_c_327_n 0.00645337f $X=2.67 $Y=2.29 $X2=0 $Y2=0
cc_171 N_Y_c_257_n N_A_161_57#_c_329_n 0.00537021f $X=2.67 $Y=2.29 $X2=0 $Y2=0
cc_172 N_Y_c_258_n N_A_161_57#_c_329_n 0.0180007f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_173 N_VGND_c_294_n N_A_161_57#_c_326_n 0.0180055f $X=0.435 $Y=0.495 $X2=0
+ $Y2=0
cc_174 N_VGND_c_295_n N_A_161_57#_c_326_n 0.016171f $X=1.455 $Y=0.48 $X2=0 $Y2=0
cc_175 N_VGND_c_296_n N_A_161_57#_c_326_n 0.021949f $X=1.29 $Y=0 $X2=0 $Y2=0
cc_176 N_VGND_c_299_n N_A_161_57#_c_326_n 0.0124703f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_177 N_VGND_c_295_n N_A_161_57#_c_327_n 0.0259275f $X=1.455 $Y=0.48 $X2=0
+ $Y2=0
cc_178 N_VGND_c_295_n N_A_161_57#_c_329_n 0.016171f $X=1.455 $Y=0.48 $X2=0 $Y2=0
cc_179 N_VGND_c_298_n N_A_161_57#_c_329_n 0.021949f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_180 N_VGND_c_299_n N_A_161_57#_c_329_n 0.0124703f $X=2.64 $Y=0 $X2=0 $Y2=0
