* File: sky130_fd_sc_lp__xnor3_1.spice
* Created: Fri Aug 28 11:35:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor3_1.pex.spice"
.subckt sky130_fd_sc_lp__xnor3_1  VNB VPB C B A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_A_81_259#_M1019_g N_X_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2767 AS=0.2352 PD=1.96667 PS=2.24 NRD=16.428 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1006 N_A_244_137#_M1006_d N_C_M1006_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.13835 PD=1.4 PS=0.983333 NRD=0 NRS=78.396 M=1 R=2.8 SA=75000.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_81_259#_M1010_d N_C_M1010_g N_A_354_109#_M1010_s VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.1792 PD=0.99 PS=1.84 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1009 N_A_355_451#_M1009_d N_A_244_137#_M1009_g N_A_81_259#_M1010_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1002 N_A_754_367#_M1002_d N_B_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.3737 PD=2.25 PS=2.74 NRD=0 NRS=17.136 M=1 R=5.6 SA=75000.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_354_109#_M1000_d N_A_754_367#_M1000_g N_A_871_373#_M1000_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.112 AS=0.3749 PD=0.99 PS=2.9 NRD=0 NRS=99.516 M=1 R=4.26667
+ SA=75000.3 SB=75002 A=0.096 P=1.58 MULT=1
MM1004 N_A_1090_373#_M1004_d N_B_M1004_g N_A_354_109#_M1000_d VNB NSHORT L=0.15
+ W=0.64 AD=0.141826 AS=0.112 PD=1.30415 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.8 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1001 N_A_355_451#_M1001_d N_A_754_367#_M1001_g N_A_1090_373#_M1004_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.101989 AS=0.0930736 PD=0.855849 PS=0.855849
+ NRD=32.856 NRS=47.592 M=1 R=2.8 SA=75001.2 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1007 N_A_871_373#_M1007_d N_B_M1007_g N_A_355_451#_M1001_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0976 AS=0.155411 PD=0.945 PS=1.30415 NRD=4.68 NRS=8.436 M=1
+ R=4.26667 SA=75001.3 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_871_373#_M1007_d VNB NSHORT L=0.15 W=0.64
+ AD=0.16 AS=0.0976 PD=1.14 PS=0.945 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1015 N_A_1090_373#_M1015_d N_A_871_373#_M1015_g N_VGND_M1003_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.16 PD=1.85 PS=1.14 NRD=0 NRS=28.116 M=1 R=4.26667
+ SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_VPWR_M1020_d N_A_81_259#_M1020_g N_X_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.342123 AS=0.3402 PD=2.37411 PS=3.06 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.5 A=0.189 P=2.82 MULT=1
MM1014 N_A_244_137#_M1014_d N_C_M1014_g N_VPWR_M1020_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1728 AS=0.173777 PD=1.82 PS=1.20589 NRD=0 NRS=78.4848 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_A_81_259#_M1011_d N_C_M1011_g N_A_355_451#_M1011_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1806 AS=0.231 PD=1.445 PS=2.23 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1016 N_A_354_109#_M1016_d N_A_244_137#_M1016_g N_A_81_259#_M1011_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2688 AS=0.1806 PD=2.32 PS=1.445 NRD=0 NRS=37.5088 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_A_754_367#_M1021_d N_B_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.3591 PD=3.09 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1012 N_A_355_451#_M1012_d N_A_754_367#_M1012_g N_A_871_373#_M1012_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.175832 AS=0.40415 PD=1.40189 PS=2.95 NRD=0
+ NRS=99.9184 M=1 R=5.6 SA=75000.3 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1017 N_A_1090_373#_M1017_d N_B_M1017_g N_A_355_451#_M1012_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.133968 PD=0.92 PS=1.06811 NRD=0 NRS=89.2607 M=1
+ R=4.26667 SA=75000.9 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1008 N_A_354_109#_M1008_d N_A_754_367#_M1008_g N_A_1090_373#_M1017_d VPB
+ PHIGHVT L=0.15 W=0.64 AD=0.158616 AS=0.0896 PD=1.15459 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001.3 SB=75002 A=0.096 P=1.58 MULT=1
MM1013 N_A_871_373#_M1013_d N_B_M1013_g N_A_354_109#_M1008_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.231411 AS=0.208184 PD=1.42435 PS=1.51541 NRD=27.3436 NRS=50.4123
+ M=1 R=5.6 SA=75001.5 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g N_A_871_373#_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1925 AS=0.275489 PD=1.385 PS=1.69565 NRD=0 NRS=22.6353 M=1 R=6.66667
+ SA=75001.8 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1005 N_A_1090_373#_M1005_d N_A_871_373#_M1005_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.285 AS=0.1925 PD=2.57 PS=1.385 NRD=0 NRS=20.685 M=1 R=6.66667
+ SA=75002.3 SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.9271 P=20.81
c_157 VPB 0 1.36914e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__xnor3_1.pxi.spice"
*
.ends
*
*
