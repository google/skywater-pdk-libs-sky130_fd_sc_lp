* File: sky130_fd_sc_lp__nor4_2.pex.spice
* Created: Fri Aug 28 10:57:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4_2%B 3 7 11 15 17 18 19 22 23 27 28 47
c80 22 0 1.30739e-19 $X=2.02 $Y=1.51
c81 15 0 1.2912e-19 $X=2 $Y=2.465
r82 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.51 $X2=0.385 $Y2=1.51
r83 28 47 8.04956 $w=4.38e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.855 $Y2=1.565
r84 28 34 5.85063 $w=6.08e-07 $l=2.5e-07 $layer=LI1_cond $X=0.635 $Y=1.565
+ $X2=0.385 $Y2=1.565
r85 27 34 3.79782 $w=4.38e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.385 $Y2=1.565
r86 23 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.02 $Y=1.51
+ $X2=2.02 $Y2=1.675
r87 23 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.02 $Y=1.51
+ $X2=2.02 $Y2=1.345
r88 22 25 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.02 $Y=1.51
+ $X2=2.02 $Y2=1.7
r89 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.02
+ $Y=1.51 $X2=2.02 $Y2=1.51
r90 19 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=1.7
+ $X2=2.02 $Y2=1.7
r91 19 47 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.855 $Y=1.7 $X2=0.855
+ $Y2=1.7
r92 17 33 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.635 $Y=1.51
+ $X2=0.385 $Y2=1.51
r93 17 18 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.635 $Y=1.51
+ $X2=0.71 $Y2=1.51
r94 15 38 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2 $Y=2.465 $X2=2
+ $Y2=1.675
r95 11 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2 $Y=0.655 $X2=2
+ $Y2=1.345
r96 5 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.71 $Y=1.675
+ $X2=0.71 $Y2=1.51
r97 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.71 $Y=1.675 $X2=0.71
+ $Y2=2.465
r98 1 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.71 $Y=1.345
+ $X2=0.71 $Y2=1.51
r99 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.71 $Y=1.345 $X2=0.71
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%A 1 3 6 8 10 13 15 22
c50 13 0 1.30739e-19 $X=1.57 $Y=2.465
c51 8 0 1.00299e-19 $X=1.57 $Y=1.185
r52 20 22 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.285 $Y=1.35
+ $X2=1.57 $Y2=1.35
r53 17 20 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.14 $Y=1.35
+ $X2=1.285 $Y2=1.35
r54 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.285
+ $Y=1.35 $X2=1.285 $Y2=1.35
r55 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.515
+ $X2=1.57 $Y2=1.35
r56 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.57 $Y=1.515
+ $X2=1.57 $Y2=2.465
r57 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.185
+ $X2=1.57 $Y2=1.35
r58 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.57 $Y=1.185
+ $X2=1.57 $Y2=0.655
r59 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.515
+ $X2=1.14 $Y2=1.35
r60 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.14 $Y=1.515 $X2=1.14
+ $Y2=2.465
r61 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.185
+ $X2=1.14 $Y2=1.35
r62 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.14 $Y=1.185 $X2=1.14
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%C 3 7 11 15 20 21 25 26 34 45
c94 34 0 3.94798e-20 $X=4 $Y=1.51
c95 3 0 7.67244e-20 $X=2.62 $Y=0.655
r96 34 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=1.51 $X2=4
+ $Y2=1.675
r97 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=1.51 $X2=4
+ $Y2=1.345
r98 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4 $Y=1.51
+ $X2=4 $Y2=1.51
r99 26 35 2.09535 $w=4.38e-07 $l=8e-08 $layer=LI1_cond $X=4.08 $Y=1.645 $X2=4
+ $Y2=1.645
r100 25 45 8.04956 $w=4.38e-07 $l=1.35e-07 $layer=LI1_cond $X=3.6 $Y=1.645
+ $X2=3.465 $Y2=1.645
r101 25 35 7.12514 $w=6.08e-07 $l=3.15e-07 $layer=LI1_cond $X=3.685 $Y=1.645
+ $X2=4 $Y2=1.645
r102 21 32 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.51
+ $X2=2.58 $Y2=1.675
r103 21 31 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.51
+ $X2=2.58 $Y2=1.345
r104 20 23 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.56 $Y=1.51
+ $X2=2.56 $Y2=1.78
r105 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.51 $X2=2.56 $Y2=1.51
r106 18 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.78
+ $X2=2.56 $Y2=1.78
r107 18 45 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.725 $Y=1.78
+ $X2=3.465 $Y2=1.78
r108 15 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.98 $Y=2.465
+ $X2=3.98 $Y2=1.675
r109 11 36 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.91 $Y=0.655
+ $X2=3.91 $Y2=1.345
r110 7 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.69 $Y=2.465
+ $X2=2.69 $Y2=1.675
r111 3 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.62 $Y=0.655
+ $X2=2.62 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%D 1 3 6 8 10 13 15 24
c54 15 0 3.94798e-20 $X=3.12 $Y=1.295
r55 23 24 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.48 $Y=1.35 $X2=3.55
+ $Y2=1.35
r56 21 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.14 $Y=1.35
+ $X2=3.48 $Y2=1.35
r57 19 21 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.12 $Y=1.35 $X2=3.14
+ $Y2=1.35
r58 17 19 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.05 $Y=1.35 $X2=3.12
+ $Y2=1.35
r59 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.14
+ $Y=1.35 $X2=3.14 $Y2=1.35
r60 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.515
+ $X2=3.55 $Y2=1.35
r61 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.55 $Y=1.515
+ $X2=3.55 $Y2=2.465
r62 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.185
+ $X2=3.48 $Y2=1.35
r63 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.48 $Y=1.185
+ $X2=3.48 $Y2=0.655
r64 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.515
+ $X2=3.12 $Y2=1.35
r65 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.12 $Y=1.515 $X2=3.12
+ $Y2=2.465
r66 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.185
+ $X2=3.05 $Y2=1.35
r67 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.05 $Y=1.185 $X2=3.05
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%A_74_367# 1 2 3 10 12 14 16 17 18 22
r50 20 22 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=4.23 $Y=2.905
+ $X2=4.23 $Y2=2.54
r51 19 29 6.34366 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=2.53 $Y=2.99
+ $X2=2.307 $Y2=2.99
r52 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.1 $Y=2.99
+ $X2=4.23 $Y2=2.905
r53 18 19 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=4.1 $Y=2.99
+ $X2=2.53 $Y2=2.99
r54 17 29 2.41799 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.307 $Y=2.905
+ $X2=2.307 $Y2=2.99
r55 16 27 2.42586 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.307 $Y=2.125
+ $X2=2.307 $Y2=2.04
r56 16 17 20.2001 $w=4.43e-07 $l=7.8e-07 $layer=LI1_cond $X=2.307 $Y=2.125
+ $X2=2.307 $Y2=2.905
r57 15 25 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.625 $Y=2.04
+ $X2=0.477 $Y2=2.04
r58 14 27 6.33579 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.085 $Y=2.04
+ $X2=2.307 $Y2=2.04
r59 14 15 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.085 $Y=2.04
+ $X2=0.625 $Y2=2.04
r60 10 25 2.72785 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.477 $Y=2.125
+ $X2=0.477 $Y2=2.04
r61 10 12 30.6667 $w=2.93e-07 $l=7.85e-07 $layer=LI1_cond $X=0.477 $Y=2.125
+ $X2=0.477 $Y2=2.91
r62 3 22 300 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_PDIFF $count=2 $X=4.055
+ $Y=1.835 $X2=4.195 $Y2=2.54
r63 2 29 400 $w=1.7e-07 $l=1.21135e-06 $layer=licon1_PDIFF $count=1 $X=2.075
+ $Y=1.835 $X2=2.365 $Y2=2.91
r64 2 27 400 $w=1.7e-07 $l=4.0835e-07 $layer=licon1_PDIFF $count=1 $X=2.075
+ $Y=1.835 $X2=2.365 $Y2=2.12
r65 1 25 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.37
+ $Y=1.835 $X2=0.495 $Y2=2.12
r66 1 12 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.37
+ $Y=1.835 $X2=0.495 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%A_157_367# 1 2 9 14 16
r15 10 14 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.02 $Y=2.38
+ $X2=0.907 $Y2=2.38
r16 9 16 3.9739 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.69 $Y=2.38 $X2=1.802
+ $Y2=2.38
r17 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.69 $Y=2.38 $X2=1.02
+ $Y2=2.38
r18 2 16 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=1.645
+ $Y=1.835 $X2=1.785 $Y2=2.46
r19 1 14 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=0.785
+ $Y=1.835 $X2=0.925 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%VPWR 1 6 8 10 20 21 24
r47 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 20 21 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 17 20 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 17 18 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.355 $Y2=3.33
r53 15 17 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 13 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=1.355 $Y2=3.33
r57 10 12 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 8 21 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.68
+ $Y2=3.33
r60 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=3.33
r61 4 6 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=2.76
r62 1 6 600 $w=1.7e-07 $l=9.92535e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.835 $X2=1.355 $Y2=2.76
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%A_553_367# 1 2 9 11 13
c22 9 0 1.2912e-19 $X=2.905 $Y=2.2
r23 11 13 38.3313 $w=2.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3 $Y=2.62 $X2=3.765
+ $Y2=2.62
r24 7 11 6.84978 $w=2.3e-07 $l=1.78466e-07 $layer=LI1_cond $X=2.87 $Y=2.505
+ $X2=3 $Y2=2.62
r25 7 9 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.87 $Y=2.505 $X2=2.87
+ $Y2=2.2
r26 2 13 600 $w=1.7e-07 $l=8.42096e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.835 $X2=3.765 $Y2=2.61
r27 1 9 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=2.765
+ $Y=1.835 $X2=2.905 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%Y 1 2 3 4 5 18 20 21 24 26 30 32 34 38 40 42
+ 46 51 54 58 59 60
c97 42 0 7.67244e-20 $X=1.785 $Y=0.955
c98 26 0 1.00299e-19 $X=2.65 $Y=1.17
r99 59 60 11.9635 $w=3.13e-07 $l=3.27e-07 $layer=LI1_cond $X=4.557 $Y=1.665
+ $X2=4.557 $Y2=1.992
r100 58 59 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=4.557 $Y=1.295
+ $X2=4.557 $Y2=1.665
r101 57 58 4.39026 $w=3.13e-07 $l=1.2e-07 $layer=LI1_cond $X=4.557 $Y=1.175
+ $X2=4.557 $Y2=1.295
r102 54 55 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=3.69 $Y=0.93
+ $X2=3.69 $Y2=1.09
r103 53 54 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=0.845
+ $X2=3.69 $Y2=0.93
r104 49 51 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=2.185
+ $X2=3.5 $Y2=2.185
r105 46 47 13.6186 $w=2.15e-07 $l=2.4e-07 $layer=LI1_cond $X=2.79 $Y=0.93
+ $X2=2.79 $Y2=1.17
r106 42 44 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.785 $Y=0.955
+ $X2=1.785 $Y2=1.17
r107 42 43 3.51899 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.955
+ $X2=1.785 $Y2=0.87
r108 41 55 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.79 $Y=1.09 $X2=3.69
+ $Y2=1.09
r109 40 57 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=4.4 $Y=1.09
+ $X2=4.557 $Y2=1.175
r110 40 41 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.4 $Y=1.09
+ $X2=3.79 $Y2=1.09
r111 38 53 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=3.695 $Y=0.42
+ $X2=3.695 $Y2=0.845
r112 34 60 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=4.4 $Y=2.12
+ $X2=4.557 $Y2=2.12
r113 34 51 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=4.4 $Y=2.12 $X2=3.5
+ $Y2=2.12
r114 33 46 2.11506 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.93 $Y=0.93
+ $X2=2.79 $Y2=0.93
r115 32 54 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.59 $Y=0.93 $X2=3.69
+ $Y2=0.93
r116 32 33 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.59 $Y=0.93
+ $X2=2.93 $Y2=0.93
r117 28 46 4.39198 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=0.845
+ $X2=2.79 $Y2=0.93
r118 28 30 17.4924 $w=2.78e-07 $l=4.25e-07 $layer=LI1_cond $X=2.79 $Y=0.845
+ $X2=2.79 $Y2=0.42
r119 27 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=1.17
+ $X2=1.785 $Y2=1.17
r120 26 47 2.11506 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.65 $Y=1.17
+ $X2=2.79 $Y2=1.17
r121 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.65 $Y=1.17 $X2=1.95
+ $Y2=1.17
r122 24 43 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=1.82 $Y=0.42
+ $X2=1.82 $Y2=0.87
r123 20 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0.955
+ $X2=1.785 $Y2=0.955
r124 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.62 $Y=0.955
+ $X2=1.01 $Y2=0.955
r125 16 21 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=0.902 $Y=0.87
+ $X2=1.01 $Y2=0.955
r126 16 18 23.5849 $w=2.13e-07 $l=4.4e-07 $layer=LI1_cond $X=0.902 $Y=0.87
+ $X2=0.902 $Y2=0.43
r127 5 49 600 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.835 $X2=3.335 $Y2=2.15
r128 4 54 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.235 $X2=3.695 $Y2=0.93
r129 4 38 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.235 $X2=3.695 $Y2=0.42
r130 3 30 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.695
+ $Y=0.235 $X2=2.835 $Y2=0.42
r131 2 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.645
+ $Y=0.235 $X2=1.785 $Y2=0.42
r132 1 18 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=0.785
+ $Y=0.235 $X2=0.925 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_2%VGND 1 2 3 4 5 18 20 24 26 30 32 36 40 42 43
+ 44 50 57 58 61 64 67 70
r72 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r73 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r74 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r75 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r76 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r77 58 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r78 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r79 55 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.125
+ $Y2=0
r80 55 57 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.56
+ $Y2=0
r81 54 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r82 54 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r83 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r84 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.265
+ $Y2=0
r85 51 53 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.6
+ $Y2=0
r86 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=4.125
+ $Y2=0
r87 50 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=3.6
+ $Y2=0
r88 48 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r89 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r90 44 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r91 44 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r92 42 47 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.33 $Y=0 $X2=0.24
+ $Y2=0
r93 42 43 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.33 $Y=0 $X2=0.477
+ $Y2=0
r94 38 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0.085
+ $X2=4.125 $Y2=0
r95 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.125 $Y=0.085
+ $X2=4.125 $Y2=0.38
r96 34 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=0.085
+ $X2=3.265 $Y2=0
r97 34 36 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.265 $Y=0.085
+ $X2=3.265 $Y2=0.55
r98 33 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.315
+ $Y2=0
r99 32 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.265
+ $Y2=0
r100 32 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.48
+ $Y2=0
r101 28 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=0.085
+ $X2=2.315 $Y2=0
r102 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.315 $Y=0.085
+ $X2=2.315 $Y2=0.38
r103 27 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.355
+ $Y2=0
r104 26 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.315
+ $Y2=0
r105 26 27 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=1.52
+ $Y2=0
r106 22 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=0.085
+ $X2=1.355 $Y2=0
r107 22 24 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.355 $Y=0.085
+ $X2=1.355 $Y2=0.575
r108 21 43 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.477 $Y2=0
r109 20 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=1.355
+ $Y2=0
r110 20 21 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=0.625
+ $Y2=0
r111 16 43 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.477 $Y=0.085
+ $X2=0.477 $Y2=0
r112 16 18 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.477 $Y=0.085
+ $X2=0.477 $Y2=0.38
r113 5 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.985
+ $Y=0.235 $X2=4.125 $Y2=0.38
r114 4 36 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.235 $X2=3.265 $Y2=0.55
r115 3 30 91 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=2 $X=2.075
+ $Y=0.235 $X2=2.315 $Y2=0.38
r116 2 24 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.235 $X2=1.355 $Y2=0.575
r117 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.37
+ $Y=0.235 $X2=0.495 $Y2=0.38
.ends

