# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 0.765000 2.280000 2.055000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.505000 0.265000 12.870000 1.095000 ;
        RECT 12.505000 1.815000 12.870000 3.065000 ;
        RECT 12.700000 1.095000 12.870000 1.815000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.010000 0.265000 11.445000 1.005000 ;
        RECT 11.085000 1.695000 11.445000 2.995000 ;
        RECT 11.275000 1.005000 11.445000 1.695000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.205000 1.180000 10.550000 1.515000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.375000 1.405000 4.705000 1.780000 ;
        RECT 4.375000 1.780000 4.675000 2.150000 ;
        RECT 8.265000 1.660000 8.560000 2.150000 ;
      LAYER mcon ;
        RECT 4.475000 1.950000 4.645000 2.120000 ;
        RECT 8.315000 1.950000 8.485000 2.120000 ;
      LAYER met1 ;
        RECT 4.415000 1.920000 4.705000 1.965000 ;
        RECT 4.415000 1.965000 8.545000 2.105000 ;
        RECT 4.415000 2.105000 4.705000 2.150000 ;
        RECT 8.255000 1.920000 8.545000 1.965000 ;
        RECT 8.255000 2.105000 8.545000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.905000 0.455000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.960000 0.085000 ;
        RECT  0.115000  0.085000  0.365000 0.725000 ;
        RECT  1.765000  0.085000  2.095000 0.585000 ;
        RECT  4.050000  0.085000  4.380000 0.875000 ;
        RECT  6.140000  0.085000  6.390000 0.580000 ;
        RECT  8.070000  0.085000  8.320000 0.765000 ;
        RECT 10.580000  0.085000 10.830000 1.000000 ;
        RECT 12.075000  0.085000 12.325000 0.935000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.960000 3.415000 ;
        RECT  0.185000 2.385000  0.515000 3.245000 ;
        RECT  1.765000 2.585000  2.095000 3.245000 ;
        RECT  4.265000 2.680000  4.595000 3.245000 ;
        RECT  5.595000 2.310000  5.925000 3.245000 ;
        RECT  8.140000 2.680000  8.470000 3.245000 ;
        RECT  9.500000 2.555000  9.830000 3.245000 ;
        RECT 10.575000 2.555000 10.905000 3.245000 ;
        RECT 12.075000 1.815000 12.325000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.545000 0.265000  0.875000 0.725000 ;
      RECT  0.695000 0.725000  0.875000 1.270000 ;
      RECT  0.695000 1.270000  1.025000 3.065000 ;
      RECT  1.105000 0.265000  1.585000 0.675000 ;
      RECT  1.255000 0.675000  1.585000 2.235000 ;
      RECT  1.255000 2.235000  2.630000 2.405000 ;
      RECT  1.255000 2.405000  1.585000 2.975000 ;
      RECT  2.460000 1.180000  2.755000 1.560000 ;
      RECT  2.460000 1.560000  3.000000 1.880000 ;
      RECT  2.460000 1.880000  2.630000 2.235000 ;
      RECT  2.630000 0.265000  2.960000 0.830000 ;
      RECT  2.630000 0.830000  3.350000 1.000000 ;
      RECT  2.810000 2.060000  3.350000 2.230000 ;
      RECT  2.810000 2.230000  3.140000 2.755000 ;
      RECT  3.140000 0.265000  3.470000 0.480000 ;
      RECT  3.140000 0.480000  3.700000 0.650000 ;
      RECT  3.180000 1.000000  3.350000 2.060000 ;
      RECT  3.320000 2.410000  3.700000 2.755000 ;
      RECT  3.530000 0.650000  3.700000 1.055000 ;
      RECT  3.530000 1.055000  5.200000 1.225000 ;
      RECT  3.530000 1.225000  3.700000 2.410000 ;
      RECT  3.880000 1.405000  4.165000 2.330000 ;
      RECT  3.880000 2.330000  5.105000 2.500000 ;
      RECT  4.560000 0.265000  5.910000 0.435000 ;
      RECT  4.560000 0.435000  4.890000 0.875000 ;
      RECT  4.855000 1.960000  6.555000 2.130000 ;
      RECT  4.855000 2.130000  5.105000 2.330000 ;
      RECT  4.855000 2.500000  5.105000 2.755000 ;
      RECT  4.915000 1.225000  5.200000 1.385000 ;
      RECT  5.070000 0.615000  5.400000 0.705000 ;
      RECT  5.070000 0.705000  5.550000 0.875000 ;
      RECT  5.380000 0.875000  5.550000 1.960000 ;
      RECT  5.580000 0.435000  5.910000 0.525000 ;
      RECT  5.730000 0.760000  6.740000 0.930000 ;
      RECT  5.730000 0.930000  6.015000 1.315000 ;
      RECT  6.225000 1.110000  6.555000 1.960000 ;
      RECT  6.570000 0.265000  7.835000 0.435000 ;
      RECT  6.570000 0.435000  6.740000 0.760000 ;
      RECT  6.640000 2.580000  7.585000 2.750000 ;
      RECT  6.640000 2.750000  6.970000 3.000000 ;
      RECT  6.805000 1.110000  7.135000 2.070000 ;
      RECT  6.805000 2.070000  7.235000 2.400000 ;
      RECT  6.960000 0.615000  7.485000 0.930000 ;
      RECT  7.315000 0.930000  7.485000 1.310000 ;
      RECT  7.315000 1.310000  8.910000 1.480000 ;
      RECT  7.415000 1.480000  7.585000 2.580000 ;
      RECT  7.665000 0.435000  7.835000 0.945000 ;
      RECT  7.665000 0.945000  8.910000 1.115000 ;
      RECT  7.765000 1.660000  8.055000 2.330000 ;
      RECT  7.765000 2.330000 10.905000 2.375000 ;
      RECT  7.765000 2.375000  8.990000 2.500000 ;
      RECT  8.500000 0.265000  9.845000 0.595000 ;
      RECT  8.740000 0.775000 10.400000 0.945000 ;
      RECT  8.740000 1.480000  8.910000 1.635000 ;
      RECT  8.740000 1.635000  9.135000 1.965000 ;
      RECT  8.740000 2.145000  9.485000 2.205000 ;
      RECT  8.740000 2.205000 10.905000 2.330000 ;
      RECT  8.740000 2.500000  8.990000 3.010000 ;
      RECT  9.090000 1.125000  9.485000 1.455000 ;
      RECT  9.315000 1.455000  9.485000 2.145000 ;
      RECT  9.680000 0.945000 10.400000 1.000000 ;
      RECT  9.680000 1.000000 10.010000 1.695000 ;
      RECT  9.680000 1.695000 10.395000 2.025000 ;
      RECT 10.070000 0.635000 10.400000 0.775000 ;
      RECT 10.735000 1.185000 11.095000 1.515000 ;
      RECT 10.735000 1.515000 10.905000 2.205000 ;
      RECT 11.645000 0.635000 11.895000 1.115000 ;
      RECT 11.645000 1.115000 12.325000 1.285000 ;
      RECT 11.645000 1.465000 12.520000 1.635000 ;
      RECT 11.645000 1.635000 11.895000 2.495000 ;
      RECT 12.155000 1.285000 12.325000 1.305000 ;
      RECT 12.155000 1.305000 12.520000 1.465000 ;
    LAYER mcon ;
      RECT 2.555000 1.210000 2.725000 1.380000 ;
      RECT 6.875000 1.210000 7.045000 1.380000 ;
    LAYER met1 ;
      RECT 2.495000 1.180000 2.785000 1.225000 ;
      RECT 2.495000 1.225000 7.105000 1.365000 ;
      RECT 2.495000 1.365000 2.785000 1.410000 ;
      RECT 6.815000 1.180000 7.105000 1.225000 ;
      RECT 6.815000 1.365000 7.105000 1.410000 ;
  END
END sky130_fd_sc_lp__dfbbp_1
