* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B1 a_43_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_43_65# B2 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 Y B2 a_43_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_43_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND A1 a_43_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_43_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_491_367# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_43_367# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR B1 a_43_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND A2 a_43_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_43_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_491_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 Y A2 a_491_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_43_65# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y B2 a_43_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR A1 a_491_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
