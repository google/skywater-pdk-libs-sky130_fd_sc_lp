* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
X0 a_251_47# a_44_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_455_367# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_251_367# a_44_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR a_44_367# a_251_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 Y A0 a_455_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_251_367# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_423_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_44_367# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND S a_423_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_455_367# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 Y A1 a_251_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y A0 a_251_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_251_47# A0 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_44_367# S VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y A1 a_423_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VGND a_44_367# a_251_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VPWR S a_455_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_423_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
