* NGSPICE file created from sky130_fd_sc_lp__or4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
M1000 a_415_391# a_196_535# a_332_391# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1001 X a_332_391# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=4.977e+11p ps=4.67e+06u
M1002 a_487_391# a_27_535# a_415_391# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1003 a_196_535# D_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1004 VGND a_27_535# a_332_391# VNB nshort w=420000u l=150000u
+  ad=6.573e+11p pd=6.8e+06u as=2.352e+11p ps=2.8e+06u
M1005 a_595_391# B a_487_391# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 VPWR A a_595_391# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_332_391# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C_N a_27_535# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1009 a_196_535# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1010 a_332_391# a_196_535# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C_N a_27_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 X a_332_391# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1013 a_332_391# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

