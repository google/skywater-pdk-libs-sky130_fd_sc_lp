* File: sky130_fd_sc_lp__or4b_m.pex.spice
* Created: Fri Aug 28 11:26:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4B_M%D_N 2 5 9 11 12 13 17 18
r34 17 19 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.412 $Y=1.655
+ $X2=0.412 $Y2=1.49
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.655 $X2=0.385 $Y2=1.655
r36 12 13 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=2.035
r37 12 18 0.365855 $w=3.13e-07 $l=1e-08 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=1.655
r38 9 11 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.53 $Y=2.73 $X2=0.53
+ $Y2=2.16
r39 5 19 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.53 $Y=0.835
+ $X2=0.53 $Y2=1.49
r40 2 11 49.2522 $w=3.85e-07 $l=1.92e-07 $layer=POLY_cond $X=0.412 $Y=1.968
+ $X2=0.412 $Y2=2.16
r41 1 17 3.9003 $w=3.85e-07 $l=2.7e-08 $layer=POLY_cond $X=0.412 $Y=1.682
+ $X2=0.412 $Y2=1.655
r42 1 2 41.3143 $w=3.85e-07 $l=2.86e-07 $layer=POLY_cond $X=0.412 $Y=1.682
+ $X2=0.412 $Y2=1.968
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%A_38_125# 1 2 9 10 11 14 17 18 21 25 27 28 29
+ 32 33 35 40
c69 29 0 1.47672e-19 $X=0.857 $Y=1.31
r70 35 40 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=0.735 $Y=2.34
+ $X2=0.735 $Y2=1.825
r71 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.98
+ $Y=1.32 $X2=0.98 $Y2=1.32
r72 30 40 9.87967 $w=4.13e-07 $l=2.07e-07 $layer=LI1_cond $X=0.857 $Y=1.618
+ $X2=0.857 $Y2=1.825
r73 30 32 8.27537 $w=4.13e-07 $l=2.98e-07 $layer=LI1_cond $X=0.857 $Y=1.618
+ $X2=0.857 $Y2=1.32
r74 29 32 0.277697 $w=4.13e-07 $l=1e-08 $layer=LI1_cond $X=0.857 $Y=1.31
+ $X2=0.857 $Y2=1.32
r75 27 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.65 $Y=2.425
+ $X2=0.735 $Y2=2.34
r76 27 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.65 $Y=2.425
+ $X2=0.4 $Y2=2.425
r77 23 28 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.305 $Y=2.51
+ $X2=0.4 $Y2=2.425
r78 23 25 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=0.305 $Y=2.51
+ $X2=0.305 $Y2=2.665
r79 19 29 35.3604 $w=1.68e-07 $l=5.42e-07 $layer=LI1_cond $X=0.315 $Y=1.225
+ $X2=0.857 $Y2=1.225
r80 19 21 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.315 $Y=1.14
+ $X2=0.315 $Y2=0.9
r81 18 33 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.98 $Y=1.675
+ $X2=0.98 $Y2=1.32
r82 17 33 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.155
+ $X2=0.98 $Y2=1.32
r83 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.615 $Y=1.825
+ $X2=1.615 $Y2=2.195
r84 11 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.145 $Y=1.75
+ $X2=0.98 $Y2=1.675
r85 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.54 $Y=1.75
+ $X2=1.615 $Y2=1.825
r86 10 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.54 $Y=1.75
+ $X2=1.145 $Y2=1.75
r87 9 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1 $Y=0.835 $X2=1
+ $Y2=1.155
r88 2 25 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=2.52 $X2=0.315 $Y2=2.665
r89 1 21 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.625 $X2=0.315 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%C 1 3 4 5 9 10 11 12 17
c44 17 0 2.40824e-19 $X=1.885 $Y=2.94
c45 1 0 1.47672e-19 $X=1.43 $Y=1.155
r46 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=2.94
+ $X2=1.885 $Y2=2.775
r47 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=2.94 $X2=1.885 $Y2=2.94
r48 12 18 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=2.16 $Y=2.857
+ $X2=1.885 $Y2=2.857
r49 11 18 7.05226 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=1.68 $Y=2.857
+ $X2=1.885 $Y2=2.857
r50 10 11 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.857
+ $X2=1.68 $Y2=2.857
r51 9 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.975 $Y=2.195
+ $X2=1.975 $Y2=2.775
r52 6 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.975 $Y=1.305
+ $X2=1.975 $Y2=2.195
r53 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.9 $Y=1.23
+ $X2=1.975 $Y2=1.305
r54 4 5 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.9 $Y=1.23 $X2=1.505
+ $Y2=1.23
r55 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.43 $Y=1.155
+ $X2=1.505 $Y2=1.23
r56 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.43 $Y=1.155 $X2=1.43
+ $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%B 3 5 7 8 12
r28 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.245 $Y=0.35
+ $X2=2.245 $Y2=0.515
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.245
+ $Y=0.35 $X2=2.245 $Y2=0.35
r30 8 13 12.1391 $w=3.73e-07 $l=3.95e-07 $layer=LI1_cond $X=2.64 $Y=0.452
+ $X2=2.245 $Y2=0.452
r31 7 13 2.6122 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.452
+ $X2=2.245 $Y2=0.452
r32 3 5 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=2.335 $Y=0.835
+ $X2=2.335 $Y2=2.195
r33 3 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.335 $Y=0.835
+ $X2=2.335 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%A 3 7 9 10 11 12 18
r39 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.66
+ $X2=2.785 $Y2=1.825
r40 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.66
+ $X2=2.785 $Y2=1.495
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=1.66 $X2=2.785 $Y2=1.66
r42 12 19 21.2312 $w=1.73e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=1.662
+ $X2=2.785 $Y2=1.662
r43 11 19 9.18961 $w=1.73e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.662
+ $X2=2.785 $Y2=1.662
r44 10 11 30.4208 $w=1.73e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.662
+ $X2=2.64 $Y2=1.662
r45 9 10 30.4208 $w=1.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.662
+ $X2=2.16 $Y2=1.662
r46 7 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.765 $Y=0.835
+ $X2=2.765 $Y2=1.495
r47 3 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.695 $Y=2.195
+ $X2=2.695 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%A_215_125# 1 2 3 10 15 18 21 23 25 26 28 32
+ 35 39 41 46 49
c107 46 0 1.62868e-19 $X=2.65 $Y=2.94
c108 35 0 7.79559e-20 $X=2.57 $Y=2.855
r109 47 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.65 $Y=2.94 $X2=2.65
+ $Y2=2.85
r110 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=2.94 $X2=2.65 $Y2=2.94
r111 37 39 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.215 $Y=0.855
+ $X2=1.33 $Y2=0.855
r112 35 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=2.855
+ $X2=2.57 $Y2=2.94
r113 34 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.57 $Y=2.335
+ $X2=2.57 $Y2=2.855
r114 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.55 $Y=1.225
+ $X2=2.55 $Y2=0.92
r115 29 43 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=2.17
+ $X2=1.33 $Y2=2.17
r116 28 34 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.485 $Y=2.17
+ $X2=2.57 $Y2=2.335
r117 28 29 37.3671 $w=3.28e-07 $l=1.07e-06 $layer=LI1_cond $X=2.485 $Y=2.17
+ $X2=1.415 $Y2=2.17
r118 27 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=1.31
+ $X2=1.33 $Y2=1.31
r119 26 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.385 $Y=1.31
+ $X2=2.55 $Y2=1.225
r120 26 27 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=2.385 $Y=1.31
+ $X2=1.415 $Y2=1.31
r121 25 43 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=2.005
+ $X2=1.33 $Y2=2.17
r122 24 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=1.395
+ $X2=1.33 $Y2=1.31
r123 24 25 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.33 $Y=1.395
+ $X2=1.33 $Y2=2.005
r124 23 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=1.225
+ $X2=1.33 $Y2=1.31
r125 22 39 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.33 $Y=0.96
+ $X2=1.33 $Y2=0.855
r126 22 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.33 $Y=0.96
+ $X2=1.33 $Y2=1.225
r127 20 21 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.245 $Y=1.725
+ $X2=3.245 $Y2=1.875
r128 18 20 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.255 $Y=0.835
+ $X2=3.255 $Y2=1.725
r129 15 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.235 $Y=2.195
+ $X2=3.235 $Y2=1.875
r130 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.235 $Y=2.775
+ $X2=3.235 $Y2=2.195
r131 11 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=2.85
+ $X2=2.65 $Y2=2.85
r132 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.16 $Y=2.85
+ $X2=3.235 $Y2=2.775
r133 10 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=3.16 $Y=2.85
+ $X2=2.815 $Y2=2.85
r134 3 43 600 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.985 $X2=1.4 $Y2=2.17
r135 2 32 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.625 $X2=2.55 $Y2=0.92
r136 1 37 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.625 $X2=1.215 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%VPWR 1 2 9 12 16 19 20 21 23 36 37 40
r45 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 31 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 30 33 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 28 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.745 $Y2=3.33
r53 28 30 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 26 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 23 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.745 $Y2=3.33
r57 23 25 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 21 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 21 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 19 33 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.08 $Y2=3.33
r62 18 36 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.08 $Y2=3.33
r64 14 16 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=3 $Y=2.26 $X2=3.08
+ $Y2=2.26
r65 12 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=3.33
r66 11 16 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.08 $Y=2.365
+ $X2=3.08 $Y2=2.26
r67 11 12 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=3.08 $Y=2.365
+ $X2=3.08 $Y2=3.245
r68 7 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=3.33
r69 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=2.795
r70 2 14 600 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.985 $X2=3 $Y2=2.26
r71 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=2.52 $X2=0.745 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%X 1 2 7 8 9 10 11 12 13 46
r16 34 46 2.2032 $w=3.38e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=2.1
+ $X2=3.515 $Y2=2.035
r17 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.515 $Y=2.405
+ $X2=3.515 $Y2=2.775
r18 12 37 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=3.515 $Y=2.405
+ $X2=3.515 $Y2=2.13
r19 11 46 0.338954 $w=3.38e-07 $l=1e-08 $layer=LI1_cond $X=3.515 $Y=2.025
+ $X2=3.515 $Y2=2.035
r20 11 44 3.40832 $w=3.38e-07 $l=9.5e-08 $layer=LI1_cond $X=3.515 $Y=2.025
+ $X2=3.515 $Y2=1.93
r21 11 37 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=3.515 $Y=2.11
+ $X2=3.515 $Y2=2.13
r22 11 34 0.338954 $w=3.38e-07 $l=1e-08 $layer=LI1_cond $X=3.515 $Y=2.11
+ $X2=3.515 $Y2=2.1
r23 10 44 10.1799 $w=2.98e-07 $l=2.65e-07 $layer=LI1_cond $X=3.535 $Y=1.665
+ $X2=3.535 $Y2=1.93
r24 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.535 $Y=1.295
+ $X2=3.535 $Y2=1.665
r25 8 9 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.535 $Y=0.925
+ $X2=3.535 $Y2=1.295
r26 8 27 5.95429 $w=2.98e-07 $l=1.55e-07 $layer=LI1_cond $X=3.535 $Y=0.925
+ $X2=3.535 $Y2=0.77
r27 7 27 8.25918 $w=2.98e-07 $l=2.15e-07 $layer=LI1_cond $X=3.535 $Y=0.555
+ $X2=3.535 $Y2=0.77
r28 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.985 $X2=3.45 $Y2=2.13
r29 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.625 $X2=3.47 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_M%VGND 1 2 3 14 18 22 25 26 27 29 39 40 43 46
r50 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r53 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r54 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r55 34 46 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.7
+ $Y2=0
r56 34 36 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=2.64
+ $Y2=0
r57 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r58 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r59 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r60 30 43 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=0.765
+ $Y2=0
r61 30 32 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=1.2
+ $Y2=0
r62 29 46 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.595 $Y=0 $X2=1.7
+ $Y2=0
r63 29 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.595 $Y=0 $X2=1.2
+ $Y2=0
r64 27 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r65 27 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r66 25 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r67 25 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.01
+ $Y2=0
r68 24 39 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.6
+ $Y2=0
r69 24 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.01
+ $Y2=0
r70 20 26 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=0.085
+ $X2=3.01 $Y2=0
r71 20 22 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=3.01 $Y=0.085
+ $X2=3.01 $Y2=0.77
r72 16 46 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r73 16 18 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.77
r74 12 43 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0
r75 12 14 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0.77
r76 3 22 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=2.84
+ $Y=0.625 $X2=3.01 $Y2=0.77
r77 2 18 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.625 $X2=1.7 $Y2=0.77
r78 1 14 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.625 $X2=0.765 $Y2=0.77
.ends

