# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o21bai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.425000 3.335000 1.930000 ;
        RECT 3.005000 1.930000 5.435000 2.100000 ;
        RECT 5.265000 1.375000 6.615000 1.760000 ;
        RECT 5.265000 1.760000 5.435000 1.930000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.425000 4.910000 1.750000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.415000 0.550000 1.760000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.881600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 1.755000 2.725000 1.925000 ;
        RECT 1.510000 1.925000 1.740000 3.075000 ;
        RECT 1.550000 0.775000 2.725000 1.185000 ;
        RECT 2.335000 1.185000 2.725000 1.755000 ;
        RECT 2.410000 1.925000 2.725000 2.280000 ;
        RECT 2.410000 2.280000 4.790000 2.530000 ;
        RECT 2.410000 2.530000 2.600000 3.075000 ;
        RECT 3.240000 2.530000 4.790000 2.610000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.255000 0.355000 1.075000 ;
      RECT 0.095000  1.075000 0.930000 1.245000 ;
      RECT 0.150000  1.930000 0.930000 2.100000 ;
      RECT 0.150000  2.100000 0.445000 3.075000 ;
      RECT 0.525000  0.085000 0.855000 0.905000 ;
      RECT 0.615000  2.270000 1.340000 3.245000 ;
      RECT 0.760000  1.245000 0.930000 1.325000 ;
      RECT 0.760000  1.325000 1.380000 1.355000 ;
      RECT 0.760000  1.355000 2.165000 1.585000 ;
      RECT 0.760000  1.585000 1.340000 1.655000 ;
      RECT 0.760000  1.655000 0.930000 1.930000 ;
      RECT 1.050000  0.255000 3.085000 0.595000 ;
      RECT 1.050000  0.595000 1.380000 0.945000 ;
      RECT 1.100000  1.825000 1.340000 2.270000 ;
      RECT 1.910000  2.105000 2.240000 3.245000 ;
      RECT 2.770000  2.700000 3.070000 3.245000 ;
      RECT 2.895000  0.595000 3.085000 1.055000 ;
      RECT 2.895000  1.055000 6.595000 1.205000 ;
      RECT 2.895000  1.205000 4.795000 1.225000 ;
      RECT 3.240000  2.790000 5.220000 3.075000 ;
      RECT 3.255000  0.085000 3.585000 0.885000 ;
      RECT 3.755000  0.255000 3.945000 1.055000 ;
      RECT 4.115000  0.085000 4.445000 0.885000 ;
      RECT 4.615000  0.255000 4.805000 1.015000 ;
      RECT 4.615000  1.015000 5.665000 1.035000 ;
      RECT 4.615000  1.035000 6.595000 1.055000 ;
      RECT 4.960000  2.270000 6.080000 2.460000 ;
      RECT 4.960000  2.460000 5.220000 2.790000 ;
      RECT 4.975000  0.085000 5.305000 0.845000 ;
      RECT 5.390000  2.630000 5.720000 3.245000 ;
      RECT 5.475000  0.255000 5.665000 1.015000 ;
      RECT 5.835000  0.085000 6.165000 0.865000 ;
      RECT 5.880000  1.930000 6.080000 2.270000 ;
      RECT 5.890000  2.460000 6.080000 3.075000 ;
      RECT 6.250000  1.930000 6.580000 3.245000 ;
      RECT 6.335000  0.255000 6.595000 1.035000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__o21bai_4
