* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4b_2 A_N B C D VGND VNB VPB VPWR X
X0 a_222_375# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR C a_222_375# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_306_125# B a_378_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_222_375# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_53_375# a_222_375# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_450_125# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_222_375# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_222_375# a_53_375# a_306_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_222_375# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_53_375# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_378_125# C a_450_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_222_375# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 X a_222_375# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND A_N a_53_375# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
