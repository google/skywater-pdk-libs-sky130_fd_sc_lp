* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__bufinv_8 A VGND VNB VPB VPWR Y
X0 Y a_82_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 Y a_82_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_82_23# a_876_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND a_82_23# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND A a_876_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Y a_82_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y a_82_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND a_82_23# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_82_23# a_876_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND a_876_23# a_82_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 Y a_82_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR a_82_23# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR a_82_23# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_82_23# a_876_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND a_82_23# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR a_82_23# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_82_23# a_876_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VGND a_82_23# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 Y a_82_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VPWR A a_876_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR a_82_23# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 Y a_82_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 Y a_82_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VPWR a_876_23# a_82_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
