* File: sky130_fd_sc_lp__nand4_2.pex.spice
* Created: Wed Sep  2 10:05:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4_2%D 3 5 7 10 12 14 15 16 25
c41 25 0 7.78649e-20 $X=1.115 $Y=1.535
r42 27 32 4.1044 $w=1.8e-07 $l=1.63e-07 $layer=LI1_cond $X=0.715 $Y=1.67
+ $X2=0.715 $Y2=1.507
r43 24 25 37.861 $w=3.31e-07 $l=2.6e-07 $layer=POLY_cond $X=0.855 $Y=1.535
+ $X2=1.115 $Y2=1.535
r44 22 24 19.6586 $w=3.31e-07 $l=1.35e-07 $layer=POLY_cond $X=0.72 $Y=1.535
+ $X2=0.855 $Y2=1.535
r45 20 22 5.09668 $w=3.31e-07 $l=3.5e-08 $layer=POLY_cond $X=0.685 $Y=1.535
+ $X2=0.72 $Y2=1.535
r46 15 32 0.190625 $w=3.2e-07 $l=5e-09 $layer=LI1_cond $X=0.72 $Y=1.507
+ $X2=0.715 $Y2=1.507
r47 15 16 20.0253 $w=1.78e-07 $l=3.25e-07 $layer=LI1_cond $X=0.715 $Y=1.71
+ $X2=0.715 $Y2=2.035
r48 15 27 2.46465 $w=1.78e-07 $l=4e-08 $layer=LI1_cond $X=0.715 $Y=1.71
+ $X2=0.715 $Y2=1.67
r49 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.51 $X2=0.72 $Y2=1.51
r50 12 25 24.7553 $w=3.31e-07 $l=2.61534e-07 $layer=POLY_cond $X=1.285 $Y=1.725
+ $X2=1.115 $Y2=1.535
r51 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.285 $Y=1.725
+ $X2=1.285 $Y2=2.465
r52 8 25 21.295 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.115 $Y=1.345
+ $X2=1.115 $Y2=1.535
r53 8 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.115 $Y=1.345
+ $X2=1.115 $Y2=0.655
r54 5 24 21.295 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.855 $Y=1.725
+ $X2=0.855 $Y2=1.535
r55 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.855 $Y=1.725
+ $X2=0.855 $Y2=2.465
r56 1 20 21.295 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.685 $Y=1.345
+ $X2=0.685 $Y2=1.535
r57 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.685 $Y=1.345
+ $X2=0.685 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%C 1 3 6 8 10 13 15 16 22
c52 16 0 2.28515e-19 $X=2.16 $Y=1.295
r53 22 24 4.36199 $w=2.21e-07 $l=2e-08 $layer=POLY_cond $X=2.145 $Y=1.335
+ $X2=2.165 $Y2=1.335
r54 21 22 30.5339 $w=2.21e-07 $l=1.4e-07 $layer=POLY_cond $X=2.005 $Y=1.335
+ $X2=2.145 $Y2=1.335
r55 16 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.35 $X2=2.165 $Y2=1.35
r56 15 16 20.4879 $w=2.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.3 $X2=2.16
+ $Y2=1.3
r57 11 22 11.8763 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.145 $Y=1.515
+ $X2=2.145 $Y2=1.335
r58 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.145 $Y=1.515
+ $X2=2.145 $Y2=2.465
r59 8 21 11.8763 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.005 $Y=1.185
+ $X2=2.005 $Y2=1.335
r60 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.005 $Y=1.185
+ $X2=2.005 $Y2=0.655
r61 4 21 63.2489 $w=2.21e-07 $l=2.9e-07 $layer=POLY_cond $X=1.715 $Y=1.335
+ $X2=2.005 $Y2=1.335
r62 4 19 30.5339 $w=2.21e-07 $l=1.4e-07 $layer=POLY_cond $X=1.715 $Y=1.335
+ $X2=1.575 $Y2=1.335
r63 4 6 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=1.715 $Y=1.335
+ $X2=1.715 $Y2=2.465
r64 1 19 11.8763 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.575 $Y=1.185
+ $X2=1.575 $Y2=1.335
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.575 $Y=1.185
+ $X2=1.575 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%B 3 5 6 9 13 17 19 24 25
c57 25 0 3.75208e-19 $X=3.17 $Y=1.51
c58 9 0 1.3307e-19 $X=2.975 $Y=0.755
c59 6 0 9.54453e-20 $X=2.73 $Y=1.42
c60 5 0 2.49271e-20 $X=2.9 $Y=1.42
r61 24 26 38.138 $w=2.97e-07 $l=2.35e-07 $layer=POLY_cond $X=3.17 $Y=1.51
+ $X2=3.405 $Y2=1.51
r62 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.51 $X2=3.17 $Y2=1.51
r63 22 24 13.7946 $w=2.97e-07 $l=8.5e-08 $layer=POLY_cond $X=3.085 $Y=1.51
+ $X2=3.17 $Y2=1.51
r64 19 25 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.17 $Y=1.665
+ $X2=3.17 $Y2=1.51
r65 15 26 18.7323 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.405 $Y=1.345
+ $X2=3.405 $Y2=1.51
r66 15 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.405 $Y=1.345
+ $X2=3.405 $Y2=0.755
r67 11 22 18.7323 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.675
+ $X2=3.085 $Y2=1.51
r68 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.085 $Y=1.675
+ $X2=3.085 $Y2=2.465
r69 7 22 17.8519 $w=2.97e-07 $l=2.13014e-07 $layer=POLY_cond $X=2.975 $Y=1.345
+ $X2=3.085 $Y2=1.51
r70 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.975 $Y=1.345
+ $X2=2.975 $Y2=0.755
r71 5 7 23.9601 $w=2.97e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.9 $Y=1.42
+ $X2=2.975 $Y2=1.345
r72 5 6 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.9 $Y=1.42 $X2=2.73
+ $Y2=1.42
r73 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.655 $Y=1.495
+ $X2=2.73 $Y2=1.42
r74 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.655 $Y=1.495
+ $X2=2.655 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%A 3 7 11 15 17 18 19 29
c44 29 0 1.76493e-19 $X=4.265 $Y=1.51
c45 3 0 1.98715e-19 $X=3.765 $Y=2.465
r46 27 29 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.195 $Y=1.51
+ $X2=4.265 $Y2=1.51
r47 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.195
+ $Y=1.51 $X2=4.195 $Y2=1.51
r48 25 27 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.835 $Y=1.51
+ $X2=4.195 $Y2=1.51
r49 23 25 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.765 $Y=1.51
+ $X2=3.835 $Y2=1.51
r50 19 28 12.9428 $w=3.23e-07 $l=3.65e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.195 $Y2=1.587
r51 18 28 4.07788 $w=3.23e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.195 $Y2=1.587
r52 17 18 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.587
+ $X2=4.08 $Y2=1.587
r53 13 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.345
+ $X2=4.265 $Y2=1.51
r54 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.265 $Y=1.345
+ $X2=4.265 $Y2=0.755
r55 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=1.675
+ $X2=4.195 $Y2=1.51
r56 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.195 $Y=1.675
+ $X2=4.195 $Y2=2.465
r57 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.345
+ $X2=3.835 $Y2=1.51
r58 5 7 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.835 $Y=1.345
+ $X2=3.835 $Y2=0.755
r59 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.675
+ $X2=3.765 $Y2=1.51
r60 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.765 $Y=1.675
+ $X2=3.765 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%VPWR 1 2 3 4 5 18 21 24 30 34 36 38 43 46 47
+ 49 50 52 53 54 66 75
r74 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 69 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 66 74 4.53846 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.522 $Y2=3.33
r79 66 68 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.08 $Y2=3.33
r80 65 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r81 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r82 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r83 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 59 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r86 56 71 7.66976 $w=1.7e-07 $l=4.03e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.402 $Y2=3.33
r87 56 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r88 54 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r89 54 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r90 52 64 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.12 $Y2=3.33
r91 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.425 $Y2=3.33
r92 51 68 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=3.425 $Y2=3.33
r94 49 61 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.24 $Y=3.33 $X2=2.16
+ $Y2=3.33
r95 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=3.33
+ $X2=2.405 $Y2=3.33
r96 48 64 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=3.12 $Y2=3.33
r97 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=2.405 $Y2=3.33
r98 46 58 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.5 $Y2=3.33
r100 45 61 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=1.5 $Y2=3.33
r102 43 44 6.22405 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.47 $Y=2.46
+ $X2=0.47 $Y2=2.295
r103 38 41 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=4.41 $Y=2.005
+ $X2=4.41 $Y2=2.95
r104 36 74 3.22771 $w=3.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.41 $Y=3.245
+ $X2=4.522 $Y2=3.33
r105 36 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.41 $Y=3.245
+ $X2=4.41 $Y2=2.95
r106 32 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=3.33
r107 32 34 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=2.38
r108 28 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=3.245
+ $X2=2.405 $Y2=3.33
r109 28 30 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=2.405 $Y=3.245
+ $X2=2.405 $Y2=2.38
r110 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.5 $Y=2.18 $X2=1.5
+ $Y2=2.95
r111 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=3.245 $X2=1.5
+ $Y2=3.33
r112 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.5 $Y=3.245
+ $X2=1.5 $Y2=2.95
r113 21 71 2.91184 $w=6.7e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.47 $Y=3.245
+ $X2=0.402 $Y2=3.33
r114 20 43 3.03483 $w=6.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.47 $Y=2.63
+ $X2=0.47 $Y2=2.46
r115 20 21 10.9789 $w=6.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.47 $Y=2.63
+ $X2=0.47 $Y2=3.245
r116 18 44 11.3444 $w=3.18e-07 $l=3.15e-07 $layer=LI1_cond $X=0.295 $Y=1.98
+ $X2=0.295 $Y2=2.295
r117 5 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.835 $X2=4.41 $Y2=2.95
r118 5 38 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.835 $X2=4.41 $Y2=2.005
r119 4 34 300 $w=1.7e-07 $l=6.64417e-07 $layer=licon1_PDIFF $count=2 $X=3.16
+ $Y=1.835 $X2=3.425 $Y2=2.38
r120 3 30 300 $w=1.7e-07 $l=6.30754e-07 $layer=licon1_PDIFF $count=2 $X=2.22
+ $Y=1.835 $X2=2.405 $Y2=2.38
r121 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.95
r122 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.18
r123 1 43 150 $w=1.7e-07 $l=8.25379e-07 $layer=licon1_PDIFF $count=4 $X=0.175
+ $Y=1.835 $X2=0.64 $Y2=2.46
r124 1 18 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.835 $X2=0.3 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%Y 1 2 3 4 5 18 22 23 26 30 32 33 34 35 36 38
+ 42 47
c92 32 0 7.45928e-20 $X=3.885 $Y=1.16
r93 57 59 6.04049 $w=4.1e-07 $l=2.70708e-07 $layer=LI1_cond $X=2.667 $Y=1.847
+ $X2=2.87 $Y2=2.005
r94 52 54 0.14878 $w=4.1e-07 $l=5e-09 $layer=LI1_cond $X=1.925 $Y=1.847 $X2=1.93
+ $Y2=1.847
r95 50 57 1.93746 $w=3.35e-07 $l=2.42e-07 $layer=LI1_cond $X=2.667 $Y=1.605
+ $X2=2.667 $Y2=1.847
r96 47 57 0.803415 $w=4.1e-07 $l=2.7e-08 $layer=LI1_cond $X=2.64 $Y=1.847
+ $X2=2.667 $Y2=1.847
r97 47 54 21.1268 $w=4.1e-07 $l=7.1e-07 $layer=LI1_cond $X=2.64 $Y=1.847
+ $X2=1.93 $Y2=1.847
r98 47 50 0.447217 $w=3.33e-07 $l=1.3e-08 $layer=LI1_cond $X=2.667 $Y=1.592
+ $X2=2.667 $Y2=1.605
r99 44 47 11.9372 $w=3.33e-07 $l=3.47e-07 $layer=LI1_cond $X=2.667 $Y=1.245
+ $X2=2.667 $Y2=1.592
r100 40 42 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.05 $Y=1.075
+ $X2=4.05 $Y2=0.68
r101 36 46 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.945 $Y=2.09
+ $X2=3.945 $Y2=2.005
r102 36 38 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=3.945 $Y=2.09
+ $X2=3.945 $Y2=2.91
r103 35 59 9.20018 $w=4.1e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=2.005
+ $X2=2.87 $Y2=2.005
r104 34 46 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.815 $Y=2.005
+ $X2=3.945 $Y2=2.005
r105 34 35 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.815 $Y=2.005
+ $X2=3.035 $Y2=2.005
r106 33 44 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=2.835 $Y=1.16
+ $X2=2.667 $Y2=1.245
r107 32 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.885 $Y=1.16
+ $X2=4.05 $Y2=1.075
r108 32 33 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.885 $Y=1.16
+ $X2=2.835 $Y2=1.16
r109 28 59 2.68093 $w=2.95e-07 $l=9.31128e-08 $layer=LI1_cond $X=2.887 $Y=2.09
+ $X2=2.87 $Y2=2.005
r110 28 30 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.887 $Y=2.09
+ $X2=2.887 $Y2=2.46
r111 24 52 5.58152 $w=1.8e-07 $l=2.43e-07 $layer=LI1_cond $X=1.925 $Y=2.09
+ $X2=1.925 $Y2=1.847
r112 24 26 21.5657 $w=1.78e-07 $l=3.5e-07 $layer=LI1_cond $X=1.925 $Y=2.09
+ $X2=1.925 $Y2=2.44
r113 22 52 6.96848 $w=4.1e-07 $l=9.34345e-08 $layer=LI1_cond $X=1.835 $Y=1.84
+ $X2=1.925 $Y2=1.847
r114 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.835 $Y=1.84
+ $X2=1.165 $Y2=1.84
r115 18 20 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.07 $Y=1.98
+ $X2=1.07 $Y2=2.91
r116 16 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.07 $Y=1.925
+ $X2=1.165 $Y2=1.84
r117 16 18 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.07 $Y=1.925
+ $X2=1.07 $Y2=1.98
r118 5 46 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.84
+ $Y=1.835 $X2=3.98 $Y2=2.085
r119 5 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.84
+ $Y=1.835 $X2=3.98 $Y2=2.91
r120 4 59 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.835 $X2=2.87 $Y2=2.005
r121 4 30 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=2.73
+ $Y=1.835 $X2=2.87 $Y2=2.46
r122 3 54 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=1.98
r123 3 26 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=2.44
r124 2 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=1.835 $X2=1.07 $Y2=2.91
r125 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=1.835 $X2=1.07 $Y2=1.98
r126 1 42 91 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=2 $X=3.91
+ $Y=0.335 $X2=4.05 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%A_69_47# 1 2 3 12 14 15 16 19 22
c35 15 0 7.78649e-20 $X=0.565 $Y=1.07
r36 20 25 2.80098 $w=2.9e-07 $l=9e-08 $layer=LI1_cond $X=1.415 $Y=0.4 $X2=1.325
+ $Y2=0.4
r37 20 22 31.9902 $w=2.88e-07 $l=8.05e-07 $layer=LI1_cond $X=1.415 $Y=0.4
+ $X2=2.22 $Y2=0.4
r38 17 19 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.325 $Y=0.985
+ $X2=1.325 $Y2=0.93
r39 16 25 4.5127 $w=1.8e-07 $l=1.45e-07 $layer=LI1_cond $X=1.325 $Y=0.545
+ $X2=1.325 $Y2=0.4
r40 16 19 23.7222 $w=1.78e-07 $l=3.85e-07 $layer=LI1_cond $X=1.325 $Y=0.545
+ $X2=1.325 $Y2=0.93
r41 14 17 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.235 $Y=1.07
+ $X2=1.325 $Y2=0.985
r42 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.235 $Y=1.07
+ $X2=0.565 $Y2=1.07
r43 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.435 $Y=0.985
+ $X2=0.565 $Y2=1.07
r44 10 12 25.0435 $w=2.58e-07 $l=5.65e-07 $layer=LI1_cond $X=0.435 $Y=0.985
+ $X2=0.435 $Y2=0.42
r45 3 22 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.235 $X2=2.22 $Y2=0.41
r46 2 25 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.19
+ $Y=0.235 $X2=1.33 $Y2=0.42
r47 2 19 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.19
+ $Y=0.235 $X2=1.33 $Y2=0.93
r48 1 12 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.345
+ $Y=0.235 $X2=0.47 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%VGND 1 6 9 10 11 21 22
r44 21 22 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r45 18 21 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r46 18 19 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r48 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 11 22 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=4.56
+ $Y2=0
r50 11 19 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r51 9 14 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.72
+ $Y2=0
r52 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.9
+ $Y2=0
r53 8 18 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.2
+ $Y2=0
r54 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.9
+ $Y2=0
r55 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0
r56 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0.36
r57 1 6 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.76
+ $Y=0.235 $X2=0.9 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%A_330_47# 1 2 9 14
c25 9 0 2.49271e-20 $X=3.19 $Y=0.81
r26 12 14 7.98846 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=0.855
+ $X2=1.955 $Y2=0.855
r27 9 14 72.0909 $w=1.88e-07 $l=1.235e-06 $layer=LI1_cond $X=3.19 $Y=0.81
+ $X2=1.955 $Y2=0.81
r28 2 9 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=3.05
+ $Y=0.335 $X2=3.19 $Y2=0.81
r29 1 12 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.235 $X2=1.79 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_2%A_523_67# 1 2 3 10 16 18 22 24
c28 1 0 7.45928e-20 $X=2.615 $Y=0.335
r29 20 22 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=4.515 $Y=0.425
+ $X2=4.515 $Y2=0.48
r30 19 24 4.39427 $w=2.3e-07 $l=1.21347e-07 $layer=LI1_cond $X=3.715 $Y=0.34
+ $X2=3.62 $Y2=0.4
r31 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.385 $Y=0.34
+ $X2=4.515 $Y2=0.425
r32 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.385 $Y=0.34
+ $X2=3.715 $Y2=0.34
r33 14 24 2.03875 $w=1.9e-07 $l=1.45e-07 $layer=LI1_cond $X=3.62 $Y=0.545
+ $X2=3.62 $Y2=0.4
r34 14 16 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.62 $Y=0.545
+ $X2=3.62 $Y2=0.74
r35 10 24 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.525 $Y=0.4 $X2=3.62
+ $Y2=0.4
r36 10 12 30.4007 $w=2.88e-07 $l=7.65e-07 $layer=LI1_cond $X=3.525 $Y=0.4
+ $X2=2.76 $Y2=0.4
r37 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.34
+ $Y=0.335 $X2=4.48 $Y2=0.48
r38 2 16 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=3.48
+ $Y=0.335 $X2=3.62 $Y2=0.74
r39 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.335 $X2=2.76 $Y2=0.46
.ends

