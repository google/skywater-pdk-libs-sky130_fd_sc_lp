* File: sky130_fd_sc_lp__o22a_1.spice
* Created: Wed Sep  2 10:19:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22a_1.pex.spice"
.subckt sky130_fd_sc_lp__o22a_1  VNB VPB B1 B2 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_80_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_80_21#_M1000_d N_B1_M1000_g N_A_265_47#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2226 PD=1.14 PS=2.21 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1001 N_A_265_47#_M1001_d N_B2_M1001_g N_A_80_21#_M1000_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1617 AS=0.126 PD=1.225 PS=1.14 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_265_47#_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.1617 PD=1.26 PS=1.225 NRD=0 NRS=15 M=1 R=5.6 SA=75001.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1002 N_A_265_47#_M1002_d N_A1_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1764 PD=2.21 PS=1.26 NRD=0 NRS=19.992 M=1 R=5.6 SA=75001.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_A_80_21#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.33075 AS=0.3339 PD=1.785 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1008 A_348_367# N_B1_M1008_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.33075 PD=1.5 PS=1.785 NRD=10.1455 NRS=38.2968 M=1 R=8.4
+ SA=75000.9 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1009 N_A_80_21#_M1009_d N_B2_M1009_g A_348_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.28035 AS=0.1512 PD=1.705 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75001.3
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1005 A_545_367# N_A2_M1005_g N_A_80_21#_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.28035 PD=1.68 PS=1.705 NRD=24.231 NRS=25.7873 M=1 R=8.4
+ SA=75001.9 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_545_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4032 AS=0.2646 PD=3.16 PS=1.68 NRD=8.5892 NRS=24.231 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o22a_1.pxi.spice"
*
.ends
*
*
