* File: sky130_fd_sc_lp__a2111o_1.spice
* Created: Fri Aug 28 09:45:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111o_1.pex.spice"
.subckt sky130_fd_sc_lp__a2111o_1  VNB VPB D1 C1 B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_105_239#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3024 AS=0.2226 PD=1.56 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1011 N_A_105_239#_M1011_d N_D1_M1011_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3024 PD=1.12 PS=1.56 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_C1_M1000_g N_A_105_239#_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1176 PD=1.23 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1003 N_A_105_239#_M1003_d N_B1_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2772 AS=0.1638 PD=1.5 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1005 A_673_49# N_A1_M1005_g N_A_105_239#_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2772 PD=1.05 PS=1.5 NRD=7.14 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g A_673_49# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75003.2 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_105_239#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 A_325_367# N_D1_M1009_g N_A_105_239#_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3339 PD=1.5 PS=3.05 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1001 A_403_367# N_C1_M1001_g A_325_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1512 PD=1.65 PS=1.5 NRD=21.8867 NRS=10.1455 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1004 N_A_511_367#_M1004_d N_B1_M1004_g A_403_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.2457 PD=1.88 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75001.1
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_511_367#_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1002 N_A_511_367#_M1002_d N_A2_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a2111o_1.pxi.spice"
*
.ends
*
*
