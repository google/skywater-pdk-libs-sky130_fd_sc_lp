* File: sky130_fd_sc_lp__mux2i_lp2.pex.spice
* Created: Fri Aug 28 10:45:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2I_LP2%S 3 5 6 9 11 13 14 16 18 20 23 26 29 31 33
+ 34 35 40 42
c112 40 0 3.31133e-20 $X=3.035 $Y=0.93
c113 14 0 9.7113e-20 $X=3.175 $Y=1.28
c114 9 0 1.57e-19 $X=1.205 $Y=0.445
c115 5 0 7.69208e-20 $X=1.13 $Y=1.15
r116 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.035
+ $Y=0.93 $X2=3.035 $Y2=0.93
r117 35 40 11.9793 $w=3.78e-07 $l=3.95e-07 $layer=LI1_cond $X=2.64 $Y=0.905
+ $X2=3.035 $Y2=0.905
r118 35 42 7.05482 $w=3.78e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=0.905
+ $X2=2.525 $Y2=0.905
r119 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.24 $X2=0.605 $Y2=1.24
r120 31 42 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=1.38 $Y=0.8
+ $X2=2.525 $Y2=0.8
r121 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.295 $Y=0.885
+ $X2=1.38 $Y2=0.8
r122 28 29 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.295 $Y=0.885
+ $X2=1.295 $Y2=1.075
r123 27 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.605 $Y2=1.16
r124 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.16
+ $X2=1.295 $Y2=1.075
r125 26 27 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.21 $Y=1.16
+ $X2=0.77 $Y2=1.16
r126 22 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.605 $Y=1.58
+ $X2=0.605 $Y2=1.24
r127 22 23 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.58
+ $X2=0.605 $Y2=1.745
r128 21 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.605 $Y=1.225
+ $X2=0.605 $Y2=1.24
r129 18 39 45.8637 $w=1.74e-07 $l=2.62857e-07 $layer=POLY_cond $X=3.33 $Y=0.765
+ $X2=3.137 $Y2=0.93
r130 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.33 $Y=0.765
+ $X2=3.33 $Y2=0.445
r131 14 39 52.2904 $w=3.49e-07 $l=3.68511e-07 $layer=POLY_cond $X=3.175 $Y=1.28
+ $X2=3.137 $Y2=0.93
r132 14 16 326.716 $w=2.5e-07 $l=1.315e-06 $layer=POLY_cond $X=3.175 $Y=1.28
+ $X2=3.175 $Y2=2.595
r133 11 39 45.8637 $w=1.74e-07 $l=2.35465e-07 $layer=POLY_cond $X=2.97 $Y=0.765
+ $X2=3.137 $Y2=0.93
r134 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.97 $Y=0.765
+ $X2=2.97 $Y2=0.445
r135 7 9 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.205 $Y=1.075
+ $X2=1.205 $Y2=0.445
r136 6 21 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.77 $Y=1.15
+ $X2=0.605 $Y2=1.225
r137 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.13 $Y=1.15
+ $X2=1.205 $Y2=1.075
r138 5 6 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.13 $Y=1.15 $X2=0.77
+ $Y2=1.15
r139 3 23 211.186 $w=2.5e-07 $l=8.5e-07 $layer=POLY_cond $X=0.615 $Y=2.595
+ $X2=0.615 $Y2=1.745
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP2%A0 3 7 9 11 12 17 19 22
c64 12 0 1.06687e-19 $X=2.075 $Y=1.23
c65 11 0 7.38896e-20 $X=2.075 $Y=1.23
c66 9 0 1.57e-19 $X=1.73 $Y=1.23
r67 22 25 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.63
+ $X2=1.145 $Y2=1.795
r68 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.145
+ $Y=1.63 $X2=1.145 $Y2=1.63
r69 17 19 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.56 $Y=1.63
+ $X2=1.145 $Y2=1.63
r70 12 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.23
+ $X2=2.075 $Y2=1.065
r71 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.075
+ $Y=1.23 $X2=2.075 $Y2=1.23
r72 9 17 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.645 $Y=1.23 $X2=1.645
+ $Y2=1.63
r73 9 11 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.73 $Y=1.23
+ $X2=2.075 $Y2=1.23
r74 7 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.035 $Y=0.445
+ $X2=2.035 $Y2=1.065
r75 3 25 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=1.105 $Y=2.595
+ $X2=1.105 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP2%A1 3 7 9 12 15
c44 12 0 6.92517e-20 $X=1.925 $Y=1.77
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.075
+ $Y=1.77 $X2=2.075 $Y2=1.77
r46 12 14 27.8077 $w=2.6e-07 $l=1.5e-07 $layer=POLY_cond $X=1.925 $Y=1.77
+ $X2=2.075 $Y2=1.77
r47 9 15 8.36705 $w=3.63e-07 $l=2.65e-07 $layer=LI1_cond $X=2.092 $Y=2.035
+ $X2=2.092 $Y2=1.77
r48 5 12 3.77112 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.935
+ $X2=1.925 $Y2=1.77
r49 5 7 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.925 $Y=1.935
+ $X2=1.925 $Y2=2.595
r50 1 12 61.1769 $w=2.6e-07 $l=4.04166e-07 $layer=POLY_cond $X=1.595 $Y=1.605
+ $X2=1.925 $Y2=1.77
r51 1 3 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=1.595 $Y=1.605
+ $X2=1.595 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP2%A_490_21# 1 2 9 14 16 17 18 21 25 29 31 33
c64 21 0 7.38896e-20 $X=2.645 $Y=1.5
c65 18 0 1.42825e-19 $X=3.275 $Y=1.5
r66 27 31 4.56101 $w=3.82e-07 $l=1.89658e-07 $layer=LI1_cond $X=3.545 $Y=1.335
+ $X2=3.492 $Y2=1.5
r67 27 29 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=3.545 $Y=1.335
+ $X2=3.545 $Y2=0.47
r68 23 31 4.56101 $w=3.82e-07 $l=1.65e-07 $layer=LI1_cond $X=3.492 $Y=1.665
+ $X2=3.492 $Y2=1.5
r69 23 25 15.2334 $w=4.33e-07 $l=5.75e-07 $layer=LI1_cond $X=3.492 $Y=1.665
+ $X2=3.492 $Y2=2.24
r70 21 34 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.5
+ $X2=2.645 $Y2=1.665
r71 21 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.5
+ $X2=2.645 $Y2=1.335
r72 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.5 $X2=2.645 $Y2=1.5
r73 18 31 1.87921 $w=3.3e-07 $l=2.17e-07 $layer=LI1_cond $X=3.275 $Y=1.5
+ $X2=3.492 $Y2=1.5
r74 18 20 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=3.275 $Y=1.5
+ $X2=2.645 $Y2=1.5
r75 17 33 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.555 $Y=0.88
+ $X2=2.555 $Y2=1.335
r76 16 17 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.54 $Y=0.73
+ $X2=2.54 $Y2=0.88
r77 14 34 231.062 $w=2.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.605 $Y=2.595
+ $X2=2.605 $Y2=1.665
r78 9 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.525 $Y=0.445
+ $X2=2.525 $Y2=0.73
r79 2 25 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.3
+ $Y=2.095 $X2=3.44 $Y2=2.24
r80 1 29 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.235 $X2=3.545 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP2%VPWR 1 2 7 9 13 18 19 20 30 31
r42 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 24 27 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 22 34 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r50 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 20 25 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 18 27 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.87 $Y2=3.33
r55 17 30 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.87 $Y2=3.33
r57 13 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.87 $Y=2.24 $X2=2.87
+ $Y2=2.95
r58 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=3.33
r59 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.87 $Y=3.245
+ $X2=2.87 $Y2=2.95
r60 7 34 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.212 $Y2=3.33
r61 7 9 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=0.3 $Y=3.245 $X2=0.3
+ $Y2=2.44
r62 2 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.095 $X2=2.87 $Y2=2.95
r63 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.095 $X2=2.87 $Y2=2.24
r64 1 9 300 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=2.095 $X2=0.34 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP2%Y 1 2 8 9 10 11 12 14 15 17 19 20 23 26 27
+ 36 44
c84 36 0 7.69208e-20 $X=0.96 $Y=2.45
r85 36 44 1.54255 $w=7.1e-07 $l=4.5e-08 $layer=LI1_cond $X=0.96 $Y=2.45 $X2=0.96
+ $Y2=2.405
r86 26 44 0.456075 $w=5.35e-07 $l=2e-08 $layer=LI1_cond $X=0.96 $Y=2.385
+ $X2=0.96 $Y2=2.405
r87 26 27 5.13808 $w=7.08e-07 $l=3.05e-07 $layer=LI1_cond $X=0.96 $Y=2.47
+ $X2=0.96 $Y2=2.775
r88 26 36 0.336923 $w=7.08e-07 $l=2e-08 $layer=LI1_cond $X=0.96 $Y=2.47 $X2=0.96
+ $Y2=2.45
r89 25 27 2.02154 $w=7.08e-07 $l=1.2e-07 $layer=LI1_cond $X=0.96 $Y=2.895
+ $X2=0.96 $Y2=2.775
r90 21 23 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.66 $Y=2.895 $X2=1.66
+ $Y2=2.495
r91 20 25 10.8756 $w=1.7e-07 $l=3.95221e-07 $layer=LI1_cond $X=1.315 $Y=2.98
+ $X2=0.96 $Y2=2.895
r92 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.495 $Y=2.98
+ $X2=1.66 $Y2=2.895
r93 19 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.495 $Y=2.98
+ $X2=1.315 $Y2=2.98
r94 15 17 33.5062 $w=2.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.03 $Y=0.4
+ $X2=1.815 $Y2=0.4
r95 13 15 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.945 $Y=0.535
+ $X2=1.03 $Y2=0.4
r96 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.945 $Y=0.535
+ $X2=0.945 $Y2=0.725
r97 11 26 8.5514 $w=5.35e-07 $l=5.23211e-07 $layer=LI1_cond $X=0.605 $Y=2.01
+ $X2=0.96 $Y2=2.385
r98 11 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.605 $Y=2.01
+ $X2=0.26 $Y2=2.01
r99 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.86 $Y=0.81
+ $X2=0.945 $Y2=0.725
r100 9 10 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.86 $Y=0.81 $X2=0.26
+ $Y2=0.81
r101 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.175 $Y=1.925
+ $X2=0.26 $Y2=2.01
r102 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.175 $Y=0.895
+ $X2=0.26 $Y2=0.81
r103 7 8 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.175 $Y=0.895
+ $X2=0.175 $Y2=1.925
r104 2 23 300 $w=1.7e-07 $l=5.97411e-07 $layer=licon1_PDIFF $count=2 $X=1.23
+ $Y=2.095 $X2=1.66 $Y2=2.495
r105 1 17 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.235 $X2=1.815 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_LP2%VGND 1 2 9 13 16 17 18 24 30 31 34
c54 30 0 9.7113e-20 $X=3.6 $Y=0
r55 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r57 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.745
+ $Y2=0
r59 28 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=3.6
+ $Y2=0
r60 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.745
+ $Y2=0
r62 24 26 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=2.58 $Y=0 $X2=0.72
+ $Y2=0
r63 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r64 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 18 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r66 18 27 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.72
+ $Y2=0
r67 16 21 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.24
+ $Y2=0
r68 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.515
+ $Y2=0
r69 15 26 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.68 $Y=0 $X2=0.72
+ $Y2=0
r70 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0 $X2=0.515
+ $Y2=0
r71 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=0.085
+ $X2=2.745 $Y2=0
r72 11 13 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.745 $Y=0.085
+ $X2=2.745 $Y2=0.415
r73 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.515 $Y=0.085
+ $X2=0.515 $Y2=0
r74 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.515 $Y=0.085
+ $X2=0.515 $Y2=0.38
r75 2 13 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.235 $X2=2.745 $Y2=0.415
r76 1 9 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.37
+ $Y=0.235 $X2=0.515 $Y2=0.38
.ends

