* File: sky130_fd_sc_lp__a2bb2oi_lp.pex.spice
* Created: Wed Sep  2 09:24:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%B1 3 7 9 10 16
r29 14 16 7.24812 $w=2.66e-07 $l=4e-08 $layer=POLY_cond $X=0.505 $Y=0.975
+ $X2=0.545 $Y2=0.975
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.505
+ $Y=0.975 $X2=0.505 $Y2=0.975
r31 10 15 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.72 $Y=0.975
+ $X2=0.505 $Y2=0.975
r32 9 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=0.975
+ $X2=0.505 $Y2=0.975
r33 5 16 41.6767 $w=2.66e-07 $l=3.01413e-07 $layer=POLY_cond $X=0.775 $Y=0.81
+ $X2=0.545 $Y2=0.975
r34 5 7 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.775 $Y=0.81
+ $X2=0.775 $Y2=0.445
r35 1 16 4.31405 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.14
+ $X2=0.545 $Y2=0.975
r36 1 3 349.077 $w=2.5e-07 $l=1.405e-06 $layer=POLY_cond $X=0.545 $Y=1.14
+ $X2=0.545 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%B2 3 7 9 10 11 16
c36 16 0 3.5105e-19 $X=1.075 $Y=1.615
c37 3 0 1.49773e-19 $X=1.075 $Y=2.545
r38 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.615
+ $X2=1.075 $Y2=1.45
r39 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.615 $X2=1.075 $Y2=1.615
r40 11 17 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.075 $Y2=1.615
r41 10 17 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=1.075 $Y2=1.615
r42 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.72 $Y2=1.615
r43 7 18 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.165 $Y=0.445
+ $X2=1.165 $Y2=1.45
r44 1 16 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.78
+ $X2=1.075 $Y2=1.615
r45 1 3 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.075 $Y=1.78
+ $X2=1.075 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_296_146# 1 2 8 11 13 15 17 18 20 22 24
+ 25 26 27 28 32 37 39 44 48 50
c102 27 0 6.45857e-20 $X=1.605 $Y=1.695
c103 11 0 8.82946e-20 $X=1.605 $Y=1.82
r104 46 48 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.97 $Y=0.43
+ $X2=3.11 $Y2=0.43
r105 40 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.01 $Y=1.29 $X2=2.01
+ $Y2=1.2
r106 39 42 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.01 $Y=1.29 $X2=2.01
+ $Y2=1.37
r107 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.01
+ $Y=1.29 $X2=2.01 $Y2=1.29
r108 37 44 3.70735 $w=2.5e-07 $l=1.54771e-07 $layer=LI1_cond $X=3.11 $Y=1.285
+ $X2=2.992 $Y2=1.37
r109 36 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=0.595
+ $X2=3.11 $Y2=0.43
r110 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.11 $Y=0.595
+ $X2=3.11 $Y2=1.285
r111 32 34 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.955 $Y=1.84
+ $X2=2.955 $Y2=2.55
r112 30 44 3.70735 $w=2.5e-07 $l=1.01833e-07 $layer=LI1_cond $X=2.955 $Y=1.455
+ $X2=2.992 $Y2=1.37
r113 30 32 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.955 $Y=1.455
+ $X2=2.955 $Y2=1.84
r114 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.37
+ $X2=2.01 $Y2=1.37
r115 28 44 2.76166 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.79 $Y=1.37
+ $X2=2.992 $Y2=1.37
r116 28 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.79 $Y=1.37
+ $X2=2.175 $Y2=1.37
r117 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.955 $Y=0.73
+ $X2=1.955 $Y2=0.445
r118 21 25 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=1.67 $Y=0.805
+ $X2=1.575 $Y2=0.805
r119 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.88 $Y=0.805
+ $X2=1.955 $Y2=0.73
r120 20 21 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.88 $Y=0.805
+ $X2=1.67 $Y2=0.805
r121 19 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.63 $Y=1.2
+ $X2=1.555 $Y2=1.2
r122 18 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.2
+ $X2=2.01 $Y2=1.2
r123 18 19 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.845 $Y=1.2
+ $X2=1.63 $Y2=1.2
r124 15 25 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=1.595 $Y=0.73
+ $X2=1.575 $Y2=0.805
r125 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.595 $Y=0.73
+ $X2=1.595 $Y2=0.445
r126 11 27 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.605 $Y=1.82
+ $X2=1.605 $Y2=1.695
r127 11 13 180.129 $w=2.5e-07 $l=7.25e-07 $layer=POLY_cond $X=1.605 $Y=1.82
+ $X2=1.605 $Y2=2.545
r128 9 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.555 $Y=1.275
+ $X2=1.555 $Y2=1.2
r129 9 27 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.555 $Y=1.275
+ $X2=1.555 $Y2=1.695
r130 8 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.555 $Y=1.125
+ $X2=1.555 $Y2=1.2
r131 7 25 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=1.555 $Y=0.88
+ $X2=1.575 $Y2=0.805
r132 7 8 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.555 $Y=0.88
+ $X2=1.555 $Y2=1.125
r133 2 34 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.695 $X2=2.955 $Y2=2.55
r134 2 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.695 $X2=2.955 $Y2=1.84
r135 1 46 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.235 $X2=2.97 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%A2_N 1 3 6 8 10 11 17
c47 17 0 1.20711e-19 $X=2.69 $Y=0.92
r48 17 18 10.8785 $w=2.88e-07 $l=6.5e-08 $layer=POLY_cond $X=2.69 $Y=0.92
+ $X2=2.755 $Y2=0.92
r49 15 17 1.67361 $w=2.88e-07 $l=1e-08 $layer=POLY_cond $X=2.68 $Y=0.92 $X2=2.69
+ $Y2=0.92
r50 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=0.94 $X2=2.68 $Y2=0.94
r51 8 18 18.0107 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=2.755 $Y=0.735
+ $X2=2.755 $Y2=0.92
r52 8 10 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.755 $Y=0.735
+ $X2=2.755 $Y2=0.445
r53 4 17 6.18571 $w=2.5e-07 $l=1.85e-07 $layer=POLY_cond $X=2.69 $Y=1.105
+ $X2=2.69 $Y2=0.92
r54 4 6 270.814 $w=2.5e-07 $l=1.09e-06 $layer=POLY_cond $X=2.69 $Y=1.105
+ $X2=2.69 $Y2=2.195
r55 1 15 47.6979 $w=2.88e-07 $l=3.65992e-07 $layer=POLY_cond $X=2.395 $Y=0.735
+ $X2=2.68 $Y2=0.92
r56 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.395 $Y=0.735
+ $X2=2.395 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%A1_N 3 5 6 9 13 16 17 18 20 27
r46 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.64
+ $Y=1.275 $X2=3.64 $Y2=1.275
r47 20 28 7.85484 $w=6.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.08 $Y=1.445
+ $X2=3.64 $Y2=1.445
r48 18 28 0.714077 $w=6.68e-07 $l=4e-08 $layer=LI1_cond $X=3.6 $Y=1.445 $X2=3.64
+ $Y2=1.445
r49 17 27 58.221 $w=3.35e-07 $l=3.38e-07 $layer=POLY_cond $X=3.637 $Y=1.613
+ $X2=3.637 $Y2=1.275
r50 15 27 2.58377 $w=3.35e-07 $l=1.5e-08 $layer=POLY_cond $X=3.637 $Y=1.26
+ $X2=3.637 $Y2=1.275
r51 15 16 13.4622 $w=2.42e-07 $l=7.5e-08 $layer=POLY_cond $X=3.637 $Y=1.26
+ $X2=3.637 $Y2=1.185
r52 11 17 47.2295 $w=2.98e-07 $l=3.56399e-07 $layer=POLY_cond $X=3.78 $Y=1.905
+ $X2=3.637 $Y2=1.613
r53 11 13 159.01 $w=2.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.78 $Y=1.905
+ $X2=3.78 $Y2=2.545
r54 7 16 13.4622 $w=2.42e-07 $l=1.23952e-07 $layer=POLY_cond $X=3.545 $Y=1.11
+ $X2=3.637 $Y2=1.185
r55 7 9 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.545 $Y=1.11
+ $X2=3.545 $Y2=0.445
r56 5 16 12.3158 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=3.47 $Y=1.185
+ $X2=3.637 $Y2=1.185
r57 5 6 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.47 $Y=1.185 $X2=3.26
+ $Y2=1.185
r58 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.185 $Y=1.11
+ $X2=3.26 $Y2=1.185
r59 1 3 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.185 $Y=1.11
+ $X2=3.185 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_27_409# 1 2 9 13 14 17
r27 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.34 $Y=2.19 $X2=1.34
+ $Y2=2.9
r28 15 17 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.34 $Y=2.155
+ $X2=1.34 $Y2=2.19
r29 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.175 $Y=2.07
+ $X2=1.34 $Y2=2.155
r30 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.175 $Y=2.07
+ $X2=0.445 $Y2=2.07
r31 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.19 $X2=0.28
+ $Y2=2.9
r32 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.155
+ $X2=0.445 $Y2=2.07
r33 7 9 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.28 $Y=2.155 $X2=0.28
+ $Y2=2.19
r34 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.9
r35 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.19
r36 1 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r37 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%VPWR 1 2 11 13 15 19 21 30 34
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r40 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r42 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 24 27 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 24 25 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 22 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r47 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 21 33 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.88 $Y=3.33 $X2=4.1
+ $Y2=3.33
r49 21 27 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.88 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 19 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 19 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.045 $Y=2.19
+ $X2=4.045 $Y2=2.9
r53 13 33 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.045 $Y=3.245
+ $X2=4.1 $Y2=3.33
r54 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.045 $Y=3.245
+ $X2=4.045 $Y2=2.9
r55 9 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245 $X2=0.81
+ $Y2=3.33
r56 9 11 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.5
r57 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=2.045 $X2=4.045 $Y2=2.9
r58 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=2.045 $X2=4.045 $Y2=2.19
r59 1 11 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.5
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%Y 1 2 8 9 11 19 20
c49 9 0 3.02033e-19 $X=1.87 $Y=1.805
c50 8 0 4.07795e-19 $X=1.58 $Y=1.635
r51 27 28 5.62167 $w=4.08e-07 $l=2e-07 $layer=LI1_cond $X=1.38 $Y=0.47 $X2=1.58
+ $Y2=0.47
r52 20 28 2.81084 $w=4.08e-07 $l=1e-07 $layer=LI1_cond $X=1.68 $Y=0.47 $X2=1.58
+ $Y2=0.47
r53 19 27 5.05951 $w=4.08e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=0.47 $X2=1.38
+ $Y2=0.47
r54 11 13 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.87 $Y=2.19 $X2=1.87
+ $Y2=2.9
r55 9 15 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.87 $Y=1.72 $X2=1.58
+ $Y2=1.72
r56 9 11 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.87 $Y=1.805
+ $X2=1.87 $Y2=2.19
r57 8 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=1.635
+ $X2=1.58 $Y2=1.72
r58 7 28 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.58 $Y=0.675
+ $X2=1.58 $Y2=0.47
r59 7 8 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.58 $Y=0.675 $X2=1.58
+ $Y2=1.635
r60 2 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=2.045 $X2=1.87 $Y2=2.9
r61 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=2.045 $X2=1.87 $Y2=2.19
r62 1 27 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.24
+ $Y=0.235 $X2=1.38 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%A_456_339# 1 2 9 13 14 15 17
c29 9 0 6.45857e-20 $X=2.425 $Y=1.84
r30 15 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.895
+ $X2=3.515 $Y2=2.98
r31 15 17 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=3.515 $Y=2.895
+ $X2=3.515 $Y2=2.19
r32 13 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.35 $Y=2.98
+ $X2=3.515 $Y2=2.98
r33 13 14 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.35 $Y=2.98
+ $X2=2.59 $Y2=2.98
r34 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.425 $Y=1.84
+ $X2=2.425 $Y2=2.55
r35 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.425 $Y=2.895
+ $X2=2.59 $Y2=2.98
r36 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.425 $Y=2.895
+ $X2=2.425 $Y2=2.55
r37 2 20 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=2.045 $X2=3.515 $Y2=2.9
r38 2 17 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=2.045 $X2=3.515 $Y2=2.19
r39 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.695 $X2=2.425 $Y2=2.55
r40 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.695 $X2=2.425 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_LP%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45
+ 48 51
r61 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r62 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r63 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r64 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r65 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.76
+ $Y2=0
r66 39 41 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.08
+ $Y2=0
r67 38 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r68 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r69 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.17
+ $Y2=0
r70 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.64
+ $Y2=0
r71 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0 $X2=3.76
+ $Y2=0
r72 34 37 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.595 $Y=0 $X2=2.64
+ $Y2=0
r73 33 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r74 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r75 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.56
+ $Y2=0
r76 30 32 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=1.68
+ $Y2=0
r77 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.17
+ $Y2=0
r78 29 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.68
+ $Y2=0
r79 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r80 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r81 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.56
+ $Y2=0
r82 24 26 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.24
+ $Y2=0
r83 22 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r84 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r85 22 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r86 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0
r87 18 20 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0.445
r88 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0
r89 14 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0.445
r90 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0
r91 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0.42
r92 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.62
+ $Y=0.235 $X2=3.76 $Y2=0.445
r93 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.03
+ $Y=0.235 $X2=2.17 $Y2=0.445
r94 1 12 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.415
+ $Y=0.235 $X2=0.56 $Y2=0.42
.ends

