* File: sky130_fd_sc_lp__decap_8.pex.spice
* Created: Wed Sep  2 09:42:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAP_8%VGND 1 12 15 17 18 22 26 30 31 41 42 45 48
r27 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r28 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r29 42 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r30 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r31 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.095
+ $Y2=0
r32 39 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.6
+ $Y2=0
r33 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r34 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r36 34 37 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r37 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r39 32 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r40 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=0 $X2=3.095
+ $Y2=0
r41 31 37 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.93 $Y=0 $X2=2.64
+ $Y2=0
r42 26 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r43 26 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r44 22 24 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.095 $Y=0.36
+ $X2=3.095 $Y2=1.04
r45 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0
r46 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0.36
r47 18 30 22.4154 $w=1.774e-06 $l=1.03959e-06 $layer=POLY_cond $X=1.395 $Y=1.77
+ $X2=1.88 $Y2=2.595
r48 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.395
+ $Y=1.77 $X2=1.395 $Y2=1.77
r49 15 17 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.98 $Y=1.77
+ $X2=1.395 $Y2=1.77
r50 12 14 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.815 $Y=0.38
+ $X2=0.815 $Y2=1.06
r51 10 15 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.98 $Y2=1.77
r52 10 14 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.815 $Y2=1.06
r53 9 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r54 9 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.38
r55 1 24 121.333 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.095 $Y2=1.04
r56 1 22 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.095 $Y2=0.36
r57 1 14 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=0.815 $Y2=1.06
r58 1 12 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=0.815 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAP_8%VPWR 1 9 13 16 24 28 29 30 33 35 48 49 52
r27 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r29 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r30 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 43 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 42 45 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 40 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r35 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.2 $Y2=3.33
r36 38 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 35 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r39 35 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 30 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 30 43 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 28 45 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.03 $Y2=3.33
r44 27 48 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.03 $Y2=3.33
r46 24 26 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.03 $Y=2.29
+ $X2=3.03 $Y2=2.97
r47 22 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=3.33
r48 22 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=2.97
r49 21 24 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.03 $Y=1.675
+ $X2=3.03 $Y2=2.29
r50 16 33 20.7068 $w=1.804e-06 $l=7.75e-07 $layer=POLY_cond $X=1.96 $Y=1.51
+ $X2=1.96 $Y2=0.735
r51 16 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=1.51 $X2=2.8 $Y2=1.51
r52 15 19 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=2.12 $Y=1.507
+ $X2=2.8 $Y2=1.507
r53 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.12
+ $Y=1.51 $X2=2.12 $Y2=1.51
r54 13 21 6.81699 $w=3.35e-07 $l=2.36525e-07 $layer=LI1_cond $X=2.865 $Y=1.507
+ $X2=3.03 $Y2=1.675
r55 13 19 2.23608 $w=3.33e-07 $l=6.5e-08 $layer=LI1_cond $X=2.865 $Y=1.507
+ $X2=2.8 $Y2=1.507
r56 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.74 $Y=2.27 $X2=0.74
+ $Y2=2.95
r57 7 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=3.33
r58 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=2.95
r59 1 26 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=3.03 $Y2=2.97
r60 1 24 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=3.03 $Y2=2.29
r61 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=0.74 $Y2=2.95
r62 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=2.095 $X2=0.74 $Y2=2.27
.ends

