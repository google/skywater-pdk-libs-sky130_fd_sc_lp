* File: sky130_fd_sc_lp__o21bai_4.pxi.spice
* Created: Wed Sep  2 10:17:43 2020
* 
x_PM_SKY130_FD_SC_LP__O21BAI_4%B1_N N_B1_N_M1009_g N_B1_N_c_108_n N_B1_N_M1024_g
+ B1_N N_B1_N_c_109_n PM_SKY130_FD_SC_LP__O21BAI_4%B1_N
x_PM_SKY130_FD_SC_LP__O21BAI_4%A_27_49# N_A_27_49#_M1009_s N_A_27_49#_M1024_s
+ N_A_27_49#_M1006_g N_A_27_49#_c_148_n N_A_27_49#_M1001_g N_A_27_49#_M1008_g
+ N_A_27_49#_c_149_n N_A_27_49#_M1003_g N_A_27_49#_M1015_g N_A_27_49#_c_150_n
+ N_A_27_49#_M1011_g N_A_27_49#_M1018_g N_A_27_49#_c_151_n N_A_27_49#_M1021_g
+ N_A_27_49#_c_141_n N_A_27_49#_c_152_n N_A_27_49#_c_153_n N_A_27_49#_c_142_n
+ N_A_27_49#_c_143_n N_A_27_49#_c_164_n N_A_27_49#_c_154_n N_A_27_49#_c_183_p
+ N_A_27_49#_c_144_n N_A_27_49#_c_208_p N_A_27_49#_c_145_n N_A_27_49#_c_146_n
+ N_A_27_49#_c_147_n PM_SKY130_FD_SC_LP__O21BAI_4%A_27_49#
x_PM_SKY130_FD_SC_LP__O21BAI_4%A1 N_A1_M1004_g N_A1_M1002_g N_A1_M1013_g
+ N_A1_M1005_g N_A1_M1019_g N_A1_M1020_g N_A1_M1023_g N_A1_M1022_g N_A1_c_278_n
+ N_A1_c_270_n N_A1_c_290_p N_A1_c_287_n N_A1_c_280_n A1 A1 A1 N_A1_c_273_n
+ PM_SKY130_FD_SC_LP__O21BAI_4%A1
x_PM_SKY130_FD_SC_LP__O21BAI_4%A2 N_A2_M1007_g N_A2_M1000_g N_A2_M1014_g
+ N_A2_M1010_g N_A2_M1017_g N_A2_M1012_g N_A2_M1025_g N_A2_M1016_g A2 A2 A2
+ N_A2_c_388_n N_A2_c_389_n PM_SKY130_FD_SC_LP__O21BAI_4%A2
x_PM_SKY130_FD_SC_LP__O21BAI_4%VPWR N_VPWR_M1024_d N_VPWR_M1003_d N_VPWR_M1021_d
+ N_VPWR_M1013_s N_VPWR_M1023_s N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n
+ N_VPWR_c_471_n N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_503_n
+ N_VPWR_c_475_n N_VPWR_c_476_n N_VPWR_c_477_n N_VPWR_c_478_n VPWR
+ N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n N_VPWR_c_482_n N_VPWR_c_483_n
+ N_VPWR_c_467_n PM_SKY130_FD_SC_LP__O21BAI_4%VPWR
x_PM_SKY130_FD_SC_LP__O21BAI_4%Y N_Y_M1006_s N_Y_M1015_s N_Y_M1001_s N_Y_M1011_s
+ N_Y_M1007_d N_Y_M1017_d N_Y_c_625_n N_Y_c_572_n N_Y_c_573_n N_Y_c_582_n
+ N_Y_c_584_n N_Y_c_591_n N_Y_c_630_n N_Y_c_592_n N_Y_c_618_n N_Y_c_593_n
+ N_Y_c_595_n N_Y_c_596_n Y Y Y N_Y_c_571_n PM_SKY130_FD_SC_LP__O21BAI_4%Y
x_PM_SKY130_FD_SC_LP__O21BAI_4%A_653_367# N_A_653_367#_M1004_d
+ N_A_653_367#_M1014_s N_A_653_367#_M1025_s N_A_653_367#_M1019_d
+ N_A_653_367#_c_655_n N_A_653_367#_c_656_n N_A_653_367#_c_669_n
+ N_A_653_367#_c_657_n N_A_653_367#_c_662_n N_A_653_367#_c_681_n
+ PM_SKY130_FD_SC_LP__O21BAI_4%A_653_367#
x_PM_SKY130_FD_SC_LP__O21BAI_4%VGND N_VGND_M1009_d N_VGND_M1002_d N_VGND_M1010_s
+ N_VGND_M1016_s N_VGND_M1020_d N_VGND_c_688_n N_VGND_c_689_n N_VGND_c_690_n
+ N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n N_VGND_c_694_n N_VGND_c_695_n
+ N_VGND_c_696_n N_VGND_c_697_n VGND N_VGND_c_698_n N_VGND_c_699_n
+ N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n N_VGND_c_704_n
+ PM_SKY130_FD_SC_LP__O21BAI_4%VGND
x_PM_SKY130_FD_SC_LP__O21BAI_4%A_218_49# N_A_218_49#_M1006_d N_A_218_49#_M1008_d
+ N_A_218_49#_M1018_d N_A_218_49#_M1000_d N_A_218_49#_M1012_d
+ N_A_218_49#_M1005_s N_A_218_49#_M1022_s N_A_218_49#_c_798_n
+ N_A_218_49#_c_854_n N_A_218_49#_c_802_n N_A_218_49#_c_787_n
+ N_A_218_49#_c_788_n N_A_218_49#_c_858_n N_A_218_49#_c_789_n
+ N_A_218_49#_c_862_n N_A_218_49#_c_790_n N_A_218_49#_c_866_n
+ N_A_218_49#_c_791_n N_A_218_49#_c_792_n N_A_218_49#_c_793_n
+ N_A_218_49#_c_794_n N_A_218_49#_c_795_n N_A_218_49#_c_796_n
+ PM_SKY130_FD_SC_LP__O21BAI_4%A_218_49#
cc_1 VNB N_B1_N_M1009_g 0.0351385f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.665
cc_2 VNB N_B1_N_c_108_n 0.0334109f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.675
cc_3 VNB N_B1_N_c_109_n 0.00973638f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_4 VNB N_A_27_49#_M1006_g 0.0276493f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_5 VNB N_A_27_49#_M1008_g 0.0219184f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.665
cc_6 VNB N_A_27_49#_M1015_g 0.0213478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_49#_M1018_g 0.0229333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_49#_c_141_n 0.0311092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_49#_c_142_n 0.0065888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_49#_c_143_n 0.011422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_49#_c_144_n 0.00229744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_49#_c_145_n 0.0102904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_49#_c_146_n 0.0409204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_49#_c_147_n 0.0638563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1002_g 0.0237103f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.465
cc_16 VNB N_A1_M1013_g 0.00123444f $X=-0.19 $Y=-0.245 $X2=0.412 $Y2=1.51
cc_17 VNB N_A1_M1005_g 0.0202052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1019_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1020_g 0.0200544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_M1023_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_M1022_g 0.0271791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_270_n 0.0255504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB A1 0.00253791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB A1 0.011363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_273_n 0.0923189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_M1000_g 0.0226534f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.465
cc_27 VNB N_A2_M1010_g 0.02243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_M1012_g 0.02243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A2_M1016_g 0.022801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_c_388_n 0.00187959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_389_n 0.0652967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_467_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_571_n 0.00545388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_688_n 0.00943014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_689_n 6.09197e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_690_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_691_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_692_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_693_n 6.09197e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_694_n 0.0556652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_695_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_696_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_697_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_698_n 0.0154417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_699_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_700_n 0.0163964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_701_n 0.338012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_702_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_703_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_704_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_218_49#_c_787_n 0.00760991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_218_49#_c_788_n 0.00604846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_218_49#_c_789_n 0.00322376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_218_49#_c_790_n 0.0101655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_218_49#_c_791_n 0.0119591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_218_49#_c_792_n 0.0296037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_218_49#_c_793_n 0.00714562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_218_49#_c_794_n 0.00152782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_218_49#_c_795_n 0.00174672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_218_49#_c_796_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VPB N_B1_N_c_108_n 0.00843721f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.675
cc_62 VPB N_B1_N_M1024_g 0.0276521f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.465
cc_63 VPB N_B1_N_c_109_n 0.00677036f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_64 VPB N_A_27_49#_c_148_n 0.0197819f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=1.51
cc_65 VPB N_A_27_49#_c_149_n 0.0152836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_27_49#_c_150_n 0.0151645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_27_49#_c_151_n 0.0160412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_27_49#_c_152_n 0.00773819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_27_49#_c_153_n 0.0374933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_27_49#_c_154_n 0.0025667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_27_49#_c_146_n 0.0199148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_27_49#_c_147_n 0.0196434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A1_M1004_g 0.0179515f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.665
cc_74 VPB N_A1_M1013_g 0.0185521f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=1.51
cc_75 VPB N_A1_M1019_g 0.0187176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A1_M1023_g 0.0245572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A1_c_278_n 0.00255692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A1_c_270_n 0.00645295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A1_c_280_n 7.51442e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB A1 9.27404e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB A1 0.0163983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A2_M1007_g 0.0183228f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.665
cc_83 VPB N_A2_M1014_g 0.0181366f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=1.51
cc_84 VPB N_A2_M1017_g 0.0181378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A2_M1025_g 0.0187401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A2_c_388_n 0.00884706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A2_c_389_n 0.0122315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_468_n 0.00715536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_469_n 0.0015455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_470_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_471_n 0.00252657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_472_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_473_n 0.0117752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_474_n 0.0478673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_475_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_476_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_477_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_478_n 0.00452958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_479_n 0.0189574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_480_n 0.0534875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_481_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_482_n 0.0139193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_483_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_467_n 0.048694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_Y_c_572_n 0.00286079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_Y_c_573_n 0.00272989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 N_B1_N_c_108_n N_A_27_49#_c_152_n 0.00130813f $X=0.53 $Y=1.675 $X2=0
+ $Y2=0
cc_108 N_B1_N_c_109_n N_A_27_49#_c_152_n 0.0231956f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_109 N_B1_N_M1009_g N_A_27_49#_c_142_n 0.0165745f $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_110 N_B1_N_c_108_n N_A_27_49#_c_142_n 0.00318784f $X=0.53 $Y=1.675 $X2=0
+ $Y2=0
cc_111 N_B1_N_c_109_n N_A_27_49#_c_142_n 0.0141065f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_112 N_B1_N_c_108_n N_A_27_49#_c_143_n 0.00342128f $X=0.53 $Y=1.675 $X2=0
+ $Y2=0
cc_113 N_B1_N_c_109_n N_A_27_49#_c_143_n 0.01718f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_114 N_B1_N_M1024_g N_A_27_49#_c_164_n 0.0159303f $X=0.53 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B1_N_c_109_n N_A_27_49#_c_164_n 0.00715924f $X=0.385 $Y=1.51 $X2=0
+ $Y2=0
cc_116 N_B1_N_M1024_g N_A_27_49#_c_154_n 0.00397226f $X=0.53 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_B1_N_M1009_g N_A_27_49#_c_145_n 0.00566885f $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_118 N_B1_N_c_108_n N_A_27_49#_c_145_n 0.00397226f $X=0.53 $Y=1.675 $X2=0
+ $Y2=0
cc_119 N_B1_N_c_109_n N_A_27_49#_c_145_n 0.0223655f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_120 N_B1_N_M1009_g N_A_27_49#_c_146_n 0.00789768f $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_121 N_B1_N_c_108_n N_A_27_49#_c_146_n 0.0143414f $X=0.53 $Y=1.675 $X2=0 $Y2=0
cc_122 N_B1_N_c_109_n N_A_27_49#_c_146_n 3.30438e-19 $X=0.385 $Y=1.51 $X2=0
+ $Y2=0
cc_123 N_B1_N_M1024_g N_VPWR_c_468_n 0.00814732f $X=0.53 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B1_N_M1024_g N_VPWR_c_469_n 0.00318901f $X=0.53 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B1_N_M1024_g N_VPWR_c_479_n 0.00585385f $X=0.53 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_N_M1024_g N_VPWR_c_467_n 0.0128027f $X=0.53 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B1_N_M1009_g N_VGND_c_688_n 0.0143488f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_128 N_B1_N_M1009_g N_VGND_c_698_n 0.00477554f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_129 N_B1_N_M1009_g N_VGND_c_701_n 0.00919076f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_130 N_B1_N_M1009_g N_A_218_49#_c_793_n 0.00122188f $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_131 N_A_27_49#_c_147_n N_A1_M1004_g 0.0429924f $X=2.72 $Y=1.525 $X2=0 $Y2=0
cc_132 N_A_27_49#_M1018_g N_A1_M1002_g 0.0178358f $X=2.72 $Y=0.665 $X2=0 $Y2=0
cc_133 N_A_27_49#_c_147_n N_A1_c_278_n 0.00295816f $X=2.72 $Y=1.525 $X2=0 $Y2=0
cc_134 N_A_27_49#_c_147_n N_A1_c_270_n 0.0222288f $X=2.72 $Y=1.525 $X2=0 $Y2=0
cc_135 N_A_27_49#_c_151_n N_A1_c_287_n 0.00134835f $X=2.72 $Y=1.725 $X2=0 $Y2=0
cc_136 N_A_27_49#_c_164_n N_VPWR_M1024_d 0.0095894f $X=0.76 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_27_49#_c_154_n N_VPWR_M1024_d 0.00210203f $X=0.845 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_27_49#_c_148_n N_VPWR_c_469_n 0.0073184f $X=1.43 $Y=1.725 $X2=0 $Y2=0
cc_139 N_A_27_49#_c_164_n N_VPWR_c_469_n 0.0141597f $X=0.76 $Y=2.015 $X2=0 $Y2=0
cc_140 N_A_27_49#_c_154_n N_VPWR_c_469_n 0.00781998f $X=0.845 $Y=1.93 $X2=0
+ $Y2=0
cc_141 N_A_27_49#_c_183_p N_VPWR_c_469_n 0.00620234f $X=1.175 $Y=1.49 $X2=0
+ $Y2=0
cc_142 N_A_27_49#_c_144_n N_VPWR_c_469_n 0.0138968f $X=1.38 $Y=1.47 $X2=0 $Y2=0
cc_143 N_A_27_49#_c_146_n N_VPWR_c_469_n 0.00626629f $X=1.355 $Y=1.525 $X2=0
+ $Y2=0
cc_144 N_A_27_49#_c_148_n N_VPWR_c_470_n 7.40567e-19 $X=1.43 $Y=1.725 $X2=0
+ $Y2=0
cc_145 N_A_27_49#_c_149_n N_VPWR_c_470_n 0.0142198f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_146 N_A_27_49#_c_150_n N_VPWR_c_470_n 0.0141063f $X=2.29 $Y=1.725 $X2=0 $Y2=0
cc_147 N_A_27_49#_c_151_n N_VPWR_c_470_n 7.55739e-19 $X=2.72 $Y=1.725 $X2=0
+ $Y2=0
cc_148 N_A_27_49#_c_150_n N_VPWR_c_471_n 5.54101e-19 $X=2.29 $Y=1.725 $X2=0
+ $Y2=0
cc_149 N_A_27_49#_c_151_n N_VPWR_c_471_n 0.00836395f $X=2.72 $Y=1.725 $X2=0
+ $Y2=0
cc_150 N_A_27_49#_c_164_n N_VPWR_c_503_n 0.023174f $X=0.76 $Y=2.015 $X2=0 $Y2=0
cc_151 N_A_27_49#_c_183_p N_VPWR_c_503_n 0.00510345f $X=1.175 $Y=1.49 $X2=0
+ $Y2=0
cc_152 N_A_27_49#_c_146_n N_VPWR_c_503_n 0.00369139f $X=1.355 $Y=1.525 $X2=0
+ $Y2=0
cc_153 N_A_27_49#_c_148_n N_VPWR_c_475_n 0.00585385f $X=1.43 $Y=1.725 $X2=0
+ $Y2=0
cc_154 N_A_27_49#_c_149_n N_VPWR_c_475_n 0.00486043f $X=1.86 $Y=1.725 $X2=0
+ $Y2=0
cc_155 N_A_27_49#_c_150_n N_VPWR_c_477_n 0.00486043f $X=2.29 $Y=1.725 $X2=0
+ $Y2=0
cc_156 N_A_27_49#_c_151_n N_VPWR_c_477_n 0.00486043f $X=2.72 $Y=1.725 $X2=0
+ $Y2=0
cc_157 N_A_27_49#_c_153_n N_VPWR_c_479_n 0.0190529f $X=0.315 $Y=2.91 $X2=0 $Y2=0
cc_158 N_A_27_49#_M1024_s N_VPWR_c_467_n 0.00249946f $X=0.19 $Y=1.835 $X2=0
+ $Y2=0
cc_159 N_A_27_49#_c_148_n N_VPWR_c_467_n 0.0118358f $X=1.43 $Y=1.725 $X2=0 $Y2=0
cc_160 N_A_27_49#_c_149_n N_VPWR_c_467_n 0.00824727f $X=1.86 $Y=1.725 $X2=0
+ $Y2=0
cc_161 N_A_27_49#_c_150_n N_VPWR_c_467_n 0.00824727f $X=2.29 $Y=1.725 $X2=0
+ $Y2=0
cc_162 N_A_27_49#_c_151_n N_VPWR_c_467_n 0.00445664f $X=2.72 $Y=1.725 $X2=0
+ $Y2=0
cc_163 N_A_27_49#_c_153_n N_VPWR_c_467_n 0.0113912f $X=0.315 $Y=2.91 $X2=0 $Y2=0
cc_164 N_A_27_49#_c_149_n N_Y_c_572_n 0.0130695f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A_27_49#_c_150_n N_Y_c_572_n 0.0114659f $X=2.29 $Y=1.725 $X2=0 $Y2=0
cc_166 N_A_27_49#_c_208_p N_Y_c_572_n 0.0304855f $X=2 $Y=1.49 $X2=0 $Y2=0
cc_167 N_A_27_49#_c_147_n N_Y_c_572_n 0.00275588f $X=2.72 $Y=1.525 $X2=0 $Y2=0
cc_168 N_A_27_49#_c_148_n N_Y_c_573_n 0.00126637f $X=1.43 $Y=1.725 $X2=0 $Y2=0
cc_169 N_A_27_49#_c_154_n N_Y_c_573_n 0.0024893f $X=0.845 $Y=1.93 $X2=0 $Y2=0
cc_170 N_A_27_49#_c_208_p N_Y_c_573_n 0.018931f $X=2 $Y=1.49 $X2=0 $Y2=0
cc_171 N_A_27_49#_c_147_n N_Y_c_573_n 0.00287268f $X=2.72 $Y=1.525 $X2=0 $Y2=0
cc_172 N_A_27_49#_M1015_g N_Y_c_582_n 0.00274244f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_173 N_A_27_49#_M1018_g N_Y_c_582_n 0.00806402f $X=2.72 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A_27_49#_M1008_g N_Y_c_584_n 6.79845e-19 $X=1.86 $Y=0.665 $X2=0 $Y2=0
cc_175 N_A_27_49#_M1015_g N_Y_c_584_n 0.00427756f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_176 N_A_27_49#_c_150_n N_Y_c_584_n 8.67912e-19 $X=2.29 $Y=1.725 $X2=0 $Y2=0
cc_177 N_A_27_49#_M1018_g N_Y_c_584_n 0.00451889f $X=2.72 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A_27_49#_c_151_n N_Y_c_584_n 7.95638e-19 $X=2.72 $Y=1.725 $X2=0 $Y2=0
cc_179 N_A_27_49#_c_208_p N_Y_c_584_n 0.0184226f $X=2 $Y=1.49 $X2=0 $Y2=0
cc_180 N_A_27_49#_c_147_n N_Y_c_584_n 0.0350987f $X=2.72 $Y=1.525 $X2=0 $Y2=0
cc_181 N_A_27_49#_c_151_n N_Y_c_591_n 0.00755601f $X=2.72 $Y=1.725 $X2=0 $Y2=0
cc_182 N_A_27_49#_c_151_n N_Y_c_592_n 2.44127e-19 $X=2.72 $Y=1.725 $X2=0 $Y2=0
cc_183 N_A_27_49#_c_150_n N_Y_c_593_n 0.00286897f $X=2.29 $Y=1.725 $X2=0 $Y2=0
cc_184 N_A_27_49#_c_151_n N_Y_c_593_n 0.00374258f $X=2.72 $Y=1.725 $X2=0 $Y2=0
cc_185 N_A_27_49#_c_151_n N_Y_c_595_n 0.0039864f $X=2.72 $Y=1.725 $X2=0 $Y2=0
cc_186 N_A_27_49#_c_151_n N_Y_c_596_n 0.00945392f $X=2.72 $Y=1.725 $X2=0 $Y2=0
cc_187 N_A_27_49#_M1006_g N_Y_c_571_n 0.00158685f $X=1.43 $Y=0.665 $X2=0 $Y2=0
cc_188 N_A_27_49#_M1008_g N_Y_c_571_n 0.0158207f $X=1.86 $Y=0.665 $X2=0 $Y2=0
cc_189 N_A_27_49#_M1015_g N_Y_c_571_n 0.0141509f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_190 N_A_27_49#_c_208_p N_Y_c_571_n 0.047654f $X=2 $Y=1.49 $X2=0 $Y2=0
cc_191 N_A_27_49#_c_145_n N_Y_c_571_n 0.0034821f $X=0.845 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_49#_c_147_n N_Y_c_571_n 0.004937f $X=2.72 $Y=1.525 $X2=0 $Y2=0
cc_193 N_A_27_49#_c_142_n N_VGND_M1009_d 0.00166619f $X=0.76 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_27_49#_c_145_n N_VGND_M1009_d 6.49503e-19 $X=0.845 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_27_49#_M1006_g N_VGND_c_688_n 0.00339428f $X=1.43 $Y=0.665 $X2=0
+ $Y2=0
cc_196 N_A_27_49#_c_142_n N_VGND_c_688_n 0.0142339f $X=0.76 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_27_49#_c_145_n N_VGND_c_688_n 0.00852287f $X=0.845 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_27_49#_M1018_g N_VGND_c_689_n 9.56276e-19 $X=2.72 $Y=0.665 $X2=0
+ $Y2=0
cc_199 N_A_27_49#_M1006_g N_VGND_c_694_n 0.00351191f $X=1.43 $Y=0.665 $X2=0
+ $Y2=0
cc_200 N_A_27_49#_M1008_g N_VGND_c_694_n 0.00351226f $X=1.86 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_27_49#_M1015_g N_VGND_c_694_n 0.00351226f $X=2.29 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_27_49#_M1018_g N_VGND_c_694_n 0.00351226f $X=2.72 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_27_49#_c_141_n N_VGND_c_698_n 0.0178111f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_204 N_A_27_49#_M1009_s N_VGND_c_701_n 0.00368844f $X=0.135 $Y=0.245 $X2=0
+ $Y2=0
cc_205 N_A_27_49#_M1006_g N_VGND_c_701_n 0.00660265f $X=1.43 $Y=0.665 $X2=0
+ $Y2=0
cc_206 N_A_27_49#_M1008_g N_VGND_c_701_n 0.00530298f $X=1.86 $Y=0.665 $X2=0
+ $Y2=0
cc_207 N_A_27_49#_M1015_g N_VGND_c_701_n 0.00530298f $X=2.29 $Y=0.665 $X2=0
+ $Y2=0
cc_208 N_A_27_49#_M1018_g N_VGND_c_701_n 0.00545544f $X=2.72 $Y=0.665 $X2=0
+ $Y2=0
cc_209 N_A_27_49#_c_141_n N_VGND_c_701_n 0.0100304f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_210 N_A_27_49#_M1006_g N_A_218_49#_c_798_n 0.0149649f $X=1.43 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_27_49#_M1008_g N_A_218_49#_c_798_n 0.0121932f $X=1.86 $Y=0.665 $X2=0
+ $Y2=0
cc_212 N_A_27_49#_M1015_g N_A_218_49#_c_798_n 0.0121919f $X=2.29 $Y=0.665 $X2=0
+ $Y2=0
cc_213 N_A_27_49#_M1018_g N_A_218_49#_c_798_n 0.0144936f $X=2.72 $Y=0.665 $X2=0
+ $Y2=0
cc_214 N_A_27_49#_M1018_g N_A_218_49#_c_802_n 0.00474001f $X=2.72 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_27_49#_M1018_g N_A_218_49#_c_788_n 0.00122473f $X=2.72 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_27_49#_M1006_g N_A_218_49#_c_793_n 0.00787138f $X=1.43 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_27_49#_M1008_g N_A_218_49#_c_793_n 8.1291e-19 $X=1.86 $Y=0.665 $X2=0
+ $Y2=0
cc_218 N_A_27_49#_c_183_p N_A_218_49#_c_793_n 0.00557517f $X=1.175 $Y=1.49 $X2=0
+ $Y2=0
cc_219 N_A_27_49#_c_144_n N_A_218_49#_c_793_n 0.00755154f $X=1.38 $Y=1.47 $X2=0
+ $Y2=0
cc_220 N_A_27_49#_c_146_n N_A_218_49#_c_793_n 0.00365098f $X=1.355 $Y=1.525
+ $X2=0 $Y2=0
cc_221 N_A1_M1004_g N_A2_M1007_g 0.0537273f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A1_c_278_n N_A2_M1007_g 0.00428619f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_223 N_A1_c_290_p N_A2_M1007_g 0.0105687f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_224 N_A1_M1002_g N_A2_M1000_g 0.0238672f $X=3.205 $Y=0.665 $X2=0 $Y2=0
cc_225 N_A1_c_290_p N_A2_M1014_g 0.0106152f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_226 N_A1_c_290_p N_A2_M1017_g 0.0106152f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_227 N_A1_M1013_g N_A2_M1025_g 0.0217381f $X=5.34 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A1_c_290_p N_A2_M1025_g 0.0165839f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_229 N_A1_c_280_n N_A2_M1025_g 0.00106841f $X=5.35 $Y=1.93 $X2=0 $Y2=0
cc_230 N_A1_M1005_g N_A2_M1016_g 0.0213791f $X=5.355 $Y=0.665 $X2=0 $Y2=0
cc_231 N_A1_c_273_n N_A2_M1016_g 0.0110658f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_232 N_A1_M1004_g N_A2_c_388_n 2.56351e-19 $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A1_c_278_n N_A2_c_388_n 0.0263984f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_234 N_A1_c_270_n N_A2_c_388_n 0.00155711f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_235 N_A1_c_290_p N_A2_c_388_n 0.0878129f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_236 A1 N_A2_c_388_n 0.0150223f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A1_c_273_n N_A2_c_388_n 3.63024e-19 $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_238 N_A1_c_278_n N_A2_c_389_n 2.88059e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_239 N_A1_c_270_n N_A2_c_389_n 0.0211345f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_240 N_A1_c_290_p N_A2_c_389_n 0.00172102f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_241 A1 N_A2_c_389_n 0.00185963f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A1_c_273_n N_A2_c_389_n 0.0217381f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_243 N_A1_c_278_n N_VPWR_M1021_d 9.53643e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_244 N_A1_c_287_n N_VPWR_M1021_d 0.00243348f $X=3.335 $Y=2.015 $X2=0 $Y2=0
cc_245 N_A1_M1004_g N_VPWR_c_471_n 0.00316025f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A1_M1013_g N_VPWR_c_472_n 0.0116361f $X=5.34 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A1_M1019_g N_VPWR_c_472_n 0.01045f $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A1_M1023_g N_VPWR_c_472_n 5.75816e-19 $X=6.2 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A1_M1019_g N_VPWR_c_474_n 6.24191e-19 $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A1_M1023_g N_VPWR_c_474_n 0.0200733f $X=6.2 $Y=2.465 $X2=0 $Y2=0
cc_251 A1 N_VPWR_c_474_n 0.0260594f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_252 N_A1_c_273_n N_VPWR_c_474_n 0.00160096f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_253 N_A1_M1004_g N_VPWR_c_480_n 0.00547467f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_254 N_A1_M1013_g N_VPWR_c_480_n 0.00486043f $X=5.34 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A1_M1019_g N_VPWR_c_481_n 0.00486043f $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A1_M1023_g N_VPWR_c_481_n 0.00486043f $X=6.2 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A1_M1004_g N_VPWR_c_467_n 0.006232f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A1_M1013_g N_VPWR_c_467_n 0.0082726f $X=5.34 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A1_M1019_g N_VPWR_c_467_n 0.00824727f $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A1_M1023_g N_VPWR_c_467_n 0.00824727f $X=6.2 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A1_c_290_p N_Y_M1007_d 0.0034149f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_262 N_A1_c_290_p N_Y_M1017_d 0.0034149f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_263 N_A1_M1002_g N_Y_c_584_n 6.58532e-19 $X=3.205 $Y=0.665 $X2=0 $Y2=0
cc_264 N_A1_c_278_n N_Y_c_584_n 0.0171216f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_265 N_A1_c_270_n N_Y_c_584_n 0.00126633f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_266 N_A1_M1004_g N_Y_c_591_n 0.00112843f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A1_c_278_n N_Y_c_591_n 2.11117e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_268 N_A1_c_287_n N_Y_c_591_n 0.00953769f $X=3.335 $Y=2.015 $X2=0 $Y2=0
cc_269 N_A1_M1004_g N_Y_c_592_n 0.00667664f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A1_c_290_p N_Y_c_592_n 0.0781986f $X=5.265 $Y=2.015 $X2=0 $Y2=0
cc_271 N_A1_c_278_n N_Y_c_593_n 0.00966175f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_272 N_A1_M1004_g N_Y_c_596_n 0.0109084f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A1_c_270_n N_Y_c_596_n 2.68118e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_274 N_A1_c_287_n N_Y_c_596_n 0.0164189f $X=3.335 $Y=2.015 $X2=0 $Y2=0
cc_275 N_A1_c_278_n N_A_653_367#_M1004_d 0.00121536f $X=3.17 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A1_c_290_p N_A_653_367#_M1004_d 0.00745857f $X=5.265 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A1_c_290_p N_A_653_367#_M1014_s 0.0034149f $X=5.265 $Y=2.015 $X2=0
+ $Y2=0
cc_278 N_A1_c_290_p N_A_653_367#_M1025_s 0.00809843f $X=5.265 $Y=2.015 $X2=0
+ $Y2=0
cc_279 N_A1_M1004_g N_A_653_367#_c_655_n 0.00344413f $X=3.19 $Y=2.465 $X2=0
+ $Y2=0
cc_280 N_A1_c_290_p N_A_653_367#_c_656_n 0.0153678f $X=5.265 $Y=2.015 $X2=0
+ $Y2=0
cc_281 N_A1_M1013_g N_A_653_367#_c_657_n 0.0128039f $X=5.34 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A1_M1019_g N_A_653_367#_c_657_n 0.0145615f $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A1_c_290_p N_A_653_367#_c_657_n 0.0114798f $X=5.265 $Y=2.015 $X2=0
+ $Y2=0
cc_284 A1 N_A_653_367#_c_657_n 0.0130175f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_285 N_A1_c_273_n N_A_653_367#_c_657_n 4.409e-19 $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_286 A1 N_A_653_367#_c_662_n 0.0159237f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_287 N_A1_c_273_n N_A_653_367#_c_662_n 5.70006e-19 $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_288 N_A1_M1002_g N_VGND_c_689_n 0.012141f $X=3.205 $Y=0.665 $X2=0 $Y2=0
cc_289 N_A1_M1005_g N_VGND_c_692_n 0.0101171f $X=5.355 $Y=0.665 $X2=0 $Y2=0
cc_290 N_A1_M1020_g N_VGND_c_692_n 5.98801e-19 $X=5.785 $Y=0.665 $X2=0 $Y2=0
cc_291 N_A1_M1005_g N_VGND_c_693_n 6.04459e-19 $X=5.355 $Y=0.665 $X2=0 $Y2=0
cc_292 N_A1_M1020_g N_VGND_c_693_n 0.0103549f $X=5.785 $Y=0.665 $X2=0 $Y2=0
cc_293 N_A1_M1022_g N_VGND_c_693_n 0.0120479f $X=6.215 $Y=0.665 $X2=0 $Y2=0
cc_294 N_A1_M1002_g N_VGND_c_694_n 0.00477554f $X=3.205 $Y=0.665 $X2=0 $Y2=0
cc_295 N_A1_M1005_g N_VGND_c_699_n 0.00477554f $X=5.355 $Y=0.665 $X2=0 $Y2=0
cc_296 N_A1_M1020_g N_VGND_c_699_n 0.00477554f $X=5.785 $Y=0.665 $X2=0 $Y2=0
cc_297 N_A1_M1022_g N_VGND_c_700_n 0.00477554f $X=6.215 $Y=0.665 $X2=0 $Y2=0
cc_298 N_A1_M1002_g N_VGND_c_701_n 0.00841061f $X=3.205 $Y=0.665 $X2=0 $Y2=0
cc_299 N_A1_M1005_g N_VGND_c_701_n 0.00825815f $X=5.355 $Y=0.665 $X2=0 $Y2=0
cc_300 N_A1_M1020_g N_VGND_c_701_n 0.00825815f $X=5.785 $Y=0.665 $X2=0 $Y2=0
cc_301 N_A1_M1022_g N_VGND_c_701_n 0.00921794f $X=6.215 $Y=0.665 $X2=0 $Y2=0
cc_302 N_A1_M1002_g N_A_218_49#_c_787_n 0.013863f $X=3.205 $Y=0.665 $X2=0 $Y2=0
cc_303 N_A1_c_278_n N_A_218_49#_c_787_n 0.0169745f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_304 N_A1_c_270_n N_A_218_49#_c_787_n 0.00249084f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_305 N_A1_c_278_n N_A_218_49#_c_788_n 0.00622313f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_306 N_A1_c_270_n N_A_218_49#_c_788_n 0.0020436f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_307 N_A1_M1005_g N_A_218_49#_c_790_n 0.0142382f $X=5.355 $Y=0.665 $X2=0 $Y2=0
cc_308 A1 N_A_218_49#_c_790_n 0.0131256f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_309 A1 N_A_218_49#_c_790_n 0.00299172f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_310 N_A1_c_273_n N_A_218_49#_c_790_n 4.34971e-19 $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_311 N_A1_M1020_g N_A_218_49#_c_791_n 0.0136937f $X=5.785 $Y=0.665 $X2=0 $Y2=0
cc_312 N_A1_M1022_g N_A_218_49#_c_791_n 0.0146684f $X=6.215 $Y=0.665 $X2=0 $Y2=0
cc_313 A1 N_A_218_49#_c_791_n 0.0719173f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_314 N_A1_c_273_n N_A_218_49#_c_791_n 0.0103115f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_315 A1 N_A_218_49#_c_796_n 0.0161952f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_316 N_A1_c_273_n N_A_218_49#_c_796_n 0.00263213f $X=6.45 $Y=1.46 $X2=0 $Y2=0
cc_317 N_A2_M1025_g N_VPWR_c_472_n 0.00125629f $X=4.91 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A2_M1007_g N_VPWR_c_480_n 0.00357877f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A2_M1014_g N_VPWR_c_480_n 0.00357877f $X=4.05 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A2_M1017_g N_VPWR_c_480_n 0.00357877f $X=4.48 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A2_M1025_g N_VPWR_c_480_n 0.00357842f $X=4.91 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A2_M1007_g N_VPWR_c_467_n 0.00540833f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_323 N_A2_M1014_g N_VPWR_c_467_n 0.00538202f $X=4.05 $Y=2.465 $X2=0 $Y2=0
cc_324 N_A2_M1017_g N_VPWR_c_467_n 0.00538202f $X=4.48 $Y=2.465 $X2=0 $Y2=0
cc_325 N_A2_M1025_g N_VPWR_c_467_n 0.00537652f $X=4.91 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A2_M1007_g N_Y_c_592_n 0.00532185f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A2_M1007_g N_Y_c_618_n 0.00735603f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_328 N_A2_M1014_g N_Y_c_618_n 0.0127377f $X=4.05 $Y=2.465 $X2=0 $Y2=0
cc_329 N_A2_M1017_g N_Y_c_618_n 0.0128286f $X=4.48 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A2_M1007_g N_A_653_367#_c_655_n 0.0107823f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A2_M1014_g N_A_653_367#_c_655_n 0.0107823f $X=4.05 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A2_M1017_g N_A_653_367#_c_655_n 0.0107038f $X=4.48 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A2_M1025_g N_A_653_367#_c_655_n 0.0135746f $X=4.91 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_M1025_g N_A_653_367#_c_656_n 0.0023782f $X=4.91 $Y=2.465 $X2=0 $Y2=0
cc_335 N_A2_M1017_g N_A_653_367#_c_669_n 8.15857e-19 $X=4.48 $Y=2.465 $X2=0
+ $Y2=0
cc_336 N_A2_M1025_g N_A_653_367#_c_669_n 0.00695201f $X=4.91 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_A2_M1000_g N_VGND_c_689_n 0.0109917f $X=3.635 $Y=0.665 $X2=0 $Y2=0
cc_338 N_A2_M1010_g N_VGND_c_689_n 6.10117e-19 $X=4.065 $Y=0.665 $X2=0 $Y2=0
cc_339 N_A2_M1000_g N_VGND_c_690_n 6.10117e-19 $X=3.635 $Y=0.665 $X2=0 $Y2=0
cc_340 N_A2_M1010_g N_VGND_c_690_n 0.0107978f $X=4.065 $Y=0.665 $X2=0 $Y2=0
cc_341 N_A2_M1012_g N_VGND_c_690_n 0.0107978f $X=4.495 $Y=0.665 $X2=0 $Y2=0
cc_342 N_A2_M1016_g N_VGND_c_690_n 6.10117e-19 $X=4.925 $Y=0.665 $X2=0 $Y2=0
cc_343 N_A2_M1012_g N_VGND_c_691_n 0.00477554f $X=4.495 $Y=0.665 $X2=0 $Y2=0
cc_344 N_A2_M1016_g N_VGND_c_691_n 0.00477554f $X=4.925 $Y=0.665 $X2=0 $Y2=0
cc_345 N_A2_M1012_g N_VGND_c_692_n 5.98801e-19 $X=4.495 $Y=0.665 $X2=0 $Y2=0
cc_346 N_A2_M1016_g N_VGND_c_692_n 0.0101171f $X=4.925 $Y=0.665 $X2=0 $Y2=0
cc_347 N_A2_M1000_g N_VGND_c_696_n 0.00477554f $X=3.635 $Y=0.665 $X2=0 $Y2=0
cc_348 N_A2_M1010_g N_VGND_c_696_n 0.00477554f $X=4.065 $Y=0.665 $X2=0 $Y2=0
cc_349 N_A2_M1000_g N_VGND_c_701_n 0.00825815f $X=3.635 $Y=0.665 $X2=0 $Y2=0
cc_350 N_A2_M1010_g N_VGND_c_701_n 0.00825815f $X=4.065 $Y=0.665 $X2=0 $Y2=0
cc_351 N_A2_M1012_g N_VGND_c_701_n 0.00825815f $X=4.495 $Y=0.665 $X2=0 $Y2=0
cc_352 N_A2_M1016_g N_VGND_c_701_n 0.00825815f $X=4.925 $Y=0.665 $X2=0 $Y2=0
cc_353 N_A2_M1000_g N_A_218_49#_c_787_n 0.0140696f $X=3.635 $Y=0.665 $X2=0 $Y2=0
cc_354 N_A2_c_388_n N_A_218_49#_c_787_n 0.01553f $X=4.745 $Y=1.51 $X2=0 $Y2=0
cc_355 N_A2_M1010_g N_A_218_49#_c_789_n 0.0141109f $X=4.065 $Y=0.665 $X2=0 $Y2=0
cc_356 N_A2_M1012_g N_A_218_49#_c_789_n 0.0140617f $X=4.495 $Y=0.665 $X2=0 $Y2=0
cc_357 N_A2_c_388_n N_A_218_49#_c_789_n 0.0433075f $X=4.745 $Y=1.51 $X2=0 $Y2=0
cc_358 N_A2_c_389_n N_A_218_49#_c_789_n 0.00247942f $X=4.91 $Y=1.51 $X2=0 $Y2=0
cc_359 N_A2_M1016_g N_A_218_49#_c_790_n 0.0170939f $X=4.925 $Y=0.665 $X2=0 $Y2=0
cc_360 N_A2_c_388_n N_A_218_49#_c_790_n 0.00628848f $X=4.745 $Y=1.51 $X2=0 $Y2=0
cc_361 N_A2_c_388_n N_A_218_49#_c_794_n 0.0141697f $X=4.745 $Y=1.51 $X2=0 $Y2=0
cc_362 N_A2_c_389_n N_A_218_49#_c_794_n 0.00259169f $X=4.91 $Y=1.51 $X2=0 $Y2=0
cc_363 N_A2_M1016_g N_A_218_49#_c_795_n 6.32871e-19 $X=4.925 $Y=0.665 $X2=0
+ $Y2=0
cc_364 N_A2_c_388_n N_A_218_49#_c_795_n 0.0141186f $X=4.745 $Y=1.51 $X2=0 $Y2=0
cc_365 N_A2_c_389_n N_A_218_49#_c_795_n 0.00259169f $X=4.91 $Y=1.51 $X2=0 $Y2=0
cc_366 N_VPWR_c_467_n N_Y_M1001_s 0.00397496f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_367 N_VPWR_c_467_n N_Y_M1011_s 0.00405781f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_368 N_VPWR_c_467_n N_Y_M1007_d 0.00225186f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_369 N_VPWR_c_467_n N_Y_M1017_d 0.00225186f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_370 N_VPWR_c_475_n N_Y_c_625_n 0.0138717f $X=1.91 $Y=3.33 $X2=0 $Y2=0
cc_371 N_VPWR_c_467_n N_Y_c_625_n 0.00886411f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_372 N_VPWR_M1003_d N_Y_c_572_n 0.00180746f $X=1.935 $Y=1.835 $X2=0 $Y2=0
cc_373 N_VPWR_c_470_n N_Y_c_572_n 0.0163514f $X=2.075 $Y=2.19 $X2=0 $Y2=0
cc_374 N_VPWR_c_469_n N_Y_c_573_n 7.77868e-19 $X=1.215 $Y=1.99 $X2=0 $Y2=0
cc_375 N_VPWR_c_477_n N_Y_c_630_n 0.0124525f $X=2.77 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_c_467_n N_Y_c_630_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPWR_c_467_n N_Y_c_595_n 0.00439337f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_378 N_VPWR_M1021_d N_Y_c_596_n 0.00881925f $X=2.795 $Y=1.835 $X2=0 $Y2=0
cc_379 N_VPWR_c_471_n N_Y_c_596_n 0.0186172f $X=2.955 $Y=2.865 $X2=0 $Y2=0
cc_380 N_VPWR_c_467_n N_Y_c_596_n 0.00775347f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_467_n N_A_653_367#_M1004_d 0.00223577f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_382 N_VPWR_c_467_n N_A_653_367#_M1014_s 0.00223577f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_467_n N_A_653_367#_M1025_s 0.00376624f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_467_n N_A_653_367#_M1019_d 0.00536646f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_480_n N_A_653_367#_c_655_n 0.0977356f $X=5.39 $Y=3.33 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_467_n N_A_653_367#_c_655_n 0.0623809f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_480_n N_A_653_367#_c_669_n 0.0157917f $X=5.39 $Y=3.33 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_467_n N_A_653_367#_c_669_n 0.00992063f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_389 N_VPWR_M1013_s N_A_653_367#_c_657_n 0.00460332f $X=5.415 $Y=1.835 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_472_n N_A_653_367#_c_657_n 0.0172078f $X=5.555 $Y=2.765 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_481_n N_A_653_367#_c_681_n 0.0124525f $X=6.25 $Y=3.33 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_467_n N_A_653_367#_c_681_n 0.00730901f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_393 N_Y_c_592_n N_A_653_367#_M1004_d 0.00362676f $X=3.57 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_394 N_Y_c_618_n N_A_653_367#_M1014_s 0.00355423f $X=4.695 $Y=2.445 $X2=0
+ $Y2=0
cc_395 N_Y_M1007_d N_A_653_367#_c_655_n 0.00342473f $X=3.695 $Y=1.835 $X2=0
+ $Y2=0
cc_396 N_Y_M1017_d N_A_653_367#_c_655_n 0.00342473f $X=4.555 $Y=1.835 $X2=0
+ $Y2=0
cc_397 N_Y_c_592_n N_A_653_367#_c_655_n 0.0801005f $X=3.57 $Y=2.445 $X2=0 $Y2=0
cc_398 N_Y_M1006_s N_VGND_c_701_n 0.00225186f $X=1.505 $Y=0.245 $X2=0 $Y2=0
cc_399 N_Y_M1015_s N_VGND_c_701_n 0.00225186f $X=2.365 $Y=0.245 $X2=0 $Y2=0
cc_400 N_Y_c_571_n N_A_218_49#_M1008_d 0.00182459f $X=2.335 $Y=0.98 $X2=0 $Y2=0
cc_401 N_Y_M1006_s N_A_218_49#_c_798_n 0.00344337f $X=1.505 $Y=0.245 $X2=0 $Y2=0
cc_402 N_Y_M1015_s N_A_218_49#_c_798_n 0.00343901f $X=2.365 $Y=0.245 $X2=0 $Y2=0
cc_403 N_Y_c_582_n N_A_218_49#_c_798_n 0.0210584f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_404 N_Y_c_571_n N_A_218_49#_c_798_n 0.0438722f $X=2.335 $Y=0.98 $X2=0 $Y2=0
cc_405 N_Y_c_582_n N_A_218_49#_c_802_n 0.0221423f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_406 N_Y_c_582_n N_A_218_49#_c_788_n 0.0115367f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_407 N_Y_c_584_n N_A_218_49#_c_788_n 0.00337337f $X=2.53 $Y=1.755 $X2=0 $Y2=0
cc_408 N_VGND_c_701_n N_A_218_49#_M1006_d 0.00212301f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_409 N_VGND_c_701_n N_A_218_49#_M1008_d 0.00223577f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_701_n N_A_218_49#_M1018_d 0.0042086f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_701_n N_A_218_49#_M1000_d 0.00536646f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_701_n N_A_218_49#_M1012_d 0.00536646f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_701_n N_A_218_49#_M1005_s 0.00536646f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_701_n N_A_218_49#_M1022_s 0.00368844f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_694_n N_A_218_49#_c_798_n 0.0869388f $X=3.255 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_701_n N_A_218_49#_c_798_n 0.0550006f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_694_n N_A_218_49#_c_854_n 0.0129414f $X=3.255 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_701_n N_A_218_49#_c_854_n 0.00738676f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_M1002_d N_A_218_49#_c_787_n 0.00176461f $X=3.28 $Y=0.245 $X2=0
+ $Y2=0
cc_420 N_VGND_c_689_n N_A_218_49#_c_787_n 0.0170777f $X=3.42 $Y=0.37 $X2=0 $Y2=0
cc_421 N_VGND_c_696_n N_A_218_49#_c_858_n 0.0124525f $X=4.115 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_701_n N_A_218_49#_c_858_n 0.00730901f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_M1010_s N_A_218_49#_c_789_n 0.00176461f $X=4.14 $Y=0.245 $X2=0
+ $Y2=0
cc_424 N_VGND_c_690_n N_A_218_49#_c_789_n 0.0170777f $X=4.28 $Y=0.39 $X2=0 $Y2=0
cc_425 N_VGND_c_691_n N_A_218_49#_c_862_n 0.0124525f $X=4.975 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_701_n N_A_218_49#_c_862_n 0.00730901f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_M1016_s N_A_218_49#_c_790_n 0.00177068f $X=5 $Y=0.245 $X2=0 $Y2=0
cc_428 N_VGND_c_692_n N_A_218_49#_c_790_n 0.0172078f $X=5.14 $Y=0.39 $X2=0 $Y2=0
cc_429 N_VGND_c_699_n N_A_218_49#_c_866_n 0.0124525f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_701_n N_A_218_49#_c_866_n 0.00730901f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_M1020_d N_A_218_49#_c_791_n 0.00176461f $X=5.86 $Y=0.245 $X2=0
+ $Y2=0
cc_432 N_VGND_c_693_n N_A_218_49#_c_791_n 0.0170777f $X=6 $Y=0.39 $X2=0 $Y2=0
cc_433 N_VGND_c_700_n N_A_218_49#_c_792_n 0.0178111f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_701_n N_A_218_49#_c_792_n 0.0100304f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_688_n N_A_218_49#_c_793_n 0.0506995f $X=0.69 $Y=0.39 $X2=0 $Y2=0
cc_436 N_VGND_c_694_n N_A_218_49#_c_793_n 0.021207f $X=3.255 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_701_n N_A_218_49#_c_793_n 0.012647f $X=6.48 $Y=0 $X2=0 $Y2=0
