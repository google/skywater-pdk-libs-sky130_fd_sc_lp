* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_0 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_1075_493# S1 a_294_506# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_31_506# S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_442_119# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1029_37# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND A1 a_642_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_685_504# S0 a_793_504# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_793_504# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_685_504# S1 a_1075_493# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_685_504# a_1029_37# a_1075_493# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR A1 a_613_504# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_613_504# a_31_506# a_685_504# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_31_506# S0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1075_493# a_1029_37# a_294_506# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_642_119# S0 a_685_504# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1029_37# S1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_270_119# a_31_506# a_294_506# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_800_119# A0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_1075_493# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VGND A2 a_270_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_294_506# S0 a_442_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR A2 a_222_506# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_222_506# S0 a_294_506# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_685_504# a_31_506# a_800_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_1075_493# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_294_506# a_31_506# a_426_504# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_426_504# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
