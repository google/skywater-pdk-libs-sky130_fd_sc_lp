# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__dfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 1.180000 2.080000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.475000 0.265000 13.830000 1.125000 ;
        RECT 13.475000 1.815000 13.830000 3.065000 ;
        RECT 13.660000 1.125000 13.830000 1.815000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.585900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.975000 0.265000 12.435000 1.005000 ;
        RECT 12.075000 1.695000 12.435000 2.995000 ;
        RECT 12.265000 1.005000 12.435000 1.695000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.165000 1.180000 11.520000 1.515000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.895000 1.550000 5.185000 1.595000 ;
        RECT 4.895000 1.595000 9.025000 1.735000 ;
        RECT 4.895000 1.735000 5.185000 1.780000 ;
        RECT 8.735000 1.550000 9.025000 1.595000 ;
        RECT 8.735000 1.735000 9.025000 1.780000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.955000 0.445000 2.150000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 13.920000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 14.110000 3.520000 ;
        RECT 10.910000 1.535000 12.475000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.110000  0.085000  0.360000 0.775000 ;
      RECT  0.115000  2.385000  0.445000 3.245000 ;
      RECT  0.540000  0.315000  0.870000 0.775000 ;
      RECT  0.625000  0.775000  0.870000 1.195000 ;
      RECT  0.625000  1.195000  1.065000 1.865000 ;
      RECT  0.625000  1.865000  0.955000 3.065000 ;
      RECT  1.085000  0.575000  1.415000 1.015000 ;
      RECT  1.205000  2.045000  1.535000 2.905000 ;
      RECT  1.245000  1.015000  1.415000 1.875000 ;
      RECT  1.245000  1.875000  2.550000 2.045000 ;
      RECT  1.595000  0.085000  1.925000 1.000000 ;
      RECT  1.715000  2.225000  2.045000 3.245000 ;
      RECT  2.275000  2.305000  2.900000 2.475000 ;
      RECT  2.275000  2.475000  2.605000 2.685000 ;
      RECT  2.290000  1.480000  2.550000 1.875000 ;
      RECT  2.410000  0.575000  2.740000 1.130000 ;
      RECT  2.410000  1.130000  2.900000 1.300000 ;
      RECT  2.730000  1.300000  2.900000 2.305000 ;
      RECT  2.920000  0.530000  3.250000 0.950000 ;
      RECT  3.080000  0.950000  3.250000 2.225000 ;
      RECT  3.080000  2.225000  3.970000 2.395000 ;
      RECT  3.080000  2.395000  3.410000 2.685000 ;
      RECT  3.430000  1.055000  4.860000 1.225000 ;
      RECT  3.430000  1.225000  3.620000 1.750000 ;
      RECT  3.800000  1.405000  4.695000 1.575000 ;
      RECT  3.800000  1.575000  3.970000 2.225000 ;
      RECT  4.150000  1.755000  4.345000 2.310000 ;
      RECT  4.150000  2.310000  6.015000 2.480000 ;
      RECT  4.180000  0.085000  4.510000 0.875000 ;
      RECT  4.525000  1.575000  4.695000 1.960000 ;
      RECT  4.525000  1.960000  5.505000 2.130000 ;
      RECT  4.605000  2.660000  4.935000 3.245000 ;
      RECT  4.690000  0.265000  6.655000 0.435000 ;
      RECT  4.690000  0.435000  4.860000 1.055000 ;
      RECT  4.875000  1.405000  5.155000 1.780000 ;
      RECT  5.040000  0.615000  6.305000 0.785000 ;
      RECT  5.040000  0.785000  5.370000 0.990000 ;
      RECT  5.335000  1.475000  5.955000 1.735000 ;
      RECT  5.335000  1.735000  5.505000 1.960000 ;
      RECT  5.550000  0.965000  5.880000 1.125000 ;
      RECT  5.550000  1.125000  6.305000 1.295000 ;
      RECT  5.685000  1.915000  6.545000 2.085000 ;
      RECT  5.685000  2.085000  6.015000 2.310000 ;
      RECT  5.685000  2.480000  6.015000 2.755000 ;
      RECT  6.135000  0.785000  6.305000 0.945000 ;
      RECT  6.135000  1.295000  6.305000 1.435000 ;
      RECT  6.135000  1.435000  7.180000 1.695000 ;
      RECT  6.375000  1.695000  6.545000 1.915000 ;
      RECT  6.485000  0.435000  6.655000 1.085000 ;
      RECT  6.485000  1.085000  7.530000 1.255000 ;
      RECT  6.725000  1.875000  7.055000 3.245000 ;
      RECT  6.835000  0.085000  7.085000 0.905000 ;
      RECT  7.360000  1.255000  7.530000 1.345000 ;
      RECT  7.360000  1.345000  7.750000 1.675000 ;
      RECT  7.360000  1.675000  7.530000 2.895000 ;
      RECT  7.360000  2.895000  8.615000 3.065000 ;
      RECT  7.710000  2.120000  8.100000 2.715000 ;
      RECT  7.930000  0.575000  8.260000 1.150000 ;
      RECT  7.930000  1.150000  9.945000 1.320000 ;
      RECT  7.930000  1.320000  8.100000 2.120000 ;
      RECT  8.320000  1.730000  8.615000 2.895000 ;
      RECT  8.795000  1.500000  9.580000 1.830000 ;
      RECT  8.860000  2.070000 10.055000 2.205000 ;
      RECT  8.860000  2.205000 11.895000 2.375000 ;
      RECT  8.860000  2.375000 10.055000 2.400000 ;
      RECT  8.945000  0.085000  9.275000 0.970000 ;
      RECT  9.215000  2.580000  9.545000 3.245000 ;
      RECT  9.455000  0.265000 10.805000 0.435000 ;
      RECT  9.455000  0.435000  9.785000 0.970000 ;
      RECT  9.725000  2.400000 10.055000 3.065000 ;
      RECT  9.775000  1.320000  9.945000 1.460000 ;
      RECT  9.775000  1.460000 10.120000 1.790000 ;
      RECT  9.965000  0.615000 10.295000 0.830000 ;
      RECT  9.965000  0.830000 10.470000 0.970000 ;
      RECT 10.125000  0.970000 10.470000 1.000000 ;
      RECT 10.300000  1.000000 10.470000 2.205000 ;
      RECT 10.475000  0.435000 10.805000 0.650000 ;
      RECT 10.515000  2.555000 10.845000 3.245000 ;
      RECT 10.650000  0.830000 11.365000 1.000000 ;
      RECT 10.650000  1.000000 10.980000 1.695000 ;
      RECT 10.650000  1.695000 11.390000 2.025000 ;
      RECT 11.035000  0.635000 11.365000 0.830000 ;
      RECT 11.545000  0.085000 11.795000 1.000000 ;
      RECT 11.565000  2.555000 11.895000 3.245000 ;
      RECT 11.725000  1.185000 12.085000 1.515000 ;
      RECT 11.725000  1.515000 11.895000 2.205000 ;
      RECT 12.615000  0.665000 12.865000 1.305000 ;
      RECT 12.615000  1.305000 13.480000 1.635000 ;
      RECT 12.615000  1.635000 12.865000 2.495000 ;
      RECT 13.045000  0.085000 13.295000 1.125000 ;
      RECT 13.045000  1.815000 13.295000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.580000  5.125000 1.750000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.580000  8.965000 1.750000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_lp__dfbbn_1
END LIBRARY
