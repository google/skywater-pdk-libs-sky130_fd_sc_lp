* File: sky130_fd_sc_lp__and4b_1.pex.spice
* Created: Wed Sep  2 09:33:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4B_1%A_N 3 7 12 13 14 17 18
c33 18 0 6.35615e-20 $X=0.385 $Y=1.09
r34 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.09 $X2=0.385 $Y2=1.09
r35 14 18 3.40061 $w=5.08e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.26
+ $X2=0.385 $Y2=1.26
r36 12 17 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.385 $Y=1.445
+ $X2=0.385 $Y2=1.09
r37 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.412 $Y=1.445
+ $X2=0.412 $Y2=1.595
r38 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=0.925
+ $X2=0.385 $Y2=1.09
r39 7 13 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.53 $Y=2.045
+ $X2=0.53 $Y2=1.595
r40 3 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.475 $Y=0.455 $X2=0.475
+ $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%A_27_49# 1 2 9 11 12 13 15 18 21 25 27 28 29
+ 30 34 35 37 38
c81 34 0 1.26847e-19 $X=0.98 $Y=0.94
c82 29 0 1.24023e-19 $X=0.76 $Y=1.78
c83 9 0 6.35615e-20 $X=1 $Y=2.045
r84 37 38 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.845 $Y=1.695
+ $X2=0.845 $Y2=1.445
r85 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.98
+ $Y=0.94 $X2=0.98 $Y2=0.94
r86 32 38 7.98337 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=0.912 $Y=1.293
+ $X2=0.912 $Y2=1.445
r87 32 34 13.3381 $w=3.03e-07 $l=3.53e-07 $layer=LI1_cond $X=0.912 $Y=1.293
+ $X2=0.912 $Y2=0.94
r88 31 34 4.34528 $w=3.03e-07 $l=1.15e-07 $layer=LI1_cond $X=0.912 $Y=0.825
+ $X2=0.912 $Y2=0.94
r89 29 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=1.78
+ $X2=0.845 $Y2=1.695
r90 29 30 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.76 $Y=1.78
+ $X2=0.43 $Y2=1.78
r91 27 31 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=0.76 $Y=0.74
+ $X2=0.912 $Y2=0.825
r92 27 28 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.76 $Y=0.74
+ $X2=0.355 $Y2=0.74
r93 23 30 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.29 $Y=1.865
+ $X2=0.43 $Y2=1.78
r94 23 25 7.40856 $w=2.78e-07 $l=1.8e-07 $layer=LI1_cond $X=0.29 $Y=1.865
+ $X2=0.29 $Y2=2.045
r95 19 28 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=0.655
+ $X2=0.355 $Y2=0.74
r96 19 21 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=0.225 $Y=0.655
+ $X2=0.225 $Y2=0.455
r97 17 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.98 $Y=1.28
+ $X2=0.98 $Y2=0.94
r98 17 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.28
+ $X2=0.98 $Y2=1.445
r99 16 35 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.98 $Y=0.925
+ $X2=0.98 $Y2=0.94
r100 13 15 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.425 $Y=0.775
+ $X2=1.425 $Y2=0.445
r101 12 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.145 $Y=0.85
+ $X2=0.98 $Y2=0.925
r102 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.35 $Y=0.85
+ $X2=1.425 $Y2=0.775
r103 11 12 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=1.35 $Y=0.85
+ $X2=1.145 $Y2=0.85
r104 9 18 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1 $Y=2.045 $X2=1
+ $Y2=1.445
r105 2 25 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.835 $X2=0.315 $Y2=2.045
r106 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%B 3 7 9 10 18
c37 7 0 1.26847e-19 $X=1.785 $Y=0.445
c38 3 0 1.24023e-19 $X=1.43 $Y=2.045
r39 16 18 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.68 $Y=1.375
+ $X2=1.785 $Y2=1.375
r40 13 16 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.43 $Y=1.375
+ $X2=1.68 $Y2=1.375
r41 9 10 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.295
+ $X2=1.717 $Y2=1.665
r42 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.375 $X2=1.68 $Y2=1.375
r43 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.21
+ $X2=1.785 $Y2=1.375
r44 5 7 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.785 $Y=1.21
+ $X2=1.785 $Y2=0.445
r45 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.54
+ $X2=1.43 $Y2=1.375
r46 1 3 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.43 $Y=1.54 $X2=1.43
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%C 3 7 9 10 15
r37 15 17 20.271 $w=3.21e-07 $l=1.35e-07 $layer=POLY_cond $X=2.235 $Y=1.517
+ $X2=2.37 $Y2=1.517
r38 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.51 $X2=2.235 $Y2=1.51
r39 13 15 13.514 $w=3.21e-07 $l=9e-08 $layer=POLY_cond $X=2.145 $Y=1.517
+ $X2=2.235 $Y2=1.517
r40 10 16 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.175 $Y=1.665
+ $X2=2.175 $Y2=1.51
r41 9 16 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.175 $Y=1.295
+ $X2=2.175 $Y2=1.51
r42 5 17 20.5661 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=2.37 $Y=1.69
+ $X2=2.37 $Y2=1.517
r43 5 7 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=2.37 $Y=1.69 $X2=2.37
+ $Y2=2.045
r44 1 13 20.5661 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.145 $Y=1.345
+ $X2=2.145 $Y2=1.517
r45 1 3 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.145 $Y=1.345 $X2=2.145
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%D 1 3 8 11 12 19
c43 8 0 1.82261e-19 $X=2.8 $Y=2.045
r44 16 19 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.64 $Y=2.79 $X2=2.8
+ $Y2=2.79
r45 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=2.79 $X2=2.64 $Y2=2.79
r46 11 12 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.632 $Y=2.405
+ $X2=2.632 $Y2=2.775
r47 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=2.625 $X2=2.8
+ $Y2=2.79
r48 6 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.8 $Y=2.625 $X2=2.8
+ $Y2=2.045
r49 5 8 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.8 $Y=1.3 $X2=2.8
+ $Y2=2.045
r50 1 5 66.1349 $w=2.15e-07 $l=4.69894e-07 $layer=POLY_cond $X=2.505 $Y=0.955
+ $X2=2.8 $Y2=1.3
r51 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.505 $Y=0.955
+ $X2=2.505 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%A_215_367# 1 2 3 12 15 17 18 20 21 24 27 31
+ 32 42 44 45 47
r100 40 42 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.215 $Y=1.96
+ $X2=1.32 $Y2=1.96
r101 32 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.35
+ $X2=3.25 $Y2=1.515
r102 32 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.35
+ $X2=3.25 $Y2=1.185
r103 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.35 $X2=3.25 $Y2=1.35
r104 29 45 0.221902 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=2.73 $Y=1.35
+ $X2=2.61 $Y2=1.35
r105 29 31 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=2.73 $Y=1.35
+ $X2=3.25 $Y2=1.35
r106 25 45 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.515
+ $X2=2.61 $Y2=1.35
r107 25 27 21.3682 $w=2.38e-07 $l=4.45e-07 $layer=LI1_cond $X=2.61 $Y=1.515
+ $X2=2.61 $Y2=1.96
r108 24 45 7.38875 $w=2.1e-07 $l=1.79374e-07 $layer=LI1_cond $X=2.58 $Y=1.185
+ $X2=2.61 $Y2=1.35
r109 23 24 9.5505 $w=1.78e-07 $l=1.55e-07 $layer=LI1_cond $X=2.58 $Y=1.03
+ $X2=2.58 $Y2=1.185
r110 22 44 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.515 $Y=0.945
+ $X2=1.375 $Y2=0.945
r111 21 23 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.49 $Y=0.945
+ $X2=2.58 $Y2=1.03
r112 21 22 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=2.49 $Y=0.945
+ $X2=1.515 $Y2=0.945
r113 20 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=1.795
+ $X2=1.32 $Y2=1.96
r114 19 44 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=1.32 $Y=1.03
+ $X2=1.375 $Y2=0.945
r115 19 20 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.32 $Y=1.03
+ $X2=1.32 $Y2=1.795
r116 18 44 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0.86
+ $X2=1.375 $Y2=0.945
r117 17 35 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.37
+ $X2=1.21 $Y2=0.37
r118 17 18 15.4345 $w=2.78e-07 $l=3.75e-07 $layer=LI1_cond $X=1.375 $Y=0.485
+ $X2=1.375 $Y2=0.86
r119 15 48 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.325 $Y=2.465
+ $X2=3.325 $Y2=1.515
r120 12 47 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.31 $Y=0.655
+ $X2=3.31 $Y2=1.185
r121 3 27 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.835 $X2=2.585 $Y2=1.96
r122 2 40 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.835 $X2=1.215 $Y2=1.96
r123 1 35 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.21 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%VPWR 1 2 3 12 16 21 23 26 28 33 38 45 46 49
+ 52 55
c46 23 0 1.82261e-19 $X=3.065 $Y=1.98
r47 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 46 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 43 55 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.105 $Y2=3.33
r53 43 45 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 39 52 14.0152 $w=1.7e-07 $l=3.68e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=1.952 $Y2=3.33
r58 39 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=3.33 $X2=2.64
+ $Y2=3.33
r59 38 55 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.105 $Y2=3.33
r60 38 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r63 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=3.33
+ $X2=0.765 $Y2=3.33
r64 34 36 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=3.33 $X2=1.2
+ $Y2=3.33
r65 33 52 14.0152 $w=1.7e-07 $l=3.67e-07 $layer=LI1_cond $X=1.585 $Y=3.33
+ $X2=1.952 $Y2=3.33
r66 33 36 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.585 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 31 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 28 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.765 $Y2=3.33
r70 28 30 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33 $X2=0.24
+ $Y2=3.33
r71 26 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 26 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 23 25 4.78309 $w=3.63e-07 $l=1.45e-07 $layer=LI1_cond $X=3.082 $Y=1.98
+ $X2=3.082 $Y2=2.125
r74 21 25 11.7045 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=3.105 $Y=2.45
+ $X2=3.105 $Y2=2.125
r75 19 55 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=3.245
+ $X2=3.105 $Y2=3.33
r76 19 21 28.631 $w=3.18e-07 $l=7.95e-07 $layer=LI1_cond $X=3.105 $Y=3.245
+ $X2=3.105 $Y2=2.45
r77 14 52 2.96355 $w=7.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.952 $Y=3.245
+ $X2=1.952 $Y2=3.33
r78 14 16 19.5278 $w=7.33e-07 $l=1.2e-06 $layer=LI1_cond $X=1.952 $Y=3.245
+ $X2=1.952 $Y2=2.045
r79 10 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=3.245
+ $X2=0.765 $Y2=3.33
r80 10 12 39.2878 $w=3.28e-07 $l=1.125e-06 $layer=LI1_cond $X=0.765 $Y=3.245
+ $X2=0.765 $Y2=2.12
r81 3 23 600 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.835 $X2=3.065 $Y2=1.98
r82 3 21 300 $w=1.7e-07 $l=7.23015e-07 $layer=licon1_PDIFF $count=2 $X=2.875
+ $Y=1.835 $X2=3.11 $Y2=2.45
r83 2 16 300 $w=1.7e-07 $l=7.47663e-07 $layer=licon1_PDIFF $count=2 $X=1.505
+ $Y=1.835 $X2=2.155 $Y2=2.045
r84 1 12 600 $w=1.7e-07 $l=3.56125e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.835 $X2=0.765 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%X 1 2 7 8 9 10 11 12 13 24 37
r20 34 37 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=3.595 $Y=1.975
+ $X2=3.595 $Y2=1.98
r21 13 44 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=3.595 $Y=2.775
+ $X2=3.595 $Y2=2.91
r22 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.595 $Y=2.405
+ $X2=3.595 $Y2=2.775
r23 11 34 0.46818 $w=3.18e-07 $l=1.3e-08 $layer=LI1_cond $X=3.595 $Y=1.962
+ $X2=3.595 $Y2=1.975
r24 11 50 5.87672 $w=3.18e-07 $l=1.47e-07 $layer=LI1_cond $X=3.595 $Y=1.962
+ $X2=3.595 $Y2=1.815
r25 11 12 12.893 $w=3.18e-07 $l=3.58e-07 $layer=LI1_cond $X=3.595 $Y=2.047
+ $X2=3.595 $Y2=2.405
r26 11 37 2.41293 $w=3.18e-07 $l=6.7e-08 $layer=LI1_cond $X=3.595 $Y=2.047
+ $X2=3.595 $Y2=1.98
r27 10 50 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=3.63 $Y=1.665
+ $X2=3.63 $Y2=1.815
r28 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.63 $Y=1.295
+ $X2=3.63 $Y2=1.665
r29 9 48 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.63 $Y=1.295
+ $X2=3.63 $Y2=1.015
r30 8 48 4.172 $w=3.93e-07 $l=9e-08 $layer=LI1_cond $X=3.557 $Y=0.925 $X2=3.557
+ $Y2=1.015
r31 8 22 3.12181 $w=3.93e-07 $l=1.07e-07 $layer=LI1_cond $X=3.557 $Y=0.925
+ $X2=3.557 $Y2=0.818
r32 7 22 7.67323 $w=3.93e-07 $l=2.63e-07 $layer=LI1_cond $X=3.557 $Y=0.555
+ $X2=3.557 $Y2=0.818
r33 7 24 4.37637 $w=3.93e-07 $l=1.5e-07 $layer=LI1_cond $X=3.557 $Y=0.555
+ $X2=3.557 $Y2=0.405
r34 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.835 $X2=3.54 $Y2=2.91
r35 2 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.835 $X2=3.54 $Y2=1.98
r36 1 24 91 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.235 $X2=3.525 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_1%VGND 1 2 9 13 15 17 22 32 33 36
r52 43 44 8.62314 $w=6.33e-07 $l=2.3e-07 $layer=LI1_cond $X=2.872 $Y=0.38
+ $X2=2.872 $Y2=0.61
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 33 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r55 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 30 32 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.6
+ $Y2=0
r57 29 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r58 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r59 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r60 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r61 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r62 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r63 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r64 22 43 7.15763 $w=6.33e-07 $l=3.8e-07 $layer=LI1_cond $X=2.872 $Y=0 $X2=2.872
+ $Y2=0.38
r65 22 30 8.68381 $w=1.7e-07 $l=3.18e-07 $layer=LI1_cond $X=2.872 $Y=0 $X2=3.19
+ $Y2=0
r66 22 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r67 22 28 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=0 $X2=2.16
+ $Y2=0
r68 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r69 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r70 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r71 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r72 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r73 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r74 13 44 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=3.06 $Y=0.85
+ $X2=3.06 $Y2=0.61
r75 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r76 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.4
r77 2 43 91 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_NDIFF $count=2 $X=2.58
+ $Y=0.235 $X2=3.095 $Y2=0.38
r78 2 13 182 $w=1.7e-07 $l=8.33637e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.235 $X2=3.095 $Y2=0.85
r79 1 9 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.245 $X2=0.69 $Y2=0.4
.ends

