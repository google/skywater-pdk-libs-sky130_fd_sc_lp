* NGSPICE file created from sky130_fd_sc_lp__o21a_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VGND A2 a_300_51# VNB nshort w=840000u l=150000u
+  ad=5.418e+11p pd=4.65e+06u as=4.578e+11p ps=4.45e+06u
M1001 a_420_367# A2 a_80_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=4.914e+11p ps=3.3e+06u
M1002 VPWR a_80_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1781e+12p pd=6.91e+06u as=3.339e+11p ps=3.05e+06u
M1003 VGND a_80_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1004 VPWR A1 a_420_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_300_51# B1 a_80_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1006 a_300_51# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_80_21# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

