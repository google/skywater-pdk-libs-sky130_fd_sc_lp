* File: sky130_fd_sc_lp__nand4bb_m.spice
* Created: Wed Sep  2 10:07:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4bb_m.pex.spice"
.subckt sky130_fd_sc_lp__nand4bb_m  VNB VPB B_N D C A_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A_N	A_N
* C	C
* D	D
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B_N_M1005_g N_A_27_151#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.11235 AS=0.1113 PD=0.955 PS=1.37 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1000 A_247_151# N_D_M1000_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.11235 PD=0.63 PS=0.955 NRD=14.28 NRS=49.992 M=1 R=2.8 SA=75000.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1011 A_319_151# N_C_M1011_g A_247_151# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75001.2 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1006 A_427_151# N_A_27_151#_M1006_g A_319_151# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_469_125#_M1001_g A_427_151# VNB NSHORT L=0.15 W=0.42
+ AD=0.1425 AS=0.0441 PD=1.64 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_469_125#_M1007_d N_A_N_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B_N_M1003_g N_A_27_151#_M1003_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1037 AS=0.1113 PD=0.93 PS=1.37 NRD=44.5417 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_D_M1009_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1037 PD=0.7 PS=0.93 NRD=0 NRS=44.5417 M=1 R=2.8 SA=75000.8
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_C_M1002_g N_Y_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.2 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1010 N_Y_M1010_d N_A_27_151#_M1010_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=18.7544 M=1 R=2.8 SA=75001.7
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_469_125#_M1004_g N_Y_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.10815 AS=0.0588 PD=0.935 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1008 N_A_469_125#_M1008_d N_A_N_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.10815 PD=1.37 PS=0.935 NRD=0 NRS=110.222 M=1 R=2.8
+ SA=75002.8 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__nand4bb_m.pxi.spice"
*
.ends
*
*
