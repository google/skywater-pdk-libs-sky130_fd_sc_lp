* File: sky130_fd_sc_lp__a2111oi_0.pxi.spice
* Created: Fri Aug 28 09:46:26 2020
* 
x_PM_SKY130_FD_SC_LP__A2111OI_0%D1 N_D1_c_79_n N_D1_c_80_n N_D1_c_81_n
+ N_D1_c_87_n N_D1_c_88_n N_D1_M1002_g N_D1_c_89_n N_D1_M1003_g N_D1_c_83_n D1
+ D1 D1 D1 N_D1_c_85_n PM_SKY130_FD_SC_LP__A2111OI_0%D1
x_PM_SKY130_FD_SC_LP__A2111OI_0%C1 N_C1_M1008_g N_C1_M1004_g N_C1_c_119_n
+ N_C1_c_124_n C1 C1 C1 C1 C1 N_C1_c_121_n PM_SKY130_FD_SC_LP__A2111OI_0%C1
x_PM_SKY130_FD_SC_LP__A2111OI_0%B1 N_B1_c_162_n N_B1_M1009_g N_B1_M1006_g
+ N_B1_c_168_n B1 B1 N_B1_c_165_n PM_SKY130_FD_SC_LP__A2111OI_0%B1
x_PM_SKY130_FD_SC_LP__A2111OI_0%A1 N_A1_M1005_g N_A1_M1000_g N_A1_c_208_n A1 A1
+ A1 N_A1_c_206_n PM_SKY130_FD_SC_LP__A2111OI_0%A1
x_PM_SKY130_FD_SC_LP__A2111OI_0%A2 N_A2_M1007_g N_A2_M1001_g N_A2_c_253_n
+ N_A2_c_254_n N_A2_c_260_n N_A2_c_261_n N_A2_c_255_n N_A2_c_256_n A2 A2 A2 A2
+ N_A2_c_258_n PM_SKY130_FD_SC_LP__A2111OI_0%A2
x_PM_SKY130_FD_SC_LP__A2111OI_0%Y N_Y_M1002_d N_Y_M1006_d N_Y_M1003_s
+ N_Y_c_302_n N_Y_c_303_n N_Y_c_297_n N_Y_c_298_n Y Y Y N_Y_c_299_n N_Y_c_300_n
+ Y N_Y_c_301_n PM_SKY130_FD_SC_LP__A2111OI_0%Y
x_PM_SKY130_FD_SC_LP__A2111OI_0%A_318_483# N_A_318_483#_M1009_d
+ N_A_318_483#_M1001_d N_A_318_483#_c_349_n N_A_318_483#_c_350_n
+ N_A_318_483#_c_351_n N_A_318_483#_c_352_n N_A_318_483#_c_353_n
+ N_A_318_483#_c_354_n PM_SKY130_FD_SC_LP__A2111OI_0%A_318_483#
x_PM_SKY130_FD_SC_LP__A2111OI_0%VPWR N_VPWR_M1005_d N_VPWR_c_385_n VPWR
+ N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_384_n N_VPWR_c_389_n
+ PM_SKY130_FD_SC_LP__A2111OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A2111OI_0%VGND N_VGND_M1002_s N_VGND_M1008_d
+ N_VGND_M1007_d N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n
+ N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n VGND N_VGND_c_421_n
+ N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n
+ PM_SKY130_FD_SC_LP__A2111OI_0%VGND
cc_1 VNB N_D1_c_79_n 0.00995287f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.14
cc_2 VNB N_D1_c_80_n 0.0255083f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.915
cc_3 VNB N_D1_c_81_n 0.0188553f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.915
cc_4 VNB N_D1_M1002_g 0.0270121f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_5 VNB N_D1_c_83_n 0.0197835f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_6 VNB D1 0.0375221f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_D1_c_85_n 0.0297019f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_8 VNB N_C1_M1008_g 0.0425445f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.915
cc_9 VNB N_C1_c_119_n 0.0182697f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.29
cc_10 VNB C1 0.00513598f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.735
cc_11 VNB N_C1_c_121_n 0.0166213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_162_n 0.0184472f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.14
cc_13 VNB N_B1_M1006_g 0.0386234f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_14 VNB B1 0.00305761f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_15 VNB N_B1_c_165_n 0.0171375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1000_g 0.0365295f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.84
cc_17 VNB A1 0.0102933f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_18 VNB N_A1_c_206_n 0.0548377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_M1007_g 0.0240704f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.915
cc_20 VNB N_A2_c_253_n 0.0541411f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.445
cc_21 VNB N_A2_c_254_n 0.00711081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_255_n 0.0089214f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_23 VNB N_A2_c_256_n 0.0185685f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_24 VNB A2 0.030873f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB N_A2_c_258_n 0.0301182f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_26 VNB N_Y_c_297_n 0.00285767f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_Y_c_298_n 0.0123837f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_28 VNB N_Y_c_299_n 0.00970304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_300_n 0.0116464f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.295
cc_30 VNB N_Y_c_301_n 0.00746138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_384_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_414_n 0.0192699f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.735
cc_33 VNB N_VGND_c_415_n 0.00497133f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_34 VNB N_VGND_c_416_n 0.0175746f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_35 VNB N_VGND_c_417_n 0.0131219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_418_n 0.00564902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_419_n 0.0165526f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_38 VNB N_VGND_c_420_n 0.00622613f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_39 VNB N_VGND_c_421_n 0.0239127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_422_n 0.0191681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_423_n 0.19698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_424_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_D1_c_79_n 0.0318507f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.14
cc_44 VPB N_D1_c_87_n 0.0355878f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.215
cc_45 VPB N_D1_c_88_n 0.01554f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.215
cc_46 VPB N_D1_c_89_n 0.0198827f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.29
cc_47 VPB D1 0.028742f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_48 VPB N_C1_M1004_g 0.0325172f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.84
cc_49 VPB N_C1_c_119_n 0.00557261f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.29
cc_50 VPB N_C1_c_124_n 0.018909f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.735
cc_51 VPB C1 0.00965929f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.735
cc_52 VPB N_B1_c_162_n 0.00155892f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.14
cc_53 VPB N_B1_M1009_g 0.038015f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.215
cc_54 VPB N_B1_c_168_n 0.0172095f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.29
cc_55 VPB B1 0.0015918f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_56 VPB N_A1_M1005_g 0.0209435f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.915
cc_57 VPB N_A1_c_208_n 0.0372045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB A1 0.00341349f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_59 VPB N_A1_c_206_n 0.0297463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A2_M1001_g 0.0241128f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.84
cc_61 VPB N_A2_c_260_n 0.0445985f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.29
cc_62 VPB N_A2_c_261_n 0.00600099f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.735
cc_63 VPB N_A2_c_255_n 0.0313335f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_64 VPB A2 0.0298016f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_65 VPB N_Y_c_302_n 0.00782248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_Y_c_303_n 0.0221704f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.735
cc_67 VPB N_Y_c_298_n 0.0128533f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_68 VPB N_A_318_483#_c_349_n 0.00389279f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.445
cc_69 VPB N_A_318_483#_c_350_n 0.00948911f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.29
cc_70 VPB N_A_318_483#_c_351_n 0.00191236f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.735
cc_71 VPB N_A_318_483#_c_352_n 0.00695802f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_72 VPB N_A_318_483#_c_353_n 0.0219878f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_73 VPB N_A_318_483#_c_354_n 0.00458706f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_74 VPB N_VPWR_c_385_n 0.00932704f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.215
cc_75 VPB N_VPWR_c_386_n 0.0588171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_387_n 0.0307594f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_77 VPB N_VPWR_c_384_n 0.0925157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_389_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 N_D1_M1002_g N_C1_M1008_g 0.0216137f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_80 N_D1_c_85_n N_C1_M1008_g 0.00165492f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_81 N_D1_c_79_n N_C1_M1004_g 0.00157508f $X=0.36 $Y=2.14 $X2=0 $Y2=0
cc_82 N_D1_c_87_n N_C1_M1004_g 0.0633708f $X=0.72 $Y=2.215 $X2=0 $Y2=0
cc_83 N_D1_c_83_n N_C1_c_119_n 0.00406453f $X=0.27 $Y=1.51 $X2=0 $Y2=0
cc_84 N_D1_c_79_n N_C1_c_124_n 0.00406453f $X=0.36 $Y=2.14 $X2=0 $Y2=0
cc_85 N_D1_c_87_n C1 0.00606041f $X=0.72 $Y=2.215 $X2=0 $Y2=0
cc_86 N_D1_c_85_n N_C1_c_121_n 0.00406453f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_87 N_D1_c_88_n N_Y_c_302_n 0.00687484f $X=0.435 $Y=2.215 $X2=0 $Y2=0
cc_88 N_D1_M1002_g N_Y_c_297_n 0.00345987f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_89 N_D1_c_80_n N_Y_c_298_n 0.00198435f $X=0.65 $Y=0.915 $X2=0 $Y2=0
cc_90 N_D1_c_87_n N_Y_c_298_n 0.0162586f $X=0.72 $Y=2.215 $X2=0 $Y2=0
cc_91 N_D1_c_89_n N_Y_c_298_n 0.00348255f $X=0.795 $Y=2.29 $X2=0 $Y2=0
cc_92 D1 N_Y_c_298_n 0.0879506f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_D1_c_85_n N_Y_c_298_n 0.00925574f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_94 N_D1_c_80_n N_Y_c_300_n 0.0132456f $X=0.65 $Y=0.915 $X2=0 $Y2=0
cc_95 N_D1_M1002_g N_Y_c_300_n 0.00590987f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_96 D1 N_Y_c_300_n 0.0193737f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_97 N_D1_c_89_n N_VPWR_c_386_n 0.00545548f $X=0.795 $Y=2.29 $X2=0 $Y2=0
cc_98 N_D1_c_89_n N_VPWR_c_384_n 0.011419f $X=0.795 $Y=2.29 $X2=0 $Y2=0
cc_99 N_D1_c_80_n N_VGND_c_414_n 5.86586e-19 $X=0.65 $Y=0.915 $X2=0 $Y2=0
cc_100 N_D1_c_81_n N_VGND_c_414_n 0.0071475f $X=0.435 $Y=0.915 $X2=0 $Y2=0
cc_101 N_D1_M1002_g N_VGND_c_414_n 0.00370983f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_102 D1 N_VGND_c_414_n 0.00163808f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_103 N_D1_M1002_g N_VGND_c_419_n 0.00585385f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_104 N_D1_M1002_g N_VGND_c_423_n 0.00735078f $X=0.725 $Y=0.445 $X2=0 $Y2=0
cc_105 D1 N_VGND_c_423_n 0.0108824f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_106 N_C1_c_121_n N_B1_c_162_n 0.0301104f $X=1.065 $Y=1.395 $X2=0 $Y2=0
cc_107 N_C1_c_124_n N_B1_M1009_g 0.0301104f $X=1.065 $Y=1.9 $X2=0 $Y2=0
cc_108 N_C1_M1008_g N_B1_M1006_g 0.02514f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_109 N_C1_c_119_n N_B1_c_168_n 0.0301104f $X=1.065 $Y=1.735 $X2=0 $Y2=0
cc_110 N_C1_M1008_g B1 5.76938e-19 $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_111 C1 B1 0.0564526f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_C1_M1008_g N_B1_c_165_n 0.0301104f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_113 C1 N_B1_c_165_n 0.0153606f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_C1_M1008_g N_Y_c_297_n 0.00193726f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_115 N_C1_M1008_g N_Y_c_298_n 0.00383459f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_116 N_C1_M1004_g N_Y_c_298_n 0.00110098f $X=1.155 $Y=2.735 $X2=0 $Y2=0
cc_117 C1 N_Y_c_298_n 0.0813282f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_C1_c_121_n N_Y_c_298_n 0.00611489f $X=1.065 $Y=1.395 $X2=0 $Y2=0
cc_119 N_C1_M1008_g N_Y_c_299_n 0.0153075f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_120 C1 N_Y_c_300_n 0.0305187f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_121 N_C1_c_121_n N_Y_c_300_n 0.00393194f $X=1.065 $Y=1.395 $X2=0 $Y2=0
cc_122 C1 A_174_483# 0.00580823f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_123 C1 A_246_483# 0.00553472f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_124 N_C1_M1004_g N_A_318_483#_c_349_n 0.00127992f $X=1.155 $Y=2.735 $X2=0
+ $Y2=0
cc_125 C1 N_A_318_483#_c_349_n 0.0459981f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_126 C1 N_A_318_483#_c_351_n 0.0127607f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 N_C1_M1004_g N_VPWR_c_386_n 0.0035749f $X=1.155 $Y=2.735 $X2=0 $Y2=0
cc_128 C1 N_VPWR_c_386_n 0.0110924f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_129 N_C1_M1004_g N_VPWR_c_384_n 0.00485911f $X=1.155 $Y=2.735 $X2=0 $Y2=0
cc_130 C1 N_VPWR_c_384_n 0.0124359f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_131 N_C1_M1008_g N_VGND_c_415_n 0.00187332f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_132 N_C1_M1008_g N_VGND_c_419_n 0.00585385f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_133 N_C1_M1008_g N_VGND_c_423_n 0.00635314f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_134 N_B1_M1006_g N_A1_M1000_g 0.0322753f $X=1.655 $Y=0.445 $X2=0 $Y2=0
cc_135 B1 N_A1_M1000_g 0.00268547f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B1_c_165_n N_A1_M1000_g 0.0217833f $X=1.635 $Y=1.355 $X2=0 $Y2=0
cc_137 N_B1_M1009_g N_A1_c_208_n 0.0196237f $X=1.515 $Y=2.735 $X2=0 $Y2=0
cc_138 B1 N_A1_c_208_n 9.37789e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_139 B1 A1 0.0534437f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B1_c_165_n A1 2.32748e-19 $X=1.635 $Y=1.355 $X2=0 $Y2=0
cc_141 N_B1_c_162_n N_A1_c_206_n 0.0217833f $X=1.62 $Y=1.68 $X2=0 $Y2=0
cc_142 N_B1_M1009_g N_A1_c_206_n 0.00719929f $X=1.515 $Y=2.735 $X2=0 $Y2=0
cc_143 B1 N_A1_c_206_n 0.0355582f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_144 N_B1_M1006_g N_Y_c_299_n 0.0129236f $X=1.655 $Y=0.445 $X2=0 $Y2=0
cc_145 B1 N_Y_c_299_n 0.0169275f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_146 N_B1_c_165_n N_Y_c_299_n 0.00515847f $X=1.635 $Y=1.355 $X2=0 $Y2=0
cc_147 N_B1_M1006_g N_Y_c_301_n 0.0036154f $X=1.655 $Y=0.445 $X2=0 $Y2=0
cc_148 B1 N_Y_c_301_n 0.0475501f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_149 N_B1_c_165_n N_Y_c_301_n 0.00171814f $X=1.635 $Y=1.355 $X2=0 $Y2=0
cc_150 N_B1_M1009_g N_A_318_483#_c_349_n 0.0122011f $X=1.515 $Y=2.735 $X2=0
+ $Y2=0
cc_151 B1 N_A_318_483#_c_350_n 0.030275f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B1_M1009_g N_A_318_483#_c_351_n 0.00470874f $X=1.515 $Y=2.735 $X2=0
+ $Y2=0
cc_153 N_B1_c_168_n N_A_318_483#_c_351_n 0.0056435f $X=1.62 $Y=1.86 $X2=0 $Y2=0
cc_154 B1 N_A_318_483#_c_351_n 0.0246944f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B1_M1009_g N_VPWR_c_386_n 0.00511657f $X=1.515 $Y=2.735 $X2=0 $Y2=0
cc_156 N_B1_M1009_g N_VPWR_c_384_n 0.00954952f $X=1.515 $Y=2.735 $X2=0 $Y2=0
cc_157 N_B1_M1006_g N_VGND_c_415_n 0.00329429f $X=1.655 $Y=0.445 $X2=0 $Y2=0
cc_158 N_B1_M1006_g N_VGND_c_421_n 0.00585385f $X=1.655 $Y=0.445 $X2=0 $Y2=0
cc_159 N_B1_M1006_g N_VGND_c_423_n 0.00639414f $X=1.655 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A1_M1000_g N_A2_M1007_g 0.0528715f $X=2.085 $Y=0.445 $X2=0 $Y2=0
cc_161 A1 N_A2_M1007_g 0.00302575f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_162 A1 N_A2_c_253_n 0.0134473f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_163 A1 N_A2_c_254_n 0.00299236f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_164 N_A1_c_206_n N_A2_c_254_n 0.0185613f $X=2.52 $Y=1.37 $X2=0 $Y2=0
cc_165 A1 N_A2_c_260_n 5.27096e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_166 N_A1_M1005_g N_A2_c_261_n 0.00890042f $X=1.945 $Y=2.735 $X2=0 $Y2=0
cc_167 N_A1_c_208_n N_A2_c_261_n 0.0089218f $X=2.1 $Y=2.1 $X2=0 $Y2=0
cc_168 A1 N_A2_c_261_n 2.75996e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_169 N_A1_c_206_n N_A2_c_261_n 0.0157226f $X=2.52 $Y=1.37 $X2=0 $Y2=0
cc_170 A1 A2 0.081463f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_171 N_A1_c_206_n A2 7.07714e-19 $X=2.52 $Y=1.37 $X2=0 $Y2=0
cc_172 A1 N_A2_c_258_n 0.00736268f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_173 N_A1_c_206_n N_A2_c_258_n 0.0343018f $X=2.52 $Y=1.37 $X2=0 $Y2=0
cc_174 N_A1_M1000_g N_Y_c_301_n 0.0217686f $X=2.085 $Y=0.445 $X2=0 $Y2=0
cc_175 A1 N_Y_c_301_n 0.0199225f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_176 N_A1_c_206_n N_Y_c_301_n 7.82016e-19 $X=2.52 $Y=1.37 $X2=0 $Y2=0
cc_177 N_A1_c_208_n N_A_318_483#_c_349_n 0.00520611f $X=2.1 $Y=2.1 $X2=0 $Y2=0
cc_178 N_A1_c_208_n N_A_318_483#_c_350_n 0.0225217f $X=2.1 $Y=2.1 $X2=0 $Y2=0
cc_179 A1 N_A_318_483#_c_350_n 0.028636f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_180 N_A1_c_206_n N_A_318_483#_c_350_n 0.00919669f $X=2.52 $Y=1.37 $X2=0 $Y2=0
cc_181 N_A1_M1005_g N_A_318_483#_c_354_n 8.39383e-19 $X=1.945 $Y=2.735 $X2=0
+ $Y2=0
cc_182 N_A1_M1005_g N_VPWR_c_385_n 0.0032248f $X=1.945 $Y=2.735 $X2=0 $Y2=0
cc_183 N_A1_c_208_n N_VPWR_c_385_n 0.00415699f $X=2.1 $Y=2.1 $X2=0 $Y2=0
cc_184 N_A1_M1005_g N_VPWR_c_386_n 0.00545548f $X=1.945 $Y=2.735 $X2=0 $Y2=0
cc_185 N_A1_M1005_g N_VPWR_c_384_n 0.010533f $X=1.945 $Y=2.735 $X2=0 $Y2=0
cc_186 N_A1_M1000_g N_VGND_c_416_n 0.00164766f $X=2.085 $Y=0.445 $X2=0 $Y2=0
cc_187 A1 N_VGND_c_416_n 0.0211278f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_188 N_A1_M1000_g N_VGND_c_421_n 0.00362854f $X=2.085 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A1_M1000_g N_VGND_c_423_n 0.00528707f $X=2.085 $Y=0.445 $X2=0 $Y2=0
cc_190 A1 N_VGND_c_423_n 0.00308656f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_191 N_A2_M1007_g N_Y_c_301_n 0.00831525f $X=2.445 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A2_c_260_n N_A_318_483#_c_350_n 0.00560586f $X=2.925 $Y=2.19 $X2=0
+ $Y2=0
cc_193 N_A2_c_261_n N_A_318_483#_c_350_n 0.00934601f $X=2.55 $Y=2.19 $X2=0 $Y2=0
cc_194 A2 N_A_318_483#_c_350_n 0.0146787f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_195 N_A2_M1001_g N_A_318_483#_c_352_n 0.00192766f $X=2.475 $Y=2.735 $X2=0
+ $Y2=0
cc_196 N_A2_c_260_n N_A_318_483#_c_352_n 0.00378417f $X=2.925 $Y=2.19 $X2=0
+ $Y2=0
cc_197 N_A2_M1001_g N_A_318_483#_c_353_n 0.00498071f $X=2.475 $Y=2.735 $X2=0
+ $Y2=0
cc_198 N_A2_M1001_g N_A_318_483#_c_354_n 0.00468641f $X=2.475 $Y=2.735 $X2=0
+ $Y2=0
cc_199 N_A2_c_260_n N_A_318_483#_c_354_n 0.00752995f $X=2.925 $Y=2.19 $X2=0
+ $Y2=0
cc_200 N_A2_c_261_n N_A_318_483#_c_354_n 6.43197e-19 $X=2.55 $Y=2.19 $X2=0 $Y2=0
cc_201 N_A2_M1001_g N_VPWR_c_385_n 0.00316252f $X=2.475 $Y=2.735 $X2=0 $Y2=0
cc_202 N_A2_M1001_g N_VPWR_c_387_n 0.00532839f $X=2.475 $Y=2.735 $X2=0 $Y2=0
cc_203 N_A2_M1001_g N_VPWR_c_384_n 0.0112072f $X=2.475 $Y=2.735 $X2=0 $Y2=0
cc_204 N_A2_M1007_g N_VGND_c_416_n 0.0110427f $X=2.445 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A2_c_253_n N_VGND_c_416_n 0.00397036f $X=2.925 $Y=0.89 $X2=0 $Y2=0
cc_206 N_A2_M1007_g N_VGND_c_421_n 0.00486043f $X=2.445 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A2_M1007_g N_VGND_c_423_n 0.00634722f $X=2.445 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A2_c_253_n N_VGND_c_423_n 0.0106198f $X=2.925 $Y=0.89 $X2=0 $Y2=0
cc_209 A2 N_VGND_c_423_n 0.0120784f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_210 N_Y_c_303_n N_VPWR_c_386_n 0.0214297f $X=0.55 $Y=2.56 $X2=0 $Y2=0
cc_211 N_Y_c_303_n N_VPWR_c_384_n 0.0123021f $X=0.55 $Y=2.56 $X2=0 $Y2=0
cc_212 N_Y_c_300_n N_VGND_c_414_n 0.00650106f $X=1.065 $Y=0.9 $X2=0 $Y2=0
cc_213 N_Y_c_299_n N_VGND_c_415_n 0.0227065f $X=1.735 $Y=0.9 $X2=0 $Y2=0
cc_214 N_Y_c_301_n N_VGND_c_416_n 0.0210845f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_215 N_Y_c_297_n N_VGND_c_419_n 0.0125251f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_216 N_Y_c_301_n N_VGND_c_421_n 0.0267527f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_217 N_Y_M1002_d N_VGND_c_423_n 0.00241536f $X=0.8 $Y=0.235 $X2=0 $Y2=0
cc_218 N_Y_M1006_d N_VGND_c_423_n 0.00228191f $X=1.73 $Y=0.235 $X2=0 $Y2=0
cc_219 N_Y_c_297_n N_VGND_c_423_n 0.00963317f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_220 N_Y_c_299_n N_VGND_c_423_n 0.00663295f $X=1.735 $Y=0.9 $X2=0 $Y2=0
cc_221 N_Y_c_300_n N_VGND_c_423_n 0.0109894f $X=1.065 $Y=0.9 $X2=0 $Y2=0
cc_222 N_Y_c_301_n N_VGND_c_423_n 0.0195699f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_223 N_Y_c_301_n A_432_47# 0.00422339f $X=1.87 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_224 N_A_318_483#_c_349_n N_VPWR_c_385_n 0.00142637f $X=1.73 $Y=2.56 $X2=0
+ $Y2=0
cc_225 N_A_318_483#_c_350_n N_VPWR_c_385_n 0.0261338f $X=2.54 $Y=2.135 $X2=0
+ $Y2=0
cc_226 N_A_318_483#_c_352_n N_VPWR_c_385_n 0.0253006f $X=2.697 $Y=2.552 $X2=0
+ $Y2=0
cc_227 N_A_318_483#_c_349_n N_VPWR_c_386_n 0.0196723f $X=1.73 $Y=2.56 $X2=0
+ $Y2=0
cc_228 N_A_318_483#_c_353_n N_VPWR_c_387_n 0.021066f $X=2.69 $Y=2.56 $X2=0 $Y2=0
cc_229 N_A_318_483#_c_349_n N_VPWR_c_384_n 0.0112265f $X=1.73 $Y=2.56 $X2=0
+ $Y2=0
cc_230 N_A_318_483#_c_353_n N_VPWR_c_384_n 0.0120681f $X=2.69 $Y=2.56 $X2=0
+ $Y2=0
cc_231 N_VGND_c_423_n A_432_47# 0.00537988f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
