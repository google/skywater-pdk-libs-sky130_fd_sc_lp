* File: sky130_fd_sc_lp__and4_4.pxi.spice
* Created: Wed Sep  2 09:32:59 2020
* 
x_PM_SKY130_FD_SC_LP__AND4_4%A N_A_c_80_n N_A_M1009_g N_A_c_81_n N_A_M1000_g A A
+ PM_SKY130_FD_SC_LP__AND4_4%A
x_PM_SKY130_FD_SC_LP__AND4_4%B N_B_M1003_g N_B_M1007_g B B N_B_c_103_n
+ N_B_c_104_n PM_SKY130_FD_SC_LP__AND4_4%B
x_PM_SKY130_FD_SC_LP__AND4_4%C N_C_M1008_g N_C_M1006_g C N_C_c_139_n
+ PM_SKY130_FD_SC_LP__AND4_4%C
x_PM_SKY130_FD_SC_LP__AND4_4%D N_D_M1015_g N_D_M1012_g D N_D_c_173_n
+ PM_SKY130_FD_SC_LP__AND4_4%D
x_PM_SKY130_FD_SC_LP__AND4_4%A_58_47# N_A_58_47#_M1009_s N_A_58_47#_M1000_d
+ N_A_58_47#_M1006_d N_A_58_47#_M1002_g N_A_58_47#_M1001_g N_A_58_47#_M1004_g
+ N_A_58_47#_M1005_g N_A_58_47#_M1011_g N_A_58_47#_M1010_g N_A_58_47#_M1014_g
+ N_A_58_47#_M1013_g N_A_58_47#_c_344_p N_A_58_47#_c_226_n N_A_58_47#_c_227_n
+ N_A_58_47#_c_233_n N_A_58_47#_c_220_n N_A_58_47#_c_221_n N_A_58_47#_c_240_n
+ N_A_58_47#_c_222_n N_A_58_47#_c_211_n N_A_58_47#_c_212_n N_A_58_47#_c_213_n
+ N_A_58_47#_c_214_n N_A_58_47#_c_225_n N_A_58_47#_c_215_n
+ PM_SKY130_FD_SC_LP__AND4_4%A_58_47#
x_PM_SKY130_FD_SC_LP__AND4_4%VPWR N_VPWR_M1000_s N_VPWR_M1007_d N_VPWR_M1012_d
+ N_VPWR_M1005_d N_VPWR_M1013_d N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n
+ N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_362_n
+ N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n VPWR N_VPWR_c_366_n
+ N_VPWR_c_367_n N_VPWR_c_354_n N_VPWR_c_369_n N_VPWR_c_370_n
+ PM_SKY130_FD_SC_LP__AND4_4%VPWR
x_PM_SKY130_FD_SC_LP__AND4_4%X N_X_M1002_s N_X_M1011_s N_X_M1001_s N_X_M1010_s
+ N_X_c_467_n N_X_c_481_p N_X_c_420_n N_X_c_421_n N_X_c_427_n N_X_c_428_n
+ N_X_c_448_n N_X_c_471_n N_X_c_429_n N_X_c_422_n N_X_c_423_n N_X_c_430_n X X X
+ X X PM_SKY130_FD_SC_LP__AND4_4%X
x_PM_SKY130_FD_SC_LP__AND4_4%VGND N_VGND_M1015_d N_VGND_M1004_d N_VGND_M1014_d
+ N_VGND_c_494_n N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n N_VGND_c_498_n
+ N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n VGND N_VGND_c_502_n
+ N_VGND_c_503_n N_VGND_c_504_n PM_SKY130_FD_SC_LP__AND4_4%VGND
cc_1 VNB N_A_c_80_n 0.0216251f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.185
cc_2 VNB N_A_c_81_n 0.0596821f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.725
cc_3 VNB A 0.0212372f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B_M1007_g 0.00816884f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_5 VNB B 0.00902078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B_c_103_n 0.0276094f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_7 VNB N_B_c_104_n 0.0169284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_C_M1008_g 0.0199015f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.655
cc_9 VNB N_C_M1006_g 0.00677949f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB C 0.00588324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_c_139_n 0.0306723f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_12 VNB N_D_M1015_g 0.0202767f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.655
cc_13 VNB N_D_M1012_g 0.0067132f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB D 0.00217658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D_c_173_n 0.0326717f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_16 VNB N_A_58_47#_M1002_g 0.0238884f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_17 VNB N_A_58_47#_M1004_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_58_47#_M1011_g 0.0222627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_58_47#_M1014_g 0.0284217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_58_47#_c_211_n 0.00256644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_58_47#_c_212_n 7.22757e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_58_47#_c_213_n 0.0015776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_58_47#_c_214_n 0.0835064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_58_47#_c_215_n 0.00130582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_354_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_420_n 0.00310505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_421_n 0.0025979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_422_n 0.0104727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_423_n 0.00190113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB X 0.0385526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB X 0.00882499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 0.0230589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_494_n 0.00503465f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_34 VNB N_VGND_c_495_n 3.31813e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_496_n 0.0149762f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.665
cc_36 VNB N_VGND_c_497_n 0.00439483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_498_n 0.0700751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_499_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_500_n 0.0167855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_501_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_502_n 0.0172686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_503_n 0.264905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_504_n 0.00442067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_A_c_81_n 0.030415f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.725
cc_45 VPB A 0.0118113f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_46 VPB N_B_M1007_g 0.0211634f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_47 VPB N_C_M1006_g 0.0211667f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_48 VPB N_D_M1012_g 0.0210539f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_49 VPB N_A_58_47#_M1001_g 0.0200496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_58_47#_M1005_g 0.0185138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_58_47#_M1010_g 0.0185219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_58_47#_M1013_g 0.0223753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_58_47#_c_220_n 0.00692389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_58_47#_c_221_n 0.00324156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_58_47#_c_222_n 0.00501441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_58_47#_c_212_n 0.001037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_58_47#_c_214_n 0.0151402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_58_47#_c_225_n 0.00768186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_355_n 0.015284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_356_n 0.0482776f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.665
cc_61 VPB N_VPWR_c_357_n 0.0155418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_358_n 0.0043916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_359_n 0.00445607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_360_n 3.23223e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_361_n 0.040815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_362_n 0.0178386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_363_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_364_n 0.0166915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_365_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_366_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_367_n 0.017577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_354_n 0.0663175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_369_n 0.00631492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_370_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_X_c_427_n 0.00316451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_X_c_428_n 0.00194676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_X_c_429_n 0.0291619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_X_c_430_n 0.00149902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.00694732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 N_A_c_81_n N_B_M1007_g 0.027572f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_81 A N_B_M1007_g 8.18048e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_c_81_n B 0.014685f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_83 A B 0.0252047f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A_c_81_n N_B_c_103_n 0.0455387f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_85 N_A_c_80_n N_B_c_104_n 0.0455387f $X=0.63 $Y=1.185 $X2=0 $Y2=0
cc_86 N_A_c_80_n N_A_58_47#_c_226_n 0.0116531f $X=0.63 $Y=1.185 $X2=0 $Y2=0
cc_87 N_A_c_81_n N_A_58_47#_c_227_n 0.00568217f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_88 A N_A_58_47#_c_227_n 0.0123784f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A_c_81_n N_A_58_47#_c_221_n 0.00253514f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_90 N_A_c_81_n N_VPWR_c_356_n 0.0258024f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_91 A N_VPWR_c_356_n 0.0184319f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A_c_81_n N_VPWR_c_357_n 0.00486043f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_93 N_A_c_81_n N_VPWR_c_354_n 0.0082726f $X=0.63 $Y=1.725 $X2=0 $Y2=0
cc_94 N_A_c_80_n N_VGND_c_498_n 0.00585385f $X=0.63 $Y=1.185 $X2=0 $Y2=0
cc_95 N_A_c_80_n N_VGND_c_503_n 0.00754594f $X=0.63 $Y=1.185 $X2=0 $Y2=0
cc_96 B N_C_M1008_g 0.00211147f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B_c_103_n N_C_M1008_g 0.0205733f $X=1.08 $Y=1.35 $X2=0 $Y2=0
cc_98 N_B_c_104_n N_C_M1008_g 0.0386968f $X=1.08 $Y=1.185 $X2=0 $Y2=0
cc_99 N_B_M1007_g N_C_M1006_g 0.0381894f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_100 B C 0.0264243f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B_c_103_n C 3.00625e-19 $X=1.08 $Y=1.35 $X2=0 $Y2=0
cc_102 N_B_M1007_g N_C_c_139_n 0.00103226f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_103 B N_A_58_47#_c_226_n 0.0466942f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B_c_103_n N_A_58_47#_c_226_n 0.00425874f $X=1.08 $Y=1.35 $X2=0 $Y2=0
cc_105 N_B_c_104_n N_A_58_47#_c_226_n 0.0121264f $X=1.08 $Y=1.185 $X2=0 $Y2=0
cc_106 N_B_M1007_g N_A_58_47#_c_233_n 0.0157033f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_107 N_B_M1007_g N_A_58_47#_c_220_n 0.0117982f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_108 B N_A_58_47#_c_220_n 0.0184104f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B_c_103_n N_A_58_47#_c_220_n 0.00235248f $X=1.08 $Y=1.35 $X2=0 $Y2=0
cc_110 N_B_M1007_g N_A_58_47#_c_221_n 0.00172707f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_111 B N_A_58_47#_c_221_n 0.0177813f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B_c_103_n N_A_58_47#_c_221_n 0.00182638f $X=1.08 $Y=1.35 $X2=0 $Y2=0
cc_113 N_B_M1007_g N_A_58_47#_c_240_n 7.5774e-19 $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B_M1007_g N_VPWR_c_356_n 8.7487e-19 $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B_M1007_g N_VPWR_c_357_n 0.00541359f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_VPWR_c_358_n 0.00777641f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B_M1007_g N_VPWR_c_354_n 0.0100974f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B_c_104_n N_VGND_c_498_n 0.00585385f $X=1.08 $Y=1.185 $X2=0 $Y2=0
cc_119 N_B_c_104_n N_VGND_c_503_n 0.00670341f $X=1.08 $Y=1.185 $X2=0 $Y2=0
cc_120 N_C_M1008_g N_D_M1015_g 0.0374157f $X=1.53 $Y=0.655 $X2=0 $Y2=0
cc_121 C N_D_M1015_g 0.00194141f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_C_M1006_g N_D_M1012_g 0.0277675f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_123 C D 0.0263443f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_124 N_C_c_139_n D 3.74634e-19 $X=1.62 $Y=1.375 $X2=0 $Y2=0
cc_125 N_C_c_139_n N_D_c_173_n 0.0206141f $X=1.62 $Y=1.375 $X2=0 $Y2=0
cc_126 N_C_M1008_g N_A_58_47#_c_226_n 0.0145802f $X=1.53 $Y=0.655 $X2=0 $Y2=0
cc_127 C N_A_58_47#_c_226_n 0.0226312f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_C_c_139_n N_A_58_47#_c_226_n 0.0011003f $X=1.62 $Y=1.375 $X2=0 $Y2=0
cc_129 N_C_M1006_g N_A_58_47#_c_233_n 7.59342e-19 $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_130 N_C_M1006_g N_A_58_47#_c_220_n 0.0116798f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_131 C N_A_58_47#_c_220_n 0.0108624f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 N_C_c_139_n N_A_58_47#_c_220_n 0.00240758f $X=1.62 $Y=1.375 $X2=0 $Y2=0
cc_133 N_C_M1006_g N_A_58_47#_c_240_n 0.016066f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_134 N_C_M1006_g N_A_58_47#_c_225_n 0.0018847f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_135 C N_A_58_47#_c_225_n 0.0102942f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_C_c_139_n N_A_58_47#_c_225_n 5.38111e-19 $X=1.62 $Y=1.375 $X2=0 $Y2=0
cc_137 N_C_M1006_g N_VPWR_c_358_n 0.00785102f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_138 N_C_M1006_g N_VPWR_c_362_n 0.00541359f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_139 N_C_M1006_g N_VPWR_c_354_n 0.0100974f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_140 N_C_M1008_g N_VGND_c_498_n 0.00585385f $X=1.53 $Y=0.655 $X2=0 $Y2=0
cc_141 N_C_M1008_g N_VGND_c_503_n 0.00715943f $X=1.53 $Y=0.655 $X2=0 $Y2=0
cc_142 N_D_M1015_g N_A_58_47#_M1002_g 0.0262256f $X=2.07 $Y=0.655 $X2=0 $Y2=0
cc_143 D N_A_58_47#_M1002_g 3.1759e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_144 N_D_c_173_n N_A_58_47#_M1002_g 0.01675f $X=2.16 $Y=1.375 $X2=0 $Y2=0
cc_145 N_D_M1015_g N_A_58_47#_c_226_n 0.0134742f $X=2.07 $Y=0.655 $X2=0 $Y2=0
cc_146 D N_A_58_47#_c_226_n 0.0168406f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_147 N_D_c_173_n N_A_58_47#_c_226_n 0.00326283f $X=2.16 $Y=1.375 $X2=0 $Y2=0
cc_148 N_D_M1012_g N_A_58_47#_c_240_n 0.01474f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_149 N_D_M1012_g N_A_58_47#_c_222_n 0.0127921f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_150 D N_A_58_47#_c_222_n 0.0149267f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_151 N_D_c_173_n N_A_58_47#_c_222_n 0.00327208f $X=2.16 $Y=1.375 $X2=0 $Y2=0
cc_152 N_D_M1015_g N_A_58_47#_c_211_n 0.00329638f $X=2.07 $Y=0.655 $X2=0 $Y2=0
cc_153 D N_A_58_47#_c_211_n 0.0158469f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_D_c_173_n N_A_58_47#_c_211_n 0.00135187f $X=2.16 $Y=1.375 $X2=0 $Y2=0
cc_155 N_D_M1012_g N_A_58_47#_c_212_n 0.00325473f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_156 N_D_M1012_g N_A_58_47#_c_214_n 0.0363947f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_157 N_D_M1012_g N_A_58_47#_c_225_n 0.00161219f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_158 D N_A_58_47#_c_225_n 5.98581e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_159 N_D_M1012_g N_A_58_47#_c_215_n 0.00114023f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_160 D N_A_58_47#_c_215_n 0.0103581f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_161 N_D_c_173_n N_A_58_47#_c_215_n 9.49874e-19 $X=2.16 $Y=1.375 $X2=0 $Y2=0
cc_162 N_D_M1012_g N_VPWR_c_359_n 0.00804301f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_163 N_D_M1012_g N_VPWR_c_362_n 0.00564131f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_164 N_D_M1012_g N_VPWR_c_354_n 0.0106023f $X=2.07 $Y=2.465 $X2=0 $Y2=0
cc_165 N_D_M1015_g N_VGND_c_494_n 0.00607613f $X=2.07 $Y=0.655 $X2=0 $Y2=0
cc_166 N_D_M1015_g N_VGND_c_498_n 0.00585385f $X=2.07 $Y=0.655 $X2=0 $Y2=0
cc_167 N_D_M1015_g N_VGND_c_503_n 0.00705709f $X=2.07 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A_58_47#_c_220_n N_VPWR_M1007_d 0.00378554f $X=1.685 $Y=1.84 $X2=0
+ $Y2=0
cc_169 N_A_58_47#_c_222_n N_VPWR_M1012_d 0.00368975f $X=2.425 $Y=1.84 $X2=0
+ $Y2=0
cc_170 N_A_58_47#_c_233_n N_VPWR_c_357_n 0.0160289f $X=0.845 $Y=1.98 $X2=0 $Y2=0
cc_171 N_A_58_47#_c_220_n N_VPWR_c_358_n 0.0246333f $X=1.685 $Y=1.84 $X2=0 $Y2=0
cc_172 N_A_58_47#_M1001_g N_VPWR_c_359_n 0.0121739f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_58_47#_c_222_n N_VPWR_c_359_n 0.0246034f $X=2.425 $Y=1.84 $X2=0 $Y2=0
cc_174 N_A_58_47#_M1001_g N_VPWR_c_360_n 7.55501e-19 $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_58_47#_M1005_g N_VPWR_c_360_n 0.0142073f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_58_47#_M1010_g N_VPWR_c_360_n 0.0140168f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_58_47#_M1013_g N_VPWR_c_360_n 7.21513e-19 $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_58_47#_M1010_g N_VPWR_c_361_n 7.21513e-19 $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_58_47#_M1013_g N_VPWR_c_361_n 0.0150803f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_58_47#_c_240_n N_VPWR_c_362_n 0.0185828f $X=1.855 $Y=1.98 $X2=0 $Y2=0
cc_181 N_A_58_47#_M1001_g N_VPWR_c_364_n 0.00585385f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_58_47#_M1005_g N_VPWR_c_364_n 0.00486043f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_58_47#_M1010_g N_VPWR_c_366_n 0.00486043f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_58_47#_M1013_g N_VPWR_c_366_n 0.00486043f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_58_47#_M1000_d N_VPWR_c_354_n 0.00380103f $X=0.705 $Y=1.835 $X2=0
+ $Y2=0
cc_186 N_A_58_47#_M1006_d N_VPWR_c_354_n 0.00223559f $X=1.715 $Y=1.835 $X2=0
+ $Y2=0
cc_187 N_A_58_47#_M1001_g N_VPWR_c_354_n 0.0111271f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_58_47#_M1005_g N_VPWR_c_354_n 0.00824727f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_58_47#_M1010_g N_VPWR_c_354_n 0.00824727f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_58_47#_M1013_g N_VPWR_c_354_n 0.00824727f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_58_47#_c_233_n N_VPWR_c_354_n 0.010019f $X=0.845 $Y=1.98 $X2=0 $Y2=0
cc_192 N_A_58_47#_c_240_n N_VPWR_c_354_n 0.0122144f $X=1.855 $Y=1.98 $X2=0 $Y2=0
cc_193 N_A_58_47#_M1004_g N_X_c_420_n 0.0137831f $X=3.075 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A_58_47#_M1011_g N_X_c_420_n 0.01419f $X=3.505 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_58_47#_c_213_n N_X_c_420_n 0.0447065f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_196 N_A_58_47#_c_214_n N_X_c_420_n 0.00244902f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_197 N_A_58_47#_M1002_g N_X_c_421_n 0.0013216f $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_198 N_A_58_47#_c_211_n N_X_c_421_n 0.0126453f $X=2.51 $Y=1.415 $X2=0 $Y2=0
cc_199 N_A_58_47#_c_213_n N_X_c_421_n 0.0139138f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_200 N_A_58_47#_c_214_n N_X_c_421_n 0.00255521f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_201 N_A_58_47#_M1005_g N_X_c_427_n 0.0129381f $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A_58_47#_M1010_g N_X_c_427_n 0.0130468f $X=3.505 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A_58_47#_c_213_n N_X_c_427_n 0.0428812f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_204 N_A_58_47#_c_214_n N_X_c_427_n 0.00243312f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_205 N_A_58_47#_M1001_g N_X_c_428_n 4.89726e-19 $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_58_47#_c_222_n N_X_c_428_n 0.00911097f $X=2.425 $Y=1.84 $X2=0 $Y2=0
cc_207 N_A_58_47#_c_213_n N_X_c_428_n 0.014105f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_208 N_A_58_47#_c_214_n N_X_c_428_n 0.00254241f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_209 N_A_58_47#_M1014_g N_X_c_448_n 0.0102503f $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A_58_47#_M1013_g N_X_c_429_n 0.0150769f $X=3.935 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_58_47#_c_213_n N_X_c_429_n 0.0286754f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_212 N_A_58_47#_c_214_n N_X_c_429_n 0.0060828f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_213 N_A_58_47#_M1014_g N_X_c_422_n 0.0146672f $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A_58_47#_c_213_n N_X_c_422_n 0.0264831f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_215 N_A_58_47#_c_214_n N_X_c_422_n 0.00612256f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_216 N_A_58_47#_M1014_g N_X_c_423_n 0.00205286f $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A_58_47#_c_213_n N_X_c_423_n 0.0185299f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_218 N_A_58_47#_c_214_n N_X_c_423_n 0.00255521f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_219 N_A_58_47#_c_213_n N_X_c_430_n 0.014105f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_220 N_A_58_47#_c_214_n N_X_c_430_n 0.00254241f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_221 N_A_58_47#_M1014_g X 0.00331729f $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A_58_47#_M1014_g X 0.00275073f $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_223 N_A_58_47#_M1013_g X 0.00302858f $X=3.935 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_58_47#_c_213_n X 0.0138877f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_225 N_A_58_47#_c_214_n X 0.00824949f $X=4.095 $Y=1.5 $X2=0 $Y2=0
cc_226 N_A_58_47#_c_226_n A_141_47# 0.00298571f $X=2.425 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_58_47#_c_226_n A_213_47# 0.0102957f $X=2.425 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_58_47#_c_226_n A_321_47# 0.0115791f $X=2.425 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_229 N_A_58_47#_c_226_n N_VGND_M1015_d 0.00889609f $X=2.425 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_230 N_A_58_47#_c_211_n N_VGND_M1015_d 5.56021e-19 $X=2.51 $Y=1.415 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A_58_47#_M1002_g N_VGND_c_494_n 0.00659056f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_232 N_A_58_47#_c_226_n N_VGND_c_494_n 0.0251446f $X=2.425 $Y=0.945 $X2=0
+ $Y2=0
cc_233 N_A_58_47#_M1002_g N_VGND_c_495_n 6.6497e-19 $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_234 N_A_58_47#_M1004_g N_VGND_c_495_n 0.0113349f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_235 N_A_58_47#_M1011_g N_VGND_c_495_n 0.0112586f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_236 N_A_58_47#_M1014_g N_VGND_c_495_n 7.0569e-19 $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_237 N_A_58_47#_M1011_g N_VGND_c_496_n 0.00486043f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_238 N_A_58_47#_M1014_g N_VGND_c_496_n 0.00579312f $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_58_47#_M1014_g N_VGND_c_497_n 0.00327527f $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_58_47#_c_344_p N_VGND_c_498_n 0.00781481f $X=0.415 $Y=0.525 $X2=0
+ $Y2=0
cc_241 N_A_58_47#_M1002_g N_VGND_c_500_n 0.00585385f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_242 N_A_58_47#_M1004_g N_VGND_c_500_n 0.00486043f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_243 N_A_58_47#_M1009_s N_VGND_c_503_n 0.003338f $X=0.29 $Y=0.235 $X2=0 $Y2=0
cc_244 N_A_58_47#_M1002_g N_VGND_c_503_n 0.0103938f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_245 N_A_58_47#_M1004_g N_VGND_c_503_n 0.00824727f $X=3.075 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_58_47#_M1011_g N_VGND_c_503_n 0.00824727f $X=3.505 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_A_58_47#_M1014_g N_VGND_c_503_n 0.0117246f $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_248 N_A_58_47#_c_344_p N_VGND_c_503_n 0.00689141f $X=0.415 $Y=0.525 $X2=0
+ $Y2=0
cc_249 N_A_58_47#_c_226_n N_VGND_c_503_n 0.0569239f $X=2.425 $Y=0.945 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_354_n N_X_M1001_s 0.00536646f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_251 N_VPWR_c_354_n N_X_M1010_s 0.00536646f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_364_n N_X_c_467_n 0.0124525f $X=3.125 $Y=3.33 $X2=0 $Y2=0
cc_253 N_VPWR_c_354_n N_X_c_467_n 0.00730901f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_254 N_VPWR_M1005_d N_X_c_427_n 0.00176461f $X=3.15 $Y=1.835 $X2=0 $Y2=0
cc_255 N_VPWR_c_360_n N_X_c_427_n 0.0170777f $X=3.29 $Y=2.2 $X2=0 $Y2=0
cc_256 N_VPWR_c_366_n N_X_c_471_n 0.0124525f $X=3.985 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_354_n N_X_c_471_n 0.00730901f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_258 N_VPWR_M1013_d N_X_c_429_n 0.0027239f $X=4.01 $Y=1.835 $X2=0 $Y2=0
cc_259 N_VPWR_c_361_n N_X_c_429_n 0.0220026f $X=4.15 $Y=2.2 $X2=0 $Y2=0
cc_260 N_X_c_420_n N_VGND_M1004_d 0.00176461f $X=3.625 $Y=1.15 $X2=0 $Y2=0
cc_261 N_X_c_422_n N_VGND_M1014_d 0.0025562f $X=4.43 $Y=1.15 $X2=0 $Y2=0
cc_262 N_X_c_420_n N_VGND_c_495_n 0.0170777f $X=3.625 $Y=1.15 $X2=0 $Y2=0
cc_263 N_X_c_448_n N_VGND_c_496_n 0.0143246f $X=3.72 $Y=0.42 $X2=0 $Y2=0
cc_264 N_X_c_422_n N_VGND_c_497_n 0.0160276f $X=4.43 $Y=1.15 $X2=0 $Y2=0
cc_265 X N_VGND_c_497_n 0.0395278f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_266 N_X_c_481_p N_VGND_c_500_n 0.0120977f $X=2.86 $Y=0.42 $X2=0 $Y2=0
cc_267 X N_VGND_c_502_n 0.0101072f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_268 N_X_M1002_s N_VGND_c_503_n 0.00571434f $X=2.72 $Y=0.235 $X2=0 $Y2=0
cc_269 N_X_M1011_s N_VGND_c_503_n 0.00380103f $X=3.58 $Y=0.235 $X2=0 $Y2=0
cc_270 N_X_c_481_p N_VGND_c_503_n 0.00691495f $X=2.86 $Y=0.42 $X2=0 $Y2=0
cc_271 N_X_c_448_n N_VGND_c_503_n 0.00916141f $X=3.72 $Y=0.42 $X2=0 $Y2=0
cc_272 X N_VGND_c_503_n 0.00947563f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_273 A_141_47# N_VGND_c_503_n 0.00314438f $X=0.705 $Y=0.235 $X2=0.415
+ $Y2=0.525
cc_274 A_213_47# N_VGND_c_503_n 0.00584965f $X=1.065 $Y=0.235 $X2=0.415
+ $Y2=0.525
cc_275 A_321_47# N_VGND_c_503_n 0.00584965f $X=1.605 $Y=0.235 $X2=0.415
+ $Y2=0.525
