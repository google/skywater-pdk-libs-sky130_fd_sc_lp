* File: sky130_fd_sc_lp__bufbuf_8.spice
* Created: Wed Sep  2 09:35:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__bufbuf_8.pex.spice"
.subckt sky130_fd_sc_lp__bufbuf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_117_265#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.5 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_117_265#_M1009_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1009_d N_A_117_265#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_117_265#_M1013_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1013_d N_A_117_265#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1020 N_VGND_M1020_d N_A_117_265#_M1020_g N_X_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1020_d N_A_117_265#_M1022_g N_X_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_A_117_265#_M1024_g N_X_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1365 AS=0.1176 PD=1.165 PS=1.12 NRD=3.564 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1004 N_A_117_265#_M1004_d N_A_837_23#_M1004_g N_VGND_M1024_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1365 PD=1.12 PS=1.165 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75003.7 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1010 N_A_117_265#_M1004_d N_A_837_23#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1018 N_A_117_265#_M1018_d N_A_837_23#_M1018_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A_1217_23#_M1007_g N_A_837_23#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1904 AS=0.2394 PD=1.67333 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75000.2 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1005 N_A_1217_23#_M1005_d N_A_M1005_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0952 PD=1.37 PS=0.836667 NRD=0 NRS=38.568 M=1 R=2.8 SA=75000.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_117_265#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1003 N_X_M1001_d N_A_117_265#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1006 N_X_M1006_d N_A_117_265#_M1006_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1008 N_X_M1006_d N_A_117_265#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1015 N_X_M1015_d N_A_117_265#_M1015_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1016 N_X_M1015_d N_A_117_265#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1021 N_X_M1021_d N_A_117_265#_M1021_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1023 N_X_M1021_d N_A_117_265#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.20475 PD=1.54 PS=1.585 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1000 N_A_117_265#_M1000_d N_A_837_23#_M1000_g N_VPWR_M1023_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.20475 PD=1.54 PS=1.585 NRD=0 NRS=7.0329 M=1 R=8.4
+ SA=75003.7 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1014 N_A_117_265#_M1000_d N_A_837_23#_M1014_g N_VPWR_M1014_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_A_117_265#_M1025_d N_A_837_23#_M1025_g N_VPWR_M1014_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A_1217_23#_M1019_g N_A_837_23#_M1019_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.268115 AS=0.3339 PD=2.16853 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1011 N_A_1217_23#_M1011_d N_A_M1011_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=30.7714 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
DX26_noxref VNB VPB NWDIODE A=14.1367 P=18.89
*
.include "sky130_fd_sc_lp__bufbuf_8.pxi.spice"
*
.ends
*
*
