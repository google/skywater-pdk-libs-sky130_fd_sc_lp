* File: sky130_fd_sc_lp__nor4_lp.spice
* Created: Wed Sep  2 10:10:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4_lp.pex.spice"
.subckt sky130_fd_sc_lp__nor4_lp  VNB VPB C D B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* D	D
* C	C
* VPB	VPB
* VNB	VNB
MM1007 A_138_57# N_C_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.9
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g A_138_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1008 A_296_57# N_D_M1008_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75002.1 A=0.063
+ P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_D_M1009_g A_296_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1002 A_454_57# N_B_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1010 N_Y_M1010_d N_B_M1010_g A_454_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1003 A_612_57# N_A_M1003_g N_Y_M1010_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g A_612_57# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_134_409#_M1005_d N_C_M1005_g N_A_27_409#_M1005_s VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_27_409#_M1000_d N_D_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1006 A_570_409# N_B_M1006_g N_A_134_409#_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g A_570_409# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.12 PD=2.57 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125000 A=0.25
+ P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.0827 P=12.53
c_42 VNB 0 1.85906e-19 $X=0 $Y=0
c_70 VPB 0 1.57071e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nor4_lp.pxi.spice"
*
.ends
*
*
