* NGSPICE file created from sky130_fd_sc_lp__o32ai_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o32ai_m A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_179_535# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_179_535# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=4.62e+11p ps=3.88e+06u
M1002 VPWR A1 a_431_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1003 a_66_82# A2 VGND VNB nshort w=420000u l=150000u
+  ad=3.801e+11p pd=4.33e+06u as=2.457e+11p ps=2.85e+06u
M1004 VGND A1 a_66_82# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_431_535# A2 a_337_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1006 VGND A3 a_66_82# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_66_82# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1008 a_337_535# A3 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_66_82# B2 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

