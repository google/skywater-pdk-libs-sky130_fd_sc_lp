* File: sky130_fd_sc_lp__and2b_4.pex.spice
* Created: Fri Aug 28 10:05:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2B_4%A_N 3 7 8 9 10 15 17
c29 15 0 1.21325e-19 $X=0.69 $Y=1.375
c30 8 0 1.37293e-20 $X=0.72 $Y=1.295
r31 15 18 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.667 $Y=1.375
+ $X2=0.667 $Y2=1.54
r32 15 17 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.667 $Y=1.375
+ $X2=0.667 $Y2=1.21
r33 9 10 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.742 $Y=1.665
+ $X2=0.742 $Y2=2.035
r34 8 9 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.742 $Y=1.295
+ $X2=0.742 $Y2=1.665
r35 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.375 $X2=0.69 $Y2=1.375
r36 7 17 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.615 $Y=0.875
+ $X2=0.615 $Y2=1.21
r37 3 18 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.555 $Y=2.045
+ $X2=0.555 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_4%A_213_23# 1 2 9 13 17 21 25 29 33 37 39 48
+ 50 51 52 53 55 59 61 68
c114 50 0 5.24654e-20 $X=2.57 $Y=1.93
c115 37 0 1.53355e-19 $X=2.43 $Y=2.465
c116 17 0 1.37293e-20 $X=1.57 $Y=0.665
r117 62 64 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.14 $Y=1.51
+ $X2=1.57 $Y2=1.51
r118 57 59 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=3.58 $Y=0.995
+ $X2=3.58 $Y2=0.39
r119 53 55 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.66 $Y=2.095
+ $X2=3.15 $Y2=2.095
r120 51 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.415 $Y=1.08
+ $X2=3.58 $Y2=0.995
r121 51 52 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.415 $Y=1.08
+ $X2=2.66 $Y2=1.08
r122 50 53 7.61292 $w=3.3e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.57 $Y=1.93
+ $X2=2.66 $Y2=2.095
r123 49 61 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=2.57 $Y=1.645
+ $X2=2.57 $Y2=1.53
r124 49 50 17.5606 $w=1.78e-07 $l=2.85e-07 $layer=LI1_cond $X=2.57 $Y=1.645
+ $X2=2.57 $Y2=1.93
r125 48 61 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=2.57 $Y=1.415
+ $X2=2.57 $Y2=1.53
r126 47 52 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.57 $Y=1.165
+ $X2=2.66 $Y2=1.08
r127 47 48 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=2.57 $Y=1.165
+ $X2=2.57 $Y2=1.415
r128 46 68 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.34 $Y=1.51 $X2=2.43
+ $Y2=1.51
r129 46 66 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.34 $Y=1.51 $X2=2
+ $Y2=1.51
r130 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.34
+ $Y=1.51 $X2=2.34 $Y2=1.51
r131 42 66 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.66 $Y=1.51 $X2=2
+ $Y2=1.51
r132 42 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.66 $Y=1.51 $X2=1.57
+ $Y2=1.51
r133 41 45 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.66 $Y=1.53
+ $X2=2.34 $Y2=1.53
r134 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.51 $X2=1.66 $Y2=1.51
r135 39 61 0.47666 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=2.48 $Y=1.53 $X2=2.57
+ $Y2=1.53
r136 39 45 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.48 $Y=1.53
+ $X2=2.34 $Y2=1.53
r137 35 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.675
+ $X2=2.43 $Y2=1.51
r138 35 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.43 $Y=1.675
+ $X2=2.43 $Y2=2.465
r139 31 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.345
+ $X2=2.43 $Y2=1.51
r140 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.43 $Y=1.345
+ $X2=2.43 $Y2=0.665
r141 27 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.675 $X2=2
+ $Y2=1.51
r142 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2 $Y=1.675 $X2=2
+ $Y2=2.465
r143 23 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.345 $X2=2
+ $Y2=1.51
r144 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2 $Y=1.345 $X2=2
+ $Y2=0.665
r145 19 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.675
+ $X2=1.57 $Y2=1.51
r146 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.57 $Y=1.675
+ $X2=1.57 $Y2=2.465
r147 15 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.345
+ $X2=1.57 $Y2=1.51
r148 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.57 $Y=1.345
+ $X2=1.57 $Y2=0.665
r149 11 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.675
+ $X2=1.14 $Y2=1.51
r150 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.14 $Y=1.675
+ $X2=1.14 $Y2=2.465
r151 7 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.345
+ $X2=1.14 $Y2=1.51
r152 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.14 $Y=1.345
+ $X2=1.14 $Y2=0.665
r153 2 55 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.835 $X2=3.15 $Y2=2.095
r154 1 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.44
+ $Y=0.245 $X2=3.58 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_4%B 3 7 9 12
c40 12 0 1.9916e-19 $X=2.915 $Y=1.51
r41 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.51
+ $X2=2.915 $Y2=1.675
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.51
+ $X2=2.915 $Y2=1.345
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.51 $X2=2.915 $Y2=1.51
r44 9 13 5.69279 $w=4.13e-07 $l=2.05e-07 $layer=LI1_cond $X=3.12 $Y=1.552
+ $X2=2.915 $Y2=1.552
r45 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.005 $Y=0.665
+ $X2=3.005 $Y2=1.345
r46 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.935 $Y=2.465
+ $X2=2.935 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_4%A_43_367# 1 2 9 13 18 19 20 22 26 29 30
c68 29 0 1.39705e-19 $X=3.55 $Y=1.46
c69 22 0 5.94552e-20 $X=3.63 $Y=2.43
r70 30 33 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.55 $Y=1.46
+ $X2=3.365 $Y2=1.46
r71 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.46 $X2=3.55 $Y2=1.46
r72 23 26 3.84148 $w=2.98e-07 $l=1e-07 $layer=LI1_cond $X=0.3 $Y=0.87 $X2=0.4
+ $Y2=0.87
r73 21 29 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.63 $Y=1.545
+ $X2=3.55 $Y2=1.46
r74 21 22 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.63 $Y=1.545
+ $X2=3.63 $Y2=2.43
r75 19 22 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.545 $Y=2.52
+ $X2=3.63 $Y2=2.43
r76 19 20 192.242 $w=1.78e-07 $l=3.12e-06 $layer=LI1_cond $X=3.545 $Y=2.52
+ $X2=0.425 $Y2=2.52
r77 16 20 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=0.3 $Y=2.43
+ $X2=0.425 $Y2=2.52
r78 16 18 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.3 $Y=2.43 $X2=0.3
+ $Y2=2.11
r79 15 23 1.80669 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=0.3 $Y=1.02 $X2=0.3
+ $Y2=0.87
r80 15 18 50.2465 $w=2.48e-07 $l=1.09e-06 $layer=LI1_cond $X=0.3 $Y=1.02 $X2=0.3
+ $Y2=2.11
r81 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.625
+ $X2=3.365 $Y2=1.46
r82 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.365 $Y=1.625
+ $X2=3.365 $Y2=2.465
r83 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.295
+ $X2=3.365 $Y2=1.46
r84 7 9 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.365 $Y=1.295
+ $X2=3.365 $Y2=0.665
r85 2 18 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.11
r86 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.665 $X2=0.4 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_4%VPWR 1 2 3 4 15 17 21 25 27 29 31 32 33 39
+ 44 50 53 57
r60 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r61 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 48 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 48 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 45 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.68 $Y2=3.33
r67 45 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 44 56 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.627 $Y2=3.33
r69 44 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 40 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=3.33
+ $X2=1.785 $Y2=3.33
r73 40 42 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.95 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 39 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.68 $Y2=3.33
r75 39 42 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 37 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 33 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r79 33 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r80 31 36 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=3.33 $X2=0.72
+ $Y2=3.33
r81 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=3.33
+ $X2=0.925 $Y2=3.33
r82 27 56 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.627 $Y2=3.33
r83 27 29 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=2.915
r84 23 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=3.33
r85 23 25 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=2.915
r86 19 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=3.245
+ $X2=1.785 $Y2=3.33
r87 19 21 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.785 $Y=3.245
+ $X2=1.785 $Y2=2.915
r88 18 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.925 $Y2=3.33
r89 17 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=3.33
+ $X2=1.785 $Y2=3.33
r90 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.62 $Y=3.33
+ $X2=1.09 $Y2=3.33
r91 13 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=3.33
r92 13 15 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=2.915
r93 4 29 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=2.915
r94 3 25 600 $w=1.7e-07 $l=1.16422e-06 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.835 $X2=2.68 $Y2=2.915
r95 2 21 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.835 $X2=1.785 $Y2=2.915
r96 1 15 600 $w=1.7e-07 $l=1.21861e-06 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.925 $Y2=2.915
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_4%X 1 2 3 4 14 17 19 20 23 28 29 30
c46 30 0 1.53355e-19 $X=2.16 $Y=2.035
c47 20 0 1.21325e-19 $X=1.45 $Y=1.16
r48 29 30 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.98
+ $X2=2.16 $Y2=1.98
r49 29 37 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.68 $Y=1.98
+ $X2=1.355 $Y2=1.98
r50 28 37 3.0582 $w=4.98e-07 $l=7e-08 $layer=LI1_cond $X=1.285 $Y=1.98 $X2=1.355
+ $Y2=1.98
r51 21 23 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.215 $Y=1.075
+ $X2=2.215 $Y2=0.42
r52 19 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.12 $Y=1.16
+ $X2=2.215 $Y2=1.075
r53 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.12 $Y=1.16
+ $X2=1.45 $Y2=1.16
r54 15 20 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.34 $Y=1.16
+ $X2=1.45 $Y2=1.16
r55 15 17 34.3114 $w=2.18e-07 $l=6.55e-07 $layer=LI1_cond $X=1.34 $Y=1.075
+ $X2=1.34 $Y2=0.42
r56 14 28 4.12218 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=1.167 $Y=1.815
+ $X2=1.167 $Y2=1.98
r57 13 15 11.2866 $w=1.68e-07 $l=1.73e-07 $layer=LI1_cond $X=1.167 $Y=1.16
+ $X2=1.34 $Y2=1.16
r58 13 14 27.9529 $w=2.33e-07 $l=5.7e-07 $layer=LI1_cond $X=1.167 $Y=1.245
+ $X2=1.167 $Y2=1.815
r59 4 30 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.075
+ $Y=1.835 $X2=2.215 $Y2=1.98
r60 3 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.835 $X2=1.355 $Y2=1.98
r61 2 23 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.075
+ $Y=0.245 $X2=2.215 $Y2=0.42
r62 1 17 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.215
+ $Y=0.245 $X2=1.355 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_4%VGND 1 2 3 12 14 18 22 24 25 26 32 39 40 43
+ 46
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r55 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 40 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r57 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 37 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.715
+ $Y2=0
r59 37 39 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r60 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r61 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 33 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=1.785
+ $Y2=0
r63 33 35 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=2.16
+ $Y2=0
r64 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.715
+ $Y2=0
r65 32 35 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.16
+ $Y2=0
r66 30 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r67 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r68 26 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r69 26 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r70 24 29 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.72
+ $Y2=0
r71 24 25 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.91
+ $Y2=0
r72 20 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0
r73 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0.37
r74 16 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0
r75 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0.39
r76 15 25 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.91
+ $Y2=0
r77 14 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.785
+ $Y2=0
r78 14 15 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.06
+ $Y2=0
r79 10 25 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=0.085 $X2=0.91
+ $Y2=0
r80 10 12 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=0.91 $Y=0.085
+ $X2=0.91 $Y2=0.39
r81 3 22 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=2.505
+ $Y=0.245 $X2=2.715 $Y2=0.37
r82 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.645
+ $Y=0.245 $X2=1.785 $Y2=0.39
r83 1 12 91 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=2 $X=0.69
+ $Y=0.665 $X2=0.925 $Y2=0.39
.ends

