* File: sky130_fd_sc_lp__o2111a_2.spice
* Created: Fri Aug 28 11:00:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111a_2.pex.spice"
.subckt sky130_fd_sc_lp__o2111a_2  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_80_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1005_d N_A_80_21#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 A_386_51# N_D1_M1001_g N_A_80_21#_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1002 A_458_51# N_C1_M1002_g A_386_51# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75000.6 SB=75001.8
+ A=0.126 P=1.98 MULT=1
MM1006 N_A_566_51#_M1006_d N_B1_M1006_g A_458_51# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=8.568 NRS=19.992 M=1 R=5.6 SA=75001.1
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_566_51#_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=5.712 NRS=7.14 M=1 R=5.6 SA=75001.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1011 N_A_566_51#_M1011_d N_A1_M1011_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_80_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A_80_21#_M1012_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4599 AS=0.1764 PD=1.99 PS=1.54 NRD=1.5563 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1003 N_A_80_21#_M1003_d N_D1_M1003_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4599 PD=1.54 PS=1.99 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_C1_M1013_g N_A_80_21#_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1764 PD=1.65 PS=1.54 NRD=9.3772 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1004 N_A_80_21#_M1004_d N_B1_M1004_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=9.3772 NRS=7.8012 M=1 R=8.4 SA=75002.5
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1010 A_674_367# N_A2_M1010_g N_A_80_21#_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75003
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_674_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75003.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o2111a_2.pxi.spice"
*
.ends
*
*
