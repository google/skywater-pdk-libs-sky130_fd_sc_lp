* File: sky130_fd_sc_lp__dlxtn_1.pex.spice
* Created: Wed Sep  2 09:48:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXTN_1%D 3 6 8 9 10 15 17
r33 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.34
+ $X2=0.585 $Y2=1.505
r34 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.34
+ $X2=0.585 $Y2=1.175
r35 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.34 $X2=0.585 $Y2=1.34
r36 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.34 $X2=1.68
+ $Y2=1.34
r37 8 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.34 $X2=1.2
+ $Y2=1.34
r38 8 16 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.34
+ $X2=0.585 $Y2=1.34
r39 6 18 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=0.635 $Y=2.725
+ $X2=0.635 $Y2=1.505
r40 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.635 $Y=0.855
+ $X2=0.635 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%GATE_N 1 3 6 8 11 12 13 14 15 20
r46 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=0.38
+ $X2=1.68 $Y2=0.545
r47 14 15 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.467
+ $X2=2.16 $Y2=0.467
r48 14 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=0.38 $X2=1.68 $Y2=0.38
r49 13 14 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.467 $X2=1.68
+ $Y2=0.467
r50 11 23 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.59 $Y=1.175
+ $X2=1.59 $Y2=0.545
r51 9 12 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.14 $Y=1.25
+ $X2=1.065 $Y2=1.25
r52 8 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.515 $Y=1.25
+ $X2=1.59 $Y2=1.175
r53 8 9 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.515 $Y=1.25
+ $X2=1.14 $Y2=1.25
r54 4 12 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.065 $Y=1.325
+ $X2=1.065 $Y2=1.25
r55 4 6 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=1.065 $Y=1.325
+ $X2=1.065 $Y2=2.725
r56 1 12 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.065 $Y=1.175
+ $X2=1.065 $Y2=1.25
r57 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.065 $Y=1.175
+ $X2=1.065 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%A_228_129# 1 2 9 11 12 15 19 23 27 28 34 36
+ 37 41 42 43 49 50 51 54 55 58 59 60
c148 49 0 1.38845e-19 $X=3.835 $Y=2.06
r149 58 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.08
+ $X2=3.655 $Y2=0.915
r150 57 60 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=3.655 $Y=1.12
+ $X2=3.795 $Y2=1.12
r151 57 59 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=1.12
+ $X2=3.49 $Y2=1.12
r152 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=1.08 $X2=3.655 $Y2=1.08
r153 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.11
+ $Y=1.08 $X2=2.11 $Y2=1.08
r154 51 54 6.04159 $w=3.28e-07 $l=1.73e-07 $layer=LI1_cond $X=2.11 $Y=0.907
+ $X2=2.11 $Y2=1.08
r155 50 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=2.06
+ $X2=3.835 $Y2=2.225
r156 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.835
+ $Y=2.06 $X2=3.835 $Y2=2.06
r157 47 49 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=3.795 $Y=2.375
+ $X2=3.795 $Y2=2.06
r158 46 60 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.795 $Y=1.245
+ $X2=3.795 $Y2=1.12
r159 46 49 37.5696 $w=2.48e-07 $l=8.15e-07 $layer=LI1_cond $X=3.795 $Y=1.245
+ $X2=3.795 $Y2=2.06
r160 45 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=1.08
+ $X2=2.11 $Y2=1.08
r161 45 59 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.275 $Y=1.08
+ $X2=3.49 $Y2=1.08
r162 42 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.67 $Y=2.46
+ $X2=3.795 $Y2=2.375
r163 42 43 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.67 $Y=2.46
+ $X2=2.27 $Y2=2.46
r164 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=2.545
+ $X2=2.27 $Y2=2.46
r165 40 41 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.185 $Y=2.545
+ $X2=2.185 $Y2=2.905
r166 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.1 $Y=2.99
+ $X2=2.185 $Y2=2.905
r167 36 37 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.1 $Y=2.99
+ $X2=1.445 $Y2=2.99
r168 32 37 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.297 $Y=2.905
+ $X2=1.445 $Y2=2.99
r169 32 34 13.8684 $w=2.93e-07 $l=3.55e-07 $layer=LI1_cond $X=1.297 $Y=2.905
+ $X2=1.297 $Y2=2.55
r170 28 51 3.83364 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0.907
+ $X2=2.11 $Y2=0.907
r171 28 30 37.8228 $w=1.93e-07 $l=6.65e-07 $layer=LI1_cond $X=1.945 $Y=0.907
+ $X2=1.28 $Y2=0.907
r172 26 55 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.11 $Y=1.42
+ $X2=2.11 $Y2=1.08
r173 26 27 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.42
+ $X2=2.11 $Y2=1.585
r174 25 55 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=2.11 $Y=0.935
+ $X2=2.11 $Y2=1.08
r175 23 68 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.745 $Y=2.615
+ $X2=3.745 $Y2=2.225
r176 19 64 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.565 $Y=0.445
+ $X2=3.565 $Y2=0.915
r177 13 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.775 $Y=0.785
+ $X2=2.775 $Y2=0.445
r178 12 25 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.275 $Y=0.86
+ $X2=2.11 $Y2=0.935
r179 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.7 $Y=0.86
+ $X2=2.775 $Y2=0.785
r180 11 12 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.7 $Y=0.86
+ $X2=2.275 $Y2=0.86
r181 9 27 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.05 $Y=2.725
+ $X2=2.05 $Y2=1.585
r182 2 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=2.405 $X2=1.28 $Y2=2.55
r183 1 30 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.645 $X2=1.28 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%A_59_129# 1 2 9 11 12 15 19 21 24 26 30 31
+ 36 38
c83 12 0 6.65831e-20 $X=2.92 $Y=1.22
r84 33 36 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.24 $Y=0.84
+ $X2=0.42 $Y2=0.84
r85 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.725
+ $Y=1.43 $X2=2.725 $Y2=1.43
r86 28 30 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.725 $Y=1.675
+ $X2=2.725 $Y2=1.43
r87 27 38 2.90107 $w=1.9e-07 $l=2e-07 $layer=LI1_cond $X=0.55 $Y=1.77 $X2=0.35
+ $Y2=1.77
r88 26 28 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=2.56 $Y=1.77
+ $X2=2.725 $Y2=1.675
r89 26 27 117.33 $w=1.88e-07 $l=2.01e-06 $layer=LI1_cond $X=2.56 $Y=1.77
+ $X2=0.55 $Y2=1.77
r90 22 38 3.58697 $w=2.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.35 $Y=1.865
+ $X2=0.35 $Y2=1.77
r91 22 24 19.7356 $w=3.98e-07 $l=6.85e-07 $layer=LI1_cond $X=0.35 $Y=1.865
+ $X2=0.35 $Y2=2.55
r92 21 38 3.58697 $w=2.9e-07 $l=1.50167e-07 $layer=LI1_cond $X=0.24 $Y=1.675
+ $X2=0.35 $Y2=1.77
r93 20 33 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.005
+ $X2=0.24 $Y2=0.84
r94 20 21 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=0.24 $Y=1.005
+ $X2=0.24 $Y2=1.675
r95 18 31 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=2.74 $Y=1.755
+ $X2=2.74 $Y2=1.43
r96 18 19 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=2.74 $Y=1.755
+ $X2=2.74 $Y2=1.935
r97 17 31 21.6391 $w=3.6e-07 $l=1.35e-07 $layer=POLY_cond $X=2.74 $Y=1.295
+ $X2=2.74 $Y2=1.43
r98 13 15 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=3.205 $Y=1.145
+ $X2=3.205 $Y2=0.445
r99 12 17 33.3473 $w=1.5e-07 $l=2.14243e-07 $layer=POLY_cond $X=2.92 $Y=1.22
+ $X2=2.74 $Y2=1.295
r100 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.13 $Y=1.22
+ $X2=3.205 $Y2=1.145
r101 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.13 $Y=1.22
+ $X2=2.92 $Y2=1.22
r102 9 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.845 $Y=2.725
+ $X2=2.845 $Y2=1.935
r103 2 24 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.295
+ $Y=2.405 $X2=0.42 $Y2=2.55
r104 1 36 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.295
+ $Y=0.645 $X2=0.42 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%A_342_481# 1 2 9 11 12 15 18 20 21 25 27 28
+ 31 33 34 37 38 42 43
c111 42 0 5.37319e-20 $X=4.195 $Y=0.93
c112 34 0 6.65831e-20 $X=2.645 $Y=0.74
r113 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.195
+ $Y=0.93 $X2=4.195 $Y2=0.93
r114 40 42 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=4.19 $Y=0.825
+ $X2=4.19 $Y2=0.93
r115 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.295
+ $Y=1.7 $X2=3.295 $Y2=1.7
r116 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.295 $Y=2.035
+ $X2=3.295 $Y2=1.7
r117 33 40 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.09 $Y=0.74
+ $X2=4.19 $Y2=0.825
r118 33 34 94.2727 $w=1.68e-07 $l=1.445e-06 $layer=LI1_cond $X=4.09 $Y=0.74
+ $X2=2.645 $Y2=0.74
r119 29 34 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.55 $Y=0.655
+ $X2=2.645 $Y2=0.74
r120 29 31 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.55 $Y=0.655
+ $X2=2.55 $Y2=0.46
r121 27 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.13 $Y=2.12
+ $X2=3.295 $Y2=2.035
r122 27 28 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=3.13 $Y=2.12
+ $X2=1.93 $Y2=2.12
r123 23 28 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.83 $Y=2.205
+ $X2=1.93 $Y2=2.12
r124 23 25 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.83 $Y=2.205
+ $X2=1.83 $Y2=2.57
r125 21 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.195 $Y=1.27
+ $X2=4.195 $Y2=0.93
r126 21 22 54.9356 $w=3.3e-07 $l=3.47419e-07 $layer=POLY_cond $X=4.195 $Y=1.27
+ $X2=4.18 $Y2=1.61
r127 20 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=0.765
+ $X2=4.195 $Y2=0.93
r128 17 38 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.295 $Y=2.04
+ $X2=3.295 $Y2=1.7
r129 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=2.04
+ $X2=3.295 $Y2=2.205
r130 16 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.295 $Y=1.685
+ $X2=3.295 $Y2=1.7
r131 15 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.105 $Y=0.445
+ $X2=4.105 $Y2=0.765
r132 12 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.46 $Y=1.61
+ $X2=3.295 $Y2=1.685
r133 11 22 11.8763 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.03 $Y=1.61
+ $X2=4.18 $Y2=1.61
r134 11 12 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.03 $Y=1.61
+ $X2=3.46 $Y2=1.61
r135 9 18 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.205 $Y=2.725
+ $X2=3.205 $Y2=2.205
r136 2 25 600 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.405 $X2=1.835 $Y2=2.57
r137 1 31 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.235 $X2=2.56 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%A_842_413# 1 2 9 13 17 20 22 26 30 33 37 40
+ 41 45 47 48 49 50 55
c95 45 0 1.92577e-19 $X=4.615 $Y=2.05
r96 45 53 5.69291 $w=2.54e-07 $l=3e-08 $layer=POLY_cond $X=4.615 $Y=2.05
+ $X2=4.645 $Y2=2.05
r97 44 47 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=2.085
+ $X2=4.78 $Y2=2.085
r98 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.615
+ $Y=2.05 $X2=4.615 $Y2=2.05
r99 41 56 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=6.122 $Y=1.42
+ $X2=6.122 $Y2=1.585
r100 41 55 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=6.122 $Y=1.42
+ $X2=6.122 $Y2=1.255
r101 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.09
+ $Y=1.42 $X2=6.09 $Y2=1.42
r102 38 50 0.067832 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=5.66 $Y=1.42
+ $X2=5.525 $Y2=1.42
r103 38 40 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.66 $Y=1.42
+ $X2=6.09 $Y2=1.42
r104 35 49 3.29812 $w=2.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=5.525 $Y=1.965
+ $X2=5.51 $Y2=2.05
r105 35 37 3.20123 $w=2.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.525 $Y=1.965
+ $X2=5.525 $Y2=1.89
r106 34 50 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.525 $Y=1.585
+ $X2=5.525 $Y2=1.42
r107 34 37 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.525 $Y=1.585
+ $X2=5.525 $Y2=1.89
r108 33 50 7.13466 $w=2.2e-07 $l=1.88348e-07 $layer=LI1_cond $X=5.475 $Y=1.255
+ $X2=5.525 $Y2=1.42
r109 33 48 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.475 $Y=1.255
+ $X2=5.475 $Y2=1.075
r110 28 49 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=2.135
+ $X2=5.51 $Y2=2.05
r111 28 30 9.41162 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=5.51 $Y=2.135
+ $X2=5.51 $Y2=2.38
r112 24 48 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=5.42 $Y=0.935
+ $X2=5.42 $Y2=1.075
r113 24 26 21.1967 $w=2.78e-07 $l=5.15e-07 $layer=LI1_cond $X=5.42 $Y=0.935
+ $X2=5.42 $Y2=0.42
r114 22 49 3.25423 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.36 $Y=2.05
+ $X2=5.51 $Y2=2.05
r115 22 47 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=5.36 $Y=2.05
+ $X2=4.78 $Y2=2.05
r116 20 56 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=6.245 $Y=2.465
+ $X2=6.245 $Y2=1.585
r117 17 55 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.245 $Y=0.725
+ $X2=6.245 $Y2=1.255
r118 11 53 15.087 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.645 $Y=1.885
+ $X2=4.645 $Y2=2.05
r119 11 13 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=4.645 $Y=1.885
+ $X2=4.645 $Y2=0.445
r120 7 45 62.622 $w=2.54e-07 $l=4.04166e-07 $layer=POLY_cond $X=4.285 $Y=2.215
+ $X2=4.615 $Y2=2.05
r121 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.285 $Y=2.215
+ $X2=4.285 $Y2=2.615
r122 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.745 $X2=5.495 $Y2=1.89
r123 2 30 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.745 $X2=5.495 $Y2=2.38
r124 1 26 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.245
+ $Y=0.235 $X2=5.385 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%A_656_481# 1 2 9 13 15 19 24 25 26 28 31 32
+ 34
r98 32 37 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.157 $Y=1.42
+ $X2=5.157 $Y2=1.585
r99 32 36 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.157 $Y=1.42
+ $X2=5.157 $Y2=1.255
r100 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.125
+ $Y=1.42 $X2=5.125 $Y2=1.42
r101 29 34 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=1.52
+ $X2=4.545 $Y2=1.52
r102 29 31 11.1709 $w=5.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.63 $Y=1.52
+ $X2=5.125 $Y2=1.52
r103 28 34 4.03347 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=4.545 $Y=1.255
+ $X2=4.545 $Y2=1.52
r104 27 28 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.545 $Y=0.465
+ $X2=4.545 $Y2=1.255
r105 25 34 2.73602 $w=3.5e-07 $l=2.18403e-07 $layer=LI1_cond $X=4.46 $Y=1.7
+ $X2=4.545 $Y2=1.52
r106 25 26 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.46 $Y=1.7
+ $X2=4.28 $Y2=1.7
r107 23 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.185 $Y=1.785
+ $X2=4.28 $Y2=1.7
r108 23 24 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.185 $Y=1.785
+ $X2=4.185 $Y2=2.715
r109 19 27 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.46 $Y=0.37
+ $X2=4.545 $Y2=0.465
r110 19 21 33.2727 $w=1.88e-07 $l=5.7e-07 $layer=LI1_cond $X=4.46 $Y=0.37
+ $X2=3.89 $Y2=0.37
r111 15 24 7.62524 $w=3.5e-07 $l=2.17371e-07 $layer=LI1_cond $X=4.09 $Y=2.89
+ $X2=4.185 $Y2=2.715
r112 15 17 22.0611 $w=3.48e-07 $l=6.7e-07 $layer=LI1_cond $X=4.09 $Y=2.89
+ $X2=3.42 $Y2=2.89
r113 13 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.28 $Y=2.375
+ $X2=5.28 $Y2=1.585
r114 9 36 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.17 $Y=0.655 $X2=5.17
+ $Y2=1.255
r115 2 17 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=2.405 $X2=3.42 $Y2=2.88
r116 1 21 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.235 $X2=3.89 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%VPWR 1 2 3 4 17 21 25 29 31 39 44 51 52 55
+ 58 65 68
r77 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r78 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 63 65 12.9421 $w=6.74e-07 $l=7.15e-07 $layer=LI1_cond $X=4.82 $Y=2.615
+ $X2=4.82 $Y2=3.33
r80 61 63 1.71958 $w=6.74e-07 $l=9.5e-08 $layer=LI1_cond $X=4.82 $Y=2.52
+ $X2=4.82 $Y2=2.615
r81 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 52 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r84 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r85 49 68 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.02 $Y2=3.33
r86 49 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.48 $Y2=3.33
r87 48 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r88 48 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r89 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 45 65 9.07283 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=5.19 $Y=3.33 $X2=4.82
+ $Y2=3.33
r91 45 47 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.19 $Y=3.33
+ $X2=5.52 $Y2=3.33
r92 44 68 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.865 $Y=3.33
+ $X2=6.02 $Y2=3.33
r93 44 47 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=3.33
+ $X2=5.52 $Y2=3.33
r94 43 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 40 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.7 $Y=3.33 $X2=2.57
+ $Y2=3.33
r97 40 42 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.7 $Y=3.33
+ $X2=4.08 $Y2=3.33
r98 39 65 9.07283 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=4.45 $Y=3.33 $X2=4.82
+ $Y2=3.33
r99 39 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.45 $Y=3.33 $X2=4.08
+ $Y2=3.33
r100 38 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r102 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r105 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r106 32 55 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.85 $Y2=3.33
r107 32 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 31 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.44 $Y=3.33
+ $X2=2.57 $Y2=3.33
r109 31 37 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 29 43 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 29 59 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 25 28 36.0603 $w=3.08e-07 $l=9.7e-07 $layer=LI1_cond $X=6.02 $Y=1.98
+ $X2=6.02 $Y2=2.95
r113 23 68 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=3.245
+ $X2=6.02 $Y2=3.33
r114 23 28 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=6.02 $Y=3.245
+ $X2=6.02 $Y2=2.95
r115 19 58 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=3.245
+ $X2=2.57 $Y2=3.33
r116 19 21 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=2.57 $Y=3.245
+ $X2=2.57 $Y2=2.88
r117 15 55 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=3.33
r118 15 17 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=2.55
r119 4 28 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.835 $X2=6.03 $Y2=2.95
r120 4 25 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.835 $X2=6.03 $Y2=1.98
r121 3 63 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.405 $X2=4.535 $Y2=2.615
r122 3 61 300 $w=1.7e-07 $l=7.60329e-07 $layer=licon1_PDIFF $count=2 $X=4.36
+ $Y=2.405 $X2=5.065 $Y2=2.52
r123 2 21 600 $w=1.7e-07 $l=6.48363e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=2.405 $X2=2.535 $Y2=2.88
r124 1 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.71
+ $Y=2.405 $X2=0.85 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%Q 1 2 7 8 9 10 11 12 13 22
r11 13 40 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=6.49 $Y=2.775
+ $X2=6.49 $Y2=2.91
r12 12 13 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=6.49 $Y=2.405
+ $X2=6.49 $Y2=2.775
r13 11 12 16.8893 $w=2.88e-07 $l=4.25e-07 $layer=LI1_cond $X=6.49 $Y=1.98
+ $X2=6.49 $Y2=2.405
r14 10 11 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=6.49 $Y=1.665
+ $X2=6.49 $Y2=1.98
r15 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=6.49 $Y=1.295
+ $X2=6.49 $Y2=1.665
r16 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=6.49 $Y=0.925 $X2=6.49
+ $Y2=1.295
r17 7 8 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=6.49 $Y=0.555 $X2=6.49
+ $Y2=0.925
r18 7 22 4.17264 $w=2.88e-07 $l=1.05e-07 $layer=LI1_cond $X=6.49 $Y=0.555
+ $X2=6.49 $Y2=0.45
r19 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.91
r20 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=1.98
r21 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.305 $X2=6.46 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_1%VGND 1 2 3 4 17 21 25 31 34 35 36 38 50 56
+ 57 60 63 66
r77 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r78 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r79 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r80 57 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r81 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r82 54 66 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=6.175 $Y=0 $X2=6.02
+ $Y2=0
r83 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.175 $Y=0 $X2=6.48
+ $Y2=0
r84 53 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r85 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r86 50 66 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=6.02
+ $Y2=0
r87 50 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=5.52
+ $Y2=0
r88 49 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r89 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r90 46 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=2.99
+ $Y2=0
r91 46 48 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=3.155 $Y=0
+ $X2=4.56 $Y2=0
r92 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r93 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r94 42 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r95 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r96 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r97 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r98 39 60 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.832
+ $Y2=0
r99 39 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r100 38 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.99
+ $Y2=0
r101 38 44 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=0
+ $X2=2.64 $Y2=0
r102 36 49 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.56
+ $Y2=0
r103 36 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r104 34 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r105 34 35 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.955
+ $Y2=0
r106 33 52 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=5.52
+ $Y2=0
r107 33 35 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=4.955
+ $Y2=0
r108 29 66 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=0.085
+ $X2=6.02 $Y2=0
r109 29 31 13.5691 $w=3.08e-07 $l=3.65e-07 $layer=LI1_cond $X=6.02 $Y=0.085
+ $X2=6.02 $Y2=0.45
r110 25 27 20.0748 $w=3.08e-07 $l=5.4e-07 $layer=LI1_cond $X=4.955 $Y=0.38
+ $X2=4.955 $Y2=0.92
r111 23 35 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.955 $Y=0.085
+ $X2=4.955 $Y2=0
r112 23 25 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.955 $Y=0.085
+ $X2=4.955 $Y2=0.38
r113 19 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0
r114 19 21 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0.385
r115 15 60 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.832 $Y=0.085
+ $X2=0.832 $Y2=0
r116 15 17 38.6709 $w=2.23e-07 $l=7.55e-07 $layer=LI1_cond $X=0.832 $Y=0.085
+ $X2=0.832 $Y2=0.84
r117 4 31 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.905
+ $Y=0.305 $X2=6.03 $Y2=0.45
r118 3 27 182 $w=1.7e-07 $l=7.93851e-07 $layer=licon1_NDIFF $count=1 $X=4.72
+ $Y=0.235 $X2=4.955 $Y2=0.92
r119 3 25 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=4.72
+ $Y=0.235 $X2=4.925 $Y2=0.38
r120 2 21 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.235 $X2=2.99 $Y2=0.385
r121 1 17 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.71
+ $Y=0.645 $X2=0.85 $Y2=0.84
.ends

