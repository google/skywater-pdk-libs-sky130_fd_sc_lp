* File: sky130_fd_sc_lp__maj3_4.pxi.spice
* Created: Wed Sep  2 09:59:38 2020
* 
x_PM_SKY130_FD_SC_LP__MAJ3_4%C N_C_M1002_g N_C_M1014_g N_C_M1016_g N_C_M1019_g
+ N_C_c_97_n N_C_c_112_p N_C_c_133_p N_C_c_98_n N_C_c_99_n N_C_c_100_n C
+ N_C_c_101_n N_C_c_102_n N_C_c_103_n PM_SKY130_FD_SC_LP__MAJ3_4%C
x_PM_SKY130_FD_SC_LP__MAJ3_4%A N_A_c_183_n N_A_M1001_g N_A_M1000_g N_A_c_185_n
+ N_A_M1010_g N_A_M1008_g A A N_A_c_188_n PM_SKY130_FD_SC_LP__MAJ3_4%A
x_PM_SKY130_FD_SC_LP__MAJ3_4%B N_B_c_228_n N_B_M1011_g N_B_M1018_g N_B_c_230_n
+ N_B_M1017_g N_B_M1009_g B N_B_c_233_n PM_SKY130_FD_SC_LP__MAJ3_4%B
x_PM_SKY130_FD_SC_LP__MAJ3_4%A_65_367# N_A_65_367#_M1002_s N_A_65_367#_M1011_d
+ N_A_65_367#_M1014_s N_A_65_367#_M1018_d N_A_65_367#_M1006_g
+ N_A_65_367#_M1003_g N_A_65_367#_M1007_g N_A_65_367#_M1004_g
+ N_A_65_367#_M1005_g N_A_65_367#_M1013_g N_A_65_367#_M1012_g
+ N_A_65_367#_M1015_g N_A_65_367#_c_291_n N_A_65_367#_c_280_n
+ N_A_65_367#_c_303_n N_A_65_367#_c_281_n N_A_65_367#_c_282_n
+ N_A_65_367#_c_293_n N_A_65_367#_c_294_n N_A_65_367#_c_310_n
+ N_A_65_367#_c_311_n N_A_65_367#_c_346_n N_A_65_367#_c_283_n
+ N_A_65_367#_c_284_n N_A_65_367#_c_373_p N_A_65_367#_c_295_n
+ N_A_65_367#_c_285_n N_A_65_367#_c_286_n PM_SKY130_FD_SC_LP__MAJ3_4%A_65_367#
x_PM_SKY130_FD_SC_LP__MAJ3_4%VPWR N_VPWR_M1000_d N_VPWR_M1019_d N_VPWR_M1007_d
+ N_VPWR_M1015_d N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n
+ N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n VPWR N_VPWR_c_449_n
+ N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_441_n
+ PM_SKY130_FD_SC_LP__MAJ3_4%VPWR
x_PM_SKY130_FD_SC_LP__MAJ3_4%X N_X_M1003_s N_X_M1005_s N_X_M1006_s N_X_M1013_s
+ N_X_c_524_n N_X_c_575_p N_X_c_519_n N_X_c_520_n N_X_c_514_n N_X_c_515_n
+ N_X_c_542_n N_X_c_544_n N_X_c_516_n N_X_c_521_n N_X_c_517_n N_X_c_522_n X X
+ PM_SKY130_FD_SC_LP__MAJ3_4%X
x_PM_SKY130_FD_SC_LP__MAJ3_4%VGND N_VGND_M1001_d N_VGND_M1016_d N_VGND_M1004_d
+ N_VGND_M1012_d N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n N_VGND_c_586_n
+ N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n
+ VGND N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n
+ PM_SKY130_FD_SC_LP__MAJ3_4%VGND
cc_1 VNB N_C_M1014_g 0.00736866f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_2 VNB N_C_M1016_g 0.0230824f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.655
cc_3 VNB N_C_M1019_g 0.00252884f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=2.465
cc_4 VNB N_C_c_97_n 0.00121704f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.225
cc_5 VNB N_C_c_98_n 9.25047e-19 $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=2.225
cc_6 VNB N_C_c_99_n 0.00677702f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.44
cc_7 VNB N_C_c_100_n 0.0291856f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.44
cc_8 VNB N_C_c_101_n 0.0362553f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_9 VNB N_C_c_102_n 0.0194471f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.185
cc_10 VNB N_C_c_103_n 0.00851341f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.347
cc_11 VNB N_A_c_183_n 0.0157298f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.185
cc_12 VNB N_A_M1000_g 0.0064729f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_13 VNB N_A_c_185_n 0.0156895f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.275
cc_14 VNB N_A_M1008_g 0.00700511f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=2.465
cc_15 VNB A 0.00333002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_c_188_n 0.0379097f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.44
cc_17 VNB N_B_c_228_n 0.0158886f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.185
cc_18 VNB N_B_M1018_g 0.00702754f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_19 VNB N_B_c_230_n 0.0159817f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=1.275
cc_20 VNB N_B_M1009_g 0.00702775f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=2.465
cc_21 VNB B 0.00377015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_233_n 0.0379466f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.44
cc_23 VNB N_A_65_367#_M1006_g 0.00281093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_65_367#_M1003_g 0.0223219f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.31
cc_25 VNB N_A_65_367#_M1007_g 0.00278413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_65_367#_M1004_g 0.0208293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_65_367#_M1005_g 0.0215603f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_28 VNB N_A_65_367#_M1013_g 0.00278265f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.44
cc_29 VNB N_A_65_367#_M1012_g 0.0247544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_65_367#_M1015_g 0.00269456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_65_367#_c_280_n 0.0216484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_65_367#_c_281_n 0.0153683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_65_367#_c_282_n 0.0107904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_65_367#_c_283_n 0.00224257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_65_367#_c_284_n 0.00449861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_65_367#_c_285_n 0.0324612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_65_367#_c_286_n 0.0915677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_441_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_514_n 0.00302036f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.44
cc_40 VNB N_X_c_515_n 0.00144547f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.44
cc_41 VNB N_X_c_516_n 0.0108933f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.605
cc_42 VNB N_X_c_517_n 0.00245859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB X 0.0284213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_583_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_584_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.31
cc_46 VNB N_VGND_c_585_n 0.00240024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_586_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.44
cc_48 VNB N_VGND_c_587_n 0.0252127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_588_n 0.0366759f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_50 VNB N_VGND_c_589_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_51 VNB N_VGND_c_590_n 0.0213653f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.185
cc_52 VNB N_VGND_c_591_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.515
cc_53 VNB N_VGND_c_592_n 0.0341884f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=1.605
cc_54 VNB N_VGND_c_593_n 0.0199813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_594_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_595_n 0.271395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VPB N_C_M1014_g 0.0225079f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_58 VPB N_C_M1019_g 0.0204327f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.465
cc_59 VPB N_C_c_97_n 0.00125361f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.225
cc_60 VPB N_C_c_98_n 0.00152602f $X=-0.19 $Y=1.655 $X2=2.57 $Y2=2.225
cc_61 VPB N_A_M1000_g 0.0189096f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_62 VPB N_A_M1008_g 0.0193877f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.465
cc_63 VPB A 0.00457738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_B_M1018_g 0.0191799f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_65 VPB N_B_M1009_g 0.0194279f $X=-0.19 $Y=1.655 $X2=2.725 $Y2=2.465
cc_66 VPB N_A_65_367#_M1006_g 0.0214239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_65_367#_M1007_g 0.0211414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_65_367#_M1013_g 0.0211375f $X=-0.19 $Y=1.655 $X2=2.815 $Y2=1.44
cc_69 VPB N_A_65_367#_M1015_g 0.0232644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_65_367#_c_291_n 0.0510126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_65_367#_c_282_n 0.0022772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_65_367#_c_293_n 4.42052e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_65_367#_c_294_n 0.00398748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_65_367#_c_295_n 0.0198114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_65_367#_c_285_n 0.00698284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_442_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_443_n 0.0149763f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.31
cc_78 VPB N_VPWR_c_444_n 0.00561774f $X=-0.19 $Y=1.655 $X2=2.815 $Y2=1.44
cc_79 VPB N_VPWR_c_445_n 0.011928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_446_n 0.0403864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_447_n 0.0424857f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.35
cc_82 VPB N_VPWR_c_448_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.185
cc_83 VPB N_VPWR_c_449_n 0.032943f $X=-0.19 $Y=1.655 $X2=2.815 $Y2=1.275
cc_84 VPB N_VPWR_c_450_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_451_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_452_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_453_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_441_n 0.0483354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_X_c_519_n 0.00342708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_X_c_520_n 0.00235119f $X=-0.19 $Y=1.655 $X2=2.815 $Y2=1.44
cc_91 VPB N_X_c_521_n 0.0124084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_X_c_522_n 0.00235119f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.347
cc_93 VPB X 0.00657223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 N_C_c_102_n N_A_c_183_n 0.0543919f $X=0.605 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_95 N_C_c_103_n N_A_c_183_n 0.0026001f $X=0.82 $Y=1.347 $X2=-0.19 $Y2=-0.245
cc_96 N_C_M1014_g N_A_M1000_g 0.0543919f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_97 N_C_c_97_n N_A_M1000_g 0.0113079f $X=0.82 $Y=2.225 $X2=0 $Y2=0
cc_98 N_C_c_112_p N_A_M1000_g 0.0170781f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_99 N_C_c_112_p N_A_M1008_g 0.0186344f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_100 N_C_M1014_g A 2.36504e-19 $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_101 N_C_c_97_n A 0.019039f $X=0.82 $Y=2.225 $X2=0 $Y2=0
cc_102 N_C_c_112_p A 0.011487f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_103 N_C_c_102_n A 2.93484e-19 $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_104 N_C_c_103_n A 0.0260326f $X=0.82 $Y=1.347 $X2=0 $Y2=0
cc_105 N_C_c_101_n N_A_c_188_n 0.0543919f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_106 N_C_c_112_p N_B_M1018_g 0.0148387f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_107 N_C_M1016_g N_B_c_230_n 0.0553222f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_108 N_C_M1019_g N_B_M1009_g 0.0553222f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_109 N_C_c_112_p N_B_M1009_g 0.0186052f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_110 N_C_c_98_n N_B_M1009_g 0.0100792f $X=2.57 $Y=2.225 $X2=0 $Y2=0
cc_111 N_C_M1016_g B 4.90383e-19 $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_112 N_C_c_99_n B 0.0188046f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_113 N_C_c_99_n N_B_c_233_n 0.00450616f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_114 N_C_c_100_n N_B_c_233_n 0.0553222f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_115 N_C_c_112_p N_A_65_367#_M1018_d 0.00814554f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_116 N_C_M1019_g N_A_65_367#_M1006_g 0.0345478f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_117 N_C_c_98_n N_A_65_367#_M1006_g 9.28419e-19 $X=2.57 $Y=2.225 $X2=0 $Y2=0
cc_118 N_C_M1016_g N_A_65_367#_M1003_g 0.0197016f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_119 N_C_c_133_p N_A_65_367#_c_291_n 0.0137433f $X=0.905 $Y=2.31 $X2=0 $Y2=0
cc_120 N_C_c_102_n N_A_65_367#_c_280_n 0.0101532f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_121 N_C_c_102_n N_A_65_367#_c_303_n 0.00837828f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_122 N_C_c_101_n N_A_65_367#_c_281_n 0.00110965f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_123 N_C_c_102_n N_A_65_367#_c_281_n 7.90452e-19 $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_124 N_C_c_103_n N_A_65_367#_c_281_n 0.0298012f $X=0.82 $Y=1.347 $X2=0 $Y2=0
cc_125 N_C_c_112_p N_A_65_367#_c_293_n 0.00982214f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_126 N_C_c_112_p N_A_65_367#_c_294_n 0.0235064f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_127 N_C_c_98_n N_A_65_367#_c_294_n 0.0171906f $X=2.57 $Y=2.225 $X2=0 $Y2=0
cc_128 N_C_M1016_g N_A_65_367#_c_310_n 0.00189708f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_129 N_C_M1016_g N_A_65_367#_c_311_n 0.0129826f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_130 N_C_c_99_n N_A_65_367#_c_311_n 0.0226991f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_131 N_C_c_100_n N_A_65_367#_c_311_n 0.00359534f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_132 N_C_M1016_g N_A_65_367#_c_283_n 0.0049452f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_133 N_C_c_99_n N_A_65_367#_c_284_n 0.0273738f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_134 N_C_c_100_n N_A_65_367#_c_284_n 0.00129212f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_135 N_C_M1014_g N_A_65_367#_c_295_n 0.0151563f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_136 N_C_c_97_n N_A_65_367#_c_295_n 0.0313056f $X=0.82 $Y=2.225 $X2=0 $Y2=0
cc_137 N_C_c_101_n N_A_65_367#_c_295_n 0.00249576f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_138 N_C_c_103_n N_A_65_367#_c_295_n 0.00663736f $X=0.82 $Y=1.347 $X2=0 $Y2=0
cc_139 N_C_M1014_g N_A_65_367#_c_285_n 0.00492468f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_140 N_C_c_97_n N_A_65_367#_c_285_n 0.00925313f $X=0.82 $Y=2.225 $X2=0 $Y2=0
cc_141 N_C_c_101_n N_A_65_367#_c_285_n 0.00229059f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_142 N_C_c_102_n N_A_65_367#_c_285_n 0.00464968f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_143 N_C_c_103_n N_A_65_367#_c_285_n 0.0247443f $X=0.82 $Y=1.347 $X2=0 $Y2=0
cc_144 N_C_c_99_n N_A_65_367#_c_286_n 3.65359e-19 $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_145 N_C_c_100_n N_A_65_367#_c_286_n 0.0182352f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_146 N_C_c_97_n A_154_367# 0.00434959f $X=0.82 $Y=2.225 $X2=-0.19 $Y2=-0.245
cc_147 N_C_c_112_p A_154_367# 0.00358662f $X=2.485 $Y=2.31 $X2=-0.19 $Y2=-0.245
cc_148 N_C_c_133_p A_154_367# 0.00347351f $X=0.905 $Y=2.31 $X2=-0.19 $Y2=-0.245
cc_149 N_C_c_112_p N_VPWR_M1000_d 0.00462185f $X=2.485 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_150 N_C_M1014_g N_VPWR_c_442_n 0.00268359f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_151 N_C_c_112_p N_VPWR_c_442_n 0.0164319f $X=2.485 $Y=2.31 $X2=0 $Y2=0
cc_152 N_C_M1019_g N_VPWR_c_443_n 0.0114176f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_153 N_C_c_98_n N_VPWR_c_443_n 0.0154459f $X=2.57 $Y=2.225 $X2=0 $Y2=0
cc_154 N_C_c_99_n N_VPWR_c_443_n 0.01117f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_155 N_C_c_100_n N_VPWR_c_443_n 0.00332104f $X=2.815 $Y=1.44 $X2=0 $Y2=0
cc_156 N_C_M1019_g N_VPWR_c_447_n 0.00585385f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_157 N_C_M1014_g N_VPWR_c_449_n 0.00585385f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_158 N_C_M1014_g N_VPWR_c_441_n 0.0118766f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_159 N_C_M1019_g N_VPWR_c_441_n 0.0110752f $X=2.725 $Y=2.465 $X2=0 $Y2=0
cc_160 N_C_c_112_p A_318_367# 0.00617953f $X=2.485 $Y=2.31 $X2=-0.19 $Y2=-0.245
cc_161 N_C_c_112_p A_482_367# 0.00612411f $X=2.485 $Y=2.31 $X2=-0.19 $Y2=-0.245
cc_162 N_C_c_98_n A_482_367# 0.00380049f $X=2.57 $Y=2.225 $X2=-0.19 $Y2=-0.245
cc_163 N_C_c_102_n N_VGND_c_583_n 0.00232625f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_164 N_C_M1016_g N_VGND_c_584_n 0.0128416f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_165 N_C_M1016_g N_VGND_c_588_n 0.00486043f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_166 N_C_c_102_n N_VGND_c_592_n 0.00549284f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_167 N_C_M1016_g N_VGND_c_595_n 0.00451716f $X=2.725 $Y=0.655 $X2=0 $Y2=0
cc_168 N_C_c_102_n N_VGND_c_595_n 0.00726776f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A_c_185_n N_B_c_228_n 0.0542833f $X=1.515 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_170 N_A_M1008_g N_B_M1018_g 0.0542833f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A_c_188_n N_B_c_233_n 0.0542833f $X=1.515 $Y=1.35 $X2=0 $Y2=0
cc_172 N_A_c_183_n N_A_65_367#_c_280_n 0.001982f $X=1.085 $Y=1.185 $X2=0 $Y2=0
cc_173 N_A_c_183_n N_A_65_367#_c_303_n 0.0138338f $X=1.085 $Y=1.185 $X2=0 $Y2=0
cc_174 N_A_c_185_n N_A_65_367#_c_303_n 0.0160666f $X=1.515 $Y=1.185 $X2=0 $Y2=0
cc_175 A N_A_65_367#_c_303_n 0.0222952f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A_c_188_n N_A_65_367#_c_303_n 6.86408e-19 $X=1.515 $Y=1.35 $X2=0 $Y2=0
cc_177 N_A_c_185_n N_A_65_367#_c_282_n 0.00796921f $X=1.515 $Y=1.185 $X2=0 $Y2=0
cc_178 A N_A_65_367#_c_282_n 0.039598f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A_M1008_g N_A_65_367#_c_293_n 0.00203125f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_c_185_n N_A_65_367#_c_310_n 0.00189708f $X=1.515 $Y=1.185 $X2=0 $Y2=0
cc_181 N_A_M1000_g N_VPWR_c_442_n 0.0161113f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_M1008_g N_VPWR_c_442_n 0.0159555f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_M1008_g N_VPWR_c_447_n 0.00486043f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_M1000_g N_VPWR_c_449_n 0.00486043f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_M1000_g N_VPWR_c_441_n 0.00827383f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_M1008_g N_VPWR_c_441_n 0.00827383f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_c_183_n N_VGND_c_583_n 0.012389f $X=1.085 $Y=1.185 $X2=0 $Y2=0
cc_188 N_A_c_185_n N_VGND_c_583_n 0.0124226f $X=1.515 $Y=1.185 $X2=0 $Y2=0
cc_189 N_A_c_185_n N_VGND_c_588_n 0.00486043f $X=1.515 $Y=1.185 $X2=0 $Y2=0
cc_190 N_A_c_183_n N_VGND_c_592_n 0.00486043f $X=1.085 $Y=1.185 $X2=0 $Y2=0
cc_191 N_A_c_183_n N_VGND_c_595_n 0.00451716f $X=1.085 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A_c_185_n N_VGND_c_595_n 0.00451716f $X=1.515 $Y=1.185 $X2=0 $Y2=0
cc_193 N_B_c_228_n N_A_65_367#_c_282_n 0.0122107f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_194 B N_A_65_367#_c_282_n 0.0240759f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_195 N_B_M1018_g N_A_65_367#_c_294_n 0.0147315f $X=1.905 $Y=2.465 $X2=0 $Y2=0
cc_196 N_B_M1009_g N_A_65_367#_c_294_n 0.0039139f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_197 B N_A_65_367#_c_294_n 0.0164526f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_198 N_B_c_233_n N_A_65_367#_c_294_n 6.60564e-19 $X=2.335 $Y=1.35 $X2=0 $Y2=0
cc_199 N_B_c_228_n N_A_65_367#_c_310_n 0.0101554f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_200 N_B_c_230_n N_A_65_367#_c_310_n 0.0101649f $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_201 N_B_c_230_n N_A_65_367#_c_311_n 0.0115716f $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_202 N_B_c_228_n N_A_65_367#_c_346_n 0.0136034f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_203 N_B_c_230_n N_A_65_367#_c_346_n 7.89477e-19 $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_204 B N_A_65_367#_c_346_n 0.0202756f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_205 N_B_c_233_n N_A_65_367#_c_346_n 6.86408e-19 $X=2.335 $Y=1.35 $X2=0 $Y2=0
cc_206 N_B_M1018_g N_VPWR_c_442_n 0.00366539f $X=1.905 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B_M1018_g N_VPWR_c_447_n 0.00585385f $X=1.905 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B_M1009_g N_VPWR_c_447_n 0.00585385f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B_M1018_g N_VPWR_c_441_n 0.0108996f $X=1.905 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B_M1009_g N_VPWR_c_441_n 0.0108996f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B_c_228_n N_VGND_c_583_n 0.00239004f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_212 N_B_c_230_n N_VGND_c_584_n 0.00239004f $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_213 N_B_c_228_n N_VGND_c_588_n 0.00550269f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_214 N_B_c_230_n N_VGND_c_588_n 0.00550269f $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_215 N_B_c_228_n N_VGND_c_595_n 0.00618469f $X=1.905 $Y=1.185 $X2=0 $Y2=0
cc_216 N_B_c_230_n N_VGND_c_595_n 0.00618469f $X=2.335 $Y=1.185 $X2=0 $Y2=0
cc_217 N_A_65_367#_c_291_n N_VPWR_c_442_n 0.014892f $X=0.47 $Y=2.9 $X2=0 $Y2=0
cc_218 N_A_65_367#_M1006_g N_VPWR_c_443_n 0.0109677f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_219 N_A_65_367#_M1007_g N_VPWR_c_444_n 0.00905986f $X=3.725 $Y=2.465 $X2=0
+ $Y2=0
cc_220 N_A_65_367#_M1013_g N_VPWR_c_444_n 0.00905986f $X=4.315 $Y=2.465 $X2=0
+ $Y2=0
cc_221 N_A_65_367#_M1015_g N_VPWR_c_446_n 0.009097f $X=4.745 $Y=2.465 $X2=0
+ $Y2=0
cc_222 N_A_65_367#_c_291_n N_VPWR_c_449_n 0.0309061f $X=0.47 $Y=2.9 $X2=0 $Y2=0
cc_223 N_A_65_367#_M1006_g N_VPWR_c_450_n 0.00549284f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_224 N_A_65_367#_M1007_g N_VPWR_c_450_n 0.00549284f $X=3.725 $Y=2.465 $X2=0
+ $Y2=0
cc_225 N_A_65_367#_M1013_g N_VPWR_c_451_n 0.00549284f $X=4.315 $Y=2.465 $X2=0
+ $Y2=0
cc_226 N_A_65_367#_M1015_g N_VPWR_c_451_n 0.00549284f $X=4.745 $Y=2.465 $X2=0
+ $Y2=0
cc_227 N_A_65_367#_M1014_s N_VPWR_c_441_n 0.00466625f $X=0.325 $Y=1.835 $X2=0
+ $Y2=0
cc_228 N_A_65_367#_M1018_d N_VPWR_c_441_n 0.0119922f $X=1.98 $Y=1.835 $X2=0
+ $Y2=0
cc_229 N_A_65_367#_M1006_g N_VPWR_c_441_n 0.0102512f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_230 N_A_65_367#_M1007_g N_VPWR_c_441_n 0.0102882f $X=3.725 $Y=2.465 $X2=0
+ $Y2=0
cc_231 N_A_65_367#_M1013_g N_VPWR_c_441_n 0.0102882f $X=4.315 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_A_65_367#_M1015_g N_VPWR_c_441_n 0.0107779f $X=4.745 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_65_367#_c_291_n N_VPWR_c_441_n 0.0179149f $X=0.47 $Y=2.9 $X2=0 $Y2=0
cc_234 N_A_65_367#_c_293_n A_318_367# 0.0014668f $X=1.795 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_65_367#_M1006_g N_X_c_524_n 0.013837f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_65_367#_M1007_g N_X_c_524_n 0.0156695f $X=3.725 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_65_367#_M1013_g N_X_c_524_n 9.96931e-19 $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_65_367#_M1007_g N_X_c_519_n 0.0120022f $X=3.725 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A_65_367#_M1013_g N_X_c_519_n 0.0120022f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_65_367#_c_373_p N_X_c_519_n 0.0486665f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_241 N_A_65_367#_c_286_n N_X_c_519_n 0.00627911f $X=4.745 $Y=1.44 $X2=0 $Y2=0
cc_242 N_A_65_367#_M1006_g N_X_c_520_n 0.0028793f $X=3.295 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A_65_367#_M1007_g N_X_c_520_n 0.00134746f $X=3.725 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A_65_367#_c_373_p N_X_c_520_n 0.0264336f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_245 N_A_65_367#_c_286_n N_X_c_520_n 0.00264974f $X=4.745 $Y=1.44 $X2=0 $Y2=0
cc_246 N_A_65_367#_M1004_g N_X_c_514_n 0.0127153f $X=3.81 $Y=0.655 $X2=0 $Y2=0
cc_247 N_A_65_367#_M1005_g N_X_c_514_n 0.0113524f $X=4.275 $Y=0.655 $X2=0 $Y2=0
cc_248 N_A_65_367#_c_373_p N_X_c_514_n 0.0453297f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_249 N_A_65_367#_c_286_n N_X_c_514_n 0.00300734f $X=4.745 $Y=1.44 $X2=0 $Y2=0
cc_250 N_A_65_367#_c_283_n N_X_c_515_n 0.00390708f $X=3.245 $Y=1.275 $X2=0 $Y2=0
cc_251 N_A_65_367#_c_373_p N_X_c_515_n 0.0137341f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_252 N_A_65_367#_c_286_n N_X_c_515_n 0.00264974f $X=4.745 $Y=1.44 $X2=0 $Y2=0
cc_253 N_A_65_367#_M1004_g N_X_c_542_n 7.53442e-19 $X=3.81 $Y=0.655 $X2=0 $Y2=0
cc_254 N_A_65_367#_M1005_g N_X_c_542_n 0.0103249f $X=4.275 $Y=0.655 $X2=0 $Y2=0
cc_255 N_A_65_367#_M1007_g N_X_c_544_n 9.96931e-19 $X=3.725 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A_65_367#_M1013_g N_X_c_544_n 0.0156695f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A_65_367#_M1015_g N_X_c_544_n 0.0200389f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_65_367#_M1012_g N_X_c_516_n 0.019292f $X=4.745 $Y=0.655 $X2=0 $Y2=0
cc_259 N_A_65_367#_c_373_p N_X_c_516_n 0.00104391f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_260 N_A_65_367#_M1015_g N_X_c_521_n 0.016399f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_65_367#_M1005_g N_X_c_517_n 0.00101275f $X=4.275 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A_65_367#_c_373_p N_X_c_517_n 0.0265471f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_263 N_A_65_367#_c_286_n N_X_c_517_n 0.00340139f $X=4.745 $Y=1.44 $X2=0 $Y2=0
cc_264 N_A_65_367#_M1013_g N_X_c_522_n 0.00134746f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A_65_367#_M1015_g N_X_c_522_n 0.00227204f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A_65_367#_c_373_p N_X_c_522_n 0.0245279f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_267 N_A_65_367#_c_286_n N_X_c_522_n 0.00231808f $X=4.745 $Y=1.44 $X2=0 $Y2=0
cc_268 N_A_65_367#_M1012_g X 0.0234984f $X=4.745 $Y=0.655 $X2=0 $Y2=0
cc_269 N_A_65_367#_c_373_p X 0.0197383f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_270 N_A_65_367#_c_303_n A_154_47# 0.00518345f $X=1.625 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_271 N_A_65_367#_c_303_n N_VGND_M1001_d 0.00335711f $X=1.625 $Y=0.915
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_65_367#_c_311_n N_VGND_M1016_d 0.0152989f $X=3.16 $Y=0.915 $X2=0
+ $Y2=0
cc_273 N_A_65_367#_c_283_n N_VGND_M1016_d 0.00100449f $X=3.245 $Y=1.275 $X2=0
+ $Y2=0
cc_274 N_A_65_367#_c_280_n N_VGND_c_583_n 0.0121971f $X=0.48 $Y=0.43 $X2=0 $Y2=0
cc_275 N_A_65_367#_c_303_n N_VGND_c_583_n 0.0159912f $X=1.625 $Y=0.915 $X2=0
+ $Y2=0
cc_276 N_A_65_367#_c_310_n N_VGND_c_583_n 0.0112466f $X=2.12 $Y=0.38 $X2=0 $Y2=0
cc_277 N_A_65_367#_M1003_g N_VGND_c_584_n 0.00706372f $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_278 N_A_65_367#_c_310_n N_VGND_c_584_n 0.0112466f $X=2.12 $Y=0.38 $X2=0 $Y2=0
cc_279 N_A_65_367#_c_311_n N_VGND_c_584_n 0.0204369f $X=3.16 $Y=0.915 $X2=0
+ $Y2=0
cc_280 N_A_65_367#_M1003_g N_VGND_c_585_n 0.00124221f $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_281 N_A_65_367#_M1004_g N_VGND_c_585_n 0.0115984f $X=3.81 $Y=0.655 $X2=0
+ $Y2=0
cc_282 N_A_65_367#_M1005_g N_VGND_c_585_n 0.00538688f $X=4.275 $Y=0.655 $X2=0
+ $Y2=0
cc_283 N_A_65_367#_M1012_g N_VGND_c_587_n 0.00729581f $X=4.745 $Y=0.655 $X2=0
+ $Y2=0
cc_284 N_A_65_367#_c_310_n N_VGND_c_588_n 0.0148925f $X=2.12 $Y=0.38 $X2=0 $Y2=0
cc_285 N_A_65_367#_M1003_g N_VGND_c_590_n 0.00585385f $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_286 N_A_65_367#_M1004_g N_VGND_c_590_n 0.00486043f $X=3.81 $Y=0.655 $X2=0
+ $Y2=0
cc_287 N_A_65_367#_c_280_n N_VGND_c_592_n 0.0195196f $X=0.48 $Y=0.43 $X2=0 $Y2=0
cc_288 N_A_65_367#_M1005_g N_VGND_c_593_n 0.00549284f $X=4.275 $Y=0.655 $X2=0
+ $Y2=0
cc_289 N_A_65_367#_M1012_g N_VGND_c_593_n 0.00585385f $X=4.745 $Y=0.655 $X2=0
+ $Y2=0
cc_290 N_A_65_367#_M1002_s N_VGND_c_595_n 0.0023218f $X=0.335 $Y=0.235 $X2=0
+ $Y2=0
cc_291 N_A_65_367#_M1011_d N_VGND_c_595_n 0.00225632f $X=1.98 $Y=0.235 $X2=0
+ $Y2=0
cc_292 N_A_65_367#_M1003_g N_VGND_c_595_n 0.0106376f $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_293 N_A_65_367#_M1004_g N_VGND_c_595_n 0.00824727f $X=3.81 $Y=0.655 $X2=0
+ $Y2=0
cc_294 N_A_65_367#_M1005_g N_VGND_c_595_n 0.0101921f $X=4.275 $Y=0.655 $X2=0
+ $Y2=0
cc_295 N_A_65_367#_M1012_g N_VGND_c_595_n 0.0118044f $X=4.745 $Y=0.655 $X2=0
+ $Y2=0
cc_296 N_A_65_367#_c_280_n N_VGND_c_595_n 0.0124452f $X=0.48 $Y=0.43 $X2=0 $Y2=0
cc_297 N_A_65_367#_c_303_n N_VGND_c_595_n 0.0317345f $X=1.625 $Y=0.915 $X2=0
+ $Y2=0
cc_298 N_A_65_367#_c_281_n N_VGND_c_595_n 0.0232101f $X=0.645 $Y=0.915 $X2=0
+ $Y2=0
cc_299 N_A_65_367#_c_310_n N_VGND_c_595_n 0.0120439f $X=2.12 $Y=0.38 $X2=0 $Y2=0
cc_300 N_A_65_367#_c_311_n N_VGND_c_595_n 0.00959099f $X=3.16 $Y=0.915 $X2=0
+ $Y2=0
cc_301 N_A_65_367#_c_282_n A_318_47# 3.7257e-19 $X=1.71 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_302 N_A_65_367#_c_346_n A_318_47# 0.00288418f $X=2.285 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_303 N_A_65_367#_c_311_n A_482_47# 0.00461646f $X=3.16 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_304 A_154_367# N_VPWR_c_441_n 0.010279f $X=0.77 $Y=1.835 $X2=0 $Y2=0
cc_305 N_VPWR_c_441_n A_318_367# 0.010279f $X=5.04 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_306 N_VPWR_c_441_n A_482_367# 0.010279f $X=5.04 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_307 N_VPWR_c_441_n N_X_M1006_s 0.00223819f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_441_n N_X_M1013_s 0.00223819f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_c_450_n N_X_c_524_n 0.0177952f $X=3.855 $Y=3.33 $X2=0 $Y2=0
cc_310 N_VPWR_c_441_n N_X_c_524_n 0.0123247f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_311 N_VPWR_M1007_d N_X_c_519_n 0.00407652f $X=3.8 $Y=1.835 $X2=0 $Y2=0
cc_312 N_VPWR_c_444_n N_X_c_519_n 0.0254128f $X=4.02 $Y=2.3 $X2=0 $Y2=0
cc_313 N_VPWR_c_443_n N_X_c_520_n 0.00800069f $X=3 $Y=1.96 $X2=0 $Y2=0
cc_314 N_VPWR_c_451_n N_X_c_544_n 0.0177952f $X=4.875 $Y=3.33 $X2=0 $Y2=0
cc_315 N_VPWR_c_441_n N_X_c_544_n 0.0123247f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_316 N_VPWR_M1015_d N_X_c_521_n 0.00324991f $X=4.82 $Y=1.835 $X2=0 $Y2=0
cc_317 N_VPWR_c_446_n N_X_c_521_n 0.0209617f $X=4.96 $Y=2.3 $X2=0 $Y2=0
cc_318 N_X_c_514_n N_VGND_M1004_d 0.00311564f $X=4.325 $Y=1.01 $X2=0 $Y2=0
cc_319 N_X_c_516_n N_VGND_M1012_d 0.00420987f $X=4.925 $Y=1.01 $X2=0 $Y2=0
cc_320 N_X_c_514_n N_VGND_c_585_n 0.0147641f $X=4.325 $Y=1.01 $X2=0 $Y2=0
cc_321 N_X_c_542_n N_VGND_c_585_n 0.0304484f $X=4.49 $Y=0.43 $X2=0 $Y2=0
cc_322 N_X_c_516_n N_VGND_c_587_n 0.0236067f $X=4.925 $Y=1.01 $X2=0 $Y2=0
cc_323 N_X_c_575_p N_VGND_c_590_n 0.0110337f $X=3.595 $Y=0.43 $X2=0 $Y2=0
cc_324 N_X_c_542_n N_VGND_c_593_n 0.0183971f $X=4.49 $Y=0.43 $X2=0 $Y2=0
cc_325 N_X_M1003_s N_VGND_c_595_n 0.00606379f $X=3.455 $Y=0.235 $X2=0 $Y2=0
cc_326 N_X_M1005_s N_VGND_c_595_n 0.00308191f $X=4.35 $Y=0.235 $X2=0 $Y2=0
cc_327 N_X_c_575_p N_VGND_c_595_n 0.00648955f $X=3.595 $Y=0.43 $X2=0 $Y2=0
cc_328 N_X_c_542_n N_VGND_c_595_n 0.012508f $X=4.49 $Y=0.43 $X2=0 $Y2=0
cc_329 A_154_47# N_VGND_c_595_n 0.003486f $X=0.77 $Y=0.235 $X2=2.12 $Y2=1.96
cc_330 N_VGND_c_595_n A_318_47# 0.003486f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_331 N_VGND_c_595_n A_482_47# 0.003486f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
