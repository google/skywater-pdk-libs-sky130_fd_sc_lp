* File: sky130_fd_sc_lp__o311ai_1.spice
* Created: Fri Aug 28 11:14:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o311ai_1  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_A_173_47#_M1000_d N_A1_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_173_47#_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1008 N_A_173_47#_M1008_d N_A3_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1512 PD=1.46 PS=1.2 NRD=0 NRS=5.712 M=1 R=5.6 SA=75001.1
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1002 A_515_47# N_B1_M1002_g N_A_173_47#_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2604 PD=1.05 PS=1.46 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g A_515_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75002.3 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1009 A_173_367# N_A1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1827 AS=0.3339 PD=1.55 PS=3.05 NRD=14.0658 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1001 A_261_367# N_A2_M1001_g A_173_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.1953
+ AS=0.1827 PD=1.57 PS=1.55 NRD=15.6221 NRS=14.0658 M=1 R=8.4 SA=75000.6
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A3_M1005_g A_261_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1953 PD=1.65 PS=1.57 NRD=8.5892 NRS=15.6221 M=1 R=8.4 SA=75001.1
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3024 AS=0.2457 PD=1.74 PS=1.65 NRD=15.6221 NRS=8.5892 M=1 R=8.4
+ SA=75001.6 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3024 PD=3.05 PS=1.74 NRD=0 NRS=15.6221 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o311ai_1.pxi.spice"
*
.ends
*
*
