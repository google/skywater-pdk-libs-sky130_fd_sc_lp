* File: sky130_fd_sc_lp__o2111ai_2.pxi.spice
* Created: Fri Aug 28 11:01:03 2020
* 
x_PM_SKY130_FD_SC_LP__O2111AI_2%D1 N_D1_c_90_n N_D1_M1012_g N_D1_M1009_g
+ N_D1_c_92_n N_D1_M1015_g N_D1_M1018_g D1 D1 N_D1_c_95_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%D1
x_PM_SKY130_FD_SC_LP__O2111AI_2%C1 N_C1_c_132_n N_C1_M1001_g N_C1_M1000_g
+ N_C1_c_134_n N_C1_M1011_g N_C1_M1010_g C1 C1 N_C1_c_137_n N_C1_c_138_n C1
+ PM_SKY130_FD_SC_LP__O2111AI_2%C1
x_PM_SKY130_FD_SC_LP__O2111AI_2%B1 N_B1_M1006_g N_B1_M1016_g N_B1_c_194_n
+ N_B1_M1005_g N_B1_c_195_n N_B1_M1017_g B1 B1 B1 N_B1_c_197_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%B1
x_PM_SKY130_FD_SC_LP__O2111AI_2%A2 N_A2_c_243_n N_A2_M1004_g N_A2_M1003_g
+ N_A2_c_245_n N_A2_M1013_g N_A2_M1014_g A2 A2 N_A2_c_248_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%A2
x_PM_SKY130_FD_SC_LP__O2111AI_2%A1 N_A1_c_291_n N_A1_M1002_g N_A1_M1007_g
+ N_A1_c_293_n N_A1_M1008_g N_A1_M1019_g A1 A1 N_A1_c_296_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%A1
x_PM_SKY130_FD_SC_LP__O2111AI_2%VPWR N_VPWR_M1009_s N_VPWR_M1018_s
+ N_VPWR_M1010_d N_VPWR_M1016_d N_VPWR_M1007_s N_VPWR_c_329_n N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n
+ VPWR N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_328_n N_VPWR_c_344_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O2111AI_2%Y N_Y_M1012_s N_Y_M1009_d N_Y_M1000_s
+ N_Y_M1006_s N_Y_M1003_s N_Y_c_417_n N_Y_c_418_n N_Y_c_412_n N_Y_c_463_n
+ N_Y_c_413_n N_Y_c_467_n N_Y_c_414_n N_Y_c_453_n N_Y_c_421_n N_Y_c_415_n
+ N_Y_c_416_n Y Y Y PM_SKY130_FD_SC_LP__O2111AI_2%Y
x_PM_SKY130_FD_SC_LP__O2111AI_2%A_694_367# N_A_694_367#_M1003_d
+ N_A_694_367#_M1014_d N_A_694_367#_M1019_d N_A_694_367#_c_483_n
+ N_A_694_367#_c_484_n N_A_694_367#_c_490_n N_A_694_367#_c_511_n
+ N_A_694_367#_c_485_n N_A_694_367#_c_481_n N_A_694_367#_c_482_n
+ N_A_694_367#_c_488_n PM_SKY130_FD_SC_LP__O2111AI_2%A_694_367#
x_PM_SKY130_FD_SC_LP__O2111AI_2%A_43_69# N_A_43_69#_M1012_d N_A_43_69#_M1015_d
+ N_A_43_69#_M1011_s N_A_43_69#_c_523_n N_A_43_69#_c_524_n N_A_43_69#_c_525_n
+ N_A_43_69#_c_532_n N_A_43_69#_c_537_n N_A_43_69#_c_526_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%A_43_69#
x_PM_SKY130_FD_SC_LP__O2111AI_2%A_298_69# N_A_298_69#_M1001_d
+ N_A_298_69#_M1005_d N_A_298_69#_c_561_n N_A_298_69#_c_559_n
+ N_A_298_69#_c_560_n N_A_298_69#_c_566_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%A_298_69#
x_PM_SKY130_FD_SC_LP__O2111AI_2%A_522_47# N_A_522_47#_M1005_s
+ N_A_522_47#_M1017_s N_A_522_47#_M1013_s N_A_522_47#_M1008_s
+ N_A_522_47#_c_585_n N_A_522_47#_c_616_p N_A_522_47#_c_593_n
+ N_A_522_47#_c_615_p N_A_522_47#_c_597_n N_A_522_47#_c_586_n
+ N_A_522_47#_c_587_n N_A_522_47#_c_592_n N_A_522_47#_c_598_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%A_522_47#
x_PM_SKY130_FD_SC_LP__O2111AI_2%VGND N_VGND_M1004_d N_VGND_M1002_d
+ N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n N_VGND_c_631_n VGND
+ N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n
+ PM_SKY130_FD_SC_LP__O2111AI_2%VGND
cc_1 VNB N_D1_c_90_n 0.019103f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.295
cc_2 VNB N_D1_M1009_g 0.00146396f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_3 VNB N_D1_c_92_n 0.0159497f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.295
cc_4 VNB N_D1_M1018_g 0.00140289f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_5 VNB D1 0.0231981f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_D1_c_95_n 0.0713621f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.46
cc_7 VNB N_C1_c_132_n 0.0164884f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.295
cc_8 VNB N_C1_M1000_g 0.00152181f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_9 VNB N_C1_c_134_n 0.0189138f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.295
cc_10 VNB N_C1_M1010_g 0.00152414f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_11 VNB C1 0.00309584f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_C1_c_137_n 0.0462109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C1_c_138_n 0.00716768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_M1006_g 0.00699606f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.765
cc_15 VNB N_B1_M1016_g 0.0111855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_194_n 0.0202392f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.765
cc_17 VNB N_B1_c_195_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_18 VNB B1 0.00735359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_197_n 0.0998978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_c_243_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.295
cc_21 VNB N_A2_M1003_g 0.0111836f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_22 VNB N_A2_c_245_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.295
cc_23 VNB N_A2_M1014_g 0.00728783f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_24 VNB A2 0.0063768f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_A2_c_248_n 0.0364761f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.46
cc_26 VNB N_A1_c_291_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.295
cc_27 VNB N_A1_M1007_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_28 VNB N_A1_c_293_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.295
cc_29 VNB N_A1_M1019_g 0.0100771f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_30 VNB A1 0.0327159f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_A1_c_296_n 0.0414337f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.46
cc_32 VNB N_VPWR_c_328_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_694_367#_c_481_n 0.0083778f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.46
cc_34 VNB N_A_694_367#_c_482_n 0.00238941f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.46
cc_35 VNB N_A_43_69#_c_523_n 0.023359f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_36 VNB N_A_43_69#_c_524_n 0.00513046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_43_69#_c_525_n 0.00935084f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_38 VNB N_A_43_69#_c_526_n 0.0132783f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.46
cc_39 VNB N_A_298_69#_c_559_n 0.0187028f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.625
cc_40 VNB N_A_298_69#_c_560_n 0.00270685f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_41 VNB N_A_522_47#_c_585_n 0.00329826f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_42 VNB N_A_522_47#_c_586_n 0.0075508f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.46
cc_43 VNB N_A_522_47#_c_587_n 0.0224525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_628_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.765
cc_45 VNB N_VGND_c_629_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_46 VNB N_VGND_c_630_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_47 VNB N_VGND_c_631_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_632_n 0.093411f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.46
cc_49 VNB N_VGND_c_633_n 0.0212629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_634_n 0.313485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_635_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_D1_M1009_g 0.02456f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_53 VPB N_D1_M1018_g 0.0186121f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_54 VPB D1 0.010012f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_55 VPB N_C1_M1000_g 0.0190736f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_56 VPB N_C1_M1010_g 0.0190778f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_57 VPB N_B1_M1006_g 0.0190608f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.765
cc_58 VPB N_B1_M1016_g 0.0234993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A2_M1003_g 0.0243601f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_60 VPB N_A2_M1014_g 0.019469f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_61 VPB N_A1_M1007_g 0.018727f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_62 VPB N_A1_M1019_g 0.0232847f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_63 VPB N_VPWR_c_329_n 0.0125627f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_64 VPB N_VPWR_c_330_n 0.0484034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_331_n 3.22457e-19 $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.46
cc_66 VPB N_VPWR_c_332_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.665
cc_67 VPB N_VPWR_c_333_n 0.0153577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_334_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_335_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_336_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_337_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_338_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_339_n 0.0401167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_340_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_341_n 0.0156522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_342_n 0.0212501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_328_n 0.0701193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_344_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_Y_c_412_n 0.00405562f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_80 VPB N_Y_c_413_n 0.00523247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_Y_c_414_n 0.0261131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_Y_c_415_n 0.00155509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_Y_c_416_n 0.00391071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_694_367#_c_483_n 0.00226522f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.765
cc_85 VPB N_A_694_367#_c_484_n 0.0103399f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_86 VPB N_A_694_367#_c_485_n 9.3142e-19 $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.46
cc_87 VPB N_A_694_367#_c_481_n 0.0110324f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.46
cc_88 VPB N_A_694_367#_c_482_n 0.00105268f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.46
cc_89 VPB N_A_694_367#_c_488_n 0.0498589f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.46
cc_90 N_D1_c_92_n N_C1_c_132_n 0.0153606f $X=0.985 $Y=1.295 $X2=-0.19 $Y2=-0.245
cc_91 N_D1_M1018_g N_C1_M1000_g 0.0219054f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_92 N_D1_c_95_n N_C1_c_137_n 0.0226329f $X=0.985 $Y=1.46 $X2=0 $Y2=0
cc_93 N_D1_c_92_n N_C1_c_138_n 0.00284524f $X=0.985 $Y=1.295 $X2=0 $Y2=0
cc_94 N_D1_M1009_g N_VPWR_c_330_n 0.00466141f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_95 D1 N_VPWR_c_330_n 0.0219561f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_96 N_D1_c_95_n N_VPWR_c_330_n 0.00144174f $X=0.985 $Y=1.46 $X2=0 $Y2=0
cc_97 N_D1_M1009_g N_VPWR_c_331_n 8.27324e-19 $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_98 N_D1_M1018_g N_VPWR_c_331_n 0.014363f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_99 N_D1_M1009_g N_VPWR_c_341_n 0.00533769f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_100 N_D1_M1018_g N_VPWR_c_341_n 0.00486043f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_101 N_D1_M1009_g N_VPWR_c_328_n 0.0104224f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_102 N_D1_M1018_g N_VPWR_c_328_n 0.00824727f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_103 N_D1_M1009_g N_Y_c_417_n 0.0147089f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_104 N_D1_c_90_n N_Y_c_418_n 0.0104429f $X=0.555 $Y=1.295 $X2=0 $Y2=0
cc_105 N_D1_c_92_n N_Y_c_418_n 0.00717238f $X=0.985 $Y=1.295 $X2=0 $Y2=0
cc_106 N_D1_M1018_g N_Y_c_412_n 0.0141566f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_107 N_D1_M1009_g N_Y_c_421_n 0.0090904f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_108 N_D1_M1018_g N_Y_c_421_n 0.00252935f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_109 N_D1_c_90_n Y 0.00471292f $X=0.555 $Y=1.295 $X2=0 $Y2=0
cc_110 N_D1_M1009_g Y 0.00295895f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_111 N_D1_c_92_n Y 0.00297999f $X=0.985 $Y=1.295 $X2=0 $Y2=0
cc_112 N_D1_M1018_g Y 0.00383878f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_113 D1 Y 0.0414577f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_114 N_D1_c_95_n Y 0.0231139f $X=0.985 $Y=1.46 $X2=0 $Y2=0
cc_115 D1 N_A_43_69#_c_523_n 0.022426f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_116 N_D1_c_95_n N_A_43_69#_c_523_n 0.0015759f $X=0.985 $Y=1.46 $X2=0 $Y2=0
cc_117 N_D1_c_90_n N_A_43_69#_c_524_n 0.0128219f $X=0.555 $Y=1.295 $X2=0 $Y2=0
cc_118 N_D1_c_92_n N_A_43_69#_c_524_n 0.0119696f $X=0.985 $Y=1.295 $X2=0 $Y2=0
cc_119 N_D1_c_90_n N_VGND_c_632_n 0.0029147f $X=0.555 $Y=1.295 $X2=0 $Y2=0
cc_120 N_D1_c_92_n N_VGND_c_632_n 0.0029147f $X=0.985 $Y=1.295 $X2=0 $Y2=0
cc_121 N_D1_c_90_n N_VGND_c_634_n 0.00421708f $X=0.555 $Y=1.295 $X2=0 $Y2=0
cc_122 N_D1_c_92_n N_VGND_c_634_n 0.00399217f $X=0.985 $Y=1.295 $X2=0 $Y2=0
cc_123 N_C1_M1010_g N_B1_M1006_g 0.0222755f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_124 N_C1_c_134_n B1 3.13738e-19 $X=1.845 $Y=1.295 $X2=0 $Y2=0
cc_125 C1 B1 0.00965239f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_C1_c_137_n B1 4.72303e-19 $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_127 N_C1_c_134_n N_B1_c_197_n 0.00274659f $X=1.845 $Y=1.295 $X2=0 $Y2=0
cc_128 C1 N_B1_c_197_n 0.00147149f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_129 N_C1_c_137_n N_B1_c_197_n 0.0203933f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_130 N_C1_M1000_g N_VPWR_c_331_n 0.0141832f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_131 N_C1_M1010_g N_VPWR_c_331_n 7.27171e-19 $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_132 N_C1_M1000_g N_VPWR_c_332_n 7.27171e-19 $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_133 N_C1_M1010_g N_VPWR_c_332_n 0.0141832f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_134 N_C1_M1000_g N_VPWR_c_335_n 0.00486043f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_135 N_C1_M1010_g N_VPWR_c_335_n 0.00486043f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_136 N_C1_M1000_g N_VPWR_c_328_n 0.00824727f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_137 N_C1_M1010_g N_VPWR_c_328_n 0.00824727f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_138 N_C1_c_132_n N_Y_c_418_n 7.66511e-19 $X=1.415 $Y=1.295 $X2=0 $Y2=0
cc_139 N_C1_M1000_g N_Y_c_412_n 0.0134064f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_140 N_C1_c_137_n N_Y_c_412_n 0.00168053f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_141 N_C1_c_138_n N_Y_c_412_n 0.027704f $X=1.608 $Y=1.377 $X2=0 $Y2=0
cc_142 N_C1_M1010_g N_Y_c_413_n 0.0134005f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_143 C1 N_Y_c_413_n 0.0158045f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_C1_c_137_n N_Y_c_413_n 0.00167966f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_145 C1 N_Y_c_415_n 0.00846419f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_C1_c_137_n N_Y_c_415_n 0.00251445f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_147 N_C1_c_138_n N_Y_c_415_n 0.00522892f $X=1.608 $Y=1.377 $X2=0 $Y2=0
cc_148 N_C1_M1000_g Y 6.26061e-19 $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_149 N_C1_c_137_n Y 4.71559e-19 $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_150 N_C1_c_138_n Y 0.0280434f $X=1.608 $Y=1.377 $X2=0 $Y2=0
cc_151 N_C1_c_132_n N_A_43_69#_c_524_n 8.02085e-19 $X=1.415 $Y=1.295 $X2=0 $Y2=0
cc_152 N_C1_c_132_n N_A_43_69#_c_532_n 0.0127342f $X=1.415 $Y=1.295 $X2=0 $Y2=0
cc_153 N_C1_c_134_n N_A_43_69#_c_532_n 0.0105779f $X=1.845 $Y=1.295 $X2=0 $Y2=0
cc_154 C1 N_A_43_69#_c_532_n 0.0171847f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_155 N_C1_c_137_n N_A_43_69#_c_532_n 5.7861e-19 $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_156 N_C1_c_138_n N_A_43_69#_c_532_n 0.0179973f $X=1.608 $Y=1.377 $X2=0 $Y2=0
cc_157 N_C1_c_137_n N_A_43_69#_c_537_n 2.80421e-19 $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_158 N_C1_c_138_n N_A_43_69#_c_537_n 0.0166693f $X=1.608 $Y=1.377 $X2=0 $Y2=0
cc_159 N_C1_c_134_n N_A_43_69#_c_526_n 5.83502e-19 $X=1.845 $Y=1.295 $X2=0 $Y2=0
cc_160 C1 N_A_43_69#_c_526_n 0.00353481f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_161 N_C1_c_137_n N_A_43_69#_c_526_n 0.00112306f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_162 N_C1_c_134_n N_A_298_69#_c_561_n 0.00786076f $X=1.845 $Y=1.295 $X2=0
+ $Y2=0
cc_163 N_C1_c_134_n N_A_298_69#_c_559_n 0.0104977f $X=1.845 $Y=1.295 $X2=0 $Y2=0
cc_164 N_C1_c_132_n N_A_298_69#_c_560_n 7.85031e-19 $X=1.415 $Y=1.295 $X2=0
+ $Y2=0
cc_165 N_C1_c_134_n N_A_298_69#_c_560_n 9.46184e-19 $X=1.845 $Y=1.295 $X2=0
+ $Y2=0
cc_166 N_C1_c_132_n N_VGND_c_632_n 0.00482246f $X=1.415 $Y=1.295 $X2=0 $Y2=0
cc_167 N_C1_c_134_n N_VGND_c_632_n 0.00291465f $X=1.845 $Y=1.295 $X2=0 $Y2=0
cc_168 N_C1_c_132_n N_VGND_c_634_n 0.00955107f $X=1.415 $Y=1.295 $X2=0 $Y2=0
cc_169 N_C1_c_134_n N_VGND_c_634_n 0.00428625f $X=1.845 $Y=1.295 $X2=0 $Y2=0
cc_170 N_B1_c_195_n N_A2_c_243_n 0.0154574f $X=3.38 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_171 B1 A2 0.022107f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_172 B1 N_A2_c_248_n 0.00515655f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_173 N_B1_c_197_n N_A2_c_248_n 0.0154574f $X=3.29 $Y=1.35 $X2=0 $Y2=0
cc_174 N_B1_M1006_g N_VPWR_c_332_n 0.0141832f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B1_M1016_g N_VPWR_c_332_n 7.27171e-19 $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_176 N_B1_M1006_g N_VPWR_c_333_n 7.6326e-19 $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_177 N_B1_M1016_g N_VPWR_c_333_n 0.0174479f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B1_M1006_g N_VPWR_c_337_n 0.00486043f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_179 N_B1_M1016_g N_VPWR_c_337_n 0.00486043f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B1_M1006_g N_VPWR_c_328_n 0.00824727f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B1_M1016_g N_VPWR_c_328_n 0.00824727f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B1_M1006_g N_Y_c_413_n 0.0158803f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B1_M1016_g N_Y_c_414_n 0.0159238f $X=2.705 $Y=2.465 $X2=0 $Y2=0
cc_184 B1 N_Y_c_414_n 0.084568f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B1_c_197_n N_Y_c_414_n 0.017025f $X=3.29 $Y=1.35 $X2=0 $Y2=0
cc_186 N_B1_M1006_g N_Y_c_416_n 0.0022704f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_187 B1 N_Y_c_416_n 0.010964f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_188 N_B1_c_197_n N_Y_c_416_n 0.00243529f $X=3.29 $Y=1.35 $X2=0 $Y2=0
cc_189 N_B1_M1016_g N_A_694_367#_c_484_n 0.00184493f $X=2.705 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_B1_c_194_n N_A_43_69#_c_526_n 0.00670191f $X=2.95 $Y=1.185 $X2=0 $Y2=0
cc_191 B1 N_A_43_69#_c_526_n 0.00159424f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_192 N_B1_c_197_n N_A_43_69#_c_526_n 0.00267246f $X=3.29 $Y=1.35 $X2=0 $Y2=0
cc_193 N_B1_c_194_n N_A_298_69#_c_559_n 0.0106146f $X=2.95 $Y=1.185 $X2=0 $Y2=0
cc_194 N_B1_c_194_n N_A_298_69#_c_566_n 0.00963096f $X=2.95 $Y=1.185 $X2=0 $Y2=0
cc_195 N_B1_c_195_n N_A_298_69#_c_566_n 0.00441544f $X=3.38 $Y=1.185 $X2=0 $Y2=0
cc_196 N_B1_c_194_n N_A_522_47#_c_585_n 0.0110927f $X=2.95 $Y=1.185 $X2=0 $Y2=0
cc_197 N_B1_c_195_n N_A_522_47#_c_585_n 0.011445f $X=3.38 $Y=1.185 $X2=0 $Y2=0
cc_198 B1 N_A_522_47#_c_585_n 0.0616182f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_199 N_B1_c_197_n N_A_522_47#_c_585_n 0.00984579f $X=3.29 $Y=1.35 $X2=0 $Y2=0
cc_200 B1 N_A_522_47#_c_592_n 0.0153941f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_201 N_B1_c_195_n N_VGND_c_628_n 0.00121106f $X=3.38 $Y=1.185 $X2=0 $Y2=0
cc_202 N_B1_c_194_n N_VGND_c_632_n 0.00359361f $X=2.95 $Y=1.185 $X2=0 $Y2=0
cc_203 N_B1_c_195_n N_VGND_c_632_n 0.0054895f $X=3.38 $Y=1.185 $X2=0 $Y2=0
cc_204 N_B1_c_194_n N_VGND_c_634_n 0.00681249f $X=2.95 $Y=1.185 $X2=0 $Y2=0
cc_205 N_B1_c_195_n N_VGND_c_634_n 0.00616748f $X=3.38 $Y=1.185 $X2=0 $Y2=0
cc_206 N_A2_c_245_n N_A1_c_291_n 0.0192951f $X=4.24 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A2_M1014_g N_A1_M1007_g 0.0192951f $X=4.24 $Y=2.465 $X2=0 $Y2=0
cc_208 A2 A1 0.0209934f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_209 A2 N_A1_c_296_n 0.0106351f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A2_c_248_n N_A1_c_296_n 0.0192951f $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_211 N_A2_M1003_g N_VPWR_c_333_n 0.00176621f $X=3.81 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A2_M1014_g N_VPWR_c_334_n 0.00109252f $X=4.24 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A2_M1003_g N_VPWR_c_339_n 0.00357877f $X=3.81 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A2_M1014_g N_VPWR_c_339_n 0.00357877f $X=4.24 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A2_M1003_g N_VPWR_c_328_n 0.00665089f $X=3.81 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A2_M1014_g N_VPWR_c_328_n 0.00537654f $X=4.24 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A2_M1003_g N_Y_c_414_n 0.0177629f $X=3.81 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A2_M1014_g N_Y_c_414_n 0.00395535f $X=4.24 $Y=2.465 $X2=0 $Y2=0
cc_219 A2 N_Y_c_414_n 0.0199733f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A2_c_248_n N_Y_c_414_n 0.00245863f $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_221 N_A2_M1003_g N_Y_c_453_n 0.0152162f $X=3.81 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A2_M1014_g N_Y_c_453_n 0.00921043f $X=4.24 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A2_M1003_g N_A_694_367#_c_490_n 0.0114565f $X=3.81 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A2_M1014_g N_A_694_367#_c_490_n 0.0115031f $X=4.24 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A2_M1014_g N_A_694_367#_c_485_n 0.00107035f $X=4.24 $Y=2.465 $X2=0
+ $Y2=0
cc_226 A2 N_A_694_367#_c_481_n 0.00904104f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_227 N_A2_M1014_g N_A_694_367#_c_482_n 0.00330334f $X=4.24 $Y=2.465 $X2=0
+ $Y2=0
cc_228 A2 N_A_694_367#_c_482_n 0.0164807f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_229 N_A2_c_243_n N_A_522_47#_c_593_n 0.0115651f $X=3.81 $Y=1.185 $X2=0 $Y2=0
cc_230 N_A2_c_245_n N_A_522_47#_c_593_n 0.00973618f $X=4.24 $Y=1.185 $X2=0 $Y2=0
cc_231 A2 N_A_522_47#_c_593_n 0.029734f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_232 N_A2_c_248_n N_A_522_47#_c_593_n 0.00224206f $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_233 A2 N_A_522_47#_c_597_n 0.00735053f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_234 A2 N_A_522_47#_c_598_n 0.0150671f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_235 N_A2_c_243_n N_VGND_c_628_n 0.0111514f $X=3.81 $Y=1.185 $X2=0 $Y2=0
cc_236 N_A2_c_245_n N_VGND_c_628_n 0.0100168f $X=4.24 $Y=1.185 $X2=0 $Y2=0
cc_237 N_A2_c_245_n N_VGND_c_629_n 5.68743e-19 $X=4.24 $Y=1.185 $X2=0 $Y2=0
cc_238 N_A2_c_245_n N_VGND_c_630_n 0.00486043f $X=4.24 $Y=1.185 $X2=0 $Y2=0
cc_239 N_A2_c_243_n N_VGND_c_632_n 0.00486043f $X=3.81 $Y=1.185 $X2=0 $Y2=0
cc_240 N_A2_c_243_n N_VGND_c_634_n 0.0045769f $X=3.81 $Y=1.185 $X2=0 $Y2=0
cc_241 N_A2_c_245_n N_VGND_c_634_n 0.0045769f $X=4.24 $Y=1.185 $X2=0 $Y2=0
cc_242 N_A1_M1007_g N_VPWR_c_334_n 0.0185929f $X=4.67 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A1_M1019_g N_VPWR_c_334_n 0.0194824f $X=5.1 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A1_M1007_g N_VPWR_c_339_n 0.00486043f $X=4.67 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A1_M1019_g N_VPWR_c_342_n 0.00486043f $X=5.1 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A1_M1007_g N_VPWR_c_328_n 0.0082726f $X=4.67 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A1_M1019_g N_VPWR_c_328_n 0.00931409f $X=5.1 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A1_M1007_g N_A_694_367#_c_485_n 0.0014373f $X=4.67 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A1_M1007_g N_A_694_367#_c_481_n 0.0148258f $X=4.67 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A1_M1019_g N_A_694_367#_c_481_n 0.0156808f $X=5.1 $Y=2.465 $X2=0 $Y2=0
cc_251 A1 N_A_694_367#_c_481_n 0.0497307f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_252 N_A1_c_296_n N_A_694_367#_c_481_n 0.00251391f $X=5.1 $Y=1.35 $X2=0 $Y2=0
cc_253 N_A1_M1019_g N_A_694_367#_c_488_n 0.0046421f $X=5.1 $Y=2.465 $X2=0 $Y2=0
cc_254 N_A1_c_291_n N_A_522_47#_c_597_n 0.0106855f $X=4.67 $Y=1.185 $X2=0 $Y2=0
cc_255 N_A1_c_293_n N_A_522_47#_c_597_n 0.00974987f $X=5.1 $Y=1.185 $X2=0 $Y2=0
cc_256 A1 N_A_522_47#_c_597_n 0.0231795f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_257 N_A1_c_296_n N_A_522_47#_c_597_n 0.00228466f $X=5.1 $Y=1.35 $X2=0 $Y2=0
cc_258 A1 N_A_522_47#_c_586_n 0.0216244f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_259 N_A1_c_291_n N_VGND_c_628_n 5.68743e-19 $X=4.67 $Y=1.185 $X2=0 $Y2=0
cc_260 N_A1_c_291_n N_VGND_c_629_n 0.0100168f $X=4.67 $Y=1.185 $X2=0 $Y2=0
cc_261 N_A1_c_293_n N_VGND_c_629_n 0.0116902f $X=5.1 $Y=1.185 $X2=0 $Y2=0
cc_262 N_A1_c_291_n N_VGND_c_630_n 0.00486043f $X=4.67 $Y=1.185 $X2=0 $Y2=0
cc_263 N_A1_c_293_n N_VGND_c_633_n 0.00486043f $X=5.1 $Y=1.185 $X2=0 $Y2=0
cc_264 N_A1_c_291_n N_VGND_c_634_n 0.0045769f $X=4.67 $Y=1.185 $X2=0 $Y2=0
cc_265 N_A1_c_293_n N_VGND_c_634_n 0.00561839f $X=5.1 $Y=1.185 $X2=0 $Y2=0
cc_266 N_VPWR_c_328_n N_Y_M1009_d 0.00380103f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_328_n N_Y_M1000_s 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_c_328_n N_Y_M1006_s 0.00571434f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_c_328_n N_Y_M1003_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_270 N_VPWR_c_341_n N_Y_c_417_n 0.0163698f $X=1.035 $Y=3.33 $X2=0 $Y2=0
cc_271 N_VPWR_c_328_n N_Y_c_417_n 0.0101905f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_M1018_s N_Y_c_412_n 0.00176461f $X=1.06 $Y=1.835 $X2=0 $Y2=0
cc_273 N_VPWR_c_331_n N_Y_c_412_n 0.0170777f $X=1.2 $Y=2.18 $X2=0 $Y2=0
cc_274 N_VPWR_c_335_n N_Y_c_463_n 0.0124525f $X=1.895 $Y=3.33 $X2=0 $Y2=0
cc_275 N_VPWR_c_328_n N_Y_c_463_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_276 N_VPWR_M1010_d N_Y_c_413_n 0.00176461f $X=1.92 $Y=1.835 $X2=0 $Y2=0
cc_277 N_VPWR_c_332_n N_Y_c_413_n 0.0170777f $X=2.06 $Y=2.18 $X2=0 $Y2=0
cc_278 N_VPWR_c_337_n N_Y_c_467_n 0.0120977f $X=2.755 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_c_328_n N_Y_c_467_n 0.00691495f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_280 N_VPWR_M1016_d N_Y_c_414_n 0.00230047f $X=2.78 $Y=1.835 $X2=0 $Y2=0
cc_281 N_VPWR_c_333_n N_Y_c_414_n 0.0220026f $X=2.92 $Y=2.11 $X2=0 $Y2=0
cc_282 N_VPWR_c_328_n N_A_694_367#_M1003_d 0.00215161f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_283 N_VPWR_c_328_n N_A_694_367#_M1014_d 0.00376627f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_328_n N_A_694_367#_M1019_d 0.00371702f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_333_n N_A_694_367#_c_483_n 0.00919722f $X=2.92 $Y=2.11 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_339_n N_A_694_367#_c_483_n 0.0179183f $X=4.72 $Y=3.33 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_328_n N_A_694_367#_c_483_n 0.0101082f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_333_n N_A_694_367#_c_484_n 0.0440921f $X=2.92 $Y=2.11 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_339_n N_A_694_367#_c_490_n 0.0361172f $X=4.72 $Y=3.33 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_328_n N_A_694_367#_c_490_n 0.023676f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_291 N_VPWR_c_339_n N_A_694_367#_c_511_n 0.0125234f $X=4.72 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_328_n N_A_694_367#_c_511_n 0.0073762f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_334_n N_A_694_367#_c_481_n 0.0216087f $X=4.885 $Y=2.03 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_342_n N_A_694_367#_c_488_n 0.0178111f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_328_n N_A_694_367#_c_488_n 0.0100304f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_296 N_Y_c_414_n N_A_694_367#_M1003_d 0.00230047f $X=3.86 $Y=1.77 $X2=-0.19
+ $Y2=1.655
cc_297 N_Y_c_414_n N_A_694_367#_c_484_n 0.0202165f $X=3.86 $Y=1.77 $X2=0 $Y2=0
cc_298 N_Y_M1003_s N_A_694_367#_c_490_n 0.00332344f $X=3.885 $Y=1.835 $X2=0
+ $Y2=0
cc_299 N_Y_c_453_n N_A_694_367#_c_490_n 0.0159805f $X=4.025 $Y=1.97 $X2=0 $Y2=0
cc_300 N_Y_c_414_n N_A_694_367#_c_485_n 0.00559861f $X=3.86 $Y=1.77 $X2=0 $Y2=0
cc_301 N_Y_c_414_n N_A_694_367#_c_482_n 0.00802274f $X=3.86 $Y=1.77 $X2=0 $Y2=0
cc_302 N_Y_M1012_s N_A_43_69#_c_524_n 0.00176461f $X=0.63 $Y=0.345 $X2=0 $Y2=0
cc_303 N_Y_c_418_n N_A_43_69#_c_524_n 0.0159805f $X=0.77 $Y=0.68 $X2=0 $Y2=0
cc_304 N_Y_c_413_n N_A_43_69#_c_526_n 0.0102092f $X=2.385 $Y=1.84 $X2=0 $Y2=0
cc_305 N_Y_c_414_n N_A_522_47#_c_593_n 0.00336914f $X=3.86 $Y=1.77 $X2=0 $Y2=0
cc_306 N_A_694_367#_c_481_n N_A_522_47#_c_597_n 0.00389734f $X=5.22 $Y=1.69
+ $X2=0 $Y2=0
cc_307 N_A_43_69#_c_532_n N_A_298_69#_M1001_d 0.00332954f $X=1.945 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_308 N_A_43_69#_c_532_n N_A_298_69#_c_561_n 0.0133061f $X=1.945 $Y=0.955 $X2=0
+ $Y2=0
cc_309 N_A_43_69#_M1011_s N_A_298_69#_c_559_n 0.0033329f $X=1.92 $Y=0.345 $X2=0
+ $Y2=0
cc_310 N_A_43_69#_c_532_n N_A_298_69#_c_559_n 0.00447792f $X=1.945 $Y=0.955
+ $X2=0 $Y2=0
cc_311 N_A_43_69#_c_526_n N_A_298_69#_c_559_n 0.022529f $X=2.11 $Y=0.68 $X2=0
+ $Y2=0
cc_312 N_A_43_69#_c_524_n N_A_298_69#_c_560_n 0.00833305f $X=1.115 $Y=0.34 $X2=0
+ $Y2=0
cc_313 N_A_43_69#_c_526_n N_A_522_47#_c_585_n 0.0143382f $X=2.11 $Y=0.68 $X2=0
+ $Y2=0
cc_314 N_A_43_69#_c_524_n N_VGND_c_632_n 0.0586439f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_315 N_A_43_69#_c_525_n N_VGND_c_632_n 0.0186386f $X=0.435 $Y=0.34 $X2=0 $Y2=0
cc_316 N_A_43_69#_c_524_n N_VGND_c_634_n 0.0327464f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_317 N_A_43_69#_c_525_n N_VGND_c_634_n 0.0101082f $X=0.435 $Y=0.34 $X2=0 $Y2=0
cc_318 N_A_298_69#_c_559_n N_A_522_47#_M1005_s 0.00585625f $X=3 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_319 N_A_298_69#_M1005_d N_A_522_47#_c_585_n 0.00330588f $X=3.025 $Y=0.235
+ $X2=0 $Y2=0
cc_320 N_A_298_69#_c_559_n N_A_522_47#_c_585_n 0.0137436f $X=3 $Y=0.34 $X2=0
+ $Y2=0
cc_321 N_A_298_69#_c_566_n N_A_522_47#_c_585_n 0.0160969f $X=3.165 $Y=0.34 $X2=0
+ $Y2=0
cc_322 N_A_298_69#_c_559_n N_VGND_c_632_n 0.0762241f $X=3 $Y=0.34 $X2=0 $Y2=0
cc_323 N_A_298_69#_c_560_n N_VGND_c_632_n 0.0187393f $X=1.775 $Y=0.34 $X2=0
+ $Y2=0
cc_324 N_A_298_69#_c_566_n N_VGND_c_632_n 0.0182958f $X=3.165 $Y=0.34 $X2=0
+ $Y2=0
cc_325 N_A_298_69#_M1005_d N_VGND_c_634_n 0.00225167f $X=3.025 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_298_69#_c_559_n N_VGND_c_634_n 0.0448252f $X=3 $Y=0.34 $X2=0 $Y2=0
cc_327 N_A_298_69#_c_560_n N_VGND_c_634_n 0.0103621f $X=1.775 $Y=0.34 $X2=0
+ $Y2=0
cc_328 N_A_298_69#_c_566_n N_VGND_c_634_n 0.0123228f $X=3.165 $Y=0.34 $X2=0
+ $Y2=0
cc_329 N_A_522_47#_c_593_n N_VGND_M1004_d 0.00328155f $X=4.36 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_330 N_A_522_47#_c_597_n N_VGND_M1002_d 0.00363794f $X=5.22 $Y=0.93 $X2=0
+ $Y2=0
cc_331 N_A_522_47#_c_593_n N_VGND_c_628_n 0.016709f $X=4.36 $Y=0.93 $X2=0 $Y2=0
cc_332 N_A_522_47#_c_597_n N_VGND_c_629_n 0.016709f $X=5.22 $Y=0.93 $X2=0 $Y2=0
cc_333 N_A_522_47#_c_615_p N_VGND_c_630_n 0.0124525f $X=4.455 $Y=0.42 $X2=0
+ $Y2=0
cc_334 N_A_522_47#_c_616_p N_VGND_c_632_n 0.0124525f $X=3.595 $Y=0.42 $X2=0
+ $Y2=0
cc_335 N_A_522_47#_c_587_n N_VGND_c_633_n 0.0178111f $X=5.315 $Y=0.42 $X2=0
+ $Y2=0
cc_336 N_A_522_47#_M1005_s N_VGND_c_634_n 0.0021598f $X=2.61 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_A_522_47#_M1017_s N_VGND_c_634_n 0.00276363f $X=3.455 $Y=0.235 $X2=0
+ $Y2=0
cc_338 N_A_522_47#_M1013_s N_VGND_c_634_n 0.00280978f $X=4.315 $Y=0.235 $X2=0
+ $Y2=0
cc_339 N_A_522_47#_M1008_s N_VGND_c_634_n 0.00243868f $X=5.175 $Y=0.235 $X2=0
+ $Y2=0
cc_340 N_A_522_47#_c_585_n N_VGND_c_634_n 0.00730497f $X=3.5 $Y=0.895 $X2=0
+ $Y2=0
cc_341 N_A_522_47#_c_616_p N_VGND_c_634_n 0.00730901f $X=3.595 $Y=0.42 $X2=0
+ $Y2=0
cc_342 N_A_522_47#_c_593_n N_VGND_c_634_n 0.0108383f $X=4.36 $Y=0.93 $X2=0 $Y2=0
cc_343 N_A_522_47#_c_615_p N_VGND_c_634_n 0.00730901f $X=4.455 $Y=0.42 $X2=0
+ $Y2=0
cc_344 N_A_522_47#_c_597_n N_VGND_c_634_n 0.0108383f $X=5.22 $Y=0.93 $X2=0 $Y2=0
cc_345 N_A_522_47#_c_587_n N_VGND_c_634_n 0.0100304f $X=5.315 $Y=0.42 $X2=0
+ $Y2=0
