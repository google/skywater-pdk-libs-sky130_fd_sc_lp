* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ha_2 A B VGND VNB VPB VPWR COUT SUM
X0 a_227_397# a_270_95# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_45_121# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A a_155_397# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 COUT a_270_95# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 COUT a_270_95# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND a_227_397# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR a_270_95# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 SUM a_227_397# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND B a_45_121# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_227_397# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 SUM a_227_397# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_155_397# B a_227_397# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_270_95# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VPWR B a_270_95# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_492_131# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_45_121# a_270_95# a_227_397# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_270_95# B a_492_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_270_95# COUT VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
