* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_921_65# A3 a_1291_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_1291_65# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_30_367# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_478_65# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR A4 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A4 a_1291_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Y A1 a_478_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_921_65# A2 a_478_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_1291_65# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_30_367# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR A2 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_921_65# A2 a_478_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_1291_65# A3 a_921_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR A1 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VPWR A1 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR A4 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_921_65# A3 a_1291_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 Y A1 a_478_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 Y B1 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_30_367# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_478_65# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 VPWR A3 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VGND A4 a_1291_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_30_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_30_367# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VPWR A2 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_30_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 VPWR A3 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_30_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_30_367# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_30_367# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_478_65# A2 a_921_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 Y B1 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 a_30_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 a_478_65# A2 a_921_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 a_1291_65# A3 a_921_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
