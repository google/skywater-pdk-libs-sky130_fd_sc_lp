* File: sky130_fd_sc_lp__o31ai_0.pxi.spice
* Created: Fri Aug 28 11:16:13 2020
* 
x_PM_SKY130_FD_SC_LP__O31AI_0%A1 N_A1_c_64_n N_A1_c_65_n N_A1_M1006_g
+ N_A1_c_71_n N_A1_M1000_g N_A1_c_66_n N_A1_c_67_n N_A1_c_72_n A1 A1 A1 A1
+ N_A1_c_69_n PM_SKY130_FD_SC_LP__O31AI_0%A1
x_PM_SKY130_FD_SC_LP__O31AI_0%A2 N_A2_c_104_n N_A2_M1007_g N_A2_M1001_g
+ N_A2_c_110_n A2 A2 A2 N_A2_c_107_n PM_SKY130_FD_SC_LP__O31AI_0%A2
x_PM_SKY130_FD_SC_LP__O31AI_0%A3 N_A3_M1005_g N_A3_M1002_g N_A3_c_155_n
+ N_A3_c_156_n A3 A3 N_A3_c_157_n N_A3_c_158_n PM_SKY130_FD_SC_LP__O31AI_0%A3
x_PM_SKY130_FD_SC_LP__O31AI_0%B1 N_B1_M1003_g N_B1_M1004_g N_B1_c_196_n
+ N_B1_c_197_n N_B1_c_204_n N_B1_c_198_n B1 B1 B1 N_B1_c_200_n N_B1_c_201_n
+ PM_SKY130_FD_SC_LP__O31AI_0%B1
x_PM_SKY130_FD_SC_LP__O31AI_0%VPWR N_VPWR_M1000_s N_VPWR_M1003_d N_VPWR_c_242_n
+ N_VPWR_c_243_n N_VPWR_c_244_n N_VPWR_c_245_n VPWR N_VPWR_c_246_n
+ N_VPWR_c_247_n N_VPWR_c_241_n N_VPWR_c_249_n PM_SKY130_FD_SC_LP__O31AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O31AI_0%Y N_Y_M1004_d N_Y_M1005_d N_Y_c_271_n N_Y_c_272_n
+ N_Y_c_291_n Y Y Y Y Y Y Y N_Y_c_270_n N_Y_c_275_n
+ PM_SKY130_FD_SC_LP__O31AI_0%Y
x_PM_SKY130_FD_SC_LP__O31AI_0%VGND N_VGND_M1006_s N_VGND_M1007_d N_VGND_c_309_n
+ N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n VGND N_VGND_c_313_n
+ N_VGND_c_314_n N_VGND_c_315_n PM_SKY130_FD_SC_LP__O31AI_0%VGND
x_PM_SKY130_FD_SC_LP__O31AI_0%A_138_65# N_A_138_65#_M1006_d N_A_138_65#_M1002_d
+ N_A_138_65#_c_341_n N_A_138_65#_c_342_n N_A_138_65#_c_343_n
+ N_A_138_65#_c_353_n PM_SKY130_FD_SC_LP__O31AI_0%A_138_65#
cc_1 VNB N_A1_c_64_n 0.00799077f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.155
cc_2 VNB N_A1_c_65_n 0.0214842f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.855
cc_3 VNB N_A1_c_66_n 0.038165f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.93
cc_4 VNB N_A1_c_67_n 0.0185672f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_5 VNB A1 0.0350324f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A1_c_69_n 0.0285686f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_7 VNB N_A2_c_104_n 0.0143645f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.155
cc_8 VNB N_A2_M1007_g 0.0394448f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.535
cc_9 VNB A2 0.00852003f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.93
cc_10 VNB N_A2_c_107_n 0.0252189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_M1002_g 0.0306653f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.735
cc_12 VNB N_A3_c_155_n 0.0218141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A3_c_156_n 0.00290425f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.93
cc_14 VNB N_A3_c_157_n 0.0157595f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.23
cc_15 VNB N_A3_c_158_n 0.00715745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_196_n 0.0229887f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.93
cc_17 VNB N_B1_c_197_n 0.00798402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_198_n 0.023686f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.23
cc_19 VNB B1 0.0028878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_200_n 0.0236289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_201_n 0.0214281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_241_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB Y 0.0552687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_270_n 0.0156072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_309_n 0.0155138f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.735
cc_26 VNB N_VGND_c_310_n 0.0206562f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.93
cc_27 VNB N_VGND_c_311_n 0.0161299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_312_n 0.00763253f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_29 VNB N_VGND_c_313_n 0.0391991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_314_n 0.182327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_315_n 0.00632158f $X=-0.19 $Y=-0.245 $X2=0.247 $Y2=0.925
cc_32 VNB N_A_138_65#_c_341_n 2.02372e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.93
cc_33 VNB N_A_138_65#_c_342_n 0.0165925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_138_65#_c_343_n 0.00342974f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.93
cc_35 VPB N_A1_c_64_n 0.0307009f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.155
cc_36 VPB N_A1_c_71_n 0.0208289f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.305
cc_37 VPB N_A1_c_72_n 0.0325993f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.23
cc_38 VPB A1 0.0293914f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_39 VPB N_A2_c_104_n 0.00284218f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.155
cc_40 VPB N_A2_M1001_g 0.0372143f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.93
cc_41 VPB N_A2_c_110_n 0.0245559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB A2 0.0130905f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.93
cc_43 VPB N_A3_M1005_g 0.0428426f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.855
cc_44 VPB N_A3_c_156_n 0.0128819f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.93
cc_45 VPB N_A3_c_158_n 0.00427395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B1_M1003_g 0.0304706f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.855
cc_47 VPB N_B1_c_197_n 0.0229891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B1_c_204_n 0.0188689f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.36
cc_49 VPB B1 0.00306061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_242_n 0.0330415f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.93
cc_51 VPB N_VPWR_c_243_n 0.0343622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_244_n 0.0108943f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.23
cc_53 VPB N_VPWR_c_245_n 0.00541171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_246_n 0.0400413f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_55 VPB N_VPWR_c_247_n 0.0223503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_241_n 0.0963799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_249_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_Y_c_271_n 0.0196844f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.735
cc_59 VPB N_Y_c_272_n 0.00229315f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.735
cc_60 VPB Y 0.00207453f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.36
cc_61 VPB Y 0.0196589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_Y_c_275_n 0.0280698f $X=-0.19 $Y=1.655 $X2=0.247 $Y2=1.665
cc_63 N_A1_c_67_n N_A2_c_104_n 0.0113397f $X=0.27 $Y=1.525 $X2=0 $Y2=0
cc_64 N_A1_c_65_n N_A2_M1007_g 0.0185935f $X=0.615 $Y=0.855 $X2=0 $Y2=0
cc_65 A1 N_A2_M1007_g 0.00176932f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_A1_c_69_n N_A2_M1007_g 0.00269168f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_67 N_A1_c_64_n N_A2_M1001_g 0.00226037f $X=0.36 $Y=2.155 $X2=0 $Y2=0
cc_68 N_A1_c_72_n N_A2_M1001_g 0.0569912f $X=0.655 $Y=2.23 $X2=0 $Y2=0
cc_69 A1 N_A2_M1001_g 3.49144e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_A1_c_64_n N_A2_c_110_n 0.0113397f $X=0.36 $Y=2.155 $X2=0 $Y2=0
cc_71 N_A1_c_72_n N_A2_c_110_n 0.00304845f $X=0.655 $Y=2.23 $X2=0 $Y2=0
cc_72 N_A1_c_66_n A2 0.00522513f $X=0.615 $Y=0.93 $X2=0 $Y2=0
cc_73 N_A1_c_72_n A2 0.0125145f $X=0.655 $Y=2.23 $X2=0 $Y2=0
cc_74 A1 A2 0.0879284f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_A1_c_69_n A2 0.00662003f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_76 N_A1_c_66_n N_A2_c_107_n 8.34398e-19 $X=0.615 $Y=0.93 $X2=0 $Y2=0
cc_77 A1 N_A2_c_107_n 6.75732e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A1_c_69_n N_A2_c_107_n 0.0113397f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_79 N_A1_c_71_n N_VPWR_c_242_n 0.018148f $X=0.655 $Y=2.305 $X2=0 $Y2=0
cc_80 N_A1_c_72_n N_VPWR_c_242_n 0.01159f $X=0.655 $Y=2.23 $X2=0 $Y2=0
cc_81 A1 N_VPWR_c_242_n 0.0118973f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_82 N_A1_c_71_n N_VPWR_c_246_n 0.00452967f $X=0.655 $Y=2.305 $X2=0 $Y2=0
cc_83 N_A1_c_71_n N_VPWR_c_241_n 0.00809218f $X=0.655 $Y=2.305 $X2=0 $Y2=0
cc_84 N_A1_c_65_n N_VGND_c_310_n 0.0105043f $X=0.615 $Y=0.855 $X2=0 $Y2=0
cc_85 N_A1_c_66_n N_VGND_c_310_n 0.00542545f $X=0.615 $Y=0.93 $X2=0 $Y2=0
cc_86 A1 N_VGND_c_310_n 0.0155813f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A1_c_65_n N_VGND_c_311_n 0.00414769f $X=0.615 $Y=0.855 $X2=0 $Y2=0
cc_88 N_A1_c_65_n N_VGND_c_314_n 0.0078848f $X=0.615 $Y=0.855 $X2=0 $Y2=0
cc_89 A1 N_VGND_c_314_n 0.00654415f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A1_c_65_n N_A_138_65#_c_341_n 5.37715e-19 $X=0.615 $Y=0.855 $X2=0 $Y2=0
cc_91 N_A1_c_65_n N_A_138_65#_c_343_n 0.00360072f $X=0.615 $Y=0.855 $X2=0 $Y2=0
cc_92 A1 N_A_138_65#_c_343_n 0.00499902f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A2_c_110_n N_A3_M1005_g 0.0277519f $X=0.897 $Y=1.915 $X2=0 $Y2=0
cc_94 N_A2_M1007_g N_A3_M1002_g 0.0174511f $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_95 N_A2_c_107_n N_A3_c_155_n 0.0277519f $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A2_c_104_n N_A3_c_156_n 0.0277519f $X=0.897 $Y=1.693 $X2=0 $Y2=0
cc_97 N_A2_M1007_g N_A3_c_157_n 0.0277519f $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_98 A2 N_A3_c_157_n 0.00363202f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A2_M1007_g N_A3_c_158_n 0.00289068f $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_100 A2 N_A3_c_158_n 0.0297701f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A2_M1001_g N_VPWR_c_242_n 0.00423267f $X=1.045 $Y=2.735 $X2=0 $Y2=0
cc_102 A2 N_VPWR_c_242_n 0.00194697f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A2_M1001_g N_VPWR_c_246_n 0.00545548f $X=1.045 $Y=2.735 $X2=0 $Y2=0
cc_104 N_A2_M1001_g N_VPWR_c_241_n 0.0104231f $X=1.045 $Y=2.735 $X2=0 $Y2=0
cc_105 N_A2_M1001_g N_Y_c_272_n 6.87277e-19 $X=1.045 $Y=2.735 $X2=0 $Y2=0
cc_106 A2 N_Y_c_272_n 0.00853699f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A2_M1001_g Y 0.00416087f $X=1.045 $Y=2.735 $X2=0 $Y2=0
cc_108 N_A2_M1007_g N_VGND_c_310_n 4.80864e-19 $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_109 N_A2_M1007_g N_VGND_c_311_n 0.00494765f $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_110 N_A2_M1007_g N_VGND_c_312_n 0.00188929f $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_111 N_A2_M1007_g N_VGND_c_314_n 0.00513371f $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_112 N_A2_M1007_g N_A_138_65#_c_341_n 0.00549053f $X=1.045 $Y=0.535 $X2=0
+ $Y2=0
cc_113 N_A2_M1007_g N_A_138_65#_c_342_n 0.0134006f $X=1.045 $Y=0.535 $X2=0 $Y2=0
cc_114 A2 N_A_138_65#_c_342_n 0.00194751f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A2_M1007_g N_A_138_65#_c_343_n 0.00165559f $X=1.045 $Y=0.535 $X2=0
+ $Y2=0
cc_116 A2 N_A_138_65#_c_343_n 0.0200718f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A2_c_107_n N_A_138_65#_c_343_n 0.00135248f $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A2_M1007_g N_A_138_65#_c_353_n 3.53389e-19 $X=1.045 $Y=0.535 $X2=0
+ $Y2=0
cc_119 N_A3_c_157_n N_B1_c_196_n 0.0114215f $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_120 N_A3_c_158_n N_B1_c_196_n 0.00582975f $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_121 N_A3_M1005_g N_B1_c_197_n 0.00763827f $X=1.435 $Y=2.735 $X2=0 $Y2=0
cc_122 N_A3_c_156_n N_B1_c_197_n 0.0114215f $X=1.525 $Y=1.775 $X2=0 $Y2=0
cc_123 N_A3_M1005_g N_B1_c_204_n 0.024421f $X=1.435 $Y=2.735 $X2=0 $Y2=0
cc_124 N_A3_c_158_n N_B1_c_204_n 7.58098e-19 $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_125 N_A3_c_155_n N_B1_c_198_n 0.0114215f $X=1.525 $Y=1.61 $X2=0 $Y2=0
cc_126 N_A3_M1002_g B1 8.83339e-19 $X=1.575 $Y=0.535 $X2=0 $Y2=0
cc_127 N_A3_c_157_n B1 4.88354e-19 $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_128 N_A3_c_158_n B1 0.0557887f $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_129 N_A3_M1002_g N_B1_c_201_n 0.0236889f $X=1.575 $Y=0.535 $X2=0 $Y2=0
cc_130 N_A3_M1005_g N_VPWR_c_246_n 0.00511657f $X=1.435 $Y=2.735 $X2=0 $Y2=0
cc_131 N_A3_M1005_g N_VPWR_c_241_n 0.00961146f $X=1.435 $Y=2.735 $X2=0 $Y2=0
cc_132 N_A3_c_158_n N_Y_c_271_n 0.00682166f $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_133 N_A3_M1005_g N_Y_c_272_n 0.00741973f $X=1.435 $Y=2.735 $X2=0 $Y2=0
cc_134 N_A3_c_156_n N_Y_c_272_n 0.00127981f $X=1.525 $Y=1.775 $X2=0 $Y2=0
cc_135 N_A3_c_158_n N_Y_c_272_n 0.0307745f $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_136 N_A3_M1005_g Y 0.0173623f $X=1.435 $Y=2.735 $X2=0 $Y2=0
cc_137 N_A3_M1002_g N_VGND_c_312_n 0.00354727f $X=1.575 $Y=0.535 $X2=0 $Y2=0
cc_138 N_A3_M1002_g N_VGND_c_313_n 0.00494765f $X=1.575 $Y=0.535 $X2=0 $Y2=0
cc_139 N_A3_M1002_g N_VGND_c_314_n 0.00513371f $X=1.575 $Y=0.535 $X2=0 $Y2=0
cc_140 N_A3_M1002_g N_A_138_65#_c_341_n 3.53562e-19 $X=1.575 $Y=0.535 $X2=0
+ $Y2=0
cc_141 N_A3_M1002_g N_A_138_65#_c_342_n 0.0115123f $X=1.575 $Y=0.535 $X2=0 $Y2=0
cc_142 N_A3_c_157_n N_A_138_65#_c_342_n 0.00127342f $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_143 N_A3_c_158_n N_A_138_65#_c_342_n 0.0450331f $X=1.525 $Y=1.27 $X2=0 $Y2=0
cc_144 N_A3_M1002_g N_A_138_65#_c_353_n 0.00549696f $X=1.575 $Y=0.535 $X2=0
+ $Y2=0
cc_145 N_B1_M1003_g N_VPWR_c_243_n 0.0049642f $X=1.865 $Y=2.735 $X2=0 $Y2=0
cc_146 N_B1_c_204_n N_VPWR_c_243_n 6.28929e-19 $X=2.005 $Y=2.09 $X2=0 $Y2=0
cc_147 N_B1_M1003_g N_VPWR_c_246_n 0.00511657f $X=1.865 $Y=2.735 $X2=0 $Y2=0
cc_148 N_B1_M1003_g N_VPWR_c_241_n 0.0105216f $X=1.865 $Y=2.735 $X2=0 $Y2=0
cc_149 N_B1_M1003_g N_Y_c_271_n 0.00779587f $X=1.865 $Y=2.735 $X2=0 $Y2=0
cc_150 N_B1_c_197_n N_Y_c_271_n 0.00824348f $X=2.005 $Y=2.015 $X2=0 $Y2=0
cc_151 N_B1_c_204_n N_Y_c_271_n 0.0111065f $X=2.005 $Y=2.09 $X2=0 $Y2=0
cc_152 N_B1_c_198_n N_Y_c_271_n 0.00290723f $X=2.127 $Y=1.525 $X2=0 $Y2=0
cc_153 B1 N_Y_c_271_n 0.0161653f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_154 N_B1_M1003_g N_Y_c_272_n 8.27236e-19 $X=1.865 $Y=2.735 $X2=0 $Y2=0
cc_155 N_B1_c_204_n N_Y_c_272_n 0.00248749f $X=2.005 $Y=2.09 $X2=0 $Y2=0
cc_156 B1 N_Y_c_291_n 0.0134831f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_157 N_B1_c_200_n N_Y_c_291_n 0.00415211f $X=2.16 $Y=1.02 $X2=0 $Y2=0
cc_158 N_B1_c_201_n N_Y_c_291_n 0.00367435f $X=2.127 $Y=0.855 $X2=0 $Y2=0
cc_159 N_B1_M1003_g Y 0.016973f $X=1.865 $Y=2.735 $X2=0 $Y2=0
cc_160 N_B1_c_197_n Y 0.00670685f $X=2.005 $Y=2.015 $X2=0 $Y2=0
cc_161 B1 Y 0.075505f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_162 N_B1_c_200_n Y 0.0172096f $X=2.16 $Y=1.02 $X2=0 $Y2=0
cc_163 N_B1_c_201_n Y 0.0029062f $X=2.127 $Y=0.855 $X2=0 $Y2=0
cc_164 N_B1_c_201_n N_VGND_c_313_n 0.00481189f $X=2.127 $Y=0.855 $X2=0 $Y2=0
cc_165 N_B1_c_201_n N_VGND_c_314_n 0.00985463f $X=2.127 $Y=0.855 $X2=0 $Y2=0
cc_166 B1 N_A_138_65#_c_342_n 0.00768488f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_167 N_B1_c_201_n N_A_138_65#_c_342_n 0.00201642f $X=2.127 $Y=0.855 $X2=0
+ $Y2=0
cc_168 N_B1_c_201_n N_A_138_65#_c_353_n 3.04752e-19 $X=2.127 $Y=0.855 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_243_n N_Y_c_271_n 0.0223462f $X=2.08 $Y=2.56 $X2=0 $Y2=0
cc_170 N_VPWR_c_243_n Y 0.0262636f $X=2.08 $Y=2.56 $X2=0 $Y2=0
cc_171 N_VPWR_c_246_n Y 0.021949f $X=1.985 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_241_n Y 0.0124703f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_173 N_Y_c_291_n N_VGND_c_313_n 0.0142842f $X=2.425 $Y=0.505 $X2=0 $Y2=0
cc_174 N_Y_c_270_n N_VGND_c_313_n 0.0166501f $X=2.607 $Y=0.67 $X2=0 $Y2=0
cc_175 N_Y_c_291_n N_VGND_c_314_n 0.0129745f $X=2.425 $Y=0.505 $X2=0 $Y2=0
cc_176 N_Y_c_270_n N_VGND_c_314_n 0.0135611f $X=2.607 $Y=0.67 $X2=0 $Y2=0
cc_177 Y N_A_138_65#_c_342_n 0.00300709f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_178 Y N_A_138_65#_c_353_n 0.00199941f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_179 N_VGND_c_311_n N_A_138_65#_c_341_n 0.00816195f $X=1.145 $Y=0 $X2=0 $Y2=0
cc_180 N_VGND_c_314_n N_A_138_65#_c_341_n 0.00859584f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_181 N_VGND_c_312_n N_A_138_65#_c_342_n 0.0235363f $X=1.31 $Y=0.49 $X2=0 $Y2=0
cc_182 N_VGND_c_314_n N_A_138_65#_c_342_n 0.0116672f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_183 N_VGND_c_313_n N_A_138_65#_c_353_n 0.00837508f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_184 N_VGND_c_314_n N_A_138_65#_c_353_n 0.00895833f $X=2.64 $Y=0 $X2=0 $Y2=0
