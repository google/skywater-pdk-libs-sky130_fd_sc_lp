* NGSPICE file created from sky130_fd_sc_lp__o31a_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VGND A2 a_355_47# VNB nshort w=840000u l=150000u
+  ad=9.786e+11p pd=7.37e+06u as=5.964e+11p ps=4.78e+06u
M1001 a_355_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=1.4364e+12p ps=9.84e+06u
M1002 VPWR a_85_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1003 a_85_21# B1 a_355_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1004 a_355_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_85_21# A3 a_427_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.914e+11p pd=3.3e+06u as=4.914e+11p ps=3.3e+06u
M1006 a_427_367# A2 a_355_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_355_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_85_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B1 a_85_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_85_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1011 X a_85_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

