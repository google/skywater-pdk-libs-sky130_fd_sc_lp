* File: sky130_fd_sc_lp__srdlstp_1.pxi.spice
* Created: Fri Aug 28 11:33:10 2020
* 
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%D N_D_c_231_n N_D_M1024_g N_D_M1028_g
+ N_D_c_234_n D D N_D_c_235_n N_D_c_236_n PM_SKY130_FD_SC_LP__SRDLSTP_1%D
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_27_400# N_A_27_400#_M1024_d
+ N_A_27_400#_M1028_s N_A_27_400#_M1005_g N_A_27_400#_c_265_n
+ N_A_27_400#_M1031_g N_A_27_400#_c_272_n N_A_27_400#_c_267_n
+ N_A_27_400#_c_273_n N_A_27_400#_c_274_n N_A_27_400#_c_268_n
+ N_A_27_400#_c_269_n N_A_27_400#_c_270_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%A_27_400#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%SET_B N_SET_B_c_332_n N_SET_B_M1025_g
+ N_SET_B_c_333_n N_SET_B_M1026_g N_SET_B_M1011_g N_SET_B_c_336_n
+ N_SET_B_c_337_n N_SET_B_c_338_n N_SET_B_c_339_n N_SET_B_c_340_n SET_B
+ N_SET_B_c_342_n PM_SKY130_FD_SC_LP__SRDLSTP_1%SET_B
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_404_353# N_A_404_353#_M1013_s
+ N_A_404_353#_M1007_d N_A_404_353#_c_431_n N_A_404_353#_M1010_g
+ N_A_404_353#_M1034_g N_A_404_353#_c_433_n N_A_404_353#_c_434_n
+ N_A_404_353#_M1033_g N_A_404_353#_M1030_g N_A_404_353#_M1029_g
+ N_A_404_353#_c_437_n N_A_404_353#_c_454_p N_A_404_353#_c_559_p
+ N_A_404_353#_c_422_n N_A_404_353#_c_455_p N_A_404_353#_c_439_n
+ N_A_404_353#_c_423_n N_A_404_353#_c_424_n N_A_404_353#_c_425_n
+ N_A_404_353#_c_426_n N_A_404_353#_c_442_n N_A_404_353#_c_443_n
+ N_A_404_353#_c_427_n N_A_404_353#_c_428_n N_A_404_353#_c_458_p
+ N_A_404_353#_c_429_n N_A_404_353#_c_430_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%A_404_353#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_434_405# N_A_434_405#_M1034_d
+ N_A_434_405#_M1010_d N_A_434_405#_c_618_n N_A_434_405#_M1019_g
+ N_A_434_405#_c_619_n N_A_434_405#_M1021_g N_A_434_405#_c_621_n
+ N_A_434_405#_M1014_g N_A_434_405#_c_622_n N_A_434_405#_c_623_n
+ N_A_434_405#_c_624_n N_A_434_405#_c_625_n N_A_434_405#_c_626_n
+ N_A_434_405#_c_633_n N_A_434_405#_c_627_n N_A_434_405#_c_628_n
+ N_A_434_405#_c_629_n PM_SKY130_FD_SC_LP__SRDLSTP_1%A_434_405#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_878_357# N_A_878_357#_M1006_d
+ N_A_878_357#_M1009_d N_A_878_357#_M1000_g N_A_878_357#_c_714_n
+ N_A_878_357#_M1012_g N_A_878_357#_c_715_n N_A_878_357#_c_716_n
+ N_A_878_357#_c_717_n N_A_878_357#_M1016_g N_A_878_357#_c_718_n
+ N_A_878_357#_c_719_n N_A_878_357#_c_725_n N_A_878_357#_c_720_n
+ N_A_878_357#_c_727_n N_A_878_357#_c_728_n N_A_878_357#_c_721_n
+ N_A_878_357#_c_722_n N_A_878_357#_c_729_n N_A_878_357#_c_723_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%A_878_357#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_1294_315# N_A_1294_315#_M1023_s
+ N_A_1294_315#_M1001_d N_A_1294_315#_M1002_g N_A_1294_315#_c_823_n
+ N_A_1294_315#_M1020_g N_A_1294_315#_c_829_n N_A_1294_315#_c_830_n
+ N_A_1294_315#_c_831_n N_A_1294_315#_c_832_n N_A_1294_315#_c_833_n
+ N_A_1294_315#_c_825_n N_A_1294_315#_c_835_n N_A_1294_315#_c_836_n
+ N_A_1294_315#_c_837_n N_A_1294_315#_c_826_n N_A_1294_315#_c_868_p
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%A_1294_315#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%GATE N_GATE_c_923_n N_GATE_c_924_n
+ N_GATE_M1007_g N_GATE_M1013_g N_GATE_c_927_n GATE GATE N_GATE_c_929_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%GATE
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%SLEEP_B N_SLEEP_B_M1004_g N_SLEEP_B_M1003_g
+ N_SLEEP_B_M1032_g N_SLEEP_B_c_970_n N_SLEEP_B_c_971_n N_SLEEP_B_M1001_g
+ N_SLEEP_B_c_973_n N_SLEEP_B_M1023_g N_SLEEP_B_M1015_g N_SLEEP_B_c_976_n
+ N_SLEEP_B_c_977_n SLEEP_B SLEEP_B N_SLEEP_B_c_978_n N_SLEEP_B_c_979_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%SLEEP_B
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_700_451# N_A_700_451#_M1021_d
+ N_A_700_451#_M1030_d N_A_700_451#_M1026_s N_A_700_451#_M1022_g
+ N_A_700_451#_M1009_g N_A_700_451#_c_1039_n N_A_700_451#_c_1040_n
+ N_A_700_451#_c_1041_n N_A_700_451#_M1006_g N_A_700_451#_M1017_g
+ N_A_700_451#_M1027_g N_A_700_451#_c_1045_n N_A_700_451#_c_1056_n
+ N_A_700_451#_c_1082_n N_A_700_451#_c_1065_n N_A_700_451#_c_1046_n
+ N_A_700_451#_c_1047_n N_A_700_451#_c_1048_n N_A_700_451#_c_1049_n
+ N_A_700_451#_c_1050_n N_A_700_451#_c_1058_n N_A_700_451#_c_1059_n
+ N_A_700_451#_c_1051_n N_A_700_451#_c_1061_n N_A_700_451#_c_1052_n
+ N_A_700_451#_c_1053_n PM_SKY130_FD_SC_LP__SRDLSTP_1%A_700_451#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_2266_367# N_A_2266_367#_M1017_d
+ N_A_2266_367#_M1027_s N_A_2266_367#_M1008_g N_A_2266_367#_M1018_g
+ N_A_2266_367#_c_1223_n N_A_2266_367#_c_1224_n N_A_2266_367#_c_1229_n
+ N_A_2266_367#_c_1225_n N_A_2266_367#_c_1226_n N_A_2266_367#_c_1227_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%A_2266_367#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%VPWR N_VPWR_M1028_d N_VPWR_M1010_s
+ N_VPWR_M1027_d N_VPWR_c_1265_n N_VPWR_c_1266_n N_VPWR_c_1267_n N_VPWR_c_1268_n
+ VPWR N_VPWR_c_1269_n N_VPWR_c_1270_n N_VPWR_c_1264_n N_VPWR_c_1272_n
+ N_VPWR_c_1273_n N_VPWR_c_1274_n PM_SKY130_FD_SC_LP__SRDLSTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_217_130# N_A_217_130#_M1031_s
+ N_A_217_130#_M1019_s N_A_217_130#_M1005_d N_A_217_130#_M1033_s
+ N_A_217_130#_c_1362_n N_A_217_130#_c_1370_n N_A_217_130#_c_1371_n
+ N_A_217_130#_c_1372_n N_A_217_130#_c_1373_n N_A_217_130#_c_1363_n
+ N_A_217_130#_c_1364_n N_A_217_130#_c_1365_n N_A_217_130#_c_1366_n
+ N_A_217_130#_c_1367_n N_A_217_130#_c_1368_n N_A_217_130#_c_1375_n
+ N_A_217_130#_c_1369_n N_A_217_130#_c_1377_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%A_217_130#
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%KAPWR N_KAPWR_M1000_d N_KAPWR_M1002_d
+ N_KAPWR_M1007_s N_KAPWR_M1003_d KAPWR N_KAPWR_c_1479_n N_KAPWR_c_1480_n
+ N_KAPWR_c_1481_n N_KAPWR_c_1482_n N_KAPWR_c_1483_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%KAPWR
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%Q N_Q_M1008_d N_Q_M1018_d Q Q Q Q Q N_Q_c_1576_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%Q
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%VGND N_VGND_M1024_s N_VGND_M1025_d
+ N_VGND_M1011_s N_VGND_M1020_d N_VGND_M1032_d N_VGND_M1015_d N_VGND_M1008_s
+ N_VGND_c_1590_n N_VGND_c_1591_n N_VGND_c_1592_n N_VGND_c_1593_n
+ N_VGND_c_1594_n N_VGND_c_1595_n N_VGND_c_1596_n N_VGND_c_1597_n
+ N_VGND_c_1598_n N_VGND_c_1599_n N_VGND_c_1600_n VGND N_VGND_c_1601_n
+ N_VGND_c_1602_n N_VGND_c_1603_n N_VGND_c_1604_n N_VGND_c_1605_n
+ N_VGND_c_1606_n N_VGND_c_1607_n N_VGND_c_1608_n N_VGND_c_1609_n
+ N_VGND_c_1610_n N_VGND_c_1611_n N_VGND_c_1612_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%VGND
x_PM_SKY130_FD_SC_LP__SRDLSTP_1%A_988_47# N_A_988_47#_M1016_d
+ N_A_988_47#_M1011_d N_A_988_47#_c_1744_n N_A_988_47#_c_1745_n
+ N_A_988_47#_c_1746_n N_A_988_47#_c_1747_n N_A_988_47#_c_1748_n
+ PM_SKY130_FD_SC_LP__SRDLSTP_1%A_988_47#
cc_1 VNB N_D_c_231_n 0.0287713f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.408
cc_2 VNB N_D_M1024_g 0.0312678f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_3 VNB N_D_M1028_g 0.00179598f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.32
cc_4 VNB N_D_c_234_n 0.0338436f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.625
cc_5 VNB N_D_c_235_n 0.0347636f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_6 VNB N_D_c_236_n 0.00544187f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_7 VNB N_A_27_400#_c_265_n 0.0276363f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.625
cc_8 VNB N_A_27_400#_M1031_g 0.0257198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_400#_c_267_n 0.0139676f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_10 VNB N_A_27_400#_c_268_n 0.0181952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_400#_c_269_n 0.0017057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_400#_c_270_n 0.0227557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SET_B_c_332_n 0.0237193f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.172
cc_14 VNB N_SET_B_c_333_n 0.0450856f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_15 VNB N_SET_B_M1026_g 0.00655175f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.32
cc_16 VNB N_SET_B_M1011_g 0.0227668f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_SET_B_c_336_n 0.0190174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SET_B_c_337_n 0.019639f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.12
cc_19 VNB N_SET_B_c_338_n 0.0170601f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_20 VNB N_SET_B_c_339_n 0.054288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SET_B_c_340_n 0.00182751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB SET_B 0.00885596f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_23 VNB N_SET_B_c_342_n 0.0419666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_404_353#_M1034_g 0.0394102f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB N_A_404_353#_M1029_g 0.0359227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_404_353#_c_422_n 0.00398045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_404_353#_c_423_n 0.011399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_404_353#_c_424_n 0.00362546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_404_353#_c_425_n 0.00349508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_404_353#_c_426_n 0.00492046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_404_353#_c_427_n 0.00572626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_404_353#_c_428_n 0.039213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_404_353#_c_429_n 0.0180514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_404_353#_c_430_n 0.00937817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_434_405#_c_618_n 0.0187875f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.625
cc_36 VNB N_A_434_405#_c_619_n 0.0102122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_434_405#_M1021_g 0.0243005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_434_405#_c_621_n 0.0131843f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_39 VNB N_A_434_405#_c_622_n 0.0366796f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_40 VNB N_A_434_405#_c_623_n 0.0107381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_434_405#_c_624_n 0.0096311f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_42 VNB N_A_434_405#_c_625_n 0.0135759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_434_405#_c_626_n 0.00707257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_434_405#_c_627_n 0.00316125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_434_405#_c_628_n 0.00454424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_434_405#_c_629_n 0.00604027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_878_357#_c_714_n 0.0138253f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.625
cc_48 VNB N_A_878_357#_c_715_n 0.00964802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_878_357#_c_716_n 0.0120875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_878_357#_c_717_n 0.0184572f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.12
cc_51 VNB N_A_878_357#_c_718_n 0.0450995f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_52 VNB N_A_878_357#_c_719_n 0.00599831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_878_357#_c_720_n 0.0094758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_878_357#_c_721_n 0.0022791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_878_357#_c_722_n 0.0230025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_878_357#_c_723_n 0.00441542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1294_315#_c_823_n 0.00822433f $X=-0.19 $Y=-0.245 $X2=0.342
+ $Y2=1.625
cc_58 VNB N_A_1294_315#_M1020_g 0.0277565f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_59 VNB N_A_1294_315#_c_825_n 0.00892285f $X=-0.19 $Y=-0.245 $X2=0.29
+ $Y2=1.665
cc_60 VNB N_A_1294_315#_c_826_n 0.00986083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_GATE_c_923_n 0.00959432f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.172
cc_62 VNB N_GATE_c_924_n 0.0185919f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.408
cc_63 VNB N_GATE_M1007_g 0.00126817f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_64 VNB N_GATE_M1013_g 0.0267564f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.32
cc_65 VNB N_GATE_c_927_n 0.00629887f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_66 VNB GATE 0.0030793f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_67 VNB N_GATE_c_929_n 0.00177503f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_68 VNB N_SLEEP_B_M1004_g 0.0172181f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.955
cc_69 VNB N_SLEEP_B_M1003_g 0.00141661f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.625
cc_70 VNB N_SLEEP_B_M1032_g 0.0224602f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.625
cc_71 VNB N_SLEEP_B_c_970_n 0.0161954f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_72 VNB N_SLEEP_B_c_971_n 0.020369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_SLEEP_B_M1001_g 0.00169989f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_74 VNB N_SLEEP_B_c_973_n 0.017703f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=0.955
cc_75 VNB N_SLEEP_B_M1023_g 0.0313268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_SLEEP_B_M1015_g 0.0291058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_SLEEP_B_c_976_n 0.0167486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_SLEEP_B_c_977_n 0.0178603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_SLEEP_B_c_978_n 0.00197347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_SLEEP_B_c_979_n 0.00139549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_700_451#_M1022_g 0.0255465f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_82 VNB N_A_700_451#_c_1039_n 0.339519f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_83 VNB N_A_700_451#_c_1040_n 0.011606f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=0.955
cc_84 VNB N_A_700_451#_c_1041_n 0.0241775f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_85 VNB N_A_700_451#_M1006_g 0.0185744f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_86 VNB N_A_700_451#_M1017_g 0.0311548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_700_451#_M1027_g 0.015654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_700_451#_c_1045_n 0.0267619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_700_451#_c_1046_n 0.00570404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_700_451#_c_1047_n 0.0111713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_700_451#_c_1048_n 0.00669064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_700_451#_c_1049_n 0.00810429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_700_451#_c_1050_n 0.0027221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_700_451#_c_1051_n 0.00756103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_700_451#_c_1052_n 0.00417998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_700_451#_c_1053_n 0.0162536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2266_367#_M1008_g 0.0293615f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.32
cc_98 VNB N_A_2266_367#_M1018_g 6.66984e-19 $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_99 VNB N_A_2266_367#_c_1223_n 0.0395372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2266_367#_c_1224_n 0.0146779f $X=-0.19 $Y=-0.245 $X2=0.342
+ $Y2=1.12
cc_101 VNB N_A_2266_367#_c_1225_n 0.0113215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2266_367#_c_1226_n 0.0140875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2266_367#_c_1227_n 0.0092713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VPWR_c_1264_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_217_130#_c_1362_n 0.0082424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_217_130#_c_1363_n 0.0123945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_217_130#_c_1364_n 0.00357801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_217_130#_c_1365_n 0.00778396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_217_130#_c_1366_n 0.00604549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_217_130#_c_1367_n 0.00399925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_217_130#_c_1368_n 0.00221419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_217_130#_c_1369_n 0.00240624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_Q_c_1576_n 0.0573238f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_114 VNB N_VGND_c_1590_n 0.01004f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_115 VNB N_VGND_c_1591_n 0.0301542f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_116 VNB N_VGND_c_1592_n 0.0142647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1593_n 0.0157676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1594_n 0.00519587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1595_n 0.00594195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1596_n 0.0431681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1597_n 0.0229267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1598_n 0.0186317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1599_n 0.0288733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1600_n 0.00360663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1601_n 0.036295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1602_n 0.0933335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1603_n 0.0187707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1604_n 0.0772482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1605_n 0.0221298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1606_n 0.0193242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1607_n 0.646871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1608_n 0.00286121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1609_n 0.00448506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1610_n 0.00536178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1611_n 0.00476075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1612_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_988_47#_c_1744_n 0.00625957f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=1.625
cc_138 VNB N_A_988_47#_c_1745_n 0.0214021f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.32
cc_139 VNB N_A_988_47#_c_1746_n 0.00506232f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_140 VNB N_A_988_47#_c_1747_n 0.00676255f $X=-0.19 $Y=-0.245 $X2=0.342
+ $Y2=1.12
cc_141 VNB N_A_988_47#_c_1748_n 0.01289f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_142 VPB N_D_M1028_g 0.039884f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.32
cc_143 VPB N_D_c_236_n 0.00747698f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_144 VPB N_A_27_400#_M1005_g 0.0269281f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.32
cc_145 VPB N_A_27_400#_c_272_n 0.00445022f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=0.955
cc_146 VPB N_A_27_400#_c_273_n 0.00333657f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.665
cc_147 VPB N_A_27_400#_c_274_n 0.033052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_27_400#_c_269_n 0.00289005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_27_400#_c_270_n 0.01775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_SET_B_M1026_g 0.0400227f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.32
cc_151 VPB N_A_404_353#_c_431_n 0.0237344f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.625
cc_152 VPB N_A_404_353#_M1034_g 0.00792129f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_153 VPB N_A_404_353#_c_433_n 0.0408374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_404_353#_c_434_n 0.0211035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_404_353#_M1033_g 0.0211799f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_156 VPB N_A_404_353#_M1030_g 0.018599f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.295
cc_157 VPB N_A_404_353#_c_437_n 0.00114233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_404_353#_c_422_n 0.00435369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_404_353#_c_439_n 0.0290789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_404_353#_c_423_n 0.0184468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_404_353#_c_426_n 0.00464402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_404_353#_c_442_n 0.00232021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_404_353#_c_443_n 0.0401422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_434_405#_M1014_g 0.0328635f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_165 VPB N_A_434_405#_c_625_n 0.0391338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_434_405#_c_626_n 2.64875e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_434_405#_c_633_n 0.00681664f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_878_357#_M1000_g 0.0282613f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.32
cc_169 VPB N_A_878_357#_c_725_n 0.00170719f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.665
cc_170 VPB N_A_878_357#_c_720_n 0.0517759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_878_357#_c_727_n 0.0158919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_878_357#_c_728_n 4.8461e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_878_357#_c_729_n 0.00566097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_878_357#_c_723_n 0.00512039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_1294_315#_M1002_g 0.0333126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_1294_315#_c_823_n 0.0250161f $X=-0.19 $Y=1.655 $X2=0.342
+ $Y2=1.625
cc_177 VPB N_A_1294_315#_c_829_n 0.094635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_1294_315#_c_830_n 0.0177998f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.12
cc_179 VPB N_A_1294_315#_c_831_n 0.00999542f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_180 VPB N_A_1294_315#_c_832_n 0.0146245f $X=-0.19 $Y=1.655 $X2=0.342
+ $Y2=0.955
cc_181 VPB N_A_1294_315#_c_833_n 0.00458704f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_182 VPB N_A_1294_315#_c_825_n 0.00121211f $X=-0.19 $Y=1.655 $X2=0.29
+ $Y2=1.665
cc_183 VPB N_A_1294_315#_c_835_n 0.00178556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1294_315#_c_836_n 0.0577431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1294_315#_c_837_n 0.00988732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_GATE_M1007_g 0.0570952f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.555
cc_187 VPB GATE 0.00271744f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_188 VPB N_GATE_c_929_n 0.0453658f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_189 VPB N_SLEEP_B_M1003_g 0.0229178f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.625
cc_190 VPB N_SLEEP_B_M1001_g 0.0323252f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_191 VPB N_SLEEP_B_c_978_n 0.0502359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_SLEEP_B_c_979_n 0.0105144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_700_451#_M1009_g 0.0262446f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.12
cc_194 VPB N_A_700_451#_M1027_g 0.0289385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_700_451#_c_1056_n 0.00300409f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_700_451#_c_1046_n 0.00665744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_700_451#_c_1058_n 0.00839184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_700_451#_c_1059_n 0.0157738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_700_451#_c_1051_n 0.0033687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_700_451#_c_1061_n 0.00815924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_700_451#_c_1052_n 0.00208702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_700_451#_c_1053_n 0.0120871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_2266_367#_M1018_g 0.0292315f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_204 VPB N_A_2266_367#_c_1229_n 0.0218142f $X=-0.19 $Y=1.655 $X2=0.342
+ $Y2=0.955
cc_205 VPB N_VPWR_c_1265_n 0.0169309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1266_n 0.0178582f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.12
cc_207 VPB N_VPWR_c_1267_n 0.0147273f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_208 VPB N_VPWR_c_1268_n 0.0212444f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.665
cc_209 VPB N_VPWR_c_1269_n 0.280265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1270_n 0.0188222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1264_n 0.0877663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1272_n 0.027469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1273_n 0.00631563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1274_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_217_130#_c_1370_n 0.00432829f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_216 VPB N_A_217_130#_c_1371_n 0.0062322f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_217 VPB N_A_217_130#_c_1372_n 0.0200129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_217_130#_c_1373_n 0.00557272f $X=-0.19 $Y=1.655 $X2=0.29
+ $Y2=1.665
cc_219 VPB N_A_217_130#_c_1368_n 0.00749009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_217_130#_c_1375_n 0.00375049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_217_130#_c_1369_n 0.0100067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_217_130#_c_1377_n 0.00894665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_KAPWR_c_1479_n 0.0168757f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=0.955
cc_224 VPB N_KAPWR_c_1480_n 0.0103531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_KAPWR_c_1481_n 0.00233841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_KAPWR_c_1482_n 0.120327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_KAPWR_c_1483_n 0.0175351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_Q_c_1576_n 0.0481696f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_229 N_D_M1028_g N_A_27_400#_M1005_g 0.0195673f $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_230 N_D_M1028_g N_A_27_400#_c_272_n 0.0117269f $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_231 N_D_c_236_n N_A_27_400#_c_272_n 0.00123997f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_232 N_D_M1024_g N_A_27_400#_c_267_n 0.00600966f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_233 N_D_c_235_n N_A_27_400#_c_267_n 0.0134909f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_234 N_D_c_236_n N_A_27_400#_c_267_n 0.0313985f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_235 N_D_M1028_g N_A_27_400#_c_273_n 0.00389575f $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_236 N_D_M1028_g N_A_27_400#_c_274_n 0.00903301f $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_237 N_D_c_234_n N_A_27_400#_c_274_n 0.00153536f $X=0.342 $Y=1.625 $X2=0 $Y2=0
cc_238 N_D_c_236_n N_A_27_400#_c_274_n 0.0255629f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_239 N_D_M1024_g N_A_27_400#_c_268_n 0.0078524f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_240 N_D_c_235_n N_A_27_400#_c_268_n 4.6035e-19 $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_241 N_D_c_234_n N_A_27_400#_c_269_n 0.00300675f $X=0.342 $Y=1.625 $X2=0 $Y2=0
cc_242 N_D_c_236_n N_A_27_400#_c_269_n 0.0193848f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_243 N_D_c_234_n N_A_27_400#_c_270_n 0.0169427f $X=0.342 $Y=1.625 $X2=0 $Y2=0
cc_244 N_D_c_236_n N_A_27_400#_c_270_n 2.66794e-19 $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_245 N_D_M1028_g N_VPWR_c_1265_n 0.00551379f $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_246 N_D_M1028_g N_VPWR_c_1264_n 7.18873e-19 $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_247 N_D_M1028_g N_VPWR_c_1272_n 0.00249171f $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_248 N_D_M1024_g N_A_217_130#_c_1362_n 3.37537e-19 $X=0.475 $Y=0.555 $X2=0
+ $Y2=0
cc_249 N_D_M1028_g N_KAPWR_c_1482_n 0.00620723f $X=0.485 $Y=2.32 $X2=0 $Y2=0
cc_250 N_D_M1024_g N_VGND_c_1591_n 0.00573369f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_251 N_D_c_235_n N_VGND_c_1591_n 0.0017067f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_252 N_D_c_236_n N_VGND_c_1591_n 0.0194357f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_253 N_D_M1024_g N_VGND_c_1601_n 0.00453398f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_254 N_D_M1024_g N_VGND_c_1607_n 0.00911701f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_255 N_A_27_400#_M1031_g N_SET_B_c_336_n 0.0514554f $X=1.425 $Y=0.97 $X2=0
+ $Y2=0
cc_256 N_A_27_400#_c_265_n N_A_434_405#_c_626_n 0.00278534f $X=1.35 $Y=1.555
+ $X2=0 $Y2=0
cc_257 N_A_27_400#_c_272_n N_VPWR_M1028_d 0.00519094f $X=0.685 $Y=2.065
+ $X2=-0.19 $Y2=-0.245
cc_258 N_A_27_400#_M1005_g N_VPWR_c_1265_n 0.0128319f $X=1.02 $Y=2.42 $X2=0
+ $Y2=0
cc_259 N_A_27_400#_c_272_n N_VPWR_c_1265_n 0.0175964f $X=0.685 $Y=2.065 $X2=0
+ $Y2=0
cc_260 N_A_27_400#_c_274_n N_VPWR_c_1265_n 0.022883f $X=0.27 $Y=2.145 $X2=0
+ $Y2=0
cc_261 N_A_27_400#_c_269_n N_VPWR_c_1265_n 0.00284724f $X=0.965 $Y=1.645 $X2=0
+ $Y2=0
cc_262 N_A_27_400#_c_270_n N_VPWR_c_1265_n 0.00164629f $X=0.965 $Y=1.555 $X2=0
+ $Y2=0
cc_263 N_A_27_400#_M1005_g N_VPWR_c_1266_n 0.00410575f $X=1.02 $Y=2.42 $X2=0
+ $Y2=0
cc_264 N_A_27_400#_M1005_g N_VPWR_c_1267_n 0.00125756f $X=1.02 $Y=2.42 $X2=0
+ $Y2=0
cc_265 N_A_27_400#_M1005_g N_VPWR_c_1264_n 0.00248276f $X=1.02 $Y=2.42 $X2=0
+ $Y2=0
cc_266 N_A_27_400#_c_274_n N_VPWR_c_1272_n 0.00518715f $X=0.27 $Y=2.145 $X2=0
+ $Y2=0
cc_267 N_A_27_400#_M1031_g N_A_217_130#_c_1362_n 0.0111083f $X=1.425 $Y=0.97
+ $X2=0 $Y2=0
cc_268 N_A_27_400#_c_268_n N_A_217_130#_c_1362_n 0.0256865f $X=0.69 $Y=0.555
+ $X2=0 $Y2=0
cc_269 N_A_27_400#_M1005_g N_A_217_130#_c_1370_n 0.00354757f $X=1.02 $Y=2.42
+ $X2=0 $Y2=0
cc_270 N_A_27_400#_c_265_n N_A_217_130#_c_1370_n 0.00315691f $X=1.35 $Y=1.555
+ $X2=0 $Y2=0
cc_271 N_A_27_400#_c_272_n N_A_217_130#_c_1370_n 0.00564875f $X=0.685 $Y=2.065
+ $X2=0 $Y2=0
cc_272 N_A_27_400#_M1005_g N_A_217_130#_c_1373_n 5.96075e-19 $X=1.02 $Y=2.42
+ $X2=0 $Y2=0
cc_273 N_A_27_400#_M1031_g N_A_217_130#_c_1367_n 0.00472019f $X=1.425 $Y=0.97
+ $X2=0 $Y2=0
cc_274 N_A_27_400#_c_267_n N_A_217_130#_c_1367_n 0.0256865f $X=0.77 $Y=1.48
+ $X2=0 $Y2=0
cc_275 N_A_27_400#_c_269_n N_A_217_130#_c_1367_n 0.007084f $X=0.965 $Y=1.645
+ $X2=0 $Y2=0
cc_276 N_A_27_400#_c_270_n N_A_217_130#_c_1367_n 0.00696536f $X=0.965 $Y=1.555
+ $X2=0 $Y2=0
cc_277 N_A_27_400#_M1005_g N_A_217_130#_c_1368_n 0.00251379f $X=1.02 $Y=2.42
+ $X2=0 $Y2=0
cc_278 N_A_27_400#_c_265_n N_A_217_130#_c_1368_n 0.0123637f $X=1.35 $Y=1.555
+ $X2=0 $Y2=0
cc_279 N_A_27_400#_M1031_g N_A_217_130#_c_1368_n 0.00849234f $X=1.425 $Y=0.97
+ $X2=0 $Y2=0
cc_280 N_A_27_400#_c_267_n N_A_217_130#_c_1368_n 0.00464631f $X=0.77 $Y=1.48
+ $X2=0 $Y2=0
cc_281 N_A_27_400#_c_273_n N_A_217_130#_c_1368_n 0.00462017f $X=0.77 $Y=1.98
+ $X2=0 $Y2=0
cc_282 N_A_27_400#_c_269_n N_A_217_130#_c_1368_n 0.0247917f $X=0.965 $Y=1.645
+ $X2=0 $Y2=0
cc_283 N_A_27_400#_c_270_n N_A_217_130#_c_1368_n 0.00126186f $X=0.965 $Y=1.555
+ $X2=0 $Y2=0
cc_284 N_A_27_400#_M1005_g N_KAPWR_c_1482_n 0.00747531f $X=1.02 $Y=2.42 $X2=0
+ $Y2=0
cc_285 N_A_27_400#_c_272_n N_KAPWR_c_1482_n 0.00703889f $X=0.685 $Y=2.065 $X2=0
+ $Y2=0
cc_286 N_A_27_400#_c_274_n N_KAPWR_c_1482_n 0.014528f $X=0.27 $Y=2.145 $X2=0
+ $Y2=0
cc_287 N_A_27_400#_c_268_n N_VGND_c_1591_n 0.0179429f $X=0.69 $Y=0.555 $X2=0
+ $Y2=0
cc_288 N_A_27_400#_M1031_g N_VGND_c_1592_n 0.00234669f $X=1.425 $Y=0.97 $X2=0
+ $Y2=0
cc_289 N_A_27_400#_M1031_g N_VGND_c_1593_n 0.00223752f $X=1.425 $Y=0.97 $X2=0
+ $Y2=0
cc_290 N_A_27_400#_M1031_g N_VGND_c_1601_n 0.00330012f $X=1.425 $Y=0.97 $X2=0
+ $Y2=0
cc_291 N_A_27_400#_c_268_n N_VGND_c_1601_n 0.0159714f $X=0.69 $Y=0.555 $X2=0
+ $Y2=0
cc_292 N_A_27_400#_M1031_g N_VGND_c_1607_n 0.00462577f $X=1.425 $Y=0.97 $X2=0
+ $Y2=0
cc_293 N_A_27_400#_c_268_n N_VGND_c_1607_n 0.0121063f $X=0.69 $Y=0.555 $X2=0
+ $Y2=0
cc_294 N_SET_B_c_332_n N_A_404_353#_M1034_g 0.0129305f $X=1.785 $Y=0.53 $X2=0
+ $Y2=0
cc_295 N_SET_B_c_338_n N_A_404_353#_M1034_g 0.00220915f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_296 N_SET_B_c_339_n N_A_404_353#_M1034_g 0.00540924f $X=2.145 $Y=0.365 $X2=0
+ $Y2=0
cc_297 N_SET_B_c_340_n N_A_404_353#_M1034_g 5.09464e-19 $X=2.31 $Y=0.365 $X2=0
+ $Y2=0
cc_298 N_SET_B_c_338_n N_A_404_353#_M1029_g 0.00968138f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_299 N_SET_B_M1026_g N_A_404_353#_c_439_n 0.0168514f $X=6.105 $Y=2.205 $X2=0
+ $Y2=0
cc_300 N_SET_B_c_338_n N_A_434_405#_c_618_n 0.0112969f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_301 N_SET_B_c_338_n N_A_434_405#_M1021_g 0.0135252f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_302 N_SET_B_c_338_n N_A_434_405#_c_622_n 0.00109887f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_303 N_SET_B_c_338_n N_A_434_405#_c_627_n 0.00626639f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_304 N_SET_B_c_332_n N_A_434_405#_c_628_n 5.71421e-19 $X=1.785 $Y=0.53 $X2=0
+ $Y2=0
cc_305 N_SET_B_c_338_n N_A_434_405#_c_629_n 0.012328f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_306 N_SET_B_c_338_n N_A_878_357#_c_714_n 0.00874071f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_307 N_SET_B_c_338_n N_A_878_357#_c_717_n 0.014766f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_308 SET_B N_A_878_357#_c_717_n 0.00169058f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_309 N_SET_B_c_342_n N_A_878_357#_c_717_n 0.00671248f $X=5.6 $Y=0.305 $X2=0
+ $Y2=0
cc_310 N_SET_B_M1026_g N_A_878_357#_c_727_n 0.0182651f $X=6.105 $Y=2.205 $X2=0
+ $Y2=0
cc_311 N_SET_B_M1026_g N_A_1294_315#_c_823_n 0.0845585f $X=6.105 $Y=2.205 $X2=0
+ $Y2=0
cc_312 N_SET_B_M1026_g N_A_1294_315#_M1020_g 9.66366e-19 $X=6.105 $Y=2.205 $X2=0
+ $Y2=0
cc_313 N_SET_B_M1011_g N_A_1294_315#_M1020_g 0.0152835f $X=6.235 $Y=0.845 $X2=0
+ $Y2=0
cc_314 N_SET_B_c_338_n N_A_700_451#_M1021_d 0.00536937f $X=5.435 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_315 N_SET_B_c_338_n N_A_700_451#_c_1065_n 0.00844204f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_316 N_SET_B_c_338_n N_A_700_451#_c_1047_n 0.0463891f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_317 N_SET_B_M1026_g N_A_700_451#_c_1059_n 0.0172798f $X=6.105 $Y=2.205 $X2=0
+ $Y2=0
cc_318 N_SET_B_c_337_n N_A_700_451#_c_1059_n 0.0021836f $X=6.145 $Y=1.315 $X2=0
+ $Y2=0
cc_319 N_SET_B_c_337_n N_A_700_451#_c_1051_n 0.00371242f $X=6.145 $Y=1.315 $X2=0
+ $Y2=0
cc_320 N_SET_B_M1026_g N_A_700_451#_c_1061_n 0.00890344f $X=6.105 $Y=2.205 $X2=0
+ $Y2=0
cc_321 N_SET_B_M1026_g N_VPWR_c_1269_n 0.00490748f $X=6.105 $Y=2.205 $X2=0 $Y2=0
cc_322 N_SET_B_M1026_g N_VPWR_c_1264_n 0.00129538f $X=6.105 $Y=2.205 $X2=0 $Y2=0
cc_323 N_SET_B_c_338_n N_A_217_130#_M1019_s 0.00474891f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_324 N_SET_B_c_332_n N_A_217_130#_c_1362_n 0.00244235f $X=1.785 $Y=0.53 $X2=0
+ $Y2=0
cc_325 N_SET_B_c_338_n N_A_217_130#_c_1365_n 0.0343911f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_326 N_SET_B_M1026_g N_KAPWR_c_1482_n 0.0102003f $X=6.105 $Y=2.205 $X2=0 $Y2=0
cc_327 N_SET_B_c_332_n N_VGND_c_1592_n 0.00599851f $X=1.785 $Y=0.53 $X2=0 $Y2=0
cc_328 N_SET_B_c_336_n N_VGND_c_1592_n 0.0168451f $X=1.86 $Y=0.365 $X2=0 $Y2=0
cc_329 N_SET_B_c_340_n N_VGND_c_1592_n 0.0163912f $X=2.31 $Y=0.365 $X2=0 $Y2=0
cc_330 N_SET_B_c_332_n N_VGND_c_1593_n 0.022124f $X=1.785 $Y=0.53 $X2=0 $Y2=0
cc_331 N_SET_B_c_339_n N_VGND_c_1593_n 0.00780505f $X=2.145 $Y=0.365 $X2=0 $Y2=0
cc_332 N_SET_B_c_340_n N_VGND_c_1593_n 0.0127862f $X=2.31 $Y=0.365 $X2=0 $Y2=0
cc_333 N_SET_B_c_333_n N_VGND_c_1594_n 0.0189858f $X=6.16 $Y=0.305 $X2=0 $Y2=0
cc_334 N_SET_B_M1011_g N_VGND_c_1594_n 0.0123122f $X=6.235 $Y=0.845 $X2=0 $Y2=0
cc_335 N_SET_B_c_337_n N_VGND_c_1594_n 0.00107698f $X=6.145 $Y=1.315 $X2=0 $Y2=0
cc_336 SET_B N_VGND_c_1594_n 0.0297716f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_337 N_SET_B_c_342_n N_VGND_c_1594_n 6.63207e-19 $X=5.6 $Y=0.305 $X2=0 $Y2=0
cc_338 N_SET_B_c_333_n N_VGND_c_1595_n 0.00507788f $X=6.16 $Y=0.305 $X2=0 $Y2=0
cc_339 N_SET_B_M1011_g N_VGND_c_1595_n 4.33145e-19 $X=6.235 $Y=0.845 $X2=0 $Y2=0
cc_340 N_SET_B_c_336_n N_VGND_c_1602_n 0.00984171f $X=1.86 $Y=0.365 $X2=0 $Y2=0
cc_341 N_SET_B_c_340_n N_VGND_c_1602_n 0.201979f $X=2.31 $Y=0.365 $X2=0 $Y2=0
cc_342 SET_B N_VGND_c_1602_n 0.0215354f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_343 N_SET_B_c_342_n N_VGND_c_1602_n 0.0105048f $X=5.6 $Y=0.305 $X2=0 $Y2=0
cc_344 N_SET_B_c_333_n N_VGND_c_1603_n 0.00389963f $X=6.16 $Y=0.305 $X2=0 $Y2=0
cc_345 N_SET_B_c_333_n N_VGND_c_1607_n 0.0169083f $X=6.16 $Y=0.305 $X2=0 $Y2=0
cc_346 N_SET_B_c_336_n N_VGND_c_1607_n 0.00135675f $X=1.86 $Y=0.365 $X2=0 $Y2=0
cc_347 N_SET_B_c_339_n N_VGND_c_1607_n 0.0116523f $X=2.145 $Y=0.365 $X2=0 $Y2=0
cc_348 N_SET_B_c_340_n N_VGND_c_1607_n 0.125045f $X=2.31 $Y=0.365 $X2=0 $Y2=0
cc_349 SET_B N_VGND_c_1607_n 0.0111266f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_350 N_SET_B_c_342_n N_VGND_c_1607_n 0.00753695f $X=5.6 $Y=0.305 $X2=0 $Y2=0
cc_351 N_SET_B_c_338_n A_667_47# 0.00192199f $X=5.435 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_352 N_SET_B_c_338_n A_844_47# 0.00192448f $X=5.435 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_353 N_SET_B_c_338_n A_916_47# 0.00187064f $X=5.435 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_354 N_SET_B_c_338_n N_A_988_47#_M1016_d 0.00867816f $X=5.435 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_355 N_SET_B_c_338_n N_A_988_47#_c_1744_n 0.00573384f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_356 SET_B N_A_988_47#_c_1744_n 0.00356706f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_357 N_SET_B_c_342_n N_A_988_47#_c_1744_n 2.39436e-19 $X=5.6 $Y=0.305 $X2=0
+ $Y2=0
cc_358 N_SET_B_M1011_g N_A_988_47#_c_1745_n 0.00829166f $X=6.235 $Y=0.845 $X2=0
+ $Y2=0
cc_359 N_SET_B_c_337_n N_A_988_47#_c_1745_n 0.0142866f $X=6.145 $Y=1.315 $X2=0
+ $Y2=0
cc_360 SET_B N_A_988_47#_c_1745_n 0.00352372f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_361 N_SET_B_c_342_n N_A_988_47#_c_1745_n 6.01923e-19 $X=5.6 $Y=0.305 $X2=0
+ $Y2=0
cc_362 N_SET_B_M1011_g N_A_988_47#_c_1746_n 0.00729227f $X=6.235 $Y=0.845 $X2=0
+ $Y2=0
cc_363 N_SET_B_c_338_n N_A_988_47#_c_1747_n 0.0181818f $X=5.435 $Y=0.34 $X2=0
+ $Y2=0
cc_364 SET_B N_A_988_47#_c_1747_n 0.00580928f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_365 N_SET_B_M1011_g N_A_988_47#_c_1748_n 0.00385524f $X=6.235 $Y=0.845 $X2=0
+ $Y2=0
cc_366 N_SET_B_c_337_n N_A_988_47#_c_1748_n 3.78473e-19 $X=6.145 $Y=1.315 $X2=0
+ $Y2=0
cc_367 SET_B N_A_988_47#_c_1748_n 0.0138555f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_368 N_SET_B_c_342_n N_A_988_47#_c_1748_n 9.85675e-19 $X=5.6 $Y=0.305 $X2=0
+ $Y2=0
cc_369 N_A_404_353#_c_443_n N_A_434_405#_c_619_n 0.00197719f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_370 N_A_404_353#_M1029_g N_A_434_405#_M1021_g 0.0279185f $X=4.145 $Y=0.445
+ $X2=0 $Y2=0
cc_371 N_A_404_353#_c_422_n N_A_434_405#_c_621_n 4.45224e-19 $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_372 N_A_404_353#_c_437_n N_A_434_405#_M1014_g 0.0010355f $X=3.27 $Y=2.905
+ $X2=0 $Y2=0
cc_373 N_A_404_353#_c_454_p N_A_434_405#_M1014_g 0.0161212f $X=4.23 $Y=2.99
+ $X2=0 $Y2=0
cc_374 N_A_404_353#_c_455_p N_A_434_405#_M1014_g 0.00524681f $X=4.315 $Y=2.905
+ $X2=0 $Y2=0
cc_375 N_A_404_353#_c_442_n N_A_434_405#_M1014_g 3.1694e-19 $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_376 N_A_404_353#_c_443_n N_A_434_405#_M1014_g 0.0312366f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_377 N_A_404_353#_c_458_p N_A_434_405#_M1014_g 0.00173488f $X=4.315 $Y=2.4
+ $X2=0 $Y2=0
cc_378 N_A_404_353#_M1034_g N_A_434_405#_c_622_n 0.00479524f $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_379 N_A_404_353#_c_433_n N_A_434_405#_c_622_n 0.00563452f $X=2.99 $Y=1.84
+ $X2=0 $Y2=0
cc_380 N_A_404_353#_c_443_n N_A_434_405#_c_623_n 0.00563452f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_381 N_A_404_353#_c_427_n N_A_434_405#_c_624_n 3.20598e-19 $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_382 N_A_404_353#_c_428_n N_A_434_405#_c_624_n 0.0103156f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_383 N_A_404_353#_c_422_n N_A_434_405#_c_625_n 0.00881654f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_384 N_A_404_353#_c_443_n N_A_434_405#_c_625_n 0.00273748f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_385 N_A_404_353#_c_427_n N_A_434_405#_c_625_n 5.99496e-19 $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_386 N_A_404_353#_c_428_n N_A_434_405#_c_625_n 0.00456405f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_387 N_A_404_353#_M1034_g N_A_434_405#_c_626_n 0.0144081f $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_388 N_A_404_353#_c_431_n N_A_434_405#_c_633_n 0.0119847f $X=2.095 $Y=1.915
+ $X2=0 $Y2=0
cc_389 N_A_404_353#_M1034_g N_A_434_405#_c_633_n 0.00460726f $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_390 N_A_404_353#_c_433_n N_A_434_405#_c_633_n 0.00960617f $X=2.99 $Y=1.84
+ $X2=0 $Y2=0
cc_391 N_A_404_353#_c_434_n N_A_434_405#_c_633_n 0.0109027f $X=2.385 $Y=1.84
+ $X2=0 $Y2=0
cc_392 N_A_404_353#_M1034_g N_A_434_405#_c_628_n 0.00886958f $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_393 N_A_404_353#_M1034_g N_A_434_405#_c_629_n 0.00586998f $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_394 N_A_404_353#_c_433_n N_A_434_405#_c_629_n 0.00538021f $X=2.99 $Y=1.84
+ $X2=0 $Y2=0
cc_395 N_A_404_353#_c_439_n N_A_878_357#_M1009_d 0.00471378f $X=7.92 $Y=2.4
+ $X2=0 $Y2=0
cc_396 N_A_404_353#_c_454_p N_A_878_357#_M1000_g 0.00447047f $X=4.23 $Y=2.99
+ $X2=0 $Y2=0
cc_397 N_A_404_353#_c_422_n N_A_878_357#_M1000_g 0.0127933f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_398 N_A_404_353#_c_455_p N_A_878_357#_M1000_g 0.0123132f $X=4.315 $Y=2.905
+ $X2=0 $Y2=0
cc_399 N_A_404_353#_c_439_n N_A_878_357#_M1000_g 0.0216577f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_400 N_A_404_353#_c_458_p N_A_878_357#_M1000_g 0.00129677f $X=4.315 $Y=2.4
+ $X2=0 $Y2=0
cc_401 N_A_404_353#_M1029_g N_A_878_357#_c_714_n 0.0531511f $X=4.145 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_404_353#_M1029_g N_A_878_357#_c_718_n 0.00264107f $X=4.145 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_404_353#_c_422_n N_A_878_357#_c_718_n 0.00404047f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_404 N_A_404_353#_c_427_n N_A_878_357#_c_718_n 2.066e-19 $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_405 N_A_404_353#_c_428_n N_A_878_357#_c_718_n 0.00827835f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_406 N_A_404_353#_c_422_n N_A_878_357#_c_725_n 0.0197009f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_407 N_A_404_353#_c_422_n N_A_878_357#_c_720_n 0.00665743f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_408 N_A_404_353#_c_439_n N_A_878_357#_c_720_n 0.00132626f $X=7.92 $Y=2.4
+ $X2=0 $Y2=0
cc_409 N_A_404_353#_c_428_n N_A_878_357#_c_720_n 3.83538e-19 $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_410 N_A_404_353#_c_439_n N_A_878_357#_c_727_n 0.150397f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_411 N_A_404_353#_c_422_n N_A_878_357#_c_728_n 0.00981726f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_412 N_A_404_353#_c_439_n N_A_878_357#_c_728_n 0.021142f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_413 N_A_404_353#_c_424_n N_A_878_357#_c_721_n 0.014132f $X=8.09 $Y=1.225
+ $X2=0 $Y2=0
cc_414 N_A_404_353#_c_429_n N_A_878_357#_c_721_n 0.00850192f $X=8.425 $Y=1.08
+ $X2=0 $Y2=0
cc_415 N_A_404_353#_c_430_n N_A_878_357#_c_721_n 0.00868033f $X=8.755 $Y=1.08
+ $X2=0 $Y2=0
cc_416 N_A_404_353#_c_439_n N_A_878_357#_c_729_n 0.0209832f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_417 N_A_404_353#_c_423_n N_A_878_357#_c_723_n 0.0645385f $X=8.005 $Y=2.315
+ $X2=0 $Y2=0
cc_418 N_A_404_353#_c_424_n N_A_878_357#_c_723_n 0.0136815f $X=8.09 $Y=1.225
+ $X2=0 $Y2=0
cc_419 N_A_404_353#_c_430_n N_A_878_357#_c_723_n 0.00452322f $X=8.755 $Y=1.08
+ $X2=0 $Y2=0
cc_420 N_A_404_353#_c_439_n N_A_1294_315#_M1002_g 0.0159706f $X=7.92 $Y=2.4
+ $X2=0 $Y2=0
cc_421 N_A_404_353#_c_439_n N_A_1294_315#_c_829_n 0.0126852f $X=7.92 $Y=2.4
+ $X2=0 $Y2=0
cc_422 N_A_404_353#_M1007_d N_A_1294_315#_c_832_n 0.00522917f $X=8.975 $Y=2.33
+ $X2=0 $Y2=0
cc_423 N_A_404_353#_c_426_n N_A_1294_315#_c_832_n 0.0211691f $X=9.23 $Y=1.985
+ $X2=0 $Y2=0
cc_424 N_A_404_353#_c_439_n N_A_1294_315#_c_833_n 0.0154601f $X=7.92 $Y=2.4
+ $X2=0 $Y2=0
cc_425 N_A_404_353#_c_439_n N_A_1294_315#_c_836_n 6.78261e-19 $X=7.92 $Y=2.4
+ $X2=0 $Y2=0
cc_426 N_A_404_353#_c_439_n N_A_1294_315#_c_837_n 0.00172338f $X=7.92 $Y=2.4
+ $X2=0 $Y2=0
cc_427 N_A_404_353#_c_425_n N_GATE_c_923_n 0.00486237f $X=9.065 $Y=1.225
+ $X2=-0.19 $Y2=-0.245
cc_428 N_A_404_353#_c_423_n N_GATE_c_924_n 0.0153174f $X=8.005 $Y=2.315 $X2=0
+ $Y2=0
cc_429 N_A_404_353#_c_429_n N_GATE_c_924_n 0.002388f $X=8.425 $Y=1.08 $X2=0
+ $Y2=0
cc_430 N_A_404_353#_c_430_n N_GATE_c_924_n 0.00486237f $X=8.755 $Y=1.08 $X2=0
+ $Y2=0
cc_431 N_A_404_353#_c_426_n N_GATE_M1007_g 0.00640341f $X=9.23 $Y=1.985 $X2=0
+ $Y2=0
cc_432 N_A_404_353#_c_425_n N_GATE_M1013_g 0.0208503f $X=9.065 $Y=1.225 $X2=0
+ $Y2=0
cc_433 N_A_404_353#_c_426_n N_GATE_M1013_g 0.0062214f $X=9.23 $Y=1.985 $X2=0
+ $Y2=0
cc_434 N_A_404_353#_c_430_n N_GATE_M1013_g 0.0117812f $X=8.755 $Y=1.08 $X2=0
+ $Y2=0
cc_435 N_A_404_353#_c_423_n GATE 0.0453865f $X=8.005 $Y=2.315 $X2=0 $Y2=0
cc_436 N_A_404_353#_c_426_n GATE 0.0255318f $X=9.23 $Y=1.985 $X2=0 $Y2=0
cc_437 N_A_404_353#_c_429_n GATE 0.027306f $X=8.425 $Y=1.08 $X2=0 $Y2=0
cc_438 N_A_404_353#_c_425_n N_SLEEP_B_M1004_g 0.0115991f $X=9.065 $Y=1.225 $X2=0
+ $Y2=0
cc_439 N_A_404_353#_c_426_n N_SLEEP_B_M1004_g 0.0037772f $X=9.23 $Y=1.985 $X2=0
+ $Y2=0
cc_440 N_A_404_353#_c_426_n N_SLEEP_B_M1003_g 0.0143005f $X=9.23 $Y=1.985 $X2=0
+ $Y2=0
cc_441 N_A_404_353#_c_425_n N_SLEEP_B_M1032_g 5.14957e-19 $X=9.065 $Y=1.225
+ $X2=0 $Y2=0
cc_442 N_A_404_353#_c_426_n N_SLEEP_B_M1032_g 0.00373667f $X=9.23 $Y=1.985 $X2=0
+ $Y2=0
cc_443 N_A_404_353#_c_426_n N_SLEEP_B_c_971_n 0.0136735f $X=9.23 $Y=1.985 $X2=0
+ $Y2=0
cc_444 N_A_404_353#_c_426_n N_SLEEP_B_M1001_g 0.00241493f $X=9.23 $Y=1.985 $X2=0
+ $Y2=0
cc_445 N_A_404_353#_c_454_p N_A_700_451#_M1030_d 0.00482454f $X=4.23 $Y=2.99
+ $X2=0 $Y2=0
cc_446 N_A_404_353#_c_439_n N_A_700_451#_M1026_s 0.0102355f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_447 N_A_404_353#_c_439_n N_A_700_451#_M1009_g 0.0158763f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_448 N_A_404_353#_c_423_n N_A_700_451#_M1009_g 0.0052097f $X=8.005 $Y=2.315
+ $X2=0 $Y2=0
cc_449 N_A_404_353#_c_430_n N_A_700_451#_c_1039_n 0.00846154f $X=8.755 $Y=1.08
+ $X2=0 $Y2=0
cc_450 N_A_404_353#_c_423_n N_A_700_451#_c_1041_n 6.79993e-19 $X=8.005 $Y=2.315
+ $X2=0 $Y2=0
cc_451 N_A_404_353#_c_424_n N_A_700_451#_M1006_g 0.00444975f $X=8.09 $Y=1.225
+ $X2=0 $Y2=0
cc_452 N_A_404_353#_c_430_n N_A_700_451#_M1006_g 0.00282113f $X=8.755 $Y=1.08
+ $X2=0 $Y2=0
cc_453 N_A_404_353#_c_422_n N_A_700_451#_c_1056_n 0.0111509f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_454 N_A_404_353#_c_442_n N_A_700_451#_c_1056_n 0.0188902f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_455 N_A_404_353#_c_443_n N_A_700_451#_c_1056_n 0.00304962f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_456 N_A_404_353#_M1030_g N_A_700_451#_c_1082_n 0.00304962f $X=3.425 $Y=2.675
+ $X2=0 $Y2=0
cc_457 N_A_404_353#_c_437_n N_A_700_451#_c_1082_n 0.0188902f $X=3.27 $Y=2.905
+ $X2=0 $Y2=0
cc_458 N_A_404_353#_c_454_p N_A_700_451#_c_1082_n 0.0210043f $X=4.23 $Y=2.99
+ $X2=0 $Y2=0
cc_459 N_A_404_353#_c_455_p N_A_700_451#_c_1082_n 0.010894f $X=4.315 $Y=2.905
+ $X2=0 $Y2=0
cc_460 N_A_404_353#_c_458_p N_A_700_451#_c_1082_n 0.00884729f $X=4.315 $Y=2.4
+ $X2=0 $Y2=0
cc_461 N_A_404_353#_M1029_g N_A_700_451#_c_1046_n 0.00681827f $X=4.145 $Y=0.445
+ $X2=0 $Y2=0
cc_462 N_A_404_353#_c_422_n N_A_700_451#_c_1046_n 0.0250387f $X=4.315 $Y=2.315
+ $X2=0 $Y2=0
cc_463 N_A_404_353#_c_442_n N_A_700_451#_c_1046_n 0.0146794f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_464 N_A_404_353#_c_443_n N_A_700_451#_c_1046_n 0.00278132f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_465 N_A_404_353#_c_427_n N_A_700_451#_c_1046_n 0.0197784f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_466 N_A_404_353#_M1029_g N_A_700_451#_c_1047_n 0.0157606f $X=4.145 $Y=0.445
+ $X2=0 $Y2=0
cc_467 N_A_404_353#_c_427_n N_A_700_451#_c_1047_n 0.0205948f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_468 N_A_404_353#_c_428_n N_A_700_451#_c_1047_n 0.00124789f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_469 N_A_404_353#_M1029_g N_A_700_451#_c_1048_n 0.00402648f $X=4.145 $Y=0.445
+ $X2=0 $Y2=0
cc_470 N_A_404_353#_c_427_n N_A_700_451#_c_1048_n 0.0119874f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_471 N_A_404_353#_c_428_n N_A_700_451#_c_1048_n 0.00120368f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_472 N_A_404_353#_c_427_n N_A_700_451#_c_1050_n 0.0141315f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_473 N_A_404_353#_c_428_n N_A_700_451#_c_1050_n 0.00140147f $X=4.235 $Y=1.29
+ $X2=0 $Y2=0
cc_474 N_A_404_353#_c_431_n N_VPWR_c_1269_n 0.00186631f $X=2.095 $Y=1.915 $X2=0
+ $Y2=0
cc_475 N_A_404_353#_M1033_g N_VPWR_c_1269_n 0.0054895f $X=3.065 $Y=2.675 $X2=0
+ $Y2=0
cc_476 N_A_404_353#_M1030_g N_VPWR_c_1269_n 0.0035787f $X=3.425 $Y=2.675 $X2=0
+ $Y2=0
cc_477 N_A_404_353#_c_454_p N_VPWR_c_1269_n 0.0597375f $X=4.23 $Y=2.99 $X2=0
+ $Y2=0
cc_478 N_A_404_353#_c_559_p N_VPWR_c_1269_n 0.00950638f $X=3.355 $Y=2.99 $X2=0
+ $Y2=0
cc_479 N_A_404_353#_c_431_n N_VPWR_c_1264_n 7.40383e-19 $X=2.095 $Y=1.915 $X2=0
+ $Y2=0
cc_480 N_A_404_353#_M1033_g N_VPWR_c_1264_n 0.00632399f $X=3.065 $Y=2.675 $X2=0
+ $Y2=0
cc_481 N_A_404_353#_M1030_g N_VPWR_c_1264_n 0.00491941f $X=3.425 $Y=2.675 $X2=0
+ $Y2=0
cc_482 N_A_404_353#_c_454_p N_VPWR_c_1264_n 0.00827896f $X=4.23 $Y=2.99 $X2=0
+ $Y2=0
cc_483 N_A_404_353#_c_559_p N_VPWR_c_1264_n 0.00158213f $X=3.355 $Y=2.99 $X2=0
+ $Y2=0
cc_484 N_A_404_353#_c_431_n N_A_217_130#_c_1370_n 0.00691294f $X=2.095 $Y=1.915
+ $X2=0 $Y2=0
cc_485 N_A_404_353#_c_431_n N_A_217_130#_c_1372_n 0.018472f $X=2.095 $Y=1.915
+ $X2=0 $Y2=0
cc_486 N_A_404_353#_c_433_n N_A_217_130#_c_1372_n 0.00378401f $X=2.99 $Y=1.84
+ $X2=0 $Y2=0
cc_487 N_A_404_353#_c_434_n N_A_217_130#_c_1372_n 7.54835e-19 $X=2.385 $Y=1.84
+ $X2=0 $Y2=0
cc_488 N_A_404_353#_c_431_n N_A_217_130#_c_1373_n 0.00151145f $X=2.095 $Y=1.915
+ $X2=0 $Y2=0
cc_489 N_A_404_353#_c_433_n N_A_217_130#_c_1363_n 0.00245853f $X=2.99 $Y=1.84
+ $X2=0 $Y2=0
cc_490 N_A_404_353#_c_442_n N_A_217_130#_c_1363_n 0.0256985f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_491 N_A_404_353#_c_443_n N_A_217_130#_c_1363_n 0.00509482f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_492 N_A_404_353#_M1034_g N_A_217_130#_c_1364_n 0.00100387f $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_493 N_A_404_353#_M1034_g N_A_217_130#_c_1365_n 0.00212033f $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_494 N_A_404_353#_c_434_n N_A_217_130#_c_1368_n 0.00691294f $X=2.385 $Y=1.84
+ $X2=0 $Y2=0
cc_495 N_A_404_353#_c_431_n N_A_217_130#_c_1375_n 0.00631383f $X=2.095 $Y=1.915
+ $X2=0 $Y2=0
cc_496 N_A_404_353#_c_433_n N_A_217_130#_c_1375_n 9.53814e-19 $X=2.99 $Y=1.84
+ $X2=0 $Y2=0
cc_497 N_A_404_353#_M1033_g N_A_217_130#_c_1375_n 0.00567922f $X=3.065 $Y=2.675
+ $X2=0 $Y2=0
cc_498 N_A_404_353#_M1030_g N_A_217_130#_c_1375_n 7.40975e-19 $X=3.425 $Y=2.675
+ $X2=0 $Y2=0
cc_499 N_A_404_353#_c_437_n N_A_217_130#_c_1375_n 0.0268941f $X=3.27 $Y=2.905
+ $X2=0 $Y2=0
cc_500 N_A_404_353#_c_431_n N_A_217_130#_c_1369_n 7.47374e-19 $X=2.095 $Y=1.915
+ $X2=0 $Y2=0
cc_501 N_A_404_353#_M1034_g N_A_217_130#_c_1369_n 8.84538e-19 $X=2.31 $Y=1.08
+ $X2=0 $Y2=0
cc_502 N_A_404_353#_c_433_n N_A_217_130#_c_1369_n 0.0138544f $X=2.99 $Y=1.84
+ $X2=0 $Y2=0
cc_503 N_A_404_353#_c_437_n N_A_217_130#_c_1369_n 0.00774201f $X=3.27 $Y=2.905
+ $X2=0 $Y2=0
cc_504 N_A_404_353#_c_442_n N_A_217_130#_c_1369_n 0.0242394f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_505 N_A_404_353#_c_443_n N_A_217_130#_c_1369_n 0.00806041f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_506 N_A_404_353#_M1033_g N_A_217_130#_c_1377_n 0.00412778f $X=3.065 $Y=2.675
+ $X2=0 $Y2=0
cc_507 N_A_404_353#_c_559_p N_A_217_130#_c_1377_n 0.00695601f $X=3.355 $Y=2.99
+ $X2=0 $Y2=0
cc_508 N_A_404_353#_c_559_p A_628_451# 9.38685e-19 $X=3.355 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_509 N_A_404_353#_c_454_p A_830_419# 0.00157878f $X=4.23 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_510 N_A_404_353#_c_422_n A_830_419# 0.00228171f $X=4.315 $Y=2.315 $X2=-0.19
+ $Y2=-0.245
cc_511 N_A_404_353#_c_455_p A_830_419# 0.00533605f $X=4.315 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_512 N_A_404_353#_c_458_p A_830_419# 0.00184923f $X=4.315 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_513 N_A_404_353#_c_439_n N_KAPWR_M1000_d 0.00511971f $X=7.92 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_514 N_A_404_353#_c_439_n N_KAPWR_M1002_d 0.0082631f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_515 N_A_404_353#_c_454_p N_KAPWR_c_1479_n 0.0109183f $X=4.23 $Y=2.99 $X2=0
+ $Y2=0
cc_516 N_A_404_353#_c_455_p N_KAPWR_c_1479_n 0.0127651f $X=4.315 $Y=2.905 $X2=0
+ $Y2=0
cc_517 N_A_404_353#_c_439_n N_KAPWR_c_1479_n 0.0349531f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_518 N_A_404_353#_c_439_n N_KAPWR_c_1480_n 0.0229025f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_519 N_A_404_353#_M1007_d N_KAPWR_c_1482_n 0.00346453f $X=8.975 $Y=2.33 $X2=0
+ $Y2=0
cc_520 N_A_404_353#_c_431_n N_KAPWR_c_1482_n 0.00750852f $X=2.095 $Y=1.915 $X2=0
+ $Y2=0
cc_521 N_A_404_353#_M1033_g N_KAPWR_c_1482_n 0.00427309f $X=3.065 $Y=2.675 $X2=0
+ $Y2=0
cc_522 N_A_404_353#_M1030_g N_KAPWR_c_1482_n 0.00849996f $X=3.425 $Y=2.675 $X2=0
+ $Y2=0
cc_523 N_A_404_353#_c_437_n N_KAPWR_c_1482_n 0.0205631f $X=3.27 $Y=2.905 $X2=0
+ $Y2=0
cc_524 N_A_404_353#_c_454_p N_KAPWR_c_1482_n 0.0282706f $X=4.23 $Y=2.99 $X2=0
+ $Y2=0
cc_525 N_A_404_353#_c_559_p N_KAPWR_c_1482_n 0.00253288f $X=3.355 $Y=2.99 $X2=0
+ $Y2=0
cc_526 N_A_404_353#_c_455_p N_KAPWR_c_1482_n 0.0225443f $X=4.315 $Y=2.905 $X2=0
+ $Y2=0
cc_527 N_A_404_353#_c_439_n N_KAPWR_c_1482_n 0.132972f $X=7.92 $Y=2.4 $X2=0
+ $Y2=0
cc_528 N_A_404_353#_c_442_n N_KAPWR_c_1482_n 0.00458104f $X=3.19 $Y=1.93 $X2=0
+ $Y2=0
cc_529 N_A_404_353#_c_439_n A_1246_341# 0.00300846f $X=7.92 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_530 N_A_404_353#_M1034_g N_VGND_c_1593_n 0.00718751f $X=2.31 $Y=1.08 $X2=0
+ $Y2=0
cc_531 N_A_404_353#_c_434_n N_VGND_c_1593_n 0.00440367f $X=2.385 $Y=1.84 $X2=0
+ $Y2=0
cc_532 N_A_404_353#_c_425_n N_VGND_c_1596_n 0.00442395f $X=9.065 $Y=1.225 $X2=0
+ $Y2=0
cc_533 N_A_404_353#_M1029_g N_VGND_c_1602_n 0.00357877f $X=4.145 $Y=0.445 $X2=0
+ $Y2=0
cc_534 N_A_404_353#_M1029_g N_VGND_c_1607_n 0.0055095f $X=4.145 $Y=0.445 $X2=0
+ $Y2=0
cc_535 N_A_404_353#_c_430_n N_VGND_c_1607_n 0.0111482f $X=8.755 $Y=1.08 $X2=0
+ $Y2=0
cc_536 N_A_404_353#_c_425_n A_1798_174# 0.00552058f $X=9.065 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_537 N_A_434_405#_M1014_g N_A_878_357#_M1000_g 0.0385944f $X=4.025 $Y=2.595
+ $X2=0 $Y2=0
cc_538 N_A_434_405#_c_625_n N_A_878_357#_c_720_n 0.0402061f $X=3.67 $Y=1.695
+ $X2=0 $Y2=0
cc_539 N_A_434_405#_M1014_g N_A_700_451#_c_1056_n 0.00517877f $X=4.025 $Y=2.595
+ $X2=0 $Y2=0
cc_540 N_A_434_405#_c_625_n N_A_700_451#_c_1056_n 0.00521563f $X=3.67 $Y=1.695
+ $X2=0 $Y2=0
cc_541 N_A_434_405#_M1014_g N_A_700_451#_c_1082_n 0.00919568f $X=4.025 $Y=2.595
+ $X2=0 $Y2=0
cc_542 N_A_434_405#_c_618_n N_A_700_451#_c_1065_n 2.29836e-19 $X=3.26 $Y=0.985
+ $X2=0 $Y2=0
cc_543 N_A_434_405#_M1021_g N_A_700_451#_c_1065_n 0.00361646f $X=3.62 $Y=0.555
+ $X2=0 $Y2=0
cc_544 N_A_434_405#_c_618_n N_A_700_451#_c_1046_n 2.05778e-19 $X=3.26 $Y=0.985
+ $X2=0 $Y2=0
cc_545 N_A_434_405#_M1021_g N_A_700_451#_c_1046_n 0.00518012f $X=3.62 $Y=0.555
+ $X2=0 $Y2=0
cc_546 N_A_434_405#_c_621_n N_A_700_451#_c_1046_n 0.00560785f $X=3.67 $Y=1.545
+ $X2=0 $Y2=0
cc_547 N_A_434_405#_M1014_g N_A_700_451#_c_1046_n 0.0029423f $X=4.025 $Y=2.595
+ $X2=0 $Y2=0
cc_548 N_A_434_405#_c_624_n N_A_700_451#_c_1046_n 0.00529177f $X=3.645 $Y=1.24
+ $X2=0 $Y2=0
cc_549 N_A_434_405#_c_625_n N_A_700_451#_c_1046_n 0.0205432f $X=3.67 $Y=1.695
+ $X2=0 $Y2=0
cc_550 N_A_434_405#_c_625_n N_A_700_451#_c_1047_n 4.6985e-19 $X=3.67 $Y=1.695
+ $X2=0 $Y2=0
cc_551 N_A_434_405#_M1014_g N_VPWR_c_1269_n 0.00596462f $X=4.025 $Y=2.595 $X2=0
+ $Y2=0
cc_552 N_A_434_405#_M1014_g N_VPWR_c_1264_n 0.00713172f $X=4.025 $Y=2.595 $X2=0
+ $Y2=0
cc_553 N_A_434_405#_c_633_n N_A_217_130#_c_1370_n 0.0119015f $X=2.31 $Y=2.17
+ $X2=0 $Y2=0
cc_554 N_A_434_405#_M1010_d N_A_217_130#_c_1372_n 0.0029807f $X=2.17 $Y=2.025
+ $X2=0 $Y2=0
cc_555 N_A_434_405#_c_633_n N_A_217_130#_c_1372_n 0.023665f $X=2.31 $Y=2.17
+ $X2=0 $Y2=0
cc_556 N_A_434_405#_c_621_n N_A_217_130#_c_1363_n 0.00383217f $X=3.67 $Y=1.545
+ $X2=0 $Y2=0
cc_557 N_A_434_405#_c_622_n N_A_217_130#_c_1363_n 0.00540278f $X=3.185 $Y=1.15
+ $X2=0 $Y2=0
cc_558 N_A_434_405#_c_627_n N_A_217_130#_c_1363_n 0.0225369f $X=2.995 $Y=1.15
+ $X2=0 $Y2=0
cc_559 N_A_434_405#_c_622_n N_A_217_130#_c_1364_n 2.55481e-19 $X=3.185 $Y=1.15
+ $X2=0 $Y2=0
cc_560 N_A_434_405#_c_628_n N_A_217_130#_c_1364_n 0.0148633f $X=2.33 $Y=1.48
+ $X2=0 $Y2=0
cc_561 N_A_434_405#_c_629_n N_A_217_130#_c_1364_n 0.0146974f $X=2.69 $Y=1.052
+ $X2=0 $Y2=0
cc_562 N_A_434_405#_c_618_n N_A_217_130#_c_1365_n 0.00993134f $X=3.26 $Y=0.985
+ $X2=0 $Y2=0
cc_563 N_A_434_405#_c_622_n N_A_217_130#_c_1365_n 0.00672631f $X=3.185 $Y=1.15
+ $X2=0 $Y2=0
cc_564 N_A_434_405#_c_627_n N_A_217_130#_c_1365_n 0.0196048f $X=2.995 $Y=1.15
+ $X2=0 $Y2=0
cc_565 N_A_434_405#_c_618_n N_A_217_130#_c_1366_n 0.00507658f $X=3.26 $Y=0.985
+ $X2=0 $Y2=0
cc_566 N_A_434_405#_c_619_n N_A_217_130#_c_1366_n 0.00749863f $X=3.545 $Y=1.24
+ $X2=0 $Y2=0
cc_567 N_A_434_405#_M1021_g N_A_217_130#_c_1366_n 0.0019792f $X=3.62 $Y=0.555
+ $X2=0 $Y2=0
cc_568 N_A_434_405#_c_621_n N_A_217_130#_c_1366_n 0.00227676f $X=3.67 $Y=1.545
+ $X2=0 $Y2=0
cc_569 N_A_434_405#_c_623_n N_A_217_130#_c_1366_n 0.00740802f $X=3.26 $Y=1.15
+ $X2=0 $Y2=0
cc_570 N_A_434_405#_c_627_n N_A_217_130#_c_1366_n 0.020415f $X=2.995 $Y=1.15
+ $X2=0 $Y2=0
cc_571 N_A_434_405#_c_629_n N_A_217_130#_c_1366_n 0.00372624f $X=2.69 $Y=1.052
+ $X2=0 $Y2=0
cc_572 N_A_434_405#_c_626_n N_A_217_130#_c_1368_n 0.0119015f $X=2.33 $Y=1.665
+ $X2=0 $Y2=0
cc_573 N_A_434_405#_c_633_n N_A_217_130#_c_1375_n 0.0290891f $X=2.31 $Y=2.17
+ $X2=0 $Y2=0
cc_574 N_A_434_405#_c_626_n N_A_217_130#_c_1369_n 0.0290891f $X=2.33 $Y=1.665
+ $X2=0 $Y2=0
cc_575 N_A_434_405#_M1014_g N_KAPWR_c_1479_n 2.97501e-19 $X=4.025 $Y=2.595 $X2=0
+ $Y2=0
cc_576 N_A_434_405#_M1014_g N_KAPWR_c_1482_n 0.0134276f $X=4.025 $Y=2.595 $X2=0
+ $Y2=0
cc_577 N_A_434_405#_c_626_n N_VGND_c_1593_n 0.00164722f $X=2.33 $Y=1.665 $X2=0
+ $Y2=0
cc_578 N_A_434_405#_c_628_n N_VGND_c_1593_n 0.00392482f $X=2.33 $Y=1.48 $X2=0
+ $Y2=0
cc_579 N_A_434_405#_c_629_n N_VGND_c_1593_n 0.0312639f $X=2.69 $Y=1.052 $X2=0
+ $Y2=0
cc_580 N_A_434_405#_c_618_n N_VGND_c_1602_n 0.00357877f $X=3.26 $Y=0.985 $X2=0
+ $Y2=0
cc_581 N_A_434_405#_M1021_g N_VGND_c_1602_n 0.00357877f $X=3.62 $Y=0.555 $X2=0
+ $Y2=0
cc_582 N_A_434_405#_c_618_n N_VGND_c_1607_n 0.0066108f $X=3.26 $Y=0.985 $X2=0
+ $Y2=0
cc_583 N_A_434_405#_M1021_g N_VGND_c_1607_n 0.00546664f $X=3.62 $Y=0.555 $X2=0
+ $Y2=0
cc_584 N_A_878_357#_c_727_n N_A_1294_315#_M1002_g 0.0170508f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_585 N_A_878_357#_c_727_n N_A_1294_315#_c_823_n 4.52366e-19 $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_586 N_A_878_357#_c_721_n N_GATE_M1013_g 0.00143855f $X=8.04 $Y=0.8 $X2=0
+ $Y2=0
cc_587 N_A_878_357#_c_722_n N_GATE_M1013_g 0.00137597f $X=8.04 $Y=0.655 $X2=0
+ $Y2=0
cc_588 N_A_878_357#_c_727_n N_A_700_451#_M1026_s 0.00940891f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_589 N_A_878_357#_c_722_n N_A_700_451#_M1022_g 0.00366272f $X=8.04 $Y=0.655
+ $X2=0 $Y2=0
cc_590 N_A_878_357#_c_723_n N_A_700_451#_M1022_g 9.90115e-19 $X=7.585 $Y=1.685
+ $X2=0 $Y2=0
cc_591 N_A_878_357#_c_727_n N_A_700_451#_M1009_g 0.0153821f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_592 N_A_878_357#_c_729_n N_A_700_451#_M1009_g 0.0167434f $X=7.585 $Y=1.915
+ $X2=0 $Y2=0
cc_593 N_A_878_357#_c_721_n N_A_700_451#_c_1039_n 0.00206157f $X=8.04 $Y=0.8
+ $X2=0 $Y2=0
cc_594 N_A_878_357#_c_722_n N_A_700_451#_c_1039_n 0.00793966f $X=8.04 $Y=0.655
+ $X2=0 $Y2=0
cc_595 N_A_878_357#_c_729_n N_A_700_451#_c_1041_n 0.00451683f $X=7.585 $Y=1.915
+ $X2=0 $Y2=0
cc_596 N_A_878_357#_c_723_n N_A_700_451#_c_1041_n 0.00948886f $X=7.585 $Y=1.685
+ $X2=0 $Y2=0
cc_597 N_A_878_357#_c_721_n N_A_700_451#_M1006_g 0.0102892f $X=8.04 $Y=0.8 $X2=0
+ $Y2=0
cc_598 N_A_878_357#_c_722_n N_A_700_451#_M1006_g 0.0119381f $X=8.04 $Y=0.655
+ $X2=0 $Y2=0
cc_599 N_A_878_357#_c_723_n N_A_700_451#_M1006_g 0.00844567f $X=7.585 $Y=1.685
+ $X2=0 $Y2=0
cc_600 N_A_878_357#_M1000_g N_A_700_451#_c_1056_n 5.26479e-19 $X=4.515 $Y=2.595
+ $X2=0 $Y2=0
cc_601 N_A_878_357#_c_714_n N_A_700_451#_c_1047_n 0.00692275f $X=4.505 $Y=0.765
+ $X2=0 $Y2=0
cc_602 N_A_878_357#_c_715_n N_A_700_451#_c_1047_n 0.00415937f $X=4.79 $Y=0.84
+ $X2=0 $Y2=0
cc_603 N_A_878_357#_c_716_n N_A_700_451#_c_1047_n 0.00844685f $X=4.58 $Y=0.84
+ $X2=0 $Y2=0
cc_604 N_A_878_357#_c_717_n N_A_700_451#_c_1047_n 0.00121257f $X=4.865 $Y=0.765
+ $X2=0 $Y2=0
cc_605 N_A_878_357#_c_715_n N_A_700_451#_c_1048_n 0.00380937f $X=4.79 $Y=0.84
+ $X2=0 $Y2=0
cc_606 N_A_878_357#_c_716_n N_A_700_451#_c_1048_n 4.76463e-19 $X=4.58 $Y=0.84
+ $X2=0 $Y2=0
cc_607 N_A_878_357#_c_718_n N_A_700_451#_c_1048_n 0.00833389f $X=4.865 $Y=1.605
+ $X2=0 $Y2=0
cc_608 N_A_878_357#_c_715_n N_A_700_451#_c_1049_n 0.00103653f $X=4.79 $Y=0.84
+ $X2=0 $Y2=0
cc_609 N_A_878_357#_c_718_n N_A_700_451#_c_1049_n 0.0160375f $X=4.865 $Y=1.605
+ $X2=0 $Y2=0
cc_610 N_A_878_357#_c_725_n N_A_700_451#_c_1049_n 0.0173158f $X=4.805 $Y=1.77
+ $X2=0 $Y2=0
cc_611 N_A_878_357#_c_720_n N_A_700_451#_c_1049_n 0.00125423f $X=4.805 $Y=1.77
+ $X2=0 $Y2=0
cc_612 N_A_878_357#_c_727_n N_A_700_451#_c_1049_n 0.00588557f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_613 N_A_878_357#_c_725_n N_A_700_451#_c_1050_n 0.00865844f $X=4.805 $Y=1.77
+ $X2=0 $Y2=0
cc_614 N_A_878_357#_c_720_n N_A_700_451#_c_1050_n 0.00407319f $X=4.805 $Y=1.77
+ $X2=0 $Y2=0
cc_615 N_A_878_357#_c_727_n N_A_700_451#_c_1058_n 0.0114256f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_616 N_A_878_357#_c_727_n N_A_700_451#_c_1059_n 0.0446024f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_617 N_A_878_357#_c_718_n N_A_700_451#_c_1051_n 0.00574809f $X=4.865 $Y=1.605
+ $X2=0 $Y2=0
cc_618 N_A_878_357#_c_720_n N_A_700_451#_c_1051_n 7.51326e-19 $X=4.805 $Y=1.77
+ $X2=0 $Y2=0
cc_619 N_A_878_357#_c_727_n N_A_700_451#_c_1051_n 0.00812318f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_620 N_A_878_357#_c_725_n N_A_700_451#_c_1061_n 0.00557104f $X=4.805 $Y=1.77
+ $X2=0 $Y2=0
cc_621 N_A_878_357#_c_720_n N_A_700_451#_c_1061_n 0.00305165f $X=4.805 $Y=1.77
+ $X2=0 $Y2=0
cc_622 N_A_878_357#_c_727_n N_A_700_451#_c_1061_n 0.0253593f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_623 N_A_878_357#_c_727_n N_A_700_451#_c_1052_n 0.0116513f $X=7.42 $Y=2.06
+ $X2=0 $Y2=0
cc_624 N_A_878_357#_c_723_n N_A_700_451#_c_1052_n 0.0299337f $X=7.585 $Y=1.685
+ $X2=0 $Y2=0
cc_625 N_A_878_357#_c_727_n N_A_700_451#_c_1053_n 3.97e-19 $X=7.42 $Y=2.06 $X2=0
+ $Y2=0
cc_626 N_A_878_357#_c_723_n N_A_700_451#_c_1053_n 0.00914197f $X=7.585 $Y=1.685
+ $X2=0 $Y2=0
cc_627 N_A_878_357#_M1000_g N_VPWR_c_1269_n 0.00922542f $X=4.515 $Y=2.595 $X2=0
+ $Y2=0
cc_628 N_A_878_357#_M1000_g N_VPWR_c_1264_n 0.00871855f $X=4.515 $Y=2.595 $X2=0
+ $Y2=0
cc_629 N_A_878_357#_c_728_n N_KAPWR_M1000_d 0.00271531f $X=4.97 $Y=2.06
+ $X2=-0.19 $Y2=-0.245
cc_630 N_A_878_357#_c_727_n N_KAPWR_M1002_d 0.00998057f $X=7.42 $Y=2.06 $X2=0
+ $Y2=0
cc_631 N_A_878_357#_M1000_g N_KAPWR_c_1479_n 0.00695659f $X=4.515 $Y=2.595 $X2=0
+ $Y2=0
cc_632 N_A_878_357#_M1009_d N_KAPWR_c_1482_n 0.00255308f $X=7.445 $Y=1.705 $X2=0
+ $Y2=0
cc_633 N_A_878_357#_M1000_g N_KAPWR_c_1482_n 0.00355816f $X=4.515 $Y=2.595 $X2=0
+ $Y2=0
cc_634 N_A_878_357#_c_727_n A_1246_341# 0.00317058f $X=7.42 $Y=2.06 $X2=-0.19
+ $Y2=-0.245
cc_635 N_A_878_357#_c_714_n N_VGND_c_1602_n 0.00357877f $X=4.505 $Y=0.765 $X2=0
+ $Y2=0
cc_636 N_A_878_357#_c_717_n N_VGND_c_1602_n 0.00357877f $X=4.865 $Y=0.765 $X2=0
+ $Y2=0
cc_637 N_A_878_357#_c_722_n N_VGND_c_1604_n 0.0148095f $X=8.04 $Y=0.655 $X2=0
+ $Y2=0
cc_638 N_A_878_357#_c_714_n N_VGND_c_1607_n 0.00504318f $X=4.505 $Y=0.765 $X2=0
+ $Y2=0
cc_639 N_A_878_357#_c_717_n N_VGND_c_1607_n 0.00651363f $X=4.865 $Y=0.765 $X2=0
+ $Y2=0
cc_640 N_A_878_357#_c_721_n N_VGND_c_1607_n 0.00898734f $X=8.04 $Y=0.8 $X2=0
+ $Y2=0
cc_641 N_A_878_357#_c_722_n N_VGND_c_1607_n 0.0107179f $X=8.04 $Y=0.655 $X2=0
+ $Y2=0
cc_642 N_A_878_357#_c_717_n N_A_988_47#_c_1747_n 0.0105019f $X=4.865 $Y=0.765
+ $X2=0 $Y2=0
cc_643 N_A_878_357#_c_718_n N_A_988_47#_c_1748_n 0.00640131f $X=4.865 $Y=1.605
+ $X2=0 $Y2=0
cc_644 N_A_1294_315#_c_832_n N_GATE_c_923_n 6.01727e-19 $X=10.255 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_645 N_A_1294_315#_c_831_n N_GATE_M1007_g 0.00418666f $X=8.345 $Y=2.745 $X2=0
+ $Y2=0
cc_646 N_A_1294_315#_c_832_n N_GATE_M1007_g 0.017405f $X=10.255 $Y=2.405 $X2=0
+ $Y2=0
cc_647 N_A_1294_315#_c_836_n N_GATE_M1007_g 0.00586674f $X=8.215 $Y=2.91 $X2=0
+ $Y2=0
cc_648 N_A_1294_315#_c_837_n N_GATE_M1007_g 0.0019821f $X=8.345 $Y=2.91 $X2=0
+ $Y2=0
cc_649 N_A_1294_315#_c_832_n N_GATE_c_927_n 3.64746e-19 $X=10.255 $Y=2.405 $X2=0
+ $Y2=0
cc_650 N_A_1294_315#_c_832_n GATE 0.0141557f $X=10.255 $Y=2.405 $X2=0 $Y2=0
cc_651 N_A_1294_315#_c_833_n GATE 0.0119858f $X=8.43 $Y=2.405 $X2=0 $Y2=0
cc_652 N_A_1294_315#_c_832_n N_GATE_c_929_n 0.00127918f $X=10.255 $Y=2.405 $X2=0
+ $Y2=0
cc_653 N_A_1294_315#_c_833_n N_GATE_c_929_n 7.95902e-19 $X=8.43 $Y=2.405 $X2=0
+ $Y2=0
cc_654 N_A_1294_315#_c_836_n N_GATE_c_929_n 0.00133251f $X=8.215 $Y=2.91 $X2=0
+ $Y2=0
cc_655 N_A_1294_315#_c_832_n N_SLEEP_B_M1003_g 0.0150945f $X=10.255 $Y=2.405
+ $X2=0 $Y2=0
cc_656 N_A_1294_315#_c_825_n N_SLEEP_B_M1032_g 0.00423479f $X=10.42 $Y=1.985
+ $X2=0 $Y2=0
cc_657 N_A_1294_315#_c_826_n N_SLEEP_B_M1032_g 0.00132871f $X=10.43 $Y=0.865
+ $X2=0 $Y2=0
cc_658 N_A_1294_315#_c_832_n N_SLEEP_B_c_971_n 0.00784383f $X=10.255 $Y=2.405
+ $X2=0 $Y2=0
cc_659 N_A_1294_315#_c_832_n N_SLEEP_B_M1001_g 0.0198546f $X=10.255 $Y=2.405
+ $X2=0 $Y2=0
cc_660 N_A_1294_315#_c_825_n N_SLEEP_B_M1001_g 0.0323005f $X=10.42 $Y=1.985
+ $X2=0 $Y2=0
cc_661 N_A_1294_315#_c_835_n N_SLEEP_B_M1001_g 0.0103821f $X=10.42 $Y=2.695
+ $X2=0 $Y2=0
cc_662 N_A_1294_315#_c_868_p N_SLEEP_B_M1001_g 3.84191e-19 $X=10.38 $Y=2.405
+ $X2=0 $Y2=0
cc_663 N_A_1294_315#_c_825_n N_SLEEP_B_c_973_n 0.0134406f $X=10.42 $Y=1.985
+ $X2=0 $Y2=0
cc_664 N_A_1294_315#_c_825_n N_SLEEP_B_M1023_g 0.0154343f $X=10.42 $Y=1.985
+ $X2=0 $Y2=0
cc_665 N_A_1294_315#_c_826_n N_SLEEP_B_M1023_g 0.0102235f $X=10.43 $Y=0.865
+ $X2=0 $Y2=0
cc_666 N_A_1294_315#_c_826_n N_SLEEP_B_M1015_g 0.00125175f $X=10.43 $Y=0.865
+ $X2=0 $Y2=0
cc_667 N_A_1294_315#_c_825_n N_SLEEP_B_c_976_n 0.00787953f $X=10.42 $Y=1.985
+ $X2=0 $Y2=0
cc_668 N_A_1294_315#_c_825_n N_SLEEP_B_c_978_n 0.00182139f $X=10.42 $Y=1.985
+ $X2=0 $Y2=0
cc_669 N_A_1294_315#_c_825_n N_SLEEP_B_c_979_n 0.0512609f $X=10.42 $Y=1.985
+ $X2=0 $Y2=0
cc_670 N_A_1294_315#_M1020_g N_A_700_451#_M1022_g 0.014405f $X=6.77 $Y=0.845
+ $X2=0 $Y2=0
cc_671 N_A_1294_315#_c_823_n N_A_700_451#_M1009_g 0.0376797f $X=6.77 $Y=1.345
+ $X2=0 $Y2=0
cc_672 N_A_1294_315#_c_829_n N_A_700_451#_M1009_g 0.0143838f $X=8.05 $Y=3.15
+ $X2=0 $Y2=0
cc_673 N_A_1294_315#_c_836_n N_A_700_451#_M1009_g 0.00148042f $X=8.215 $Y=2.91
+ $X2=0 $Y2=0
cc_674 N_A_1294_315#_c_837_n N_A_700_451#_M1009_g 5.6599e-19 $X=8.345 $Y=2.91
+ $X2=0 $Y2=0
cc_675 N_A_1294_315#_c_826_n N_A_700_451#_c_1039_n 0.00635386f $X=10.43 $Y=0.865
+ $X2=0 $Y2=0
cc_676 N_A_1294_315#_c_823_n N_A_700_451#_c_1059_n 0.0256105f $X=6.77 $Y=1.345
+ $X2=0 $Y2=0
cc_677 N_A_1294_315#_M1020_g N_A_700_451#_c_1052_n 0.00446736f $X=6.77 $Y=0.845
+ $X2=0 $Y2=0
cc_678 N_A_1294_315#_c_823_n N_A_700_451#_c_1053_n 6.35235e-19 $X=6.77 $Y=1.345
+ $X2=0 $Y2=0
cc_679 N_A_1294_315#_M1020_g N_A_700_451#_c_1053_n 0.0160708f $X=6.77 $Y=0.845
+ $X2=0 $Y2=0
cc_680 N_A_1294_315#_c_830_n N_VPWR_c_1269_n 0.0602576f $X=6.72 $Y=3.15 $X2=0
+ $Y2=0
cc_681 N_A_1294_315#_c_835_n N_VPWR_c_1269_n 0.0077512f $X=10.42 $Y=2.695 $X2=0
+ $Y2=0
cc_682 N_A_1294_315#_c_837_n N_VPWR_c_1269_n 0.0246005f $X=8.345 $Y=2.91 $X2=0
+ $Y2=0
cc_683 N_A_1294_315#_c_829_n N_VPWR_c_1264_n 0.0252569f $X=8.05 $Y=3.15 $X2=0
+ $Y2=0
cc_684 N_A_1294_315#_c_830_n N_VPWR_c_1264_n 0.00807098f $X=6.72 $Y=3.15 $X2=0
+ $Y2=0
cc_685 N_A_1294_315#_c_835_n N_VPWR_c_1264_n 9.54636e-19 $X=10.42 $Y=2.695 $X2=0
+ $Y2=0
cc_686 N_A_1294_315#_c_836_n N_VPWR_c_1264_n 0.00905989f $X=8.215 $Y=2.91 $X2=0
+ $Y2=0
cc_687 N_A_1294_315#_c_837_n N_VPWR_c_1264_n 0.0029545f $X=8.345 $Y=2.91 $X2=0
+ $Y2=0
cc_688 N_A_1294_315#_c_832_n N_KAPWR_M1007_s 0.00334554f $X=10.255 $Y=2.405
+ $X2=0 $Y2=0
cc_689 N_A_1294_315#_c_832_n N_KAPWR_M1003_d 0.0132937f $X=10.255 $Y=2.405 $X2=0
+ $Y2=0
cc_690 N_A_1294_315#_M1002_g N_KAPWR_c_1480_n 0.00953766f $X=6.595 $Y=2.205
+ $X2=0 $Y2=0
cc_691 N_A_1294_315#_c_829_n N_KAPWR_c_1480_n 0.0075395f $X=8.05 $Y=3.15 $X2=0
+ $Y2=0
cc_692 N_A_1294_315#_c_831_n N_KAPWR_c_1481_n 0.00605644f $X=8.345 $Y=2.745
+ $X2=0 $Y2=0
cc_693 N_A_1294_315#_c_832_n N_KAPWR_c_1481_n 0.0214598f $X=10.255 $Y=2.405
+ $X2=0 $Y2=0
cc_694 N_A_1294_315#_c_836_n N_KAPWR_c_1481_n 7.24985e-19 $X=8.215 $Y=2.91 $X2=0
+ $Y2=0
cc_695 N_A_1294_315#_c_837_n N_KAPWR_c_1481_n 0.0180827f $X=8.345 $Y=2.91 $X2=0
+ $Y2=0
cc_696 N_A_1294_315#_M1001_d N_KAPWR_c_1482_n 0.00246912f $X=10.28 $Y=1.84 $X2=0
+ $Y2=0
cc_697 N_A_1294_315#_M1002_g N_KAPWR_c_1482_n 0.0128108f $X=6.595 $Y=2.205 $X2=0
+ $Y2=0
cc_698 N_A_1294_315#_c_829_n N_KAPWR_c_1482_n 0.00790518f $X=8.05 $Y=3.15 $X2=0
+ $Y2=0
cc_699 N_A_1294_315#_c_831_n N_KAPWR_c_1482_n 0.00830564f $X=8.345 $Y=2.745
+ $X2=0 $Y2=0
cc_700 N_A_1294_315#_c_832_n N_KAPWR_c_1482_n 0.0411052f $X=10.255 $Y=2.405
+ $X2=0 $Y2=0
cc_701 N_A_1294_315#_c_835_n N_KAPWR_c_1482_n 0.0301878f $X=10.42 $Y=2.695 $X2=0
+ $Y2=0
cc_702 N_A_1294_315#_c_836_n N_KAPWR_c_1482_n 0.00472287f $X=8.215 $Y=2.91 $X2=0
+ $Y2=0
cc_703 N_A_1294_315#_c_837_n N_KAPWR_c_1482_n 0.021665f $X=8.345 $Y=2.91 $X2=0
+ $Y2=0
cc_704 N_A_1294_315#_c_832_n N_KAPWR_c_1483_n 0.0490226f $X=10.255 $Y=2.405
+ $X2=0 $Y2=0
cc_705 N_A_1294_315#_c_835_n N_KAPWR_c_1483_n 0.00711861f $X=10.42 $Y=2.695
+ $X2=0 $Y2=0
cc_706 N_A_1294_315#_M1020_g N_VGND_c_1594_n 4.28038e-19 $X=6.77 $Y=0.845 $X2=0
+ $Y2=0
cc_707 N_A_1294_315#_M1020_g N_VGND_c_1595_n 0.00908647f $X=6.77 $Y=0.845 $X2=0
+ $Y2=0
cc_708 N_A_1294_315#_c_826_n N_VGND_c_1596_n 0.0481932f $X=10.43 $Y=0.865 $X2=0
+ $Y2=0
cc_709 N_A_1294_315#_c_826_n N_VGND_c_1597_n 0.0151051f $X=10.43 $Y=0.865 $X2=0
+ $Y2=0
cc_710 N_A_1294_315#_c_826_n N_VGND_c_1599_n 0.00672647f $X=10.43 $Y=0.865 $X2=0
+ $Y2=0
cc_711 N_A_1294_315#_M1020_g N_VGND_c_1603_n 0.00340865f $X=6.77 $Y=0.845 $X2=0
+ $Y2=0
cc_712 N_A_1294_315#_M1020_g N_VGND_c_1607_n 0.00392009f $X=6.77 $Y=0.845 $X2=0
+ $Y2=0
cc_713 N_A_1294_315#_c_826_n N_VGND_c_1607_n 0.00885163f $X=10.43 $Y=0.865 $X2=0
+ $Y2=0
cc_714 N_A_1294_315#_c_823_n N_A_988_47#_c_1745_n 0.0027514f $X=6.77 $Y=1.345
+ $X2=0 $Y2=0
cc_715 N_A_1294_315#_M1020_g N_A_988_47#_c_1745_n 0.00374919f $X=6.77 $Y=0.845
+ $X2=0 $Y2=0
cc_716 N_A_1294_315#_M1020_g N_A_988_47#_c_1746_n 0.00191582f $X=6.77 $Y=0.845
+ $X2=0 $Y2=0
cc_717 N_GATE_M1013_g N_SLEEP_B_M1004_g 0.0240436f $X=8.915 $Y=1.08 $X2=0 $Y2=0
cc_718 N_GATE_M1007_g N_SLEEP_B_M1003_g 0.0234594f $X=8.9 $Y=2.65 $X2=0 $Y2=0
cc_719 N_GATE_c_927_n N_SLEEP_B_c_971_n 0.0240436f $X=8.907 $Y=1.555 $X2=0 $Y2=0
cc_720 N_GATE_M1013_g N_A_700_451#_c_1039_n 0.00470938f $X=8.915 $Y=1.08 $X2=0
+ $Y2=0
cc_721 N_GATE_M1007_g N_VPWR_c_1269_n 0.00295805f $X=8.9 $Y=2.65 $X2=0 $Y2=0
cc_722 N_GATE_M1007_g N_VPWR_c_1264_n 0.00332551f $X=8.9 $Y=2.65 $X2=0 $Y2=0
cc_723 N_GATE_M1007_g N_KAPWR_c_1481_n 0.01305f $X=8.9 $Y=2.65 $X2=0 $Y2=0
cc_724 GATE N_KAPWR_c_1482_n 8.41632e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_725 N_GATE_M1007_g N_KAPWR_c_1483_n 0.00203298f $X=8.9 $Y=2.65 $X2=0 $Y2=0
cc_726 N_GATE_M1013_g N_VGND_c_1607_n 9.3892e-19 $X=8.915 $Y=1.08 $X2=0 $Y2=0
cc_727 N_SLEEP_B_M1004_g N_A_700_451#_c_1039_n 0.00470938f $X=9.305 $Y=1.08
+ $X2=0 $Y2=0
cc_728 N_SLEEP_B_M1032_g N_A_700_451#_c_1039_n 0.00450393f $X=9.665 $Y=1.08
+ $X2=0 $Y2=0
cc_729 N_SLEEP_B_M1023_g N_A_700_451#_c_1039_n 0.0090052f $X=10.645 $Y=0.865
+ $X2=0 $Y2=0
cc_730 N_SLEEP_B_M1015_g N_A_700_451#_c_1039_n 0.00899129f $X=11.005 $Y=0.865
+ $X2=0 $Y2=0
cc_731 N_SLEEP_B_M1015_g N_A_700_451#_M1017_g 0.0187369f $X=11.005 $Y=0.865
+ $X2=0 $Y2=0
cc_732 N_SLEEP_B_M1015_g N_A_700_451#_M1027_g 0.00496133f $X=11.005 $Y=0.865
+ $X2=0 $Y2=0
cc_733 N_SLEEP_B_c_978_n N_A_700_451#_M1027_g 0.0054572f $X=10.89 $Y=1.645 $X2=0
+ $Y2=0
cc_734 N_SLEEP_B_c_979_n N_A_700_451#_M1027_g 3.89402e-19 $X=10.89 $Y=1.645
+ $X2=0 $Y2=0
cc_735 N_SLEEP_B_c_978_n N_A_2266_367#_c_1229_n 0.00470824f $X=10.89 $Y=1.645
+ $X2=0 $Y2=0
cc_736 N_SLEEP_B_c_979_n N_A_2266_367#_c_1229_n 0.02976f $X=10.89 $Y=1.645 $X2=0
+ $Y2=0
cc_737 N_SLEEP_B_M1015_g N_A_2266_367#_c_1225_n 0.00123641f $X=11.005 $Y=0.865
+ $X2=0 $Y2=0
cc_738 N_SLEEP_B_M1015_g N_A_2266_367#_c_1227_n 0.00511395f $X=11.005 $Y=0.865
+ $X2=0 $Y2=0
cc_739 N_SLEEP_B_c_979_n N_A_2266_367#_c_1227_n 0.0103351f $X=10.89 $Y=1.645
+ $X2=0 $Y2=0
cc_740 N_SLEEP_B_M1001_g N_VPWR_c_1269_n 0.00802751f $X=10.155 $Y=2.34 $X2=0
+ $Y2=0
cc_741 N_SLEEP_B_M1001_g N_VPWR_c_1264_n 0.00492612f $X=10.155 $Y=2.34 $X2=0
+ $Y2=0
cc_742 N_SLEEP_B_M1001_g N_KAPWR_c_1482_n 0.0100121f $X=10.155 $Y=2.34 $X2=0
+ $Y2=0
cc_743 N_SLEEP_B_c_979_n N_KAPWR_c_1482_n 0.0132757f $X=10.89 $Y=1.645 $X2=0
+ $Y2=0
cc_744 N_SLEEP_B_M1003_g N_KAPWR_c_1483_n 0.00462278f $X=9.445 $Y=2.16 $X2=0
+ $Y2=0
cc_745 N_SLEEP_B_M1001_g N_KAPWR_c_1483_n 0.00842459f $X=10.155 $Y=2.34 $X2=0
+ $Y2=0
cc_746 N_SLEEP_B_M1004_g N_VGND_c_1596_n 0.00218253f $X=9.305 $Y=1.08 $X2=0
+ $Y2=0
cc_747 N_SLEEP_B_M1032_g N_VGND_c_1596_n 0.0143572f $X=9.665 $Y=1.08 $X2=0 $Y2=0
cc_748 N_SLEEP_B_c_970_n N_VGND_c_1596_n 0.00952978f $X=10.03 $Y=1.555 $X2=0
+ $Y2=0
cc_749 N_SLEEP_B_M1023_g N_VGND_c_1596_n 0.00371696f $X=10.645 $Y=0.865 $X2=0
+ $Y2=0
cc_750 N_SLEEP_B_M1023_g N_VGND_c_1597_n 0.00180891f $X=10.645 $Y=0.865 $X2=0
+ $Y2=0
cc_751 N_SLEEP_B_M1015_g N_VGND_c_1597_n 0.0122465f $X=11.005 $Y=0.865 $X2=0
+ $Y2=0
cc_752 N_SLEEP_B_M1004_g N_VGND_c_1607_n 9.3892e-19 $X=9.305 $Y=1.08 $X2=0 $Y2=0
cc_753 N_SLEEP_B_M1032_g N_VGND_c_1607_n 7.88693e-19 $X=9.665 $Y=1.08 $X2=0
+ $Y2=0
cc_754 N_SLEEP_B_M1023_g N_VGND_c_1607_n 9.15004e-19 $X=10.645 $Y=0.865 $X2=0
+ $Y2=0
cc_755 N_SLEEP_B_M1015_g N_VGND_c_1607_n 7.68603e-19 $X=11.005 $Y=0.865 $X2=0
+ $Y2=0
cc_756 N_A_700_451#_c_1045_n N_A_2266_367#_M1008_g 0.00177536f $X=11.69 $Y=1.26
+ $X2=0 $Y2=0
cc_757 N_A_700_451#_M1027_g N_A_2266_367#_M1018_g 0.0125703f $X=11.69 $Y=2.155
+ $X2=0 $Y2=0
cc_758 N_A_700_451#_c_1045_n N_A_2266_367#_c_1223_n 0.018115f $X=11.69 $Y=1.26
+ $X2=0 $Y2=0
cc_759 N_A_700_451#_M1027_g N_A_2266_367#_c_1229_n 0.0216548f $X=11.69 $Y=2.155
+ $X2=0 $Y2=0
cc_760 N_A_700_451#_M1017_g N_A_2266_367#_c_1225_n 0.0101466f $X=11.435 $Y=0.865
+ $X2=0 $Y2=0
cc_761 N_A_700_451#_c_1045_n N_A_2266_367#_c_1225_n 0.0126396f $X=11.69 $Y=1.26
+ $X2=0 $Y2=0
cc_762 N_A_700_451#_M1027_g N_A_2266_367#_c_1227_n 0.0181785f $X=11.69 $Y=2.155
+ $X2=0 $Y2=0
cc_763 N_A_700_451#_c_1045_n N_A_2266_367#_c_1227_n 0.0104902f $X=11.69 $Y=1.26
+ $X2=0 $Y2=0
cc_764 N_A_700_451#_M1027_g N_VPWR_c_1268_n 0.0095853f $X=11.69 $Y=2.155 $X2=0
+ $Y2=0
cc_765 N_A_700_451#_M1027_g N_VPWR_c_1269_n 0.00312414f $X=11.69 $Y=2.155 $X2=0
+ $Y2=0
cc_766 N_A_700_451#_M1030_d N_VPWR_c_1264_n 0.00164553f $X=3.5 $Y=2.255 $X2=0
+ $Y2=0
cc_767 N_A_700_451#_M1009_g N_VPWR_c_1264_n 2.39862e-19 $X=7.32 $Y=2.205 $X2=0
+ $Y2=0
cc_768 N_A_700_451#_c_1046_n N_A_217_130#_c_1363_n 0.0136807f $X=3.755 $Y=2.075
+ $X2=0 $Y2=0
cc_769 N_A_700_451#_c_1065_n N_A_217_130#_c_1366_n 0.00408777f $X=3.755 $Y=0.895
+ $X2=0 $Y2=0
cc_770 N_A_700_451#_c_1046_n N_A_217_130#_c_1366_n 0.0372034f $X=3.755 $Y=2.075
+ $X2=0 $Y2=0
cc_771 N_A_700_451#_M1009_g N_KAPWR_c_1480_n 0.00373577f $X=7.32 $Y=2.205 $X2=0
+ $Y2=0
cc_772 N_A_700_451#_M1030_d N_KAPWR_c_1482_n 0.00368344f $X=3.5 $Y=2.255 $X2=0
+ $Y2=0
cc_773 N_A_700_451#_M1026_s N_KAPWR_c_1482_n 0.00365653f $X=5.58 $Y=1.575 $X2=0
+ $Y2=0
cc_774 N_A_700_451#_M1009_g N_KAPWR_c_1482_n 0.00771391f $X=7.32 $Y=2.205 $X2=0
+ $Y2=0
cc_775 N_A_700_451#_M1027_g N_KAPWR_c_1482_n 0.00480838f $X=11.69 $Y=2.155 $X2=0
+ $Y2=0
cc_776 N_A_700_451#_c_1082_n N_KAPWR_c_1482_n 0.0254614f $X=3.755 $Y=2.405 $X2=0
+ $Y2=0
cc_777 N_A_700_451#_M1022_g N_VGND_c_1595_n 0.0256038f $X=7.2 $Y=0.845 $X2=0
+ $Y2=0
cc_778 N_A_700_451#_c_1040_n N_VGND_c_1595_n 0.00836149f $X=7.275 $Y=0.21 $X2=0
+ $Y2=0
cc_779 N_A_700_451#_M1006_g N_VGND_c_1595_n 0.00160495f $X=7.71 $Y=0.845 $X2=0
+ $Y2=0
cc_780 N_A_700_451#_c_1059_n N_VGND_c_1595_n 0.00910389f $X=7.08 $Y=1.54 $X2=0
+ $Y2=0
cc_781 N_A_700_451#_c_1052_n N_VGND_c_1595_n 0.00377041f $X=7.25 $Y=1.35 $X2=0
+ $Y2=0
cc_782 N_A_700_451#_c_1039_n N_VGND_c_1596_n 0.0275976f $X=11.36 $Y=0.21 $X2=0
+ $Y2=0
cc_783 N_A_700_451#_c_1039_n N_VGND_c_1597_n 0.021354f $X=11.36 $Y=0.21 $X2=0
+ $Y2=0
cc_784 N_A_700_451#_M1017_g N_VGND_c_1597_n 0.0129762f $X=11.435 $Y=0.865 $X2=0
+ $Y2=0
cc_785 N_A_700_451#_c_1039_n N_VGND_c_1598_n 0.0111258f $X=11.36 $Y=0.21 $X2=0
+ $Y2=0
cc_786 N_A_700_451#_M1017_g N_VGND_c_1598_n 0.00113454f $X=11.435 $Y=0.865 $X2=0
+ $Y2=0
cc_787 N_A_700_451#_c_1039_n N_VGND_c_1599_n 0.0302951f $X=11.36 $Y=0.21 $X2=0
+ $Y2=0
cc_788 N_A_700_451#_c_1040_n N_VGND_c_1604_n 0.0821843f $X=7.275 $Y=0.21 $X2=0
+ $Y2=0
cc_789 N_A_700_451#_c_1039_n N_VGND_c_1605_n 0.00730371f $X=11.36 $Y=0.21 $X2=0
+ $Y2=0
cc_790 N_A_700_451#_M1021_d N_VGND_c_1607_n 0.00301588f $X=3.695 $Y=0.235 $X2=0
+ $Y2=0
cc_791 N_A_700_451#_c_1039_n N_VGND_c_1607_n 0.153232f $X=11.36 $Y=0.21 $X2=0
+ $Y2=0
cc_792 N_A_700_451#_c_1040_n N_VGND_c_1607_n 0.00752871f $X=7.275 $Y=0.21 $X2=0
+ $Y2=0
cc_793 N_A_700_451#_M1006_g N_VGND_c_1607_n 9.07789e-19 $X=7.71 $Y=0.845 $X2=0
+ $Y2=0
cc_794 N_A_700_451#_c_1047_n A_844_47# 9.92258e-19 $X=4.57 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_795 N_A_700_451#_c_1047_n A_916_47# 0.00101497f $X=4.57 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_796 N_A_700_451#_c_1058_n N_A_988_47#_c_1744_n 0.00658433f $X=5.56 $Y=1.54
+ $X2=0 $Y2=0
cc_797 N_A_700_451#_c_1051_n N_A_988_47#_c_1744_n 0.00251096f $X=5.225 $Y=1.37
+ $X2=0 $Y2=0
cc_798 N_A_700_451#_c_1059_n N_A_988_47#_c_1745_n 0.0562537f $X=7.08 $Y=1.54
+ $X2=0 $Y2=0
cc_799 N_A_700_451#_c_1061_n N_A_988_47#_c_1745_n 0.0191264f $X=5.725 $Y=1.54
+ $X2=0 $Y2=0
cc_800 N_A_700_451#_c_1052_n N_A_988_47#_c_1745_n 0.00455712f $X=7.25 $Y=1.35
+ $X2=0 $Y2=0
cc_801 N_A_700_451#_c_1047_n N_A_988_47#_c_1747_n 0.0158347f $X=4.57 $Y=0.745
+ $X2=0 $Y2=0
cc_802 N_A_700_451#_c_1048_n N_A_988_47#_c_1747_n 0.00627339f $X=4.655 $Y=1.285
+ $X2=0 $Y2=0
cc_803 N_A_700_451#_c_1049_n N_A_988_47#_c_1747_n 0.0071897f $X=5.14 $Y=1.37
+ $X2=0 $Y2=0
cc_804 N_A_700_451#_c_1051_n N_A_988_47#_c_1747_n 0.00752223f $X=5.225 $Y=1.37
+ $X2=0 $Y2=0
cc_805 N_A_700_451#_c_1058_n N_A_988_47#_c_1748_n 0.00644474f $X=5.56 $Y=1.54
+ $X2=0 $Y2=0
cc_806 N_A_700_451#_c_1061_n N_A_988_47#_c_1748_n 0.00759895f $X=5.725 $Y=1.54
+ $X2=0 $Y2=0
cc_807 N_A_2266_367#_M1018_g N_VPWR_c_1268_n 0.0203269f $X=12.455 $Y=2.465 $X2=0
+ $Y2=0
cc_808 N_A_2266_367#_c_1223_n N_VPWR_c_1268_n 0.00764098f $X=12.38 $Y=1.48 $X2=0
+ $Y2=0
cc_809 N_A_2266_367#_c_1229_n N_VPWR_c_1268_n 0.02942f $X=11.475 $Y=1.98 $X2=0
+ $Y2=0
cc_810 N_A_2266_367#_c_1226_n N_VPWR_c_1268_n 0.0276613f $X=12.17 $Y=1.48 $X2=0
+ $Y2=0
cc_811 N_A_2266_367#_M1018_g N_VPWR_c_1270_n 0.0054895f $X=12.455 $Y=2.465 $X2=0
+ $Y2=0
cc_812 N_A_2266_367#_M1018_g N_VPWR_c_1264_n 0.00744693f $X=12.455 $Y=2.465
+ $X2=0 $Y2=0
cc_813 N_A_2266_367#_M1018_g N_KAPWR_c_1482_n 0.0106059f $X=12.455 $Y=2.465
+ $X2=0 $Y2=0
cc_814 N_A_2266_367#_c_1229_n N_KAPWR_c_1482_n 0.0179983f $X=11.475 $Y=1.98
+ $X2=0 $Y2=0
cc_815 N_A_2266_367#_M1008_g N_Q_c_1576_n 0.0245583f $X=12.455 $Y=0.705 $X2=0
+ $Y2=0
cc_816 N_A_2266_367#_M1018_g N_Q_c_1576_n 0.0267812f $X=12.455 $Y=2.465 $X2=0
+ $Y2=0
cc_817 N_A_2266_367#_c_1224_n N_Q_c_1576_n 0.0120152f $X=12.455 $Y=1.48 $X2=0
+ $Y2=0
cc_818 N_A_2266_367#_c_1226_n N_Q_c_1576_n 0.0261825f $X=12.17 $Y=1.48 $X2=0
+ $Y2=0
cc_819 N_A_2266_367#_c_1225_n N_VGND_c_1597_n 0.0179429f $X=11.65 $Y=0.865 $X2=0
+ $Y2=0
cc_820 N_A_2266_367#_M1008_g N_VGND_c_1598_n 0.00782598f $X=12.455 $Y=0.705
+ $X2=0 $Y2=0
cc_821 N_A_2266_367#_c_1223_n N_VGND_c_1598_n 0.00577732f $X=12.38 $Y=1.48 $X2=0
+ $Y2=0
cc_822 N_A_2266_367#_c_1225_n N_VGND_c_1598_n 0.0309466f $X=11.65 $Y=0.865 $X2=0
+ $Y2=0
cc_823 N_A_2266_367#_c_1226_n N_VGND_c_1598_n 0.0209147f $X=12.17 $Y=1.48 $X2=0
+ $Y2=0
cc_824 N_A_2266_367#_c_1225_n N_VGND_c_1605_n 0.00658678f $X=11.65 $Y=0.865
+ $X2=0 $Y2=0
cc_825 N_A_2266_367#_M1008_g N_VGND_c_1606_n 0.00502664f $X=12.455 $Y=0.705
+ $X2=0 $Y2=0
cc_826 N_A_2266_367#_M1008_g N_VGND_c_1607_n 0.0109827f $X=12.455 $Y=0.705 $X2=0
+ $Y2=0
cc_827 N_A_2266_367#_c_1225_n N_VGND_c_1607_n 0.00983014f $X=11.65 $Y=0.865
+ $X2=0 $Y2=0
cc_828 N_VPWR_c_1264_n N_A_217_130#_M1033_s 0.00114985f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_829 N_VPWR_M1010_s N_A_217_130#_c_1372_n 0.0167135f $X=1.64 $Y=2.025 $X2=0
+ $Y2=0
cc_830 N_VPWR_c_1266_n N_A_217_130#_c_1372_n 0.00210567f $X=1.61 $Y=3.33 $X2=0
+ $Y2=0
cc_831 N_VPWR_c_1267_n N_A_217_130#_c_1372_n 0.0210468f $X=1.775 $Y=3.01 $X2=0
+ $Y2=0
cc_832 N_VPWR_c_1269_n N_A_217_130#_c_1372_n 0.011074f $X=12.005 $Y=3.33 $X2=0
+ $Y2=0
cc_833 N_VPWR_c_1265_n N_A_217_130#_c_1373_n 0.0152792f $X=0.805 $Y=2.59 $X2=0
+ $Y2=0
cc_834 N_VPWR_c_1266_n N_A_217_130#_c_1373_n 0.0092435f $X=1.61 $Y=3.33 $X2=0
+ $Y2=0
cc_835 N_VPWR_c_1267_n N_A_217_130#_c_1373_n 8.77885e-19 $X=1.775 $Y=3.01 $X2=0
+ $Y2=0
cc_836 N_VPWR_c_1264_n N_A_217_130#_c_1373_n 0.00108438f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_837 N_VPWR_c_1269_n N_A_217_130#_c_1377_n 0.0210329f $X=12.005 $Y=3.33 $X2=0
+ $Y2=0
cc_838 N_VPWR_c_1264_n N_A_217_130#_c_1377_n 0.00303861f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_839 N_VPWR_c_1264_n A_628_451# 0.00103828f $X=12.72 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_840 N_VPWR_c_1264_n A_830_419# 9.79211e-19 $X=12.72 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_841 N_VPWR_c_1264_n N_KAPWR_M1000_d 0.00117608f $X=12.72 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_842 N_VPWR_c_1269_n N_KAPWR_c_1479_n 0.0348327f $X=12.005 $Y=3.33 $X2=0 $Y2=0
cc_843 N_VPWR_c_1264_n N_KAPWR_c_1479_n 0.00479366f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_844 N_VPWR_c_1269_n N_KAPWR_c_1480_n 0.0141969f $X=12.005 $Y=3.33 $X2=0 $Y2=0
cc_845 N_VPWR_c_1264_n N_KAPWR_c_1480_n 0.00282749f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_846 N_VPWR_c_1269_n N_KAPWR_c_1481_n 0.0169477f $X=12.005 $Y=3.33 $X2=0 $Y2=0
cc_847 N_VPWR_c_1264_n N_KAPWR_c_1481_n 0.0033753f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_848 N_VPWR_M1010_s N_KAPWR_c_1482_n 0.00252192f $X=1.64 $Y=2.025 $X2=0 $Y2=0
cc_849 N_VPWR_M1027_d N_KAPWR_c_1482_n 0.00199666f $X=11.765 $Y=1.835 $X2=0
+ $Y2=0
cc_850 N_VPWR_c_1265_n N_KAPWR_c_1482_n 0.036794f $X=0.805 $Y=2.59 $X2=0 $Y2=0
cc_851 N_VPWR_c_1266_n N_KAPWR_c_1482_n 0.00229555f $X=1.61 $Y=3.33 $X2=0 $Y2=0
cc_852 N_VPWR_c_1267_n N_KAPWR_c_1482_n 0.0163658f $X=1.775 $Y=3.01 $X2=0 $Y2=0
cc_853 N_VPWR_c_1268_n N_KAPWR_c_1482_n 0.0448539f $X=12.17 $Y=1.98 $X2=0 $Y2=0
cc_854 N_VPWR_c_1269_n N_KAPWR_c_1482_n 0.0334805f $X=12.005 $Y=3.33 $X2=0 $Y2=0
cc_855 N_VPWR_c_1270_n N_KAPWR_c_1482_n 0.00138894f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_856 N_VPWR_c_1264_n N_KAPWR_c_1482_n 1.3659f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_857 N_VPWR_c_1272_n N_KAPWR_c_1482_n 0.00234064f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_858 N_VPWR_c_1269_n N_KAPWR_c_1483_n 0.030543f $X=12.005 $Y=3.33 $X2=0 $Y2=0
cc_859 N_VPWR_c_1264_n N_KAPWR_c_1483_n 0.00626082f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_860 N_VPWR_c_1264_n N_Q_M1018_d 0.00119401f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_861 N_VPWR_c_1268_n N_Q_c_1576_n 0.0516088f $X=12.17 $Y=1.98 $X2=0 $Y2=0
cc_862 N_VPWR_c_1270_n N_Q_c_1576_n 0.0210192f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_863 N_VPWR_c_1264_n N_Q_c_1576_n 0.00303861f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_864 N_A_217_130#_M1005_d N_KAPWR_c_1482_n 0.0021453f $X=1.095 $Y=2 $X2=0
+ $Y2=0
cc_865 N_A_217_130#_c_1372_n N_KAPWR_c_1482_n 0.0474253f $X=2.685 $Y=2.59 $X2=0
+ $Y2=0
cc_866 N_A_217_130#_c_1373_n N_KAPWR_c_1482_n 0.0328365f $X=1.47 $Y=2.59 $X2=0
+ $Y2=0
cc_867 N_A_217_130#_c_1375_n N_KAPWR_c_1482_n 0.0175689f $X=2.85 $Y=2.43 $X2=0
+ $Y2=0
cc_868 N_A_217_130#_c_1377_n N_KAPWR_c_1482_n 0.0243552f $X=2.85 $Y=2.59 $X2=0
+ $Y2=0
cc_869 N_A_217_130#_c_1362_n N_VGND_c_1592_n 0.00114952f $X=1.21 $Y=0.795 $X2=0
+ $Y2=0
cc_870 N_A_217_130#_c_1362_n N_VGND_c_1593_n 0.03433f $X=1.21 $Y=0.795 $X2=0
+ $Y2=0
cc_871 N_A_217_130#_c_1362_n N_VGND_c_1601_n 0.00837847f $X=1.21 $Y=0.795 $X2=0
+ $Y2=0
cc_872 N_A_217_130#_M1019_s N_VGND_c_1607_n 0.0021598f $X=2.92 $Y=0.235 $X2=0
+ $Y2=0
cc_873 N_A_217_130#_c_1362_n N_VGND_c_1607_n 0.0127401f $X=1.21 $Y=0.795 $X2=0
+ $Y2=0
cc_874 N_A_217_130#_c_1365_n A_667_47# 0.00101497f $X=3.33 $Y=0.705 $X2=-0.19
+ $Y2=-0.245
cc_875 A_628_451# N_KAPWR_c_1482_n 8.15929e-19 $X=3.14 $Y=2.255 $X2=4.315
+ $Y2=2.485
cc_876 A_830_419# N_KAPWR_c_1482_n 0.00327867f $X=4.15 $Y=2.095 $X2=4.315
+ $Y2=2.485
cc_877 N_KAPWR_c_1482_n A_1246_341# 0.00206078f $X=9.36 $Y=2.82 $X2=-0.19
+ $Y2=1.655
cc_878 N_KAPWR_c_1482_n N_Q_c_1576_n 0.039348f $X=9.36 $Y=2.82 $X2=0 $Y2=0
cc_879 N_Q_c_1576_n N_VGND_c_1598_n 0.0329963f $X=12.67 $Y=0.43 $X2=0 $Y2=0
cc_880 N_Q_c_1576_n N_VGND_c_1606_n 0.0220321f $X=12.67 $Y=0.43 $X2=0 $Y2=0
cc_881 N_Q_c_1576_n N_VGND_c_1607_n 0.0125808f $X=12.67 $Y=0.43 $X2=0 $Y2=0
cc_882 N_VGND_c_1593_n A_300_130# 0.00190018f $X=2 $Y=0.815 $X2=-0.19 $Y2=-0.245
cc_883 N_VGND_c_1607_n A_667_47# 0.00168889f $X=12.72 $Y=0 $X2=-0.19 $Y2=-0.245
cc_884 N_VGND_c_1607_n A_844_47# 0.00168889f $X=12.72 $Y=0 $X2=-0.19 $Y2=-0.245
cc_885 N_VGND_c_1607_n A_916_47# 0.00168889f $X=12.72 $Y=0 $X2=-0.19 $Y2=-0.245
cc_886 N_VGND_c_1607_n N_A_988_47#_M1016_d 0.00313365f $X=12.72 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_887 N_VGND_c_1594_n N_A_988_47#_c_1745_n 0.0177502f $X=6.02 $Y=0.78 $X2=0
+ $Y2=0
cc_888 N_VGND_c_1594_n N_A_988_47#_c_1746_n 0.0212973f $X=6.02 $Y=0.78 $X2=0
+ $Y2=0
cc_889 N_VGND_c_1595_n N_A_988_47#_c_1746_n 0.0150645f $X=6.985 $Y=0.815 $X2=0
+ $Y2=0
cc_890 N_VGND_c_1603_n N_A_988_47#_c_1746_n 0.00523206f $X=6.82 $Y=0 $X2=0 $Y2=0
cc_891 N_VGND_c_1607_n N_A_988_47#_c_1746_n 0.00763213f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_892 N_VGND_c_1594_n N_A_988_47#_c_1747_n 0.00465615f $X=6.02 $Y=0.78 $X2=0
+ $Y2=0
cc_893 N_VGND_c_1594_n N_A_988_47#_c_1748_n 0.00552422f $X=6.02 $Y=0.78 $X2=0
+ $Y2=0
