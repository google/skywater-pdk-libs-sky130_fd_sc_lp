* File: sky130_fd_sc_lp__or2_4.pxi.spice
* Created: Wed Sep  2 10:29:12 2020
* 
x_PM_SKY130_FD_SC_LP__OR2_4%B N_B_M1003_g N_B_M1011_g N_B_c_68_n N_B_c_69_n
+ N_B_c_70_n B B N_B_c_72_n PM_SKY130_FD_SC_LP__OR2_4%B
x_PM_SKY130_FD_SC_LP__OR2_4%A N_A_M1009_g N_A_M1008_g A N_A_c_100_n N_A_c_101_n
+ PM_SKY130_FD_SC_LP__OR2_4%A
x_PM_SKY130_FD_SC_LP__OR2_4%A_27_367# N_A_27_367#_M1003_d N_A_27_367#_M1011_s
+ N_A_27_367#_M1001_g N_A_27_367#_M1000_g N_A_27_367#_M1002_g
+ N_A_27_367#_M1004_g N_A_27_367#_M1005_g N_A_27_367#_M1006_g
+ N_A_27_367#_M1007_g N_A_27_367#_M1010_g N_A_27_367#_c_158_n
+ N_A_27_367#_c_159_n N_A_27_367#_c_165_n N_A_27_367#_c_167_n
+ N_A_27_367#_c_148_n N_A_27_367#_c_149_n N_A_27_367#_c_150_n
+ N_A_27_367#_c_151_n N_A_27_367#_c_215_p N_A_27_367#_c_152_n
+ N_A_27_367#_c_153_n PM_SKY130_FD_SC_LP__OR2_4%A_27_367#
x_PM_SKY130_FD_SC_LP__OR2_4%VPWR N_VPWR_M1009_d N_VPWR_M1004_d N_VPWR_M1010_d
+ N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n
+ N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n VPWR N_VPWR_c_273_n
+ N_VPWR_c_264_n N_VPWR_c_275_n PM_SKY130_FD_SC_LP__OR2_4%VPWR
x_PM_SKY130_FD_SC_LP__OR2_4%X N_X_M1001_d N_X_M1005_d N_X_M1000_s N_X_M1006_s
+ N_X_c_367_p N_X_c_353_n N_X_c_313_n N_X_c_314_n N_X_c_319_n N_X_c_320_n
+ N_X_c_368_p N_X_c_357_n N_X_c_315_n N_X_c_321_n N_X_c_316_n N_X_c_322_n X X
+ N_X_c_317_n X PM_SKY130_FD_SC_LP__OR2_4%X
x_PM_SKY130_FD_SC_LP__OR2_4%VGND N_VGND_M1003_s N_VGND_M1008_d N_VGND_M1002_s
+ N_VGND_M1007_s N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n
+ N_VGND_c_382_n VGND N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n
+ PM_SKY130_FD_SC_LP__OR2_4%VGND
cc_1 VNB N_B_c_68_n 0.0215538f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.185
cc_2 VNB N_B_c_69_n 0.0193601f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.335
cc_3 VNB N_B_c_70_n 0.00714147f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.725
cc_4 VNB B 0.0180081f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_B_c_72_n 0.0193771f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.375
cc_6 VNB N_A_M1008_g 0.0252108f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.335
cc_7 VNB N_A_c_100_n 0.0244101f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.725
cc_8 VNB N_A_c_101_n 0.00321979f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A_27_367#_M1001_g 0.0236193f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.335
cc_10 VNB N_A_27_367#_M1002_g 0.0221725f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.375
cc_11 VNB N_A_27_367#_M1005_g 0.0221584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_367#_M1007_g 0.0270724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_367#_c_148_n 0.00436375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_367#_c_149_n 0.003071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_367#_c_150_n 0.00204814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_367#_c_151_n 4.02988e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_367#_c_152_n 0.00101481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_367#_c_153_n 0.0677107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_264_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_313_n 0.0030484f $X=-0.19 $Y=-0.245 $X2=0.262 $Y2=1.375
cc_21 VNB N_X_c_314_n 0.00270083f $X=-0.19 $Y=-0.245 $X2=0.262 $Y2=1.665
cc_22 VNB N_X_c_315_n 0.00141276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_316_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_317_n 0.017778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB X 0.0244868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_373_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_VGND_c_374_n 0.0340332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_375_n 0.0043131f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.375
cc_29 VNB N_VGND_c_376_n 3.14366e-19 $X=-0.19 $Y=-0.245 $X2=0.262 $Y2=1.375
cc_30 VNB N_VGND_c_377_n 0.0284267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_378_n 0.01489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_379_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_380_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_381_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_382_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_383_n 0.0150851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_384_n 0.194919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_385_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_B_c_70_n 0.0328235f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.725
cc_40 VPB B 0.00715364f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_41 VPB N_A_M1009_g 0.0190187f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_42 VPB N_A_c_100_n 0.00619087f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.725
cc_43 VPB N_A_c_101_n 0.00354907f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_44 VPB N_A_27_367#_M1000_g 0.0200036f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_45 VPB N_A_27_367#_M1004_g 0.018348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_27_367#_M1006_g 0.0183339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_27_367#_M1010_g 0.0218662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_27_367#_c_158_n 0.00755006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_27_367#_c_159_n 0.0379885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_27_367#_c_151_n 0.00146669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_27_367#_c_153_n 0.00888213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_265_n 0.00500785f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.725
cc_53 VPB N_VPWR_c_266_n 3.20903e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_267_n 0.0408143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_268_n 0.0163082f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_269_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_270_n 0.0110534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_271_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_272_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_273_n 0.0294792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_264_n 0.0517506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_275_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_X_c_319_n 0.00305125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_X_c_320_n 0.00194123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_X_c_321_n 0.0193617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_X_c_322_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB X 0.00598057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 N_B_c_70_n N_A_M1009_g 0.0500028f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_69 N_B_c_68_n N_A_M1008_g 0.0207542f $X=0.37 $Y=1.185 $X2=0 $Y2=0
cc_70 B N_A_M1008_g 6.68712e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_B_c_72_n N_A_M1008_g 3.38491e-19 $X=0.355 $Y=1.375 $X2=0 $Y2=0
cc_72 N_B_c_70_n N_A_c_100_n 0.0500028f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_73 B N_A_c_100_n 3.3617e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B_c_72_n N_A_c_100_n 0.0119695f $X=0.355 $Y=1.375 $X2=0 $Y2=0
cc_75 N_B_c_70_n N_A_c_101_n 0.00128223f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_76 B N_A_c_101_n 0.033107f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_B_c_72_n N_A_c_101_n 0.0016557f $X=0.355 $Y=1.375 $X2=0 $Y2=0
cc_78 N_B_c_70_n N_A_27_367#_c_158_n 0.0020691f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_79 B N_A_27_367#_c_158_n 0.0271311f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B_c_70_n N_A_27_367#_c_159_n 0.0197729f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_81 N_B_c_70_n N_A_27_367#_c_165_n 0.013271f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_82 B N_A_27_367#_c_165_n 0.00101367f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_B_c_68_n N_A_27_367#_c_167_n 0.00282096f $X=0.37 $Y=1.185 $X2=0 $Y2=0
cc_84 N_B_c_68_n N_A_27_367#_c_149_n 0.00434622f $X=0.37 $Y=1.185 $X2=0 $Y2=0
cc_85 N_B_c_70_n N_VPWR_c_273_n 0.0054895f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_86 N_B_c_70_n N_VPWR_c_264_n 0.0107853f $X=0.37 $Y=1.725 $X2=0 $Y2=0
cc_87 N_B_c_68_n N_VGND_c_374_n 0.0169427f $X=0.37 $Y=1.185 $X2=0 $Y2=0
cc_88 N_B_c_69_n N_VGND_c_374_n 0.00537586f $X=0.37 $Y=1.335 $X2=0 $Y2=0
cc_89 B N_VGND_c_374_n 0.0260321f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_90 N_B_c_68_n N_VGND_c_383_n 0.00486043f $X=0.37 $Y=1.185 $X2=0 $Y2=0
cc_91 N_B_c_68_n N_VGND_c_384_n 0.00830854f $X=0.37 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A_M1008_g N_A_27_367#_M1001_g 0.0191727f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_93 N_A_M1009_g N_A_27_367#_M1000_g 0.0349889f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_c_101_n N_A_27_367#_M1000_g 2.27373e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_95 N_A_M1009_g N_A_27_367#_c_159_n 0.00313204f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A_M1009_g N_A_27_367#_c_165_n 0.0152716f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_c_100_n N_A_27_367#_c_165_n 0.00291213f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_98 N_A_c_101_n N_A_27_367#_c_165_n 0.0268001f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_99 N_A_M1008_g N_A_27_367#_c_148_n 0.01489f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_100 N_A_c_100_n N_A_27_367#_c_148_n 0.00361714f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_101 N_A_c_101_n N_A_27_367#_c_148_n 0.0140341f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_102 N_A_c_100_n N_A_27_367#_c_149_n 0.00190679f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A_c_101_n N_A_27_367#_c_149_n 0.0194709f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A_M1008_g N_A_27_367#_c_150_n 0.00349105f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_105 N_A_c_100_n N_A_27_367#_c_150_n 4.752e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_106 N_A_c_101_n N_A_27_367#_c_150_n 0.00526056f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_107 N_A_M1009_g N_A_27_367#_c_151_n 0.0035991f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_c_100_n N_A_27_367#_c_151_n 5.90868e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A_c_101_n N_A_27_367#_c_151_n 0.0132745f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_110 N_A_c_100_n N_A_27_367#_c_152_n 0.00128858f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_111 N_A_c_101_n N_A_27_367#_c_152_n 0.0146217f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_112 N_A_c_100_n N_A_27_367#_c_153_n 0.0168017f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A_c_101_n N_A_27_367#_c_153_n 2.89103e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_114 N_A_M1009_g N_VPWR_c_265_n 0.00814344f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_M1009_g N_VPWR_c_273_n 0.00585385f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_M1009_g N_VPWR_c_264_n 0.0110396f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_M1008_g N_VGND_c_374_n 6.75007e-19 $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_118 N_A_M1008_g N_VGND_c_375_n 0.00175212f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_119 N_A_M1008_g N_VGND_c_383_n 0.00585385f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_120 N_A_M1008_g N_VGND_c_384_n 0.0107334f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A_27_367#_c_165_n A_110_367# 0.00466597f $X=1.19 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_27_367#_c_165_n N_VPWR_M1009_d 0.00903334f $X=1.19 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_27_367#_c_151_n N_VPWR_M1009_d 0.00118786f $X=1.275 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_27_367#_M1000_g N_VPWR_c_265_n 0.00677703f $X=1.41 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_27_367#_c_165_n N_VPWR_c_265_n 0.0259956f $X=1.19 $Y=2.015 $X2=0
+ $Y2=0
cc_126 N_A_27_367#_M1000_g N_VPWR_c_266_n 7.49636e-19 $X=1.41 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_A_27_367#_M1004_g N_VPWR_c_266_n 0.0142954f $X=1.84 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_A_27_367#_M1006_g N_VPWR_c_266_n 0.0141372f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_27_367#_M1010_g N_VPWR_c_266_n 7.21513e-19 $X=2.7 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_27_367#_M1006_g N_VPWR_c_267_n 7.21513e-19 $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_27_367#_M1010_g N_VPWR_c_267_n 0.0150803f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_27_367#_M1000_g N_VPWR_c_268_n 0.00585385f $X=1.41 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_27_367#_M1004_g N_VPWR_c_268_n 0.00486043f $X=1.84 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_27_367#_M1006_g N_VPWR_c_271_n 0.00486043f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_27_367#_M1010_g N_VPWR_c_271_n 0.00486043f $X=2.7 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_27_367#_c_159_n N_VPWR_c_273_n 0.0210467f $X=0.26 $Y=2.95 $X2=0 $Y2=0
cc_137 N_A_27_367#_M1011_s N_VPWR_c_264_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_138 N_A_27_367#_M1000_g N_VPWR_c_264_n 0.0110861f $X=1.41 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_27_367#_M1004_g N_VPWR_c_264_n 0.00824727f $X=1.84 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_27_367#_M1006_g N_VPWR_c_264_n 0.00824727f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A_27_367#_M1010_g N_VPWR_c_264_n 0.00824727f $X=2.7 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_27_367#_c_159_n N_VPWR_c_264_n 0.0125689f $X=0.26 $Y=2.95 $X2=0 $Y2=0
cc_143 N_A_27_367#_M1002_g N_X_c_313_n 0.0141485f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_144 N_A_27_367#_M1005_g N_X_c_313_n 0.0145488f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_145 N_A_27_367#_c_215_p N_X_c_313_n 0.0469373f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_146 N_A_27_367#_c_153_n N_X_c_313_n 0.00246815f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_147 N_A_27_367#_M1001_g N_X_c_314_n 0.00139624f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_148 N_A_27_367#_c_148_n N_X_c_314_n 0.00929059f $X=1.19 $Y=1.08 $X2=0 $Y2=0
cc_149 N_A_27_367#_c_150_n N_X_c_314_n 0.00561291f $X=1.275 $Y=1.415 $X2=0 $Y2=0
cc_150 N_A_27_367#_c_215_p N_X_c_314_n 0.0153308f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_151 N_A_27_367#_c_153_n N_X_c_314_n 0.00256759f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_152 N_A_27_367#_M1004_g N_X_c_319_n 0.0135912f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_27_367#_M1006_g N_X_c_319_n 0.0137629f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_27_367#_c_215_p N_X_c_319_n 0.0471383f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_155 N_A_27_367#_c_153_n N_X_c_319_n 0.00247143f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_156 N_A_27_367#_M1000_g N_X_c_320_n 6.58764e-19 $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_27_367#_c_151_n N_X_c_320_n 0.00919426f $X=1.275 $Y=1.93 $X2=0 $Y2=0
cc_158 N_A_27_367#_c_215_p N_X_c_320_n 0.0145237f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_159 N_A_27_367#_c_153_n N_X_c_320_n 0.00256759f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_160 N_A_27_367#_M1007_g N_X_c_315_n 0.0174278f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A_27_367#_c_215_p N_X_c_315_n 0.00728094f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_162 N_A_27_367#_M1010_g N_X_c_321_n 0.0167476f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_27_367#_c_215_p N_X_c_321_n 0.00731186f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_164 N_A_27_367#_c_215_p N_X_c_316_n 0.0153308f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_165 N_A_27_367#_c_153_n N_X_c_316_n 0.00256759f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_166 N_A_27_367#_c_215_p N_X_c_322_n 0.0153308f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_167 N_A_27_367#_c_153_n N_X_c_322_n 0.00256759f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_168 N_A_27_367#_M1007_g X 0.0206605f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A_27_367#_c_215_p X 0.0143568f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_170 N_A_27_367#_c_148_n N_VGND_M1008_d 0.00243517f $X=1.19 $Y=1.08 $X2=0
+ $Y2=0
cc_171 N_A_27_367#_c_167_n N_VGND_c_374_n 0.0514364f $X=0.705 $Y=0.42 $X2=0
+ $Y2=0
cc_172 N_A_27_367#_c_149_n N_VGND_c_374_n 0.00425399f $X=0.83 $Y=1.08 $X2=0
+ $Y2=0
cc_173 N_A_27_367#_M1001_g N_VGND_c_375_n 0.00173015f $X=1.41 $Y=0.655 $X2=0
+ $Y2=0
cc_174 N_A_27_367#_c_148_n N_VGND_c_375_n 0.0192093f $X=1.19 $Y=1.08 $X2=0 $Y2=0
cc_175 N_A_27_367#_M1001_g N_VGND_c_376_n 6.4319e-19 $X=1.41 $Y=0.655 $X2=0
+ $Y2=0
cc_176 N_A_27_367#_M1002_g N_VGND_c_376_n 0.0113341f $X=1.84 $Y=0.655 $X2=0
+ $Y2=0
cc_177 N_A_27_367#_M1005_g N_VGND_c_376_n 0.0112648f $X=2.27 $Y=0.655 $X2=0
+ $Y2=0
cc_178 N_A_27_367#_M1007_g N_VGND_c_376_n 6.30983e-19 $X=2.7 $Y=0.655 $X2=0
+ $Y2=0
cc_179 N_A_27_367#_M1005_g N_VGND_c_377_n 6.30983e-19 $X=2.27 $Y=0.655 $X2=0
+ $Y2=0
cc_180 N_A_27_367#_M1007_g N_VGND_c_377_n 0.0126581f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_181 N_A_27_367#_M1001_g N_VGND_c_378_n 0.00585385f $X=1.41 $Y=0.655 $X2=0
+ $Y2=0
cc_182 N_A_27_367#_M1002_g N_VGND_c_378_n 0.00486043f $X=1.84 $Y=0.655 $X2=0
+ $Y2=0
cc_183 N_A_27_367#_M1005_g N_VGND_c_381_n 0.00486043f $X=2.27 $Y=0.655 $X2=0
+ $Y2=0
cc_184 N_A_27_367#_M1007_g N_VGND_c_381_n 0.00486043f $X=2.7 $Y=0.655 $X2=0
+ $Y2=0
cc_185 N_A_27_367#_c_167_n N_VGND_c_383_n 0.0139f $X=0.705 $Y=0.42 $X2=0 $Y2=0
cc_186 N_A_27_367#_M1003_d N_VGND_c_384_n 0.00496528f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_187 N_A_27_367#_M1001_g N_VGND_c_384_n 0.0106721f $X=1.41 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A_27_367#_M1002_g N_VGND_c_384_n 0.00824727f $X=1.84 $Y=0.655 $X2=0
+ $Y2=0
cc_189 N_A_27_367#_M1005_g N_VGND_c_384_n 0.00824727f $X=2.27 $Y=0.655 $X2=0
+ $Y2=0
cc_190 N_A_27_367#_M1007_g N_VGND_c_384_n 0.00824727f $X=2.7 $Y=0.655 $X2=0
+ $Y2=0
cc_191 N_A_27_367#_c_167_n N_VGND_c_384_n 0.00847534f $X=0.705 $Y=0.42 $X2=0
+ $Y2=0
cc_192 A_110_367# N_VPWR_c_264_n 0.00899413f $X=0.55 $Y=1.835 $X2=0 $Y2=0
cc_193 N_VPWR_c_264_n N_X_M1000_s 0.00571434f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_264_n N_X_M1006_s 0.00536646f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_268_n N_X_c_353_n 0.0120977f $X=1.89 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_264_n N_X_c_353_n 0.00691495f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_M1004_d N_X_c_319_n 0.00177068f $X=1.915 $Y=1.835 $X2=0 $Y2=0
cc_198 N_VPWR_c_266_n N_X_c_319_n 0.0172078f $X=2.055 $Y=2.2 $X2=0 $Y2=0
cc_199 N_VPWR_c_271_n N_X_c_357_n 0.0124525f $X=2.75 $Y=3.33 $X2=0 $Y2=0
cc_200 N_VPWR_c_264_n N_X_c_357_n 0.00730901f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_M1010_d N_X_c_321_n 0.00279945f $X=2.775 $Y=1.835 $X2=0 $Y2=0
cc_202 N_VPWR_c_267_n N_X_c_321_n 0.0239826f $X=2.915 $Y=2.2 $X2=0 $Y2=0
cc_203 N_X_c_313_n N_VGND_M1002_s 0.00176773f $X=2.39 $Y=1.155 $X2=0 $Y2=0
cc_204 N_X_c_315_n N_VGND_M1007_s 2.34277e-19 $X=2.855 $Y=1.155 $X2=0 $Y2=0
cc_205 N_X_c_317_n N_VGND_M1007_s 0.0020943f $X=3.065 $Y=1.245 $X2=0 $Y2=0
cc_206 N_X_c_313_n N_VGND_c_376_n 0.0171443f $X=2.39 $Y=1.155 $X2=0 $Y2=0
cc_207 N_X_c_315_n N_VGND_c_377_n 0.00363499f $X=2.855 $Y=1.155 $X2=0 $Y2=0
cc_208 N_X_c_317_n N_VGND_c_377_n 0.0203341f $X=3.065 $Y=1.245 $X2=0 $Y2=0
cc_209 N_X_c_367_p N_VGND_c_378_n 0.0124525f $X=1.625 $Y=0.42 $X2=0 $Y2=0
cc_210 N_X_c_368_p N_VGND_c_381_n 0.0124525f $X=2.485 $Y=0.42 $X2=0 $Y2=0
cc_211 N_X_M1001_d N_VGND_c_384_n 0.00536646f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_212 N_X_M1005_d N_VGND_c_384_n 0.00536646f $X=2.345 $Y=0.235 $X2=0 $Y2=0
cc_213 N_X_c_367_p N_VGND_c_384_n 0.00730901f $X=1.625 $Y=0.42 $X2=0 $Y2=0
cc_214 N_X_c_368_p N_VGND_c_384_n 0.00730901f $X=2.485 $Y=0.42 $X2=0 $Y2=0
