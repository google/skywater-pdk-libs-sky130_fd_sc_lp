* File: sky130_fd_sc_lp__nor4_1.pxi.spice
* Created: Wed Sep  2 10:10:18 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4_1%A N_A_M1002_g N_A_M1007_g A N_A_c_50_n N_A_c_51_n
+ PM_SKY130_FD_SC_LP__NOR4_1%A
x_PM_SKY130_FD_SC_LP__NOR4_1%B N_B_M1004_g N_B_M1003_g B B B B N_B_c_73_n
+ N_B_c_74_n B PM_SKY130_FD_SC_LP__NOR4_1%B
x_PM_SKY130_FD_SC_LP__NOR4_1%C N_C_M1006_g N_C_M1005_g C C C C N_C_c_116_n
+ N_C_c_117_n C PM_SKY130_FD_SC_LP__NOR4_1%C
x_PM_SKY130_FD_SC_LP__NOR4_1%D N_D_M1000_g N_D_M1001_g N_D_c_161_n D D
+ N_D_c_163_n PM_SKY130_FD_SC_LP__NOR4_1%D
x_PM_SKY130_FD_SC_LP__NOR4_1%VPWR N_VPWR_M1007_s N_VPWR_c_192_n N_VPWR_c_193_n
+ VPWR N_VPWR_c_194_n N_VPWR_c_191_n PM_SKY130_FD_SC_LP__NOR4_1%VPWR
x_PM_SKY130_FD_SC_LP__NOR4_1%Y N_Y_M1002_d N_Y_M1005_d N_Y_M1001_d N_Y_c_233_n
+ N_Y_c_225_n N_Y_c_226_n N_Y_c_240_n N_Y_c_227_n Y Y Y N_Y_c_228_n
+ PM_SKY130_FD_SC_LP__NOR4_1%Y
x_PM_SKY130_FD_SC_LP__NOR4_1%VGND N_VGND_M1002_s N_VGND_M1004_d N_VGND_M1000_d
+ N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n N_VGND_c_283_n VGND
+ N_VGND_c_284_n N_VGND_c_285_n N_VGND_c_286_n N_VGND_c_287_n N_VGND_c_288_n
+ N_VGND_c_289_n PM_SKY130_FD_SC_LP__NOR4_1%VGND
cc_1 VNB N_A_M1002_g 0.0341449f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_c_50_n 0.0306254f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.51
cc_3 VNB N_A_c_51_n 0.0153958f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.51
cc_4 VNB N_B_M1004_g 0.0262849f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_5 VNB N_B_c_73_n 0.0225277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B_c_74_n 0.00410584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_C_M1005_g 0.0262562f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_8 VNB N_C_c_116_n 0.0250741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_c_117_n 0.00274515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_D_M1000_g 0.0201996f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_11 VNB N_D_M1001_g 0.00723175f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_12 VNB N_D_c_161_n 0.0116475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB D 0.039743f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.51
cc_14 VNB N_D_c_163_n 0.052241f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.51
cc_15 VNB N_VPWR_c_191_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.665
cc_16 VNB N_Y_c_225_n 0.00978884f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.345
cc_17 VNB N_Y_c_226_n 0.00506483f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.675
cc_18 VNB N_Y_c_227_n 0.0074262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_228_n 0.00105645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_280_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_281_n 0.0384945f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.51
cc_22 VNB N_VGND_c_282_n 0.00451132f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.51
cc_23 VNB N_VGND_c_283_n 0.028337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_284_n 0.016701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_285_n 0.016701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_286_n 0.0185316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_287_n 0.184737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_288_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_289_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A_M1007_g 0.0246658f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_31 VPB N_A_c_50_n 0.00705623f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=1.51
cc_32 VPB N_A_c_51_n 0.00680852f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=1.51
cc_33 VPB N_B_M1003_g 0.0187111f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_34 VPB N_B_c_73_n 0.00625094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_B_c_74_n 0.0028192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_C_M1006_g 0.019981f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_37 VPB C 7.45203e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_38 VPB N_C_c_116_n 0.00641098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_C_c_117_n 0.00310035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_D_M1001_g 0.0258358f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_41 VPB D 0.0208843f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=1.51
cc_42 VPB N_VPWR_c_192_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_193_n 0.0484529f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_44 VPB N_VPWR_c_194_n 0.070444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_191_n 0.0615298f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.665
cc_46 VPB Y 0.00872429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB Y 0.0374549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_Y_c_228_n 0.00350675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 N_A_M1002_g N_B_M1004_g 0.0232676f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_50 N_A_M1007_g N_B_M1003_g 0.0519998f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_51 N_A_c_50_n N_B_c_73_n 0.0209994f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_52 N_A_c_51_n N_B_c_73_n 6.81522e-19 $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_53 N_A_c_50_n N_B_c_74_n 0.00711472f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_54 N_A_c_51_n N_B_c_74_n 0.0267457f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_55 N_A_M1007_g N_VPWR_c_193_n 0.0231427f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_c_50_n N_VPWR_c_193_n 0.0010888f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_57 N_A_c_51_n N_VPWR_c_193_n 0.0262906f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_58 N_A_M1007_g N_VPWR_c_194_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_M1007_g N_VPWR_c_191_n 0.00850736f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_Y_c_226_n 0.00464605f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_VGND_c_281_n 0.0178346f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_62 N_A_c_50_n N_VGND_c_281_n 0.00143487f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_63 N_A_c_51_n N_VGND_c_281_n 0.0214934f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_64 N_A_M1002_g N_VGND_c_284_n 0.00486043f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_65 N_A_M1002_g N_VGND_c_287_n 0.0082726f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_66 N_B_M1003_g N_C_M1006_g 0.0519713f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_67 B N_C_M1006_g 0.00251309f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_68 N_B_c_74_n N_C_M1006_g 0.00203836f $X=0.757 $Y=2.082 $X2=0 $Y2=0
cc_69 N_B_M1004_g N_C_M1005_g 0.0229413f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_70 N_B_M1003_g C 0.00371915f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_71 B C 0.0263643f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_72 N_B_c_74_n C 0.015402f $X=0.757 $Y=2.082 $X2=0 $Y2=0
cc_73 N_B_c_73_n N_C_c_116_n 0.0216702f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_74 N_B_c_74_n N_C_c_116_n 8.70728e-19 $X=0.757 $Y=2.082 $X2=0 $Y2=0
cc_75 N_B_c_73_n N_C_c_117_n 3.1437e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_76 N_B_c_74_n N_C_c_117_n 0.0194055f $X=0.757 $Y=2.082 $X2=0 $Y2=0
cc_77 N_B_M1003_g N_VPWR_c_193_n 0.00255019f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_78 N_B_M1003_g N_VPWR_c_194_n 0.0053453f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_79 B N_VPWR_c_194_n 0.00975276f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_80 N_B_M1003_g N_VPWR_c_191_n 0.00990261f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_81 B N_VPWR_c_191_n 0.0112198f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_82 B A_110_367# 0.00715904f $X=0.635 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_83 N_B_c_74_n A_110_367# 0.00332604f $X=0.757 $Y=2.082 $X2=-0.19 $Y2=-0.245
cc_84 N_B_c_74_n A_206_367# 7.5961e-19 $X=0.757 $Y=2.082 $X2=-0.19 $Y2=-0.245
cc_85 N_B_M1004_g N_Y_c_233_n 0.0121556f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_86 N_B_M1004_g N_Y_c_225_n 0.0121909f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_87 N_B_c_73_n N_Y_c_225_n 0.00288524f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_88 N_B_c_74_n N_Y_c_225_n 0.0164043f $X=0.757 $Y=2.082 $X2=0 $Y2=0
cc_89 N_B_M1004_g N_Y_c_226_n 0.00225587f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_90 N_B_c_73_n N_Y_c_226_n 0.0017784f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_91 N_B_c_74_n N_Y_c_226_n 0.0184894f $X=0.757 $Y=2.082 $X2=0 $Y2=0
cc_92 N_B_M1004_g N_Y_c_240_n 8.74336e-19 $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_93 N_B_M1004_g N_VGND_c_281_n 7.94728e-19 $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_94 N_B_M1004_g N_VGND_c_282_n 0.00843609f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_95 N_B_M1004_g N_VGND_c_284_n 0.0054895f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_96 N_B_M1004_g N_VGND_c_287_n 0.0105093f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_97 N_C_M1005_g N_D_M1000_g 0.0194859f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_98 N_C_M1006_g N_D_M1001_g 0.0416987f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_99 C N_D_M1001_g 0.00551876f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_100 N_C_c_116_n N_D_c_161_n 0.0194859f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_101 N_C_c_117_n N_D_c_161_n 0.00551876f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_102 N_C_M1006_g N_VPWR_c_194_n 0.00443252f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_103 C N_VPWR_c_194_n 0.0109912f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_104 N_C_M1006_g N_VPWR_c_191_n 0.0075139f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_105 C N_VPWR_c_191_n 0.0121098f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_106 C A_304_367# 0.0152615f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_107 N_C_M1005_g N_Y_c_233_n 8.72471e-19 $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_108 N_C_M1005_g N_Y_c_225_n 0.0121909f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_109 N_C_c_116_n N_Y_c_225_n 0.00485559f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_110 N_C_c_117_n N_Y_c_225_n 0.0338914f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_111 N_C_M1005_g N_Y_c_240_n 0.0122491f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_112 N_C_M1005_g N_Y_c_227_n 0.00267203f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_113 C Y 0.0583222f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_114 N_C_M1006_g Y 9.00209e-19 $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_115 N_C_M1006_g N_Y_c_228_n 0.00106206f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_116 N_C_M1005_g N_Y_c_228_n 0.00116544f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_117 N_C_c_116_n N_Y_c_228_n 2.40175e-19 $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_118 N_C_c_117_n N_Y_c_228_n 0.0583222f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_119 N_C_M1005_g N_VGND_c_282_n 0.00843609f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_120 N_C_M1005_g N_VGND_c_283_n 7.29111e-19 $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_121 N_C_M1005_g N_VGND_c_285_n 0.0054895f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_122 N_C_M1005_g N_VGND_c_287_n 0.0105093f $X=1.555 $Y=0.655 $X2=0 $Y2=0
cc_123 N_D_M1001_g N_VPWR_c_194_n 0.00404729f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_124 N_D_M1001_g N_VPWR_c_191_n 0.00808772f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_125 N_D_M1000_g N_Y_c_227_n 0.0115758f $X=1.985 $Y=0.655 $X2=0 $Y2=0
cc_126 N_D_c_161_n N_Y_c_227_n 0.00237158f $X=1.985 $Y=1.375 $X2=0 $Y2=0
cc_127 D N_Y_c_227_n 0.014492f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_128 N_D_c_163_n N_Y_c_227_n 0.00145441f $X=2.365 $Y=1.375 $X2=0 $Y2=0
cc_129 N_D_M1001_g Y 0.00350209f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_130 D Y 0.00771178f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_131 N_D_c_163_n Y 0.00628324f $X=2.365 $Y=1.375 $X2=0 $Y2=0
cc_132 N_D_M1001_g Y 0.0213444f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_133 N_D_M1001_g N_Y_c_228_n 0.0108142f $X=1.985 $Y=2.465 $X2=0 $Y2=0
cc_134 N_D_c_161_n N_Y_c_228_n 0.00691476f $X=1.985 $Y=1.375 $X2=0 $Y2=0
cc_135 D N_Y_c_228_n 0.0401797f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_136 N_D_c_163_n N_Y_c_228_n 0.00688609f $X=2.365 $Y=1.375 $X2=0 $Y2=0
cc_137 D N_VGND_M1000_d 5.6606e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_138 N_D_M1000_g N_VGND_c_283_n 0.0123942f $X=1.985 $Y=0.655 $X2=0 $Y2=0
cc_139 D N_VGND_c_283_n 0.00763351f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_140 N_D_c_163_n N_VGND_c_283_n 0.00682786f $X=2.365 $Y=1.375 $X2=0 $Y2=0
cc_141 N_D_M1000_g N_VGND_c_285_n 0.00486043f $X=1.985 $Y=0.655 $X2=0 $Y2=0
cc_142 N_D_M1000_g N_VGND_c_287_n 0.0082726f $X=1.985 $Y=0.655 $X2=0 $Y2=0
cc_143 N_VPWR_c_191_n A_110_367# 0.0045059f $X=2.64 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_144 N_VPWR_c_191_n A_206_367# 0.0145619f $X=2.64 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_145 N_VPWR_c_191_n A_304_367# 0.00827225f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_146 N_VPWR_c_191_n N_Y_M1001_d 0.00215158f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_147 N_VPWR_c_194_n Y 0.027523f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_148 N_VPWR_c_191_n Y 0.015817f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_149 N_Y_c_225_n N_VGND_M1004_d 0.00576947f $X=1.605 $Y=1.15 $X2=0 $Y2=0
cc_150 N_Y_c_226_n N_VGND_c_281_n 0.00201679f $X=0.855 $Y=1.15 $X2=0 $Y2=0
cc_151 N_Y_c_233_n N_VGND_c_282_n 0.0415005f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_152 N_Y_c_225_n N_VGND_c_282_n 0.0266856f $X=1.605 $Y=1.15 $X2=0 $Y2=0
cc_153 N_Y_c_240_n N_VGND_c_282_n 0.0415005f $X=1.77 $Y=0.42 $X2=0 $Y2=0
cc_154 N_Y_c_227_n N_VGND_c_283_n 0.00178608f $X=2.025 $Y=1.15 $X2=0 $Y2=0
cc_155 N_Y_c_233_n N_VGND_c_284_n 0.015688f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_156 N_Y_c_240_n N_VGND_c_285_n 0.015688f $X=1.77 $Y=0.42 $X2=0 $Y2=0
cc_157 N_Y_M1002_d N_VGND_c_287_n 0.00380103f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_158 N_Y_M1005_d N_VGND_c_287_n 0.00380103f $X=1.63 $Y=0.235 $X2=0 $Y2=0
cc_159 N_Y_c_233_n N_VGND_c_287_n 0.00984745f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_160 N_Y_c_240_n N_VGND_c_287_n 0.00984745f $X=1.77 $Y=0.42 $X2=0 $Y2=0
