* NGSPICE file created from sky130_fd_sc_lp__and4b_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4b_m A_N B C D VGND VNB VPB VPWR X
M1000 X a_240_73# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=4.179e+11p ps=4.51e+06u
M1001 VPWR B a_240_73# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.499e+11p ps=2.87e+06u
M1002 a_323_73# a_27_55# a_240_73# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1003 a_395_73# B a_323_73# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_467_73# C a_395_73# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1005 a_240_73# C VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR D a_240_73# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_27_55# VNB nshort w=420000u l=150000u
+  ad=2.751e+11p pd=2.99e+06u as=1.113e+11p ps=1.37e+06u
M1008 VPWR A_N a_27_55# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 VGND D a_467_73# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_240_73# a_27_55# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_240_73# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

