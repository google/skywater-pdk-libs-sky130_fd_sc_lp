* File: sky130_fd_sc_lp__a22o_lp.pex.spice
* Created: Wed Sep  2 09:22:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22O_LP%A1 3 7 9 10 12 16 18 19 23
c61 16 0 1.92583e-19 $X=1.96 $Y=1.02
c62 12 0 1.07725e-19 $X=1.96 $Y=0.94
r63 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.42
+ $Y=1.285 $X2=0.42 $Y2=1.285
r64 18 19 11.9735 $w=3.77e-07 $l=3.7e-07 $layer=LI1_cond $X=0.355 $Y=1.295
+ $X2=0.355 $Y2=1.665
r65 18 24 0.323607 $w=3.77e-07 $l=1e-08 $layer=LI1_cond $X=0.355 $Y=1.295
+ $X2=0.355 $Y2=1.285
r66 16 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.02
+ $X2=1.96 $Y2=0.855
r67 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.02 $X2=1.96 $Y2=1.02
r68 12 15 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.96 $Y=0.94 $X2=1.96
+ $Y2=1.02
r69 11 24 11.1645 $w=3.77e-07 $l=4.45393e-07 $layer=LI1_cond $X=0.585 $Y=0.94
+ $X2=0.355 $Y2=1.285
r70 10 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0.94
+ $X2=1.96 $Y2=0.94
r71 10 11 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=1.795 $Y=0.94
+ $X2=0.585 $Y2=0.94
r72 9 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.42 $Y=1.625
+ $X2=0.42 $Y2=1.285
r73 7 27 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.87 $Y=0.445
+ $X2=1.87 $Y2=0.855
r74 1 9 47.383 $w=2.95e-07 $l=3.53129e-07 $layer=POLY_cond $X=0.56 $Y=1.915
+ $X2=0.42 $Y2=1.625
r75 1 3 156.526 $w=2.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.56 $Y=1.915 $X2=0.56
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%B2 3 7 11 12 13 16
r45 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.06
+ $Y=1.37 $X2=1.06 $Y2=1.37
r46 13 17 2.49927 $w=6.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.54 $X2=1.06
+ $Y2=1.54
r47 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.06 $Y=1.71
+ $X2=1.06 $Y2=1.37
r48 11 12 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.71
+ $X2=1.06 $Y2=1.875
r49 10 16 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.205
+ $X2=1.06 $Y2=1.37
r50 7 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.05 $Y=0.445
+ $X2=1.05 $Y2=1.205
r51 3 12 166.464 $w=2.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.09 $Y=2.545
+ $X2=1.09 $Y2=1.875
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%B1 3 5 8 10 11 12 13 18
c51 11 0 1.07725e-19 $X=1.475 $Y=0.88
c52 10 0 2.10144e-20 $X=1.475 $Y=0.73
r53 18 20 24.7179 $w=2.73e-07 $l=1.4e-07 $layer=POLY_cond $X=1.785 $Y=1.677
+ $X2=1.925 $Y2=1.677
r54 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.785
+ $Y=1.615 $X2=1.785 $Y2=1.615
r55 13 19 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=1.785 $Y2=1.615
r56 12 19 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=1.785 $Y2=1.615
r57 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.475 $Y=0.73
+ $X2=1.475 $Y2=0.88
r58 6 20 4.92893 $w=2.5e-07 $l=2.28e-07 $layer=POLY_cond $X=1.925 $Y=1.905
+ $X2=1.925 $Y2=1.677
r59 6 8 159.01 $w=2.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.925 $Y=1.905
+ $X2=1.925 $Y2=2.545
r60 5 18 48.5531 $w=2.73e-07 $l=3.71551e-07 $layer=POLY_cond $X=1.51 $Y=1.45
+ $X2=1.785 $Y2=1.677
r61 5 11 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.51 $Y=1.45 $X2=1.51
+ $Y2=0.88
r62 3 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.44 $Y=0.445 $X2=1.44
+ $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%A2 1 3 6 9 10 11 15
c47 10 0 1.92583e-19 $X=2.64 $Y=1.295
r48 15 17 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.29
+ $X2=2.575 $Y2=1.125
r49 10 11 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.62 $Y=1.29
+ $X2=2.62 $Y2=1.665
r50 10 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.62
+ $Y=1.29 $X2=2.62 $Y2=1.29
r51 8 15 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=2.575 $Y=1.335
+ $X2=2.575 $Y2=1.29
r52 8 9 33.1044 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=2.575 $Y=1.335
+ $X2=2.575 $Y2=1.585
r53 6 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.44 $Y=0.445
+ $X2=2.44 $Y2=1.125
r54 1 9 45.3567 $w=3.56e-07 $l=3.90416e-07 $layer=POLY_cond $X=2.455 $Y=1.92
+ $X2=2.575 $Y2=1.585
r55 1 3 120.5 $w=2.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.455 $Y=1.92 $X2=2.455
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%A_243_409# 1 2 7 9 12 16 19 21 24 26 28 29
+ 30 32 33 35 37 41 47 48
c102 26 0 2.10144e-20 $X=2.305 $Y=0.59
r103 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.21
+ $Y=0.94 $X2=3.21 $Y2=0.94
r104 41 43 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.39 $Y=0.59
+ $X2=2.39 $Y2=0.86
r105 37 39 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.655 $Y=0.445
+ $X2=1.655 $Y2=0.59
r106 35 48 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.05 $Y=1.975
+ $X2=3.05 $Y2=1.445
r107 33 48 9.81506 $w=4.08e-07 $l=2.05e-07 $layer=LI1_cond $X=3.17 $Y=1.24
+ $X2=3.17 $Y2=1.445
r108 32 46 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=0.945
+ $X2=3.17 $Y2=0.86
r109 32 33 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.17 $Y=0.945
+ $X2=3.17 $Y2=1.24
r110 31 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.86
+ $X2=2.39 $Y2=0.86
r111 30 46 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.965 $Y=0.86
+ $X2=3.17 $Y2=0.86
r112 30 31 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.965 $Y=0.86
+ $X2=2.475 $Y2=0.86
r113 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.965 $Y=2.06
+ $X2=3.05 $Y2=1.975
r114 28 29 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.965 $Y=2.06
+ $X2=1.825 $Y2=2.06
r115 27 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=0.59
+ $X2=1.655 $Y2=0.59
r116 26 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0.59
+ $X2=2.39 $Y2=0.59
r117 26 27 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.305 $Y=0.59
+ $X2=1.82 $Y2=0.59
r118 22 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.66 $Y=2.145
+ $X2=1.825 $Y2=2.06
r119 22 24 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.66 $Y=2.145
+ $X2=1.66 $Y2=2.19
r120 20 47 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=3.232 $Y=1.258
+ $X2=3.232 $Y2=0.94
r121 20 21 31.3347 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=3.232 $Y=1.258
+ $X2=3.232 $Y2=1.445
r122 19 47 8.15692 $w=3.75e-07 $l=5.5e-08 $layer=POLY_cond $X=3.232 $Y=0.885
+ $X2=3.232 $Y2=0.94
r123 12 21 273.299 $w=2.5e-07 $l=1.1e-06 $layer=POLY_cond $X=3.215 $Y=2.545
+ $X2=3.215 $Y2=1.445
r124 7 19 24.6308 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=3.15 $Y=0.735
+ $X2=3.15 $Y2=0.885
r125 7 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.345 $Y=0.735
+ $X2=3.345 $Y2=0.445
r126 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.955 $Y=0.735
+ $X2=2.955 $Y2=0.445
r127 2 24 300 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=2 $X=1.215
+ $Y=2.045 $X2=1.66 $Y2=2.19
r128 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.235 $X2=1.655 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%VPWR 1 2 7 9 15 17 19 29 30 36
r38 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=3.33
+ $X2=2.72 $Y2=3.33
r43 27 29 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.885 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 20 33 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r50 20 22 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.72 $Y2=3.33
r52 19 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 17 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 17 23 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=3.245
+ $X2=2.72 $Y2=3.33
r56 13 15 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=2.72 $Y=3.245
+ $X2=2.72 $Y2=2.49
r57 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.295 $Y=2.19
+ $X2=0.295 $Y2=2.9
r58 7 33 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r59 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.9
r60 2 15 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=2.045 $X2=2.72 $Y2=2.49
r61 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.9
r62 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%A_137_409# 1 2 7 9 11 15
r28 13 15 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.19 $Y=2.895
+ $X2=2.19 $Y2=2.49
r29 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=2.98
+ $X2=0.825 $Y2=2.98
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.025 $Y=2.98
+ $X2=2.19 $Y2=2.895
r31 11 12 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.025 $Y=2.98
+ $X2=0.99 $Y2=2.98
r32 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=2.895
+ $X2=0.825 $Y2=2.98
r33 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.825 $Y=2.895
+ $X2=0.825 $Y2=2.22
r34 2 15 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=2.045 $X2=2.19 $Y2=2.49
r35 1 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.825 $Y2=2.9
r36 1 9 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.045 $X2=0.825 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%X 1 2 8 10 13 14 15 19
r24 19 30 1.4685 $w=4.1e-07 $l=4e-08 $layer=LI1_cond $X=3.52 $Y=2.23 $X2=3.52
+ $Y2=2.19
r25 15 25 3.51355 $w=4.08e-07 $l=1.25e-07 $layer=LI1_cond $X=3.52 $Y=2.775
+ $X2=3.52 $Y2=2.9
r26 14 15 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.52 $Y=2.405
+ $X2=3.52 $Y2=2.775
r27 14 19 4.91896 $w=4.08e-07 $l=1.75e-07 $layer=LI1_cond $X=3.52 $Y=2.405
+ $X2=3.52 $Y2=2.23
r28 13 30 5.37216 $w=3.52e-07 $l=1.55e-07 $layer=LI1_cond $X=3.52 $Y=2.035
+ $X2=3.52 $Y2=2.19
r29 10 12 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=0.43
+ $X2=3.56 $Y2=0.595
r30 8 13 7.25742 $w=3.52e-07 $l=1.67929e-07 $layer=LI1_cond $X=3.64 $Y=1.92
+ $X2=3.52 $Y2=2.035
r31 8 12 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.64 $Y=1.92
+ $X2=3.64 $Y2=0.595
r32 2 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.045 $X2=3.48 $Y2=2.19
r33 2 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.045 $X2=3.48 $Y2=2.9
r34 1 10 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.235 $X2=3.56 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_LP%VGND 1 2 11 15 18 19 20 30 31 34
r46 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r48 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r49 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r52 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.835
+ $Y2=0
r54 22 24 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.2 $Y2=0
r55 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r56 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r57 18 27 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.64
+ $Y2=0
r58 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.78
+ $Y2=0
r59 17 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.6
+ $Y2=0
r60 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.78
+ $Y2=0
r61 13 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r62 13 15 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.405
r63 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.085
+ $X2=0.835 $Y2=0
r64 9 11 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.835 $Y=0.085
+ $X2=0.835 $Y2=0.445
r65 2 15 182 $w=1.7e-07 $l=2.98119e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.235 $X2=2.74 $Y2=0.405
r66 1 11 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.235 $X2=0.835 $Y2=0.445
.ends

