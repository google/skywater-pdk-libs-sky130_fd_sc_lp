* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_260_341# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_481# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VPWR a_218_131# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND B1 a_146_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_218_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_146_131# B2 a_218_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_218_131# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 X a_218_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR B2 a_27_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_218_131# a_260_341# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND A2_N a_260_341# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_27_481# a_260_341# a_218_131# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_260_341# A2_N a_480_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_480_367# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
