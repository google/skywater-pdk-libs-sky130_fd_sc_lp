* File: sky130_fd_sc_lp__mux2_lp2.pex.spice
* Created: Fri Aug 28 10:44:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%A_84_259# 1 2 7 9 13 17 19 25 27 29 30 32
+ 34 36 37
r87 36 37 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.66 $Y=0.535
+ $X2=2.495 $Y2=0.535
r88 30 32 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.59 $Y=2.15
+ $X2=2.16 $Y2=2.15
r89 29 37 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.59 $Y=0.43
+ $X2=2.495 $Y2=0.43
r90 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=2.065
+ $X2=1.59 $Y2=2.15
r91 26 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.235
+ $X2=1.505 $Y2=1.07
r92 26 27 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.505 $Y=1.235
+ $X2=1.505 $Y2=2.065
r93 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=0.905
+ $X2=1.505 $Y2=1.07
r94 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=0.515
+ $X2=1.59 $Y2=0.43
r95 24 25 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.505 $Y=0.515
+ $X2=1.505 $Y2=0.905
r96 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.795
+ $Y=1.07 $X2=0.795 $Y2=1.07
r97 19 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=1.07
+ $X2=1.505 $Y2=1.07
r98 19 21 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=1.42 $Y=1.07
+ $X2=0.795 $Y2=1.07
r99 15 22 41.6532 $w=1.93e-07 $l=2.38642e-07 $layer=POLY_cond $X=0.86 $Y=0.905
+ $X2=0.69 $Y2=1.07
r100 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.86 $Y=0.905
+ $X2=0.86 $Y2=0.495
r101 11 22 41.6532 $w=1.93e-07 $l=2.59711e-07 $layer=POLY_cond $X=0.5 $Y=0.905
+ $X2=0.69 $Y2=1.07
r102 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.5 $Y=0.905
+ $X2=0.5 $Y2=0.495
r103 7 22 49.619 $w=3.87e-07 $l=4.16233e-07 $layer=POLY_cond $X=0.545 $Y=1.42
+ $X2=0.69 $Y2=1.07
r104 7 9 269.572 $w=2.5e-07 $l=1.085e-06 $layer=POLY_cond $X=0.545 $Y=1.42
+ $X2=0.545 $Y2=2.505
r105 2 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.02
+ $Y=2.005 $X2=2.16 $Y2=2.15
r106 1 36 182 $w=1.7e-07 $l=6.21188e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.285 $X2=2.66 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%A_182_303# 1 2 9 12 13 15 16 17 20 24 27 28
+ 29 30 33 35 38 41 43
r105 43 45 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.38 $Y=0.495
+ $X2=4.38 $Y2=0.725
r106 38 45 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=4.46 $Y=1.985
+ $X2=4.46 $Y2=0.725
r107 36 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=2.07
+ $X2=3.75 $Y2=2.07
r108 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.375 $Y=2.07
+ $X2=4.46 $Y2=1.985
r109 35 36 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.375 $Y=2.07
+ $X2=3.915 $Y2=2.07
r110 31 41 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=2.585
+ $X2=3.75 $Y2=2.5
r111 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.75 $Y=2.585
+ $X2=3.75 $Y2=2.86
r112 30 41 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=2.415
+ $X2=3.75 $Y2=2.5
r113 29 40 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=2.155
+ $X2=3.75 $Y2=2.07
r114 29 30 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=3.75 $Y=2.155
+ $X2=3.75 $Y2=2.415
r115 27 41 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=2.5
+ $X2=3.75 $Y2=2.5
r116 27 28 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=3.585 $Y=2.5
+ $X2=1.24 $Y2=2.5
r117 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.68 $X2=1.075 $Y2=1.68
r118 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.075 $Y=2.415
+ $X2=1.24 $Y2=2.5
r119 22 24 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=1.075 $Y=2.415
+ $X2=1.075 $Y2=1.68
r120 18 20 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.455 $Y=0.855
+ $X2=1.67 $Y2=0.855
r121 16 25 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.28 $Y=1.68
+ $X2=1.075 $Y2=1.68
r122 16 17 1.50692 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.28 $Y=1.68
+ $X2=1.405 $Y2=1.68
r123 13 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.67 $Y=0.78
+ $X2=1.67 $Y2=0.855
r124 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.67 $Y=0.78
+ $X2=1.67 $Y2=0.495
r125 12 17 30.2679 $w=2e-07 $l=1.88348e-07 $layer=POLY_cond $X=1.455 $Y=1.515
+ $X2=1.405 $Y2=1.68
r126 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.455 $Y=0.93
+ $X2=1.455 $Y2=0.855
r127 11 12 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=1.455 $Y=0.93
+ $X2=1.455 $Y2=1.515
r128 7 17 30.2679 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.845
+ $X2=1.405 $Y2=1.68
r129 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.405 $Y=1.845
+ $X2=1.405 $Y2=2.505
r130 2 40 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=2.005 $X2=3.75 $Y2=2.15
r131 2 33 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=2.005 $X2=3.75 $Y2=2.86
r132 1 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.24
+ $Y=0.285 $X2=4.38 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%A1 3 7 9 12 15 16 17 20 21 22 32
c67 20 0 1.80374e-19 $X=2.895 $Y=1.07
r68 22 32 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.07
+ $X2=3.12 $Y2=0.905
r69 22 32 1.65351 $w=2.28e-07 $l=3.3e-08 $layer=LI1_cond $X=3.12 $Y=0.872
+ $X2=3.12 $Y2=0.905
r70 21 22 15.8837 $w=2.28e-07 $l=3.17e-07 $layer=LI1_cond $X=3.12 $Y=0.555
+ $X2=3.12 $Y2=0.872
r71 20 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.895 $Y=1.07
+ $X2=2.895 $Y2=0.905
r72 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.895
+ $Y=1.07 $X2=2.895 $Y2=1.07
r73 17 19 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.665 $Y=1.07
+ $X2=2.895 $Y2=1.07
r74 16 22 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=1.07
+ $X2=3.12 $Y2=1.07
r75 16 19 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.005 $Y=1.07
+ $X2=2.895 $Y2=1.07
r76 14 17 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.58 $Y=1.235
+ $X2=2.665 $Y2=1.07
r77 14 15 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.58 $Y=1.235
+ $X2=2.58 $Y2=1.515
r78 12 28 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.68
+ $X2=1.935 $Y2=1.845
r79 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.68 $X2=1.935 $Y2=1.68
r80 9 15 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.495 $Y=1.68
+ $X2=2.58 $Y2=1.515
r81 9 11 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.495 $Y=1.68
+ $X2=1.935 $Y2=1.68
r82 7 30 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.875 $Y=0.495
+ $X2=2.875 $Y2=0.905
r83 3 28 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.895 $Y=2.505
+ $X2=1.895 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%A0 1 3 6 8 10 11 15
c45 11 0 1.80374e-19 $X=2.16 $Y=0.925
r46 13 15 16.2472 $w=2.67e-07 $l=9e-08 $layer=POLY_cond $X=2.06 $Y=0.98 $X2=2.15
+ $Y2=0.98
r47 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=0.98 $X2=2.15 $Y2=0.98
r48 6 10 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.465 $Y=1.6
+ $X2=2.465 $Y2=1.475
r49 6 8 224.851 $w=2.5e-07 $l=9.05e-07 $layer=POLY_cond $X=2.465 $Y=1.6
+ $X2=2.465 $Y2=2.505
r50 4 15 47.839 $w=2.67e-07 $l=3.37565e-07 $layer=POLY_cond $X=2.415 $Y=1.145
+ $X2=2.15 $Y2=0.98
r51 4 10 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.415 $Y=1.145
+ $X2=2.415 $Y2=1.475
r52 1 13 16.2448 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=0.815
+ $X2=2.06 $Y2=0.98
r53 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.06 $Y=0.815 $X2=2.06
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%S 3 7 11 15 19 21 22 23 38
r60 36 38 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.03 $Y=1.64
+ $X2=4.165 $Y2=1.64
r61 34 36 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.805 $Y=1.64
+ $X2=4.03 $Y2=1.64
r62 33 34 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=3.485 $Y=1.64
+ $X2=3.805 $Y2=1.64
r63 32 33 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.375 $Y=1.64
+ $X2=3.485 $Y2=1.64
r64 30 32 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=3.01 $Y=1.64
+ $X2=3.375 $Y2=1.64
r65 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.01
+ $Y=1.64 $X2=3.01 $Y2=1.64
r66 27 30 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.955 $Y=1.64
+ $X2=3.01 $Y2=1.64
r67 23 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.03
+ $Y=1.64 $X2=4.03 $Y2=1.64
r68 22 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.64 $X2=4.03
+ $Y2=1.64
r69 21 22 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.64 $X2=3.6
+ $Y2=1.64
r70 21 31 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.12 $Y=1.64
+ $X2=3.01 $Y2=1.64
r71 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.165 $Y=1.475
+ $X2=4.165 $Y2=1.64
r72 17 19 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.165 $Y=1.475
+ $X2=4.165 $Y2=0.495
r73 13 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.475
+ $X2=3.805 $Y2=1.64
r74 13 15 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.805 $Y=1.475
+ $X2=3.805 $Y2=0.495
r75 9 33 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.805
+ $X2=3.485 $Y2=1.64
r76 9 11 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.485 $Y=1.805
+ $X2=3.485 $Y2=2.505
r77 5 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.475
+ $X2=3.375 $Y2=1.64
r78 5 7 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.375 $Y=1.475
+ $X2=3.375 $Y2=0.495
r79 1 27 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.805
+ $X2=2.955 $Y2=1.64
r80 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.955 $Y=1.805 $X2=2.955
+ $Y2=2.505
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%X 1 2 9 11 12 13 14 15 16 41
r21 24 41 1.78887 $w=3.33e-07 $l=5.2e-08 $layer=LI1_cond $X=0.282 $Y=2.353
+ $X2=0.282 $Y2=2.405
r22 16 43 3.40573 $w=3.33e-07 $l=9.9e-08 $layer=LI1_cond $X=0.282 $Y=2.421
+ $X2=0.282 $Y2=2.52
r23 16 41 0.550421 $w=3.33e-07 $l=1.6e-08 $layer=LI1_cond $X=0.282 $Y=2.421
+ $X2=0.282 $Y2=2.405
r24 16 24 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=0.282 $Y=2.336
+ $X2=0.282 $Y2=2.353
r25 16 38 6.39864 $w=3.33e-07 $l=1.86e-07 $layer=LI1_cond $X=0.282 $Y=2.336
+ $X2=0.282 $Y2=2.15
r26 15 38 3.95615 $w=3.33e-07 $l=1.15e-07 $layer=LI1_cond $X=0.282 $Y=2.035
+ $X2=0.282 $Y2=2.15
r27 14 15 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=2.035
r28 13 14 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=1.295
+ $X2=0.282 $Y2=1.665
r29 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.282 $Y=0.925
+ $X2=0.282 $Y2=1.295
r30 11 12 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=0.282 $Y=0.495
+ $X2=0.282 $Y2=0.925
r31 9 43 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.28 $Y=2.86 $X2=0.28
+ $Y2=2.52
r32 2 38 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.005 $X2=0.28 $Y2=2.15
r33 2 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.005 $X2=0.28 $Y2=2.86
r34 1 11 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.285 $X2=0.285 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%VPWR 1 2 11 15 17 19 29 30 33 36
r41 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r44 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r45 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r47 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r48 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.22 $Y2=3.33
r49 24 26 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.6 $Y2=3.33
r50 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r53 20 22 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=3.22 $Y2=3.33
r55 19 22 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 17 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 17 23 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=3.245
+ $X2=3.22 $Y2=3.33
r59 13 15 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.22 $Y=3.245
+ $X2=3.22 $Y2=2.855
r60 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245 $X2=0.81
+ $Y2=3.33
r61 9 11 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.855
r62 2 15 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=2.005 $X2=3.22 $Y2=2.855
r63 1 11 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.005 $X2=0.81 $Y2=2.855
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP2%VGND 1 2 9 13 15 17 22 29 30 33 36
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r54 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r56 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r57 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.59
+ $Y2=0
r58 27 29 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=4.56
+ $Y2=0
r59 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r60 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.075
+ $Y2=0
r62 23 25 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=1.24 $Y=0 $X2=3.12
+ $Y2=0
r63 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.59
+ $Y2=0
r64 22 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.12
+ $Y2=0
r65 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r66 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.075
+ $Y2=0
r68 17 19 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.72
+ $Y2=0
r69 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r70 15 34 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r71 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=0.085
+ $X2=3.59 $Y2=0
r72 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.59 $Y=0.085
+ $X2=3.59 $Y2=0.495
r73 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.075 $Y=0.085
+ $X2=1.075 $Y2=0
r74 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.075 $Y=0.085
+ $X2=1.075 $Y2=0.495
r75 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.285 $X2=3.59 $Y2=0.495
r76 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.285 $X2=1.075 $Y2=0.495
.ends

