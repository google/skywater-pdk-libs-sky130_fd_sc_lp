* File: sky130_fd_sc_lp__o21bai_1.spice
* Created: Wed Sep  2 10:17:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21bai_1.pex.spice"
.subckt sky130_fd_sc_lp__o21bai_1  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B1_N_M1005_g N_A_27_69#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_310_47#_M1006_d N_A_27_69#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1197 AS=0.2352 PD=1.125 PS=2.24 NRD=0.708 NRS=2.136 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_310_47#_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1449 AS=0.1197 PD=1.185 PS=1.125 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1004 N_A_310_47#_M1004_d N_A1_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1449 PD=2.21 PS=1.185 NRD=0 NRS=6.42 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_B1_N_M1000_g N_A_27_69#_M1000_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=46.886 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_27_69#_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.285075 PD=1.68 PS=2.4525 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 A_424_367# N_A2_M1007_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.2646 PD=1.47 PS=1.68 NRD=7.8012 NRS=10.9335 M=1 R=8.4 SA=75000.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_424_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__o21bai_1.pxi.spice"
*
.ends
*
*
