* File: sky130_fd_sc_lp__o32ai_1.spice
* Created: Fri Aug 28 11:18:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o32ai_1  VNB VPB B1 B2 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_Y_M1009_d N_B1_M1009_g N_A_76_69#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1386 AS=0.2226 PD=1.17 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_76_69#_M1001_d N_B2_M1001_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.1386 PD=1.14 PS=1.17 NRD=2.856 NRS=7.14 M=1 R=5.6 SA=75000.7
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A3_M1003_g N_A_76_69#_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.126 PD=1.46 PS=1.14 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75001.4
+ A=0.126 P=1.98 MULT=1
MM1007 N_A_76_69#_M1007_d N_A2_M1007_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A1_M1002_g N_A_76_69#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 A_159_367# N_B1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g A_159_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.4347
+ AS=0.1323 PD=1.95 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6 SB=75001.9
+ A=0.189 P=2.82 MULT=1
MM1006 A_399_367# N_A3_M1006_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.4347 PD=1.56 PS=1.95 NRD=14.8341 NRS=0 M=1 R=8.4 SA=75001.4 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1008 A_489_367# N_A2_M1008_g A_399_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.189 PD=1.56 PS=1.56 NRD=14.8341 NRS=14.8341 M=1 R=8.4 SA=75001.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_489_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.189 PD=3.05 PS=1.56 NRD=0 NRS=14.8341 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o32ai_1.pxi.spice"
*
.ends
*
*
