* File: sky130_fd_sc_lp__srsdfrtn_1.pxi.spice
* Created: Wed Sep  2 10:39:07 2020
* 
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%SCE N_SCE_M1001_g N_SCE_M1016_g N_SCE_c_363_n
+ N_SCE_c_364_n N_SCE_M1025_g N_SCE_c_365_n N_SCE_M1023_g N_SCE_c_366_n
+ N_SCE_c_367_n SCE SCE N_SCE_c_368_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%SCE
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%D N_D_M1026_g N_D_M1040_g D D N_D_c_421_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%D
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_27_55# N_A_27_55#_M1001_s N_A_27_55#_M1016_s
+ N_A_27_55#_c_468_n N_A_27_55#_M1004_g N_A_27_55#_c_464_n N_A_27_55#_M1003_g
+ N_A_27_55#_c_466_n N_A_27_55#_c_467_n N_A_27_55#_c_472_n N_A_27_55#_c_473_n
+ N_A_27_55#_c_474_n N_A_27_55#_c_475_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_27_55#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%SCD N_SCD_M1052_g N_SCD_M1022_g N_SCD_c_544_n
+ N_SCD_c_549_n SCD N_SCD_c_545_n N_SCD_c_546_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%SCD
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%RESET_B N_RESET_B_c_584_n N_RESET_B_M1028_g
+ N_RESET_B_M1049_g N_RESET_B_c_586_n N_RESET_B_M1011_g N_RESET_B_M1007_g
+ N_RESET_B_c_601_n N_RESET_B_c_602_n N_RESET_B_M1008_g N_RESET_B_c_589_n
+ N_RESET_B_c_590_n N_RESET_B_M1005_g N_RESET_B_c_592_n N_RESET_B_c_593_n
+ N_RESET_B_c_594_n N_RESET_B_c_595_n N_RESET_B_c_596_n N_RESET_B_c_597_n
+ N_RESET_B_c_607_n N_RESET_B_c_608_n RESET_B N_RESET_B_c_598_n
+ N_RESET_B_c_610_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%RESET_B
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_742_63# N_A_742_63#_M1038_s
+ N_A_742_63#_M1042_d N_A_742_63#_M1018_g N_A_742_63#_M1021_g
+ N_A_742_63#_c_781_n N_A_742_63#_c_782_n N_A_742_63#_M1000_g
+ N_A_742_63#_c_784_n N_A_742_63#_M1037_g N_A_742_63#_c_767_n
+ N_A_742_63#_M1041_g N_A_742_63#_M1050_g N_A_742_63#_c_768_n
+ N_A_742_63#_c_769_n N_A_742_63#_M1030_g N_A_742_63#_c_770_n
+ N_A_742_63#_M1044_g N_A_742_63#_c_789_n N_A_742_63#_c_771_n
+ N_A_742_63#_c_772_n N_A_742_63#_c_791_n N_A_742_63#_c_792_n
+ N_A_742_63#_c_793_n N_A_742_63#_c_853_p N_A_742_63#_c_794_n
+ N_A_742_63#_c_842_p N_A_742_63#_c_795_n N_A_742_63#_c_796_n
+ N_A_742_63#_c_797_n N_A_742_63#_c_773_n N_A_742_63#_c_798_n
+ N_A_742_63#_c_799_n N_A_742_63#_c_800_n N_A_742_63#_c_774_n
+ N_A_742_63#_c_802_n N_A_742_63#_c_803_n N_A_742_63#_c_804_n
+ N_A_742_63#_c_805_n N_A_742_63#_c_865_p N_A_742_63#_c_775_n
+ N_A_742_63#_c_776_n N_A_742_63#_c_777_n N_A_742_63#_c_778_n
+ N_A_742_63#_c_779_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_742_63#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_666_89# N_A_666_89#_M1018_s
+ N_A_666_89#_M1021_s N_A_666_89#_c_1066_n N_A_666_89#_M1045_g
+ N_A_666_89#_M1053_g N_A_666_89#_c_1067_n N_A_666_89#_M1034_g
+ N_A_666_89#_c_1068_n N_A_666_89#_M1015_g N_A_666_89#_M1013_g
+ N_A_666_89#_c_1070_n N_A_666_89#_M1002_g N_A_666_89#_c_1072_n
+ N_A_666_89#_c_1073_n N_A_666_89#_c_1080_n N_A_666_89#_c_1081_n
+ N_A_666_89#_c_1082_n N_A_666_89#_c_1083_n N_A_666_89#_c_1074_n
+ N_A_666_89#_c_1128_p N_A_666_89#_c_1085_n N_A_666_89#_c_1075_n
+ N_A_666_89#_c_1076_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_666_89#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1343_51# N_A_1343_51#_M1032_d
+ N_A_1343_51#_M1044_s N_A_1343_51#_M1029_d N_A_1343_51#_M1015_d
+ N_A_1343_51#_M1012_g N_A_1343_51#_c_1263_n N_A_1343_51#_M1010_g
+ N_A_1343_51#_M1035_g N_A_1343_51#_c_1266_n N_A_1343_51#_c_1267_n
+ N_A_1343_51#_c_1268_n N_A_1343_51#_c_1269_n N_A_1343_51#_c_1270_n
+ N_A_1343_51#_c_1271_n N_A_1343_51#_c_1272_n N_A_1343_51#_c_1315_n
+ N_A_1343_51#_c_1273_n N_A_1343_51#_c_1274_n N_A_1343_51#_c_1275_n
+ N_A_1343_51#_c_1276_n N_A_1343_51#_c_1366_p N_A_1343_51#_c_1367_p
+ N_A_1343_51#_c_1277_n N_A_1343_51#_c_1278_n N_A_1343_51#_c_1279_n
+ N_A_1343_51#_c_1340_n N_A_1343_51#_c_1280_n N_A_1343_51#_c_1281_n
+ N_A_1343_51#_c_1288_n N_A_1343_51#_c_1289_n N_A_1343_51#_c_1282_n
+ N_A_1343_51#_c_1283_n N_A_1343_51#_c_1290_n N_A_1343_51#_c_1284_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1343_51#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1724_21# N_A_1724_21#_M1020_d
+ N_A_1724_21#_M1017_d N_A_1724_21#_M1027_g N_A_1724_21#_M1014_g
+ N_A_1724_21#_c_1481_n N_A_1724_21#_c_1482_n N_A_1724_21#_c_1483_n
+ N_A_1724_21#_c_1484_n N_A_1724_21#_c_1485_n N_A_1724_21#_c_1486_n
+ N_A_1724_21#_c_1487_n N_A_1724_21#_c_1495_n N_A_1724_21#_c_1496_n
+ N_A_1724_21#_c_1497_n N_A_1724_21#_c_1488_n N_A_1724_21#_c_1489_n
+ N_A_1724_21#_c_1490_n N_A_1724_21#_c_1491_n N_A_1724_21#_c_1492_n
+ N_A_1724_21#_c_1493_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1724_21#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1113_419# N_A_1113_419#_M1041_d
+ N_A_1113_419#_M1037_d N_A_1113_419#_M1011_s N_A_1113_419#_c_1634_n
+ N_A_1113_419#_M1048_g N_A_1113_419#_M1029_g N_A_1113_419#_c_1636_n
+ N_A_1113_419#_M1032_g N_A_1113_419#_c_1637_n N_A_1113_419#_c_1638_n
+ N_A_1113_419#_c_1639_n N_A_1113_419#_c_1642_n N_A_1113_419#_c_1668_n
+ N_A_1113_419#_c_1672_n N_A_1113_419#_c_1699_n N_A_1113_419#_c_1643_n
+ N_A_1113_419#_c_1653_n N_A_1113_419#_c_1644_n N_A_1113_419#_c_1645_n
+ N_A_1113_419#_c_1646_n N_A_1113_419#_c_1656_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1113_419#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%CLK_N N_CLK_N_M1038_g N_CLK_N_c_1779_n
+ N_CLK_N_M1042_g N_CLK_N_c_1780_n CLK_N N_CLK_N_c_1781_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%CLK_N
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%SLEEP_B N_SLEEP_B_c_1826_n N_SLEEP_B_M1039_g
+ N_SLEEP_B_M1019_g N_SLEEP_B_c_1828_n N_SLEEP_B_M1043_g N_SLEEP_B_c_1835_n
+ N_SLEEP_B_M1017_g N_SLEEP_B_c_1829_n N_SLEEP_B_M1006_g N_SLEEP_B_c_1830_n
+ N_SLEEP_B_c_1831_n N_SLEEP_B_c_1832_n N_SLEEP_B_M1020_g SLEEP_B
+ N_SLEEP_B_c_1833_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%SLEEP_B
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2999_73# N_A_2999_73#_M1009_d
+ N_A_2999_73#_M1005_d N_A_2999_73#_M1051_g N_A_2999_73#_M1031_g
+ N_A_2999_73#_c_1928_n N_A_2999_73#_c_1929_n N_A_2999_73#_c_1924_n
+ N_A_2999_73#_c_1931_n N_A_2999_73#_c_1925_n N_A_2999_73#_c_1932_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2999_73#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2717_427# N_A_2717_427#_M1044_d
+ N_A_2717_427#_M1030_d N_A_2717_427#_c_1997_n N_A_2717_427#_M1009_g
+ N_A_2717_427#_c_1998_n N_A_2717_427#_c_1999_n N_A_2717_427#_M1046_g
+ N_A_2717_427#_c_2001_n N_A_2717_427#_c_2002_n N_A_2717_427#_c_2017_n
+ N_A_2717_427#_c_2018_n N_A_2717_427#_M1036_g N_A_2717_427#_M1047_g
+ N_A_2717_427#_c_2004_n N_A_2717_427#_c_2005_n N_A_2717_427#_c_2021_n
+ N_A_2717_427#_c_2022_n N_A_2717_427#_c_2023_n N_A_2717_427#_c_2006_n
+ N_A_2717_427#_c_2007_n N_A_2717_427#_c_2008_n N_A_2717_427#_c_2009_n
+ N_A_2717_427#_c_2010_n N_A_2717_427#_c_2011_n N_A_2717_427#_c_2012_n
+ N_A_2717_427#_c_2025_n N_A_2717_427#_c_2013_n N_A_2717_427#_c_2014_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2717_427#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_3368_57# N_A_3368_57#_M1036_s
+ N_A_3368_57#_M1047_s N_A_3368_57#_M1033_g N_A_3368_57#_M1024_g
+ N_A_3368_57#_c_2158_n N_A_3368_57#_c_2159_n N_A_3368_57#_c_2166_n
+ N_A_3368_57#_c_2167_n N_A_3368_57#_c_2160_n N_A_3368_57#_c_2161_n
+ N_A_3368_57#_c_2162_n N_A_3368_57#_c_2163_n N_A_3368_57#_c_2164_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_3368_57#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%VPWR N_VPWR_M1016_d N_VPWR_M1052_d
+ N_VPWR_M1021_d N_VPWR_M1031_d N_VPWR_M1046_d N_VPWR_M1047_d N_VPWR_c_2221_n
+ N_VPWR_c_2222_n N_VPWR_c_2223_n N_VPWR_c_2224_n N_VPWR_c_2225_n
+ N_VPWR_c_2226_n N_VPWR_c_2227_n N_VPWR_c_2228_n N_VPWR_c_2229_n
+ N_VPWR_c_2230_n N_VPWR_c_2231_n N_VPWR_c_2232_n N_VPWR_c_2233_n
+ N_VPWR_c_2234_n VPWR N_VPWR_c_2235_n N_VPWR_c_2236_n N_VPWR_c_2237_n
+ N_VPWR_c_2220_n N_VPWR_c_2239_n N_VPWR_c_2240_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%VPWR
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_305_97# N_A_305_97#_M1023_d
+ N_A_305_97#_M1034_d N_A_305_97#_M1026_d N_A_305_97#_M1049_d
+ N_A_305_97#_c_2391_n N_A_305_97#_c_2415_n N_A_305_97#_c_2404_n
+ N_A_305_97#_c_2405_n N_A_305_97#_c_2392_n N_A_305_97#_c_2393_n
+ N_A_305_97#_c_2394_n N_A_305_97#_c_2395_n N_A_305_97#_c_2407_n
+ N_A_305_97#_c_2408_n N_A_305_97#_c_2409_n N_A_305_97#_c_2410_n
+ N_A_305_97#_c_2396_n N_A_305_97#_c_2397_n N_A_305_97#_c_2398_n
+ N_A_305_97#_c_2458_n N_A_305_97#_c_2411_n N_A_305_97#_c_2399_n
+ N_A_305_97#_c_2461_n N_A_305_97#_c_2463_n N_A_305_97#_c_2400_n
+ N_A_305_97#_c_2401_n N_A_305_97#_c_2412_n N_A_305_97#_c_2402_n
+ N_A_305_97#_c_2413_n N_A_305_97#_c_2403_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_305_97#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%KAPWR N_KAPWR_M1010_d N_KAPWR_M1014_d
+ N_KAPWR_M1042_s N_KAPWR_M1019_d N_KAPWR_c_2586_n N_KAPWR_c_2587_n
+ N_KAPWR_c_2588_n KAPWR N_KAPWR_c_2590_n N_KAPWR_c_2591_n N_KAPWR_c_2592_n
+ N_KAPWR_c_2593_n N_KAPWR_c_2594_n KAPWR N_KAPWR_c_2595_n N_KAPWR_c_2659_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%KAPWR
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2562_427# N_A_2562_427#_M1050_s
+ N_A_2562_427#_M1031_s N_A_2562_427#_c_2779_n N_A_2562_427#_c_2780_n
+ N_A_2562_427#_c_2781_n N_A_2562_427#_c_2782_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2562_427#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%Q N_Q_M1033_d N_Q_M1024_d Q Q Q Q Q
+ N_Q_c_2814_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%Q
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%VGND N_VGND_M1001_d N_VGND_M1018_d
+ N_VGND_M1007_s N_VGND_M1027_d N_VGND_M1043_d N_VGND_M1051_d N_VGND_M1036_d
+ N_VGND_c_2830_n N_VGND_c_2831_n N_VGND_c_2832_n N_VGND_c_2833_n
+ N_VGND_c_2834_n N_VGND_c_2835_n N_VGND_c_2836_n N_VGND_c_2837_n
+ N_VGND_c_2838_n VGND N_VGND_c_2839_n N_VGND_c_2840_n N_VGND_c_2841_n
+ N_VGND_c_2842_n N_VGND_c_2843_n N_VGND_c_2844_n N_VGND_c_2845_n
+ N_VGND_c_2846_n N_VGND_c_2847_n N_VGND_c_2848_n N_VGND_c_2849_n
+ N_VGND_c_2850_n N_VGND_c_2851_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%VGND
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%noxref_30 N_noxref_30_M1023_s
+ N_noxref_30_M1022_d N_noxref_30_c_2991_n N_noxref_30_c_2992_n
+ N_noxref_30_c_2993_n N_noxref_30_c_2994_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%noxref_30
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%noxref_32 N_noxref_32_M1003_d
+ N_noxref_32_M1028_d N_noxref_32_c_3021_n N_noxref_32_c_3022_n
+ N_noxref_32_c_3023_n N_noxref_32_c_3024_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%noxref_32
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1009_107# N_A_1009_107#_M1041_s
+ N_A_1009_107#_M1012_s N_A_1009_107#_c_3056_n
+ PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1009_107#
x_PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1453_77# N_A_1453_77#_M1035_d
+ N_A_1453_77#_M1007_d N_A_1453_77#_c_3075_n N_A_1453_77#_c_3076_n
+ N_A_1453_77#_c_3077_n PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1453_77#
cc_1 VNB N_SCE_M1001_g 0.0375416f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.485
cc_2 VNB N_SCE_c_363_n 0.0386169f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.09
cc_3 VNB N_SCE_c_364_n 0.00865403f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.69
cc_4 VNB N_SCE_c_365_n 0.0199839f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.015
cc_5 VNB N_SCE_c_366_n 0.030387f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.09
cc_6 VNB N_SCE_c_367_n 0.00247672f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_7 VNB N_SCE_c_368_n 0.0343515f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_8 VNB N_D_M1040_g 0.0366899f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_9 VNB D 0.0120547f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.69
cc_10 VNB N_D_c_421_n 0.0344073f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.695
cc_11 VNB N_A_27_55#_c_464_n 0.0144384f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.69
cc_12 VNB N_A_27_55#_M1003_g 0.0264456f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.775
cc_13 VNB N_A_27_55#_c_466_n 0.00950552f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.695
cc_14 VNB N_A_27_55#_c_467_n 0.0693295f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.09
cc_15 VNB N_SCD_M1022_g 0.0576195f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_16 VNB N_SCD_c_544_n 0.00673706f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.09
cc_17 VNB N_SCD_c_545_n 0.0140078f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.015
cc_18 VNB N_SCD_c_546_n 0.00235078f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.695
cc_19 VNB N_RESET_B_c_584_n 0.018081f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.015
cc_20 VNB N_RESET_B_M1049_g 0.0415463f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_21 VNB N_RESET_B_c_586_n 0.0448942f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.09
cc_22 VNB N_RESET_B_M1007_g 0.050938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_RESET_B_M1008_g 0.0369473f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.615
cc_24 VNB N_RESET_B_c_589_n 0.0198714f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_25 VNB N_RESET_B_c_590_n 0.008402f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_26 VNB N_RESET_B_M1005_g 0.00317395f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_27 VNB N_RESET_B_c_592_n 0.0398677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_RESET_B_c_593_n 0.0203426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_RESET_B_c_594_n 0.0109855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_RESET_B_c_595_n 0.0413035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_RESET_B_c_596_n 0.0510812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_RESET_B_c_597_n 0.00845028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_c_598_n 0.00457752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_742_63#_M1018_g 0.0922719f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.09
cc_35 VNB N_A_742_63#_c_767_n 0.0171436f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_36 VNB N_A_742_63#_c_768_n 0.00918763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_742_63#_c_769_n 0.0157788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_742_63#_c_770_n 0.0227394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_742_63#_c_771_n 0.026469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_742_63#_c_772_n 0.00526036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_742_63#_c_773_n 0.0107483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_742_63#_c_774_n 0.0025136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_742_63#_c_775_n 0.00305859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_742_63#_c_776_n 0.00438232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_742_63#_c_777_n 0.00879077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_742_63#_c_778_n 0.0400396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_742_63#_c_779_n 0.0213644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_666_89#_c_1066_n 0.0140922f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_49 VNB N_A_666_89#_c_1067_n 0.0153644f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.775
cc_50 VNB N_A_666_89#_c_1068_n 0.0416464f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.015
cc_51 VNB N_A_666_89#_M1013_g 0.0220541f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_52 VNB N_A_666_89#_c_1070_n 0.0220245f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_53 VNB N_A_666_89#_M1002_g 0.0189645f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_54 VNB N_A_666_89#_c_1072_n 0.00448011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_666_89#_c_1073_n 0.00440585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_666_89#_c_1074_n 0.00338152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_666_89#_c_1075_n 0.0346839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_666_89#_c_1076_n 0.00463183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1343_51#_c_1263_n 0.0126036f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.015
cc_60 VNB N_A_1343_51#_M1010_g 0.0369257f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.165
cc_61 VNB N_A_1343_51#_M1035_g 0.0313245f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_62 VNB N_A_1343_51#_c_1266_n 0.0197839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1343_51#_c_1267_n 0.0094458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1343_51#_c_1268_n 9.88085e-19 $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_65 VNB N_A_1343_51#_c_1269_n 0.0139291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1343_51#_c_1270_n 0.00309434f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.665
cc_67 VNB N_A_1343_51#_c_1271_n 0.00545342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1343_51#_c_1272_n 0.0108356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1343_51#_c_1273_n 0.00941569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1343_51#_c_1274_n 0.0327528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1343_51#_c_1275_n 2.71348e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1343_51#_c_1276_n 5.5124e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1343_51#_c_1277_n 0.00101683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1343_51#_c_1278_n 0.00304019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1343_51#_c_1279_n 0.0158183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1343_51#_c_1280_n 0.00634049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1343_51#_c_1281_n 0.00159323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1343_51#_c_1282_n 0.0142433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1343_51#_c_1283_n 0.00558319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1343_51#_c_1284_n 0.0453998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1724_21#_M1027_g 0.0396181f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.09
cc_82 VNB N_A_1724_21#_c_1481_n 0.0180885f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.775
cc_83 VNB N_A_1724_21#_c_1482_n 0.00578298f $X=-0.19 $Y=-0.245 $X2=1.45
+ $Y2=0.695
cc_84 VNB N_A_1724_21#_c_1483_n 0.0107593f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.695
cc_85 VNB N_A_1724_21#_c_1484_n 0.00351845f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.165
cc_86 VNB N_A_1724_21#_c_1485_n 4.01303e-19 $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.615
cc_87 VNB N_A_1724_21#_c_1486_n 0.00996167f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_88 VNB N_A_1724_21#_c_1487_n 0.00137663f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_89 VNB N_A_1724_21#_c_1488_n 0.00528483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1724_21#_c_1489_n 0.00893064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1724_21#_c_1490_n 0.00802614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1724_21#_c_1491_n 0.024563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1724_21#_c_1492_n 5.13554e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1724_21#_c_1493_n 0.0031054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1113_419#_c_1634_n 0.015322f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.09
cc_96 VNB N_A_1113_419#_M1029_g 0.0244342f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.775
cc_97 VNB N_A_1113_419#_c_1636_n 0.0193001f $X=-0.19 $Y=-0.245 $X2=1.45
+ $Y2=1.015
cc_98 VNB N_A_1113_419#_c_1637_n 0.0356626f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.165
cc_99 VNB N_A_1113_419#_c_1638_n 0.0308257f $X=-0.19 $Y=-0.245 $X2=0.662
+ $Y2=1.09
cc_100 VNB N_A_1113_419#_c_1639_n 0.0286803f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.69
cc_101 VNB N_CLK_N_M1038_g 0.047446f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.485
cc_102 VNB N_CLK_N_c_1779_n 0.00370131f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.765
cc_103 VNB N_CLK_N_c_1780_n 0.0224327f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.09
cc_104 VNB N_CLK_N_c_1781_n 0.00627578f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.775
cc_105 VNB N_SLEEP_B_c_1826_n 0.0140611f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.015
cc_106 VNB N_SLEEP_B_M1019_g 8.393e-19 $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.775
cc_107 VNB N_SLEEP_B_c_1828_n 0.0163877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_SLEEP_B_c_1829_n 0.0171996f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.775
cc_109 VNB N_SLEEP_B_c_1830_n 0.0218977f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.015
cc_110 VNB N_SLEEP_B_c_1831_n 0.109673f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.695
cc_111 VNB N_SLEEP_B_c_1832_n 0.0180564f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.695
cc_112 VNB N_SLEEP_B_c_1833_n 0.00254511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2999_73#_M1051_g 0.051887f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.09
cc_114 VNB N_A_2999_73#_c_1924_n 0.00650515f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_115 VNB N_A_2999_73#_c_1925_n 0.00156783f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.26
cc_116 VNB N_A_2717_427#_c_1997_n 0.0182289f $X=-0.19 $Y=-0.245 $X2=0.66
+ $Y2=2.775
cc_117 VNB N_A_2717_427#_c_1998_n 0.0158153f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.09
cc_118 VNB N_A_2717_427#_c_1999_n 0.00901392f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.69
cc_119 VNB N_A_2717_427#_M1046_g 0.00438762f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=2.775
cc_120 VNB N_A_2717_427#_c_2001_n 0.00537274f $X=-0.19 $Y=-0.245 $X2=1.45
+ $Y2=1.015
cc_121 VNB N_A_2717_427#_c_2002_n 0.0337829f $X=-0.19 $Y=-0.245 $X2=1.45
+ $Y2=0.695
cc_122 VNB N_A_2717_427#_M1036_g 0.0266548f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_123 VNB N_A_2717_427#_c_2004_n 0.0051639f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.26
cc_124 VNB N_A_2717_427#_c_2005_n 0.00854107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2717_427#_c_2006_n 0.00286233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2717_427#_c_2007_n 0.0107535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_2717_427#_c_2008_n 0.00611235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_2717_427#_c_2009_n 0.00416261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_2717_427#_c_2010_n 0.0168433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_2717_427#_c_2011_n 0.00266269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_2717_427#_c_2012_n 0.0106997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_2717_427#_c_2013_n 0.00979795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_2717_427#_c_2014_n 0.0889665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_3368_57#_M1033_g 0.0278682f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.09
cc_135 VNB N_A_3368_57#_M1024_g 6.56926e-19 $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=1.765
cc_136 VNB N_A_3368_57#_c_2158_n 0.0443189f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=2.775
cc_137 VNB N_A_3368_57#_c_2159_n 0.0158658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_3368_57#_c_2160_n 0.00713609f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.615
cc_139 VNB N_A_3368_57#_c_2161_n 0.00327839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_3368_57#_c_2162_n 0.0086727f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_141 VNB N_A_3368_57#_c_2163_n 2.35235e-19 $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.665
cc_142 VNB N_A_3368_57#_c_2164_n 0.00418528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VPWR_c_2220_n 0.760753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_305_97#_c_2391_n 0.00309576f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=1.765
cc_145 VNB N_A_305_97#_c_2392_n 0.00549919f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_146 VNB N_A_305_97#_c_2393_n 0.0255696f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_147 VNB N_A_305_97#_c_2394_n 0.00290025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_A_305_97#_c_2395_n 0.0102718f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_149 VNB N_A_305_97#_c_2396_n 0.00996669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_A_305_97#_c_2397_n 0.00503025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_A_305_97#_c_2398_n 0.00331057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_A_305_97#_c_2399_n 0.00661983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_305_97#_c_2400_n 0.00882927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_305_97#_c_2401_n 6.0718e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_A_305_97#_c_2402_n 0.00122144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_A_305_97#_c_2403_n 0.00782529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_Q_c_2814_n 0.0577541f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.695
cc_158 VNB N_VGND_c_2830_n 0.0121964f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_159 VNB N_VGND_c_2831_n 0.0127389f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_160 VNB N_VGND_c_2832_n 0.0182829f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.26
cc_161 VNB N_VGND_c_2833_n 0.00432763f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.665
cc_162 VNB N_VGND_c_2834_n 0.00552922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2835_n 0.0111723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2836_n 0.0116956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2837_n 0.0676497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2838_n 0.00477645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2839_n 0.0160515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2840_n 0.0755706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2841_n 0.0867356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2842_n 0.0713912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2843_n 0.0481722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2844_n 0.0189138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2845_n 0.982109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2846_n 0.0054376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2847_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2848_n 0.0134666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2849_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2850_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2851_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_noxref_30_c_2991_n 0.00851461f $X=-0.19 $Y=-0.245 $X2=1.375
+ $Y2=1.09
cc_181 VNB N_noxref_30_c_2992_n 0.022606f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.69
cc_182 VNB N_noxref_30_c_2993_n 0.00391982f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.69
cc_183 VNB N_noxref_30_c_2994_n 0.0131651f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.765
cc_184 VNB N_noxref_32_c_3021_n 3.12925e-19 $X=-0.19 $Y=-0.245 $X2=1.375
+ $Y2=1.09
cc_185 VNB N_noxref_32_c_3022_n 0.036729f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.69
cc_186 VNB N_noxref_32_c_3023_n 0.0029575f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.69
cc_187 VNB N_noxref_32_c_3024_n 0.0113059f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.775
cc_188 VNB N_A_1009_107#_c_3056_n 0.0266399f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.69
cc_189 VNB N_A_1453_77#_c_3075_n 0.00969341f $X=-0.19 $Y=-0.245 $X2=0.66
+ $Y2=2.775
cc_190 VNB N_A_1453_77#_c_3076_n 0.00631975f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.09
cc_191 VNB N_A_1453_77#_c_3077_n 0.00249901f $X=-0.19 $Y=-0.245 $X2=1.16
+ $Y2=2.775
cc_192 VPB N_SCE_M1016_g 0.0564316f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_193 VPB N_SCE_c_364_n 0.00676271f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.69
cc_194 VPB N_SCE_M1025_g 0.0456733f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.775
cc_195 VPB N_SCE_c_367_n 0.00935095f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.69
cc_196 VPB SCE 0.00176604f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_197 VPB N_D_M1026_g 0.0489795f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.485
cc_198 VPB D 0.00502394f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.69
cc_199 VPB N_D_c_421_n 0.011916f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_200 VPB N_A_27_55#_c_468_n 0.049437f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_201 VPB N_A_27_55#_M1004_g 0.0224687f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=1.09
cc_202 VPB N_A_27_55#_c_464_n 0.00612843f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.69
cc_203 VPB N_A_27_55#_c_467_n 0.0159236f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.09
cc_204 VPB N_A_27_55#_c_472_n 0.0398957f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_205 VPB N_A_27_55#_c_473_n 0.0181773f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_206 VPB N_A_27_55#_c_474_n 0.00225859f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_207 VPB N_A_27_55#_c_475_n 0.0206961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_SCD_M1052_g 0.0233028f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.485
cc_209 VPB N_SCD_c_544_n 0.0203101f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.09
cc_210 VPB N_SCD_c_549_n 0.0163755f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.69
cc_211 VPB N_SCD_c_545_n 0.00273741f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=1.015
cc_212 VPB N_SCD_c_546_n 0.0055139f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_213 VPB N_RESET_B_M1049_g 0.0197869f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_214 VPB N_RESET_B_M1011_g 0.0395261f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.765
cc_215 VPB N_RESET_B_c_601_n 0.540985f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_216 VPB N_RESET_B_c_602_n 0.0177998f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_217 VPB N_RESET_B_M1005_g 0.0505697f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_218 VPB N_RESET_B_c_593_n 0.0170954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_RESET_B_c_594_n 0.00421923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_RESET_B_c_597_n 0.00529045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_RESET_B_c_607_n 0.0157369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_RESET_B_c_608_n 6.90525e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_RESET_B_c_598_n 0.00638557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_RESET_B_c_610_n 0.00145355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_742_63#_M1018_g 0.0378247f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=1.09
cc_226 VPB N_A_742_63#_c_781_n 0.0853014f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.765
cc_227 VPB N_A_742_63#_c_782_n 0.012806f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.775
cc_228 VPB N_A_742_63#_M1000_g 0.0347761f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_229 VPB N_A_742_63#_c_784_n 0.0214815f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_230 VPB N_A_742_63#_M1037_g 0.0301509f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_231 VPB N_A_742_63#_M1050_g 0.032848f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_232 VPB N_A_742_63#_c_768_n 8.30539e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_742_63#_M1030_g 0.0366085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_742_63#_c_789_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_742_63#_c_772_n 6.09015e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_742_63#_c_791_n 0.00982946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_742_63#_c_792_n 0.00183425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_742_63#_c_793_n 0.00476816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_742_63#_c_794_n 0.00575043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_742_63#_c_795_n 2.30474e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_742_63#_c_796_n 0.0201547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_742_63#_c_797_n 0.00125024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_742_63#_c_798_n 0.0140695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_742_63#_c_799_n 0.00396194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_742_63#_c_800_n 0.00237991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_742_63#_c_774_n 0.00195643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_742_63#_c_802_n 5.67166e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_742_63#_c_803_n 0.00366156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_742_63#_c_804_n 0.00210016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_742_63#_c_805_n 8.87845e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_742_63#_c_776_n 0.00236325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_742_63#_c_778_n 0.00306983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_742_63#_c_779_n 0.0204516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_666_89#_M1053_g 0.0272671f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.69
cc_255 VPB N_A_666_89#_c_1068_n 0.0141435f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=1.015
cc_256 VPB N_A_666_89#_M1015_g 0.0204433f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_257 VPB N_A_666_89#_c_1080_n 0.00947399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_666_89#_c_1081_n 0.00173447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_666_89#_c_1082_n 0.0304812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_666_89#_c_1083_n 0.0011951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_666_89#_c_1074_n 0.00181249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_666_89#_c_1085_n 0.00148634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_666_89#_c_1075_n 0.00954177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_666_89#_c_1076_n 9.34293e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_1343_51#_M1010_g 0.033676f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.165
cc_266 VPB N_A_1343_51#_c_1271_n 0.00196742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_1343_51#_c_1280_n 0.00229163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_1343_51#_c_1288_n 0.00591233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_1343_51#_c_1289_n 0.00632228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_1343_51#_c_1290_n 0.00620028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_1343_51#_c_1284_n 0.0169708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_1724_21#_M1014_g 0.0220573f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.765
cc_273 VPB N_A_1724_21#_c_1495_n 0.00535614f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.58
cc_274 VPB N_A_1724_21#_c_1496_n 0.00926337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_1724_21#_c_1497_n 0.0153426f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_276 VPB N_A_1724_21#_c_1490_n 0.00260425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_1724_21#_c_1491_n 0.0104223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_1724_21#_c_1492_n 7.8745e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_1113_419#_M1029_g 0.0321176f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.775
cc_280 VPB N_A_1113_419#_c_1639_n 0.0410517f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.69
cc_281 VPB N_A_1113_419#_c_1642_n 3.75833e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_A_1113_419#_c_1643_n 0.0141025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_1113_419#_c_1644_n 0.00347342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_1113_419#_c_1645_n 0.00188761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_A_1113_419#_c_1646_n 0.0485527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_CLK_N_c_1779_n 0.04913f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.765
cc_287 VPB N_CLK_N_c_1780_n 0.0363833f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=1.09
cc_288 VPB N_CLK_N_c_1781_n 0.00199098f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.775
cc_289 VPB N_SLEEP_B_M1019_g 0.0320902f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.775
cc_290 VPB N_SLEEP_B_c_1835_n 0.0201318f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.69
cc_291 VPB N_SLEEP_B_c_1831_n 0.0127644f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_292 VPB N_SLEEP_B_c_1833_n 0.0030218f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_A_2999_73#_M1051_g 0.0109766f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=1.09
cc_294 VPB N_A_2999_73#_M1031_g 0.0206023f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.765
cc_295 VPB N_A_2999_73#_c_1928_n 0.00433844f $X=-0.19 $Y=1.655 $X2=1.16
+ $Y2=2.775
cc_296 VPB N_A_2999_73#_c_1929_n 0.00219715f $X=-0.19 $Y=1.655 $X2=0.75
+ $Y2=1.615
cc_297 VPB N_A_2999_73#_c_1924_n 0.00139922f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.58
cc_298 VPB N_A_2999_73#_c_1931_n 0.00229455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_A_2999_73#_c_1932_n 0.055139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_A_2717_427#_M1046_g 0.0487441f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.775
cc_301 VPB N_A_2717_427#_c_2001_n 0.0113122f $X=-0.19 $Y=1.655 $X2=1.45
+ $Y2=1.015
cc_302 VPB N_A_2717_427#_c_2017_n 0.0358718f $X=-0.19 $Y=1.655 $X2=0.75
+ $Y2=1.165
cc_303 VPB N_A_2717_427#_c_2018_n 0.0118181f $X=-0.19 $Y=1.655 $X2=0.662
+ $Y2=1.09
cc_304 VPB N_A_2717_427#_M1047_g 0.0418064f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_305 VPB N_A_2717_427#_c_2005_n 0.00679575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_A_2717_427#_c_2021_n 0.0228296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_A_2717_427#_c_2022_n 0.0031471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_A_2717_427#_c_2023_n 0.0105906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_309 VPB N_A_2717_427#_c_2006_n 0.00349455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_A_2717_427#_c_2025_n 0.00750082f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_A_3368_57#_M1024_g 0.0268182f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.765
cc_312 VPB N_A_3368_57#_c_2166_n 0.00343529f $X=-0.19 $Y=1.655 $X2=1.45
+ $Y2=1.015
cc_313 VPB N_A_3368_57#_c_2167_n 0.00367448f $X=-0.19 $Y=1.655 $X2=1.45
+ $Y2=0.695
cc_314 VPB N_A_3368_57#_c_2163_n 0.0105628f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.665
cc_315 VPB N_VPWR_c_2221_n 0.00626187f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.09
cc_316 VPB N_VPWR_c_2222_n 0.00240024f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_317 VPB N_VPWR_c_2223_n 0.0081958f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_318 VPB N_VPWR_c_2224_n 0.0103201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_2225_n 0.0294251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_2226_n 0.011762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_2227_n 0.0221079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_2228_n 0.00510509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_2229_n 0.0413582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_2230_n 0.00356769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2231_n 0.031889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_2232_n 0.00223798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_2233_n 0.0192019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2234_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_2235_n 0.267649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_2236_n 0.0202711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2237_n 0.0184065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_2220_n 0.0577153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_2239_n 0.00330333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2240_n 0.00477947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_A_305_97#_c_2404_n 0.0165463f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.09
cc_336 VPB N_A_305_97#_c_2405_n 0.0033919f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.615
cc_337 VPB N_A_305_97#_c_2395_n 0.0112312f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_338 VPB N_A_305_97#_c_2407_n 0.00716897f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_339 VPB N_A_305_97#_c_2408_n 0.0119562f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_340 VPB N_A_305_97#_c_2409_n 0.00333638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_A_305_97#_c_2410_n 0.00651509f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.665
cc_342 VPB N_A_305_97#_c_2411_n 0.00406246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_343 VPB N_A_305_97#_c_2412_n 0.00530346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_344 VPB N_A_305_97#_c_2413_n 0.00129007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_345 VPB N_KAPWR_c_2586_n 0.00322005f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.775
cc_346 VPB N_KAPWR_c_2587_n 0.0176974f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=1.015
cc_347 VPB N_KAPWR_c_2588_n 0.00688137f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_348 VPB KAPWR 0.0324494f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.165
cc_349 VPB N_KAPWR_c_2590_n 0.0116888f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.26
cc_350 VPB N_KAPWR_c_2591_n 0.00919158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_351 VPB N_KAPWR_c_2592_n 9.47438e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_352 VPB N_KAPWR_c_2593_n 0.0291736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_353 VPB N_KAPWR_c_2594_n 0.0012903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_354 VPB N_KAPWR_c_2595_n 0.0157473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_355 VPB N_A_2562_427#_c_2779_n 0.0106727f $X=-0.19 $Y=1.655 $X2=1.375
+ $Y2=1.09
cc_356 VPB N_A_2562_427#_c_2780_n 0.0372314f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.69
cc_357 VPB N_A_2562_427#_c_2781_n 0.0078874f $X=-0.19 $Y=1.655 $X2=0.915
+ $Y2=1.69
cc_358 VPB N_A_2562_427#_c_2782_n 0.00559087f $X=-0.19 $Y=1.655 $X2=1.16
+ $Y2=2.775
cc_359 VPB N_Q_c_2814_n 0.0488589f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=0.695
cc_360 N_SCE_M1025_g N_D_M1026_g 0.044806f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_361 N_SCE_c_365_n N_D_M1040_g 0.022411f $X=1.45 $Y=1.015 $X2=0 $Y2=0
cc_362 N_SCE_c_363_n D 0.0141595f $X=1.375 $Y=1.09 $X2=0 $Y2=0
cc_363 N_SCE_c_364_n D 0.00819333f $X=1.085 $Y=1.69 $X2=0 $Y2=0
cc_364 N_SCE_M1025_g D 0.00248486f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_365 SCE D 0.0499073f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_366 N_SCE_c_368_n D 0.00433538f $X=0.75 $Y=1.26 $X2=0 $Y2=0
cc_367 N_SCE_c_363_n N_D_c_421_n 0.00327785f $X=1.375 $Y=1.09 $X2=0 $Y2=0
cc_368 N_SCE_c_364_n N_D_c_421_n 0.044806f $X=1.085 $Y=1.69 $X2=0 $Y2=0
cc_369 SCE N_D_c_421_n 3.80952e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_370 N_SCE_c_368_n N_D_c_421_n 0.00223401f $X=0.75 $Y=1.26 $X2=0 $Y2=0
cc_371 N_SCE_M1001_g N_A_27_55#_c_467_n 0.0197422f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_372 SCE N_A_27_55#_c_467_n 0.0422236f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_373 N_SCE_c_368_n N_A_27_55#_c_467_n 0.0201206f $X=0.75 $Y=1.26 $X2=0 $Y2=0
cc_374 N_SCE_M1016_g N_A_27_55#_c_472_n 0.0248184f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_375 N_SCE_M1025_g N_A_27_55#_c_472_n 0.00172721f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_376 N_SCE_M1016_g N_A_27_55#_c_473_n 0.00454477f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_377 SCE N_A_27_55#_c_473_n 0.00203275f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_378 N_SCE_M1016_g N_A_27_55#_c_475_n 0.00893655f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_379 N_SCE_M1025_g N_A_27_55#_c_475_n 0.0119202f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_380 N_SCE_c_367_n N_A_27_55#_c_475_n 0.00331183f $X=0.75 $Y=1.69 $X2=0 $Y2=0
cc_381 SCE N_A_27_55#_c_475_n 0.0246201f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_382 N_SCE_M1016_g N_VPWR_c_2221_n 0.00673401f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_383 N_SCE_M1025_g N_VPWR_c_2221_n 0.0153739f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_384 N_SCE_M1016_g N_VPWR_c_2227_n 0.0054895f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_385 N_SCE_M1025_g N_VPWR_c_2229_n 0.00486043f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_386 N_SCE_M1016_g N_VPWR_c_2220_n 0.00648738f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_387 N_SCE_M1025_g N_VPWR_c_2220_n 0.00358042f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_388 N_SCE_c_365_n N_A_305_97#_c_2391_n 0.00444704f $X=1.45 $Y=1.015 $X2=0
+ $Y2=0
cc_389 N_SCE_M1025_g N_A_305_97#_c_2415_n 0.00141858f $X=1.16 $Y=2.775 $X2=0
+ $Y2=0
cc_390 N_SCE_M1025_g N_A_305_97#_c_2405_n 4.79243e-19 $X=1.16 $Y=2.775 $X2=0
+ $Y2=0
cc_391 N_SCE_M1016_g N_KAPWR_c_2593_n 0.00463272f $X=0.66 $Y=2.775 $X2=0 $Y2=0
cc_392 N_SCE_M1025_g N_KAPWR_c_2593_n 0.0044442f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_393 N_SCE_M1001_g N_VGND_c_2830_n 0.0128648f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_394 N_SCE_c_365_n N_VGND_c_2830_n 7.54732e-19 $X=1.45 $Y=1.015 $X2=0 $Y2=0
cc_395 N_SCE_c_366_n N_VGND_c_2830_n 0.00555605f $X=0.662 $Y=1.09 $X2=0 $Y2=0
cc_396 SCE N_VGND_c_2830_n 0.0135635f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_397 N_SCE_M1001_g N_VGND_c_2839_n 0.00452967f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_398 N_SCE_c_365_n N_VGND_c_2840_n 7.35405e-19 $X=1.45 $Y=1.015 $X2=0 $Y2=0
cc_399 N_SCE_M1001_g N_VGND_c_2845_n 0.00887478f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_400 N_SCE_M1001_g N_noxref_30_c_2991_n 0.00579352f $X=0.485 $Y=0.485 $X2=0
+ $Y2=0
cc_401 N_SCE_c_363_n N_noxref_30_c_2991_n 0.00533227f $X=1.375 $Y=1.09 $X2=0
+ $Y2=0
cc_402 N_SCE_c_365_n N_noxref_30_c_2991_n 0.00343185f $X=1.45 $Y=1.015 $X2=0
+ $Y2=0
cc_403 N_SCE_c_365_n N_noxref_30_c_2992_n 0.0114775f $X=1.45 $Y=1.015 $X2=0
+ $Y2=0
cc_404 N_SCE_M1001_g N_noxref_30_c_2993_n 4.10117e-19 $X=0.485 $Y=0.485 $X2=0
+ $Y2=0
cc_405 N_D_M1026_g N_A_27_55#_c_468_n 0.0475325f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_406 D N_A_27_55#_c_468_n 3.38944e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_407 N_D_c_421_n N_A_27_55#_c_468_n 0.00214419f $X=1.64 $Y=1.54 $X2=0 $Y2=0
cc_408 N_D_M1026_g N_A_27_55#_c_464_n 9.38065e-19 $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_409 D N_A_27_55#_c_464_n 0.00280695f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_410 N_D_c_421_n N_A_27_55#_c_464_n 0.0191672f $X=1.64 $Y=1.54 $X2=0 $Y2=0
cc_411 N_D_M1040_g N_A_27_55#_M1003_g 0.042454f $X=1.88 $Y=0.695 $X2=0 $Y2=0
cc_412 N_D_M1040_g N_A_27_55#_c_466_n 0.00942719f $X=1.88 $Y=0.695 $X2=0 $Y2=0
cc_413 N_D_M1026_g N_A_27_55#_c_474_n 8.36255e-19 $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_414 N_D_M1026_g N_A_27_55#_c_475_n 0.011465f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_415 D N_A_27_55#_c_475_n 0.0574518f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_416 N_D_c_421_n N_A_27_55#_c_475_n 0.00522383f $X=1.64 $Y=1.54 $X2=0 $Y2=0
cc_417 N_D_M1026_g N_VPWR_c_2221_n 0.00313684f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_418 N_D_M1026_g N_VPWR_c_2229_n 0.0054895f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_419 N_D_M1026_g N_VPWR_c_2220_n 0.00524789f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_420 N_D_M1040_g N_A_305_97#_c_2391_n 0.0163782f $X=1.88 $Y=0.695 $X2=0 $Y2=0
cc_421 D N_A_305_97#_c_2391_n 0.0199468f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_422 N_D_c_421_n N_A_305_97#_c_2391_n 0.00132771f $X=1.64 $Y=1.54 $X2=0 $Y2=0
cc_423 N_D_M1026_g N_A_305_97#_c_2415_n 0.00808669f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_424 N_D_M1026_g N_A_305_97#_c_2405_n 0.00473299f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_425 N_D_M1040_g N_A_305_97#_c_2392_n 0.00677786f $X=1.88 $Y=0.695 $X2=0 $Y2=0
cc_426 D N_A_305_97#_c_2392_n 0.0067051f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_427 N_D_M1040_g N_A_305_97#_c_2394_n 0.00136078f $X=1.88 $Y=0.695 $X2=0 $Y2=0
cc_428 D N_A_305_97#_c_2394_n 0.015174f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_429 N_D_M1026_g N_KAPWR_c_2593_n 0.00445017f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_430 N_D_M1040_g N_VGND_c_2840_n 7.35405e-19 $X=1.88 $Y=0.695 $X2=0 $Y2=0
cc_431 D N_noxref_30_c_2991_n 0.0162369f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_432 N_D_M1040_g N_noxref_30_c_2992_n 0.00696817f $X=1.88 $Y=0.695 $X2=0 $Y2=0
cc_433 N_A_27_55#_c_464_n N_SCD_M1022_g 0.010606f $X=2.24 $Y=1.765 $X2=0 $Y2=0
cc_434 N_A_27_55#_M1003_g N_SCD_M1022_g 0.0294313f $X=2.27 $Y=0.695 $X2=0 $Y2=0
cc_435 N_A_27_55#_c_468_n N_SCD_c_544_n 0.0201693f $X=1.98 $Y=2.275 $X2=0 $Y2=0
cc_436 N_A_27_55#_c_474_n N_SCD_c_544_n 2.51429e-19 $X=2.14 $Y=2.11 $X2=0 $Y2=0
cc_437 N_A_27_55#_c_468_n N_SCD_c_549_n 0.00661432f $X=1.98 $Y=2.275 $X2=0 $Y2=0
cc_438 N_A_27_55#_M1004_g N_SCD_c_549_n 0.0237313f $X=1.98 $Y=2.775 $X2=0 $Y2=0
cc_439 N_A_27_55#_c_464_n N_SCD_c_545_n 0.00777222f $X=2.24 $Y=1.765 $X2=0 $Y2=0
cc_440 N_A_27_55#_c_468_n N_SCD_c_546_n 0.00188289f $X=1.98 $Y=2.275 $X2=0 $Y2=0
cc_441 N_A_27_55#_c_464_n N_SCD_c_546_n 0.0068958f $X=2.24 $Y=1.765 $X2=0 $Y2=0
cc_442 N_A_27_55#_c_474_n N_SCD_c_546_n 0.0221902f $X=2.14 $Y=2.11 $X2=0 $Y2=0
cc_443 N_A_27_55#_c_472_n N_VPWR_c_2221_n 0.0293093f $X=0.445 $Y=2.755 $X2=0
+ $Y2=0
cc_444 N_A_27_55#_c_475_n N_VPWR_c_2221_n 0.0161382f $X=1.975 $Y=2.11 $X2=0
+ $Y2=0
cc_445 N_A_27_55#_M1004_g N_VPWR_c_2222_n 0.0023154f $X=1.98 $Y=2.775 $X2=0
+ $Y2=0
cc_446 N_A_27_55#_c_472_n N_VPWR_c_2227_n 0.0335644f $X=0.445 $Y=2.755 $X2=0
+ $Y2=0
cc_447 N_A_27_55#_M1004_g N_VPWR_c_2229_n 0.00424868f $X=1.98 $Y=2.775 $X2=0
+ $Y2=0
cc_448 N_A_27_55#_M1016_s N_VPWR_c_2220_n 0.00119809f $X=0.3 $Y=2.455 $X2=0
+ $Y2=0
cc_449 N_A_27_55#_M1004_g N_VPWR_c_2220_n 0.00554203f $X=1.98 $Y=2.775 $X2=0
+ $Y2=0
cc_450 N_A_27_55#_c_472_n N_VPWR_c_2220_n 0.00469612f $X=0.445 $Y=2.755 $X2=0
+ $Y2=0
cc_451 N_A_27_55#_M1003_g N_A_305_97#_c_2391_n 0.00133065f $X=2.27 $Y=0.695
+ $X2=0 $Y2=0
cc_452 N_A_27_55#_M1004_g N_A_305_97#_c_2415_n 0.0114565f $X=1.98 $Y=2.775 $X2=0
+ $Y2=0
cc_453 N_A_27_55#_c_468_n N_A_305_97#_c_2404_n 0.00646272f $X=1.98 $Y=2.275
+ $X2=0 $Y2=0
cc_454 N_A_27_55#_M1004_g N_A_305_97#_c_2404_n 0.00960371f $X=1.98 $Y=2.775
+ $X2=0 $Y2=0
cc_455 N_A_27_55#_c_474_n N_A_305_97#_c_2404_n 0.02326f $X=2.14 $Y=2.11 $X2=0
+ $Y2=0
cc_456 N_A_27_55#_c_475_n N_A_305_97#_c_2404_n 0.00157687f $X=1.975 $Y=2.11
+ $X2=0 $Y2=0
cc_457 N_A_27_55#_M1004_g N_A_305_97#_c_2405_n 0.00229015f $X=1.98 $Y=2.775
+ $X2=0 $Y2=0
cc_458 N_A_27_55#_c_475_n N_A_305_97#_c_2405_n 0.0154984f $X=1.975 $Y=2.11 $X2=0
+ $Y2=0
cc_459 N_A_27_55#_M1003_g N_A_305_97#_c_2392_n 0.00412467f $X=2.27 $Y=0.695
+ $X2=0 $Y2=0
cc_460 N_A_27_55#_c_466_n N_A_305_97#_c_2392_n 0.0011837f $X=2.255 $Y=1.365
+ $X2=0 $Y2=0
cc_461 N_A_27_55#_c_468_n N_A_305_97#_c_2393_n 4.01537e-19 $X=1.98 $Y=2.275
+ $X2=0 $Y2=0
cc_462 N_A_27_55#_c_464_n N_A_305_97#_c_2393_n 0.00619064f $X=2.24 $Y=1.765
+ $X2=0 $Y2=0
cc_463 N_A_27_55#_c_466_n N_A_305_97#_c_2393_n 0.0117004f $X=2.255 $Y=1.365
+ $X2=0 $Y2=0
cc_464 N_A_27_55#_c_474_n N_A_305_97#_c_2393_n 0.00471681f $X=2.14 $Y=2.11 $X2=0
+ $Y2=0
cc_465 N_A_27_55#_c_468_n N_A_305_97#_c_2394_n 0.00338216f $X=1.98 $Y=2.275
+ $X2=0 $Y2=0
cc_466 N_A_27_55#_c_474_n N_A_305_97#_c_2394_n 0.00629974f $X=2.14 $Y=2.11 $X2=0
+ $Y2=0
cc_467 N_A_27_55#_M1004_g N_KAPWR_c_2593_n 0.00474211f $X=1.98 $Y=2.775 $X2=0
+ $Y2=0
cc_468 N_A_27_55#_c_472_n N_KAPWR_c_2593_n 0.0556013f $X=0.445 $Y=2.755 $X2=0
+ $Y2=0
cc_469 N_A_27_55#_c_475_n N_KAPWR_c_2593_n 0.0227376f $X=1.975 $Y=2.11 $X2=0
+ $Y2=0
cc_470 N_A_27_55#_c_467_n N_VGND_c_2830_n 0.0179429f $X=0.27 $Y=0.485 $X2=0
+ $Y2=0
cc_471 N_A_27_55#_c_467_n N_VGND_c_2839_n 0.0177783f $X=0.27 $Y=0.485 $X2=0
+ $Y2=0
cc_472 N_A_27_55#_M1003_g N_VGND_c_2840_n 7.35405e-19 $X=2.27 $Y=0.695 $X2=0
+ $Y2=0
cc_473 N_A_27_55#_c_467_n N_VGND_c_2845_n 0.00964167f $X=0.27 $Y=0.485 $X2=0
+ $Y2=0
cc_474 N_A_27_55#_M1003_g N_noxref_30_c_2992_n 0.0115494f $X=2.27 $Y=0.695 $X2=0
+ $Y2=0
cc_475 N_A_27_55#_M1003_g N_noxref_30_c_2994_n 8.48223e-19 $X=2.27 $Y=0.695
+ $X2=0 $Y2=0
cc_476 N_A_27_55#_M1003_g N_noxref_32_c_3023_n 0.00166409f $X=2.27 $Y=0.695
+ $X2=0 $Y2=0
cc_477 N_SCD_M1022_g N_A_666_89#_c_1072_n 7.27045e-19 $X=2.7 $Y=0.695 $X2=0
+ $Y2=0
cc_478 N_SCD_M1052_g N_VPWR_c_2222_n 0.0123962f $X=2.62 $Y=2.775 $X2=0 $Y2=0
cc_479 N_SCD_M1052_g N_VPWR_c_2229_n 0.00362954f $X=2.62 $Y=2.775 $X2=0 $Y2=0
cc_480 N_SCD_M1052_g N_VPWR_c_2220_n 0.00388137f $X=2.62 $Y=2.775 $X2=0 $Y2=0
cc_481 N_SCD_M1052_g N_A_305_97#_c_2415_n 0.00239045f $X=2.62 $Y=2.775 $X2=0
+ $Y2=0
cc_482 N_SCD_M1052_g N_A_305_97#_c_2404_n 0.0143131f $X=2.62 $Y=2.775 $X2=0
+ $Y2=0
cc_483 N_SCD_c_549_n N_A_305_97#_c_2404_n 0.00541557f $X=2.715 $Y=2.305 $X2=0
+ $Y2=0
cc_484 N_SCD_c_546_n N_A_305_97#_c_2404_n 0.025463f $X=2.72 $Y=1.77 $X2=0 $Y2=0
cc_485 N_SCD_M1022_g N_A_305_97#_c_2393_n 0.0121532f $X=2.7 $Y=0.695 $X2=0 $Y2=0
cc_486 N_SCD_c_545_n N_A_305_97#_c_2393_n 0.00180261f $X=2.72 $Y=1.77 $X2=0
+ $Y2=0
cc_487 N_SCD_c_546_n N_A_305_97#_c_2393_n 0.026915f $X=2.72 $Y=1.77 $X2=0 $Y2=0
cc_488 N_SCD_M1052_g N_A_305_97#_c_2395_n 0.00395034f $X=2.62 $Y=2.775 $X2=0
+ $Y2=0
cc_489 N_SCD_M1022_g N_A_305_97#_c_2395_n 0.00522589f $X=2.7 $Y=0.695 $X2=0
+ $Y2=0
cc_490 N_SCD_c_545_n N_A_305_97#_c_2395_n 0.0164136f $X=2.72 $Y=1.77 $X2=0 $Y2=0
cc_491 N_SCD_c_546_n N_A_305_97#_c_2395_n 0.0500012f $X=2.72 $Y=1.77 $X2=0 $Y2=0
cc_492 N_SCD_M1052_g N_A_305_97#_c_2407_n 0.00333878f $X=2.62 $Y=2.775 $X2=0
+ $Y2=0
cc_493 N_SCD_M1052_g N_KAPWR_c_2593_n 0.00629054f $X=2.62 $Y=2.775 $X2=0 $Y2=0
cc_494 N_SCD_M1022_g N_VGND_c_2840_n 7.30329e-19 $X=2.7 $Y=0.695 $X2=0 $Y2=0
cc_495 N_SCD_M1022_g N_noxref_30_c_2992_n 0.00695764f $X=2.7 $Y=0.695 $X2=0
+ $Y2=0
cc_496 N_SCD_M1022_g N_noxref_30_c_2994_n 0.00847066f $X=2.7 $Y=0.695 $X2=0
+ $Y2=0
cc_497 N_SCD_M1022_g N_noxref_32_c_3021_n 4.37993e-19 $X=2.7 $Y=0.695 $X2=0
+ $Y2=0
cc_498 N_SCD_M1022_g N_noxref_32_c_3022_n 0.013407f $X=2.7 $Y=0.695 $X2=0 $Y2=0
cc_499 N_RESET_B_c_584_n N_A_742_63#_M1018_g 0.0212669f $X=4.32 $Y=1.145 $X2=0
+ $Y2=0
cc_500 N_RESET_B_M1049_g N_A_742_63#_M1018_g 0.0202886f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_501 N_RESET_B_M1049_g N_A_742_63#_c_781_n 0.0101003f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_502 N_RESET_B_M1049_g N_A_742_63#_M1000_g 0.0199872f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_503 N_RESET_B_c_586_n N_A_742_63#_c_767_n 0.00622075f $X=4.86 $Y=1.145 $X2=0
+ $Y2=0
cc_504 N_RESET_B_c_601_n N_A_742_63#_M1050_g 0.00431758f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_601_n N_A_742_63#_M1030_g 0.00430817f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_506 N_RESET_B_M1049_g N_A_742_63#_c_791_n 3.4555e-19 $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_507 N_RESET_B_M1011_g N_A_742_63#_c_794_n 0.0164471f $X=8.285 $Y=2.205 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_601_n N_A_742_63#_c_794_n 0.0016365f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_509 N_RESET_B_c_601_n N_A_742_63#_c_796_n 0.0173045f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_510 N_RESET_B_c_601_n N_A_742_63#_c_797_n 0.00139796f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_511 N_RESET_B_M1049_g N_A_742_63#_c_775_n 3.50857e-19 $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_512 N_RESET_B_M1049_g N_A_742_63#_c_778_n 0.00935303f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_513 N_RESET_B_c_597_n N_A_666_89#_c_1067_n 7.25259e-19 $X=6.985 $Y=1.61 $X2=0
+ $Y2=0
cc_514 N_RESET_B_c_601_n N_A_666_89#_M1015_g 0.00378029f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_515 N_RESET_B_M1049_g N_A_666_89#_c_1080_n 0.0076481f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_516 N_RESET_B_M1011_g N_A_666_89#_c_1082_n 0.00767335f $X=8.285 $Y=2.205
+ $X2=0 $Y2=0
cc_517 N_RESET_B_c_607_n N_A_666_89#_c_1082_n 0.00550332f $X=7.805 $Y=1.695
+ $X2=0 $Y2=0
cc_518 N_RESET_B_c_608_n N_A_666_89#_c_1082_n 0.00137976f $X=7.07 $Y=1.695 $X2=0
+ $Y2=0
cc_519 N_RESET_B_c_610_n N_A_666_89#_c_1082_n 0.00275732f $X=7.972 $Y=1.61 $X2=0
+ $Y2=0
cc_520 N_RESET_B_c_597_n N_A_666_89#_c_1076_n 2.12906e-19 $X=6.985 $Y=1.61 $X2=0
+ $Y2=0
cc_521 N_RESET_B_c_608_n N_A_666_89#_c_1076_n 0.00872066f $X=7.07 $Y=1.695 $X2=0
+ $Y2=0
cc_522 N_RESET_B_c_597_n N_A_1343_51#_M1010_g 0.00605633f $X=6.985 $Y=1.61 $X2=0
+ $Y2=0
cc_523 N_RESET_B_c_608_n N_A_1343_51#_M1010_g 0.00848994f $X=7.07 $Y=1.695 $X2=0
+ $Y2=0
cc_524 N_RESET_B_c_595_n N_A_1343_51#_M1035_g 0.00378728f $X=6.9 $Y=0.34 $X2=0
+ $Y2=0
cc_525 N_RESET_B_c_597_n N_A_1343_51#_M1035_g 0.00616162f $X=6.985 $Y=1.61 $X2=0
+ $Y2=0
cc_526 N_RESET_B_c_595_n N_A_1343_51#_c_1266_n 0.0146065f $X=6.9 $Y=0.34 $X2=0
+ $Y2=0
cc_527 N_RESET_B_c_597_n N_A_1343_51#_c_1266_n 0.00413113f $X=6.985 $Y=1.61
+ $X2=0 $Y2=0
cc_528 N_RESET_B_c_597_n N_A_1343_51#_c_1267_n 0.00337134f $X=6.985 $Y=1.61
+ $X2=0 $Y2=0
cc_529 N_RESET_B_M1007_g N_A_1343_51#_c_1268_n 0.00201303f $X=8.265 $Y=0.445
+ $X2=0 $Y2=0
cc_530 N_RESET_B_c_593_n N_A_1343_51#_c_1268_n 2.83785e-19 $X=8.16 $Y=1.38 $X2=0
+ $Y2=0
cc_531 N_RESET_B_c_597_n N_A_1343_51#_c_1268_n 0.0291036f $X=6.985 $Y=1.61 $X2=0
+ $Y2=0
cc_532 N_RESET_B_c_607_n N_A_1343_51#_c_1268_n 0.0249705f $X=7.805 $Y=1.695
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_598_n N_A_1343_51#_c_1268_n 0.0140029f $X=7.975 $Y=1.38 $X2=0
+ $Y2=0
cc_534 N_RESET_B_M1007_g N_A_1343_51#_c_1269_n 0.0170531f $X=8.265 $Y=0.445
+ $X2=0 $Y2=0
cc_535 N_RESET_B_c_593_n N_A_1343_51#_c_1269_n 0.00433313f $X=8.16 $Y=1.38 $X2=0
+ $Y2=0
cc_536 N_RESET_B_c_594_n N_A_1343_51#_c_1269_n 4.99796e-19 $X=8.16 $Y=1.215
+ $X2=0 $Y2=0
cc_537 N_RESET_B_c_607_n N_A_1343_51#_c_1269_n 0.00765796f $X=7.805 $Y=1.695
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_598_n N_A_1343_51#_c_1269_n 0.0262398f $X=7.975 $Y=1.38 $X2=0
+ $Y2=0
cc_539 N_RESET_B_c_597_n N_A_1343_51#_c_1270_n 0.0135839f $X=6.985 $Y=1.61 $X2=0
+ $Y2=0
cc_540 N_RESET_B_M1011_g N_A_1343_51#_c_1271_n 0.00259624f $X=8.285 $Y=2.205
+ $X2=0 $Y2=0
cc_541 N_RESET_B_M1007_g N_A_1343_51#_c_1271_n 0.00601762f $X=8.265 $Y=0.445
+ $X2=0 $Y2=0
cc_542 N_RESET_B_c_594_n N_A_1343_51#_c_1271_n 0.00502111f $X=8.16 $Y=1.215
+ $X2=0 $Y2=0
cc_543 N_RESET_B_c_598_n N_A_1343_51#_c_1271_n 0.024302f $X=7.975 $Y=1.38 $X2=0
+ $Y2=0
cc_544 N_RESET_B_c_610_n N_A_1343_51#_c_1271_n 0.00403295f $X=7.972 $Y=1.61
+ $X2=0 $Y2=0
cc_545 N_RESET_B_M1011_g N_A_1343_51#_c_1315_n 0.00714232f $X=8.285 $Y=2.205
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_610_n N_A_1343_51#_c_1315_n 0.00519791f $X=7.972 $Y=1.61
+ $X2=0 $Y2=0
cc_547 N_RESET_B_M1007_g N_A_1343_51#_c_1284_n 0.00227902f $X=8.265 $Y=0.445
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_593_n N_A_1343_51#_c_1284_n 0.0134348f $X=8.16 $Y=1.38 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_597_n N_A_1343_51#_c_1284_n 0.00996268f $X=6.985 $Y=1.61
+ $X2=0 $Y2=0
cc_550 N_RESET_B_c_607_n N_A_1343_51#_c_1284_n 0.0148746f $X=7.805 $Y=1.695
+ $X2=0 $Y2=0
cc_551 N_RESET_B_c_598_n N_A_1343_51#_c_1284_n 0.001814f $X=7.975 $Y=1.38 $X2=0
+ $Y2=0
cc_552 N_RESET_B_M1007_g N_A_1724_21#_M1027_g 0.0200812f $X=8.265 $Y=0.445 $X2=0
+ $Y2=0
cc_553 N_RESET_B_M1011_g N_A_1724_21#_M1014_g 0.0477671f $X=8.285 $Y=2.205 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_601_n N_A_1724_21#_M1014_g 0.0123562f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_601_n N_A_1724_21#_c_1496_n 0.00557408f $X=15.75 $Y=3.15
+ $X2=0 $Y2=0
cc_556 N_RESET_B_c_594_n N_A_1724_21#_c_1491_n 0.0678484f $X=8.16 $Y=1.215 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_610_n N_A_1113_419#_M1011_s 0.00266412f $X=7.972 $Y=1.61
+ $X2=0 $Y2=0
cc_558 N_RESET_B_c_601_n N_A_1113_419#_M1029_g 0.0132492f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_593_n N_A_1113_419#_c_1643_n 0.0013319f $X=8.16 $Y=1.38 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_607_n N_A_1113_419#_c_1643_n 0.0515041f $X=7.805 $Y=1.695
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_608_n N_A_1113_419#_c_1643_n 0.0122579f $X=7.07 $Y=1.695
+ $X2=0 $Y2=0
cc_562 N_RESET_B_c_610_n N_A_1113_419#_c_1643_n 0.0221933f $X=7.972 $Y=1.61
+ $X2=0 $Y2=0
cc_563 N_RESET_B_c_608_n N_A_1113_419#_c_1653_n 3.431e-19 $X=7.07 $Y=1.695 $X2=0
+ $Y2=0
cc_564 N_RESET_B_M1011_g N_A_1113_419#_c_1644_n 0.0125669f $X=8.285 $Y=2.205
+ $X2=0 $Y2=0
cc_565 N_RESET_B_c_601_n N_A_1113_419#_c_1646_n 0.00659944f $X=15.75 $Y=3.15
+ $X2=0 $Y2=0
cc_566 N_RESET_B_M1011_g N_A_1113_419#_c_1656_n 0.00313884f $X=8.285 $Y=2.205
+ $X2=0 $Y2=0
cc_567 N_RESET_B_c_601_n N_CLK_N_c_1779_n 0.00933385f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_601_n N_SLEEP_B_M1019_g 0.00934735f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_601_n N_SLEEP_B_c_1835_n 0.0168173f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_570 N_RESET_B_M1008_g N_A_2999_73#_M1051_g 0.0373581f $X=15.5 $Y=0.705 $X2=0
+ $Y2=0
cc_571 N_RESET_B_M1005_g N_A_2999_73#_M1051_g 0.00373923f $X=15.825 $Y=2.525
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_601_n N_A_2999_73#_M1031_g 0.0101105f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_573 N_RESET_B_M1005_g N_A_2999_73#_M1031_g 0.0156077f $X=15.825 $Y=2.525
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_590_n N_A_2999_73#_c_1928_n 0.00533409f $X=15.575 $Y=1.49
+ $X2=0 $Y2=0
cc_575 N_RESET_B_M1005_g N_A_2999_73#_c_1928_n 0.0130522f $X=15.825 $Y=2.525
+ $X2=0 $Y2=0
cc_576 N_RESET_B_M1005_g N_A_2999_73#_c_1929_n 0.0105803f $X=15.825 $Y=2.525
+ $X2=0 $Y2=0
cc_577 N_RESET_B_M1008_g N_A_2999_73#_c_1924_n 0.00266195f $X=15.5 $Y=0.705
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_589_n N_A_2999_73#_c_1924_n 0.00869622f $X=15.75 $Y=1.49
+ $X2=0 $Y2=0
cc_579 N_RESET_B_M1005_g N_A_2999_73#_c_1931_n 0.00519244f $X=15.825 $Y=2.525
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_590_n N_A_2999_73#_c_1932_n 0.00685224f $X=15.575 $Y=1.49
+ $X2=0 $Y2=0
cc_581 N_RESET_B_M1005_g N_A_2999_73#_c_1932_n 0.021398f $X=15.825 $Y=2.525
+ $X2=0 $Y2=0
cc_582 N_RESET_B_M1008_g N_A_2717_427#_c_1997_n 0.0366517f $X=15.5 $Y=0.705
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_589_n N_A_2717_427#_c_1999_n 0.00600628f $X=15.75 $Y=1.49
+ $X2=0 $Y2=0
cc_584 N_RESET_B_M1005_g N_A_2717_427#_M1046_g 0.0237171f $X=15.825 $Y=2.525
+ $X2=0 $Y2=0
cc_585 N_RESET_B_M1008_g N_A_2717_427#_c_2006_n 0.0015782f $X=15.5 $Y=0.705
+ $X2=0 $Y2=0
cc_586 N_RESET_B_M1008_g N_A_2717_427#_c_2007_n 0.015096f $X=15.5 $Y=0.705 $X2=0
+ $Y2=0
cc_587 N_RESET_B_c_589_n N_A_2717_427#_c_2007_n 0.00578455f $X=15.75 $Y=1.49
+ $X2=0 $Y2=0
cc_588 N_RESET_B_M1008_g N_A_2717_427#_c_2009_n 0.00615371f $X=15.5 $Y=0.705
+ $X2=0 $Y2=0
cc_589 N_RESET_B_M1008_g N_A_2717_427#_c_2011_n 4.61872e-19 $X=15.5 $Y=0.705
+ $X2=0 $Y2=0
cc_590 N_RESET_B_M1008_g N_A_2717_427#_c_2014_n 0.00323349f $X=15.5 $Y=0.705
+ $X2=0 $Y2=0
cc_591 N_RESET_B_c_589_n N_A_2717_427#_c_2014_n 0.0237171f $X=15.75 $Y=1.49
+ $X2=0 $Y2=0
cc_592 N_RESET_B_M1049_g N_VPWR_c_2223_n 0.00310437f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_601_n N_VPWR_c_2224_n 0.019904f $X=15.75 $Y=3.15 $X2=0 $Y2=0
cc_594 N_RESET_B_M1005_g N_VPWR_c_2224_n 0.00706539f $X=15.825 $Y=2.525 $X2=0
+ $Y2=0
cc_595 N_RESET_B_M1005_g N_VPWR_c_2225_n 0.00797886f $X=15.825 $Y=2.525 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_601_n N_VPWR_c_2233_n 0.00768994f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_597 N_RESET_B_c_602_n N_VPWR_c_2235_n 0.168512f $X=8.41 $Y=3.15 $X2=0 $Y2=0
cc_598 N_RESET_B_c_601_n N_VPWR_c_2220_n 0.133393f $X=15.75 $Y=3.15 $X2=0 $Y2=0
cc_599 N_RESET_B_c_602_n N_VPWR_c_2220_n 0.00778506f $X=8.41 $Y=3.15 $X2=0 $Y2=0
cc_600 N_RESET_B_M1049_g N_A_305_97#_c_2410_n 0.00216264f $X=4.585 $Y=2.415
+ $X2=0 $Y2=0
cc_601 N_RESET_B_M1049_g N_A_305_97#_c_2396_n 0.0102329f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_602 N_RESET_B_c_592_n N_A_305_97#_c_2396_n 0.00582679f $X=4.86 $Y=1.22 $X2=0
+ $Y2=0
cc_603 N_RESET_B_M1049_g N_A_305_97#_c_2398_n 0.0161754f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_604 N_RESET_B_M1049_g N_A_305_97#_c_2458_n 0.00348611f $X=4.585 $Y=2.415
+ $X2=0 $Y2=0
cc_605 N_RESET_B_M1049_g N_A_305_97#_c_2411_n 0.00689128f $X=4.585 $Y=2.415
+ $X2=0 $Y2=0
cc_606 N_RESET_B_c_592_n N_A_305_97#_c_2399_n 0.00873939f $X=4.86 $Y=1.22 $X2=0
+ $Y2=0
cc_607 N_RESET_B_M1049_g N_A_305_97#_c_2461_n 0.00990508f $X=4.585 $Y=2.415
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_592_n N_A_305_97#_c_2461_n 0.0115242f $X=4.86 $Y=1.22 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_586_n N_A_305_97#_c_2463_n 0.00337907f $X=4.86 $Y=1.145 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_586_n N_A_305_97#_c_2401_n 0.00213866f $X=4.86 $Y=1.145 $X2=0
+ $Y2=0
cc_611 N_RESET_B_M1049_g N_A_305_97#_c_2402_n 0.00203166f $X=4.585 $Y=2.415
+ $X2=0 $Y2=0
cc_612 N_RESET_B_M1049_g N_A_305_97#_c_2413_n 0.00468205f $X=4.585 $Y=2.415
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_597_n N_A_305_97#_c_2403_n 0.0315538f $X=6.985 $Y=1.61 $X2=0
+ $Y2=0
cc_614 N_RESET_B_c_601_n N_KAPWR_c_2587_n 0.0193742f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_615 N_RESET_B_c_601_n N_KAPWR_c_2588_n 0.00420304f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_616 N_RESET_B_M1005_g KAPWR 0.00730875f $X=15.825 $Y=2.525 $X2=0 $Y2=0
cc_617 N_RESET_B_M1011_g N_KAPWR_c_2590_n 0.0090303f $X=8.285 $Y=2.205 $X2=0
+ $Y2=0
cc_618 N_RESET_B_M1011_g N_KAPWR_c_2591_n 0.0142741f $X=8.285 $Y=2.205 $X2=0
+ $Y2=0
cc_619 N_RESET_B_c_601_n N_KAPWR_c_2591_n 0.0133905f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_620 N_RESET_B_M1049_g N_KAPWR_c_2593_n 0.00788983f $X=4.585 $Y=2.415 $X2=0
+ $Y2=0
cc_621 N_RESET_B_M1011_g N_KAPWR_c_2594_n 0.00815124f $X=8.285 $Y=2.205 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_601_n N_KAPWR_c_2595_n 0.0225774f $X=15.75 $Y=3.15 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_601_n N_A_2562_427#_c_2780_n 0.0450577f $X=15.75 $Y=3.15
+ $X2=0 $Y2=0
cc_624 N_RESET_B_c_601_n N_A_2562_427#_c_2781_n 0.00780634f $X=15.75 $Y=3.15
+ $X2=0 $Y2=0
cc_625 N_RESET_B_c_584_n N_VGND_c_2831_n 0.00445474f $X=4.32 $Y=1.145 $X2=0
+ $Y2=0
cc_626 N_RESET_B_c_595_n N_VGND_c_2831_n 0.00689732f $X=6.9 $Y=0.34 $X2=0 $Y2=0
cc_627 N_RESET_B_c_596_n N_VGND_c_2831_n 0.0045552f $X=4.77 $Y=0.34 $X2=0 $Y2=0
cc_628 N_RESET_B_M1007_g N_VGND_c_2832_n 0.0040248f $X=8.265 $Y=0.445 $X2=0
+ $Y2=0
cc_629 N_RESET_B_M1008_g N_VGND_c_2835_n 0.00869547f $X=15.5 $Y=0.705 $X2=0
+ $Y2=0
cc_630 N_RESET_B_c_584_n N_VGND_c_2841_n 0.00404905f $X=4.32 $Y=1.145 $X2=0
+ $Y2=0
cc_631 N_RESET_B_c_595_n N_VGND_c_2841_n 0.1586f $X=6.9 $Y=0.34 $X2=0 $Y2=0
cc_632 N_RESET_B_c_596_n N_VGND_c_2841_n 0.00659816f $X=4.77 $Y=0.34 $X2=0 $Y2=0
cc_633 N_RESET_B_M1008_g N_VGND_c_2843_n 0.00407914f $X=15.5 $Y=0.705 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_584_n N_VGND_c_2845_n 0.00472204f $X=4.32 $Y=1.145 $X2=0
+ $Y2=0
cc_635 N_RESET_B_M1007_g N_VGND_c_2845_n 0.00709767f $X=8.265 $Y=0.445 $X2=0
+ $Y2=0
cc_636 N_RESET_B_M1008_g N_VGND_c_2845_n 0.00425776f $X=15.5 $Y=0.705 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_595_n N_VGND_c_2845_n 0.0913057f $X=6.9 $Y=0.34 $X2=0 $Y2=0
cc_638 N_RESET_B_c_596_n N_VGND_c_2845_n 0.0104196f $X=4.77 $Y=0.34 $X2=0 $Y2=0
cc_639 N_RESET_B_M1007_g N_VGND_c_2848_n 0.00749764f $X=8.265 $Y=0.445 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_584_n N_noxref_32_c_3022_n 0.0132915f $X=4.32 $Y=1.145 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_584_n N_noxref_32_c_3024_n 0.00833495f $X=4.32 $Y=1.145 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_586_n N_noxref_32_c_3024_n 0.00858726f $X=4.86 $Y=1.145 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_592_n N_noxref_32_c_3024_n 0.00592695f $X=4.86 $Y=1.22 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_595_n N_noxref_32_c_3024_n 0.00689632f $X=6.9 $Y=0.34 $X2=0
+ $Y2=0
cc_645 N_RESET_B_c_596_n N_noxref_32_c_3024_n 0.00123572f $X=4.77 $Y=0.34 $X2=0
+ $Y2=0
cc_646 N_RESET_B_c_595_n N_A_1009_107#_M1012_s 0.0027844f $X=6.9 $Y=0.34 $X2=0
+ $Y2=0
cc_647 N_RESET_B_c_586_n N_A_1009_107#_c_3056_n 0.00420455f $X=4.86 $Y=1.145
+ $X2=0 $Y2=0
cc_648 N_RESET_B_c_595_n N_A_1009_107#_c_3056_n 0.116433f $X=6.9 $Y=0.34 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_597_n A_1373_77# 0.00164114f $X=6.985 $Y=1.61 $X2=-0.19
+ $Y2=-0.245
cc_650 N_RESET_B_M1007_g N_A_1453_77#_c_3075_n 0.0105795f $X=8.265 $Y=0.445
+ $X2=0 $Y2=0
cc_651 N_RESET_B_M1007_g N_A_1453_77#_c_3076_n 0.00430107f $X=8.265 $Y=0.445
+ $X2=0 $Y2=0
cc_652 N_RESET_B_c_595_n N_A_1453_77#_c_3076_n 0.00314781f $X=6.9 $Y=0.34 $X2=0
+ $Y2=0
cc_653 N_RESET_B_M1007_g N_A_1453_77#_c_3077_n 0.0108788f $X=8.265 $Y=0.445
+ $X2=0 $Y2=0
cc_654 N_A_742_63#_c_767_n N_A_666_89#_c_1066_n 0.0108692f $X=5.5 $Y=1.605 $X2=0
+ $Y2=0
cc_655 N_A_742_63#_M1037_g N_A_666_89#_M1053_g 0.0330693f $X=5.49 $Y=2.305 $X2=0
+ $Y2=0
cc_656 N_A_742_63#_c_791_n N_A_666_89#_M1053_g 2.29953e-19 $X=5.295 $Y=2.905
+ $X2=0 $Y2=0
cc_657 N_A_742_63#_c_792_n N_A_666_89#_M1053_g 0.015459f $X=7.075 $Y=2.99 $X2=0
+ $Y2=0
cc_658 N_A_742_63#_c_769_n N_A_666_89#_c_1068_n 0.00425451f $X=13.51 $Y=1.405
+ $X2=0 $Y2=0
cc_659 N_A_742_63#_c_771_n N_A_666_89#_c_1068_n 0.00277848f $X=13.74 $Y=1.1
+ $X2=0 $Y2=0
cc_660 N_A_742_63#_c_772_n N_A_666_89#_c_1068_n 0.0118167f $X=13.51 $Y=1.48
+ $X2=0 $Y2=0
cc_661 N_A_742_63#_M1030_g N_A_666_89#_M1015_g 0.0118167f $X=13.51 $Y=2.345
+ $X2=0 $Y2=0
cc_662 N_A_742_63#_c_770_n N_A_666_89#_M1013_g 0.0138207f $X=13.74 $Y=1.025
+ $X2=0 $Y2=0
cc_663 N_A_742_63#_M1018_g N_A_666_89#_c_1072_n 0.0208711f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_664 N_A_742_63#_M1018_g N_A_666_89#_c_1080_n 0.0110317f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_665 N_A_742_63#_M1000_g N_A_666_89#_c_1080_n 0.00913564f $X=5.13 $Y=2.305
+ $X2=0 $Y2=0
cc_666 N_A_742_63#_M1037_g N_A_666_89#_c_1080_n 0.0115018f $X=5.49 $Y=2.305
+ $X2=0 $Y2=0
cc_667 N_A_742_63#_c_791_n N_A_666_89#_c_1080_n 0.0187682f $X=5.295 $Y=2.905
+ $X2=0 $Y2=0
cc_668 N_A_742_63#_c_775_n N_A_666_89#_c_1080_n 0.007751f $X=5.215 $Y=1.77 $X2=0
+ $Y2=0
cc_669 N_A_742_63#_M1018_g N_A_666_89#_c_1081_n 0.00142008f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_670 N_A_742_63#_M1050_g N_A_666_89#_c_1082_n 0.00601177f $X=13.15 $Y=2.345
+ $X2=0 $Y2=0
cc_671 N_A_742_63#_M1030_g N_A_666_89#_c_1082_n 0.0115226f $X=13.51 $Y=2.345
+ $X2=0 $Y2=0
cc_672 N_A_742_63#_c_794_n N_A_666_89#_c_1082_n 0.0132002f $X=9.41 $Y=2.435
+ $X2=0 $Y2=0
cc_673 N_A_742_63#_c_842_p N_A_666_89#_c_1082_n 0.00122109f $X=7.245 $Y=2.435
+ $X2=0 $Y2=0
cc_674 N_A_742_63#_c_799_n N_A_666_89#_c_1082_n 0.012822f $X=10.855 $Y=2.095
+ $X2=0 $Y2=0
cc_675 N_A_742_63#_c_800_n N_A_666_89#_c_1082_n 0.0123261f $X=10.675 $Y=2.095
+ $X2=0 $Y2=0
cc_676 N_A_742_63#_c_774_n N_A_666_89#_c_1082_n 0.0115699f $X=10.94 $Y=2.01
+ $X2=0 $Y2=0
cc_677 N_A_742_63#_c_803_n N_A_666_89#_c_1082_n 0.0461197f $X=11.91 $Y=2.035
+ $X2=0 $Y2=0
cc_678 N_A_742_63#_c_804_n N_A_666_89#_c_1082_n 0.0364553f $X=11.445 $Y=2.035
+ $X2=0 $Y2=0
cc_679 N_A_742_63#_c_776_n N_A_666_89#_c_1082_n 0.00262818f $X=12.98 $Y=1.57
+ $X2=0 $Y2=0
cc_680 N_A_742_63#_c_777_n N_A_666_89#_c_1082_n 0.00738198f $X=12.75 $Y=1.555
+ $X2=0 $Y2=0
cc_681 N_A_742_63#_M1018_g N_A_666_89#_c_1074_n 0.0306805f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_682 N_A_742_63#_c_778_n N_A_666_89#_c_1075_n 0.0162069f $X=5.5 $Y=1.77 $X2=0
+ $Y2=0
cc_683 N_A_742_63#_c_792_n N_A_1343_51#_M1010_g 0.0169103f $X=7.075 $Y=2.99
+ $X2=0 $Y2=0
cc_684 N_A_742_63#_c_853_p N_A_1343_51#_M1010_g 0.0133194f $X=7.16 $Y=2.905
+ $X2=0 $Y2=0
cc_685 N_A_742_63#_c_842_p N_A_1343_51#_M1010_g 0.00475869f $X=7.245 $Y=2.435
+ $X2=0 $Y2=0
cc_686 N_A_742_63#_c_770_n N_A_1343_51#_c_1279_n 0.0105825f $X=13.74 $Y=1.025
+ $X2=0 $Y2=0
cc_687 N_A_742_63#_c_771_n N_A_1343_51#_c_1283_n 0.00504675f $X=13.74 $Y=1.1
+ $X2=0 $Y2=0
cc_688 N_A_742_63#_c_794_n N_A_1724_21#_M1014_g 0.0147138f $X=9.41 $Y=2.435
+ $X2=0 $Y2=0
cc_689 N_A_742_63#_c_795_n N_A_1724_21#_M1014_g 9.13735e-19 $X=9.495 $Y=2.725
+ $X2=0 $Y2=0
cc_690 N_A_742_63#_c_773_n N_A_1724_21#_c_1481_n 0.00385328f $X=10.855 $Y=1.1
+ $X2=0 $Y2=0
cc_691 N_A_742_63#_c_774_n N_A_1724_21#_c_1481_n 0.0035088f $X=10.94 $Y=2.01
+ $X2=0 $Y2=0
cc_692 N_A_742_63#_c_773_n N_A_1724_21#_c_1482_n 0.0197451f $X=10.855 $Y=1.1
+ $X2=0 $Y2=0
cc_693 N_A_742_63#_M1038_s N_A_1724_21#_c_1483_n 0.00918457f $X=10.44 $Y=0.485
+ $X2=0 $Y2=0
cc_694 N_A_742_63#_c_773_n N_A_1724_21#_c_1483_n 0.0432029f $X=10.855 $Y=1.1
+ $X2=0 $Y2=0
cc_695 N_A_742_63#_c_773_n N_A_1724_21#_c_1485_n 0.00163541f $X=10.855 $Y=1.1
+ $X2=0 $Y2=0
cc_696 N_A_742_63#_c_865_p N_A_1724_21#_c_1486_n 0.00950132f $X=12.08 $Y=1.46
+ $X2=0 $Y2=0
cc_697 N_A_742_63#_c_777_n N_A_1724_21#_c_1486_n 0.0359284f $X=12.75 $Y=1.555
+ $X2=0 $Y2=0
cc_698 N_A_742_63#_c_773_n N_A_1724_21#_c_1487_n 0.0157846f $X=10.855 $Y=1.1
+ $X2=0 $Y2=0
cc_699 N_A_742_63#_M1050_g N_A_1724_21#_c_1495_n 0.0044803f $X=13.15 $Y=2.345
+ $X2=0 $Y2=0
cc_700 N_A_742_63#_c_803_n N_A_1724_21#_c_1495_n 0.00858679f $X=11.91 $Y=2.035
+ $X2=0 $Y2=0
cc_701 N_A_742_63#_c_805_n N_A_1724_21#_c_1495_n 0.0170333f $X=11.995 $Y=1.95
+ $X2=0 $Y2=0
cc_702 N_A_742_63#_c_776_n N_A_1724_21#_c_1495_n 0.00161853f $X=12.98 $Y=1.57
+ $X2=0 $Y2=0
cc_703 N_A_742_63#_c_777_n N_A_1724_21#_c_1495_n 0.0265194f $X=12.75 $Y=1.555
+ $X2=0 $Y2=0
cc_704 N_A_742_63#_M1050_g N_A_1724_21#_c_1496_n 0.0047852f $X=13.15 $Y=2.345
+ $X2=0 $Y2=0
cc_705 N_A_742_63#_c_803_n N_A_1724_21#_c_1496_n 0.00314096f $X=11.91 $Y=2.035
+ $X2=0 $Y2=0
cc_706 N_A_742_63#_M1050_g N_A_1724_21#_c_1497_n 0.0153748f $X=13.15 $Y=2.345
+ $X2=0 $Y2=0
cc_707 N_A_742_63#_M1030_g N_A_1724_21#_c_1497_n 0.00436029f $X=13.51 $Y=2.345
+ $X2=0 $Y2=0
cc_708 N_A_742_63#_c_776_n N_A_1724_21#_c_1497_n 0.027362f $X=12.98 $Y=1.57
+ $X2=0 $Y2=0
cc_709 N_A_742_63#_c_777_n N_A_1724_21#_c_1497_n 0.00634566f $X=12.75 $Y=1.555
+ $X2=0 $Y2=0
cc_710 N_A_742_63#_c_779_n N_A_1724_21#_c_1497_n 0.00582934f $X=13.02 $Y=1.48
+ $X2=0 $Y2=0
cc_711 N_A_742_63#_c_770_n N_A_1724_21#_c_1488_n 0.00499804f $X=13.74 $Y=1.025
+ $X2=0 $Y2=0
cc_712 N_A_742_63#_c_770_n N_A_1724_21#_c_1489_n 5.5335e-19 $X=13.74 $Y=1.025
+ $X2=0 $Y2=0
cc_713 N_A_742_63#_c_771_n N_A_1724_21#_c_1489_n 0.00472408f $X=13.74 $Y=1.1
+ $X2=0 $Y2=0
cc_714 N_A_742_63#_c_776_n N_A_1724_21#_c_1489_n 0.00302183f $X=12.98 $Y=1.57
+ $X2=0 $Y2=0
cc_715 N_A_742_63#_c_779_n N_A_1724_21#_c_1489_n 0.00653368f $X=13.02 $Y=1.48
+ $X2=0 $Y2=0
cc_716 N_A_742_63#_c_768_n N_A_1724_21#_c_1490_n 0.00697312f $X=13.435 $Y=1.48
+ $X2=0 $Y2=0
cc_717 N_A_742_63#_c_769_n N_A_1724_21#_c_1490_n 0.00657496f $X=13.51 $Y=1.405
+ $X2=0 $Y2=0
cc_718 N_A_742_63#_M1030_g N_A_1724_21#_c_1490_n 0.00588428f $X=13.51 $Y=2.345
+ $X2=0 $Y2=0
cc_719 N_A_742_63#_c_771_n N_A_1724_21#_c_1490_n 0.00153336f $X=13.74 $Y=1.1
+ $X2=0 $Y2=0
cc_720 N_A_742_63#_c_772_n N_A_1724_21#_c_1490_n 0.00180745f $X=13.51 $Y=1.48
+ $X2=0 $Y2=0
cc_721 N_A_742_63#_c_776_n N_A_1724_21#_c_1490_n 0.0275473f $X=12.98 $Y=1.57
+ $X2=0 $Y2=0
cc_722 N_A_742_63#_c_779_n N_A_1724_21#_c_1490_n 0.00487092f $X=13.02 $Y=1.48
+ $X2=0 $Y2=0
cc_723 N_A_742_63#_c_776_n N_A_1724_21#_c_1493_n 0.0218734f $X=12.98 $Y=1.57
+ $X2=0 $Y2=0
cc_724 N_A_742_63#_c_779_n N_A_1724_21#_c_1493_n 0.00191505f $X=13.02 $Y=1.48
+ $X2=0 $Y2=0
cc_725 N_A_742_63#_c_792_n N_A_1113_419#_M1037_d 0.00354099f $X=7.075 $Y=2.99
+ $X2=0 $Y2=0
cc_726 N_A_742_63#_c_794_n N_A_1113_419#_M1011_s 0.00505428f $X=9.41 $Y=2.435
+ $X2=0 $Y2=0
cc_727 N_A_742_63#_c_794_n N_A_1113_419#_M1029_g 0.0118871f $X=9.41 $Y=2.435
+ $X2=0 $Y2=0
cc_728 N_A_742_63#_c_795_n N_A_1113_419#_M1029_g 0.00846735f $X=9.495 $Y=2.725
+ $X2=0 $Y2=0
cc_729 N_A_742_63#_c_797_n N_A_1113_419#_M1029_g 0.00525093f $X=9.58 $Y=2.81
+ $X2=0 $Y2=0
cc_730 N_A_742_63#_c_773_n N_A_1113_419#_c_1637_n 0.00144168f $X=10.855 $Y=1.1
+ $X2=0 $Y2=0
cc_731 N_A_742_63#_c_798_n N_A_1113_419#_c_1639_n 2.11433e-19 $X=10.59 $Y=2.725
+ $X2=0 $Y2=0
cc_732 N_A_742_63#_c_800_n N_A_1113_419#_c_1639_n 7.9343e-19 $X=10.675 $Y=2.095
+ $X2=0 $Y2=0
cc_733 N_A_742_63#_M1037_g N_A_1113_419#_c_1642_n 0.0101313f $X=5.49 $Y=2.305
+ $X2=0 $Y2=0
cc_734 N_A_742_63#_c_791_n N_A_1113_419#_c_1642_n 0.024553f $X=5.295 $Y=2.905
+ $X2=0 $Y2=0
cc_735 N_A_742_63#_c_792_n N_A_1113_419#_c_1642_n 0.0286898f $X=7.075 $Y=2.99
+ $X2=0 $Y2=0
cc_736 N_A_742_63#_M1037_g N_A_1113_419#_c_1668_n 0.00933555f $X=5.49 $Y=2.305
+ $X2=0 $Y2=0
cc_737 N_A_742_63#_c_767_n N_A_1113_419#_c_1668_n 0.0108519f $X=5.5 $Y=1.605
+ $X2=0 $Y2=0
cc_738 N_A_742_63#_c_775_n N_A_1113_419#_c_1668_n 0.0452248f $X=5.215 $Y=1.77
+ $X2=0 $Y2=0
cc_739 N_A_742_63#_c_778_n N_A_1113_419#_c_1668_n 0.0102249f $X=5.5 $Y=1.77
+ $X2=0 $Y2=0
cc_740 N_A_742_63#_c_792_n N_A_1113_419#_c_1672_n 0.0176867f $X=7.075 $Y=2.99
+ $X2=0 $Y2=0
cc_741 N_A_742_63#_c_842_p N_A_1113_419#_c_1672_n 0.0122365f $X=7.245 $Y=2.435
+ $X2=0 $Y2=0
cc_742 N_A_742_63#_c_794_n N_A_1113_419#_c_1643_n 0.119963f $X=9.41 $Y=2.435
+ $X2=0 $Y2=0
cc_743 N_A_742_63#_c_842_p N_A_1113_419#_c_1643_n 0.0124504f $X=7.245 $Y=2.435
+ $X2=0 $Y2=0
cc_744 N_A_742_63#_c_794_n N_A_1113_419#_c_1644_n 0.0098878f $X=9.41 $Y=2.435
+ $X2=0 $Y2=0
cc_745 N_A_742_63#_c_796_n N_A_1113_419#_c_1644_n 0.00887562f $X=10.505 $Y=2.81
+ $X2=0 $Y2=0
cc_746 N_A_742_63#_c_800_n N_A_1113_419#_c_1644_n 0.0141113f $X=10.675 $Y=2.095
+ $X2=0 $Y2=0
cc_747 N_A_742_63#_c_796_n N_A_1113_419#_c_1645_n 0.0171718f $X=10.505 $Y=2.81
+ $X2=0 $Y2=0
cc_748 N_A_742_63#_c_798_n N_A_1113_419#_c_1645_n 0.0277379f $X=10.59 $Y=2.725
+ $X2=0 $Y2=0
cc_749 N_A_742_63#_c_796_n N_A_1113_419#_c_1646_n 0.00351548f $X=10.505 $Y=2.81
+ $X2=0 $Y2=0
cc_750 N_A_742_63#_c_798_n N_A_1113_419#_c_1646_n 0.00411566f $X=10.59 $Y=2.725
+ $X2=0 $Y2=0
cc_751 N_A_742_63#_c_773_n N_CLK_N_M1038_g 0.0145164f $X=10.855 $Y=1.1 $X2=0
+ $Y2=0
cc_752 N_A_742_63#_c_774_n N_CLK_N_M1038_g 0.0114024f $X=10.94 $Y=2.01 $X2=0
+ $Y2=0
cc_753 N_A_742_63#_c_798_n N_CLK_N_c_1779_n 0.00234905f $X=10.59 $Y=2.725 $X2=0
+ $Y2=0
cc_754 N_A_742_63#_c_774_n N_CLK_N_c_1779_n 0.0254565f $X=10.94 $Y=2.01 $X2=0
+ $Y2=0
cc_755 N_A_742_63#_c_802_n N_CLK_N_c_1779_n 0.00884018f $X=11.36 $Y=2.405 $X2=0
+ $Y2=0
cc_756 N_A_742_63#_c_804_n N_CLK_N_c_1779_n 0.016451f $X=11.445 $Y=2.035 $X2=0
+ $Y2=0
cc_757 N_A_742_63#_c_773_n N_CLK_N_c_1780_n 0.0119805f $X=10.855 $Y=1.1 $X2=0
+ $Y2=0
cc_758 N_A_742_63#_c_799_n N_CLK_N_c_1780_n 0.00658177f $X=10.855 $Y=2.095 $X2=0
+ $Y2=0
cc_759 N_A_742_63#_c_800_n N_CLK_N_c_1780_n 0.00391179f $X=10.675 $Y=2.095 $X2=0
+ $Y2=0
cc_760 N_A_742_63#_c_773_n N_CLK_N_c_1781_n 0.0139537f $X=10.855 $Y=1.1 $X2=0
+ $Y2=0
cc_761 N_A_742_63#_c_799_n N_CLK_N_c_1781_n 6.09209e-19 $X=10.855 $Y=2.095 $X2=0
+ $Y2=0
cc_762 N_A_742_63#_c_800_n N_CLK_N_c_1781_n 0.0112962f $X=10.675 $Y=2.095 $X2=0
+ $Y2=0
cc_763 N_A_742_63#_c_774_n N_CLK_N_c_1781_n 0.0209422f $X=10.94 $Y=2.01 $X2=0
+ $Y2=0
cc_764 N_A_742_63#_c_773_n N_SLEEP_B_c_1826_n 6.56102e-19 $X=10.855 $Y=1.1
+ $X2=-0.19 $Y2=-0.245
cc_765 N_A_742_63#_c_774_n N_SLEEP_B_M1019_g 0.00169115f $X=10.94 $Y=2.01 $X2=0
+ $Y2=0
cc_766 N_A_742_63#_c_802_n N_SLEEP_B_M1019_g 7.45316e-19 $X=11.36 $Y=2.405 $X2=0
+ $Y2=0
cc_767 N_A_742_63#_c_803_n N_SLEEP_B_M1019_g 0.0150711f $X=11.91 $Y=2.035 $X2=0
+ $Y2=0
cc_768 N_A_742_63#_c_805_n N_SLEEP_B_M1019_g 0.00438947f $X=11.995 $Y=1.95 $X2=0
+ $Y2=0
cc_769 N_A_742_63#_c_803_n N_SLEEP_B_c_1835_n 0.00607149f $X=11.91 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_A_742_63#_c_805_n N_SLEEP_B_c_1835_n 0.00951161f $X=11.995 $Y=1.95
+ $X2=0 $Y2=0
cc_771 N_A_742_63#_c_771_n N_SLEEP_B_c_1830_n 0.0017449f $X=13.74 $Y=1.1 $X2=0
+ $Y2=0
cc_772 N_A_742_63#_c_776_n N_SLEEP_B_c_1830_n 0.00648042f $X=12.98 $Y=1.57 $X2=0
+ $Y2=0
cc_773 N_A_742_63#_c_773_n N_SLEEP_B_c_1831_n 0.00368018f $X=10.855 $Y=1.1 $X2=0
+ $Y2=0
cc_774 N_A_742_63#_c_774_n N_SLEEP_B_c_1831_n 0.00151126f $X=10.94 $Y=2.01 $X2=0
+ $Y2=0
cc_775 N_A_742_63#_c_803_n N_SLEEP_B_c_1831_n 0.00616665f $X=11.91 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_A_742_63#_c_804_n N_SLEEP_B_c_1831_n 0.00116113f $X=11.445 $Y=2.035
+ $X2=0 $Y2=0
cc_777 N_A_742_63#_c_805_n N_SLEEP_B_c_1831_n 0.00510513f $X=11.995 $Y=1.95
+ $X2=0 $Y2=0
cc_778 N_A_742_63#_c_865_p N_SLEEP_B_c_1831_n 0.00942043f $X=12.08 $Y=1.46 $X2=0
+ $Y2=0
cc_779 N_A_742_63#_c_776_n N_SLEEP_B_c_1831_n 0.00160484f $X=12.98 $Y=1.57 $X2=0
+ $Y2=0
cc_780 N_A_742_63#_c_777_n N_SLEEP_B_c_1831_n 0.0199428f $X=12.75 $Y=1.555 $X2=0
+ $Y2=0
cc_781 N_A_742_63#_c_779_n N_SLEEP_B_c_1831_n 0.00578733f $X=13.02 $Y=1.48 $X2=0
+ $Y2=0
cc_782 N_A_742_63#_c_774_n N_SLEEP_B_c_1833_n 0.0387523f $X=10.94 $Y=2.01 $X2=0
+ $Y2=0
cc_783 N_A_742_63#_c_803_n N_SLEEP_B_c_1833_n 0.00797561f $X=11.91 $Y=2.035
+ $X2=0 $Y2=0
cc_784 N_A_742_63#_c_804_n N_SLEEP_B_c_1833_n 0.0206428f $X=11.445 $Y=2.035
+ $X2=0 $Y2=0
cc_785 N_A_742_63#_c_805_n N_SLEEP_B_c_1833_n 0.00996665f $X=11.995 $Y=1.95
+ $X2=0 $Y2=0
cc_786 N_A_742_63#_c_865_p N_SLEEP_B_c_1833_n 0.00764136f $X=12.08 $Y=1.46 $X2=0
+ $Y2=0
cc_787 N_A_742_63#_c_770_n N_A_2717_427#_c_2004_n 0.00854431f $X=13.74 $Y=1.025
+ $X2=0 $Y2=0
cc_788 N_A_742_63#_c_769_n N_A_2717_427#_c_2005_n 0.016425f $X=13.51 $Y=1.405
+ $X2=0 $Y2=0
cc_789 N_A_742_63#_c_770_n N_A_2717_427#_c_2005_n 0.00250863f $X=13.74 $Y=1.025
+ $X2=0 $Y2=0
cc_790 N_A_742_63#_c_771_n N_A_2717_427#_c_2005_n 0.0096103f $X=13.74 $Y=1.1
+ $X2=0 $Y2=0
cc_791 N_A_742_63#_M1030_g N_A_2717_427#_c_2022_n 0.0018396f $X=13.51 $Y=2.345
+ $X2=0 $Y2=0
cc_792 N_A_742_63#_M1018_g N_VPWR_c_2223_n 0.00167339f $X=3.785 $Y=0.655 $X2=0
+ $Y2=0
cc_793 N_A_742_63#_c_781_n N_VPWR_c_2223_n 0.0169604f $X=5.055 $Y=3.15 $X2=0
+ $Y2=0
cc_794 N_A_742_63#_M1000_g N_VPWR_c_2223_n 0.00430004f $X=5.13 $Y=2.305 $X2=0
+ $Y2=0
cc_795 N_A_742_63#_c_782_n N_VPWR_c_2231_n 0.0150071f $X=3.86 $Y=3.15 $X2=0
+ $Y2=0
cc_796 N_A_742_63#_c_781_n N_VPWR_c_2235_n 0.03213f $X=5.055 $Y=3.15 $X2=0 $Y2=0
cc_797 N_A_742_63#_c_792_n N_VPWR_c_2235_n 0.111853f $X=7.075 $Y=2.99 $X2=0
+ $Y2=0
cc_798 N_A_742_63#_c_793_n N_VPWR_c_2235_n 0.0115893f $X=5.38 $Y=2.99 $X2=0
+ $Y2=0
cc_799 N_A_742_63#_c_796_n N_VPWR_c_2235_n 0.0376753f $X=10.505 $Y=2.81 $X2=0
+ $Y2=0
cc_800 N_A_742_63#_c_797_n N_VPWR_c_2235_n 0.00595471f $X=9.58 $Y=2.81 $X2=0
+ $Y2=0
cc_801 N_A_742_63#_c_781_n N_VPWR_c_2220_n 0.0190823f $X=5.055 $Y=3.15 $X2=0
+ $Y2=0
cc_802 N_A_742_63#_c_782_n N_VPWR_c_2220_n 0.00544415f $X=3.86 $Y=3.15 $X2=0
+ $Y2=0
cc_803 N_A_742_63#_c_784_n N_VPWR_c_2220_n 0.00848318f $X=5.415 $Y=3.15 $X2=0
+ $Y2=0
cc_804 N_A_742_63#_c_789_n N_VPWR_c_2220_n 0.00367996f $X=5.13 $Y=3.15 $X2=0
+ $Y2=0
cc_805 N_A_742_63#_c_792_n N_VPWR_c_2220_n 0.0146878f $X=7.075 $Y=2.99 $X2=0
+ $Y2=0
cc_806 N_A_742_63#_c_793_n N_VPWR_c_2220_n 0.00141402f $X=5.38 $Y=2.99 $X2=0
+ $Y2=0
cc_807 N_A_742_63#_c_796_n N_VPWR_c_2220_n 0.0038467f $X=10.505 $Y=2.81 $X2=0
+ $Y2=0
cc_808 N_A_742_63#_c_797_n N_VPWR_c_2220_n 5.96303e-19 $X=9.58 $Y=2.81 $X2=0
+ $Y2=0
cc_809 N_A_742_63#_M1018_g N_A_305_97#_c_2393_n 6.77363e-19 $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_810 N_A_742_63#_M1018_g N_A_305_97#_c_2395_n 0.0035825f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_811 N_A_742_63#_M1018_g N_A_305_97#_c_2407_n 0.00327479f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_812 N_A_742_63#_M1018_g N_A_305_97#_c_2408_n 0.0140623f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_813 N_A_742_63#_c_781_n N_A_305_97#_c_2408_n 0.00543107f $X=5.055 $Y=3.15
+ $X2=0 $Y2=0
cc_814 N_A_742_63#_M1018_g N_A_305_97#_c_2410_n 0.0130144f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_815 N_A_742_63#_M1018_g N_A_305_97#_c_2397_n 0.0020967f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_816 N_A_742_63#_c_767_n N_A_305_97#_c_2398_n 0.00363022f $X=5.5 $Y=1.605
+ $X2=0 $Y2=0
cc_817 N_A_742_63#_c_775_n N_A_305_97#_c_2398_n 0.00740486f $X=5.215 $Y=1.77
+ $X2=0 $Y2=0
cc_818 N_A_742_63#_c_778_n N_A_305_97#_c_2398_n 0.0010121f $X=5.5 $Y=1.77 $X2=0
+ $Y2=0
cc_819 N_A_742_63#_M1000_g N_A_305_97#_c_2458_n 0.00600217f $X=5.13 $Y=2.305
+ $X2=0 $Y2=0
cc_820 N_A_742_63#_c_791_n N_A_305_97#_c_2458_n 0.0262999f $X=5.295 $Y=2.905
+ $X2=0 $Y2=0
cc_821 N_A_742_63#_c_781_n N_A_305_97#_c_2411_n 0.00556695f $X=5.055 $Y=3.15
+ $X2=0 $Y2=0
cc_822 N_A_742_63#_c_775_n N_A_305_97#_c_2399_n 0.0249444f $X=5.215 $Y=1.77
+ $X2=0 $Y2=0
cc_823 N_A_742_63#_c_778_n N_A_305_97#_c_2399_n 0.002357f $X=5.5 $Y=1.77 $X2=0
+ $Y2=0
cc_824 N_A_742_63#_c_767_n N_A_305_97#_c_2400_n 0.0141389f $X=5.5 $Y=1.605 $X2=0
+ $Y2=0
cc_825 N_A_742_63#_M1018_g N_A_305_97#_c_2412_n 4.37323e-19 $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_826 N_A_742_63#_c_775_n N_A_305_97#_c_2402_n 0.0109141f $X=5.215 $Y=1.77
+ $X2=0 $Y2=0
cc_827 N_A_742_63#_c_778_n N_A_305_97#_c_2402_n 0.00150476f $X=5.5 $Y=1.77 $X2=0
+ $Y2=0
cc_828 N_A_742_63#_M1000_g N_A_305_97#_c_2413_n 0.00113268f $X=5.13 $Y=2.305
+ $X2=0 $Y2=0
cc_829 N_A_742_63#_c_791_n N_A_305_97#_c_2413_n 0.00518663f $X=5.295 $Y=2.905
+ $X2=0 $Y2=0
cc_830 N_A_742_63#_c_775_n N_A_305_97#_c_2413_n 0.00168638f $X=5.215 $Y=1.77
+ $X2=0 $Y2=0
cc_831 N_A_742_63#_c_778_n N_A_305_97#_c_2413_n 2.31524e-19 $X=5.5 $Y=1.77 $X2=0
+ $Y2=0
cc_832 N_A_742_63#_c_791_n A_1041_419# 0.00212545f $X=5.295 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_833 N_A_742_63#_c_792_n A_1242_419# 0.00923461f $X=7.075 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_834 N_A_742_63#_c_792_n N_KAPWR_M1010_d 0.00523469f $X=7.075 $Y=2.99
+ $X2=-0.19 $Y2=-0.245
cc_835 N_A_742_63#_c_853_p N_KAPWR_M1010_d 0.0151934f $X=7.16 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_836 N_A_742_63#_c_794_n N_KAPWR_M1010_d 0.0114548f $X=9.41 $Y=2.435 $X2=-0.19
+ $Y2=-0.245
cc_837 N_A_742_63#_c_842_p N_KAPWR_M1010_d 0.0048087f $X=7.245 $Y=2.435
+ $X2=-0.19 $Y2=-0.245
cc_838 N_A_742_63#_c_794_n N_KAPWR_M1014_d 0.00676128f $X=9.41 $Y=2.435 $X2=0
+ $Y2=0
cc_839 N_A_742_63#_c_799_n N_KAPWR_M1042_s 0.00125621f $X=10.855 $Y=2.095 $X2=0
+ $Y2=0
cc_840 N_A_742_63#_c_804_n N_KAPWR_M1042_s 0.00173711f $X=11.445 $Y=2.035 $X2=0
+ $Y2=0
cc_841 N_A_742_63#_c_803_n N_KAPWR_M1019_d 0.00478541f $X=11.91 $Y=2.035 $X2=0
+ $Y2=0
cc_842 N_A_742_63#_c_805_n N_KAPWR_M1019_d 0.00262563f $X=11.995 $Y=1.95 $X2=0
+ $Y2=0
cc_843 N_A_742_63#_c_796_n N_KAPWR_c_2586_n 0.0123245f $X=10.505 $Y=2.81 $X2=0
+ $Y2=0
cc_844 N_A_742_63#_c_798_n N_KAPWR_c_2586_n 0.0274894f $X=10.59 $Y=2.725 $X2=0
+ $Y2=0
cc_845 N_A_742_63#_c_799_n N_KAPWR_c_2586_n 6.11119e-19 $X=10.855 $Y=2.095 $X2=0
+ $Y2=0
cc_846 N_A_742_63#_c_802_n N_KAPWR_c_2586_n 0.0139955f $X=11.36 $Y=2.405 $X2=0
+ $Y2=0
cc_847 N_A_742_63#_c_804_n N_KAPWR_c_2586_n 0.0126311f $X=11.445 $Y=2.035 $X2=0
+ $Y2=0
cc_848 N_A_742_63#_c_802_n N_KAPWR_c_2587_n 0.0165853f $X=11.36 $Y=2.405 $X2=0
+ $Y2=0
cc_849 N_A_742_63#_M1050_g KAPWR 0.00257315f $X=13.15 $Y=2.345 $X2=0 $Y2=0
cc_850 N_A_742_63#_M1030_g KAPWR 0.00597578f $X=13.51 $Y=2.345 $X2=0 $Y2=0
cc_851 N_A_742_63#_c_803_n KAPWR 0.00150017f $X=11.91 $Y=2.035 $X2=0 $Y2=0
cc_852 N_A_742_63#_c_792_n N_KAPWR_c_2590_n 0.0144104f $X=7.075 $Y=2.99 $X2=0
+ $Y2=0
cc_853 N_A_742_63#_c_853_p N_KAPWR_c_2590_n 0.0149762f $X=7.16 $Y=2.905 $X2=0
+ $Y2=0
cc_854 N_A_742_63#_c_794_n N_KAPWR_c_2590_n 0.0403835f $X=9.41 $Y=2.435 $X2=0
+ $Y2=0
cc_855 N_A_742_63#_c_794_n N_KAPWR_c_2591_n 0.0517346f $X=9.41 $Y=2.435 $X2=0
+ $Y2=0
cc_856 N_A_742_63#_c_795_n N_KAPWR_c_2591_n 0.00231666f $X=9.495 $Y=2.725 $X2=0
+ $Y2=0
cc_857 N_A_742_63#_c_797_n N_KAPWR_c_2591_n 0.0122342f $X=9.58 $Y=2.81 $X2=0
+ $Y2=0
cc_858 N_A_742_63#_c_802_n N_KAPWR_c_2592_n 0.0155367f $X=11.36 $Y=2.405 $X2=0
+ $Y2=0
cc_859 N_A_742_63#_c_803_n N_KAPWR_c_2592_n 0.0210027f $X=11.91 $Y=2.035 $X2=0
+ $Y2=0
cc_860 N_A_742_63#_M1018_g N_KAPWR_c_2593_n 0.0107974f $X=3.785 $Y=0.655 $X2=0
+ $Y2=0
cc_861 N_A_742_63#_c_781_n N_KAPWR_c_2593_n 0.00706281f $X=5.055 $Y=3.15 $X2=0
+ $Y2=0
cc_862 N_A_742_63#_M1000_g N_KAPWR_c_2593_n 0.0121474f $X=5.13 $Y=2.305 $X2=0
+ $Y2=0
cc_863 N_A_742_63#_M1037_g N_KAPWR_c_2593_n 0.00836769f $X=5.49 $Y=2.305 $X2=0
+ $Y2=0
cc_864 N_A_742_63#_c_791_n N_KAPWR_c_2593_n 0.0262856f $X=5.295 $Y=2.905 $X2=0
+ $Y2=0
cc_865 N_A_742_63#_c_792_n N_KAPWR_c_2593_n 0.0482977f $X=7.075 $Y=2.99 $X2=0
+ $Y2=0
cc_866 N_A_742_63#_c_793_n N_KAPWR_c_2593_n 0.00352305f $X=5.38 $Y=2.99 $X2=0
+ $Y2=0
cc_867 N_A_742_63#_c_853_p N_KAPWR_c_2593_n 0.0169664f $X=7.16 $Y=2.905 $X2=0
+ $Y2=0
cc_868 N_A_742_63#_c_794_n N_KAPWR_c_2593_n 0.0186595f $X=9.41 $Y=2.435 $X2=0
+ $Y2=0
cc_869 N_A_742_63#_c_853_p N_KAPWR_c_2594_n 5.19653e-19 $X=7.16 $Y=2.905 $X2=0
+ $Y2=0
cc_870 N_A_742_63#_c_794_n N_KAPWR_c_2594_n 0.0168163f $X=9.41 $Y=2.435 $X2=0
+ $Y2=0
cc_871 N_A_742_63#_M1042_d N_KAPWR_c_2595_n 7.18337e-19 $X=11.22 $Y=2.095 $X2=0
+ $Y2=0
cc_872 N_A_742_63#_c_794_n N_KAPWR_c_2595_n 0.0264403f $X=9.41 $Y=2.435 $X2=0
+ $Y2=0
cc_873 N_A_742_63#_c_795_n N_KAPWR_c_2595_n 0.00637078f $X=9.495 $Y=2.725 $X2=0
+ $Y2=0
cc_874 N_A_742_63#_c_796_n N_KAPWR_c_2595_n 0.0410679f $X=10.505 $Y=2.81 $X2=0
+ $Y2=0
cc_875 N_A_742_63#_c_797_n N_KAPWR_c_2595_n 0.00617041f $X=9.58 $Y=2.81 $X2=0
+ $Y2=0
cc_876 N_A_742_63#_c_798_n N_KAPWR_c_2595_n 0.0125398f $X=10.59 $Y=2.725 $X2=0
+ $Y2=0
cc_877 N_A_742_63#_c_799_n N_KAPWR_c_2595_n 0.00608531f $X=10.855 $Y=2.095 $X2=0
+ $Y2=0
cc_878 N_A_742_63#_c_802_n N_KAPWR_c_2595_n 0.0192704f $X=11.36 $Y=2.405 $X2=0
+ $Y2=0
cc_879 N_A_742_63#_c_803_n N_KAPWR_c_2595_n 0.00486381f $X=11.91 $Y=2.035 $X2=0
+ $Y2=0
cc_880 N_A_742_63#_c_804_n N_KAPWR_c_2595_n 0.00622322f $X=11.445 $Y=2.035 $X2=0
+ $Y2=0
cc_881 N_A_742_63#_c_802_n N_KAPWR_c_2659_n 3.8211e-19 $X=11.36 $Y=2.405 $X2=0
+ $Y2=0
cc_882 N_A_742_63#_c_803_n N_KAPWR_c_2659_n 0.00105888f $X=11.91 $Y=2.035 $X2=0
+ $Y2=0
cc_883 N_A_742_63#_c_794_n A_1682_341# 0.00181239f $X=9.41 $Y=2.435 $X2=-0.19
+ $Y2=-0.245
cc_884 N_A_742_63#_M1050_g N_A_2562_427#_c_2779_n 0.0109499f $X=13.15 $Y=2.345
+ $X2=0 $Y2=0
cc_885 N_A_742_63#_M1030_g N_A_2562_427#_c_2779_n 0.00126733f $X=13.51 $Y=2.345
+ $X2=0 $Y2=0
cc_886 N_A_742_63#_M1050_g N_A_2562_427#_c_2780_n 0.00202281f $X=13.15 $Y=2.345
+ $X2=0 $Y2=0
cc_887 N_A_742_63#_M1030_g N_A_2562_427#_c_2780_n 0.00244237f $X=13.51 $Y=2.345
+ $X2=0 $Y2=0
cc_888 N_A_742_63#_M1018_g N_VGND_c_2831_n 0.0225355f $X=3.785 $Y=0.655 $X2=0
+ $Y2=0
cc_889 N_A_742_63#_M1018_g N_VGND_c_2840_n 0.00435433f $X=3.785 $Y=0.655 $X2=0
+ $Y2=0
cc_890 N_A_742_63#_c_770_n N_VGND_c_2842_n 0.00332046f $X=13.74 $Y=1.025 $X2=0
+ $Y2=0
cc_891 N_A_742_63#_M1018_g N_VGND_c_2845_n 0.0043858f $X=3.785 $Y=0.655 $X2=0
+ $Y2=0
cc_892 N_A_742_63#_c_770_n N_VGND_c_2845_n 0.00697981f $X=13.74 $Y=1.025 $X2=0
+ $Y2=0
cc_893 N_A_742_63#_M1018_g N_noxref_30_c_2994_n 0.0101402f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_894 N_A_742_63#_M1018_g N_noxref_32_c_3022_n 0.0205108f $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_895 N_A_742_63#_M1018_g N_noxref_32_c_3024_n 8.00494e-19 $X=3.785 $Y=0.655
+ $X2=0 $Y2=0
cc_896 N_A_742_63#_c_767_n N_A_1009_107#_c_3056_n 0.00101497f $X=5.5 $Y=1.605
+ $X2=0 $Y2=0
cc_897 N_A_666_89#_c_1082_n N_A_1343_51#_M1029_d 0.00272255f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_898 N_A_666_89#_c_1128_p N_A_1343_51#_M1015_d 0.00381504f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_899 N_A_666_89#_c_1085_n N_A_1343_51#_M1015_d 0.0040282f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_900 N_A_666_89#_c_1067_n N_A_1343_51#_c_1263_n 0.0113185f $X=6.29 $Y=1.605
+ $X2=0 $Y2=0
cc_901 N_A_666_89#_M1053_g N_A_1343_51#_M1010_g 0.0300902f $X=6.085 $Y=2.595
+ $X2=0 $Y2=0
cc_902 N_A_666_89#_c_1082_n N_A_1343_51#_M1010_g 0.00189766f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_903 N_A_666_89#_c_1083_n N_A_1343_51#_M1010_g 0.00161271f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_904 N_A_666_89#_c_1075_n N_A_1343_51#_M1010_g 0.017069f $X=6.29 $Y=1.77 $X2=0
+ $Y2=0
cc_905 N_A_666_89#_c_1076_n N_A_1343_51#_M1010_g 0.00700991f $X=6.32 $Y=1.77
+ $X2=0 $Y2=0
cc_906 N_A_666_89#_c_1067_n N_A_1343_51#_c_1267_n 0.00353474f $X=6.29 $Y=1.605
+ $X2=0 $Y2=0
cc_907 N_A_666_89#_c_1082_n N_A_1343_51#_c_1315_n 0.00444489f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_908 N_A_666_89#_M1013_g N_A_1343_51#_c_1279_n 0.0114202f $X=14.32 $Y=0.705
+ $X2=0 $Y2=0
cc_909 N_A_666_89#_M1002_g N_A_1343_51#_c_1279_n 0.00331974f $X=14.68 $Y=0.705
+ $X2=0 $Y2=0
cc_910 N_A_666_89#_M1015_g N_A_1343_51#_c_1340_n 0.00649957f $X=14.035 $Y=2.135
+ $X2=0 $Y2=0
cc_911 N_A_666_89#_c_1128_p N_A_1343_51#_c_1340_n 0.00772757f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_912 N_A_666_89#_c_1085_n N_A_1343_51#_c_1340_n 0.0236074f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_913 N_A_666_89#_c_1068_n N_A_1343_51#_c_1280_n 0.0032784f $X=14.035 $Y=1.565
+ $X2=0 $Y2=0
cc_914 N_A_666_89#_M1015_g N_A_1343_51#_c_1280_n 2.91251e-19 $X=14.035 $Y=2.135
+ $X2=0 $Y2=0
cc_915 N_A_666_89#_M1013_g N_A_1343_51#_c_1280_n 0.00790625f $X=14.32 $Y=0.705
+ $X2=0 $Y2=0
cc_916 N_A_666_89#_c_1070_n N_A_1343_51#_c_1280_n 0.00878495f $X=14.605 $Y=1.2
+ $X2=0 $Y2=0
cc_917 N_A_666_89#_M1002_g N_A_1343_51#_c_1280_n 0.0167481f $X=14.68 $Y=0.705
+ $X2=0 $Y2=0
cc_918 N_A_666_89#_c_1073_n N_A_1343_51#_c_1280_n 0.0239645f $X=14.22 $Y=1.29
+ $X2=0 $Y2=0
cc_919 N_A_666_89#_c_1085_n N_A_1343_51#_c_1280_n 0.00848817f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_920 N_A_666_89#_c_1082_n N_A_1343_51#_c_1289_n 0.0360498f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_921 N_A_666_89#_M1015_g N_A_1343_51#_c_1290_n 8.95332e-19 $X=14.035 $Y=2.135
+ $X2=0 $Y2=0
cc_922 N_A_666_89#_c_1070_n N_A_1343_51#_c_1290_n 0.00429463f $X=14.605 $Y=1.2
+ $X2=0 $Y2=0
cc_923 N_A_666_89#_c_1085_n N_A_1343_51#_c_1290_n 0.0130058f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_924 N_A_666_89#_c_1082_n N_A_1724_21#_M1014_g 0.0027536f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_925 N_A_666_89#_c_1082_n N_A_1724_21#_c_1481_n 0.00627708f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_926 N_A_666_89#_c_1082_n N_A_1724_21#_c_1495_n 0.0102504f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_927 N_A_666_89#_c_1082_n N_A_1724_21#_c_1496_n 0.0198668f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_928 N_A_666_89#_c_1082_n N_A_1724_21#_c_1497_n 0.0455982f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_929 N_A_666_89#_c_1082_n N_A_1113_419#_M1029_g 0.00292375f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_930 N_A_666_89#_c_1082_n N_A_1113_419#_c_1639_n 0.00307547f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_931 N_A_666_89#_M1053_g N_A_1113_419#_c_1642_n 0.0125393f $X=6.085 $Y=2.595
+ $X2=0 $Y2=0
cc_932 N_A_666_89#_c_1066_n N_A_1113_419#_c_1668_n 0.0108349f $X=5.93 $Y=1.605
+ $X2=0 $Y2=0
cc_933 N_A_666_89#_M1053_g N_A_1113_419#_c_1668_n 0.0145362f $X=6.085 $Y=2.595
+ $X2=0 $Y2=0
cc_934 N_A_666_89#_c_1067_n N_A_1113_419#_c_1668_n 0.00158258f $X=6.29 $Y=1.605
+ $X2=0 $Y2=0
cc_935 N_A_666_89#_c_1080_n N_A_1113_419#_c_1668_n 0.0526139f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_936 N_A_666_89#_c_1083_n N_A_1113_419#_c_1668_n 4.42833e-19 $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_937 N_A_666_89#_c_1075_n N_A_1113_419#_c_1668_n 0.014098f $X=6.29 $Y=1.77
+ $X2=0 $Y2=0
cc_938 N_A_666_89#_c_1076_n N_A_1113_419#_c_1668_n 0.0402273f $X=6.32 $Y=1.77
+ $X2=0 $Y2=0
cc_939 N_A_666_89#_M1053_g N_A_1113_419#_c_1672_n 0.0146958f $X=6.085 $Y=2.595
+ $X2=0 $Y2=0
cc_940 N_A_666_89#_c_1080_n N_A_1113_419#_c_1672_n 0.00734964f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_941 N_A_666_89#_c_1082_n N_A_1113_419#_c_1672_n 0.00466214f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_942 N_A_666_89#_c_1083_n N_A_1113_419#_c_1672_n 0.00295045f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_943 N_A_666_89#_c_1075_n N_A_1113_419#_c_1672_n 0.00108496f $X=6.29 $Y=1.77
+ $X2=0 $Y2=0
cc_944 N_A_666_89#_c_1076_n N_A_1113_419#_c_1672_n 0.0233029f $X=6.32 $Y=1.77
+ $X2=0 $Y2=0
cc_945 N_A_666_89#_M1053_g N_A_1113_419#_c_1699_n 7.82509e-19 $X=6.085 $Y=2.595
+ $X2=0 $Y2=0
cc_946 N_A_666_89#_c_1082_n N_A_1113_419#_c_1643_n 0.0509494f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_947 N_A_666_89#_M1053_g N_A_1113_419#_c_1653_n 3.65661e-19 $X=6.085 $Y=2.595
+ $X2=0 $Y2=0
cc_948 N_A_666_89#_c_1082_n N_A_1113_419#_c_1653_n 0.0191111f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_949 N_A_666_89#_c_1083_n N_A_1113_419#_c_1653_n 0.00186601f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_950 N_A_666_89#_c_1076_n N_A_1113_419#_c_1653_n 0.0138544f $X=6.32 $Y=1.77
+ $X2=0 $Y2=0
cc_951 N_A_666_89#_c_1082_n N_A_1113_419#_c_1644_n 0.0807862f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_952 N_A_666_89#_c_1082_n N_A_1113_419#_c_1646_n 0.00124435f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_953 N_A_666_89#_c_1082_n N_A_1113_419#_c_1656_n 0.0066373f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_954 N_A_666_89#_c_1082_n N_CLK_N_c_1779_n 0.00777589f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_955 N_A_666_89#_c_1082_n N_CLK_N_c_1780_n 0.0127393f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_956 N_A_666_89#_c_1082_n N_CLK_N_c_1781_n 0.014943f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_957 N_A_666_89#_c_1082_n N_SLEEP_B_c_1835_n 0.00908361f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_958 N_A_666_89#_c_1082_n N_SLEEP_B_c_1833_n 0.00291975f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_959 N_A_666_89#_c_1068_n N_A_2999_73#_M1051_g 0.00378616f $X=14.035 $Y=1.565
+ $X2=0 $Y2=0
cc_960 N_A_666_89#_M1002_g N_A_2999_73#_M1051_g 0.0453921f $X=14.68 $Y=0.705
+ $X2=0 $Y2=0
cc_961 N_A_666_89#_c_1082_n N_A_2717_427#_M1030_d 0.0026227f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_962 N_A_666_89#_c_1068_n N_A_2717_427#_c_2004_n 0.00466674f $X=14.035
+ $Y=1.565 $X2=0 $Y2=0
cc_963 N_A_666_89#_M1013_g N_A_2717_427#_c_2004_n 0.00432874f $X=14.32 $Y=0.705
+ $X2=0 $Y2=0
cc_964 N_A_666_89#_c_1073_n N_A_2717_427#_c_2004_n 0.00670583f $X=14.22 $Y=1.29
+ $X2=0 $Y2=0
cc_965 N_A_666_89#_c_1068_n N_A_2717_427#_c_2005_n 0.00660294f $X=14.035
+ $Y=1.565 $X2=0 $Y2=0
cc_966 N_A_666_89#_M1013_g N_A_2717_427#_c_2005_n 0.00152143f $X=14.32 $Y=0.705
+ $X2=0 $Y2=0
cc_967 N_A_666_89#_c_1073_n N_A_2717_427#_c_2005_n 0.06126f $X=14.22 $Y=1.29
+ $X2=0 $Y2=0
cc_968 N_A_666_89#_c_1082_n N_A_2717_427#_c_2005_n 0.0339651f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_969 N_A_666_89#_c_1128_p N_A_2717_427#_c_2005_n 0.00242593f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_970 N_A_666_89#_M1015_g N_A_2717_427#_c_2021_n 0.0102103f $X=14.035 $Y=2.135
+ $X2=0 $Y2=0
cc_971 N_A_666_89#_c_1082_n N_A_2717_427#_c_2021_n 0.00334833f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_972 N_A_666_89#_c_1128_p N_A_2717_427#_c_2021_n 0.00341592f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_973 N_A_666_89#_c_1085_n N_A_2717_427#_c_2021_n 0.00385038f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_974 N_A_666_89#_M1015_g N_A_2717_427#_c_2023_n 0.0037818f $X=14.035 $Y=2.135
+ $X2=0 $Y2=0
cc_975 N_A_666_89#_M1002_g N_A_2717_427#_c_2008_n 0.00133354f $X=14.68 $Y=0.705
+ $X2=0 $Y2=0
cc_976 N_A_666_89#_c_1080_n N_VPWR_M1021_d 0.0118289f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_977 N_A_666_89#_c_1080_n N_VPWR_c_2223_n 0.011034f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_978 N_A_666_89#_M1053_g N_VPWR_c_2235_n 0.00596462f $X=6.085 $Y=2.595 $X2=0
+ $Y2=0
cc_979 N_A_666_89#_M1053_g N_VPWR_c_2220_n 0.00773412f $X=6.085 $Y=2.595 $X2=0
+ $Y2=0
cc_980 N_A_666_89#_c_1080_n N_A_305_97#_M1049_d 0.00346118f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_981 N_A_666_89#_c_1072_n N_A_305_97#_c_2393_n 0.0148538f $X=3.465 $Y=1.43
+ $X2=0 $Y2=0
cc_982 N_A_666_89#_c_1072_n N_A_305_97#_c_2395_n 0.0125045f $X=3.465 $Y=1.43
+ $X2=0 $Y2=0
cc_983 N_A_666_89#_c_1081_n N_A_305_97#_c_2395_n 0.00699295f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_984 N_A_666_89#_c_1074_n N_A_305_97#_c_2395_n 0.0431836f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_985 N_A_666_89#_c_1074_n N_A_305_97#_c_2407_n 0.00686879f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_986 N_A_666_89#_c_1074_n N_A_305_97#_c_2408_n 0.0165161f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_987 N_A_666_89#_c_1080_n N_A_305_97#_c_2410_n 0.0237732f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_988 N_A_666_89#_c_1081_n N_A_305_97#_c_2410_n 0.00219752f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_989 N_A_666_89#_c_1074_n N_A_305_97#_c_2410_n 0.0484381f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_990 N_A_666_89#_c_1080_n N_A_305_97#_c_2396_n 0.0216996f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_991 N_A_666_89#_c_1074_n N_A_305_97#_c_2397_n 0.0120086f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_992 N_A_666_89#_c_1080_n N_A_305_97#_c_2458_n 0.0198305f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_993 N_A_666_89#_c_1080_n N_A_305_97#_c_2399_n 0.00709076f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_994 N_A_666_89#_c_1066_n N_A_305_97#_c_2400_n 0.0103345f $X=5.93 $Y=1.605
+ $X2=0 $Y2=0
cc_995 N_A_666_89#_c_1067_n N_A_305_97#_c_2400_n 0.00863658f $X=6.29 $Y=1.605
+ $X2=0 $Y2=0
cc_996 N_A_666_89#_c_1075_n N_A_305_97#_c_2400_n 8.80967e-19 $X=6.29 $Y=1.77
+ $X2=0 $Y2=0
cc_997 N_A_666_89#_c_1076_n N_A_305_97#_c_2400_n 0.00489394f $X=6.32 $Y=1.77
+ $X2=0 $Y2=0
cc_998 N_A_666_89#_c_1074_n N_A_305_97#_c_2412_n 0.0118473f $X=3.6 $Y=2.035
+ $X2=0 $Y2=0
cc_999 N_A_666_89#_c_1080_n N_A_305_97#_c_2413_n 0.0168935f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_1000 N_A_666_89#_c_1066_n N_A_305_97#_c_2403_n 0.00133388f $X=5.93 $Y=1.605
+ $X2=0 $Y2=0
cc_1001 N_A_666_89#_c_1067_n N_A_305_97#_c_2403_n 0.00823305f $X=6.29 $Y=1.605
+ $X2=0 $Y2=0
cc_1002 N_A_666_89#_c_1082_n N_A_305_97#_c_2403_n 0.00157445f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_1003 N_A_666_89#_c_1083_n N_A_305_97#_c_2403_n 0.003346f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_1004 N_A_666_89#_c_1075_n N_A_305_97#_c_2403_n 7.61794e-19 $X=6.29 $Y=1.77
+ $X2=0 $Y2=0
cc_1005 N_A_666_89#_c_1076_n N_A_305_97#_c_2403_n 0.0160056f $X=6.32 $Y=1.77
+ $X2=0 $Y2=0
cc_1006 N_A_666_89#_c_1080_n A_1041_419# 0.00129319f $X=6.335 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_1007 N_A_666_89#_c_1082_n A_1242_419# 8.21967e-19 $X=14.015 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_1008 N_A_666_89#_c_1083_n A_1242_419# 0.00239346f $X=6.625 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_1009 N_A_666_89#_c_1076_n A_1242_419# 0.00239124f $X=6.32 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_1010 N_A_666_89#_c_1082_n N_KAPWR_M1014_d 0.00332756f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_1011 N_A_666_89#_c_1082_n N_KAPWR_c_2586_n 0.00119666f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_1012 N_A_666_89#_c_1128_p KAPWR 0.0126511f $X=14.16 $Y=2.035 $X2=0 $Y2=0
cc_1013 N_A_666_89#_c_1085_n KAPWR 2.21315e-19 $X=14.16 $Y=2.035 $X2=0 $Y2=0
cc_1014 N_A_666_89#_c_1082_n N_KAPWR_c_2592_n 0.00257171f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_1015 N_A_666_89#_M1021_s N_KAPWR_c_2593_n 0.00165097f $X=3.425 $Y=2.095 $X2=0
+ $Y2=0
cc_1016 N_A_666_89#_M1053_g N_KAPWR_c_2593_n 0.00657926f $X=6.085 $Y=2.595 $X2=0
+ $Y2=0
cc_1017 N_A_666_89#_c_1081_n N_KAPWR_c_2593_n 0.0125132f $X=3.745 $Y=2.035 $X2=0
+ $Y2=0
cc_1018 N_A_666_89#_c_1083_n N_KAPWR_c_2593_n 0.0137398f $X=6.625 $Y=2.035 $X2=0
+ $Y2=0
cc_1019 N_A_666_89#_c_1074_n N_KAPWR_c_2593_n 0.0125124f $X=3.6 $Y=2.035 $X2=0
+ $Y2=0
cc_1020 N_A_666_89#_c_1082_n N_KAPWR_c_2594_n 0.0250226f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_1021 N_A_666_89#_c_1082_n N_KAPWR_c_2659_n 0.0113202f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_1022 N_A_666_89#_c_1082_n A_1682_341# 0.00158741f $X=14.015 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_1023 N_A_666_89#_c_1082_n N_A_2562_427#_c_2779_n 0.00876898f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_1024 N_A_666_89#_M1015_g N_A_2562_427#_c_2780_n 3.82123e-19 $X=14.035
+ $Y=2.135 $X2=0 $Y2=0
cc_1025 N_A_666_89#_M1002_g N_VGND_c_2835_n 0.00155595f $X=14.68 $Y=0.705 $X2=0
+ $Y2=0
cc_1026 N_A_666_89#_M1013_g N_VGND_c_2842_n 7.17276e-19 $X=14.32 $Y=0.705 $X2=0
+ $Y2=0
cc_1027 N_A_666_89#_M1002_g N_VGND_c_2842_n 0.00225337f $X=14.68 $Y=0.705 $X2=0
+ $Y2=0
cc_1028 N_A_666_89#_M1002_g N_VGND_c_2845_n 0.00185855f $X=14.68 $Y=0.705 $X2=0
+ $Y2=0
cc_1029 N_A_666_89#_M1018_s N_noxref_32_c_3022_n 0.0164357f $X=3.33 $Y=0.445
+ $X2=0 $Y2=0
cc_1030 N_A_666_89#_c_1072_n N_noxref_32_c_3022_n 0.0284617f $X=3.465 $Y=1.43
+ $X2=0 $Y2=0
cc_1031 N_A_666_89#_c_1066_n N_A_1009_107#_c_3056_n 0.00101497f $X=5.93 $Y=1.605
+ $X2=0 $Y2=0
cc_1032 N_A_666_89#_c_1067_n N_A_1009_107#_c_3056_n 0.00100792f $X=6.29 $Y=1.605
+ $X2=0 $Y2=0
cc_1033 N_A_1343_51#_c_1271_n N_A_1724_21#_M1027_g 0.00964111f $X=8.44 $Y=1.67
+ $X2=0 $Y2=0
cc_1034 N_A_1343_51#_c_1272_n N_A_1724_21#_M1027_g 0.0161292f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1035 N_A_1343_51#_c_1289_n N_A_1724_21#_M1014_g 0.0159438f $X=9.63 $Y=1.715
+ $X2=0 $Y2=0
cc_1036 N_A_1343_51#_c_1272_n N_A_1724_21#_c_1481_n 0.0261955f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1037 N_A_1343_51#_c_1288_n N_A_1724_21#_c_1481_n 0.0215052f $X=9.795 $Y=1.755
+ $X2=0 $Y2=0
cc_1038 N_A_1343_51#_c_1289_n N_A_1724_21#_c_1481_n 0.02728f $X=9.63 $Y=1.715
+ $X2=0 $Y2=0
cc_1039 N_A_1343_51#_c_1272_n N_A_1724_21#_c_1482_n 0.0132812f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1040 N_A_1343_51#_c_1273_n N_A_1724_21#_c_1482_n 0.00864203f $X=9.7 $Y=0.465
+ $X2=0 $Y2=0
cc_1041 N_A_1343_51#_c_1274_n N_A_1724_21#_c_1483_n 0.0747432f $X=11.535 $Y=0.34
+ $X2=0 $Y2=0
cc_1042 N_A_1343_51#_c_1273_n N_A_1724_21#_c_1484_n 0.0150383f $X=9.7 $Y=0.465
+ $X2=0 $Y2=0
cc_1043 N_A_1343_51#_c_1274_n N_A_1724_21#_c_1484_n 0.0134313f $X=11.535 $Y=0.34
+ $X2=0 $Y2=0
cc_1044 N_A_1343_51#_c_1274_n N_A_1724_21#_c_1486_n 0.00567979f $X=11.535
+ $Y=0.34 $X2=0 $Y2=0
cc_1045 N_A_1343_51#_c_1366_p N_A_1724_21#_c_1486_n 0.0589068f $X=12.425 $Y=0.7
+ $X2=0 $Y2=0
cc_1046 N_A_1343_51#_c_1367_p N_A_1724_21#_c_1486_n 0.0106593f $X=11.705 $Y=0.7
+ $X2=0 $Y2=0
cc_1047 N_A_1343_51#_c_1282_n N_A_1724_21#_c_1486_n 0.00485081f $X=13.325
+ $Y=0.435 $X2=0 $Y2=0
cc_1048 N_A_1343_51#_c_1282_n N_A_1724_21#_c_1488_n 0.0225977f $X=13.325
+ $Y=0.435 $X2=0 $Y2=0
cc_1049 N_A_1343_51#_c_1283_n N_A_1724_21#_c_1488_n 0.00128541f $X=13.655
+ $Y=0.435 $X2=0 $Y2=0
cc_1050 N_A_1343_51#_c_1282_n N_A_1724_21#_c_1489_n 0.00786824f $X=13.325
+ $Y=0.435 $X2=0 $Y2=0
cc_1051 N_A_1343_51#_c_1283_n N_A_1724_21#_c_1489_n 0.00855967f $X=13.655
+ $Y=0.435 $X2=0 $Y2=0
cc_1052 N_A_1343_51#_c_1272_n N_A_1724_21#_c_1491_n 0.00629234f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1053 N_A_1343_51#_c_1289_n N_A_1724_21#_c_1491_n 0.00355769f $X=9.63 $Y=1.715
+ $X2=0 $Y2=0
cc_1054 N_A_1343_51#_c_1271_n N_A_1724_21#_c_1492_n 0.0221138f $X=8.44 $Y=1.67
+ $X2=0 $Y2=0
cc_1055 N_A_1343_51#_c_1272_n N_A_1724_21#_c_1492_n 0.0608836f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1056 N_A_1343_51#_c_1289_n N_A_1724_21#_c_1492_n 0.0228999f $X=9.63 $Y=1.715
+ $X2=0 $Y2=0
cc_1057 N_A_1343_51#_c_1273_n N_A_1113_419#_c_1634_n 0.00112601f $X=9.7 $Y=0.465
+ $X2=0 $Y2=0
cc_1058 N_A_1343_51#_c_1275_n N_A_1113_419#_c_1634_n 4.60652e-19 $X=9.865
+ $Y=0.34 $X2=0 $Y2=0
cc_1059 N_A_1343_51#_c_1288_n N_A_1113_419#_M1029_g 0.0023126f $X=9.795 $Y=1.755
+ $X2=0 $Y2=0
cc_1060 N_A_1343_51#_c_1289_n N_A_1113_419#_M1029_g 0.0170082f $X=9.63 $Y=1.715
+ $X2=0 $Y2=0
cc_1061 N_A_1343_51#_c_1273_n N_A_1113_419#_c_1636_n 0.00769324f $X=9.7 $Y=0.465
+ $X2=0 $Y2=0
cc_1062 N_A_1343_51#_c_1275_n N_A_1113_419#_c_1636_n 0.00329177f $X=9.865
+ $Y=0.34 $X2=0 $Y2=0
cc_1063 N_A_1343_51#_c_1272_n N_A_1113_419#_c_1637_n 0.0152295f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1064 N_A_1343_51#_c_1274_n N_A_1113_419#_c_1637_n 0.00520355f $X=11.535
+ $Y=0.34 $X2=0 $Y2=0
cc_1065 N_A_1343_51#_c_1272_n N_A_1113_419#_c_1638_n 0.0369177f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1066 N_A_1343_51#_c_1273_n N_A_1113_419#_c_1638_n 0.00733755f $X=9.7 $Y=0.465
+ $X2=0 $Y2=0
cc_1067 N_A_1343_51#_c_1288_n N_A_1113_419#_c_1639_n 0.00289859f $X=9.795
+ $Y=1.755 $X2=0 $Y2=0
cc_1068 N_A_1343_51#_M1010_g N_A_1113_419#_c_1672_n 0.012125f $X=6.85 $Y=2.595
+ $X2=0 $Y2=0
cc_1069 N_A_1343_51#_M1010_g N_A_1113_419#_c_1699_n 0.00953687f $X=6.85 $Y=2.595
+ $X2=0 $Y2=0
cc_1070 N_A_1343_51#_M1010_g N_A_1113_419#_c_1643_n 0.00957708f $X=6.85 $Y=2.595
+ $X2=0 $Y2=0
cc_1071 N_A_1343_51#_c_1284_n N_A_1113_419#_c_1643_n 0.00100043f $X=7.19
+ $Y=1.282 $X2=0 $Y2=0
cc_1072 N_A_1343_51#_M1010_g N_A_1113_419#_c_1653_n 0.0129624f $X=6.85 $Y=2.595
+ $X2=0 $Y2=0
cc_1073 N_A_1343_51#_M1029_d N_A_1113_419#_c_1644_n 0.00754484f $X=9.56 $Y=1.705
+ $X2=0 $Y2=0
cc_1074 N_A_1343_51#_c_1315_n N_A_1113_419#_c_1644_n 0.00870478f $X=8.525
+ $Y=1.755 $X2=0 $Y2=0
cc_1075 N_A_1343_51#_c_1289_n N_A_1113_419#_c_1644_n 0.079081f $X=9.63 $Y=1.715
+ $X2=0 $Y2=0
cc_1076 N_A_1343_51#_c_1274_n N_CLK_N_M1038_g 0.00782537f $X=11.535 $Y=0.34
+ $X2=0 $Y2=0
cc_1077 N_A_1343_51#_c_1288_n N_CLK_N_c_1781_n 0.0171813f $X=9.795 $Y=1.755
+ $X2=0 $Y2=0
cc_1078 N_A_1343_51#_c_1274_n N_SLEEP_B_c_1826_n 0.00696485f $X=11.535 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_1079 N_A_1343_51#_c_1276_n N_SLEEP_B_c_1826_n 0.0015257f $X=11.62 $Y=0.615
+ $X2=-0.19 $Y2=-0.245
cc_1080 N_A_1343_51#_c_1274_n N_SLEEP_B_c_1828_n 0.00371788f $X=11.535 $Y=0.34
+ $X2=0 $Y2=0
cc_1081 N_A_1343_51#_c_1276_n N_SLEEP_B_c_1828_n 0.00545448f $X=11.62 $Y=0.615
+ $X2=0 $Y2=0
cc_1082 N_A_1343_51#_c_1366_p N_SLEEP_B_c_1828_n 0.00471953f $X=12.425 $Y=0.7
+ $X2=0 $Y2=0
cc_1083 N_A_1343_51#_c_1367_p N_SLEEP_B_c_1828_n 0.00399764f $X=11.705 $Y=0.7
+ $X2=0 $Y2=0
cc_1084 N_A_1343_51#_c_1276_n N_SLEEP_B_c_1829_n 8.61234e-19 $X=11.62 $Y=0.615
+ $X2=0 $Y2=0
cc_1085 N_A_1343_51#_c_1366_p N_SLEEP_B_c_1829_n 0.0115442f $X=12.425 $Y=0.7
+ $X2=0 $Y2=0
cc_1086 N_A_1343_51#_c_1277_n N_SLEEP_B_c_1829_n 0.00161884f $X=12.51 $Y=0.615
+ $X2=0 $Y2=0
cc_1087 N_A_1343_51#_c_1278_n N_SLEEP_B_c_1829_n 7.03875e-19 $X=12.595 $Y=0.34
+ $X2=0 $Y2=0
cc_1088 N_A_1343_51#_c_1366_p N_SLEEP_B_c_1830_n 4.00046e-19 $X=12.425 $Y=0.7
+ $X2=0 $Y2=0
cc_1089 N_A_1343_51#_c_1366_p N_SLEEP_B_c_1831_n 0.00195584f $X=12.425 $Y=0.7
+ $X2=0 $Y2=0
cc_1090 N_A_1343_51#_c_1277_n N_SLEEP_B_c_1832_n 0.00186466f $X=12.51 $Y=0.615
+ $X2=0 $Y2=0
cc_1091 N_A_1343_51#_c_1282_n N_SLEEP_B_c_1832_n 0.00913631f $X=13.325 $Y=0.435
+ $X2=0 $Y2=0
cc_1092 N_A_1343_51#_c_1283_n N_SLEEP_B_c_1832_n 0.00396769f $X=13.655 $Y=0.435
+ $X2=0 $Y2=0
cc_1093 N_A_1343_51#_c_1340_n N_A_2999_73#_M1051_g 8.3168e-19 $X=14.5 $Y=1.86
+ $X2=0 $Y2=0
cc_1094 N_A_1343_51#_c_1280_n N_A_2999_73#_M1051_g 0.00392929f $X=14.615
+ $Y=1.625 $X2=0 $Y2=0
cc_1095 N_A_1343_51#_c_1290_n N_A_2999_73#_M1051_g 9.14966e-19 $X=14.615 $Y=1.71
+ $X2=0 $Y2=0
cc_1096 N_A_1343_51#_c_1340_n N_A_2999_73#_c_1932_n 6.79371e-19 $X=14.5 $Y=1.86
+ $X2=0 $Y2=0
cc_1097 N_A_1343_51#_c_1279_n N_A_2717_427#_M1044_d 0.00337304f $X=14.53 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_1098 N_A_1343_51#_c_1279_n N_A_2717_427#_c_2004_n 0.0259673f $X=14.53 $Y=0.34
+ $X2=0 $Y2=0
cc_1099 N_A_1343_51#_c_1280_n N_A_2717_427#_c_2004_n 0.0157621f $X=14.615
+ $Y=1.625 $X2=0 $Y2=0
cc_1100 N_A_1343_51#_c_1280_n N_A_2717_427#_c_2005_n 0.00525316f $X=14.615
+ $Y=1.625 $X2=0 $Y2=0
cc_1101 N_A_1343_51#_c_1340_n N_A_2717_427#_c_2021_n 0.0126871f $X=14.5 $Y=1.86
+ $X2=0 $Y2=0
cc_1102 N_A_1343_51#_c_1340_n N_A_2717_427#_c_2023_n 0.0191837f $X=14.5 $Y=1.86
+ $X2=0 $Y2=0
cc_1103 N_A_1343_51#_c_1340_n N_A_2717_427#_c_2006_n 0.00848349f $X=14.5 $Y=1.86
+ $X2=0 $Y2=0
cc_1104 N_A_1343_51#_c_1280_n N_A_2717_427#_c_2006_n 0.0263153f $X=14.615
+ $Y=1.625 $X2=0 $Y2=0
cc_1105 N_A_1343_51#_c_1290_n N_A_2717_427#_c_2006_n 0.0132277f $X=14.615
+ $Y=1.71 $X2=0 $Y2=0
cc_1106 N_A_1343_51#_c_1280_n N_A_2717_427#_c_2008_n 0.0136811f $X=14.615
+ $Y=1.625 $X2=0 $Y2=0
cc_1107 N_A_1343_51#_c_1340_n N_A_2717_427#_c_2025_n 0.0124299f $X=14.5 $Y=1.86
+ $X2=0 $Y2=0
cc_1108 N_A_1343_51#_M1010_g N_VPWR_c_2235_n 0.00596462f $X=6.85 $Y=2.595 $X2=0
+ $Y2=0
cc_1109 N_A_1343_51#_M1010_g N_VPWR_c_2220_n 0.00885411f $X=6.85 $Y=2.595 $X2=0
+ $Y2=0
cc_1110 N_A_1343_51#_c_1263_n N_A_305_97#_c_2403_n 0.00379199f $X=6.8 $Y=1.305
+ $X2=0 $Y2=0
cc_1111 N_A_1343_51#_c_1267_n N_A_305_97#_c_2403_n 0.00139622f $X=6.795 $Y=1.065
+ $X2=0 $Y2=0
cc_1112 N_A_1343_51#_c_1289_n N_KAPWR_M1014_d 0.00370871f $X=9.63 $Y=1.715 $X2=0
+ $Y2=0
cc_1113 N_A_1343_51#_c_1340_n KAPWR 0.00107507f $X=14.5 $Y=1.86 $X2=0 $Y2=0
cc_1114 N_A_1343_51#_M1010_g N_KAPWR_c_2590_n 9.22952e-19 $X=6.85 $Y=2.595 $X2=0
+ $Y2=0
cc_1115 N_A_1343_51#_M1010_g N_KAPWR_c_2593_n 0.0101976f $X=6.85 $Y=2.595 $X2=0
+ $Y2=0
cc_1116 N_A_1343_51#_M1029_d N_KAPWR_c_2595_n 0.00422144f $X=9.56 $Y=1.705 $X2=0
+ $Y2=0
cc_1117 N_A_1343_51#_c_1315_n A_1682_341# 5.76994e-19 $X=8.525 $Y=1.755
+ $X2=-0.19 $Y2=-0.245
cc_1118 N_A_1343_51#_c_1289_n A_1682_341# 3.53584e-19 $X=9.63 $Y=1.715 $X2=-0.19
+ $Y2=-0.245
cc_1119 N_A_1343_51#_c_1366_p N_VGND_M1043_d 0.00991913f $X=12.425 $Y=0.7 $X2=0
+ $Y2=0
cc_1120 N_A_1343_51#_c_1272_n N_VGND_c_2833_n 0.0184719f $X=9.535 $Y=0.96 $X2=0
+ $Y2=0
cc_1121 N_A_1343_51#_c_1273_n N_VGND_c_2833_n 0.00817341f $X=9.7 $Y=0.465 $X2=0
+ $Y2=0
cc_1122 N_A_1343_51#_c_1275_n N_VGND_c_2833_n 0.00591401f $X=9.865 $Y=0.34 $X2=0
+ $Y2=0
cc_1123 N_A_1343_51#_c_1274_n N_VGND_c_2834_n 0.0123391f $X=11.535 $Y=0.34 $X2=0
+ $Y2=0
cc_1124 N_A_1343_51#_c_1276_n N_VGND_c_2834_n 0.00122418f $X=11.62 $Y=0.615
+ $X2=0 $Y2=0
cc_1125 N_A_1343_51#_c_1366_p N_VGND_c_2834_n 0.0188164f $X=12.425 $Y=0.7 $X2=0
+ $Y2=0
cc_1126 N_A_1343_51#_c_1277_n N_VGND_c_2834_n 0.0011095f $X=12.51 $Y=0.615 $X2=0
+ $Y2=0
cc_1127 N_A_1343_51#_c_1278_n N_VGND_c_2834_n 0.0108033f $X=12.595 $Y=0.34 $X2=0
+ $Y2=0
cc_1128 N_A_1343_51#_c_1279_n N_VGND_c_2835_n 0.00749734f $X=14.53 $Y=0.34 $X2=0
+ $Y2=0
cc_1129 N_A_1343_51#_c_1280_n N_VGND_c_2835_n 0.0175266f $X=14.615 $Y=1.625
+ $X2=0 $Y2=0
cc_1130 N_A_1343_51#_c_1274_n N_VGND_c_2837_n 0.119481f $X=11.535 $Y=0.34 $X2=0
+ $Y2=0
cc_1131 N_A_1343_51#_c_1275_n N_VGND_c_2837_n 0.0211917f $X=9.865 $Y=0.34 $X2=0
+ $Y2=0
cc_1132 N_A_1343_51#_c_1366_p N_VGND_c_2837_n 0.00323373f $X=12.425 $Y=0.7 $X2=0
+ $Y2=0
cc_1133 N_A_1343_51#_M1035_g N_VGND_c_2841_n 0.00540915f $X=7.19 $Y=0.595 $X2=0
+ $Y2=0
cc_1134 N_A_1343_51#_c_1266_n N_VGND_c_2841_n 0.00388395f $X=6.795 $Y=0.915
+ $X2=0 $Y2=0
cc_1135 N_A_1343_51#_c_1366_p N_VGND_c_2842_n 0.00400574f $X=12.425 $Y=0.7 $X2=0
+ $Y2=0
cc_1136 N_A_1343_51#_c_1278_n N_VGND_c_2842_n 0.0119604f $X=12.595 $Y=0.34 $X2=0
+ $Y2=0
cc_1137 N_A_1343_51#_c_1279_n N_VGND_c_2842_n 0.0121867f $X=14.53 $Y=0.34 $X2=0
+ $Y2=0
cc_1138 N_A_1343_51#_c_1282_n N_VGND_c_2842_n 0.125255f $X=13.325 $Y=0.435 $X2=0
+ $Y2=0
cc_1139 N_A_1343_51#_M1032_d N_VGND_c_2845_n 0.00232718f $X=9.56 $Y=0.235 $X2=0
+ $Y2=0
cc_1140 N_A_1343_51#_M1035_g N_VGND_c_2845_n 0.0054106f $X=7.19 $Y=0.595 $X2=0
+ $Y2=0
cc_1141 N_A_1343_51#_c_1266_n N_VGND_c_2845_n 0.0054106f $X=6.795 $Y=0.915 $X2=0
+ $Y2=0
cc_1142 N_A_1343_51#_c_1274_n N_VGND_c_2845_n 0.069347f $X=11.535 $Y=0.34 $X2=0
+ $Y2=0
cc_1143 N_A_1343_51#_c_1275_n N_VGND_c_2845_n 0.0127152f $X=9.865 $Y=0.34 $X2=0
+ $Y2=0
cc_1144 N_A_1343_51#_c_1366_p N_VGND_c_2845_n 0.0146704f $X=12.425 $Y=0.7 $X2=0
+ $Y2=0
cc_1145 N_A_1343_51#_c_1278_n N_VGND_c_2845_n 0.00656672f $X=12.595 $Y=0.34
+ $X2=0 $Y2=0
cc_1146 N_A_1343_51#_c_1279_n N_VGND_c_2845_n 0.00660921f $X=14.53 $Y=0.34 $X2=0
+ $Y2=0
cc_1147 N_A_1343_51#_c_1282_n N_VGND_c_2845_n 0.0722643f $X=13.325 $Y=0.435
+ $X2=0 $Y2=0
cc_1148 N_A_1343_51#_M1035_g N_VGND_c_2848_n 0.00284344f $X=7.19 $Y=0.595 $X2=0
+ $Y2=0
cc_1149 N_A_1343_51#_c_1266_n N_A_1009_107#_c_3056_n 0.00235098f $X=6.795
+ $Y=0.915 $X2=0 $Y2=0
cc_1150 N_A_1343_51#_c_1269_n N_A_1453_77#_c_3075_n 0.0551213f $X=8.355 $Y=0.96
+ $X2=0 $Y2=0
cc_1151 N_A_1343_51#_M1035_g N_A_1453_77#_c_3076_n 0.00436134f $X=7.19 $Y=0.595
+ $X2=0 $Y2=0
cc_1152 N_A_1343_51#_c_1270_n N_A_1453_77#_c_3076_n 0.025806f $X=7.57 $Y=0.96
+ $X2=0 $Y2=0
cc_1153 N_A_1343_51#_c_1284_n N_A_1453_77#_c_3076_n 0.00123101f $X=7.19 $Y=1.282
+ $X2=0 $Y2=0
cc_1154 N_A_1343_51#_c_1269_n N_A_1453_77#_c_3077_n 0.00295363f $X=8.355 $Y=0.96
+ $X2=0 $Y2=0
cc_1155 N_A_1343_51#_c_1272_n N_A_1453_77#_c_3077_n 0.00948583f $X=9.535 $Y=0.96
+ $X2=0 $Y2=0
cc_1156 N_A_1343_51#_c_1281_n N_A_1453_77#_c_3077_n 0.0154492f $X=8.44 $Y=0.96
+ $X2=0 $Y2=0
cc_1157 N_A_1343_51#_c_1366_p A_2480_97# 0.00128354f $X=12.425 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_1158 N_A_1343_51#_c_1280_n A_2879_99# 0.00480249f $X=14.615 $Y=1.625
+ $X2=-0.19 $Y2=-0.245
cc_1159 N_A_1724_21#_M1027_g N_A_1113_419#_c_1634_n 0.0206434f $X=8.695 $Y=0.445
+ $X2=0 $Y2=0
cc_1160 N_A_1724_21#_M1014_g N_A_1113_419#_M1029_g 0.0390064f $X=8.745 $Y=2.205
+ $X2=0 $Y2=0
cc_1161 N_A_1724_21#_c_1481_n N_A_1113_419#_M1029_g 0.0166142f $X=10.035 $Y=1.3
+ $X2=0 $Y2=0
cc_1162 N_A_1724_21#_c_1482_n N_A_1113_419#_M1029_g 8.34208e-19 $X=10.12
+ $Y=1.215 $X2=0 $Y2=0
cc_1163 N_A_1724_21#_c_1491_n N_A_1113_419#_M1029_g 0.0149607f $X=8.86 $Y=1.355
+ $X2=0 $Y2=0
cc_1164 N_A_1724_21#_c_1492_n N_A_1113_419#_M1029_g 7.51638e-19 $X=9.025
+ $Y=1.357 $X2=0 $Y2=0
cc_1165 N_A_1724_21#_c_1484_n N_A_1113_419#_c_1636_n 5.59254e-19 $X=10.205
+ $Y=0.68 $X2=0 $Y2=0
cc_1166 N_A_1724_21#_c_1481_n N_A_1113_419#_c_1637_n 0.0056001f $X=10.035 $Y=1.3
+ $X2=0 $Y2=0
cc_1167 N_A_1724_21#_c_1482_n N_A_1113_419#_c_1637_n 0.00815228f $X=10.12
+ $Y=1.215 $X2=0 $Y2=0
cc_1168 N_A_1724_21#_M1027_g N_A_1113_419#_c_1638_n 0.00642855f $X=8.695
+ $Y=0.445 $X2=0 $Y2=0
cc_1169 N_A_1724_21#_c_1481_n N_A_1113_419#_c_1638_n 0.00131154f $X=10.035
+ $Y=1.3 $X2=0 $Y2=0
cc_1170 N_A_1724_21#_c_1482_n N_A_1113_419#_c_1638_n 5.52585e-19 $X=10.12
+ $Y=1.215 $X2=0 $Y2=0
cc_1171 N_A_1724_21#_c_1481_n N_A_1113_419#_c_1639_n 0.0129201f $X=10.035 $Y=1.3
+ $X2=0 $Y2=0
cc_1172 N_A_1724_21#_c_1482_n N_A_1113_419#_c_1639_n 0.00550182f $X=10.12
+ $Y=1.215 $X2=0 $Y2=0
cc_1173 N_A_1724_21#_M1014_g N_A_1113_419#_c_1644_n 0.0135207f $X=8.745 $Y=2.205
+ $X2=0 $Y2=0
cc_1174 N_A_1724_21#_c_1481_n N_A_1113_419#_c_1644_n 0.0035521f $X=10.035 $Y=1.3
+ $X2=0 $Y2=0
cc_1175 N_A_1724_21#_M1014_g N_A_1113_419#_c_1656_n 3.97083e-19 $X=8.745
+ $Y=2.205 $X2=0 $Y2=0
cc_1176 N_A_1724_21#_c_1481_n N_CLK_N_M1038_g 0.00105344f $X=10.035 $Y=1.3 $X2=0
+ $Y2=0
cc_1177 N_A_1724_21#_c_1482_n N_CLK_N_M1038_g 0.00394902f $X=10.12 $Y=1.215
+ $X2=0 $Y2=0
cc_1178 N_A_1724_21#_c_1483_n N_CLK_N_M1038_g 0.0121998f $X=11.195 $Y=0.68 $X2=0
+ $Y2=0
cc_1179 N_A_1724_21#_c_1485_n N_CLK_N_M1038_g 9.99211e-19 $X=11.28 $Y=0.955
+ $X2=0 $Y2=0
cc_1180 N_A_1724_21#_c_1487_n N_CLK_N_M1038_g 6.07096e-19 $X=11.365 $Y=1.04
+ $X2=0 $Y2=0
cc_1181 N_A_1724_21#_c_1483_n N_SLEEP_B_c_1826_n 0.0065832f $X=11.195 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_1182 N_A_1724_21#_c_1485_n N_SLEEP_B_c_1826_n 0.00510565f $X=11.28 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_1183 N_A_1724_21#_c_1486_n N_SLEEP_B_c_1826_n 9.63172e-19 $X=12.765 $Y=1.04
+ $X2=-0.19 $Y2=-0.245
cc_1184 N_A_1724_21#_c_1487_n N_SLEEP_B_c_1826_n 9.32883e-19 $X=11.365 $Y=1.04
+ $X2=-0.19 $Y2=-0.245
cc_1185 N_A_1724_21#_c_1496_n N_SLEEP_B_M1019_g 9.92583e-19 $X=12.415 $Y=2.59
+ $X2=0 $Y2=0
cc_1186 N_A_1724_21#_c_1485_n N_SLEEP_B_c_1828_n 0.0011203f $X=11.28 $Y=0.955
+ $X2=0 $Y2=0
cc_1187 N_A_1724_21#_c_1486_n N_SLEEP_B_c_1828_n 0.00444505f $X=12.765 $Y=1.04
+ $X2=0 $Y2=0
cc_1188 N_A_1724_21#_c_1495_n N_SLEEP_B_c_1835_n 0.00569139f $X=12.415 $Y=2.075
+ $X2=0 $Y2=0
cc_1189 N_A_1724_21#_c_1496_n N_SLEEP_B_c_1835_n 0.012232f $X=12.415 $Y=2.59
+ $X2=0 $Y2=0
cc_1190 N_A_1724_21#_c_1486_n N_SLEEP_B_c_1829_n 0.00453317f $X=12.765 $Y=1.04
+ $X2=0 $Y2=0
cc_1191 N_A_1724_21#_c_1488_n N_SLEEP_B_c_1829_n 9.77449e-19 $X=12.93 $Y=0.76
+ $X2=0 $Y2=0
cc_1192 N_A_1724_21#_c_1486_n N_SLEEP_B_c_1830_n 0.00758921f $X=12.765 $Y=1.04
+ $X2=0 $Y2=0
cc_1193 N_A_1724_21#_c_1490_n N_SLEEP_B_c_1830_n 6.7576e-19 $X=13.4 $Y=1.905
+ $X2=0 $Y2=0
cc_1194 N_A_1724_21#_c_1493_n N_SLEEP_B_c_1830_n 0.00274048f $X=12.93 $Y=1.04
+ $X2=0 $Y2=0
cc_1195 N_A_1724_21#_c_1486_n N_SLEEP_B_c_1831_n 0.0409663f $X=12.765 $Y=1.04
+ $X2=0 $Y2=0
cc_1196 N_A_1724_21#_c_1487_n N_SLEEP_B_c_1831_n 0.00366943f $X=11.365 $Y=1.04
+ $X2=0 $Y2=0
cc_1197 N_A_1724_21#_c_1486_n N_SLEEP_B_c_1832_n 0.00444921f $X=12.765 $Y=1.04
+ $X2=0 $Y2=0
cc_1198 N_A_1724_21#_c_1488_n N_SLEEP_B_c_1832_n 0.00617657f $X=12.93 $Y=0.76
+ $X2=0 $Y2=0
cc_1199 N_A_1724_21#_c_1493_n N_SLEEP_B_c_1832_n 0.00154151f $X=12.93 $Y=1.04
+ $X2=0 $Y2=0
cc_1200 N_A_1724_21#_c_1486_n N_SLEEP_B_c_1833_n 0.0143343f $X=12.765 $Y=1.04
+ $X2=0 $Y2=0
cc_1201 N_A_1724_21#_c_1487_n N_SLEEP_B_c_1833_n 0.013977f $X=11.365 $Y=1.04
+ $X2=0 $Y2=0
cc_1202 N_A_1724_21#_c_1488_n N_A_2717_427#_c_2004_n 0.00383661f $X=12.93
+ $Y=0.76 $X2=0 $Y2=0
cc_1203 N_A_1724_21#_c_1497_n N_A_2717_427#_c_2005_n 0.0123973f $X=13.315
+ $Y=1.99 $X2=0 $Y2=0
cc_1204 N_A_1724_21#_c_1489_n N_A_2717_427#_c_2005_n 0.0138559f $X=13.315
+ $Y=1.04 $X2=0 $Y2=0
cc_1205 N_A_1724_21#_c_1490_n N_A_2717_427#_c_2005_n 0.0571856f $X=13.4 $Y=1.905
+ $X2=0 $Y2=0
cc_1206 N_A_1724_21#_c_1496_n N_VPWR_c_2235_n 0.00762755f $X=12.415 $Y=2.59
+ $X2=0 $Y2=0
cc_1207 N_A_1724_21#_c_1496_n N_VPWR_c_2220_n 9.33125e-19 $X=12.415 $Y=2.59
+ $X2=0 $Y2=0
cc_1208 N_A_1724_21#_c_1496_n KAPWR 0.028071f $X=12.415 $Y=2.59 $X2=0 $Y2=0
cc_1209 N_A_1724_21#_c_1497_n KAPWR 0.0118878f $X=13.315 $Y=1.99 $X2=0 $Y2=0
cc_1210 N_A_1724_21#_M1014_g N_KAPWR_c_2591_n 0.0104874f $X=8.745 $Y=2.205 $X2=0
+ $Y2=0
cc_1211 N_A_1724_21#_c_1496_n N_KAPWR_c_2592_n 0.0300531f $X=12.415 $Y=2.59
+ $X2=0 $Y2=0
cc_1212 N_A_1724_21#_M1014_g N_KAPWR_c_2594_n 2.41362e-19 $X=8.745 $Y=2.205
+ $X2=0 $Y2=0
cc_1213 N_A_1724_21#_M1014_g N_KAPWR_c_2595_n 0.00253459f $X=8.745 $Y=2.205
+ $X2=0 $Y2=0
cc_1214 N_A_1724_21#_c_1496_n N_A_2562_427#_c_2779_n 0.0382716f $X=12.415
+ $Y=2.59 $X2=0 $Y2=0
cc_1215 N_A_1724_21#_c_1497_n N_A_2562_427#_c_2779_n 0.0212889f $X=13.315
+ $Y=1.99 $X2=0 $Y2=0
cc_1216 N_A_1724_21#_M1027_g N_VGND_c_2832_n 0.0054895f $X=8.695 $Y=0.445 $X2=0
+ $Y2=0
cc_1217 N_A_1724_21#_M1027_g N_VGND_c_2833_n 0.00309362f $X=8.695 $Y=0.445 $X2=0
+ $Y2=0
cc_1218 N_A_1724_21#_M1027_g N_VGND_c_2845_n 0.0100257f $X=8.695 $Y=0.445 $X2=0
+ $Y2=0
cc_1219 N_A_1724_21#_M1027_g N_A_1453_77#_c_3077_n 0.00617706f $X=8.695 $Y=0.445
+ $X2=0 $Y2=0
cc_1220 N_A_1724_21#_c_1483_n A_2198_97# 0.00608736f $X=11.195 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_1221 N_A_1113_419#_c_1637_n N_CLK_N_M1038_g 0.00794864f $X=9.995 $Y=0.99
+ $X2=0 $Y2=0
cc_1222 N_A_1113_419#_c_1646_n N_CLK_N_c_1779_n 0.00246743f $X=10.245 $Y=2.39
+ $X2=0 $Y2=0
cc_1223 N_A_1113_419#_c_1639_n N_CLK_N_c_1780_n 0.0293702f $X=10.07 $Y=2.225
+ $X2=0 $Y2=0
cc_1224 N_A_1113_419#_c_1646_n N_CLK_N_c_1780_n 0.00321041f $X=10.245 $Y=2.39
+ $X2=0 $Y2=0
cc_1225 N_A_1113_419#_c_1639_n N_CLK_N_c_1781_n 0.00298164f $X=10.07 $Y=2.225
+ $X2=0 $Y2=0
cc_1226 N_A_1113_419#_c_1644_n N_CLK_N_c_1781_n 0.00902255f $X=10.08 $Y=2.095
+ $X2=0 $Y2=0
cc_1227 N_A_1113_419#_c_1646_n N_CLK_N_c_1781_n 0.00151011f $X=10.245 $Y=2.39
+ $X2=0 $Y2=0
cc_1228 N_A_1113_419#_M1037_d N_VPWR_c_2220_n 0.00117463f $X=5.565 $Y=2.095
+ $X2=0 $Y2=0
cc_1229 N_A_1113_419#_M1041_d N_A_305_97#_c_2400_n 0.00176461f $X=5.575 $Y=1.075
+ $X2=0 $Y2=0
cc_1230 N_A_1113_419#_c_1668_n N_A_305_97#_c_2400_n 0.0250761f $X=5.715 $Y=1.36
+ $X2=0 $Y2=0
cc_1231 N_A_1113_419#_c_1668_n N_A_305_97#_c_2403_n 0.00679304f $X=5.715 $Y=1.36
+ $X2=0 $Y2=0
cc_1232 N_A_1113_419#_c_1672_n A_1242_419# 0.0110747f $X=6.735 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_1233 N_A_1113_419#_c_1643_n N_KAPWR_M1010_d 0.00875759f $X=8.07 $Y=2.065
+ $X2=-0.19 $Y2=-0.245
cc_1234 N_A_1113_419#_c_1644_n N_KAPWR_M1014_d 0.00568296f $X=10.08 $Y=2.095
+ $X2=0 $Y2=0
cc_1235 N_A_1113_419#_M1011_s N_KAPWR_c_2590_n 8.41857e-19 $X=7.895 $Y=1.705
+ $X2=0 $Y2=0
cc_1236 N_A_1113_419#_M1029_g N_KAPWR_c_2591_n 0.00117347f $X=9.435 $Y=2.205
+ $X2=0 $Y2=0
cc_1237 N_A_1113_419#_c_1642_n N_KAPWR_c_2593_n 0.0337818f $X=5.767 $Y=2.32
+ $X2=0 $Y2=0
cc_1238 N_A_1113_419#_c_1672_n N_KAPWR_c_2593_n 0.0222028f $X=6.735 $Y=2.405
+ $X2=0 $Y2=0
cc_1239 N_A_1113_419#_c_1643_n N_KAPWR_c_2593_n 0.00731921f $X=8.07 $Y=2.065
+ $X2=0 $Y2=0
cc_1240 N_A_1113_419#_M1011_s N_KAPWR_c_2594_n 0.00205659f $X=7.895 $Y=1.705
+ $X2=0 $Y2=0
cc_1241 N_A_1113_419#_M1029_g N_KAPWR_c_2595_n 0.00244946f $X=9.435 $Y=2.205
+ $X2=0 $Y2=0
cc_1242 N_A_1113_419#_c_1644_n N_KAPWR_c_2595_n 0.013457f $X=10.08 $Y=2.095
+ $X2=0 $Y2=0
cc_1243 N_A_1113_419#_c_1645_n N_KAPWR_c_2595_n 0.00763946f $X=10.245 $Y=2.39
+ $X2=0 $Y2=0
cc_1244 N_A_1113_419#_c_1646_n N_KAPWR_c_2595_n 0.00305416f $X=10.245 $Y=2.39
+ $X2=0 $Y2=0
cc_1245 N_A_1113_419#_c_1644_n A_1682_341# 0.00145127f $X=10.08 $Y=2.095
+ $X2=-0.19 $Y2=-0.245
cc_1246 N_A_1113_419#_c_1634_n N_VGND_c_2833_n 0.0123156f $X=9.125 $Y=0.765
+ $X2=0 $Y2=0
cc_1247 N_A_1113_419#_c_1636_n N_VGND_c_2833_n 0.00235279f $X=9.485 $Y=0.765
+ $X2=0 $Y2=0
cc_1248 N_A_1113_419#_c_1634_n N_VGND_c_2837_n 0.00486043f $X=9.125 $Y=0.765
+ $X2=0 $Y2=0
cc_1249 N_A_1113_419#_c_1636_n N_VGND_c_2837_n 0.00547432f $X=9.485 $Y=0.765
+ $X2=0 $Y2=0
cc_1250 N_A_1113_419#_c_1638_n N_VGND_c_2837_n 5.09538e-19 $X=9.56 $Y=0.99 $X2=0
+ $Y2=0
cc_1251 N_A_1113_419#_c_1634_n N_VGND_c_2845_n 0.00814425f $X=9.125 $Y=0.765
+ $X2=0 $Y2=0
cc_1252 N_A_1113_419#_c_1636_n N_VGND_c_2845_n 0.0112432f $X=9.485 $Y=0.765
+ $X2=0 $Y2=0
cc_1253 N_A_1113_419#_c_1638_n N_VGND_c_2845_n 6.93005e-19 $X=9.56 $Y=0.99 $X2=0
+ $Y2=0
cc_1254 N_A_1113_419#_c_1634_n N_A_1453_77#_c_3077_n 2.87516e-19 $X=9.125
+ $Y=0.765 $X2=0 $Y2=0
cc_1255 N_CLK_N_M1038_g N_SLEEP_B_c_1826_n 0.0345091f $X=10.915 $Y=0.695
+ $X2=-0.19 $Y2=-0.245
cc_1256 N_CLK_N_c_1779_n N_SLEEP_B_M1019_g 0.0332333f $X=11.145 $Y=1.985 $X2=0
+ $Y2=0
cc_1257 N_CLK_N_c_1779_n N_SLEEP_B_c_1831_n 0.0345091f $X=11.145 $Y=1.985 $X2=0
+ $Y2=0
cc_1258 N_CLK_N_M1038_g N_SLEEP_B_c_1833_n 0.00163816f $X=10.915 $Y=0.695 $X2=0
+ $Y2=0
cc_1259 N_CLK_N_c_1779_n N_SLEEP_B_c_1833_n 7.42423e-19 $X=11.145 $Y=1.985 $X2=0
+ $Y2=0
cc_1260 N_CLK_N_c_1779_n N_KAPWR_c_2586_n 0.00400757f $X=11.145 $Y=1.985 $X2=0
+ $Y2=0
cc_1261 N_CLK_N_c_1779_n N_KAPWR_c_2587_n 0.00275107f $X=11.145 $Y=1.985 $X2=0
+ $Y2=0
cc_1262 N_CLK_N_c_1779_n N_KAPWR_c_2592_n 6.7079e-19 $X=11.145 $Y=1.985 $X2=0
+ $Y2=0
cc_1263 N_CLK_N_c_1779_n N_KAPWR_c_2595_n 0.00464942f $X=11.145 $Y=1.985 $X2=0
+ $Y2=0
cc_1264 N_CLK_N_M1038_g N_VGND_c_2837_n 7.35405e-19 $X=10.915 $Y=0.695 $X2=0
+ $Y2=0
cc_1265 N_SLEEP_B_c_1835_n N_VPWR_c_2220_n 2.134e-19 $X=12.15 $Y=1.625 $X2=0
+ $Y2=0
cc_1266 N_SLEEP_B_M1019_g N_KAPWR_c_2587_n 0.00298751f $X=11.575 $Y=2.415 $X2=0
+ $Y2=0
cc_1267 N_SLEEP_B_c_1835_n KAPWR 0.00979592f $X=12.15 $Y=1.625 $X2=0 $Y2=0
cc_1268 N_SLEEP_B_M1019_g N_KAPWR_c_2592_n 0.0143243f $X=11.575 $Y=2.415 $X2=0
+ $Y2=0
cc_1269 N_SLEEP_B_c_1835_n N_KAPWR_c_2592_n 0.0135335f $X=12.15 $Y=1.625 $X2=0
+ $Y2=0
cc_1270 N_SLEEP_B_c_1831_n N_KAPWR_c_2592_n 3.00546e-19 $X=12.4 $Y=1.09 $X2=0
+ $Y2=0
cc_1271 N_SLEEP_B_M1019_g N_KAPWR_c_2595_n 0.00292036f $X=11.575 $Y=2.415 $X2=0
+ $Y2=0
cc_1272 N_SLEEP_B_M1019_g N_KAPWR_c_2659_n 5.14879e-19 $X=11.575 $Y=2.415 $X2=0
+ $Y2=0
cc_1273 N_SLEEP_B_c_1835_n N_A_2562_427#_c_2779_n 0.00259553f $X=12.15 $Y=1.625
+ $X2=0 $Y2=0
cc_1274 N_SLEEP_B_c_1828_n N_VGND_c_2834_n 7.57836e-19 $X=11.665 $Y=1.015 $X2=0
+ $Y2=0
cc_1275 N_SLEEP_B_c_1829_n N_VGND_c_2834_n 9.63362e-19 $X=12.325 $Y=1.015 $X2=0
+ $Y2=0
cc_1276 N_SLEEP_B_c_1826_n N_VGND_c_2837_n 7.35405e-19 $X=11.305 $Y=1.015 $X2=0
+ $Y2=0
cc_1277 N_SLEEP_B_c_1828_n N_VGND_c_2837_n 0.00144978f $X=11.665 $Y=1.015 $X2=0
+ $Y2=0
cc_1278 N_SLEEP_B_c_1829_n N_VGND_c_2842_n 0.0038006f $X=12.325 $Y=1.015 $X2=0
+ $Y2=0
cc_1279 N_SLEEP_B_c_1832_n N_VGND_c_2842_n 7.35405e-19 $X=12.715 $Y=1.015 $X2=0
+ $Y2=0
cc_1280 N_SLEEP_B_c_1828_n N_VGND_c_2845_n 0.00118974f $X=11.665 $Y=1.015 $X2=0
+ $Y2=0
cc_1281 N_SLEEP_B_c_1829_n N_VGND_c_2845_n 0.00509887f $X=12.325 $Y=1.015 $X2=0
+ $Y2=0
cc_1282 N_A_2999_73#_c_1924_n N_A_2717_427#_c_1997_n 9.43567e-19 $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1283 N_A_2999_73#_c_1925_n N_A_2717_427#_c_1997_n 0.00731455f $X=16.22
+ $Y=0.765 $X2=0 $Y2=0
cc_1284 N_A_2999_73#_c_1924_n N_A_2717_427#_c_1998_n 0.00951172f $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1285 N_A_2999_73#_c_1925_n N_A_2717_427#_c_1998_n 0.00116788f $X=16.22
+ $Y=0.765 $X2=0 $Y2=0
cc_1286 N_A_2999_73#_c_1928_n N_A_2717_427#_c_1999_n 2.1846e-19 $X=15.875
+ $Y=1.97 $X2=0 $Y2=0
cc_1287 N_A_2999_73#_c_1931_n N_A_2717_427#_c_1999_n 0.00382177f $X=16.04
+ $Y=1.97 $X2=0 $Y2=0
cc_1288 N_A_2999_73#_c_1929_n N_A_2717_427#_M1046_g 0.014528f $X=16.04 $Y=2.525
+ $X2=0 $Y2=0
cc_1289 N_A_2999_73#_c_1924_n N_A_2717_427#_M1046_g 0.00602636f $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1290 N_A_2999_73#_c_1931_n N_A_2717_427#_M1046_g 0.0133756f $X=16.04 $Y=1.97
+ $X2=0 $Y2=0
cc_1291 N_A_2999_73#_c_1924_n N_A_2717_427#_c_2001_n 0.0011494f $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1292 N_A_2999_73#_c_1931_n N_A_2717_427#_c_2001_n 0.00129166f $X=16.04
+ $Y=1.97 $X2=0 $Y2=0
cc_1293 N_A_2999_73#_M1031_g N_A_2717_427#_c_2023_n 0.0049442f $X=15.395
+ $Y=2.525 $X2=0 $Y2=0
cc_1294 N_A_2999_73#_M1051_g N_A_2717_427#_c_2006_n 0.0229615f $X=15.07 $Y=0.705
+ $X2=0 $Y2=0
cc_1295 N_A_2999_73#_c_1928_n N_A_2717_427#_c_2006_n 0.0121119f $X=15.875
+ $Y=1.97 $X2=0 $Y2=0
cc_1296 N_A_2999_73#_c_1932_n N_A_2717_427#_c_2006_n 0.00579137f $X=15.395
+ $Y=1.97 $X2=0 $Y2=0
cc_1297 N_A_2999_73#_M1051_g N_A_2717_427#_c_2007_n 0.012071f $X=15.07 $Y=0.705
+ $X2=0 $Y2=0
cc_1298 N_A_2999_73#_c_1928_n N_A_2717_427#_c_2007_n 0.0194173f $X=15.875
+ $Y=1.97 $X2=0 $Y2=0
cc_1299 N_A_2999_73#_c_1924_n N_A_2717_427#_c_2007_n 0.0108378f $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1300 N_A_2999_73#_c_1932_n N_A_2717_427#_c_2007_n 0.00591712f $X=15.395
+ $Y=1.97 $X2=0 $Y2=0
cc_1301 N_A_2999_73#_M1051_g N_A_2717_427#_c_2008_n 0.00404451f $X=15.07
+ $Y=0.705 $X2=0 $Y2=0
cc_1302 N_A_2999_73#_c_1924_n N_A_2717_427#_c_2009_n 0.00957046f $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1303 N_A_2999_73#_c_1925_n N_A_2717_427#_c_2009_n 0.0106413f $X=16.22
+ $Y=0.765 $X2=0 $Y2=0
cc_1304 N_A_2999_73#_c_1925_n N_A_2717_427#_c_2010_n 0.0197592f $X=16.22
+ $Y=0.765 $X2=0 $Y2=0
cc_1305 N_A_2999_73#_c_1924_n N_A_2717_427#_c_2012_n 0.0309558f $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1306 N_A_2999_73#_c_1928_n N_A_2717_427#_c_2025_n 0.01334f $X=15.875 $Y=1.97
+ $X2=0 $Y2=0
cc_1307 N_A_2999_73#_c_1932_n N_A_2717_427#_c_2025_n 0.007234f $X=15.395 $Y=1.97
+ $X2=0 $Y2=0
cc_1308 N_A_2999_73#_c_1925_n N_A_2717_427#_c_2013_n 0.025445f $X=16.22 $Y=0.765
+ $X2=0 $Y2=0
cc_1309 N_A_2999_73#_c_1924_n N_A_2717_427#_c_2014_n 0.0161974f $X=16.12
+ $Y=1.805 $X2=0 $Y2=0
cc_1310 N_A_2999_73#_c_1925_n N_A_2717_427#_c_2014_n 0.00531173f $X=16.22
+ $Y=0.765 $X2=0 $Y2=0
cc_1311 N_A_2999_73#_M1031_g N_VPWR_c_2224_n 0.00749759f $X=15.395 $Y=2.525
+ $X2=0 $Y2=0
cc_1312 N_A_2999_73#_c_1928_n N_VPWR_c_2224_n 0.0208418f $X=15.875 $Y=1.97 $X2=0
+ $Y2=0
cc_1313 N_A_2999_73#_c_1929_n N_VPWR_c_2224_n 0.0177248f $X=16.04 $Y=2.525 $X2=0
+ $Y2=0
cc_1314 N_A_2999_73#_c_1932_n N_VPWR_c_2224_n 0.0016307f $X=15.395 $Y=1.97 $X2=0
+ $Y2=0
cc_1315 N_A_2999_73#_c_1929_n N_VPWR_c_2225_n 0.0184663f $X=16.04 $Y=2.525 $X2=0
+ $Y2=0
cc_1316 N_A_2999_73#_c_1929_n N_VPWR_c_2233_n 0.00753442f $X=16.04 $Y=2.525
+ $X2=0 $Y2=0
cc_1317 N_A_2999_73#_c_1929_n N_VPWR_c_2220_n 0.00110772f $X=16.04 $Y=2.525
+ $X2=0 $Y2=0
cc_1318 N_A_2999_73#_M1031_g KAPWR 0.00410062f $X=15.395 $Y=2.525 $X2=0 $Y2=0
cc_1319 N_A_2999_73#_c_1928_n KAPWR 0.0120972f $X=15.875 $Y=1.97 $X2=0 $Y2=0
cc_1320 N_A_2999_73#_c_1929_n KAPWR 0.0278727f $X=16.04 $Y=2.525 $X2=0 $Y2=0
cc_1321 N_A_2999_73#_c_1932_n KAPWR 0.00362046f $X=15.395 $Y=1.97 $X2=0 $Y2=0
cc_1322 N_A_2999_73#_M1031_g N_A_2562_427#_c_2782_n 0.00330488f $X=15.395
+ $Y=2.525 $X2=0 $Y2=0
cc_1323 N_A_2999_73#_c_1928_n N_A_2562_427#_c_2782_n 0.00443155f $X=15.875
+ $Y=1.97 $X2=0 $Y2=0
cc_1324 N_A_2999_73#_c_1932_n N_A_2562_427#_c_2782_n 0.00651754f $X=15.395
+ $Y=1.97 $X2=0 $Y2=0
cc_1325 N_A_2999_73#_M1051_g N_VGND_c_2835_n 0.011731f $X=15.07 $Y=0.705 $X2=0
+ $Y2=0
cc_1326 N_A_2999_73#_M1051_g N_VGND_c_2842_n 0.00407914f $X=15.07 $Y=0.705 $X2=0
+ $Y2=0
cc_1327 N_A_2999_73#_M1051_g N_VGND_c_2845_n 0.00425776f $X=15.07 $Y=0.705 $X2=0
+ $Y2=0
cc_1328 N_A_2717_427#_M1036_g N_A_3368_57#_M1033_g 0.0140011f $X=17.2 $Y=0.495
+ $X2=0 $Y2=0
cc_1329 N_A_2717_427#_c_2017_n N_A_3368_57#_M1024_g 0.022623f $X=17.145 $Y=1.96
+ $X2=0 $Y2=0
cc_1330 N_A_2717_427#_c_2014_n N_A_3368_57#_c_2158_n 0.0068075f $X=16.502 $Y=1.1
+ $X2=0 $Y2=0
cc_1331 N_A_2717_427#_c_2017_n N_A_3368_57#_c_2166_n 0.00440904f $X=17.145
+ $Y=1.96 $X2=0 $Y2=0
cc_1332 N_A_2717_427#_M1047_g N_A_3368_57#_c_2166_n 0.00436686f $X=17.22
+ $Y=2.775 $X2=0 $Y2=0
cc_1333 N_A_2717_427#_M1047_g N_A_3368_57#_c_2167_n 0.00701467f $X=17.22
+ $Y=2.775 $X2=0 $Y2=0
cc_1334 N_A_2717_427#_c_2002_n N_A_3368_57#_c_2160_n 0.0131916f $X=17.125
+ $Y=0.97 $X2=0 $Y2=0
cc_1335 N_A_2717_427#_M1036_g N_A_3368_57#_c_2160_n 0.00481865f $X=17.2 $Y=0.495
+ $X2=0 $Y2=0
cc_1336 N_A_2717_427#_c_2012_n N_A_3368_57#_c_2160_n 0.0309302f $X=16.645
+ $Y=1.06 $X2=0 $Y2=0
cc_1337 N_A_2717_427#_c_2013_n N_A_3368_57#_c_2160_n 0.00804039f $X=16.645
+ $Y=0.895 $X2=0 $Y2=0
cc_1338 N_A_2717_427#_c_2014_n N_A_3368_57#_c_2160_n 0.00474061f $X=16.502
+ $Y=1.1 $X2=0 $Y2=0
cc_1339 N_A_2717_427#_c_2002_n N_A_3368_57#_c_2161_n 0.00416697f $X=17.125
+ $Y=0.97 $X2=0 $Y2=0
cc_1340 N_A_2717_427#_c_2017_n N_A_3368_57#_c_2161_n 0.00512525f $X=17.145
+ $Y=1.96 $X2=0 $Y2=0
cc_1341 N_A_2717_427#_M1036_g N_A_3368_57#_c_2162_n 0.00683105f $X=17.2 $Y=0.495
+ $X2=0 $Y2=0
cc_1342 N_A_2717_427#_c_2010_n N_A_3368_57#_c_2162_n 0.0141537f $X=16.48 $Y=0.34
+ $X2=0 $Y2=0
cc_1343 N_A_2717_427#_c_2013_n N_A_3368_57#_c_2162_n 0.0237477f $X=16.645
+ $Y=0.895 $X2=0 $Y2=0
cc_1344 N_A_2717_427#_c_2014_n N_A_3368_57#_c_2162_n 0.00617466f $X=16.502
+ $Y=1.1 $X2=0 $Y2=0
cc_1345 N_A_2717_427#_M1046_g N_A_3368_57#_c_2163_n 0.00767267f $X=16.255
+ $Y=2.525 $X2=0 $Y2=0
cc_1346 N_A_2717_427#_c_2001_n N_A_3368_57#_c_2163_n 0.00527014f $X=16.75
+ $Y=1.885 $X2=0 $Y2=0
cc_1347 N_A_2717_427#_c_2017_n N_A_3368_57#_c_2163_n 0.0153246f $X=17.145
+ $Y=1.96 $X2=0 $Y2=0
cc_1348 N_A_2717_427#_M1047_g N_A_3368_57#_c_2163_n 0.0114836f $X=17.22 $Y=2.775
+ $X2=0 $Y2=0
cc_1349 N_A_2717_427#_c_2002_n N_A_3368_57#_c_2164_n 8.69385e-19 $X=17.125
+ $Y=0.97 $X2=0 $Y2=0
cc_1350 N_A_2717_427#_c_2012_n N_A_3368_57#_c_2164_n 0.020991f $X=16.645 $Y=1.06
+ $X2=0 $Y2=0
cc_1351 N_A_2717_427#_c_2014_n N_A_3368_57#_c_2164_n 0.00498654f $X=16.502
+ $Y=1.1 $X2=0 $Y2=0
cc_1352 N_A_2717_427#_M1046_g N_VPWR_c_2225_n 0.00517795f $X=16.255 $Y=2.525
+ $X2=0 $Y2=0
cc_1353 N_A_2717_427#_M1047_g N_VPWR_c_2225_n 0.00444034f $X=17.22 $Y=2.775
+ $X2=0 $Y2=0
cc_1354 N_A_2717_427#_c_2017_n N_VPWR_c_2226_n 0.0134605f $X=17.145 $Y=1.96
+ $X2=0 $Y2=0
cc_1355 N_A_2717_427#_M1046_g N_VPWR_c_2233_n 0.00294013f $X=16.255 $Y=2.525
+ $X2=0 $Y2=0
cc_1356 N_A_2717_427#_M1047_g N_VPWR_c_2236_n 0.0054895f $X=17.22 $Y=2.775 $X2=0
+ $Y2=0
cc_1357 N_A_2717_427#_M1046_g N_VPWR_c_2220_n 8.07163e-19 $X=16.255 $Y=2.525
+ $X2=0 $Y2=0
cc_1358 N_A_2717_427#_M1047_g N_VPWR_c_2220_n 0.00692684f $X=17.22 $Y=2.775
+ $X2=0 $Y2=0
cc_1359 N_A_2717_427#_M1046_g KAPWR 0.00994481f $X=16.255 $Y=2.525 $X2=0 $Y2=0
cc_1360 N_A_2717_427#_c_2018_n KAPWR 0.00372991f $X=16.825 $Y=1.96 $X2=0 $Y2=0
cc_1361 N_A_2717_427#_M1047_g KAPWR 0.00852607f $X=17.22 $Y=2.775 $X2=0 $Y2=0
cc_1362 N_A_2717_427#_c_2021_n KAPWR 0.0463576f $X=14.755 $Y=2.65 $X2=0 $Y2=0
cc_1363 N_A_2717_427#_c_2022_n KAPWR 0.0196794f $X=13.905 $Y=2.65 $X2=0 $Y2=0
cc_1364 N_A_2717_427#_c_2025_n KAPWR 0.00413317f $X=14.955 $Y=2.05 $X2=0 $Y2=0
cc_1365 N_A_2717_427#_c_2005_n N_A_2562_427#_c_2779_n 0.00960597f $X=13.82
+ $Y=1.86 $X2=0 $Y2=0
cc_1366 N_A_2717_427#_c_2022_n N_A_2562_427#_c_2779_n 0.00495027f $X=13.905
+ $Y=2.65 $X2=0 $Y2=0
cc_1367 N_A_2717_427#_c_2021_n N_A_2562_427#_c_2780_n 0.0721995f $X=14.755
+ $Y=2.65 $X2=0 $Y2=0
cc_1368 N_A_2717_427#_c_2022_n N_A_2562_427#_c_2780_n 0.0181362f $X=13.905
+ $Y=2.65 $X2=0 $Y2=0
cc_1369 N_A_2717_427#_c_2021_n N_A_2562_427#_c_2782_n 0.0134475f $X=14.755
+ $Y=2.65 $X2=0 $Y2=0
cc_1370 N_A_2717_427#_c_2023_n N_A_2562_427#_c_2782_n 0.0192066f $X=14.84
+ $Y=2.565 $X2=0 $Y2=0
cc_1371 N_A_2717_427#_c_1997_n N_VGND_c_2835_n 2.08046e-19 $X=15.89 $Y=1.025
+ $X2=0 $Y2=0
cc_1372 N_A_2717_427#_c_2007_n N_VGND_c_2835_n 0.0273053f $X=15.62 $Y=1.19 $X2=0
+ $Y2=0
cc_1373 N_A_2717_427#_c_2009_n N_VGND_c_2835_n 0.0224097f $X=15.705 $Y=1.105
+ $X2=0 $Y2=0
cc_1374 N_A_2717_427#_c_2011_n N_VGND_c_2835_n 0.01479f $X=15.79 $Y=0.34 $X2=0
+ $Y2=0
cc_1375 N_A_2717_427#_M1036_g N_VGND_c_2836_n 0.00957493f $X=17.2 $Y=0.495 $X2=0
+ $Y2=0
cc_1376 N_A_2717_427#_c_1997_n N_VGND_c_2843_n 7.17276e-19 $X=15.89 $Y=1.025
+ $X2=0 $Y2=0
cc_1377 N_A_2717_427#_M1036_g N_VGND_c_2843_n 0.00502664f $X=17.2 $Y=0.495 $X2=0
+ $Y2=0
cc_1378 N_A_2717_427#_c_2010_n N_VGND_c_2843_n 0.0565771f $X=16.48 $Y=0.34 $X2=0
+ $Y2=0
cc_1379 N_A_2717_427#_c_2011_n N_VGND_c_2843_n 0.0121867f $X=15.79 $Y=0.34 $X2=0
+ $Y2=0
cc_1380 N_A_2717_427#_M1036_g N_VGND_c_2845_n 0.0106059f $X=17.2 $Y=0.495 $X2=0
+ $Y2=0
cc_1381 N_A_2717_427#_c_2010_n N_VGND_c_2845_n 0.0325436f $X=16.48 $Y=0.34 $X2=0
+ $Y2=0
cc_1382 N_A_2717_427#_c_2011_n N_VGND_c_2845_n 0.00660921f $X=15.79 $Y=0.34
+ $X2=0 $Y2=0
cc_1383 N_A_2717_427#_c_2009_n A_3115_99# 0.00218706f $X=15.705 $Y=1.105
+ $X2=-0.19 $Y2=-0.245
cc_1384 N_A_3368_57#_c_2166_n N_VPWR_c_2225_n 0.0425257f $X=17.005 $Y=2.6 $X2=0
+ $Y2=0
cc_1385 N_A_3368_57#_c_2163_n N_VPWR_c_2225_n 0.00668737f $X=17.005 $Y=2.435
+ $X2=0 $Y2=0
cc_1386 N_A_3368_57#_M1024_g N_VPWR_c_2226_n 0.00474211f $X=17.755 $Y=2.465
+ $X2=0 $Y2=0
cc_1387 N_A_3368_57#_c_2158_n N_VPWR_c_2226_n 0.00577732f $X=17.67 $Y=1.48 $X2=0
+ $Y2=0
cc_1388 N_A_3368_57#_c_2161_n N_VPWR_c_2226_n 0.0209147f $X=17.46 $Y=1.48 $X2=0
+ $Y2=0
cc_1389 N_A_3368_57#_c_2163_n N_VPWR_c_2226_n 0.0795154f $X=17.005 $Y=2.435
+ $X2=0 $Y2=0
cc_1390 N_A_3368_57#_c_2167_n N_VPWR_c_2236_n 0.0210218f $X=17.005 $Y=2.755
+ $X2=0 $Y2=0
cc_1391 N_A_3368_57#_M1024_g N_VPWR_c_2237_n 0.00533769f $X=17.755 $Y=2.465
+ $X2=0 $Y2=0
cc_1392 N_A_3368_57#_M1047_s N_VPWR_c_2220_n 0.00115393f $X=16.87 $Y=2.455 $X2=0
+ $Y2=0
cc_1393 N_A_3368_57#_M1024_g N_VPWR_c_2220_n 0.00620599f $X=17.755 $Y=2.465
+ $X2=0 $Y2=0
cc_1394 N_A_3368_57#_c_2167_n N_VPWR_c_2220_n 0.00304772f $X=17.005 $Y=2.755
+ $X2=0 $Y2=0
cc_1395 N_A_3368_57#_M1024_g KAPWR 0.00639997f $X=17.755 $Y=2.465 $X2=0 $Y2=0
cc_1396 N_A_3368_57#_c_2167_n KAPWR 0.0291035f $X=17.005 $Y=2.755 $X2=0 $Y2=0
cc_1397 N_A_3368_57#_M1033_g N_Q_c_2814_n 0.0206781f $X=17.745 $Y=0.705 $X2=0
+ $Y2=0
cc_1398 N_A_3368_57#_M1024_g N_Q_c_2814_n 0.0237754f $X=17.755 $Y=2.465 $X2=0
+ $Y2=0
cc_1399 N_A_3368_57#_c_2159_n N_Q_c_2814_n 0.0125833f $X=17.75 $Y=1.48 $X2=0
+ $Y2=0
cc_1400 N_A_3368_57#_c_2160_n N_Q_c_2814_n 0.00460418f $X=17.065 $Y=1.315 $X2=0
+ $Y2=0
cc_1401 N_A_3368_57#_c_2161_n N_Q_c_2814_n 0.0261285f $X=17.46 $Y=1.48 $X2=0
+ $Y2=0
cc_1402 N_A_3368_57#_c_2163_n N_Q_c_2814_n 0.00476989f $X=17.005 $Y=2.435 $X2=0
+ $Y2=0
cc_1403 N_A_3368_57#_M1033_g N_VGND_c_2836_n 0.0040812f $X=17.745 $Y=0.705 $X2=0
+ $Y2=0
cc_1404 N_A_3368_57#_c_2158_n N_VGND_c_2836_n 0.00577732f $X=17.67 $Y=1.48 $X2=0
+ $Y2=0
cc_1405 N_A_3368_57#_c_2161_n N_VGND_c_2836_n 0.0209147f $X=17.46 $Y=1.48 $X2=0
+ $Y2=0
cc_1406 N_A_3368_57#_c_2162_n N_VGND_c_2836_n 0.0555785f $X=16.985 $Y=0.495
+ $X2=0 $Y2=0
cc_1407 N_A_3368_57#_c_2162_n N_VGND_c_2843_n 0.0217243f $X=16.985 $Y=0.495
+ $X2=0 $Y2=0
cc_1408 N_A_3368_57#_M1033_g N_VGND_c_2844_n 0.00502664f $X=17.745 $Y=0.705
+ $X2=0 $Y2=0
cc_1409 N_A_3368_57#_M1033_g N_VGND_c_2845_n 0.0102688f $X=17.745 $Y=0.705 $X2=0
+ $Y2=0
cc_1410 N_A_3368_57#_c_2162_n N_VGND_c_2845_n 0.0125174f $X=16.985 $Y=0.495
+ $X2=0 $Y2=0
cc_1411 N_VPWR_c_2220_n A_247_491# 0.00194712f $X=18 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1412 N_VPWR_c_2220_n N_A_305_97#_M1026_d 0.00114239f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1413 N_VPWR_c_2221_n N_A_305_97#_c_2415_n 0.0103595f $X=0.945 $Y=2.6 $X2=0
+ $Y2=0
cc_1414 N_VPWR_c_2229_n N_A_305_97#_c_2415_n 0.0189058f $X=2.67 $Y=3.33 $X2=0
+ $Y2=0
cc_1415 N_VPWR_c_2220_n N_A_305_97#_c_2415_n 0.00300491f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1416 N_VPWR_M1052_d N_A_305_97#_c_2404_n 0.00346753f $X=2.695 $Y=2.455 $X2=0
+ $Y2=0
cc_1417 N_VPWR_c_2222_n N_A_305_97#_c_2404_n 0.0131931f $X=2.835 $Y=2.95 $X2=0
+ $Y2=0
cc_1418 N_VPWR_c_2229_n N_A_305_97#_c_2404_n 0.00856086f $X=2.67 $Y=3.33 $X2=0
+ $Y2=0
cc_1419 N_VPWR_c_2231_n N_A_305_97#_c_2404_n 0.00152246f $X=4.285 $Y=3.33 $X2=0
+ $Y2=0
cc_1420 N_VPWR_c_2221_n N_A_305_97#_c_2405_n 0.00571183f $X=0.945 $Y=2.6 $X2=0
+ $Y2=0
cc_1421 N_VPWR_c_2222_n N_A_305_97#_c_2407_n 0.00836003f $X=2.835 $Y=2.95 $X2=0
+ $Y2=0
cc_1422 N_VPWR_c_2223_n N_A_305_97#_c_2408_n 0.0138815f $X=4.37 $Y=2.24 $X2=0
+ $Y2=0
cc_1423 N_VPWR_c_2231_n N_A_305_97#_c_2408_n 0.0552209f $X=4.285 $Y=3.33 $X2=0
+ $Y2=0
cc_1424 N_VPWR_c_2220_n N_A_305_97#_c_2408_n 0.00678137f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1425 N_VPWR_c_2222_n N_A_305_97#_c_2409_n 0.0139672f $X=2.835 $Y=2.95 $X2=0
+ $Y2=0
cc_1426 N_VPWR_c_2231_n N_A_305_97#_c_2409_n 0.0121661f $X=4.285 $Y=3.33 $X2=0
+ $Y2=0
cc_1427 N_VPWR_c_2220_n N_A_305_97#_c_2409_n 0.0015936f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1428 N_VPWR_M1021_d N_A_305_97#_c_2410_n 0.0168682f $X=3.86 $Y=2.095 $X2=0
+ $Y2=0
cc_1429 N_VPWR_c_2223_n N_A_305_97#_c_2410_n 0.0594917f $X=4.37 $Y=2.24 $X2=0
+ $Y2=0
cc_1430 N_VPWR_c_2223_n N_A_305_97#_c_2396_n 0.0111887f $X=4.37 $Y=2.24 $X2=0
+ $Y2=0
cc_1431 N_VPWR_c_2235_n N_A_305_97#_c_2411_n 0.00762486f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1432 N_VPWR_c_2220_n N_A_305_97#_c_2411_n 9.33528e-19 $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1433 N_VPWR_c_2231_n N_A_305_97#_c_2412_n 7.07575e-19 $X=4.285 $Y=3.33 $X2=0
+ $Y2=0
cc_1434 N_VPWR_c_2223_n N_A_305_97#_c_2413_n 0.0261915f $X=4.37 $Y=2.24 $X2=0
+ $Y2=0
cc_1435 N_VPWR_c_2220_n A_411_491# 0.00281409f $X=18 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1436 N_VPWR_c_2220_n A_1242_419# 0.00215342f $X=18 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1437 N_VPWR_c_2220_n N_KAPWR_M1010_d 0.00314054f $X=18 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1438 N_VPWR_c_2235_n N_KAPWR_c_2587_n 0.0681214f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1439 N_VPWR_c_2220_n N_KAPWR_c_2587_n 0.00818404f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1440 N_VPWR_c_2235_n N_KAPWR_c_2588_n 0.0115893f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1441 N_VPWR_c_2220_n N_KAPWR_c_2588_n 0.00141402f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1442 N_VPWR_M1031_d KAPWR 6.93765e-19 $X=15.47 $Y=2.315 $X2=0 $Y2=0
cc_1443 N_VPWR_M1046_d KAPWR 0.0021453f $X=16.33 $Y=2.315 $X2=0 $Y2=0
cc_1444 N_VPWR_M1047_d KAPWR 0.00611632f $X=17.295 $Y=2.455 $X2=0 $Y2=0
cc_1445 N_VPWR_c_2224_n KAPWR 0.0256535f $X=15.61 $Y=2.53 $X2=0 $Y2=0
cc_1446 N_VPWR_c_2225_n KAPWR 0.0338613f $X=16.47 $Y=2.525 $X2=0 $Y2=0
cc_1447 N_VPWR_c_2226_n KAPWR 0.0305691f $X=17.54 $Y=1.98 $X2=0 $Y2=0
cc_1448 N_VPWR_c_2233_n KAPWR 0.00287988f $X=16.385 $Y=3.33 $X2=0 $Y2=0
cc_1449 N_VPWR_c_2235_n KAPWR 0.00573463f $X=15.445 $Y=3.33 $X2=0 $Y2=0
cc_1450 N_VPWR_c_2236_n KAPWR 0.00238178f $X=17.375 $Y=3.33 $X2=0 $Y2=0
cc_1451 N_VPWR_c_2237_n KAPWR 0.00128789f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1452 N_VPWR_c_2235_n N_KAPWR_c_2590_n 0.0420664f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1453 N_VPWR_c_2220_n N_KAPWR_c_2590_n 0.0054843f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1454 N_VPWR_c_2235_n N_KAPWR_c_2591_n 0.0475137f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1455 N_VPWR_c_2220_n N_KAPWR_c_2591_n 0.00800923f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1456 N_VPWR_M1016_d N_KAPWR_c_2593_n 8.0097e-19 $X=0.735 $Y=2.455 $X2=0 $Y2=0
cc_1457 N_VPWR_M1052_d N_KAPWR_c_2593_n 0.00252562f $X=2.695 $Y=2.455 $X2=0
+ $Y2=0
cc_1458 N_VPWR_M1021_d N_KAPWR_c_2593_n 0.0125885f $X=3.86 $Y=2.095 $X2=0 $Y2=0
cc_1459 N_VPWR_c_2221_n N_KAPWR_c_2593_n 0.0287558f $X=0.945 $Y=2.6 $X2=0 $Y2=0
cc_1460 N_VPWR_c_2222_n N_KAPWR_c_2593_n 0.0149168f $X=2.835 $Y=2.95 $X2=0 $Y2=0
cc_1461 N_VPWR_c_2223_n N_KAPWR_c_2593_n 0.0267419f $X=4.37 $Y=2.24 $X2=0 $Y2=0
cc_1462 N_VPWR_c_2227_n N_KAPWR_c_2593_n 0.00139837f $X=0.78 $Y=3.33 $X2=0 $Y2=0
cc_1463 N_VPWR_c_2229_n N_KAPWR_c_2593_n 0.00508663f $X=2.67 $Y=3.33 $X2=0 $Y2=0
cc_1464 N_VPWR_c_2231_n N_KAPWR_c_2593_n 0.00214705f $X=4.285 $Y=3.33 $X2=0
+ $Y2=0
cc_1465 N_VPWR_c_2235_n N_KAPWR_c_2593_n 0.0059229f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1466 N_VPWR_c_2220_n N_KAPWR_c_2593_n 1.88996f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1467 N_VPWR_c_2235_n N_KAPWR_c_2594_n 0.0020449f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1468 N_VPWR_c_2235_n N_KAPWR_c_2595_n 0.0061641f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1469 N_VPWR_c_2224_n N_A_2562_427#_c_2780_n 0.0135846f $X=15.61 $Y=2.53 $X2=0
+ $Y2=0
cc_1470 N_VPWR_c_2235_n N_A_2562_427#_c_2780_n 0.140002f $X=15.445 $Y=3.33 $X2=0
+ $Y2=0
cc_1471 N_VPWR_c_2220_n N_A_2562_427#_c_2780_n 0.0166801f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1472 N_VPWR_c_2235_n N_A_2562_427#_c_2781_n 0.0224969f $X=15.445 $Y=3.33
+ $X2=0 $Y2=0
cc_1473 N_VPWR_c_2220_n N_A_2562_427#_c_2781_n 0.00274486f $X=18 $Y=3.33 $X2=0
+ $Y2=0
cc_1474 N_VPWR_c_2224_n N_A_2562_427#_c_2782_n 0.0268003f $X=15.61 $Y=2.53 $X2=0
+ $Y2=0
cc_1475 N_VPWR_c_2220_n N_Q_M1024_d 0.00114985f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1476 N_VPWR_c_2226_n N_Q_c_2814_n 0.0517063f $X=17.54 $Y=1.98 $X2=0 $Y2=0
cc_1477 N_VPWR_c_2237_n N_Q_c_2814_n 0.0217146f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1478 N_VPWR_c_2220_n N_Q_c_2814_n 0.00312179f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1479 A_247_491# N_KAPWR_c_2593_n 0.00436893f $X=1.235 $Y=2.455 $X2=0.78
+ $Y2=3.33
cc_1480 N_A_305_97#_c_2404_n A_411_491# 0.00723448f $X=3.04 $Y=2.53 $X2=-0.19
+ $Y2=-0.245
cc_1481 N_A_305_97#_c_2415_n N_KAPWR_c_2593_n 0.0315476f $X=1.765 $Y=2.76 $X2=0
+ $Y2=0
cc_1482 N_A_305_97#_c_2404_n N_KAPWR_c_2593_n 0.0404149f $X=3.04 $Y=2.53 $X2=0
+ $Y2=0
cc_1483 N_A_305_97#_c_2407_n N_KAPWR_c_2593_n 0.0248396f $X=3.175 $Y=2.905 $X2=0
+ $Y2=0
cc_1484 N_A_305_97#_c_2408_n N_KAPWR_c_2593_n 0.0246924f $X=3.945 $Y=2.99 $X2=0
+ $Y2=0
cc_1485 N_A_305_97#_c_2409_n N_KAPWR_c_2593_n 0.00253288f $X=3.26 $Y=2.99 $X2=0
+ $Y2=0
cc_1486 N_A_305_97#_c_2410_n N_KAPWR_c_2593_n 0.0224956f $X=4.03 $Y=2.905 $X2=0
+ $Y2=0
cc_1487 N_A_305_97#_c_2411_n N_KAPWR_c_2593_n 0.0281754f $X=4.8 $Y=2.43 $X2=0
+ $Y2=0
cc_1488 N_A_305_97#_c_2412_n N_KAPWR_c_2593_n 0.0021304f $X=3.15 $Y=2.53 $X2=0
+ $Y2=0
cc_1489 N_A_305_97#_c_2391_n N_noxref_30_c_2991_n 0.0137808f $X=1.975 $Y=0.76
+ $X2=0 $Y2=0
cc_1490 N_A_305_97#_c_2391_n N_noxref_30_c_2992_n 0.0402451f $X=1.975 $Y=0.76
+ $X2=0 $Y2=0
cc_1491 N_A_305_97#_c_2391_n noxref_31 0.00138213f $X=1.975 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_1492 N_A_305_97#_c_2391_n N_noxref_32_c_3021_n 0.00117269f $X=1.975 $Y=0.76
+ $X2=0 $Y2=0
cc_1493 N_A_305_97#_c_2393_n N_noxref_32_c_3022_n 0.0484785f $X=3.04 $Y=1.35
+ $X2=0 $Y2=0
cc_1494 N_A_305_97#_c_2396_n N_noxref_32_c_3022_n 0.00713749f $X=4.635 $Y=1.82
+ $X2=0 $Y2=0
cc_1495 N_A_305_97#_c_2397_n N_noxref_32_c_3022_n 0.00568183f $X=4.115 $Y=1.82
+ $X2=0 $Y2=0
cc_1496 N_A_305_97#_c_2392_n N_noxref_32_c_3023_n 0.010763f $X=2.06 $Y=1.265
+ $X2=0 $Y2=0
cc_1497 N_A_305_97#_c_2393_n N_noxref_32_c_3023_n 0.0140042f $X=3.04 $Y=1.35
+ $X2=0 $Y2=0
cc_1498 N_A_305_97#_c_2396_n N_noxref_32_c_3024_n 0.00796732f $X=4.635 $Y=1.82
+ $X2=0 $Y2=0
cc_1499 N_A_305_97#_c_2461_n N_noxref_32_c_3024_n 0.00556983f $X=4.805 $Y=1.35
+ $X2=0 $Y2=0
cc_1500 N_A_305_97#_c_2401_n N_noxref_32_c_3024_n 0.00625201f $X=5.38 $Y=1.02
+ $X2=0 $Y2=0
cc_1501 N_A_305_97#_c_2399_n N_A_1009_107#_M1041_s 0.00779325f $X=5.21 $Y=1.35
+ $X2=-0.19 $Y2=-0.245
cc_1502 N_A_305_97#_c_2463_n N_A_1009_107#_M1041_s 0.00228537f $X=5.295 $Y=1.265
+ $X2=-0.19 $Y2=-0.245
cc_1503 N_A_305_97#_c_2401_n N_A_1009_107#_M1041_s 0.00395797f $X=5.38 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_1504 N_A_305_97#_c_2399_n N_A_1009_107#_c_3056_n 0.00644517f $X=5.21 $Y=1.35
+ $X2=0 $Y2=0
cc_1505 N_A_305_97#_c_2400_n N_A_1009_107#_c_3056_n 0.0722448f $X=6.34 $Y=1.02
+ $X2=0 $Y2=0
cc_1506 N_A_305_97#_c_2401_n N_A_1009_107#_c_3056_n 0.0136855f $X=5.38 $Y=1.02
+ $X2=0 $Y2=0
cc_1507 N_A_305_97#_c_2403_n N_A_1009_107#_c_3056_n 0.0262786f $X=6.505 $Y=1.02
+ $X2=0 $Y2=0
cc_1508 N_A_305_97#_c_2400_n A_1201_215# 0.00290409f $X=6.34 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_1509 A_411_491# N_KAPWR_c_2593_n 0.0073577f $X=2.055 $Y=2.455 $X2=0.78
+ $Y2=3.33
cc_1510 A_1242_419# N_KAPWR_c_2593_n 0.00466677f $X=6.21 $Y=2.095 $X2=13.74
+ $Y2=1.1
cc_1511 N_KAPWR_c_2591_n A_1682_341# 4.51141e-19 $X=9.075 $Y=2.855 $X2=-0.19
+ $Y2=1.655
cc_1512 N_KAPWR_c_2594_n A_1682_341# 0.00120124f $X=8.545 $Y=2.81 $X2=-0.19
+ $Y2=1.655
cc_1513 N_KAPWR_c_2595_n A_1682_341# 6.12362e-19 $X=11.615 $Y=2.802 $X2=-0.19
+ $Y2=1.655
cc_1514 KAPWR N_A_2562_427#_M1031_s 0.00181385f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1515 KAPWR N_A_2562_427#_c_2779_n 0.0285525f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1516 KAPWR N_A_2562_427#_c_2780_n 0.0607205f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1517 KAPWR N_A_2562_427#_c_2781_n 0.00552945f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1518 KAPWR N_A_2562_427#_c_2782_n 0.0171944f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1519 KAPWR N_Q_c_2814_n 0.039908f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1520 N_Q_c_2814_n N_VGND_c_2836_n 0.0331408f $X=17.96 $Y=0.43 $X2=0 $Y2=0
cc_1521 N_Q_c_2814_n N_VGND_c_2844_n 0.0227064f $X=17.96 $Y=0.43 $X2=0 $Y2=0
cc_1522 N_Q_c_2814_n N_VGND_c_2845_n 0.0129677f $X=17.96 $Y=0.43 $X2=0 $Y2=0
cc_1523 N_VGND_c_2830_n N_noxref_30_c_2991_n 0.0207056f $X=0.7 $Y=0.485 $X2=0
+ $Y2=0
cc_1524 N_VGND_c_2840_n N_noxref_30_c_2992_n 0.092089f $X=3.835 $Y=0 $X2=0 $Y2=0
cc_1525 N_VGND_c_2845_n N_noxref_30_c_2992_n 0.0537609f $X=18 $Y=0 $X2=0 $Y2=0
cc_1526 N_VGND_c_2830_n N_noxref_30_c_2993_n 0.0131778f $X=0.7 $Y=0.485 $X2=0
+ $Y2=0
cc_1527 N_VGND_c_2840_n N_noxref_30_c_2993_n 0.0179017f $X=3.835 $Y=0 $X2=0
+ $Y2=0
cc_1528 N_VGND_c_2845_n N_noxref_30_c_2993_n 0.00971565f $X=18 $Y=0 $X2=0 $Y2=0
cc_1529 N_VGND_c_2840_n N_noxref_30_c_2994_n 0.0229767f $X=3.835 $Y=0 $X2=0
+ $Y2=0
cc_1530 N_VGND_c_2845_n N_noxref_30_c_2994_n 0.0126513f $X=18 $Y=0 $X2=0 $Y2=0
cc_1531 N_VGND_M1018_d N_noxref_32_c_3022_n 0.00286307f $X=3.86 $Y=0.445 $X2=0
+ $Y2=0
cc_1532 N_VGND_c_2831_n N_noxref_32_c_3022_n 0.0241405f $X=4 $Y=0.59 $X2=0 $Y2=0
cc_1533 N_VGND_c_2831_n N_noxref_32_c_3024_n 0.010785f $X=4 $Y=0.59 $X2=0 $Y2=0
cc_1534 N_VGND_c_2841_n N_noxref_32_c_3024_n 0.00498848f $X=7.78 $Y=0 $X2=0
+ $Y2=0
cc_1535 N_VGND_c_2845_n N_noxref_32_c_3024_n 0.00742854f $X=18 $Y=0 $X2=0 $Y2=0
cc_1536 N_VGND_c_2845_n N_A_1453_77#_M1007_d 0.00225167f $X=18 $Y=0 $X2=0 $Y2=0
cc_1537 N_VGND_M1007_s N_A_1453_77#_c_3075_n 0.00465618f $X=7.81 $Y=0.135 $X2=0
+ $Y2=0
cc_1538 N_VGND_c_2832_n N_A_1453_77#_c_3075_n 0.00385152f $X=8.825 $Y=0 $X2=0
+ $Y2=0
cc_1539 N_VGND_c_2841_n N_A_1453_77#_c_3075_n 0.00480994f $X=7.78 $Y=0 $X2=0
+ $Y2=0
cc_1540 N_VGND_c_2845_n N_A_1453_77#_c_3075_n 0.0140696f $X=18 $Y=0 $X2=0 $Y2=0
cc_1541 N_VGND_c_2848_n N_A_1453_77#_c_3075_n 0.0242212f $X=7.92 $Y=0 $X2=0
+ $Y2=0
cc_1542 N_VGND_c_2841_n N_A_1453_77#_c_3076_n 0.0130784f $X=7.78 $Y=0 $X2=0
+ $Y2=0
cc_1543 N_VGND_c_2845_n N_A_1453_77#_c_3076_n 0.0117103f $X=18 $Y=0 $X2=0 $Y2=0
cc_1544 N_VGND_c_2832_n N_A_1453_77#_c_3077_n 0.01855f $X=8.825 $Y=0 $X2=0 $Y2=0
cc_1545 N_VGND_c_2833_n N_A_1453_77#_c_3077_n 0.0157813f $X=8.91 $Y=0.445 $X2=0
+ $Y2=0
cc_1546 N_VGND_c_2845_n N_A_1453_77#_c_3077_n 0.0123988f $X=18 $Y=0 $X2=0 $Y2=0
cc_1547 N_VGND_c_2848_n N_A_1453_77#_c_3077_n 0.00739317f $X=7.92 $Y=0 $X2=0
+ $Y2=0
cc_1548 N_VGND_c_2845_n A_1840_47# 0.00830268f $X=18 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1549 N_noxref_30_c_2992_n N_noxref_32_c_3021_n 0.012638f $X=2.75 $Y=0.34
+ $X2=0 $Y2=0
cc_1550 N_noxref_30_c_2992_n N_noxref_32_c_3022_n 0.00546119f $X=2.75 $Y=0.34
+ $X2=0 $Y2=0
cc_1551 N_noxref_30_c_2994_n N_noxref_32_c_3022_n 0.0238586f $X=2.915 $Y=0.34
+ $X2=0 $Y2=0
cc_1552 N_noxref_32_c_3024_n N_A_1009_107#_c_3056_n 0.00964716f $X=4.535
+ $Y=0.825 $X2=0 $Y2=0
