* File: sky130_fd_sc_lp__srsdfrtp_1.spice
* Created: Wed Sep  2 10:39:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__srsdfrtp_1.pex.spice"
.subckt sky130_fd_sc_lp__srsdfrtp_1  VNB VPB SCE D SCD RESET_B CLK SLEEP_B VPWR
+ KAPWR Q VGND
* 
* VGND	VGND
* Q	Q
* KAPWR	KAPWR
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_SCE_M1003_g N_A_27_110#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.1155 PD=1.38 PS=1.39 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1040 N_A_332_136#_M1040_d N_SCE_M1040_g N_noxref_29_M1040_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1253 AS=0.1722 PD=1.065 PS=1.66 NRD=34.284 NRS=38.568 M=1 R=2.8
+ SA=75000.3 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1021 noxref_30 N_D_M1021_g N_A_332_136#_M1040_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1253 PD=0.63 PS=1.065 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75001
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1010 N_noxref_31_M1010_d N_A_27_110#_M1010_g noxref_30 VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_noxref_29_M1019_d N_SCD_M1019_g N_noxref_31_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.0588 PD=1.39 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_noxref_31_M1023_d N_RESET_B_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.1155 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 N_A_999_424#_M1033_d N_A_969_318#_M1033_g N_A_929_152#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.2093 PD=0.77 PS=1.88 NRD=19.992 NRS=52.848 M=1
+ R=2.8 SA=75000.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1032 N_A_332_136#_M1032_d N_A_1098_271#_M1032_g N_A_999_424#_M1033_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.1134 AS=0.0735 PD=1.38 PS=0.77 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1050 A_1343_119# N_A_1176_349#_M1050_g N_A_929_152#_M1050_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1042 N_VGND_M1042_d N_RESET_B_M1042_g A_1343_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0441 PD=1.39 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1046 N_VGND_M1046_d N_A_999_424#_M1046_g N_A_1176_349#_M1046_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.134158 AS=0.176 PD=1.23774 PS=1.83 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1029 N_A_969_318#_M1029_d N_A_1098_271#_M1029_g N_VGND_M1046_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.2703 AS=0.0880415 PD=2.42 PS=0.812264 NRD=168.156
+ NRS=31.428 M=1 R=2.8 SA=75000.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1035 A_1931_125# N_A_969_318#_M1035_g N_A_1176_349#_M1035_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0672 AS=0.176 PD=0.85 PS=1.83 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1026 N_A_1982_397#_M1026_d N_A_969_318#_M1026_g A_1931_125# VNB NSHORT L=0.15
+ W=0.64 AD=0.180528 AS=0.0672 PD=1.38264 PS=0.85 NRD=22.488 NRS=9.372 M=1
+ R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1018 A_2134_125# N_A_1098_271#_M1018_g N_A_1982_397#_M1026_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.118472 PD=0.63 PS=0.907358 NRD=14.28 NRS=30.708 M=1
+ R=2.8 SA=75001.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1011 A_2206_125# N_A_2176_99#_M1011_g A_2134_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_2176_99#_M1002_g A_2206_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0441 PD=1.39 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_2472_119# N_A_1982_397#_M1006_g N_A_2176_99#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1044 N_A_2544_119#_M1044_d N_A_1982_397#_M1044_g A_2472_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1047 N_VGND_M1047_d N_A_2586_249#_M1047_g N_A_2544_119#_M1044_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_2544_119#_M1007_d N_RESET_B_M1007_g N_VGND_M1047_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0672 PD=1.41 PS=0.74 NRD=0 NRS=11.424 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1048 A_3335_97# N_CLK_M1048_g N_A_1098_271#_M1048_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.168 PD=0.63 PS=1.64 NRD=14.28 NRS=32.856 M=1 R=2.8 SA=75000.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1028 A_3407_97# N_SLEEP_B_M1028_g A_3335_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_SLEEP_B_M1030_g A_3407_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.21765 AS=0.0441 PD=2.03 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1012 A_3694_73# N_SLEEP_B_M1012_g N_A_2586_249#_M1012_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SLEEP_B_M1014_g A_3694_73# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1031 N_A_3751_367#_M1031_d N_A_1982_397#_M1031_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=1.39 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1049 N_Q_M1049_d N_A_3751_367#_M1049_g N_VGND_M1049_s VNB NSHORT L=0.15 W=0.84
+ AD=0.231 AS=0.231 PD=2.23 PS=2.23 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1034 N_VPWR_M1034_d N_SCE_M1034_g N_A_27_110#_M1034_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.248 AS=0.1824 PD=1.415 PS=1.85 NRD=1.5366 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.8 A=0.096 P=1.58 MULT=1
MM1017 A_313_466# N_SCE_M1017_g N_VPWR_M1034_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.248 PD=0.88 PS=1.415 NRD=19.9955 NRS=150.823 M=1 R=4.26667
+ SA=75001.1 SB=75003.9 A=0.096 P=1.58 MULT=1
MM1039 N_A_332_136#_M1039_d N_D_M1039_g A_313_466# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2096 AS=0.0768 PD=1.295 PS=0.88 NRD=115.422 NRS=19.9955 M=1 R=4.26667
+ SA=75001.5 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1008 A_552_466# N_A_27_110#_M1008_g N_A_332_136#_M1039_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.2096 PD=1 PS=1.295 NRD=38.4741 NRS=0 M=1 R=4.26667
+ SA=75002.3 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_SCD_M1009_g A_552_466# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.3296 AS=0.1152 PD=1.67 PS=1 NRD=0 NRS=38.4741 M=1 R=4.26667 SA=75002.8
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1045 N_A_332_136#_M1045_d N_RESET_B_M1045_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.155774 AS=0.3296 PD=1.5034 PS=1.67 NRD=0 NRS=230.845 M=1 R=4.26667
+ SA=75004 SB=75001 A=0.096 P=1.58 MULT=1
MM1000 N_A_999_424#_M1000_d N_A_969_318#_M1000_g N_A_332_136#_M1045_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.10395 AS=0.102226 PD=0.915 PS=0.986604 NRD=100.844
+ NRS=56.2829 M=1 R=2.8 SA=75002.4 SB=75002 A=0.063 P=1.14 MULT=1
MM1004 A_1128_424# N_A_1098_271#_M1004_g N_A_999_424#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.10395 PD=0.66 PS=0.915 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75003 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_1176_349#_M1020_g A_1128_424# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1738 AS=0.0504 PD=1.39 PS=0.66 NRD=168.297 NRS=30.4759 M=1 R=2.8
+ SA=75003.4 SB=75001 A=0.063 P=1.14 MULT=1
MM1043 N_A_999_424#_M1043_d N_RESET_B_M1043_g N_VPWR_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.2173 AS=0.1738 PD=1.98 PS=1.39 NRD=56.2829 NRS=168.297 M=1 R=2.8
+ SA=75004.1 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_999_424#_M1001_g N_A_1176_349#_M1001_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.248538 AS=0.2394 PD=1.73108 PS=2.25 NRD=56.4799 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1013 N_A_969_318#_M1013_d N_A_1098_271#_M1013_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.189362 PD=1.85 PS=1.31892 NRD=0 NRS=36.9375 M=1
+ R=4.26667 SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1037 A_2069_397# N_A_1098_271#_M1037_g N_A_1982_397#_M1037_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1038 N_A_1176_349#_M1038_d N_A_1098_271#_M1038_g A_2069_397# VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 A_2836_390# N_A_969_318#_M1005_g N_A_1982_397#_M1005_s VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1022 N_KAPWR_M1022_d N_A_2176_99#_M1022_g A_2836_390# VPB PHIGHVT L=0.25 W=1
+ AD=0.1975 AS=0.12 PD=1.395 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1036 A_3063_390# N_A_2586_249#_M1036_g N_KAPWR_M1022_d VPB PHIGHVT L=0.25 W=1
+ AD=0.105 AS=0.1975 PD=1.21 PS=1.395 NRD=9.8303 NRS=22.6353 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1041 N_A_2176_99#_M1041_d N_RESET_B_M1041_g A_3063_390# VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125002 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1015 N_KAPWR_M1015_d N_A_1982_397#_M1015_g N_A_2176_99#_M1041_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.216707 AS=0.14 PD=1.70122 PS=1.28 NRD=0 NRS=0 M=1 R=4
+ SA=125002 SB=125001 A=0.25 P=2.5 MULT=1
MM1024 N_A_1098_271#_M1024_d N_CLK_M1024_g N_KAPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0992 AS=0.138693 PD=0.95 PS=1.08878 NRD=9.2196 NRS=49.7622 M=1
+ R=4.26667 SA=75003 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1027 N_KAPWR_M1027_d N_SLEEP_B_M1027_g N_A_1098_271#_M1024_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.189795 AS=0.0992 PD=1.22146 PS=0.95 NRD=74.3478 NRS=0 M=1
+ R=4.26667 SA=75003.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1025 N_A_2586_249#_M1025_d N_SLEEP_B_M1025_g N_KAPWR_M1027_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.4232 AS=0.296555 PD=2.96 PS=1.90854 NRD=23.64 NRS=22.6353 M=1
+ R=4 SA=125003 SB=125000 A=0.25 P=2.5 MULT=1
MM1051 N_VPWR_M1051_d N_A_1982_397#_M1051_g N_A_3751_367#_M1051_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.220733 AS=0.1824 PD=1.30695 PS=1.85 NRD=102.341 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1016 N_Q_M1016_d N_A_3751_367#_M1016_g N_VPWR_M1051_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.434567 PD=3.09 PS=2.57305 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75000.7 SB=75000.2 A=0.189 P=2.82 MULT=1
DX52_noxref VNB VPB NWDIODE A=38.7832 P=46.43
c_206 VNB 0 1.20173e-19 $X=0 $Y=0
c_358 VPB 0 1.73039e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__srsdfrtp_1.pxi.spice"
*
.ends
*
*
