* File: sky130_fd_sc_lp__o211a_m.pex.spice
* Created: Wed Sep  2 10:14:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211A_M%A_80_60# 1 2 3 12 16 20 21 23 24 27 29 32 33
+ 39 43 45
c76 12 0 1.47362e-19 $X=0.475 $Y=0.64
r77 40 43 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.54 $Y=0.495 $X2=2.94
+ $Y2=0.495
r78 35 37 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=3.025 $Y=1.865
+ $X2=3.025 $Y2=2
r79 34 45 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=2.625 $Y=1.78
+ $X2=2.54 $Y2=1.77
r80 33 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.93 $Y=1.78
+ $X2=3.025 $Y2=1.865
r81 33 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.93 $Y=1.78
+ $X2=2.625 $Y2=1.78
r82 32 45 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=1.675
+ $X2=2.54 $Y2=1.77
r83 31 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0.66
+ $X2=2.54 $Y2=0.495
r84 31 32 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=2.54 $Y=0.66
+ $X2=2.54 $Y2=1.675
r85 30 39 5.86152 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.105 $Y=1.77 $X2=2
+ $Y2=1.77
r86 29 45 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=1.77
+ $X2=2.54 $Y2=1.77
r87 29 30 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=2.455 $Y=1.77
+ $X2=2.105 $Y2=1.77
r88 25 39 0.793806 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=2 $Y=1.865 $X2=2
+ $Y2=1.77
r89 25 27 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2 $Y=1.865 $X2=2
+ $Y2=2
r90 23 39 5.86152 $w=1.8e-07 $l=1.09886e-07 $layer=LI1_cond $X=1.895 $Y=1.76
+ $X2=2 $Y2=1.77
r91 23 24 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=1.895 $Y=1.76
+ $X2=0.795 $Y2=1.76
r92 21 48 87.4515 $w=4.75e-07 $l=5.05e-07 $layer=POLY_cond $X=0.637 $Y=1.19
+ $X2=0.637 $Y2=1.695
r93 21 47 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.637 $Y=1.19
+ $X2=0.637 $Y2=1.025
r94 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=1.19 $X2=0.71 $Y2=1.19
r95 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=1.675
+ $X2=0.795 $Y2=1.76
r96 18 20 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.71 $Y=1.675
+ $X2=0.71 $Y2=1.19
r97 16 48 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.8 $Y=2.065 $X2=0.8
+ $Y2=1.695
r98 12 47 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=0.64
+ $X2=0.475 $Y2=1.025
r99 3 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.855 $X2=3.015 $Y2=2
r100 2 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.855 $X2=2 $Y2=2
r101 1 43 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.245 $X2=2.94 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%A1 3 7 11 14 15 18 19
c40 19 0 1.47362e-19 $X=1.25 $Y=1.07
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.25
+ $Y=1.07 $X2=1.25 $Y2=1.07
r42 15 19 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.25 $Y=1.295
+ $X2=1.25 $Y2=1.07
r43 13 18 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.25 $Y=1.425
+ $X2=1.25 $Y2=1.07
r44 13 14 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.292 $Y=1.425
+ $X2=1.292 $Y2=1.575
r45 11 18 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.25 $Y=1.055
+ $X2=1.25 $Y2=1.07
r46 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.292 $Y=0.905
+ $X2=1.292 $Y2=1.055
r47 7 14 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.425 $Y=2.065
+ $X2=1.425 $Y2=1.575
r48 3 10 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.425 $Y=0.455
+ $X2=1.425 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%A2 3 7 11 12 13 16 17
r36 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.875
+ $Y=1.07 $X2=1.875 $Y2=1.07
r37 13 17 4.57324 $w=5.08e-07 $l=1.95e-07 $layer=LI1_cond $X=1.68 $Y=1.24
+ $X2=1.875 $Y2=1.24
r38 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.875 $Y=1.41
+ $X2=1.875 $Y2=1.07
r39 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.41
+ $X2=1.875 $Y2=1.575
r40 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=0.905
+ $X2=1.875 $Y2=1.07
r41 7 10 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.935 $Y=0.455
+ $X2=1.935 $Y2=0.905
r42 3 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.785 $Y=2.065
+ $X2=1.785 $Y2=1.575
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%B1 4 7 12 13 14 18 19
r35 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.235
+ $Y=2.6 $X2=2.235 $Y2=2.6
r36 14 19 1.75894 $w=5.08e-07 $l=7.5e-08 $layer=LI1_cond $X=2.16 $Y=2.77
+ $X2=2.235 $Y2=2.77
r37 13 14 11.2572 $w=5.08e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.77
+ $X2=2.16 $Y2=2.77
r38 11 12 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=2.345 $Y=1.595
+ $X2=2.345 $Y2=1.745
r39 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=2.435
+ $X2=2.235 $Y2=2.6
r40 7 11 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.365 $Y=0.455
+ $X2=2.365 $Y2=1.595
r41 4 10 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.325 $Y=2.065
+ $X2=2.325 $Y2=2.435
r42 4 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.325 $Y=2.065
+ $X2=2.325 $Y2=1.745
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%C1 3 6 9 11 12 13 17
r25 17 19 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.852 $Y=1.005
+ $X2=2.852 $Y2=0.84
r26 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.89
+ $Y=1.005 $X2=2.89 $Y2=1.005
r27 13 18 8.35521 $w=3.98e-07 $l=2.9e-07 $layer=LI1_cond $X=3.005 $Y=1.295
+ $X2=3.005 $Y2=1.005
r28 12 18 2.30489 $w=3.98e-07 $l=8e-08 $layer=LI1_cond $X=3.005 $Y=0.925
+ $X2=3.005 $Y2=1.005
r29 9 11 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.8 $Y=2.065 $X2=2.8
+ $Y2=1.51
r30 6 11 42.3036 $w=4.05e-07 $l=2.02e-07 $layer=POLY_cond $X=2.852 $Y=1.308
+ $X2=2.852 $Y2=1.51
r31 5 17 5.08091 $w=4.05e-07 $l=3.7e-08 $layer=POLY_cond $X=2.852 $Y=1.042
+ $X2=2.852 $Y2=1.005
r32 5 6 36.5276 $w=4.05e-07 $l=2.66e-07 $layer=POLY_cond $X=2.852 $Y=1.042
+ $X2=2.852 $Y2=1.308
r33 3 19 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.725 $Y=0.455
+ $X2=2.725 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%X 1 2 7 8 9 10 11 12 13 35
r18 35 36 3.12317 $w=6.53e-07 $l=1e-08 $layer=LI1_cond $X=0.422 $Y=2.035
+ $X2=0.422 $Y2=2.025
r19 12 13 6.75647 $w=6.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.422 $Y=2.405
+ $X2=0.422 $Y2=2.775
r20 12 39 5.0217 $w=6.53e-07 $l=2.75e-07 $layer=LI1_cond $X=0.422 $Y=2.405
+ $X2=0.422 $Y2=2.13
r21 11 39 1.05912 $w=6.53e-07 $l=5.8e-08 $layer=LI1_cond $X=0.422 $Y=2.072
+ $X2=0.422 $Y2=2.13
r22 11 35 0.675647 $w=6.53e-07 $l=3.7e-08 $layer=LI1_cond $X=0.422 $Y=2.072
+ $X2=0.422 $Y2=2.035
r23 11 36 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=0.26 $Y=1.987
+ $X2=0.26 $Y2=2.025
r24 10 11 11.245 $w=3.28e-07 $l=3.22e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.987
r25 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r26 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.925 $X2=0.26
+ $Y2=1.295
r27 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.555 $X2=0.26
+ $Y2=0.925
r28 2 39 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.46
+ $Y=1.855 $X2=0.585 $Y2=2.13
r29 1 7 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.43 $X2=0.26 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%VPWR 1 2 9 11 14 18 20 22 29 30 33 36
r29 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r33 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.665 $Y2=3.33
r34 27 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.75 $Y=3.33 $X2=3.12
+ $Y2=3.33
r35 25 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r36 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 22 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.11 $Y2=3.33
r38 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 20 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 16 18 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.585 $Y=2.15
+ $X2=2.665 $Y2=2.15
r42 14 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=3.245
+ $X2=2.665 $Y2=3.33
r43 13 18 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.665 $Y=2.255
+ $X2=2.665 $Y2=2.15
r44 13 14 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.665 $Y=2.255
+ $X2=2.665 $Y2=3.245
r45 12 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=3.33
+ $X2=1.11 $Y2=3.33
r46 11 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=3.33
+ $X2=2.665 $Y2=3.33
r47 11 12 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=2.58 $Y=3.33
+ $X2=1.275 $Y2=3.33
r48 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=3.245 $X2=1.11
+ $Y2=3.33
r49 7 9 38.9386 $w=3.28e-07 $l=1.115e-06 $layer=LI1_cond $X=1.11 $Y=3.245
+ $X2=1.11 $Y2=2.13
r50 2 16 600 $w=1.7e-07 $l=3.76298e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.855 $X2=2.585 $Y2=2.15
r51 1 9 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=0.875
+ $Y=1.855 $X2=1.11 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%VGND 1 2 9 13 16 17 18 24 33 34 37
r44 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r46 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r47 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.64
+ $Y2=0
r49 28 30 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=2.16
+ $Y2=0
r50 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.64
+ $Y2=0
r52 24 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r53 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r54 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r56 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r57 18 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 16 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r59 16 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.7
+ $Y2=0
r60 15 26 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r61 15 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.7
+ $Y2=0
r62 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0
r63 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0.37
r64 7 17 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r65 7 9 28.6029 $w=1.88e-07 $l=4.9e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.575
r66 2 13 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.245 $X2=1.64 $Y2=0.37
r67 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.43 $X2=0.69 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_M%A_217_49# 1 2 9 11 12 15
r27 13 15 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.15 $Y=0.635
+ $X2=2.15 $Y2=0.52
r28 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.045 $Y=0.72
+ $X2=2.15 $Y2=0.635
r29 11 12 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.045 $Y=0.72
+ $X2=1.295 $Y2=0.72
r30 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.2 $Y=0.635
+ $X2=1.295 $Y2=0.72
r31 7 9 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=0.635 $X2=1.2
+ $Y2=0.52
r32 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.245 $X2=2.15 $Y2=0.52
r33 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.245 $X2=1.21 $Y2=0.52
.ends

