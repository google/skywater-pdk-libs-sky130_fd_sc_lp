* File: sky130_fd_sc_lp__buflp_4.spice
* Created: Wed Sep  2 09:36:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buflp_4.pex.spice"
.subckt sky130_fd_sc_lp__buflp_4  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_84_21#_M1003_g N_A_114_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.5 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_84_21#_M1004_g N_A_114_47#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1004_d N_A_84_21#_M1014_g N_A_114_47#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1001 N_X_M1001_d N_A_84_21#_M1001_g N_A_114_47#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1002 N_X_M1001_d N_A_84_21#_M1002_g N_A_114_47#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1009 N_X_M1009_d N_A_84_21#_M1009_g N_A_114_47#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1015 N_X_M1009_d N_A_84_21#_M1015_g N_A_114_47#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_A_84_21#_M1016_g N_A_114_47#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.294 AS=0.1176 PD=1.54 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1005 A_886_47# N_A_M1005_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.294 PD=1.08 PS=1.54 NRD=9.276 NRS=49.992 M=1 R=5.6 SA=75004.1 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1006 N_A_84_21#_M1006_d N_A_M1006_g A_886_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1008 PD=2.25 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75004.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_84_21#_M1000_g N_A_114_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_84_21#_M1011_g N_A_114_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1011_d N_A_84_21#_M1012_g N_A_114_367#_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1007 N_X_M1007_d N_A_84_21#_M1007_g N_A_114_367#_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.1764 PD=1.61 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1010 N_X_M1007_d N_A_84_21#_M1010_g N_A_114_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75002 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1013 N_X_M1013_d N_A_84_21#_M1013_g N_A_114_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75002.5 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1017 N_X_M1013_d N_A_84_21#_M1017_g N_A_114_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75003 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A_84_21#_M1019_g N_A_114_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2646 AS=0.2205 PD=1.68 PS=1.61 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75003.5 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1018 A_886_367# N_A_M1018_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1512
+ AS=0.2646 PD=1.5 PS=1.68 NRD=10.1455 NRS=10.9335 M=1 R=8.4 SA=75004.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_A_84_21#_M1008_d N_A_M1008_g A_886_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1512 PD=3.09 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75004.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.5559 P=15.05
*
.include "sky130_fd_sc_lp__buflp_4.pxi.spice"
*
.ends
*
*
