* File: sky130_fd_sc_lp__dlxtn_1.pxi.spice
* Created: Wed Sep  2 09:48:24 2020
* 
x_PM_SKY130_FD_SC_LP__DLXTN_1%D N_D_M1009_g N_D_M1001_g D D D N_D_c_131_n
+ N_D_c_132_n PM_SKY130_FD_SC_LP__DLXTN_1%D
x_PM_SKY130_FD_SC_LP__DLXTN_1%GATE_N N_GATE_N_c_162_n N_GATE_N_M1004_g
+ N_GATE_N_M1005_g N_GATE_N_c_164_n N_GATE_N_c_165_n N_GATE_N_c_166_n GATE_N
+ GATE_N GATE_N N_GATE_N_c_168_n PM_SKY130_FD_SC_LP__DLXTN_1%GATE_N
x_PM_SKY130_FD_SC_LP__DLXTN_1%A_228_129# N_A_228_129#_M1004_d
+ N_A_228_129#_M1005_d N_A_228_129#_M1000_g N_A_228_129#_c_209_n
+ N_A_228_129#_c_210_n N_A_228_129#_M1011_g N_A_228_129#_M1016_g
+ N_A_228_129#_M1002_g N_A_228_129#_c_213_n N_A_228_129#_c_214_n
+ N_A_228_129#_c_222_n N_A_228_129#_c_223_n N_A_228_129#_c_224_n
+ N_A_228_129#_c_247_p N_A_228_129#_c_225_n N_A_228_129#_c_226_n
+ N_A_228_129#_c_215_n N_A_228_129#_c_228_n N_A_228_129#_c_241_n
+ N_A_228_129#_c_230_n N_A_228_129#_c_216_n N_A_228_129#_c_217_n
+ N_A_228_129#_c_218_n N_A_228_129#_c_219_n
+ PM_SKY130_FD_SC_LP__DLXTN_1%A_228_129#
x_PM_SKY130_FD_SC_LP__DLXTN_1%A_59_129# N_A_59_129#_M1009_s N_A_59_129#_M1001_s
+ N_A_59_129#_M1012_g N_A_59_129#_c_356_n N_A_59_129#_c_357_n
+ N_A_59_129#_M1003_g N_A_59_129#_c_363_n N_A_59_129#_c_359_n
+ N_A_59_129#_c_365_n N_A_59_129#_c_366_n N_A_59_129#_c_403_n
+ N_A_59_129#_c_360_n N_A_59_129#_c_361_n N_A_59_129#_c_368_n
+ PM_SKY130_FD_SC_LP__DLXTN_1%A_59_129#
x_PM_SKY130_FD_SC_LP__DLXTN_1%A_342_481# N_A_342_481#_M1011_s
+ N_A_342_481#_M1000_s N_A_342_481#_M1013_g N_A_342_481#_c_439_n
+ N_A_342_481#_c_440_n N_A_342_481#_M1008_g N_A_342_481#_c_451_n
+ N_A_342_481#_c_441_n N_A_342_481#_c_442_n N_A_342_481#_c_453_n
+ N_A_342_481#_c_454_n N_A_342_481#_c_455_n N_A_342_481#_c_459_n
+ N_A_342_481#_c_443_n N_A_342_481#_c_444_n N_A_342_481#_c_445_n
+ N_A_342_481#_c_456_n N_A_342_481#_c_446_n N_A_342_481#_c_447_n
+ PM_SKY130_FD_SC_LP__DLXTN_1%A_342_481#
x_PM_SKY130_FD_SC_LP__DLXTN_1%A_842_413# N_A_842_413#_M1017_d
+ N_A_842_413#_M1010_d N_A_842_413#_M1007_g N_A_842_413#_M1014_g
+ N_A_842_413#_M1006_g N_A_842_413#_M1015_g N_A_842_413#_c_562_n
+ N_A_842_413#_c_552_n N_A_842_413#_c_563_n N_A_842_413#_c_553_n
+ N_A_842_413#_c_564_n N_A_842_413#_c_554_n N_A_842_413#_c_555_n
+ N_A_842_413#_c_566_n N_A_842_413#_c_567_n N_A_842_413#_c_556_n
+ N_A_842_413#_c_568_n N_A_842_413#_c_557_n N_A_842_413#_c_558_n
+ PM_SKY130_FD_SC_LP__DLXTN_1%A_842_413#
x_PM_SKY130_FD_SC_LP__DLXTN_1%A_656_481# N_A_656_481#_M1016_d
+ N_A_656_481#_M1013_d N_A_656_481#_M1017_g N_A_656_481#_M1010_g
+ N_A_656_481#_c_653_n N_A_656_481#_c_664_n N_A_656_481#_c_654_n
+ N_A_656_481#_c_646_n N_A_656_481#_c_647_n N_A_656_481#_c_648_n
+ N_A_656_481#_c_649_n N_A_656_481#_c_650_n N_A_656_481#_c_651_n
+ PM_SKY130_FD_SC_LP__DLXTN_1%A_656_481#
x_PM_SKY130_FD_SC_LP__DLXTN_1%VPWR N_VPWR_M1001_d N_VPWR_M1000_d N_VPWR_M1007_d
+ N_VPWR_M1015_s N_VPWR_c_744_n N_VPWR_c_745_n N_VPWR_c_746_n VPWR
+ N_VPWR_c_747_n N_VPWR_c_748_n N_VPWR_c_749_n N_VPWR_c_750_n N_VPWR_c_743_n
+ N_VPWR_c_752_n N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_755_n
+ PM_SKY130_FD_SC_LP__DLXTN_1%VPWR
x_PM_SKY130_FD_SC_LP__DLXTN_1%Q N_Q_M1006_d N_Q_M1015_d Q Q Q Q Q Q Q
+ N_Q_c_824_n PM_SKY130_FD_SC_LP__DLXTN_1%Q
x_PM_SKY130_FD_SC_LP__DLXTN_1%VGND N_VGND_M1009_d N_VGND_M1011_d N_VGND_M1014_d
+ N_VGND_M1006_s N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n
+ N_VGND_c_839_n N_VGND_c_840_n VGND N_VGND_c_841_n N_VGND_c_842_n
+ N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n
+ PM_SKY130_FD_SC_LP__DLXTN_1%VGND
cc_1 VNB N_D_M1001_g 0.00867796f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.725
cc_2 VNB D 0.014503f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_3 VNB N_D_c_131_n 0.0323087f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.34
cc_4 VNB N_D_c_132_n 0.0217107f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.175
cc_5 VNB N_GATE_N_c_162_n 0.0175076f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.175
cc_6 VNB N_GATE_N_M1005_g 0.022388f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.725
cc_7 VNB N_GATE_N_c_164_n 0.0296013f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_GATE_N_c_165_n 0.0378746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_GATE_N_c_166_n 0.00411253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB GATE_N 0.0224024f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.34
cc_11 VNB N_GATE_N_c_168_n 0.0480663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_228_129#_M1000_g 0.00602625f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_13 VNB N_A_228_129#_c_209_n 0.0358487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_228_129#_c_210_n 0.0159451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_228_129#_M1011_g 0.0205495f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.34
cc_16 VNB N_A_228_129#_M1016_g 0.0231485f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.34
cc_17 VNB N_A_228_129#_c_213_n 0.0197203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_228_129#_c_214_n 0.00772859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_228_129#_c_215_n 0.0115536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_228_129#_c_216_n 0.0389609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_228_129#_c_217_n 0.029213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_228_129#_c_218_n 0.0144857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_228_129#_c_219_n 0.00348687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_59_129#_c_356_n 0.0272312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_59_129#_c_357_n 0.0135593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_59_129#_M1003_g 0.0354416f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.34
cc_27 VNB N_A_59_129#_c_359_n 0.0314467f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.34
cc_28 VNB N_A_59_129#_c_360_n 0.0354847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_59_129#_c_361_n 0.016679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_342_481#_c_439_n 0.0215515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_342_481#_c_440_n 0.0130747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_342_481#_c_441_n 0.0172819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_342_481#_c_442_n 0.0508653f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.34
cc_34 VNB N_A_342_481#_c_443_n 0.0199204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_342_481#_c_444_n 0.00529457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_342_481#_c_445_n 0.00355104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_342_481#_c_446_n 9.01994e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_342_481#_c_447_n 0.0170528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_842_413#_M1014_g 0.058651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_842_413#_M1015_g 0.00452122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_842_413#_c_552_n 0.00792576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_842_413#_c_553_n 0.00523393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_842_413#_c_554_n 0.0122175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_842_413#_c_555_n 0.040711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_842_413#_c_556_n 0.0035929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_842_413#_c_557_n 0.00902034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_842_413#_c_558_n 0.0227221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_656_481#_M1017_g 0.0243559f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_49 VNB N_A_656_481#_c_646_n 0.00417946f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.34
cc_50 VNB N_A_656_481#_c_647_n 6.26511e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_656_481#_c_648_n 0.00355265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_656_481#_c_649_n 0.00468552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_656_481#_c_650_n 0.0323792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_656_481#_c_651_n 0.00287281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VPWR_c_743_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Q_c_824_n 0.0632177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_835_n 0.022504f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.175
cc_58 VNB N_VGND_c_836_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.34
cc_59 VNB N_VGND_c_837_n 0.00792333f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.34
cc_60 VNB N_VGND_c_838_n 0.0136234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_839_n 0.0406327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_840_n 0.00480879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_841_n 0.0461429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_842_n 0.0202998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_843_n 0.0163452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_844_n 0.36761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_845_n 0.0277418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_846_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_847_n 0.00534695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VPB N_D_M1001_g 0.0560599f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.725
cc_71 VPB N_GATE_N_M1005_g 0.0638032f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.725
cc_72 VPB N_A_228_129#_M1000_g 0.0686151f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_73 VPB N_A_228_129#_M1002_g 0.0206294f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.34
cc_74 VPB N_A_228_129#_c_222_n 0.010433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_228_129#_c_223_n 0.0158432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_228_129#_c_224_n 0.002837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_228_129#_c_225_n 0.0107921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_228_129#_c_226_n 0.0013623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_228_129#_c_215_n 0.00395455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_228_129#_c_228_n 0.0331926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_59_129#_M1012_g 0.0387345f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_82 VPB N_A_59_129#_c_363_n 0.0189918f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.34
cc_83 VPB N_A_59_129#_c_359_n 9.68173e-19 $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.34
cc_84 VPB N_A_59_129#_c_365_n 0.0646414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_59_129#_c_366_n 0.0446785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_59_129#_c_360_n 0.00739944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_59_129#_c_368_n 0.0117247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_342_481#_M1013_g 0.0239155f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_89 VPB N_A_342_481#_c_439_n 0.013686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_342_481#_c_440_n 0.00156028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_342_481#_c_451_n 0.0142743f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.505
cc_92 VPB N_A_342_481#_c_442_n 0.00687896f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.34
cc_93 VPB N_A_342_481#_c_453_n 0.0050118f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.34
cc_94 VPB N_A_342_481#_c_454_n 0.0262364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_342_481#_c_455_n 0.00506389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_342_481#_c_456_n 0.025682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_842_413#_M1007_g 0.0247264f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_98 VPB N_A_842_413#_M1014_g 0.0145818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_842_413#_M1015_g 0.0268579f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_842_413#_c_562_n 0.00334129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_842_413#_c_563_n 0.0108134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_842_413#_c_564_n 0.00711083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_842_413#_c_554_n 0.00523936f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_842_413#_c_566_n 0.0504072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_842_413#_c_567_n 0.00163076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_842_413#_c_568_n 0.00158047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_842_413#_c_557_n 3.19586e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_656_481#_M1010_g 0.0234132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_656_481#_c_653_n 0.00866035f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.34
cc_110 VPB N_A_656_481#_c_654_n 0.00643104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_656_481#_c_646_n 0.00195715f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.34
cc_112 VPB N_A_656_481#_c_647_n 7.75896e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_656_481#_c_649_n 0.00190261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_656_481#_c_650_n 0.00862416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_656_481#_c_651_n 6.57797e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_744_n 0.0108791f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.175
cc_117 VPB N_VPWR_c_745_n 0.00666604f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.34
cc_118 VPB N_VPWR_c_746_n 0.0166386f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.34
cc_119 VPB N_VPWR_c_747_n 0.0357068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_748_n 0.0461836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_749_n 0.0188738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_750_n 0.0157301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_743_n 0.0894838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_752_n 0.0263585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_753_n 0.00497591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_754_n 0.0307582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_755_n 0.00484208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_Q_c_824_n 0.0582069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 N_D_c_132_n N_GATE_N_c_162_n 0.0111679f $X=0.585 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_130 N_D_M1001_g N_GATE_N_M1005_g 0.0471663f $X=0.635 $Y=2.725 $X2=0 $Y2=0
cc_131 D N_GATE_N_M1005_g 0.0106183f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 D N_GATE_N_c_164_n 0.0232363f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_133 D N_GATE_N_c_166_n 0.00976792f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_D_c_131_n N_GATE_N_c_166_n 0.0181306f $X=0.585 $Y=1.34 $X2=0 $Y2=0
cc_135 D N_A_228_129#_c_214_n 0.0473328f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 D N_A_228_129#_c_230_n 0.0276236f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 D N_A_228_129#_c_216_n 0.00520054f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_138 N_D_M1001_g N_A_59_129#_c_359_n 0.00546105f $X=0.635 $Y=2.725 $X2=0 $Y2=0
cc_139 D N_A_59_129#_c_359_n 0.0263181f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_140 N_D_c_131_n N_A_59_129#_c_359_n 0.00817336f $X=0.585 $Y=1.34 $X2=0 $Y2=0
cc_141 N_D_c_132_n N_A_59_129#_c_359_n 0.00500228f $X=0.585 $Y=1.175 $X2=0 $Y2=0
cc_142 N_D_M1001_g N_A_59_129#_c_365_n 0.0244678f $X=0.635 $Y=2.725 $X2=0 $Y2=0
cc_143 N_D_M1001_g N_A_59_129#_c_366_n 0.017695f $X=0.635 $Y=2.725 $X2=0 $Y2=0
cc_144 D N_A_59_129#_c_366_n 0.0952857f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_145 N_D_c_131_n N_A_59_129#_c_366_n 0.00112163f $X=0.585 $Y=1.34 $X2=0 $Y2=0
cc_146 D N_A_59_129#_c_361_n 0.00199643f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_D_c_131_n N_A_59_129#_c_361_n 0.00329974f $X=0.585 $Y=1.34 $X2=0 $Y2=0
cc_148 D N_A_59_129#_c_368_n 0.00421666f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_149 N_D_c_131_n N_A_59_129#_c_368_n 0.00357888f $X=0.585 $Y=1.34 $X2=0 $Y2=0
cc_150 N_D_M1001_g N_VPWR_c_744_n 0.0029463f $X=0.635 $Y=2.725 $X2=0 $Y2=0
cc_151 N_D_M1001_g N_VPWR_c_743_n 0.010931f $X=0.635 $Y=2.725 $X2=0 $Y2=0
cc_152 N_D_M1001_g N_VPWR_c_752_n 0.0053602f $X=0.635 $Y=2.725 $X2=0 $Y2=0
cc_153 D N_VGND_c_835_n 0.0166546f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_D_c_132_n N_VGND_c_835_n 0.00344399f $X=0.585 $Y=1.175 $X2=0 $Y2=0
cc_155 N_D_c_132_n N_VGND_c_844_n 0.0046394f $X=0.585 $Y=1.175 $X2=0 $Y2=0
cc_156 N_D_c_132_n N_VGND_c_845_n 0.00404937f $X=0.585 $Y=1.175 $X2=0 $Y2=0
cc_157 N_GATE_N_c_165_n N_A_228_129#_c_210_n 0.012419f $X=1.59 $Y=1.175 $X2=0
+ $Y2=0
cc_158 GATE_N N_A_228_129#_c_210_n 0.00932997f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_159 N_GATE_N_c_162_n N_A_228_129#_c_214_n 0.00261884f $X=1.065 $Y=1.175 $X2=0
+ $Y2=0
cc_160 N_GATE_N_c_164_n N_A_228_129#_c_214_n 0.00373649f $X=1.515 $Y=1.25 $X2=0
+ $Y2=0
cc_161 N_GATE_N_c_165_n N_A_228_129#_c_214_n 0.0120004f $X=1.59 $Y=1.175 $X2=0
+ $Y2=0
cc_162 GATE_N N_A_228_129#_c_214_n 0.0611915f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_163 N_GATE_N_c_168_n N_A_228_129#_c_214_n 0.00100346f $X=1.68 $Y=0.38 $X2=0
+ $Y2=0
cc_164 N_GATE_N_M1005_g N_A_228_129#_c_222_n 4.68635e-19 $X=1.065 $Y=2.725 $X2=0
+ $Y2=0
cc_165 N_GATE_N_M1005_g N_A_228_129#_c_224_n 7.27903e-19 $X=1.065 $Y=2.725 $X2=0
+ $Y2=0
cc_166 N_GATE_N_c_165_n N_A_228_129#_c_241_n 6.63187e-19 $X=1.59 $Y=1.175 $X2=0
+ $Y2=0
cc_167 GATE_N N_A_228_129#_c_241_n 0.0268997f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_168 N_GATE_N_c_164_n N_A_228_129#_c_230_n 6.9094e-19 $X=1.515 $Y=1.25 $X2=0
+ $Y2=0
cc_169 N_GATE_N_c_164_n N_A_228_129#_c_216_n 0.012419f $X=1.515 $Y=1.25 $X2=0
+ $Y2=0
cc_170 GATE_N N_A_228_129#_c_218_n 4.76459e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_171 N_GATE_N_M1005_g N_A_59_129#_c_366_n 0.0181614f $X=1.065 $Y=2.725 $X2=0
+ $Y2=0
cc_172 N_GATE_N_c_164_n N_A_59_129#_c_366_n 0.00241877f $X=1.515 $Y=1.25 $X2=0
+ $Y2=0
cc_173 N_GATE_N_M1005_g N_A_342_481#_c_453_n 0.00465082f $X=1.065 $Y=2.725 $X2=0
+ $Y2=0
cc_174 N_GATE_N_M1005_g N_A_342_481#_c_455_n 0.00451651f $X=1.065 $Y=2.725 $X2=0
+ $Y2=0
cc_175 GATE_N N_A_342_481#_c_459_n 0.0287231f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_176 N_GATE_N_c_168_n N_A_342_481#_c_459_n 7.24385e-19 $X=1.68 $Y=0.38 $X2=0
+ $Y2=0
cc_177 N_GATE_N_M1005_g N_VPWR_c_744_n 0.00275171f $X=1.065 $Y=2.725 $X2=0 $Y2=0
cc_178 N_GATE_N_M1005_g N_VPWR_c_747_n 0.0053602f $X=1.065 $Y=2.725 $X2=0 $Y2=0
cc_179 N_GATE_N_M1005_g N_VPWR_c_743_n 0.0111019f $X=1.065 $Y=2.725 $X2=0 $Y2=0
cc_180 N_GATE_N_c_162_n N_VGND_c_835_n 0.00103802f $X=1.065 $Y=1.175 $X2=0 $Y2=0
cc_181 GATE_N N_VGND_c_835_n 0.028969f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_182 N_GATE_N_c_168_n N_VGND_c_835_n 0.00246916f $X=1.68 $Y=0.38 $X2=0 $Y2=0
cc_183 N_GATE_N_c_162_n N_VGND_c_841_n 0.00346478f $X=1.065 $Y=1.175 $X2=0 $Y2=0
cc_184 GATE_N N_VGND_c_841_n 0.0623353f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_185 N_GATE_N_c_168_n N_VGND_c_841_n 0.00625935f $X=1.68 $Y=0.38 $X2=0 $Y2=0
cc_186 N_GATE_N_c_162_n N_VGND_c_844_n 0.00386616f $X=1.065 $Y=1.175 $X2=0 $Y2=0
cc_187 GATE_N N_VGND_c_844_n 0.042156f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_188 N_GATE_N_c_168_n N_VGND_c_844_n 0.00876757f $X=1.68 $Y=0.38 $X2=0 $Y2=0
cc_189 N_A_228_129#_M1000_g N_A_59_129#_M1012_g 0.0178075f $X=2.05 $Y=2.725
+ $X2=0 $Y2=0
cc_190 N_A_228_129#_c_247_p N_A_59_129#_M1012_g 0.00294614f $X=2.185 $Y=2.905
+ $X2=0 $Y2=0
cc_191 N_A_228_129#_c_225_n N_A_59_129#_M1012_g 0.0126033f $X=3.67 $Y=2.46 $X2=0
+ $Y2=0
cc_192 N_A_228_129#_c_215_n N_A_59_129#_c_356_n 0.00170756f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_193 N_A_228_129#_c_217_n N_A_59_129#_c_356_n 0.0368611f $X=3.655 $Y=1.08
+ $X2=0 $Y2=0
cc_194 N_A_228_129#_c_218_n N_A_59_129#_c_356_n 0.0141948f $X=3.49 $Y=1.12 $X2=0
+ $Y2=0
cc_195 N_A_228_129#_c_219_n N_A_59_129#_c_356_n 6.06746e-19 $X=3.795 $Y=1.12
+ $X2=0 $Y2=0
cc_196 N_A_228_129#_c_209_n N_A_59_129#_c_357_n 0.0180476f $X=2.7 $Y=0.86 $X2=0
+ $Y2=0
cc_197 N_A_228_129#_c_241_n N_A_59_129#_c_357_n 9.68786e-19 $X=2.11 $Y=0.907
+ $X2=0 $Y2=0
cc_198 N_A_228_129#_c_216_n N_A_59_129#_c_357_n 0.0103451f $X=2.11 $Y=1.08 $X2=0
+ $Y2=0
cc_199 N_A_228_129#_c_218_n N_A_59_129#_c_357_n 0.00956935f $X=3.49 $Y=1.12
+ $X2=0 $Y2=0
cc_200 N_A_228_129#_M1011_g N_A_59_129#_M1003_g 0.0233286f $X=2.775 $Y=0.445
+ $X2=0 $Y2=0
cc_201 N_A_228_129#_M1016_g N_A_59_129#_M1003_g 0.0368611f $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_202 N_A_228_129#_c_218_n N_A_59_129#_M1003_g 0.00903469f $X=3.49 $Y=1.12
+ $X2=0 $Y2=0
cc_203 N_A_228_129#_M1000_g N_A_59_129#_c_366_n 0.0143433f $X=2.05 $Y=2.725
+ $X2=0 $Y2=0
cc_204 N_A_228_129#_c_213_n N_A_59_129#_c_366_n 0.0052532f $X=2.11 $Y=1.585
+ $X2=0 $Y2=0
cc_205 N_A_228_129#_c_214_n N_A_59_129#_c_366_n 0.0050048f $X=1.945 $Y=0.907
+ $X2=0 $Y2=0
cc_206 N_A_228_129#_c_222_n N_A_59_129#_c_366_n 0.0114801f $X=1.28 $Y=2.55 $X2=0
+ $Y2=0
cc_207 N_A_228_129#_c_230_n N_A_59_129#_c_366_n 0.0258988f $X=2.11 $Y=1.08 $X2=0
+ $Y2=0
cc_208 N_A_228_129#_c_218_n N_A_59_129#_c_366_n 0.0101007f $X=3.49 $Y=1.12 $X2=0
+ $Y2=0
cc_209 N_A_228_129#_M1000_g N_A_59_129#_c_403_n 4.98752e-19 $X=2.05 $Y=2.725
+ $X2=0 $Y2=0
cc_210 N_A_228_129#_c_230_n N_A_59_129#_c_403_n 0.00841641f $X=2.11 $Y=1.08
+ $X2=0 $Y2=0
cc_211 N_A_228_129#_c_216_n N_A_59_129#_c_403_n 0.00120379f $X=2.11 $Y=1.08
+ $X2=0 $Y2=0
cc_212 N_A_228_129#_c_218_n N_A_59_129#_c_403_n 0.0244713f $X=3.49 $Y=1.12 $X2=0
+ $Y2=0
cc_213 N_A_228_129#_M1000_g N_A_59_129#_c_360_n 0.00992651f $X=2.05 $Y=2.725
+ $X2=0 $Y2=0
cc_214 N_A_228_129#_c_213_n N_A_59_129#_c_360_n 0.0103451f $X=2.11 $Y=1.585
+ $X2=0 $Y2=0
cc_215 N_A_228_129#_c_230_n N_A_59_129#_c_360_n 9.56785e-19 $X=2.11 $Y=1.08
+ $X2=0 $Y2=0
cc_216 N_A_228_129#_c_223_n N_A_342_481#_M1000_s 0.00344308f $X=2.1 $Y=2.99
+ $X2=0 $Y2=0
cc_217 N_A_228_129#_c_225_n N_A_342_481#_M1013_g 0.0115575f $X=3.67 $Y=2.46
+ $X2=0 $Y2=0
cc_218 N_A_228_129#_c_215_n N_A_342_481#_M1013_g 9.77864e-19 $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_219 N_A_228_129#_c_228_n N_A_342_481#_M1013_g 0.0195488f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_220 N_A_228_129#_c_225_n N_A_342_481#_c_439_n 0.00419203f $X=3.67 $Y=2.46
+ $X2=0 $Y2=0
cc_221 N_A_228_129#_c_215_n N_A_342_481#_c_439_n 0.0142964f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_222 N_A_228_129#_c_228_n N_A_342_481#_c_439_n 0.0218211f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_223 N_A_228_129#_c_217_n N_A_342_481#_c_439_n 0.0152752f $X=3.655 $Y=1.08
+ $X2=0 $Y2=0
cc_224 N_A_228_129#_c_219_n N_A_342_481#_c_439_n 0.00157973f $X=3.795 $Y=1.12
+ $X2=0 $Y2=0
cc_225 N_A_228_129#_c_218_n N_A_342_481#_c_440_n 0.00204968f $X=3.49 $Y=1.12
+ $X2=0 $Y2=0
cc_226 N_A_228_129#_c_225_n N_A_342_481#_c_451_n 0.00125351f $X=3.67 $Y=2.46
+ $X2=0 $Y2=0
cc_227 N_A_228_129#_M1016_g N_A_342_481#_c_441_n 0.0207144f $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_228 N_A_228_129#_c_215_n N_A_342_481#_c_442_n 0.00713357f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_229 N_A_228_129#_c_219_n N_A_342_481#_c_442_n 0.0016865f $X=3.795 $Y=1.12
+ $X2=0 $Y2=0
cc_230 N_A_228_129#_M1000_g N_A_342_481#_c_453_n 0.00744548f $X=2.05 $Y=2.725
+ $X2=0 $Y2=0
cc_231 N_A_228_129#_c_222_n N_A_342_481#_c_453_n 0.018945f $X=1.28 $Y=2.55 $X2=0
+ $Y2=0
cc_232 N_A_228_129#_c_223_n N_A_342_481#_c_453_n 0.0142651f $X=2.1 $Y=2.99 $X2=0
+ $Y2=0
cc_233 N_A_228_129#_c_226_n N_A_342_481#_c_453_n 0.00828416f $X=2.27 $Y=2.46
+ $X2=0 $Y2=0
cc_234 N_A_228_129#_M1000_g N_A_342_481#_c_454_n 0.0168783f $X=2.05 $Y=2.725
+ $X2=0 $Y2=0
cc_235 N_A_228_129#_c_225_n N_A_342_481#_c_454_n 0.0893352f $X=3.67 $Y=2.46
+ $X2=0 $Y2=0
cc_236 N_A_228_129#_c_226_n N_A_342_481#_c_454_n 0.0141853f $X=2.27 $Y=2.46
+ $X2=0 $Y2=0
cc_237 N_A_228_129#_c_215_n N_A_342_481#_c_454_n 0.0111883f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_238 N_A_228_129#_c_228_n N_A_342_481#_c_454_n 5.90248e-19 $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_239 N_A_228_129#_c_209_n N_A_342_481#_c_443_n 0.00361466f $X=2.7 $Y=0.86
+ $X2=0 $Y2=0
cc_240 N_A_228_129#_M1011_g N_A_342_481#_c_443_n 0.00901476f $X=2.775 $Y=0.445
+ $X2=0 $Y2=0
cc_241 N_A_228_129#_M1016_g N_A_342_481#_c_443_n 0.0119732f $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_242 N_A_228_129#_c_217_n N_A_342_481#_c_443_n 0.0044365f $X=3.655 $Y=1.08
+ $X2=0 $Y2=0
cc_243 N_A_228_129#_c_218_n N_A_342_481#_c_443_n 0.0930983f $X=3.49 $Y=1.12
+ $X2=0 $Y2=0
cc_244 N_A_228_129#_c_209_n N_A_342_481#_c_444_n 0.00781278f $X=2.7 $Y=0.86
+ $X2=0 $Y2=0
cc_245 N_A_228_129#_c_241_n N_A_342_481#_c_444_n 0.00114341f $X=2.11 $Y=0.907
+ $X2=0 $Y2=0
cc_246 N_A_228_129#_c_218_n N_A_342_481#_c_444_n 0.0148874f $X=3.49 $Y=1.12
+ $X2=0 $Y2=0
cc_247 N_A_228_129#_c_215_n N_A_342_481#_c_445_n 0.0318122f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_248 N_A_228_129#_c_228_n N_A_342_481#_c_445_n 4.86971e-19 $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_249 N_A_228_129#_c_218_n N_A_342_481#_c_445_n 0.0140115f $X=3.49 $Y=1.12
+ $X2=0 $Y2=0
cc_250 N_A_228_129#_c_215_n N_A_342_481#_c_456_n 0.00531734f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_251 N_A_228_129#_c_228_n N_A_342_481#_c_456_n 0.0191927f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_252 N_A_228_129#_M1016_g N_A_342_481#_c_446_n 4.64362e-19 $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_253 N_A_228_129#_c_215_n N_A_342_481#_c_446_n 0.014148f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_254 N_A_228_129#_c_217_n N_A_342_481#_c_446_n 7.33069e-19 $X=3.655 $Y=1.08
+ $X2=0 $Y2=0
cc_255 N_A_228_129#_c_219_n N_A_342_481#_c_446_n 0.0199763f $X=3.795 $Y=1.12
+ $X2=0 $Y2=0
cc_256 N_A_228_129#_c_217_n N_A_342_481#_c_447_n 0.0209488f $X=3.655 $Y=1.08
+ $X2=0 $Y2=0
cc_257 N_A_228_129#_M1002_g N_A_842_413#_M1007_g 0.0205128f $X=3.745 $Y=2.615
+ $X2=0 $Y2=0
cc_258 N_A_228_129#_c_225_n N_A_842_413#_M1007_g 5.55633e-19 $X=3.67 $Y=2.46
+ $X2=0 $Y2=0
cc_259 N_A_228_129#_c_215_n N_A_842_413#_M1007_g 4.10796e-19 $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_260 N_A_228_129#_c_215_n N_A_842_413#_M1014_g 3.81179e-19 $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_261 N_A_228_129#_c_228_n N_A_842_413#_c_566_n 0.0134162f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_262 N_A_228_129#_c_225_n N_A_656_481#_M1013_d 0.00311814f $X=3.67 $Y=2.46
+ $X2=0 $Y2=0
cc_263 N_A_228_129#_M1002_g N_A_656_481#_c_653_n 0.0151308f $X=3.745 $Y=2.615
+ $X2=0 $Y2=0
cc_264 N_A_228_129#_c_225_n N_A_656_481#_c_653_n 0.037408f $X=3.67 $Y=2.46 $X2=0
+ $Y2=0
cc_265 N_A_228_129#_c_228_n N_A_656_481#_c_653_n 0.00263246f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_266 N_A_228_129#_M1016_g N_A_656_481#_c_664_n 0.00292613f $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_267 N_A_228_129#_M1002_g N_A_656_481#_c_654_n 0.00421355f $X=3.745 $Y=2.615
+ $X2=0 $Y2=0
cc_268 N_A_228_129#_c_225_n N_A_656_481#_c_654_n 0.0140286f $X=3.67 $Y=2.46
+ $X2=0 $Y2=0
cc_269 N_A_228_129#_c_215_n N_A_656_481#_c_654_n 0.0447503f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_270 N_A_228_129#_c_228_n N_A_656_481#_c_654_n 0.00264918f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_271 N_A_228_129#_c_215_n N_A_656_481#_c_647_n 0.0141518f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_272 N_A_228_129#_c_215_n N_A_656_481#_c_651_n 0.00662931f $X=3.835 $Y=2.06
+ $X2=0 $Y2=0
cc_273 N_A_228_129#_c_223_n N_VPWR_M1000_d 0.00138006f $X=2.1 $Y=2.99 $X2=0
+ $Y2=0
cc_274 N_A_228_129#_c_247_p N_VPWR_M1000_d 0.00439327f $X=2.185 $Y=2.905 $X2=0
+ $Y2=0
cc_275 N_A_228_129#_c_225_n N_VPWR_M1000_d 0.00840917f $X=3.67 $Y=2.46 $X2=0
+ $Y2=0
cc_276 N_A_228_129#_c_222_n N_VPWR_c_744_n 0.00153963f $X=1.28 $Y=2.55 $X2=0
+ $Y2=0
cc_277 N_A_228_129#_c_224_n N_VPWR_c_744_n 0.00252055f $X=1.445 $Y=2.99 $X2=0
+ $Y2=0
cc_278 N_A_228_129#_M1000_g N_VPWR_c_745_n 0.00264791f $X=2.05 $Y=2.725 $X2=0
+ $Y2=0
cc_279 N_A_228_129#_c_223_n N_VPWR_c_745_n 0.0143348f $X=2.1 $Y=2.99 $X2=0 $Y2=0
cc_280 N_A_228_129#_c_247_p N_VPWR_c_745_n 0.0142172f $X=2.185 $Y=2.905 $X2=0
+ $Y2=0
cc_281 N_A_228_129#_c_225_n N_VPWR_c_745_n 0.0204744f $X=3.67 $Y=2.46 $X2=0
+ $Y2=0
cc_282 N_A_228_129#_M1000_g N_VPWR_c_747_n 0.00325872f $X=2.05 $Y=2.725 $X2=0
+ $Y2=0
cc_283 N_A_228_129#_c_223_n N_VPWR_c_747_n 0.0539002f $X=2.1 $Y=2.99 $X2=0 $Y2=0
cc_284 N_A_228_129#_c_224_n N_VPWR_c_747_n 0.0211709f $X=1.445 $Y=2.99 $X2=0
+ $Y2=0
cc_285 N_A_228_129#_M1002_g N_VPWR_c_748_n 7.10185e-19 $X=3.745 $Y=2.615 $X2=0
+ $Y2=0
cc_286 N_A_228_129#_M1000_g N_VPWR_c_743_n 0.00623479f $X=2.05 $Y=2.725 $X2=0
+ $Y2=0
cc_287 N_A_228_129#_c_223_n N_VPWR_c_743_n 0.0305501f $X=2.1 $Y=2.99 $X2=0 $Y2=0
cc_288 N_A_228_129#_c_224_n N_VPWR_c_743_n 0.0114733f $X=1.445 $Y=2.99 $X2=0
+ $Y2=0
cc_289 N_A_228_129#_c_225_n N_VPWR_c_743_n 0.0258868f $X=3.67 $Y=2.46 $X2=0
+ $Y2=0
cc_290 N_A_228_129#_c_225_n A_584_481# 0.00183853f $X=3.67 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_228_129#_c_225_n A_764_481# 0.00174488f $X=3.67 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_228_129#_M1011_g N_VGND_c_836_n 0.00951069f $X=2.775 $Y=0.445 $X2=0
+ $Y2=0
cc_293 N_A_228_129#_M1016_g N_VGND_c_836_n 0.00198488f $X=3.565 $Y=0.445 $X2=0
+ $Y2=0
cc_294 N_A_228_129#_M1016_g N_VGND_c_839_n 0.00428022f $X=3.565 $Y=0.445 $X2=0
+ $Y2=0
cc_295 N_A_228_129#_M1011_g N_VGND_c_841_n 0.00355956f $X=2.775 $Y=0.445 $X2=0
+ $Y2=0
cc_296 N_A_228_129#_c_209_n N_VGND_c_844_n 0.00361074f $X=2.7 $Y=0.86 $X2=0
+ $Y2=0
cc_297 N_A_228_129#_M1011_g N_VGND_c_844_n 0.00563228f $X=2.775 $Y=0.445 $X2=0
+ $Y2=0
cc_298 N_A_228_129#_M1016_g N_VGND_c_844_n 0.00619329f $X=3.565 $Y=0.445 $X2=0
+ $Y2=0
cc_299 N_A_59_129#_c_356_n N_A_342_481#_c_440_n 0.00854253f $X=3.13 $Y=1.22
+ $X2=0 $Y2=0
cc_300 N_A_59_129#_c_366_n N_A_342_481#_c_440_n 6.3326e-19 $X=2.56 $Y=1.77 $X2=0
+ $Y2=0
cc_301 N_A_59_129#_c_403_n N_A_342_481#_c_440_n 5.38893e-19 $X=2.725 $Y=1.43
+ $X2=0 $Y2=0
cc_302 N_A_59_129#_c_360_n N_A_342_481#_c_440_n 0.034646f $X=2.725 $Y=1.43 $X2=0
+ $Y2=0
cc_303 N_A_59_129#_M1012_g N_A_342_481#_c_451_n 0.034646f $X=2.845 $Y=2.725
+ $X2=0 $Y2=0
cc_304 N_A_59_129#_M1012_g N_A_342_481#_c_454_n 0.0122495f $X=2.845 $Y=2.725
+ $X2=0 $Y2=0
cc_305 N_A_59_129#_c_363_n N_A_342_481#_c_454_n 0.00600429f $X=2.74 $Y=1.935
+ $X2=0 $Y2=0
cc_306 N_A_59_129#_c_366_n N_A_342_481#_c_454_n 0.0720391f $X=2.56 $Y=1.77 $X2=0
+ $Y2=0
cc_307 N_A_59_129#_c_366_n N_A_342_481#_c_455_n 0.0170614f $X=2.56 $Y=1.77 $X2=0
+ $Y2=0
cc_308 N_A_59_129#_c_357_n N_A_342_481#_c_443_n 0.00153254f $X=2.92 $Y=1.22
+ $X2=0 $Y2=0
cc_309 N_A_59_129#_M1003_g N_A_342_481#_c_443_n 0.0111448f $X=3.205 $Y=0.445
+ $X2=0 $Y2=0
cc_310 N_A_59_129#_c_356_n N_A_342_481#_c_445_n 6.80268e-19 $X=3.13 $Y=1.22
+ $X2=0 $Y2=0
cc_311 N_A_59_129#_c_366_n N_A_342_481#_c_445_n 0.0114372f $X=2.56 $Y=1.77 $X2=0
+ $Y2=0
cc_312 N_A_59_129#_c_403_n N_A_342_481#_c_445_n 0.00794738f $X=2.725 $Y=1.43
+ $X2=0 $Y2=0
cc_313 N_A_59_129#_c_360_n N_A_342_481#_c_445_n 0.00235462f $X=2.725 $Y=1.43
+ $X2=0 $Y2=0
cc_314 N_A_59_129#_c_363_n N_A_342_481#_c_456_n 0.034646f $X=2.74 $Y=1.935 $X2=0
+ $Y2=0
cc_315 N_A_59_129#_M1012_g N_A_656_481#_c_653_n 9.91921e-19 $X=2.845 $Y=2.725
+ $X2=0 $Y2=0
cc_316 N_A_59_129#_c_365_n N_VPWR_c_744_n 0.00315252f $X=0.42 $Y=2.55 $X2=0
+ $Y2=0
cc_317 N_A_59_129#_c_366_n N_VPWR_c_744_n 0.0100966f $X=2.56 $Y=1.77 $X2=0 $Y2=0
cc_318 N_A_59_129#_M1012_g N_VPWR_c_745_n 0.00848238f $X=2.845 $Y=2.725 $X2=0
+ $Y2=0
cc_319 N_A_59_129#_M1012_g N_VPWR_c_748_n 0.0053602f $X=2.845 $Y=2.725 $X2=0
+ $Y2=0
cc_320 N_A_59_129#_M1012_g N_VPWR_c_743_n 0.00612193f $X=2.845 $Y=2.725 $X2=0
+ $Y2=0
cc_321 N_A_59_129#_c_365_n N_VPWR_c_743_n 0.0153999f $X=0.42 $Y=2.55 $X2=0 $Y2=0
cc_322 N_A_59_129#_c_365_n N_VPWR_c_752_n 0.0268349f $X=0.42 $Y=2.55 $X2=0 $Y2=0
cc_323 N_A_59_129#_M1003_g N_VGND_c_836_n 0.00951109f $X=3.205 $Y=0.445 $X2=0
+ $Y2=0
cc_324 N_A_59_129#_M1003_g N_VGND_c_839_n 0.00355956f $X=3.205 $Y=0.445 $X2=0
+ $Y2=0
cc_325 N_A_59_129#_M1003_g N_VGND_c_844_n 0.00406467f $X=3.205 $Y=0.445 $X2=0
+ $Y2=0
cc_326 N_A_59_129#_c_361_n N_VGND_c_844_n 0.0113896f $X=0.42 $Y=0.84 $X2=0 $Y2=0
cc_327 N_A_59_129#_c_361_n N_VGND_c_845_n 0.00645798f $X=0.42 $Y=0.84 $X2=0
+ $Y2=0
cc_328 N_A_342_481#_c_441_n N_A_842_413#_M1014_g 0.0194147f $X=4.195 $Y=0.765
+ $X2=0 $Y2=0
cc_329 N_A_342_481#_c_442_n N_A_842_413#_M1014_g 0.00699351f $X=4.195 $Y=1.27
+ $X2=0 $Y2=0
cc_330 N_A_342_481#_c_443_n N_A_842_413#_M1014_g 4.21897e-19 $X=4.09 $Y=0.74
+ $X2=0 $Y2=0
cc_331 N_A_342_481#_c_446_n N_A_842_413#_M1014_g 5.59411e-19 $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_332 N_A_342_481#_c_447_n N_A_842_413#_M1014_g 0.0412721f $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_333 N_A_342_481#_c_442_n N_A_842_413#_c_566_n 0.00194462f $X=4.195 $Y=1.27
+ $X2=0 $Y2=0
cc_334 N_A_342_481#_M1013_g N_A_656_481#_c_653_n 0.0070696f $X=3.205 $Y=2.725
+ $X2=0 $Y2=0
cc_335 N_A_342_481#_c_441_n N_A_656_481#_c_664_n 0.00905063f $X=4.195 $Y=0.765
+ $X2=0 $Y2=0
cc_336 N_A_342_481#_c_443_n N_A_656_481#_c_664_n 0.0328879f $X=4.09 $Y=0.74
+ $X2=0 $Y2=0
cc_337 N_A_342_481#_c_447_n N_A_656_481#_c_664_n 0.0030012f $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_338 N_A_342_481#_c_442_n N_A_656_481#_c_646_n 0.0018996f $X=4.195 $Y=1.27
+ $X2=0 $Y2=0
cc_339 N_A_342_481#_c_446_n N_A_656_481#_c_646_n 6.52347e-19 $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_340 N_A_342_481#_c_442_n N_A_656_481#_c_647_n 0.00685352f $X=4.195 $Y=1.27
+ $X2=0 $Y2=0
cc_341 N_A_342_481#_c_446_n N_A_656_481#_c_647_n 0.0157287f $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_342 N_A_342_481#_c_441_n N_A_656_481#_c_648_n 0.00389315f $X=4.195 $Y=0.765
+ $X2=0 $Y2=0
cc_343 N_A_342_481#_c_443_n N_A_656_481#_c_648_n 0.0140835f $X=4.09 $Y=0.74
+ $X2=0 $Y2=0
cc_344 N_A_342_481#_c_446_n N_A_656_481#_c_648_n 0.0310144f $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_345 N_A_342_481#_c_447_n N_A_656_481#_c_648_n 0.00296965f $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_346 N_A_342_481#_c_442_n N_A_656_481#_c_651_n 0.00328452f $X=4.195 $Y=1.27
+ $X2=0 $Y2=0
cc_347 N_A_342_481#_c_446_n N_A_656_481#_c_651_n 0.0146418f $X=4.195 $Y=0.93
+ $X2=0 $Y2=0
cc_348 N_A_342_481#_M1013_g N_VPWR_c_748_n 0.00501304f $X=3.205 $Y=2.725 $X2=0
+ $Y2=0
cc_349 N_A_342_481#_M1013_g N_VPWR_c_743_n 0.00647292f $X=3.205 $Y=2.725 $X2=0
+ $Y2=0
cc_350 N_A_342_481#_c_443_n N_VGND_c_836_n 0.0201955f $X=4.09 $Y=0.74 $X2=0
+ $Y2=0
cc_351 N_A_342_481#_c_441_n N_VGND_c_839_n 0.00362032f $X=4.195 $Y=0.765 $X2=0
+ $Y2=0
cc_352 N_A_342_481#_c_443_n N_VGND_c_839_n 0.00943729f $X=4.09 $Y=0.74 $X2=0
+ $Y2=0
cc_353 N_A_342_481#_c_459_n N_VGND_c_841_n 0.0102922f $X=2.56 $Y=0.46 $X2=0
+ $Y2=0
cc_354 N_A_342_481#_c_443_n N_VGND_c_841_n 0.00289361f $X=4.09 $Y=0.74 $X2=0
+ $Y2=0
cc_355 N_A_342_481#_M1011_s N_VGND_c_844_n 0.00262842f $X=2.435 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_A_342_481#_c_441_n N_VGND_c_844_n 0.00591116f $X=4.195 $Y=0.765 $X2=0
+ $Y2=0
cc_357 N_A_342_481#_c_459_n N_VGND_c_844_n 0.00710598f $X=2.56 $Y=0.46 $X2=0
+ $Y2=0
cc_358 N_A_342_481#_c_443_n N_VGND_c_844_n 0.0213008f $X=4.09 $Y=0.74 $X2=0
+ $Y2=0
cc_359 N_A_342_481#_c_443_n A_836_47# 0.00123175f $X=4.09 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_360 N_A_842_413#_M1014_g N_A_656_481#_M1017_g 0.0215302f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_361 N_A_842_413#_c_553_n N_A_656_481#_M1017_g 0.00615097f $X=5.475 $Y=1.255
+ $X2=0 $Y2=0
cc_362 N_A_842_413#_M1014_g N_A_656_481#_M1010_g 0.00667285f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_363 N_A_842_413#_c_562_n N_A_656_481#_M1010_g 0.019101f $X=5.36 $Y=2.05 $X2=0
+ $Y2=0
cc_364 N_A_842_413#_c_563_n N_A_656_481#_M1010_g 0.00330549f $X=5.495 $Y=2.38
+ $X2=0 $Y2=0
cc_365 N_A_842_413#_c_564_n N_A_656_481#_M1010_g 0.00364773f $X=5.495 $Y=1.89
+ $X2=0 $Y2=0
cc_366 N_A_842_413#_c_566_n N_A_656_481#_M1010_g 0.00874013f $X=4.615 $Y=2.05
+ $X2=0 $Y2=0
cc_367 N_A_842_413#_c_567_n N_A_656_481#_M1010_g 3.3804e-19 $X=4.78 $Y=2.085
+ $X2=0 $Y2=0
cc_368 N_A_842_413#_M1007_g N_A_656_481#_c_653_n 0.00807099f $X=4.285 $Y=2.615
+ $X2=0 $Y2=0
cc_369 N_A_842_413#_M1014_g N_A_656_481#_c_664_n 0.0058488f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_370 N_A_842_413#_M1007_g N_A_656_481#_c_654_n 0.0157031f $X=4.285 $Y=2.615
+ $X2=0 $Y2=0
cc_371 N_A_842_413#_M1014_g N_A_656_481#_c_654_n 0.00302047f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_372 N_A_842_413#_c_566_n N_A_656_481#_c_654_n 0.00723224f $X=4.615 $Y=2.05
+ $X2=0 $Y2=0
cc_373 N_A_842_413#_c_567_n N_A_656_481#_c_654_n 0.0198326f $X=4.78 $Y=2.085
+ $X2=0 $Y2=0
cc_374 N_A_842_413#_c_566_n N_A_656_481#_c_646_n 0.00481766f $X=4.615 $Y=2.05
+ $X2=0 $Y2=0
cc_375 N_A_842_413#_c_567_n N_A_656_481#_c_646_n 7.00411e-19 $X=4.78 $Y=2.085
+ $X2=0 $Y2=0
cc_376 N_A_842_413#_M1014_g N_A_656_481#_c_648_n 0.0162531f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_377 N_A_842_413#_M1014_g N_A_656_481#_c_649_n 0.0169783f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_378 N_A_842_413#_c_562_n N_A_656_481#_c_649_n 0.0287973f $X=5.36 $Y=2.05
+ $X2=0 $Y2=0
cc_379 N_A_842_413#_c_564_n N_A_656_481#_c_649_n 0.0141133f $X=5.495 $Y=1.89
+ $X2=0 $Y2=0
cc_380 N_A_842_413#_c_566_n N_A_656_481#_c_649_n 0.00150655f $X=4.615 $Y=2.05
+ $X2=0 $Y2=0
cc_381 N_A_842_413#_c_567_n N_A_656_481#_c_649_n 0.0116987f $X=4.78 $Y=2.085
+ $X2=0 $Y2=0
cc_382 N_A_842_413#_c_557_n N_A_656_481#_c_649_n 0.0280792f $X=5.525 $Y=1.42
+ $X2=0 $Y2=0
cc_383 N_A_842_413#_M1014_g N_A_656_481#_c_650_n 0.0181029f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_384 N_A_842_413#_c_562_n N_A_656_481#_c_650_n 9.85223e-19 $X=5.36 $Y=2.05
+ $X2=0 $Y2=0
cc_385 N_A_842_413#_c_555_n N_A_656_481#_c_650_n 0.00471626f $X=6.09 $Y=1.42
+ $X2=0 $Y2=0
cc_386 N_A_842_413#_c_556_n N_A_656_481#_c_650_n 0.00303948f $X=5.42 $Y=1.075
+ $X2=0 $Y2=0
cc_387 N_A_842_413#_c_557_n N_A_656_481#_c_650_n 0.00467462f $X=5.525 $Y=1.42
+ $X2=0 $Y2=0
cc_388 N_A_842_413#_M1014_g N_A_656_481#_c_651_n 0.00954559f $X=4.645 $Y=0.445
+ $X2=0 $Y2=0
cc_389 N_A_842_413#_c_566_n N_A_656_481#_c_651_n 0.00278981f $X=4.615 $Y=2.05
+ $X2=0 $Y2=0
cc_390 N_A_842_413#_c_567_n N_A_656_481#_c_651_n 0.0138353f $X=4.78 $Y=2.085
+ $X2=0 $Y2=0
cc_391 N_A_842_413#_c_562_n N_VPWR_M1007_d 0.00481403f $X=5.36 $Y=2.05 $X2=0
+ $Y2=0
cc_392 N_A_842_413#_M1015_g N_VPWR_c_746_n 0.0217339f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_393 N_A_842_413#_c_563_n N_VPWR_c_746_n 0.0641828f $X=5.495 $Y=2.38 $X2=0
+ $Y2=0
cc_394 N_A_842_413#_c_564_n N_VPWR_c_746_n 0.0107025f $X=5.495 $Y=1.89 $X2=0
+ $Y2=0
cc_395 N_A_842_413#_c_554_n N_VPWR_c_746_n 0.0209545f $X=6.09 $Y=1.42 $X2=0
+ $Y2=0
cc_396 N_A_842_413#_c_555_n N_VPWR_c_746_n 0.00552801f $X=6.09 $Y=1.42 $X2=0
+ $Y2=0
cc_397 N_A_842_413#_c_568_n N_VPWR_c_746_n 0.0131191f $X=5.51 $Y=2.05 $X2=0
+ $Y2=0
cc_398 N_A_842_413#_M1007_g N_VPWR_c_748_n 0.00291497f $X=4.285 $Y=2.615 $X2=0
+ $Y2=0
cc_399 N_A_842_413#_c_563_n N_VPWR_c_749_n 0.0162117f $X=5.495 $Y=2.38 $X2=0
+ $Y2=0
cc_400 N_A_842_413#_M1015_g N_VPWR_c_750_n 0.00564095f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_842_413#_M1007_g N_VPWR_c_743_n 0.00268739f $X=4.285 $Y=2.615 $X2=0
+ $Y2=0
cc_402 N_A_842_413#_M1015_g N_VPWR_c_743_n 0.0104155f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_842_413#_c_563_n N_VPWR_c_743_n 0.0112946f $X=5.495 $Y=2.38 $X2=0
+ $Y2=0
cc_404 N_A_842_413#_M1007_g N_VPWR_c_754_n 0.00629044f $X=4.285 $Y=2.615 $X2=0
+ $Y2=0
cc_405 N_A_842_413#_c_562_n N_VPWR_c_754_n 0.0250929f $X=5.36 $Y=2.05 $X2=0
+ $Y2=0
cc_406 N_A_842_413#_c_563_n N_VPWR_c_754_n 0.00166817f $X=5.495 $Y=2.38 $X2=0
+ $Y2=0
cc_407 N_A_842_413#_c_566_n N_VPWR_c_754_n 0.00797612f $X=4.615 $Y=2.05 $X2=0
+ $Y2=0
cc_408 N_A_842_413#_c_567_n N_VPWR_c_754_n 0.0208952f $X=4.78 $Y=2.085 $X2=0
+ $Y2=0
cc_409 N_A_842_413#_c_554_n N_Q_c_824_n 0.0272547f $X=6.09 $Y=1.42 $X2=0 $Y2=0
cc_410 N_A_842_413#_c_558_n N_Q_c_824_n 0.0303311f $X=6.122 $Y=1.255 $X2=0 $Y2=0
cc_411 N_A_842_413#_M1014_g N_VGND_c_837_n 0.0104544f $X=4.645 $Y=0.445 $X2=0
+ $Y2=0
cc_412 N_A_842_413#_c_553_n N_VGND_c_837_n 4.88634e-19 $X=5.475 $Y=1.255 $X2=0
+ $Y2=0
cc_413 N_A_842_413#_c_552_n N_VGND_c_838_n 0.0452356f $X=5.385 $Y=0.42 $X2=0
+ $Y2=0
cc_414 N_A_842_413#_c_554_n N_VGND_c_838_n 0.0231351f $X=6.09 $Y=1.42 $X2=0
+ $Y2=0
cc_415 N_A_842_413#_c_555_n N_VGND_c_838_n 0.00553375f $X=6.09 $Y=1.42 $X2=0
+ $Y2=0
cc_416 N_A_842_413#_c_558_n N_VGND_c_838_n 0.0147033f $X=6.122 $Y=1.255 $X2=0
+ $Y2=0
cc_417 N_A_842_413#_M1014_g N_VGND_c_839_n 0.00495961f $X=4.645 $Y=0.445 $X2=0
+ $Y2=0
cc_418 N_A_842_413#_c_552_n N_VGND_c_842_n 0.0188828f $X=5.385 $Y=0.42 $X2=0
+ $Y2=0
cc_419 N_A_842_413#_c_558_n N_VGND_c_843_n 0.0049864f $X=6.122 $Y=1.255 $X2=0
+ $Y2=0
cc_420 N_A_842_413#_M1017_d N_VGND_c_844_n 0.00336915f $X=5.245 $Y=0.235 $X2=0
+ $Y2=0
cc_421 N_A_842_413#_M1014_g N_VGND_c_844_n 0.00925052f $X=4.645 $Y=0.445 $X2=0
+ $Y2=0
cc_422 N_A_842_413#_c_552_n N_VGND_c_844_n 0.010808f $X=5.385 $Y=0.42 $X2=0
+ $Y2=0
cc_423 N_A_842_413#_c_558_n N_VGND_c_844_n 0.00974208f $X=6.122 $Y=1.255 $X2=0
+ $Y2=0
cc_424 N_A_656_481#_c_649_n N_VPWR_M1007_d 0.00243167f $X=5.125 $Y=1.42 $X2=0
+ $Y2=0
cc_425 N_A_656_481#_c_653_n N_VPWR_c_745_n 0.0111063f $X=4.09 $Y=2.89 $X2=0
+ $Y2=0
cc_426 N_A_656_481#_M1010_g N_VPWR_c_746_n 0.00330902f $X=5.28 $Y=2.375 $X2=0
+ $Y2=0
cc_427 N_A_656_481#_c_653_n N_VPWR_c_748_n 0.0659705f $X=4.09 $Y=2.89 $X2=0
+ $Y2=0
cc_428 N_A_656_481#_M1010_g N_VPWR_c_749_n 0.00499542f $X=5.28 $Y=2.375 $X2=0
+ $Y2=0
cc_429 N_A_656_481#_M1010_g N_VPWR_c_743_n 0.010715f $X=5.28 $Y=2.375 $X2=0
+ $Y2=0
cc_430 N_A_656_481#_c_653_n N_VPWR_c_743_n 0.0389676f $X=4.09 $Y=2.89 $X2=0
+ $Y2=0
cc_431 N_A_656_481#_M1010_g N_VPWR_c_754_n 0.00427156f $X=5.28 $Y=2.375 $X2=0
+ $Y2=0
cc_432 N_A_656_481#_c_653_n N_VPWR_c_754_n 0.03151f $X=4.09 $Y=2.89 $X2=0 $Y2=0
cc_433 N_A_656_481#_c_654_n N_VPWR_c_754_n 0.0246056f $X=4.185 $Y=2.715 $X2=0
+ $Y2=0
cc_434 N_A_656_481#_c_653_n A_764_481# 0.00562367f $X=4.09 $Y=2.89 $X2=-0.19
+ $Y2=-0.245
cc_435 N_A_656_481#_c_654_n A_764_481# 0.0033642f $X=4.185 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_436 N_A_656_481#_c_664_n N_VGND_c_836_n 0.00599705f $X=4.46 $Y=0.37 $X2=0
+ $Y2=0
cc_437 N_A_656_481#_M1017_g N_VGND_c_837_n 0.0156537f $X=5.17 $Y=0.655 $X2=0
+ $Y2=0
cc_438 N_A_656_481#_c_664_n N_VGND_c_837_n 0.0155855f $X=4.46 $Y=0.37 $X2=0
+ $Y2=0
cc_439 N_A_656_481#_c_648_n N_VGND_c_837_n 0.0462495f $X=4.545 $Y=1.255 $X2=0
+ $Y2=0
cc_440 N_A_656_481#_c_649_n N_VGND_c_837_n 0.0274833f $X=5.125 $Y=1.42 $X2=0
+ $Y2=0
cc_441 N_A_656_481#_c_650_n N_VGND_c_837_n 0.00314491f $X=5.125 $Y=1.42 $X2=0
+ $Y2=0
cc_442 N_A_656_481#_M1017_g N_VGND_c_838_n 0.00344871f $X=5.17 $Y=0.655 $X2=0
+ $Y2=0
cc_443 N_A_656_481#_c_664_n N_VGND_c_839_n 0.047193f $X=4.46 $Y=0.37 $X2=0 $Y2=0
cc_444 N_A_656_481#_M1017_g N_VGND_c_842_n 0.00525069f $X=5.17 $Y=0.655 $X2=0
+ $Y2=0
cc_445 N_A_656_481#_M1016_d N_VGND_c_844_n 0.00347599f $X=3.64 $Y=0.235 $X2=0
+ $Y2=0
cc_446 N_A_656_481#_M1017_g N_VGND_c_844_n 0.0101648f $X=5.17 $Y=0.655 $X2=0
+ $Y2=0
cc_447 N_A_656_481#_c_664_n N_VGND_c_844_n 0.0328731f $X=4.46 $Y=0.37 $X2=0
+ $Y2=0
cc_448 N_A_656_481#_c_664_n A_836_47# 0.00826676f $X=4.46 $Y=0.37 $X2=-0.19
+ $Y2=-0.245
cc_449 N_A_656_481#_c_648_n A_836_47# 0.00238836f $X=4.545 $Y=1.255 $X2=-0.19
+ $Y2=-0.245
cc_450 N_VPWR_c_743_n N_Q_M1015_d 0.00302127f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_451 N_VPWR_c_746_n N_Q_c_824_n 0.0476029f $X=6.03 $Y=1.98 $X2=0 $Y2=0
cc_452 N_VPWR_c_750_n N_Q_c_824_n 0.0192376f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_453 N_VPWR_c_743_n N_Q_c_824_n 0.0111968f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_454 N_Q_c_824_n N_VGND_c_838_n 0.0305071f $X=6.46 $Y=0.45 $X2=0 $Y2=0
cc_455 N_Q_c_824_n N_VGND_c_843_n 0.0173469f $X=6.46 $Y=0.45 $X2=0 $Y2=0
cc_456 N_Q_c_824_n N_VGND_c_844_n 0.0110324f $X=6.46 $Y=0.45 $X2=0 $Y2=0
cc_457 N_VGND_c_844_n A_656_47# 0.00250288f $X=6.48 $Y=0 $X2=-0.19 $Y2=-0.245
cc_458 N_VGND_c_844_n A_836_47# 0.00315661f $X=6.48 $Y=0 $X2=-0.19 $Y2=-0.245
