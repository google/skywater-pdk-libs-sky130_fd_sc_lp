* File: sky130_fd_sc_lp__xor3_lp.pxi.spice
* Created: Fri Aug 28 11:37:11 2020
* 
x_PM_SKY130_FD_SC_LP__XOR3_LP%A N_A_M1002_g N_A_M1023_g N_A_M1025_g A
+ N_A_c_194_n N_A_c_195_n PM_SKY130_FD_SC_LP__XOR3_LP%A
x_PM_SKY130_FD_SC_LP__XOR3_LP%A_57_113# N_A_57_113#_M1002_s N_A_57_113#_M1006_d
+ N_A_57_113#_M1023_s N_A_57_113#_M1019_d N_A_57_113#_M1003_g
+ N_A_57_113#_c_233_n N_A_57_113#_M1000_g N_A_57_113#_c_234_n
+ N_A_57_113#_c_235_n N_A_57_113#_c_236_n N_A_57_113#_M1013_g
+ N_A_57_113#_c_237_n N_A_57_113#_c_238_n N_A_57_113#_c_239_n
+ N_A_57_113#_c_263_n N_A_57_113#_c_266_n N_A_57_113#_c_270_p
+ N_A_57_113#_c_292_p N_A_57_113#_c_240_n N_A_57_113#_c_241_n
+ N_A_57_113#_c_242_n N_A_57_113#_c_272_p N_A_57_113#_c_243_n
+ N_A_57_113#_c_247_n N_A_57_113#_c_244_n PM_SKY130_FD_SC_LP__XOR3_LP%A_57_113#
x_PM_SKY130_FD_SC_LP__XOR3_LP%B N_B_M1017_g N_B_M1006_g N_B_M1020_g N_B_c_367_n
+ N_B_c_368_n N_B_c_369_n N_B_M1016_g N_B_c_370_n N_B_M1014_g N_B_M1015_g
+ N_B_c_373_n N_B_M1010_g N_B_c_375_n N_B_c_376_n N_B_c_377_n N_B_c_378_n
+ N_B_c_379_n N_B_c_380_n N_B_c_381_n N_B_c_382_n N_B_c_394_n B N_B_c_383_n
+ N_B_c_384_n N_B_c_385_n N_B_c_386_n PM_SKY130_FD_SC_LP__XOR3_LP%B
x_PM_SKY130_FD_SC_LP__XOR3_LP%A_580_21# N_A_580_21#_M1015_s N_A_580_21#_M1014_s
+ N_A_580_21#_M1009_g N_A_580_21#_c_539_n N_A_580_21#_c_540_n
+ N_A_580_21#_c_541_n N_A_580_21#_c_542_n N_A_580_21#_M1019_g
+ N_A_580_21#_c_543_n N_A_580_21#_M1018_g N_A_580_21#_c_544_n
+ N_A_580_21#_c_555_n N_A_580_21#_M1007_g N_A_580_21#_c_545_n
+ N_A_580_21#_c_546_n N_A_580_21#_c_547_n N_A_580_21#_c_559_n
+ N_A_580_21#_c_548_n N_A_580_21#_c_560_n N_A_580_21#_c_561_n
+ N_A_580_21#_c_549_n N_A_580_21#_c_550_n N_A_580_21#_c_551_n
+ N_A_580_21#_c_552_n N_A_580_21#_c_553_n PM_SKY130_FD_SC_LP__XOR3_LP%A_580_21#
x_PM_SKY130_FD_SC_LP__XOR3_LP%A_1393_300# N_A_1393_300#_M1008_s
+ N_A_1393_300#_M1026_s N_A_1393_300#_M1024_g N_A_1393_300#_M1022_g
+ N_A_1393_300#_c_686_n N_A_1393_300#_c_687_n N_A_1393_300#_c_688_n
+ N_A_1393_300#_c_689_n N_A_1393_300#_c_690_n N_A_1393_300#_c_691_n
+ N_A_1393_300#_c_692_n N_A_1393_300#_c_693_n
+ PM_SKY130_FD_SC_LP__XOR3_LP%A_1393_300#
x_PM_SKY130_FD_SC_LP__XOR3_LP%C N_C_M1005_g N_C_c_770_n N_C_c_779_n N_C_M1012_g
+ N_C_c_780_n N_C_c_781_n N_C_M1026_g N_C_c_771_n N_C_M1008_g N_C_c_772_n
+ N_C_c_773_n N_C_M1001_g N_C_c_774_n N_C_c_775_n N_C_c_783_n N_C_c_784_n C C
+ N_C_c_777_n PM_SKY130_FD_SC_LP__XOR3_LP%C
x_PM_SKY130_FD_SC_LP__XOR3_LP%A_1459_406# N_A_1459_406#_M1005_d
+ N_A_1459_406#_M1024_d N_A_1459_406#_M1021_g N_A_1459_406#_M1011_g
+ N_A_1459_406#_c_861_n N_A_1459_406#_M1004_g N_A_1459_406#_c_869_n
+ N_A_1459_406#_c_870_n N_A_1459_406#_c_871_n N_A_1459_406#_c_862_n
+ N_A_1459_406#_c_863_n N_A_1459_406#_c_864_n N_A_1459_406#_c_872_n
+ N_A_1459_406#_c_873_n N_A_1459_406#_c_874_n N_A_1459_406#_c_865_n
+ N_A_1459_406#_c_866_n N_A_1459_406#_c_867_n
+ PM_SKY130_FD_SC_LP__XOR3_LP%A_1459_406#
x_PM_SKY130_FD_SC_LP__XOR3_LP%VPWR N_VPWR_M1023_d N_VPWR_M1014_d N_VPWR_M1026_d
+ N_VPWR_c_971_n N_VPWR_c_972_n N_VPWR_c_973_n N_VPWR_c_974_n N_VPWR_c_975_n
+ N_VPWR_c_976_n N_VPWR_c_977_n VPWR N_VPWR_c_978_n N_VPWR_c_979_n
+ N_VPWR_c_970_n N_VPWR_c_981_n PM_SKY130_FD_SC_LP__XOR3_LP%VPWR
x_PM_SKY130_FD_SC_LP__XOR3_LP%A_388_419# N_A_388_419#_M1013_d
+ N_A_388_419#_M1016_d N_A_388_419#_M1003_d N_A_388_419#_M1007_d
+ N_A_388_419#_c_1071_n N_A_388_419#_c_1058_n N_A_388_419#_c_1059_n
+ N_A_388_419#_c_1060_n N_A_388_419#_c_1066_n N_A_388_419#_c_1067_n
+ N_A_388_419#_c_1061_n N_A_388_419#_c_1062_n N_A_388_419#_c_1063_n
+ N_A_388_419#_c_1064_n N_A_388_419#_c_1065_n
+ PM_SKY130_FD_SC_LP__XOR3_LP%A_388_419#
x_PM_SKY130_FD_SC_LP__XOR3_LP%A_494_419# N_A_494_419#_M1009_d
+ N_A_494_419#_M1005_s N_A_494_419#_M1017_d N_A_494_419#_M1024_s
+ N_A_494_419#_c_1175_n N_A_494_419#_c_1194_n N_A_494_419#_c_1176_n
+ N_A_494_419#_c_1177_n N_A_494_419#_c_1185_n N_A_494_419#_c_1178_n
+ N_A_494_419#_c_1204_n N_A_494_419#_c_1186_n N_A_494_419#_c_1206_n
+ N_A_494_419#_c_1230_n N_A_494_419#_c_1179_n N_A_494_419#_c_1234_n
+ N_A_494_419#_c_1187_n N_A_494_419#_c_1180_n N_A_494_419#_c_1188_n
+ N_A_494_419#_c_1181_n N_A_494_419#_c_1189_n N_A_494_419#_c_1182_n
+ N_A_494_419#_c_1183_n PM_SKY130_FD_SC_LP__XOR3_LP%A_494_419#
x_PM_SKY130_FD_SC_LP__XOR3_LP%A_855_66# N_A_855_66#_M1018_d N_A_855_66#_M1022_d
+ N_A_855_66#_M1020_d N_A_855_66#_M1012_d N_A_855_66#_c_1320_n
+ N_A_855_66#_c_1321_n N_A_855_66#_c_1322_n N_A_855_66#_c_1323_n
+ N_A_855_66#_c_1324_n N_A_855_66#_c_1325_n N_A_855_66#_c_1326_n
+ N_A_855_66#_c_1329_n N_A_855_66#_c_1353_n N_A_855_66#_c_1380_n
+ PM_SKY130_FD_SC_LP__XOR3_LP%A_855_66#
x_PM_SKY130_FD_SC_LP__XOR3_LP%X N_X_M1004_d N_X_M1021_d N_X_c_1426_n
+ N_X_c_1427_n X X X X X N_X_c_1425_n X PM_SKY130_FD_SC_LP__XOR3_LP%X
x_PM_SKY130_FD_SC_LP__XOR3_LP%VGND N_VGND_M1025_d N_VGND_M1010_d N_VGND_M1001_d
+ N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1496_n N_VGND_c_1451_n
+ N_VGND_c_1452_n N_VGND_c_1453_n N_VGND_c_1454_n N_VGND_c_1455_n VGND
+ N_VGND_c_1456_n N_VGND_c_1457_n N_VGND_c_1458_n N_VGND_c_1459_n
+ PM_SKY130_FD_SC_LP__XOR3_LP%VGND
cc_1 VNB N_A_M1002_g 0.0490716f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.775
cc_2 VNB N_A_M1025_g 0.0426267f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.775
cc_3 VNB N_A_c_194_n 0.00278114f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_4 VNB N_A_c_195_n 0.00873535f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.77
cc_5 VNB N_A_57_113#_M1003_g 0.0179631f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.77
cc_6 VNB N_A_57_113#_c_233_n 0.0169428f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.77
cc_7 VNB N_A_57_113#_c_234_n 0.0182224f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_8 VNB N_A_57_113#_c_235_n 0.071974f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.77
cc_9 VNB N_A_57_113#_c_236_n 0.0162942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_57_113#_c_237_n 0.0249086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_57_113#_c_238_n 0.0097611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_57_113#_c_239_n 0.0213267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_57_113#_c_240_n 0.0101816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_57_113#_c_241_n 0.0404234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_57_113#_c_242_n 0.00395629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_57_113#_c_243_n 0.0149658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_57_113#_c_244_n 0.00615609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_367_n 0.0133726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_c_368_n 0.00953029f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.77
cc_20 VNB N_B_c_369_n 0.0154866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_370_n 0.0624677f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_22 VNB N_B_M1014_g 0.0315532f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.77
cc_23 VNB N_B_M1015_g 0.0233487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_373_n 0.0219075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_M1010_g 0.0249549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_375_n 0.00850143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_376_n 0.00616337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_377_n 0.0113645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_c_378_n 0.0036702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_379_n 0.00376304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_c_380_n 0.038607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_c_381_n 0.00351256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_c_382_n 0.0141208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_383_n 0.0190043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_c_384_n 0.0182877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_c_385_n 0.0198298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_386_n 0.00347574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_580_21#_M1009_g 0.026811f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.775
cc_39 VNB N_A_580_21#_c_539_n 0.0717118f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.775
cc_40 VNB N_A_580_21#_c_540_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_580_21#_c_541_n 0.0231852f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_42 VNB N_A_580_21#_c_542_n 0.00772884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_580_21#_c_543_n 0.0181827f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.77
cc_44 VNB N_A_580_21#_c_544_n 0.0974874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_580_21#_c_545_n 0.00819154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_580_21#_c_546_n 0.004539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_580_21#_c_547_n 0.0232032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_580_21#_c_548_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_580_21#_c_549_n 0.00875234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_580_21#_c_550_n 0.0196991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_580_21#_c_551_n 0.00313656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_580_21#_c_552_n 0.034009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_580_21#_c_553_n 0.0269405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1393_300#_M1022_g 0.0253694f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_55 VNB N_A_1393_300#_c_686_n 0.00464884f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=1.77
cc_56 VNB N_A_1393_300#_c_687_n 0.0199386f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_57 VNB N_A_1393_300#_c_688_n 0.00731168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1393_300#_c_689_n 0.00652155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1393_300#_c_690_n 0.0146308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1393_300#_c_691_n 0.0428055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1393_300#_c_692_n 0.0302023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1393_300#_c_693_n 0.0219154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_C_c_770_n 0.0205956f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.935
cc_64 VNB N_C_c_771_n 0.0177338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_C_c_772_n 0.00566598f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_66 VNB N_C_c_773_n 0.0161613f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_67 VNB N_C_c_774_n 0.0172926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_C_c_775_n 0.0108827f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.77
cc_69 VNB C 0.018789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_C_c_777_n 0.0341801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1459_406#_M1011_g 0.0120894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1459_406#_c_861_n 0.0197276f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.77
cc_73 VNB N_A_1459_406#_c_862_n 0.00845072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1459_406#_c_863_n 0.0622176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1459_406#_c_864_n 0.0104579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1459_406#_c_865_n 6.33388e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1459_406#_c_866_n 0.0595729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1459_406#_c_867_n 0.0476324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VPWR_c_970_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_388_419#_c_1058_n 0.00483482f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.77
cc_81 VNB N_A_388_419#_c_1059_n 0.00192574f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=1.77
cc_82 VNB N_A_388_419#_c_1060_n 0.00912451f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_83 VNB N_A_388_419#_c_1061_n 0.00250318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_388_419#_c_1062_n 0.00798806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_388_419#_c_1063_n 0.00702498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_388_419#_c_1064_n 0.00142512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_388_419#_c_1065_n 0.0044279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_494_419#_c_1175_n 0.00448859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_494_419#_c_1176_n 0.00935506f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_90 VNB N_A_494_419#_c_1177_n 0.00124356f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_91 VNB N_A_494_419#_c_1178_n 0.00320931f $X=-0.19 $Y=-0.245 $X2=1.075
+ $Y2=2.035
cc_92 VNB N_A_494_419#_c_1179_n 0.0140958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_494_419#_c_1180_n 0.0181799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_494_419#_c_1181_n 0.00201017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_494_419#_c_1182_n 0.0118705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_494_419#_c_1183_n 0.0185873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_855_66#_c_1320_n 0.00729583f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.77
cc_98 VNB N_A_855_66#_c_1321_n 0.00259406f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_99 VNB N_A_855_66#_c_1322_n 0.0057969f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.77
cc_100 VNB N_A_855_66#_c_1323_n 0.00772733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_855_66#_c_1324_n 0.00299627f $X=-0.19 $Y=-0.245 $X2=1.075
+ $Y2=1.77
cc_102 VNB N_A_855_66#_c_1325_n 0.0075397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_855_66#_c_1326_n 0.00974428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_X_c_1425_n 0.0476328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1449_n 0.0180096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1450_n 0.0254842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1451_n 0.0209833f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.77
cc_108 VNB N_VGND_c_1452_n 0.130384f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=2.035
cc_109 VNB N_VGND_c_1453_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1454_n 0.0844883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1455_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1456_n 0.03397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1457_n 0.0184869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1458_n 0.61498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1459_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VPB N_A_M1023_g 0.0331287f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.595
cc_117 VPB N_A_c_194_n 0.00483106f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.77
cc_118 VPB N_A_c_195_n 0.041327f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.77
cc_119 VPB N_A_57_113#_M1003_g 0.0476265f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.77
cc_120 VPB N_A_57_113#_c_238_n 0.0283397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_57_113#_c_247_n 0.0311137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_B_M1017_g 0.031702f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=0.775
cc_123 VPB N_B_M1020_g 0.0320864f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.775
cc_124 VPB N_B_M1014_g 0.0443603f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=1.77
cc_125 VPB N_B_c_375_n 0.00956014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_B_c_378_n 0.00121269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_B_c_381_n 0.00222327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_B_c_382_n 0.0216022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_B_c_394_n 0.00511653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_B_c_383_n 0.0315257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_B_c_386_n 0.00180147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_580_21#_M1019_g 0.0382916f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.77
cc_133 VPB N_A_580_21#_c_555_n 0.0294724f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_580_21#_c_545_n 0.0146686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_580_21#_c_546_n 0.00458778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_580_21#_c_547_n 0.00377826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_580_21#_c_559_n 0.0139351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_580_21#_c_560_n 0.00997894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_580_21#_c_561_n 0.0096356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_580_21#_c_550_n 0.0170501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_580_21#_c_551_n 0.00101737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_1393_300#_M1024_g 0.0316797f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=1.605
cc_143 VPB N_A_1393_300#_c_686_n 0.00352117f $X=-0.19 $Y=1.655 $X2=0.755
+ $Y2=1.77
cc_144 VPB N_A_1393_300#_c_687_n 0.0148173f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.77
cc_145 VPB N_A_1393_300#_c_688_n 6.39457e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_1393_300#_c_690_n 0.012601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_C_c_770_n 0.00855652f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.935
cc_148 VPB N_C_c_779_n 0.0237038f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.595
cc_149 VPB N_C_c_780_n 0.0717079f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.605
cc_150 VPB N_C_c_781_n 0.0280988f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.775
cc_151 VPB N_C_c_772_n 0.0094127f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.77
cc_152 VPB N_C_c_783_n 0.0114128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_C_c_784_n 0.0246847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_1459_406#_M1021_g 0.0327175f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=1.605
cc_155 VPB N_A_1459_406#_c_869_n 0.00242135f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.77
cc_156 VPB N_A_1459_406#_c_870_n 0.0219343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_1459_406#_c_871_n 0.00206712f $X=-0.19 $Y=1.655 $X2=1.075
+ $Y2=2.035
cc_158 VPB N_A_1459_406#_c_872_n 0.00139216f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_1459_406#_c_873_n 0.0152745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_1459_406#_c_874_n 0.00116256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_1459_406#_c_866_n 0.0360628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_971_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_972_n 0.010695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_973_n 0.00373081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_974_n 0.0247247f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.035
cc_166 VPB N_VPWR_c_975_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_976_n 0.119654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_977_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_978_n 0.0768151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_979_n 0.032126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_970_n 0.110693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_981_n 0.00533588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_388_419#_c_1066_n 0.00492578f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=1.77
cc_174 VPB N_A_388_419#_c_1067_n 0.00516398f $X=-0.19 $Y=1.655 $X2=1.075
+ $Y2=1.77
cc_175 VPB N_A_388_419#_c_1062_n 0.00324606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_494_419#_c_1175_n 0.00269364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_494_419#_c_1185_n 0.00944235f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=1.77
cc_178 VPB N_A_494_419#_c_1186_n 0.0106471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_494_419#_c_1187_n 0.013188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_494_419#_c_1188_n 0.0021268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_494_419#_c_1189_n 0.0108102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_494_419#_c_1182_n 0.00840161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_855_66#_c_1322_n 0.00586542f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.77
cc_184 VPB N_A_855_66#_c_1323_n 0.0269475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_855_66#_c_1329_n 0.0140193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_X_c_1426_n 0.016079f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.605
cc_187 VPB N_X_c_1427_n 0.0138923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB X 0.0084956f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.77
cc_189 VPB X 0.0343752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_X_c_1425_n 0.0240255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 N_A_M1025_g N_A_57_113#_M1003_g 0.00462012f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_192 N_A_c_194_n N_A_57_113#_M1003_g 0.00789644f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_193 N_A_c_195_n N_A_57_113#_M1003_g 0.00579484f $X=1.005 $Y=1.77 $X2=0 $Y2=0
cc_194 N_A_M1025_g N_A_57_113#_c_235_n 0.0123566f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_195 N_A_M1002_g N_A_57_113#_c_237_n 0.0125582f $X=0.645 $Y=0.775 $X2=0 $Y2=0
cc_196 N_A_M1025_g N_A_57_113#_c_237_n 0.00190675f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_197 N_A_M1002_g N_A_57_113#_c_238_n 0.00755569f $X=0.645 $Y=0.775 $X2=0 $Y2=0
cc_198 N_A_M1023_g N_A_57_113#_c_238_n 0.015055f $X=0.755 $Y=2.595 $X2=0 $Y2=0
cc_199 N_A_M1025_g N_A_57_113#_c_238_n 0.00101457f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_200 N_A_c_194_n N_A_57_113#_c_238_n 0.0406502f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_201 N_A_c_195_n N_A_57_113#_c_238_n 0.0156041f $X=1.005 $Y=1.77 $X2=0 $Y2=0
cc_202 N_A_M1002_g N_A_57_113#_c_239_n 0.0109723f $X=0.645 $Y=0.775 $X2=0 $Y2=0
cc_203 N_A_M1025_g N_A_57_113#_c_239_n 0.0202109f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_204 N_A_c_194_n N_A_57_113#_c_239_n 0.0378199f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_205 N_A_c_195_n N_A_57_113#_c_239_n 0.00176452f $X=1.005 $Y=1.77 $X2=0 $Y2=0
cc_206 N_A_M1023_g N_A_57_113#_c_263_n 0.0211933f $X=0.755 $Y=2.595 $X2=0 $Y2=0
cc_207 N_A_c_194_n N_A_57_113#_c_263_n 0.032007f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_208 N_A_c_195_n N_A_57_113#_c_263_n 0.00112162f $X=1.005 $Y=1.77 $X2=0 $Y2=0
cc_209 N_A_M1023_g N_A_57_113#_c_266_n 0.00500804f $X=0.755 $Y=2.595 $X2=0 $Y2=0
cc_210 N_A_M1025_g N_A_57_113#_c_240_n 0.00522197f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_211 N_A_M1002_g N_A_57_113#_c_243_n 0.0123038f $X=0.645 $Y=0.775 $X2=0 $Y2=0
cc_212 N_A_M1023_g N_A_57_113#_c_247_n 0.0211842f $X=0.755 $Y=2.595 $X2=0 $Y2=0
cc_213 N_A_c_194_n N_VPWR_M1023_d 0.005638f $X=1 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_214 N_A_M1023_g N_VPWR_c_971_n 0.0147781f $X=0.755 $Y=2.595 $X2=0 $Y2=0
cc_215 N_A_M1023_g N_VPWR_c_974_n 0.00840199f $X=0.755 $Y=2.595 $X2=0 $Y2=0
cc_216 N_A_M1023_g N_VPWR_c_970_n 0.00862397f $X=0.755 $Y=2.595 $X2=0 $Y2=0
cc_217 N_A_c_194_n N_A_388_419#_c_1058_n 0.0170572f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_218 N_A_M1002_g N_VGND_c_1449_n 0.0015588f $X=0.645 $Y=0.775 $X2=0 $Y2=0
cc_219 N_A_M1025_g N_VGND_c_1449_n 0.0112965f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_220 N_A_M1002_g N_VGND_c_1456_n 0.00430863f $X=0.645 $Y=0.775 $X2=0 $Y2=0
cc_221 N_A_M1025_g N_VGND_c_1456_n 0.00372658f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_222 N_A_M1002_g N_VGND_c_1458_n 0.00486331f $X=0.645 $Y=0.775 $X2=0 $Y2=0
cc_223 N_A_M1025_g N_VGND_c_1458_n 0.00408518f $X=1.005 $Y=0.775 $X2=0 $Y2=0
cc_224 N_A_57_113#_c_270_p N_B_M1017_g 0.0212532f $X=3.51 $Y=2.98 $X2=0 $Y2=0
cc_225 N_A_57_113#_c_270_p N_B_M1020_g 6.06832e-19 $X=3.51 $Y=2.98 $X2=0 $Y2=0
cc_226 N_A_57_113#_c_272_p N_B_M1020_g 0.00150006f $X=3.675 $Y=2.745 $X2=0 $Y2=0
cc_227 N_A_57_113#_M1003_g N_B_c_375_n 0.0597371f $X=1.815 $Y=2.595 $X2=0 $Y2=0
cc_228 N_A_57_113#_c_234_n N_B_c_375_n 0.0143106f $X=2.39 $Y=1.17 $X2=0 $Y2=0
cc_229 N_A_57_113#_c_244_n N_B_c_379_n 0.00211868f $X=3.985 $Y=0.35 $X2=0 $Y2=0
cc_230 N_A_57_113#_c_244_n N_B_c_380_n 7.69799e-19 $X=3.985 $Y=0.35 $X2=0 $Y2=0
cc_231 N_A_57_113#_c_241_n N_B_c_384_n 0.00371137f $X=3.82 $Y=0.35 $X2=0 $Y2=0
cc_232 N_A_57_113#_c_244_n N_B_c_384_n 0.00380153f $X=3.985 $Y=0.35 $X2=0 $Y2=0
cc_233 N_A_57_113#_c_236_n N_A_580_21#_M1009_g 0.0107801f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_234 N_A_57_113#_c_241_n N_A_580_21#_M1009_g 0.0130696f $X=3.82 $Y=0.35 $X2=0
+ $Y2=0
cc_235 N_A_57_113#_c_241_n N_A_580_21#_c_539_n 0.013467f $X=3.82 $Y=0.35 $X2=0
+ $Y2=0
cc_236 N_A_57_113#_c_244_n N_A_580_21#_c_539_n 0.00516063f $X=3.985 $Y=0.35
+ $X2=0 $Y2=0
cc_237 N_A_57_113#_c_241_n N_A_580_21#_c_541_n 0.00189786f $X=3.82 $Y=0.35 $X2=0
+ $Y2=0
cc_238 N_A_57_113#_c_234_n N_A_580_21#_c_542_n 0.0107801f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_239 N_A_57_113#_c_270_p N_A_580_21#_M1019_g 0.0186796f $X=3.51 $Y=2.98 $X2=0
+ $Y2=0
cc_240 N_A_57_113#_c_272_p N_A_580_21#_M1019_g 0.0232836f $X=3.675 $Y=2.745
+ $X2=0 $Y2=0
cc_241 N_A_57_113#_c_241_n N_A_580_21#_c_543_n 2.21879e-19 $X=3.82 $Y=0.35 $X2=0
+ $Y2=0
cc_242 N_A_57_113#_c_244_n N_A_580_21#_c_543_n 0.00781411f $X=3.985 $Y=0.35
+ $X2=0 $Y2=0
cc_243 N_A_57_113#_c_263_n N_VPWR_M1023_d 0.0260509f $X=1.365 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_244 N_A_57_113#_c_266_n N_VPWR_M1023_d 0.0127439f $X=1.45 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_245 N_A_57_113#_c_270_p N_VPWR_M1023_d 0.00463221f $X=3.51 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_246 N_A_57_113#_c_292_p N_VPWR_M1023_d 0.00476969f $X=1.535 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_57_113#_M1003_g N_VPWR_c_971_n 0.00377986f $X=1.815 $Y=2.595 $X2=0
+ $Y2=0
cc_248 N_A_57_113#_c_263_n N_VPWR_c_971_n 0.0204369f $X=1.365 $Y=2.415 $X2=0
+ $Y2=0
cc_249 N_A_57_113#_c_266_n N_VPWR_c_971_n 0.0157123f $X=1.45 $Y=2.895 $X2=0
+ $Y2=0
cc_250 N_A_57_113#_c_292_p N_VPWR_c_971_n 0.0138719f $X=1.535 $Y=2.98 $X2=0
+ $Y2=0
cc_251 N_A_57_113#_c_247_n N_VPWR_c_971_n 0.0256963f $X=0.46 $Y=2.415 $X2=0
+ $Y2=0
cc_252 N_A_57_113#_c_247_n N_VPWR_c_974_n 0.0238035f $X=0.46 $Y=2.415 $X2=0
+ $Y2=0
cc_253 N_A_57_113#_M1003_g N_VPWR_c_976_n 0.00599941f $X=1.815 $Y=2.595 $X2=0
+ $Y2=0
cc_254 N_A_57_113#_c_270_p N_VPWR_c_976_n 0.12864f $X=3.51 $Y=2.98 $X2=0 $Y2=0
cc_255 N_A_57_113#_c_292_p N_VPWR_c_976_n 0.011231f $X=1.535 $Y=2.98 $X2=0 $Y2=0
cc_256 N_A_57_113#_M1023_s N_VPWR_c_970_n 0.0023218f $X=0.345 $Y=2.095 $X2=0
+ $Y2=0
cc_257 N_A_57_113#_M1019_d N_VPWR_c_970_n 0.0113391f $X=3.535 $Y=2.095 $X2=0
+ $Y2=0
cc_258 N_A_57_113#_M1003_g N_VPWR_c_970_n 0.00935477f $X=1.815 $Y=2.595 $X2=0
+ $Y2=0
cc_259 N_A_57_113#_c_263_n N_VPWR_c_970_n 0.0129302f $X=1.365 $Y=2.415 $X2=0
+ $Y2=0
cc_260 N_A_57_113#_c_270_p N_VPWR_c_970_n 0.0831141f $X=3.51 $Y=2.98 $X2=0 $Y2=0
cc_261 N_A_57_113#_c_292_p N_VPWR_c_970_n 0.00657784f $X=1.535 $Y=2.98 $X2=0
+ $Y2=0
cc_262 N_A_57_113#_c_247_n N_VPWR_c_970_n 0.0148296f $X=0.46 $Y=2.415 $X2=0
+ $Y2=0
cc_263 N_A_57_113#_c_270_p N_A_388_419#_M1003_d 0.00340092f $X=3.51 $Y=2.98
+ $X2=0 $Y2=0
cc_264 N_A_57_113#_c_233_n N_A_388_419#_c_1071_n 0.0100848f $X=2.075 $Y=1.095
+ $X2=0 $Y2=0
cc_265 N_A_57_113#_c_240_n N_A_388_419#_c_1071_n 0.0140162f $X=1.65 $Y=1.095
+ $X2=0 $Y2=0
cc_266 N_A_57_113#_c_241_n N_A_388_419#_c_1071_n 0.00888218f $X=3.82 $Y=0.35
+ $X2=0 $Y2=0
cc_267 N_A_57_113#_M1003_g N_A_388_419#_c_1058_n 0.0477782f $X=1.815 $Y=2.595
+ $X2=0 $Y2=0
cc_268 N_A_57_113#_c_233_n N_A_388_419#_c_1058_n 0.00307528f $X=2.075 $Y=1.095
+ $X2=0 $Y2=0
cc_269 N_A_57_113#_c_234_n N_A_388_419#_c_1058_n 0.00601776f $X=2.39 $Y=1.17
+ $X2=0 $Y2=0
cc_270 N_A_57_113#_c_235_n N_A_388_419#_c_1058_n 0.0190074f $X=2.15 $Y=1.17
+ $X2=0 $Y2=0
cc_271 N_A_57_113#_c_236_n N_A_388_419#_c_1058_n 0.00193958f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_272 N_A_57_113#_c_263_n N_A_388_419#_c_1058_n 0.00755511f $X=1.365 $Y=2.415
+ $X2=0 $Y2=0
cc_273 N_A_57_113#_c_266_n N_A_388_419#_c_1058_n 0.00852076f $X=1.45 $Y=2.895
+ $X2=0 $Y2=0
cc_274 N_A_57_113#_c_270_p N_A_388_419#_c_1058_n 0.0153084f $X=3.51 $Y=2.98
+ $X2=0 $Y2=0
cc_275 N_A_57_113#_c_240_n N_A_388_419#_c_1058_n 0.0317277f $X=1.65 $Y=1.095
+ $X2=0 $Y2=0
cc_276 N_A_57_113#_c_234_n N_A_388_419#_c_1059_n 0.00187676f $X=2.39 $Y=1.17
+ $X2=0 $Y2=0
cc_277 N_A_57_113#_c_236_n N_A_388_419#_c_1059_n 0.00851322f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_278 N_A_57_113#_c_241_n N_A_388_419#_c_1059_n 0.00681218f $X=3.82 $Y=0.35
+ $X2=0 $Y2=0
cc_279 N_A_57_113#_c_233_n N_A_388_419#_c_1061_n 0.00100945f $X=2.075 $Y=1.095
+ $X2=0 $Y2=0
cc_280 N_A_57_113#_c_236_n N_A_388_419#_c_1061_n 0.00485703f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_281 N_A_57_113#_c_241_n N_A_388_419#_c_1061_n 0.0188733f $X=3.82 $Y=0.35
+ $X2=0 $Y2=0
cc_282 N_A_57_113#_M1006_d N_A_388_419#_c_1063_n 0.00440588f $X=3.765 $Y=0.625
+ $X2=0 $Y2=0
cc_283 N_A_57_113#_c_241_n N_A_388_419#_c_1063_n 0.0258311f $X=3.82 $Y=0.35
+ $X2=0 $Y2=0
cc_284 N_A_57_113#_c_244_n N_A_388_419#_c_1063_n 0.0137981f $X=3.985 $Y=0.35
+ $X2=0 $Y2=0
cc_285 N_A_57_113#_c_233_n N_A_388_419#_c_1064_n 0.00144221f $X=2.075 $Y=1.095
+ $X2=0 $Y2=0
cc_286 N_A_57_113#_c_234_n N_A_388_419#_c_1064_n 0.00137405f $X=2.39 $Y=1.17
+ $X2=0 $Y2=0
cc_287 N_A_57_113#_c_236_n N_A_388_419#_c_1064_n 5.72254e-19 $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_288 N_A_57_113#_c_240_n N_A_388_419#_c_1064_n 0.00131136f $X=1.65 $Y=1.095
+ $X2=0 $Y2=0
cc_289 N_A_57_113#_c_241_n N_A_388_419#_c_1064_n 0.0030356f $X=3.82 $Y=0.35
+ $X2=0 $Y2=0
cc_290 N_A_57_113#_c_270_p N_A_494_419#_M1017_d 0.0230583f $X=3.51 $Y=2.98 $X2=0
+ $Y2=0
cc_291 N_A_57_113#_M1003_g N_A_494_419#_c_1175_n 3.11561e-19 $X=1.815 $Y=2.595
+ $X2=0 $Y2=0
cc_292 N_A_57_113#_c_235_n N_A_494_419#_c_1175_n 7.59242e-19 $X=2.15 $Y=1.17
+ $X2=0 $Y2=0
cc_293 N_A_57_113#_c_270_p N_A_494_419#_c_1194_n 0.0208598f $X=3.51 $Y=2.98
+ $X2=0 $Y2=0
cc_294 N_A_57_113#_c_234_n N_A_494_419#_c_1177_n 0.00559204f $X=2.39 $Y=1.17
+ $X2=0 $Y2=0
cc_295 N_A_57_113#_c_235_n N_A_494_419#_c_1177_n 4.52039e-19 $X=2.15 $Y=1.17
+ $X2=0 $Y2=0
cc_296 N_A_57_113#_M1019_d N_A_494_419#_c_1185_n 0.0117017f $X=3.535 $Y=2.095
+ $X2=0 $Y2=0
cc_297 N_A_57_113#_c_270_p N_A_494_419#_c_1185_n 0.0169719f $X=3.51 $Y=2.98
+ $X2=0 $Y2=0
cc_298 N_A_57_113#_c_272_p N_A_494_419#_c_1185_n 0.0208964f $X=3.675 $Y=2.745
+ $X2=0 $Y2=0
cc_299 N_A_57_113#_c_234_n N_A_494_419#_c_1178_n 3.2296e-19 $X=2.39 $Y=1.17
+ $X2=0 $Y2=0
cc_300 N_A_57_113#_c_236_n N_A_494_419#_c_1178_n 0.00146273f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_301 N_A_57_113#_c_241_n N_A_494_419#_c_1178_n 0.023002f $X=3.82 $Y=0.35 $X2=0
+ $Y2=0
cc_302 N_A_57_113#_c_244_n N_A_494_419#_c_1178_n 0.00176513f $X=3.985 $Y=0.35
+ $X2=0 $Y2=0
cc_303 N_A_57_113#_M1019_d N_A_494_419#_c_1204_n 0.00724135f $X=3.535 $Y=2.095
+ $X2=0 $Y2=0
cc_304 N_A_57_113#_c_272_p N_A_494_419#_c_1204_n 0.0341205f $X=3.675 $Y=2.745
+ $X2=0 $Y2=0
cc_305 N_A_57_113#_M1019_d N_A_494_419#_c_1206_n 0.00248178f $X=3.535 $Y=2.095
+ $X2=0 $Y2=0
cc_306 N_A_57_113#_c_270_p N_A_494_419#_c_1206_n 0.014682f $X=3.51 $Y=2.98 $X2=0
+ $Y2=0
cc_307 N_A_57_113#_c_244_n N_A_855_66#_c_1320_n 0.0141997f $X=3.985 $Y=0.35
+ $X2=0 $Y2=0
cc_308 N_A_57_113#_c_240_n N_VGND_M1025_d 0.0121884f $X=1.65 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_309 N_A_57_113#_c_237_n N_VGND_c_1449_n 0.0123792f $X=0.43 $Y=0.775 $X2=0
+ $Y2=0
cc_310 N_A_57_113#_c_239_n N_VGND_c_1449_n 0.0246161f $X=1.565 $Y=1.26 $X2=0
+ $Y2=0
cc_311 N_A_57_113#_c_240_n N_VGND_c_1449_n 0.0354987f $X=1.65 $Y=1.095 $X2=0
+ $Y2=0
cc_312 N_A_57_113#_c_242_n N_VGND_c_1449_n 0.0144411f $X=1.735 $Y=0.35 $X2=0
+ $Y2=0
cc_313 N_A_57_113#_c_241_n N_VGND_c_1452_n 0.125951f $X=3.82 $Y=0.35 $X2=0 $Y2=0
cc_314 N_A_57_113#_c_242_n N_VGND_c_1452_n 0.0114622f $X=1.735 $Y=0.35 $X2=0
+ $Y2=0
cc_315 N_A_57_113#_c_244_n N_VGND_c_1452_n 0.0212541f $X=3.985 $Y=0.35 $X2=0
+ $Y2=0
cc_316 N_A_57_113#_c_237_n N_VGND_c_1456_n 0.00805126f $X=0.43 $Y=0.775 $X2=0
+ $Y2=0
cc_317 N_A_57_113#_c_237_n N_VGND_c_1458_n 0.0106012f $X=0.43 $Y=0.775 $X2=0
+ $Y2=0
cc_318 N_A_57_113#_c_241_n N_VGND_c_1458_n 0.0741314f $X=3.82 $Y=0.35 $X2=0
+ $Y2=0
cc_319 N_A_57_113#_c_242_n N_VGND_c_1458_n 0.00657784f $X=1.735 $Y=0.35 $X2=0
+ $Y2=0
cc_320 N_A_57_113#_c_244_n N_VGND_c_1458_n 0.0111793f $X=3.985 $Y=0.35 $X2=0
+ $Y2=0
cc_321 N_B_c_384_n N_A_580_21#_M1009_g 0.00946658f $X=3.78 $Y=1.155 $X2=0 $Y2=0
cc_322 N_B_c_384_n N_A_580_21#_c_539_n 0.00737233f $X=3.78 $Y=1.155 $X2=0 $Y2=0
cc_323 N_B_c_379_n N_A_580_21#_c_541_n 2.38084e-19 $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_324 N_B_c_384_n N_A_580_21#_c_541_n 0.0114393f $X=3.78 $Y=1.155 $X2=0 $Y2=0
cc_325 N_B_c_383_n N_A_580_21#_c_542_n 0.00618171f $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_326 N_B_c_386_n N_A_580_21#_c_542_n 0.0015841f $X=3.235 $Y=1.722 $X2=0 $Y2=0
cc_327 N_B_M1020_g N_A_580_21#_M1019_g 0.0101603f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_328 N_B_c_378_n N_A_580_21#_M1019_g 0.00459218f $X=3.615 $Y=1.73 $X2=0 $Y2=0
cc_329 N_B_c_383_n N_A_580_21#_M1019_g 0.00108894f $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_330 N_B_c_369_n N_A_580_21#_c_543_n 0.00762566f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_331 N_B_c_381_n N_A_580_21#_c_543_n 9.94976e-19 $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_332 N_B_c_382_n N_A_580_21#_c_543_n 0.00212288f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_333 N_B_c_384_n N_A_580_21#_c_543_n 0.00863061f $X=3.78 $Y=1.155 $X2=0 $Y2=0
cc_334 N_B_c_369_n N_A_580_21#_c_544_n 0.0102019f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_335 N_B_M1020_g N_A_580_21#_c_555_n 0.0390431f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_336 N_B_c_367_n N_A_580_21#_c_555_n 0.00128586f $X=4.715 $Y=1.165 $X2=0 $Y2=0
cc_337 N_B_c_370_n N_A_580_21#_c_545_n 0.00908257f $X=5.875 $Y=1.165 $X2=0 $Y2=0
cc_338 N_B_c_376_n N_A_580_21#_c_546_n 0.00908257f $X=4.79 $Y=1.165 $X2=0 $Y2=0
cc_339 N_B_c_382_n N_A_580_21#_c_546_n 0.00914448f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_340 N_B_c_378_n N_A_580_21#_c_547_n 0.00979864f $X=3.615 $Y=1.73 $X2=0 $Y2=0
cc_341 N_B_c_379_n N_A_580_21#_c_547_n 0.00350138f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_342 N_B_c_380_n N_A_580_21#_c_547_n 0.0114393f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_343 N_B_c_383_n N_A_580_21#_c_547_n 0.0201143f $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_344 N_B_c_386_n N_A_580_21#_c_547_n 3.85829e-19 $X=3.235 $Y=1.722 $X2=0 $Y2=0
cc_345 N_B_c_378_n N_A_580_21#_c_559_n 0.010993f $X=3.615 $Y=1.73 $X2=0 $Y2=0
cc_346 N_B_c_382_n N_A_580_21#_c_559_n 0.0101603f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_347 N_B_M1020_g N_A_580_21#_c_560_n 0.00134555f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_348 N_B_M1014_g N_A_580_21#_c_561_n 0.0200019f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_349 N_B_c_369_n N_A_580_21#_c_549_n 3.36415e-19 $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_350 N_B_c_370_n N_A_580_21#_c_549_n 0.0154005f $X=5.875 $Y=1.165 $X2=0 $Y2=0
cc_351 N_B_M1014_g N_A_580_21#_c_549_n 0.00458638f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_352 N_B_M1015_g N_A_580_21#_c_549_n 0.00579762f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_353 N_B_c_370_n N_A_580_21#_c_550_n 0.0212171f $X=5.875 $Y=1.165 $X2=0 $Y2=0
cc_354 N_B_M1014_g N_A_580_21#_c_550_n 0.0170391f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_355 N_B_c_370_n N_A_580_21#_c_551_n 0.00216696f $X=5.875 $Y=1.165 $X2=0 $Y2=0
cc_356 N_B_M1014_g N_A_580_21#_c_551_n 0.00211019f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_357 N_B_c_369_n N_A_580_21#_c_552_n 0.00260557f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_358 N_B_c_370_n N_A_580_21#_c_552_n 0.00644864f $X=5.875 $Y=1.165 $X2=0 $Y2=0
cc_359 N_B_M1015_g N_A_580_21#_c_552_n 0.00580119f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_360 N_B_c_369_n N_A_580_21#_c_553_n 0.00133673f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_361 N_B_c_370_n N_A_580_21#_c_553_n 0.0107366f $X=5.875 $Y=1.165 $X2=0 $Y2=0
cc_362 N_B_M1015_g N_A_580_21#_c_553_n 0.0116901f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_363 N_B_M1010_g N_A_580_21#_c_553_n 0.0012482f $X=6.51 $Y=0.655 $X2=0 $Y2=0
cc_364 N_B_M1014_g N_VPWR_c_972_n 0.0253327f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_365 N_B_M1017_g N_VPWR_c_976_n 0.00599941f $X=2.345 $Y=2.595 $X2=0 $Y2=0
cc_366 N_B_M1020_g N_VPWR_c_976_n 0.00599892f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_367 N_B_M1014_g N_VPWR_c_976_n 0.00539993f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_368 N_B_M1017_g N_VPWR_c_970_n 0.00935477f $X=2.345 $Y=2.595 $X2=0 $Y2=0
cc_369 N_B_M1020_g N_VPWR_c_970_n 0.00865575f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_370 N_B_M1014_g N_VPWR_c_970_n 0.00846827f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_371 N_B_M1017_g N_A_388_419#_c_1058_n 0.0190902f $X=2.345 $Y=2.595 $X2=0
+ $Y2=0
cc_372 N_B_c_375_n N_A_388_419#_c_1058_n 0.00978604f $X=2.47 $Y=1.73 $X2=0 $Y2=0
cc_373 N_B_c_375_n N_A_388_419#_c_1059_n 0.00165457f $X=2.47 $Y=1.73 $X2=0 $Y2=0
cc_374 N_B_c_369_n N_A_388_419#_c_1060_n 0.00664478f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_375 N_B_c_370_n N_A_388_419#_c_1060_n 0.0017289f $X=5.875 $Y=1.165 $X2=0
+ $Y2=0
cc_376 N_B_c_383_n N_A_388_419#_c_1061_n 4.58149e-19 $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_377 N_B_c_369_n N_A_388_419#_c_1062_n 0.00120249f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_378 N_B_c_370_n N_A_388_419#_c_1062_n 0.015422f $X=5.875 $Y=1.165 $X2=0 $Y2=0
cc_379 N_B_c_385_n N_A_388_419#_c_1062_n 8.90097e-19 $X=4.32 $Y=1.565 $X2=0
+ $Y2=0
cc_380 N_B_c_367_n N_A_388_419#_c_1063_n 0.00122525f $X=4.715 $Y=1.165 $X2=0
+ $Y2=0
cc_381 N_B_c_369_n N_A_388_419#_c_1063_n 0.00639141f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_382 N_B_c_378_n N_A_388_419#_c_1063_n 0.00674079f $X=3.615 $Y=1.73 $X2=0
+ $Y2=0
cc_383 N_B_c_379_n N_A_388_419#_c_1063_n 0.0133185f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_384 N_B_c_381_n N_A_388_419#_c_1063_n 0.0121827f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_385 N_B_c_382_n N_A_388_419#_c_1063_n 0.00274583f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_386 N_B_c_384_n N_A_388_419#_c_1063_n 0.00727252f $X=3.78 $Y=1.155 $X2=0
+ $Y2=0
cc_387 N_B_c_386_n N_A_388_419#_c_1063_n 0.00105075f $X=3.235 $Y=1.722 $X2=0
+ $Y2=0
cc_388 N_B_c_370_n N_A_388_419#_c_1065_n 3.9213e-19 $X=5.875 $Y=1.165 $X2=0
+ $Y2=0
cc_389 N_B_M1017_g N_A_494_419#_c_1175_n 0.00610891f $X=2.345 $Y=2.595 $X2=0
+ $Y2=0
cc_390 N_B_c_375_n N_A_494_419#_c_1175_n 0.00637055f $X=2.47 $Y=1.73 $X2=0 $Y2=0
cc_391 N_B_c_383_n N_A_494_419#_c_1175_n 0.013381f $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_392 N_B_c_386_n N_A_494_419#_c_1175_n 0.025032f $X=3.235 $Y=1.722 $X2=0 $Y2=0
cc_393 N_B_M1017_g N_A_494_419#_c_1194_n 0.0115598f $X=2.345 $Y=2.595 $X2=0
+ $Y2=0
cc_394 N_B_c_378_n N_A_494_419#_c_1176_n 0.0132656f $X=3.615 $Y=1.73 $X2=0 $Y2=0
cc_395 N_B_c_379_n N_A_494_419#_c_1176_n 0.0137327f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_396 N_B_c_380_n N_A_494_419#_c_1176_n 0.00104973f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_397 N_B_c_383_n N_A_494_419#_c_1176_n 0.0077418f $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_398 N_B_c_386_n N_A_494_419#_c_1176_n 0.0328229f $X=3.235 $Y=1.722 $X2=0
+ $Y2=0
cc_399 N_B_M1020_g N_A_494_419#_c_1185_n 0.0070659f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_400 N_B_c_380_n N_A_494_419#_c_1185_n 9.89875e-19 $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_401 N_B_c_381_n N_A_494_419#_c_1185_n 0.0197713f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_402 N_B_c_394_n N_A_494_419#_c_1185_n 0.0267647f $X=3.78 $Y=1.73 $X2=0 $Y2=0
cc_403 N_B_c_383_n N_A_494_419#_c_1185_n 0.00601241f $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_404 N_B_c_386_n N_A_494_419#_c_1185_n 0.0608605f $X=3.235 $Y=1.722 $X2=0
+ $Y2=0
cc_405 N_B_c_379_n N_A_494_419#_c_1178_n 0.00223444f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_406 N_B_c_384_n N_A_494_419#_c_1178_n 0.0130485f $X=3.78 $Y=1.155 $X2=0 $Y2=0
cc_407 N_B_M1020_g N_A_494_419#_c_1204_n 0.0199184f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_408 N_B_M1020_g N_A_494_419#_c_1186_n 0.0163735f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_409 N_B_M1014_g N_A_494_419#_c_1186_n 0.0103926f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_410 N_B_M1020_g N_A_494_419#_c_1206_n 0.00305008f $X=4.28 $Y=2.595 $X2=0
+ $Y2=0
cc_411 N_B_M1014_g N_A_494_419#_c_1230_n 0.0545171f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_412 N_B_M1014_g N_A_494_419#_c_1179_n 0.00417452f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_413 N_B_c_373_n N_A_494_419#_c_1179_n 0.0257359f $X=6.435 $Y=1.165 $X2=0
+ $Y2=0
cc_414 N_B_c_377_n N_A_494_419#_c_1179_n 0.00863921f $X=6.05 $Y=1.165 $X2=0
+ $Y2=0
cc_415 N_B_M1014_g N_A_494_419#_c_1234_n 0.00174827f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_416 N_B_c_377_n N_A_494_419#_c_1234_n 0.0052134f $X=6.05 $Y=1.165 $X2=0 $Y2=0
cc_417 N_B_M1017_g N_A_494_419#_c_1188_n 0.0061793f $X=2.345 $Y=2.595 $X2=0
+ $Y2=0
cc_418 N_B_c_383_n N_A_494_419#_c_1188_n 0.00779995f $X=2.88 $Y=1.73 $X2=0 $Y2=0
cc_419 N_B_M1014_g N_A_494_419#_c_1182_n 0.0125381f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_420 N_B_M1010_g N_A_494_419#_c_1183_n 0.00740689f $X=6.51 $Y=0.655 $X2=0
+ $Y2=0
cc_421 N_B_c_369_n N_A_855_66#_c_1320_n 0.00804057f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_422 N_B_c_367_n N_A_855_66#_c_1321_n 0.00346016f $X=4.715 $Y=1.165 $X2=0
+ $Y2=0
cc_423 N_B_c_368_n N_A_855_66#_c_1321_n 0.0068546f $X=4.485 $Y=1.165 $X2=0 $Y2=0
cc_424 N_B_c_369_n N_A_855_66#_c_1321_n 0.00112909f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_425 N_B_c_379_n N_A_855_66#_c_1321_n 0.00244935f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_426 N_B_c_380_n N_A_855_66#_c_1321_n 4.00543e-19 $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_427 N_B_M1020_g N_A_855_66#_c_1322_n 0.0130664f $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_428 N_B_c_367_n N_A_855_66#_c_1322_n 6.70359e-19 $X=4.715 $Y=1.165 $X2=0
+ $Y2=0
cc_429 N_B_c_379_n N_A_855_66#_c_1322_n 0.00505748f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_430 N_B_c_381_n N_A_855_66#_c_1322_n 0.0260181f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_431 N_B_c_382_n N_A_855_66#_c_1322_n 0.00191313f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_432 N_B_c_385_n N_A_855_66#_c_1322_n 0.00812108f $X=4.32 $Y=1.565 $X2=0 $Y2=0
cc_433 N_B_c_367_n N_A_855_66#_c_1324_n 0.00431458f $X=4.715 $Y=1.165 $X2=0
+ $Y2=0
cc_434 N_B_c_384_n N_A_855_66#_c_1324_n 0.00516811f $X=3.78 $Y=1.155 $X2=0 $Y2=0
cc_435 N_B_c_367_n N_A_855_66#_c_1325_n 0.00501037f $X=4.715 $Y=1.165 $X2=0
+ $Y2=0
cc_436 N_B_c_368_n N_A_855_66#_c_1325_n 9.32595e-19 $X=4.485 $Y=1.165 $X2=0
+ $Y2=0
cc_437 N_B_c_376_n N_A_855_66#_c_1325_n 0.0023011f $X=4.79 $Y=1.165 $X2=0 $Y2=0
cc_438 N_B_c_379_n N_A_855_66#_c_1325_n 0.00743934f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_439 N_B_c_380_n N_A_855_66#_c_1325_n 0.00125059f $X=3.78 $Y=1.32 $X2=0 $Y2=0
cc_440 N_B_c_381_n N_A_855_66#_c_1325_n 0.00628078f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_441 N_B_c_385_n N_A_855_66#_c_1325_n 0.00941298f $X=4.32 $Y=1.565 $X2=0 $Y2=0
cc_442 N_B_M1014_g N_A_855_66#_c_1329_n 0.0102474f $X=6 $Y=2.48 $X2=0 $Y2=0
cc_443 N_B_M1020_g N_A_855_66#_c_1353_n 3.42756e-19 $X=4.28 $Y=2.595 $X2=0 $Y2=0
cc_444 N_B_c_381_n N_A_855_66#_c_1353_n 2.38241e-19 $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_445 N_B_c_382_n N_A_855_66#_c_1353_n 0.0018149f $X=4.32 $Y=1.73 $X2=0 $Y2=0
cc_446 N_B_M1015_g N_VGND_c_1450_n 0.00180305f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_447 N_B_M1010_g N_VGND_c_1450_n 0.0138255f $X=6.51 $Y=0.655 $X2=0 $Y2=0
cc_448 N_B_M1015_g N_VGND_c_1452_n 0.00500171f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_449 N_B_M1010_g N_VGND_c_1452_n 0.00435433f $X=6.51 $Y=0.655 $X2=0 $Y2=0
cc_450 N_B_c_369_n N_VGND_c_1458_n 9.39239e-19 $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_451 N_B_M1015_g N_VGND_c_1458_n 0.0052212f $X=6.15 $Y=0.655 $X2=0 $Y2=0
cc_452 N_B_M1010_g N_VGND_c_1458_n 0.0043858f $X=6.51 $Y=0.655 $X2=0 $Y2=0
cc_453 N_A_580_21#_M1019_g N_VPWR_c_976_n 0.00599906f $X=3.41 $Y=2.595 $X2=0
+ $Y2=0
cc_454 N_A_580_21#_c_555_n N_VPWR_c_976_n 0.00599941f $X=4.82 $Y=2.08 $X2=0
+ $Y2=0
cc_455 N_A_580_21#_M1019_g N_VPWR_c_970_n 0.010023f $X=3.41 $Y=2.595 $X2=0 $Y2=0
cc_456 N_A_580_21#_c_555_n N_VPWR_c_970_n 0.00938086f $X=4.82 $Y=2.08 $X2=0
+ $Y2=0
cc_457 N_A_580_21#_M1009_g N_A_388_419#_c_1058_n 3.76604e-19 $X=2.975 $Y=0.775
+ $X2=0 $Y2=0
cc_458 N_A_580_21#_c_544_n N_A_388_419#_c_1060_n 0.00619022f $X=5.35 $Y=0.18
+ $X2=0 $Y2=0
cc_459 N_A_580_21#_c_546_n N_A_388_419#_c_1060_n 0.0012462f $X=4.945 $Y=1.705
+ $X2=0 $Y2=0
cc_460 N_A_580_21#_c_549_n N_A_388_419#_c_1060_n 0.00445175f $X=5.645 $Y=1.45
+ $X2=0 $Y2=0
cc_461 N_A_580_21#_c_553_n N_A_388_419#_c_1060_n 0.0144944f $X=5.645 $Y=0.575
+ $X2=0 $Y2=0
cc_462 N_A_580_21#_c_555_n N_A_388_419#_c_1066_n 0.00655352f $X=4.82 $Y=2.08
+ $X2=0 $Y2=0
cc_463 N_A_580_21#_c_545_n N_A_388_419#_c_1066_n 0.00504266f $X=5.305 $Y=1.705
+ $X2=0 $Y2=0
cc_464 N_A_580_21#_c_561_n N_A_388_419#_c_1066_n 0.0476794f $X=5.645 $Y=2.125
+ $X2=0 $Y2=0
cc_465 N_A_580_21#_M1009_g N_A_388_419#_c_1061_n 0.00221303f $X=2.975 $Y=0.775
+ $X2=0 $Y2=0
cc_466 N_A_580_21#_c_545_n N_A_388_419#_c_1062_n 0.0124048f $X=5.305 $Y=1.705
+ $X2=0 $Y2=0
cc_467 N_A_580_21#_c_560_n N_A_388_419#_c_1062_n 0.00655352f $X=4.82 $Y=1.955
+ $X2=0 $Y2=0
cc_468 N_A_580_21#_c_561_n N_A_388_419#_c_1062_n 0.0083691f $X=5.645 $Y=2.125
+ $X2=0 $Y2=0
cc_469 N_A_580_21#_c_549_n N_A_388_419#_c_1062_n 0.0149659f $X=5.645 $Y=1.45
+ $X2=0 $Y2=0
cc_470 N_A_580_21#_c_550_n N_A_388_419#_c_1062_n 0.00124625f $X=5.47 $Y=1.615
+ $X2=0 $Y2=0
cc_471 N_A_580_21#_c_551_n N_A_388_419#_c_1062_n 0.0236241f $X=5.645 $Y=1.615
+ $X2=0 $Y2=0
cc_472 N_A_580_21#_M1009_g N_A_388_419#_c_1063_n 0.0059639f $X=2.975 $Y=0.775
+ $X2=0 $Y2=0
cc_473 N_A_580_21#_c_541_n N_A_388_419#_c_1063_n 0.00120735f $X=3.255 $Y=1.195
+ $X2=0 $Y2=0
cc_474 N_A_580_21#_c_543_n N_A_388_419#_c_1063_n 0.00685902f $X=4.2 $Y=0.255
+ $X2=0 $Y2=0
cc_475 N_A_580_21#_c_544_n N_A_388_419#_c_1063_n 0.00131951f $X=5.35 $Y=0.18
+ $X2=0 $Y2=0
cc_476 N_A_580_21#_c_546_n N_A_388_419#_c_1063_n 2.17538e-19 $X=4.945 $Y=1.705
+ $X2=0 $Y2=0
cc_477 N_A_580_21#_c_544_n N_A_388_419#_c_1065_n 2.74426e-19 $X=5.35 $Y=0.18
+ $X2=0 $Y2=0
cc_478 N_A_580_21#_c_546_n N_A_388_419#_c_1065_n 7.4876e-19 $X=4.945 $Y=1.705
+ $X2=0 $Y2=0
cc_479 N_A_580_21#_c_549_n N_A_388_419#_c_1065_n 0.00433625f $X=5.645 $Y=1.45
+ $X2=0 $Y2=0
cc_480 N_A_580_21#_c_553_n N_A_388_419#_c_1065_n 0.00209528f $X=5.645 $Y=0.575
+ $X2=0 $Y2=0
cc_481 N_A_580_21#_M1019_g N_A_494_419#_c_1175_n 0.00382691f $X=3.41 $Y=2.595
+ $X2=0 $Y2=0
cc_482 N_A_580_21#_c_547_n N_A_494_419#_c_1175_n 0.00415929f $X=3.395 $Y=1.725
+ $X2=0 $Y2=0
cc_483 N_A_580_21#_M1019_g N_A_494_419#_c_1194_n 0.0129743f $X=3.41 $Y=2.595
+ $X2=0 $Y2=0
cc_484 N_A_580_21#_c_541_n N_A_494_419#_c_1176_n 0.00691538f $X=3.255 $Y=1.195
+ $X2=0 $Y2=0
cc_485 N_A_580_21#_c_542_n N_A_494_419#_c_1176_n 0.00593351f $X=3.05 $Y=1.195
+ $X2=0 $Y2=0
cc_486 N_A_580_21#_c_547_n N_A_494_419#_c_1176_n 0.00582176f $X=3.395 $Y=1.725
+ $X2=0 $Y2=0
cc_487 N_A_580_21#_M1019_g N_A_494_419#_c_1185_n 0.0216421f $X=3.41 $Y=2.595
+ $X2=0 $Y2=0
cc_488 N_A_580_21#_M1009_g N_A_494_419#_c_1178_n 0.0038831f $X=2.975 $Y=0.775
+ $X2=0 $Y2=0
cc_489 N_A_580_21#_c_541_n N_A_494_419#_c_1178_n 0.00986743f $X=3.255 $Y=1.195
+ $X2=0 $Y2=0
cc_490 N_A_580_21#_M1019_g N_A_494_419#_c_1204_n 0.00369099f $X=3.41 $Y=2.595
+ $X2=0 $Y2=0
cc_491 N_A_580_21#_c_555_n N_A_494_419#_c_1204_n 9.59622e-19 $X=4.82 $Y=2.08
+ $X2=0 $Y2=0
cc_492 N_A_580_21#_M1014_s N_A_494_419#_c_1186_n 0.00482786f $X=5.5 $Y=1.98
+ $X2=0 $Y2=0
cc_493 N_A_580_21#_c_555_n N_A_494_419#_c_1186_n 0.0169238f $X=4.82 $Y=2.08
+ $X2=0 $Y2=0
cc_494 N_A_580_21#_c_561_n N_A_494_419#_c_1186_n 0.0171499f $X=5.645 $Y=2.125
+ $X2=0 $Y2=0
cc_495 N_A_580_21#_M1019_g N_A_494_419#_c_1206_n 3.95188e-19 $X=3.41 $Y=2.595
+ $X2=0 $Y2=0
cc_496 N_A_580_21#_c_561_n N_A_494_419#_c_1230_n 0.0641776f $X=5.645 $Y=2.125
+ $X2=0 $Y2=0
cc_497 N_A_580_21#_c_549_n N_A_494_419#_c_1230_n 0.0088746f $X=5.645 $Y=1.45
+ $X2=0 $Y2=0
cc_498 N_A_580_21#_c_550_n N_A_494_419#_c_1230_n 3.2979e-19 $X=5.47 $Y=1.615
+ $X2=0 $Y2=0
cc_499 N_A_580_21#_c_551_n N_A_494_419#_c_1230_n 0.0243494f $X=5.645 $Y=1.615
+ $X2=0 $Y2=0
cc_500 N_A_580_21#_c_553_n N_A_494_419#_c_1179_n 0.00100885f $X=5.645 $Y=0.575
+ $X2=0 $Y2=0
cc_501 N_A_580_21#_c_549_n N_A_494_419#_c_1234_n 0.0126275f $X=5.645 $Y=1.45
+ $X2=0 $Y2=0
cc_502 N_A_580_21#_c_553_n N_A_494_419#_c_1234_n 0.0105021f $X=5.645 $Y=0.575
+ $X2=0 $Y2=0
cc_503 N_A_580_21#_c_543_n N_A_855_66#_c_1320_n 0.00839544f $X=4.2 $Y=0.255
+ $X2=0 $Y2=0
cc_504 N_A_580_21#_c_544_n N_A_855_66#_c_1320_n 0.00710251f $X=5.35 $Y=0.18
+ $X2=0 $Y2=0
cc_505 N_A_580_21#_c_552_n N_A_855_66#_c_1320_n 0.00213517f $X=5.515 $Y=0.43
+ $X2=0 $Y2=0
cc_506 N_A_580_21#_c_555_n N_A_855_66#_c_1322_n 0.0179471f $X=4.82 $Y=2.08 $X2=0
+ $Y2=0
cc_507 N_A_580_21#_c_546_n N_A_855_66#_c_1322_n 0.00300536f $X=4.945 $Y=1.705
+ $X2=0 $Y2=0
cc_508 N_A_580_21#_M1014_s N_A_855_66#_c_1329_n 0.00711734f $X=5.5 $Y=1.98 $X2=0
+ $Y2=0
cc_509 N_A_580_21#_c_555_n N_A_855_66#_c_1329_n 0.00890454f $X=4.82 $Y=2.08
+ $X2=0 $Y2=0
cc_510 N_A_580_21#_c_545_n N_A_855_66#_c_1329_n 0.00448991f $X=5.305 $Y=1.705
+ $X2=0 $Y2=0
cc_511 N_A_580_21#_c_561_n N_A_855_66#_c_1329_n 0.0157692f $X=5.645 $Y=2.125
+ $X2=0 $Y2=0
cc_512 N_A_580_21#_c_551_n N_A_855_66#_c_1329_n 0.00581477f $X=5.645 $Y=1.615
+ $X2=0 $Y2=0
cc_513 N_A_580_21#_c_553_n N_VGND_c_1450_n 0.0161365f $X=5.645 $Y=0.575 $X2=0
+ $Y2=0
cc_514 N_A_580_21#_c_540_n N_VGND_c_1452_n 0.0692241f $X=3.05 $Y=0.18 $X2=0
+ $Y2=0
cc_515 N_A_580_21#_c_553_n N_VGND_c_1452_n 0.0360686f $X=5.645 $Y=0.575 $X2=0
+ $Y2=0
cc_516 N_A_580_21#_c_539_n N_VGND_c_1458_n 0.0252586f $X=4.125 $Y=0.18 $X2=0
+ $Y2=0
cc_517 N_A_580_21#_c_540_n N_VGND_c_1458_n 0.00604685f $X=3.05 $Y=0.18 $X2=0
+ $Y2=0
cc_518 N_A_580_21#_c_544_n N_VGND_c_1458_n 0.0473659f $X=5.35 $Y=0.18 $X2=0
+ $Y2=0
cc_519 N_A_580_21#_c_548_n N_VGND_c_1458_n 0.00837817f $X=4.2 $Y=0.18 $X2=0
+ $Y2=0
cc_520 N_A_580_21#_c_553_n N_VGND_c_1458_n 0.0258529f $X=5.645 $Y=0.575 $X2=0
+ $Y2=0
cc_521 N_A_1393_300#_c_686_n N_C_c_770_n 6.39723e-19 $X=7.47 $Y=1.665 $X2=0
+ $Y2=0
cc_522 N_A_1393_300#_c_687_n N_C_c_770_n 0.0154798f $X=7.13 $Y=1.665 $X2=0 $Y2=0
cc_523 N_A_1393_300#_c_688_n N_C_c_770_n 0.0160826f $X=7.64 $Y=1.4 $X2=0 $Y2=0
cc_524 N_A_1393_300#_c_689_n N_C_c_770_n 0.00480316f $X=8.03 $Y=1.4 $X2=0 $Y2=0
cc_525 N_A_1393_300#_M1024_g N_C_c_779_n 0.0104115f $X=7.17 $Y=2.53 $X2=0 $Y2=0
cc_526 N_A_1393_300#_c_689_n N_C_c_780_n 0.0010383f $X=8.03 $Y=1.4 $X2=0 $Y2=0
cc_527 N_A_1393_300#_c_690_n N_C_c_780_n 0.0195723f $X=8.9 $Y=0.915 $X2=0 $Y2=0
cc_528 N_A_1393_300#_c_691_n N_C_c_780_n 0.0234569f $X=8.775 $Y=1.4 $X2=0 $Y2=0
cc_529 N_A_1393_300#_c_692_n N_C_c_780_n 0.0180925f $X=8.195 $Y=1.4 $X2=0 $Y2=0
cc_530 N_A_1393_300#_c_693_n N_C_c_780_n 0.00961025f $X=8.53 $Y=1.4 $X2=0 $Y2=0
cc_531 N_A_1393_300#_c_690_n N_C_c_781_n 0.0153642f $X=8.9 $Y=0.915 $X2=0 $Y2=0
cc_532 N_A_1393_300#_c_690_n N_C_c_771_n 0.0229455f $X=8.9 $Y=0.915 $X2=0 $Y2=0
cc_533 N_A_1393_300#_c_690_n N_C_c_772_n 3.61934e-19 $X=8.9 $Y=0.915 $X2=0 $Y2=0
cc_534 N_A_1393_300#_M1022_g N_C_c_774_n 0.00841328f $X=8.01 $Y=0.825 $X2=0
+ $Y2=0
cc_535 N_A_1393_300#_M1022_g N_C_c_775_n 0.0056288f $X=8.01 $Y=0.825 $X2=0 $Y2=0
cc_536 N_A_1393_300#_c_688_n N_C_c_775_n 0.00949705f $X=7.64 $Y=1.4 $X2=0 $Y2=0
cc_537 N_A_1393_300#_c_689_n N_C_c_775_n 4.5594e-19 $X=8.03 $Y=1.4 $X2=0 $Y2=0
cc_538 N_A_1393_300#_c_692_n N_C_c_775_n 0.0213489f $X=8.195 $Y=1.4 $X2=0 $Y2=0
cc_539 N_A_1393_300#_M1024_g N_C_c_783_n 0.0154798f $X=7.17 $Y=2.53 $X2=0 $Y2=0
cc_540 N_A_1393_300#_c_688_n N_C_c_783_n 0.00307765f $X=7.64 $Y=1.4 $X2=0 $Y2=0
cc_541 N_A_1393_300#_c_689_n N_C_c_783_n 0.00403946f $X=8.03 $Y=1.4 $X2=0 $Y2=0
cc_542 N_A_1393_300#_c_690_n N_C_c_784_n 0.00311796f $X=8.9 $Y=0.915 $X2=0 $Y2=0
cc_543 N_A_1393_300#_c_690_n C 0.0321122f $X=8.9 $Y=0.915 $X2=0 $Y2=0
cc_544 N_A_1393_300#_c_691_n C 7.09837e-19 $X=8.775 $Y=1.4 $X2=0 $Y2=0
cc_545 N_A_1393_300#_c_690_n N_C_c_777_n 0.00676586f $X=8.9 $Y=0.915 $X2=0 $Y2=0
cc_546 N_A_1393_300#_c_691_n N_C_c_777_n 0.014837f $X=8.775 $Y=1.4 $X2=0 $Y2=0
cc_547 N_A_1393_300#_M1024_g N_A_1459_406#_c_869_n 0.0151425f $X=7.17 $Y=2.53
+ $X2=0 $Y2=0
cc_548 N_A_1393_300#_c_686_n N_A_1459_406#_c_869_n 0.0160691f $X=7.47 $Y=1.665
+ $X2=0 $Y2=0
cc_549 N_A_1393_300#_c_688_n N_A_1459_406#_c_869_n 0.0104555f $X=7.64 $Y=1.4
+ $X2=0 $Y2=0
cc_550 N_A_1393_300#_M1026_s N_A_1459_406#_c_870_n 0.00564752f $X=8.755 $Y=2.065
+ $X2=0 $Y2=0
cc_551 N_A_1393_300#_c_690_n N_A_1459_406#_c_870_n 0.0248743f $X=8.9 $Y=0.915
+ $X2=0 $Y2=0
cc_552 N_A_1393_300#_M1024_g N_A_1459_406#_c_871_n 0.00411254f $X=7.17 $Y=2.53
+ $X2=0 $Y2=0
cc_553 N_A_1393_300#_M1022_g N_A_1459_406#_c_862_n 0.0132682f $X=8.01 $Y=0.825
+ $X2=0 $Y2=0
cc_554 N_A_1393_300#_c_688_n N_A_1459_406#_c_862_n 6.76284e-19 $X=7.64 $Y=1.4
+ $X2=0 $Y2=0
cc_555 N_A_1393_300#_c_689_n N_A_1459_406#_c_862_n 0.0265345f $X=8.03 $Y=1.4
+ $X2=0 $Y2=0
cc_556 N_A_1393_300#_c_692_n N_A_1459_406#_c_862_n 0.00162266f $X=8.195 $Y=1.4
+ $X2=0 $Y2=0
cc_557 N_A_1393_300#_M1022_g N_A_1459_406#_c_863_n 0.00589429f $X=8.01 $Y=0.825
+ $X2=0 $Y2=0
cc_558 N_A_1393_300#_c_690_n N_A_1459_406#_c_863_n 0.0229821f $X=8.9 $Y=0.915
+ $X2=0 $Y2=0
cc_559 N_A_1393_300#_c_690_n N_A_1459_406#_c_872_n 0.0553255f $X=8.9 $Y=0.915
+ $X2=0 $Y2=0
cc_560 N_A_1393_300#_c_690_n N_A_1459_406#_c_874_n 0.0136707f $X=8.9 $Y=0.915
+ $X2=0 $Y2=0
cc_561 N_A_1393_300#_M1024_g N_VPWR_c_972_n 0.00287879f $X=7.17 $Y=2.53 $X2=0
+ $Y2=0
cc_562 N_A_1393_300#_M1024_g N_VPWR_c_978_n 0.00803988f $X=7.17 $Y=2.53 $X2=0
+ $Y2=0
cc_563 N_A_1393_300#_M1024_g N_VPWR_c_970_n 0.0154548f $X=7.17 $Y=2.53 $X2=0
+ $Y2=0
cc_564 N_A_1393_300#_M1024_g N_A_494_419#_c_1187_n 0.0135444f $X=7.17 $Y=2.53
+ $X2=0 $Y2=0
cc_565 N_A_1393_300#_c_686_n N_A_494_419#_c_1180_n 0.0111221f $X=7.47 $Y=1.665
+ $X2=0 $Y2=0
cc_566 N_A_1393_300#_c_687_n N_A_494_419#_c_1180_n 0.00374292f $X=7.13 $Y=1.665
+ $X2=0 $Y2=0
cc_567 N_A_1393_300#_M1024_g N_A_494_419#_c_1189_n 0.00462278f $X=7.17 $Y=2.53
+ $X2=0 $Y2=0
cc_568 N_A_1393_300#_c_686_n N_A_494_419#_c_1189_n 0.00799475f $X=7.47 $Y=1.665
+ $X2=0 $Y2=0
cc_569 N_A_1393_300#_c_687_n N_A_494_419#_c_1189_n 0.00185447f $X=7.13 $Y=1.665
+ $X2=0 $Y2=0
cc_570 N_A_1393_300#_M1024_g N_A_494_419#_c_1182_n 0.00590404f $X=7.17 $Y=2.53
+ $X2=0 $Y2=0
cc_571 N_A_1393_300#_c_686_n N_A_494_419#_c_1182_n 0.0245129f $X=7.47 $Y=1.665
+ $X2=0 $Y2=0
cc_572 N_A_1393_300#_c_687_n N_A_494_419#_c_1182_n 0.00228363f $X=7.13 $Y=1.665
+ $X2=0 $Y2=0
cc_573 N_A_1393_300#_c_686_n N_A_494_419#_c_1183_n 0.0207542f $X=7.47 $Y=1.665
+ $X2=0 $Y2=0
cc_574 N_A_1393_300#_c_687_n N_A_494_419#_c_1183_n 0.00471432f $X=7.13 $Y=1.665
+ $X2=0 $Y2=0
cc_575 N_A_1393_300#_c_688_n N_A_494_419#_c_1183_n 0.00689247f $X=7.64 $Y=1.4
+ $X2=0 $Y2=0
cc_576 N_A_1393_300#_M1024_g N_A_855_66#_c_1323_n 2.69749e-19 $X=7.17 $Y=2.53
+ $X2=0 $Y2=0
cc_577 N_A_1393_300#_M1022_g N_A_855_66#_c_1323_n 0.00574556f $X=8.01 $Y=0.825
+ $X2=0 $Y2=0
cc_578 N_A_1393_300#_c_688_n N_A_855_66#_c_1323_n 0.00658057f $X=7.64 $Y=1.4
+ $X2=0 $Y2=0
cc_579 N_A_1393_300#_c_689_n N_A_855_66#_c_1323_n 0.0378297f $X=8.03 $Y=1.4
+ $X2=0 $Y2=0
cc_580 N_A_1393_300#_c_690_n N_A_855_66#_c_1323_n 0.0600463f $X=8.9 $Y=0.915
+ $X2=0 $Y2=0
cc_581 N_A_1393_300#_c_691_n N_A_855_66#_c_1323_n 0.00167515f $X=8.775 $Y=1.4
+ $X2=0 $Y2=0
cc_582 N_A_1393_300#_c_692_n N_A_855_66#_c_1323_n 0.00236261f $X=8.195 $Y=1.4
+ $X2=0 $Y2=0
cc_583 N_A_1393_300#_c_693_n N_A_855_66#_c_1323_n 0.0130557f $X=8.53 $Y=1.4
+ $X2=0 $Y2=0
cc_584 N_A_1393_300#_M1022_g N_A_855_66#_c_1326_n 0.00849368f $X=8.01 $Y=0.825
+ $X2=0 $Y2=0
cc_585 N_A_1393_300#_c_690_n N_A_855_66#_c_1326_n 0.100761f $X=8.9 $Y=0.915
+ $X2=0 $Y2=0
cc_586 N_A_1393_300#_c_692_n N_A_855_66#_c_1326_n 0.0067948f $X=8.195 $Y=1.4
+ $X2=0 $Y2=0
cc_587 N_A_1393_300#_M1024_g N_A_855_66#_c_1329_n 0.0110101f $X=7.17 $Y=2.53
+ $X2=0 $Y2=0
cc_588 N_A_1393_300#_c_686_n N_A_855_66#_c_1329_n 0.00691814f $X=7.47 $Y=1.665
+ $X2=0 $Y2=0
cc_589 N_A_1393_300#_c_688_n N_A_855_66#_c_1329_n 0.00174396f $X=7.64 $Y=1.4
+ $X2=0 $Y2=0
cc_590 N_A_1393_300#_c_690_n N_A_855_66#_c_1380_n 8.11873e-19 $X=8.9 $Y=0.915
+ $X2=0 $Y2=0
cc_591 N_A_1393_300#_M1022_g N_VGND_c_1454_n 2.33881e-19 $X=8.01 $Y=0.825 $X2=0
+ $Y2=0
cc_592 N_C_c_781_n N_A_1459_406#_M1021_g 0.0119202f $X=9.165 $Y=1.955 $X2=0
+ $Y2=0
cc_593 N_C_c_784_n N_A_1459_406#_M1021_g 0.00603868f $X=9.405 $Y=1.88 $X2=0
+ $Y2=0
cc_594 N_C_c_773_n N_A_1459_406#_M1011_g 0.0126622f $X=9.585 $Y=1.235 $X2=0
+ $Y2=0
cc_595 C N_A_1459_406#_M1011_g 0.00164264f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_596 N_C_c_779_n N_A_1459_406#_c_869_n 0.0199211f $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_597 N_C_c_783_n N_A_1459_406#_c_869_n 0.00220314f $X=7.665 $Y=1.88 $X2=0
+ $Y2=0
cc_598 N_C_c_779_n N_A_1459_406#_c_870_n 0.0137158f $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_599 N_C_c_781_n N_A_1459_406#_c_870_n 0.0205357f $X=9.165 $Y=1.955 $X2=0
+ $Y2=0
cc_600 N_C_c_779_n N_A_1459_406#_c_871_n 9.73778e-19 $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_601 N_C_c_774_n N_A_1459_406#_c_862_n 0.00372443f $X=7.565 $Y=1.11 $X2=0
+ $Y2=0
cc_602 N_C_c_775_n N_A_1459_406#_c_862_n 7.79053e-19 $X=7.565 $Y=1.26 $X2=0
+ $Y2=0
cc_603 N_C_c_771_n N_A_1459_406#_c_863_n 0.00643157f $X=9.225 $Y=1.235 $X2=0
+ $Y2=0
cc_604 N_C_c_773_n N_A_1459_406#_c_863_n 0.00643157f $X=9.585 $Y=1.235 $X2=0
+ $Y2=0
cc_605 N_C_c_781_n N_A_1459_406#_c_872_n 0.0331964f $X=9.165 $Y=1.955 $X2=0
+ $Y2=0
cc_606 N_C_c_784_n N_A_1459_406#_c_872_n 0.00489502f $X=9.405 $Y=1.88 $X2=0
+ $Y2=0
cc_607 N_C_c_772_n N_A_1459_406#_c_873_n 0.00216834f $X=9.405 $Y=1.805 $X2=0
+ $Y2=0
cc_608 N_C_c_784_n N_A_1459_406#_c_873_n 0.00479098f $X=9.405 $Y=1.88 $X2=0
+ $Y2=0
cc_609 C N_A_1459_406#_c_873_n 0.0398713f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_610 N_C_c_777_n N_A_1459_406#_c_873_n 0.00471135f $X=9.495 $Y=1.4 $X2=0 $Y2=0
cc_611 N_C_c_772_n N_A_1459_406#_c_874_n 0.00267888f $X=9.405 $Y=1.805 $X2=0
+ $Y2=0
cc_612 N_C_c_784_n N_A_1459_406#_c_874_n 0.00340342f $X=9.405 $Y=1.88 $X2=0
+ $Y2=0
cc_613 C N_A_1459_406#_c_874_n 0.013853f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_614 N_C_c_777_n N_A_1459_406#_c_874_n 4.38616e-19 $X=9.495 $Y=1.4 $X2=0 $Y2=0
cc_615 N_C_c_772_n N_A_1459_406#_c_865_n 6.84637e-19 $X=9.405 $Y=1.805 $X2=0
+ $Y2=0
cc_616 C N_A_1459_406#_c_865_n 0.0251661f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_617 N_C_c_772_n N_A_1459_406#_c_866_n 0.00603868f $X=9.405 $Y=1.805 $X2=0
+ $Y2=0
cc_618 C N_A_1459_406#_c_866_n 0.0114453f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_619 N_C_c_777_n N_A_1459_406#_c_866_n 0.0182439f $X=9.495 $Y=1.4 $X2=0 $Y2=0
cc_620 N_C_c_773_n N_A_1459_406#_c_867_n 0.00129382f $X=9.585 $Y=1.235 $X2=0
+ $Y2=0
cc_621 N_C_c_781_n N_VPWR_c_973_n 0.00532643f $X=9.165 $Y=1.955 $X2=0 $Y2=0
cc_622 N_C_c_779_n N_VPWR_c_978_n 0.00531075f $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_623 N_C_c_781_n N_VPWR_c_978_n 0.00567004f $X=9.165 $Y=1.955 $X2=0 $Y2=0
cc_624 N_C_c_779_n N_VPWR_c_970_n 0.0080075f $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_625 N_C_c_781_n N_VPWR_c_970_n 0.00924973f $X=9.165 $Y=1.955 $X2=0 $Y2=0
cc_626 N_C_c_779_n N_A_494_419#_c_1189_n 3.26157e-19 $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_627 N_C_c_770_n N_A_494_419#_c_1183_n 4.31446e-19 $X=7.58 $Y=1.805 $X2=0
+ $Y2=0
cc_628 N_C_c_774_n N_A_494_419#_c_1183_n 0.00824332f $X=7.565 $Y=1.11 $X2=0
+ $Y2=0
cc_629 N_C_c_770_n N_A_855_66#_c_1323_n 0.00319617f $X=7.58 $Y=1.805 $X2=0 $Y2=0
cc_630 N_C_c_779_n N_A_855_66#_c_1323_n 0.0133438f $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_631 N_C_c_780_n N_A_855_66#_c_1323_n 0.0320204f $X=9.04 $Y=1.88 $X2=0 $Y2=0
cc_632 N_C_c_781_n N_A_855_66#_c_1323_n 0.00121965f $X=9.165 $Y=1.955 $X2=0
+ $Y2=0
cc_633 N_C_c_771_n N_A_855_66#_c_1326_n 0.00215563f $X=9.225 $Y=1.235 $X2=0
+ $Y2=0
cc_634 N_C_c_779_n N_A_855_66#_c_1329_n 0.00808014f $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_635 N_C_c_779_n N_A_855_66#_c_1380_n 0.00202215f $X=7.7 $Y=1.955 $X2=0 $Y2=0
cc_636 N_C_c_774_n N_VGND_c_1450_n 0.00311193f $X=7.565 $Y=1.11 $X2=0 $Y2=0
cc_637 N_C_c_773_n N_VGND_c_1496_n 0.00690783f $X=9.585 $Y=1.235 $X2=0 $Y2=0
cc_638 C N_VGND_c_1496_n 0.0139019f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_639 N_C_c_774_n N_VGND_c_1454_n 0.00420632f $X=7.565 $Y=1.11 $X2=0 $Y2=0
cc_640 N_C_c_774_n N_VGND_c_1458_n 0.00472204f $X=7.565 $Y=1.11 $X2=0 $Y2=0
cc_641 N_A_1459_406#_c_870_n N_VPWR_M1026_d 0.00238559f $X=9.245 $Y=2.98 $X2=0
+ $Y2=0
cc_642 N_A_1459_406#_c_872_n N_VPWR_M1026_d 0.00815676f $X=9.33 $Y=2.895 $X2=0
+ $Y2=0
cc_643 N_A_1459_406#_M1021_g N_VPWR_c_973_n 0.0276073f $X=10.025 $Y=2.565 $X2=0
+ $Y2=0
cc_644 N_A_1459_406#_c_870_n N_VPWR_c_973_n 0.0138718f $X=9.245 $Y=2.98 $X2=0
+ $Y2=0
cc_645 N_A_1459_406#_c_872_n N_VPWR_c_973_n 0.0585588f $X=9.33 $Y=2.895 $X2=0
+ $Y2=0
cc_646 N_A_1459_406#_c_873_n N_VPWR_c_973_n 0.0233644f $X=10.135 $Y=1.83 $X2=0
+ $Y2=0
cc_647 N_A_1459_406#_c_870_n N_VPWR_c_978_n 0.105922f $X=9.245 $Y=2.98 $X2=0
+ $Y2=0
cc_648 N_A_1459_406#_c_871_n N_VPWR_c_978_n 0.022043f $X=7.6 $Y=2.98 $X2=0 $Y2=0
cc_649 N_A_1459_406#_M1021_g N_VPWR_c_979_n 0.0079675f $X=10.025 $Y=2.565 $X2=0
+ $Y2=0
cc_650 N_A_1459_406#_M1021_g N_VPWR_c_970_n 0.0146353f $X=10.025 $Y=2.565 $X2=0
+ $Y2=0
cc_651 N_A_1459_406#_c_870_n N_VPWR_c_970_n 0.0658688f $X=9.245 $Y=2.98 $X2=0
+ $Y2=0
cc_652 N_A_1459_406#_c_871_n N_VPWR_c_970_n 0.012533f $X=7.6 $Y=2.98 $X2=0 $Y2=0
cc_653 N_A_1459_406#_c_871_n N_A_494_419#_c_1187_n 0.0111138f $X=7.6 $Y=2.98
+ $X2=0 $Y2=0
cc_654 N_A_1459_406#_c_869_n N_A_494_419#_c_1189_n 0.0578954f $X=7.435 $Y=2.175
+ $X2=0 $Y2=0
cc_655 N_A_1459_406#_c_862_n N_A_494_419#_c_1183_n 0.00305012f $X=7.795 $Y=0.825
+ $X2=0 $Y2=0
cc_656 N_A_1459_406#_c_870_n N_A_855_66#_M1012_d 0.00318153f $X=9.245 $Y=2.98
+ $X2=0 $Y2=0
cc_657 N_A_1459_406#_c_869_n N_A_855_66#_c_1323_n 0.0455877f $X=7.435 $Y=2.175
+ $X2=0 $Y2=0
cc_658 N_A_1459_406#_c_870_n N_A_855_66#_c_1323_n 0.0455332f $X=9.245 $Y=2.98
+ $X2=0 $Y2=0
cc_659 N_A_1459_406#_c_862_n N_A_855_66#_c_1326_n 0.0165345f $X=7.795 $Y=0.825
+ $X2=0 $Y2=0
cc_660 N_A_1459_406#_c_863_n N_A_855_66#_c_1326_n 0.0249842f $X=9.87 $Y=0.35
+ $X2=0 $Y2=0
cc_661 N_A_1459_406#_c_869_n N_A_855_66#_c_1329_n 0.0314235f $X=7.435 $Y=2.175
+ $X2=0 $Y2=0
cc_662 N_A_1459_406#_c_870_n N_A_855_66#_c_1329_n 0.00497991f $X=9.245 $Y=2.98
+ $X2=0 $Y2=0
cc_663 N_A_1459_406#_c_869_n N_A_855_66#_c_1380_n 0.00224349f $X=7.435 $Y=2.175
+ $X2=0 $Y2=0
cc_664 N_A_1459_406#_c_870_n N_A_855_66#_c_1380_n 0.00207384f $X=9.245 $Y=2.98
+ $X2=0 $Y2=0
cc_665 N_A_1459_406#_c_873_n N_X_c_1426_n 7.74607e-19 $X=10.135 $Y=1.83 $X2=0
+ $Y2=0
cc_666 N_A_1459_406#_M1021_g N_X_c_1427_n 0.0226737f $X=10.025 $Y=2.565 $X2=0
+ $Y2=0
cc_667 N_A_1459_406#_c_873_n N_X_c_1427_n 0.0263289f $X=10.135 $Y=1.83 $X2=0
+ $Y2=0
cc_668 N_A_1459_406#_c_866_n N_X_c_1427_n 0.00212986f $X=10.3 $Y=1.4 $X2=0 $Y2=0
cc_669 N_A_1459_406#_M1021_g X 0.00154119f $X=10.025 $Y=2.565 $X2=0 $Y2=0
cc_670 N_A_1459_406#_M1021_g N_X_c_1425_n 0.00433944f $X=10.025 $Y=2.565 $X2=0
+ $Y2=0
cc_671 N_A_1459_406#_c_861_n N_X_c_1425_n 0.0101094f $X=10.545 $Y=1.235 $X2=0
+ $Y2=0
cc_672 N_A_1459_406#_c_873_n N_X_c_1425_n 0.0119574f $X=10.135 $Y=1.83 $X2=0
+ $Y2=0
cc_673 N_A_1459_406#_c_865_n N_X_c_1425_n 0.0336737f $X=10.3 $Y=1.4 $X2=0 $Y2=0
cc_674 N_A_1459_406#_c_866_n N_X_c_1425_n 0.00995914f $X=10.3 $Y=1.4 $X2=0 $Y2=0
cc_675 N_A_1459_406#_M1011_g N_VGND_c_1496_n 0.0123037f $X=10.155 $Y=0.915 $X2=0
+ $Y2=0
cc_676 N_A_1459_406#_c_861_n N_VGND_c_1496_n 0.00588592f $X=10.545 $Y=1.235
+ $X2=0 $Y2=0
cc_677 N_A_1459_406#_c_863_n N_VGND_c_1496_n 0.0207938f $X=9.87 $Y=0.35 $X2=0
+ $Y2=0
cc_678 N_A_1459_406#_c_865_n N_VGND_c_1496_n 0.0174319f $X=10.3 $Y=1.4 $X2=0
+ $Y2=0
cc_679 N_A_1459_406#_c_866_n N_VGND_c_1496_n 0.00287738f $X=10.3 $Y=1.4 $X2=0
+ $Y2=0
cc_680 N_A_1459_406#_c_867_n N_VGND_c_1496_n 8.34782e-19 $X=10.155 $Y=0.43 $X2=0
+ $Y2=0
cc_681 N_A_1459_406#_c_861_n N_VGND_c_1451_n 0.00723923f $X=10.545 $Y=1.235
+ $X2=0 $Y2=0
cc_682 N_A_1459_406#_c_863_n N_VGND_c_1451_n 0.0234275f $X=9.87 $Y=0.35 $X2=0
+ $Y2=0
cc_683 N_A_1459_406#_c_867_n N_VGND_c_1451_n 0.0118826f $X=10.155 $Y=0.43 $X2=0
+ $Y2=0
cc_684 N_A_1459_406#_c_863_n N_VGND_c_1454_n 0.13238f $X=9.87 $Y=0.35 $X2=0
+ $Y2=0
cc_685 N_A_1459_406#_c_864_n N_VGND_c_1454_n 0.0222501f $X=7.96 $Y=0.35 $X2=0
+ $Y2=0
cc_686 N_A_1459_406#_c_867_n N_VGND_c_1454_n 0.00496932f $X=10.155 $Y=0.43 $X2=0
+ $Y2=0
cc_687 N_A_1459_406#_c_861_n N_VGND_c_1457_n 0.0031218f $X=10.545 $Y=1.235 $X2=0
+ $Y2=0
cc_688 N_A_1459_406#_c_861_n N_VGND_c_1458_n 0.00376215f $X=10.545 $Y=1.235
+ $X2=0 $Y2=0
cc_689 N_A_1459_406#_c_863_n N_VGND_c_1458_n 0.0815813f $X=9.87 $Y=0.35 $X2=0
+ $Y2=0
cc_690 N_A_1459_406#_c_864_n N_VGND_c_1458_n 0.0127687f $X=7.96 $Y=0.35 $X2=0
+ $Y2=0
cc_691 N_A_1459_406#_c_867_n N_VGND_c_1458_n 0.00311548f $X=10.155 $Y=0.43 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_970_n N_A_388_419#_M1003_d 0.00225465f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_970_n N_A_388_419#_M1007_d 0.00233022f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_970_n N_A_494_419#_M1017_d 0.00671563f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_972_n N_A_494_419#_c_1186_n 0.0128931f $X=6.345 $Y=2.125 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_976_n N_A_494_419#_c_1186_n 0.108574f $X=6.26 $Y=3.33 $X2=0
+ $Y2=0
cc_697 N_VPWR_c_970_n N_A_494_419#_c_1186_n 0.0677768f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_698 N_VPWR_c_976_n N_A_494_419#_c_1206_n 0.0093013f $X=6.26 $Y=3.33 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_970_n N_A_494_419#_c_1206_n 0.00641662f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_700 N_VPWR_c_972_n N_A_494_419#_c_1230_n 0.0622048f $X=6.345 $Y=2.125 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_972_n N_A_494_419#_c_1179_n 0.00561498f $X=6.345 $Y=2.125 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_978_n N_A_494_419#_c_1187_n 0.0279532f $X=9.595 $Y=3.33 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_970_n N_A_494_419#_c_1187_n 0.0172861f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_972_n N_A_494_419#_c_1182_n 0.0803807f $X=6.345 $Y=2.125 $X2=0
+ $Y2=0
cc_705 N_VPWR_c_970_n N_A_855_66#_M1020_d 0.00233518f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_706 N_VPWR_M1014_d N_A_855_66#_c_1329_n 0.0149858f $X=6.125 $Y=1.98 $X2=0
+ $Y2=0
cc_707 N_VPWR_c_972_n N_A_855_66#_c_1329_n 0.022485f $X=6.345 $Y=2.125 $X2=0
+ $Y2=0
cc_708 N_VPWR_c_973_n N_X_c_1427_n 0.0645857f $X=9.76 $Y=2.26 $X2=0 $Y2=0
cc_709 N_VPWR_c_979_n N_X_c_1427_n 0.019758f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_710 N_VPWR_c_970_n N_X_c_1427_n 0.0125705f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_711 N_VPWR_c_979_n X 0.00810947f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_712 N_VPWR_c_970_n X 0.00864691f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_713 N_A_388_419#_c_1063_n N_A_494_419#_M1009_d 0.00481641f $X=4.895 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_714 N_A_388_419#_c_1058_n N_A_494_419#_c_1175_n 0.0506443f $X=2.08 $Y=2.395
+ $X2=0 $Y2=0
cc_715 N_A_388_419#_c_1058_n N_A_494_419#_c_1194_n 0.0338071f $X=2.08 $Y=2.395
+ $X2=0 $Y2=0
cc_716 N_A_388_419#_c_1061_n N_A_494_419#_c_1176_n 0.0174439f $X=2.68 $Y=0.775
+ $X2=0 $Y2=0
cc_717 N_A_388_419#_c_1063_n N_A_494_419#_c_1176_n 0.0121353f $X=4.895 $Y=0.925
+ $X2=0 $Y2=0
cc_718 N_A_388_419#_c_1058_n N_A_494_419#_c_1177_n 0.0139178f $X=2.08 $Y=2.395
+ $X2=0 $Y2=0
cc_719 N_A_388_419#_c_1059_n N_A_494_419#_c_1177_n 0.00589195f $X=2.515 $Y=0.907
+ $X2=0 $Y2=0
cc_720 N_A_388_419#_c_1061_n N_A_494_419#_c_1177_n 0.00592132f $X=2.68 $Y=0.775
+ $X2=0 $Y2=0
cc_721 N_A_388_419#_c_1063_n N_A_494_419#_c_1177_n 0.00136924f $X=4.895 $Y=0.925
+ $X2=0 $Y2=0
cc_722 N_A_388_419#_c_1061_n N_A_494_419#_c_1178_n 0.00415811f $X=2.68 $Y=0.775
+ $X2=0 $Y2=0
cc_723 N_A_388_419#_c_1063_n N_A_494_419#_c_1178_n 0.022761f $X=4.895 $Y=0.925
+ $X2=0 $Y2=0
cc_724 N_A_388_419#_M1007_d N_A_494_419#_c_1186_n 0.00556169f $X=4.945 $Y=2.095
+ $X2=0 $Y2=0
cc_725 N_A_388_419#_c_1067_n N_A_494_419#_c_1186_n 0.017081f $X=5.085 $Y=2.395
+ $X2=0 $Y2=0
cc_726 N_A_388_419#_c_1058_n N_A_494_419#_c_1188_n 0.0129587f $X=2.08 $Y=2.395
+ $X2=0 $Y2=0
cc_727 N_A_388_419#_c_1063_n N_A_855_66#_M1018_d 0.00142845f $X=4.895 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_728 N_A_388_419#_c_1060_n N_A_855_66#_c_1320_n 0.0196097f $X=5.04 $Y=1.04
+ $X2=0 $Y2=0
cc_729 N_A_388_419#_c_1063_n N_A_855_66#_c_1320_n 0.0108627f $X=4.895 $Y=0.925
+ $X2=0 $Y2=0
cc_730 N_A_388_419#_c_1065_n N_A_855_66#_c_1320_n 3.08449e-19 $X=5.04 $Y=0.925
+ $X2=0 $Y2=0
cc_731 N_A_388_419#_c_1062_n N_A_855_66#_c_1321_n 0.00569024f $X=5.102 $Y=1.96
+ $X2=0 $Y2=0
cc_732 N_A_388_419#_c_1067_n N_A_855_66#_c_1322_n 0.0164068f $X=5.085 $Y=2.395
+ $X2=0 $Y2=0
cc_733 N_A_388_419#_c_1062_n N_A_855_66#_c_1322_n 0.0575109f $X=5.102 $Y=1.96
+ $X2=0 $Y2=0
cc_734 N_A_388_419#_c_1063_n N_A_855_66#_c_1324_n 0.0140429f $X=4.895 $Y=0.925
+ $X2=0 $Y2=0
cc_735 N_A_388_419#_c_1065_n N_A_855_66#_c_1324_n 2.74177e-19 $X=5.04 $Y=0.925
+ $X2=0 $Y2=0
cc_736 N_A_388_419#_c_1062_n N_A_855_66#_c_1325_n 0.0129661f $X=5.102 $Y=1.96
+ $X2=0 $Y2=0
cc_737 N_A_388_419#_c_1063_n N_A_855_66#_c_1325_n 0.00605049f $X=4.895 $Y=0.925
+ $X2=0 $Y2=0
cc_738 N_A_388_419#_M1007_d N_A_855_66#_c_1329_n 2.28076e-19 $X=4.945 $Y=2.095
+ $X2=0 $Y2=0
cc_739 N_A_388_419#_c_1067_n N_A_855_66#_c_1329_n 0.0205661f $X=5.085 $Y=2.395
+ $X2=0 $Y2=0
cc_740 N_A_388_419#_c_1067_n N_A_855_66#_c_1353_n 5.83106e-19 $X=5.085 $Y=2.395
+ $X2=0 $Y2=0
cc_741 N_A_388_419#_c_1071_n N_VGND_M1025_d 0.00241065f $X=2.08 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_742 N_A_388_419#_c_1060_n N_VGND_c_1452_n 0.00743721f $X=5.04 $Y=1.04 $X2=0
+ $Y2=0
cc_743 N_A_388_419#_c_1060_n N_VGND_c_1458_n 0.00904202f $X=5.04 $Y=1.04 $X2=0
+ $Y2=0
cc_744 N_A_388_419#_c_1071_n A_430_113# 3.56716e-19 $X=2.08 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_745 N_A_388_419#_c_1059_n A_430_113# 9.76475e-19 $X=2.515 $Y=0.907 $X2=-0.19
+ $Y2=-0.245
cc_746 N_A_388_419#_c_1064_n A_430_113# 0.00104121f $X=2.305 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_747 N_A_494_419#_c_1186_n N_A_855_66#_M1020_d 0.00352795f $X=5.91 $Y=2.98
+ $X2=0 $Y2=0
cc_748 N_A_494_419#_c_1185_n N_A_855_66#_c_1322_n 0.00670537f $X=4.02 $Y=2.16
+ $X2=0 $Y2=0
cc_749 N_A_494_419#_c_1204_n N_A_855_66#_c_1322_n 0.0263441f $X=4.105 $Y=2.895
+ $X2=0 $Y2=0
cc_750 N_A_494_419#_c_1186_n N_A_855_66#_c_1322_n 0.0172821f $X=5.91 $Y=2.98
+ $X2=0 $Y2=0
cc_751 N_A_494_419#_c_1186_n N_A_855_66#_c_1329_n 0.0224095f $X=5.91 $Y=2.98
+ $X2=0 $Y2=0
cc_752 N_A_494_419#_c_1230_n N_A_855_66#_c_1329_n 0.0233148f $X=5.995 $Y=2.895
+ $X2=0 $Y2=0
cc_753 N_A_494_419#_c_1187_n N_A_855_66#_c_1329_n 0.0537586f $X=6.905 $Y=2.885
+ $X2=0 $Y2=0
cc_754 N_A_494_419#_c_1204_n N_A_855_66#_c_1353_n 0.00188527f $X=4.105 $Y=2.895
+ $X2=0 $Y2=0
cc_755 N_A_494_419#_c_1186_n N_A_855_66#_c_1353_n 0.00140769f $X=5.91 $Y=2.98
+ $X2=0 $Y2=0
cc_756 N_A_494_419#_c_1179_n N_VGND_c_1450_n 0.00311024f $X=6.615 $Y=1.235 $X2=0
+ $Y2=0
cc_757 N_A_494_419#_c_1180_n N_VGND_c_1450_n 0.00641281f $X=7.12 $Y=1.235 $X2=0
+ $Y2=0
cc_758 N_A_494_419#_c_1181_n N_VGND_c_1450_n 0.0116607f $X=6.7 $Y=1.235 $X2=0
+ $Y2=0
cc_759 N_A_494_419#_c_1183_n N_VGND_c_1450_n 0.0196195f $X=7.285 $Y=0.825 $X2=0
+ $Y2=0
cc_760 N_A_494_419#_c_1183_n N_VGND_c_1454_n 0.00717615f $X=7.285 $Y=0.825 $X2=0
+ $Y2=0
cc_761 N_A_494_419#_c_1183_n N_VGND_c_1458_n 0.0102262f $X=7.285 $Y=0.825 $X2=0
+ $Y2=0
cc_762 N_A_855_66#_c_1320_n N_VGND_c_1452_n 0.0174108f $X=4.495 $Y=0.475 $X2=0
+ $Y2=0
cc_763 N_A_855_66#_c_1320_n N_VGND_c_1458_n 0.0110845f $X=4.495 $Y=0.475 $X2=0
+ $Y2=0
cc_764 N_X_c_1425_n N_VGND_c_1451_n 0.00360907f $X=10.76 $Y=0.915 $X2=0 $Y2=0
cc_765 N_X_c_1425_n N_VGND_c_1457_n 0.00454326f $X=10.76 $Y=0.915 $X2=0 $Y2=0
cc_766 N_X_c_1425_n N_VGND_c_1458_n 0.00725286f $X=10.76 $Y=0.915 $X2=0 $Y2=0
cc_767 N_VGND_c_1496_n A_2046_141# 0.00210431f $X=10.325 $Y=0.887 $X2=-0.19
+ $Y2=-0.245
cc_768 N_VGND_c_1451_n A_2046_141# 7.68185e-19 $X=10.41 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
