* File: sky130_fd_sc_lp__a211o_1.pex.spice
* Created: Wed Sep  2 09:17:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211O_1%A_80_237# 1 2 3 12 14 16 20 21 22 23 24 25
+ 28 30 34 40 43
c87 12 0 1.27104e-19 $X=0.475 $Y=2.465
r88 44 46 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.475 $Y=1.35
+ $X2=0.515 $Y2=1.35
r89 38 40 16.7104 $w=2.98e-07 $l=4.35e-07 $layer=LI1_cond $X=3.095 $Y=0.855
+ $X2=3.095 $Y2=0.42
r90 34 36 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=3.08 $Y=1.98
+ $X2=3.08 $Y2=2.91
r91 32 34 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.08 $Y=1.865
+ $X2=3.08 $Y2=1.98
r92 31 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0.94
+ $X2=2.07 $Y2=0.94
r93 30 38 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.945 $Y=0.94
+ $X2=3.095 $Y2=0.855
r94 30 31 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.945 $Y=0.94
+ $X2=2.235 $Y2=0.94
r95 26 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.855
+ $X2=2.07 $Y2=0.94
r96 26 28 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.07 $Y=0.855
+ $X2=2.07 $Y2=0.375
r97 24 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.915 $Y=1.78
+ $X2=3.08 $Y2=1.865
r98 24 25 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=2.915 $Y=1.78
+ $X2=0.915 $Y2=1.78
r99 22 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0.94
+ $X2=2.07 $Y2=0.94
r100 22 23 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.905 $Y=0.94
+ $X2=0.915 $Y2=0.94
r101 21 46 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.75 $Y=1.35
+ $X2=0.515 $Y2=1.35
r102 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.35 $X2=0.75 $Y2=1.35
r103 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.75 $Y=1.695
+ $X2=0.915 $Y2=1.78
r104 18 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.75 $Y=1.695
+ $X2=0.75 $Y2=1.35
r105 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.75 $Y=1.025
+ $X2=0.915 $Y2=0.94
r106 17 20 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.75 $Y=1.025
+ $X2=0.75 $Y2=1.35
r107 14 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.185
+ $X2=0.515 $Y2=1.35
r108 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.515 $Y=1.185
+ $X2=0.515 $Y2=0.655
r109 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=1.35
r110 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=2.465
r111 3 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=2.91
r112 3 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=1.98
r113 2 40 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.42
r114 1 43 182 $w=1.7e-07 $l=8.03166e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=2.07 $Y2=0.94
r115 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=2.07 $Y2=0.375
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%A2 1 3 4 6 8 12
c32 12 0 6.00056e-21 $X=1.305 $Y=1.36
c33 4 0 1.27104e-19 $X=1.425 $Y=1.525
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.305
+ $Y=1.36 $X2=1.305 $Y2=1.36
r35 8 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.36
+ $X2=1.305 $Y2=1.36
r36 4 11 38.7084 $w=3.43e-07 $l=2.11069e-07 $layer=POLY_cond $X=1.425 $Y=1.525
+ $X2=1.32 $Y2=1.36
r37 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.425 $Y=1.525 $X2=1.425
+ $Y2=2.465
r38 1 11 38.7084 $w=3.43e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.395 $Y=1.195
+ $X2=1.32 $Y2=1.36
r39 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.395 $Y=1.195
+ $X2=1.395 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%A1 3 6 8 11 12 13
c31 12 0 2.79301e-20 $X=1.875 $Y=1.35
c32 6 0 3.99686e-20 $X=1.935 $Y=2.465
r33 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.35
+ $X2=1.875 $Y2=1.515
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.35
+ $X2=1.875 $Y2=1.185
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.875
+ $Y=1.35 $X2=1.875 $Y2=1.35
r36 8 12 7.13417 $w=3.13e-07 $l=1.95e-07 $layer=LI1_cond $X=1.68 $Y=1.367
+ $X2=1.875 $Y2=1.367
r37 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.935 $Y=2.465
+ $X2=1.935 $Y2=1.515
r38 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.785 $Y=0.655
+ $X2=1.785 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%B1 3 6 8 11 13
c29 8 0 3.3968e-20 $X=2.64 $Y=1.295
c30 6 0 3.40175e-20 $X=2.445 $Y=2.465
r31 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.515
r32 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.185
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.35 $X2=2.415 $Y2=1.35
r34 8 12 8.23174 $w=3.13e-07 $l=2.25e-07 $layer=LI1_cond $X=2.64 $Y=1.367
+ $X2=2.415 $Y2=1.367
r35 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.445 $Y=2.465
+ $X2=2.445 $Y2=1.515
r36 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.355 $Y=0.655
+ $X2=2.355 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%C1 1 3 6 8 13
c23 8 0 6.08738e-21 $X=3.12 $Y=1.295
r24 10 13 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.865 $Y=1.35
+ $X2=3.07 $Y2=1.35
r25 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.35 $X2=3.07 $Y2=1.35
r26 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.515
+ $X2=2.865 $Y2=1.35
r27 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.865 $Y=1.515
+ $X2=2.865 $Y2=2.465
r28 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.185
+ $X2=2.865 $Y2=1.35
r29 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.865 $Y=1.185
+ $X2=2.865 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%X 1 2 7 8 9 10 11 12 13 22
r14 13 40 5.0187 $w=3.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.25 $Y=2.775
+ $X2=0.25 $Y2=2.91
r15 12 13 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.405
+ $X2=0.25 $Y2=2.775
r16 11 12 14.4985 $w=3.08e-07 $l=3.9e-07 $layer=LI1_cond $X=0.25 $Y=2.015
+ $X2=0.25 $Y2=2.405
r17 10 11 13.0115 $w=3.08e-07 $l=3.5e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=2.015
r18 9 10 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295 $X2=0.25
+ $Y2=1.665
r19 8 9 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=0.925 $X2=0.25
+ $Y2=1.295
r20 7 8 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=0.555 $X2=0.25
+ $Y2=0.925
r21 7 22 5.0187 $w=3.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.25 $Y=0.555
+ $X2=0.25 $Y2=0.42
r22 2 40 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r23 2 11 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.015
r24 1 22 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%VPWR 1 2 9 15 17 19 24 34 35 38 41
r44 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r48 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 29 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 25 38 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.715 $Y2=3.33
r54 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 24 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 19 38 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.715 $Y2=3.33
r60 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 17 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 17 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=3.33
r65 13 15 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=2.5
r66 9 12 30.4574 $w=2.78e-07 $l=7.4e-07 $layer=LI1_cond $X=0.715 $Y=2.21
+ $X2=0.715 $Y2=2.95
r67 7 38 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=3.33
r68 7 12 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=2.95
r69 2 15 300 $w=1.7e-07 $l=7.49617e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.835 $X2=1.68 $Y2=2.5
r70 1 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
r71 1 9 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%A_217_367# 1 2 7 9 11 13 15
r20 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=2.205
+ $X2=2.195 $Y2=2.12
r21 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.195 $Y=2.205
+ $X2=2.195 $Y2=2.56
r22 12 18 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.345 $Y=2.12
+ $X2=1.195 $Y2=2.12
r23 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=2.12
+ $X2=2.195 $Y2=2.12
r24 11 12 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.03 $Y=2.12
+ $X2=1.345 $Y2=2.12
r25 7 18 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=2.205 $X2=1.195
+ $Y2=2.12
r26 7 9 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=1.195 $Y=2.205
+ $X2=1.195 $Y2=2.56
r27 2 20 600 $w=1.7e-07 $l=3.65992e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.195 $Y2=2.12
r28 2 15 300 $w=1.7e-07 $l=8.1225e-07 $layer=licon1_PDIFF $count=2 $X=2.01
+ $Y=1.835 $X2=2.195 $Y2=2.56
r29 1 18 600 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=2.12
r30 1 9 300 $w=1.7e-07 $l=7.85016e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_1%VGND 1 2 9 11 18 25 26 31 37 39
r43 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 35 37 10.9376 $w=7.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=0.3
+ $X2=1.345 $Y2=0.3
r45 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 33 35 0.31067 $w=7.68e-07 $l=2e-08 $layer=LI1_cond $X=1.18 $Y=0.3 $X2=1.2
+ $Y2=0.3
r47 30 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r48 29 33 7.1454 $w=7.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.72 $Y=0.3 $X2=1.18
+ $Y2=0.3
r49 29 31 10.9376 $w=7.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.72 $Y=0.3
+ $X2=0.575 $Y2=0.3
r50 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 26 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r52 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 23 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.61
+ $Y2=0
r54 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=3.12
+ $Y2=0
r55 22 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r56 21 37 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.345
+ $Y2=0
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r58 18 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.61
+ $Y2=0
r59 18 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.16
+ $Y2=0
r60 16 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r61 15 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.575
+ $Y2=0
r62 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 11 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r64 11 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r65 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085 $X2=2.61
+ $Y2=0
r66 7 9 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.56
r67 2 9 182 $w=1.7e-07 $l=4.05123e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.235 $X2=2.61 $Y2=0.56
r68 1 33 91 $w=1.7e-07 $l=7.34745e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.235 $X2=1.18 $Y2=0.56
.ends

