* File: sky130_fd_sc_lp__nor3b_4.pxi.spice
* Created: Wed Sep  2 10:09:49 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3B_4%C_N N_C_N_M1013_g N_C_N_c_105_n N_C_N_M1007_g C_N
+ N_C_N_c_107_n PM_SKY130_FD_SC_LP__NOR3B_4%C_N
x_PM_SKY130_FD_SC_LP__NOR3B_4%A N_A_c_141_n N_A_M1001_g N_A_M1005_g N_A_c_142_n
+ N_A_M1014_g N_A_M1016_g N_A_c_143_n N_A_M1020_g N_A_M1017_g N_A_c_144_n
+ N_A_M1021_g N_A_M1025_g N_A_c_136_n N_A_c_137_n N_A_c_138_n N_A_c_139_n A A
+ PM_SKY130_FD_SC_LP__NOR3B_4%A
x_PM_SKY130_FD_SC_LP__NOR3B_4%A_38_367# N_A_38_367#_M1007_s N_A_38_367#_M1013_s
+ N_A_38_367#_M1002_g N_A_38_367#_c_233_n N_A_38_367#_M1006_g
+ N_A_38_367#_M1003_g N_A_38_367#_c_234_n N_A_38_367#_M1011_g
+ N_A_38_367#_M1015_g N_A_38_367#_c_235_n N_A_38_367#_M1018_g
+ N_A_38_367#_M1022_g N_A_38_367#_c_236_n N_A_38_367#_M1023_g
+ N_A_38_367#_c_226_n N_A_38_367#_c_227_n N_A_38_367#_c_238_n
+ N_A_38_367#_c_239_n N_A_38_367#_c_228_n N_A_38_367#_c_229_n
+ N_A_38_367#_c_230_n N_A_38_367#_c_231_n N_A_38_367#_c_232_n
+ N_A_38_367#_c_242_n PM_SKY130_FD_SC_LP__NOR3B_4%A_38_367#
x_PM_SKY130_FD_SC_LP__NOR3B_4%B N_B_M1004_g N_B_M1000_g N_B_M1009_g N_B_M1008_g
+ N_B_M1010_g N_B_M1012_g N_B_M1019_g N_B_M1024_g N_B_c_412_p B B N_B_c_365_n
+ N_B_c_366_n B N_B_c_367_n PM_SKY130_FD_SC_LP__NOR3B_4%B
x_PM_SKY130_FD_SC_LP__NOR3B_4%VPWR N_VPWR_M1013_d N_VPWR_M1014_s N_VPWR_M1021_s
+ N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n VPWR N_VPWR_c_447_n
+ N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_443_n N_VPWR_c_452_n
+ N_VPWR_c_453_n N_VPWR_c_454_n PM_SKY130_FD_SC_LP__NOR3B_4%VPWR
x_PM_SKY130_FD_SC_LP__NOR3B_4%A_211_367# N_A_211_367#_M1001_d
+ N_A_211_367#_M1020_d N_A_211_367#_M1000_s N_A_211_367#_M1012_s
+ N_A_211_367#_c_529_n N_A_211_367#_c_562_n N_A_211_367#_c_530_n
+ N_A_211_367#_c_566_n N_A_211_367#_c_528_n N_A_211_367#_c_550_n
+ N_A_211_367#_c_535_n N_A_211_367#_c_548_n N_A_211_367#_c_555_n
+ PM_SKY130_FD_SC_LP__NOR3B_4%A_211_367#
x_PM_SKY130_FD_SC_LP__NOR3B_4%A_576_367# N_A_576_367#_M1006_s
+ N_A_576_367#_M1011_s N_A_576_367#_M1023_s N_A_576_367#_M1008_d
+ N_A_576_367#_M1024_d N_A_576_367#_c_595_n N_A_576_367#_c_599_n
+ N_A_576_367#_c_630_n N_A_576_367#_c_605_n N_A_576_367#_c_593_n
+ N_A_576_367#_c_594_n N_A_576_367#_c_601_n N_A_576_367#_c_619_n
+ PM_SKY130_FD_SC_LP__NOR3B_4%A_576_367#
x_PM_SKY130_FD_SC_LP__NOR3B_4%Y N_Y_M1005_d N_Y_M1017_d N_Y_M1002_s N_Y_M1015_s
+ N_Y_M1004_d N_Y_M1010_d N_Y_M1006_d N_Y_M1018_d N_Y_c_753_p N_Y_c_651_n
+ N_Y_c_656_n N_Y_c_747_p N_Y_c_640_n N_Y_c_754_p N_Y_c_641_n N_Y_c_648_n
+ N_Y_c_681_n N_Y_c_682_n N_Y_c_649_n N_Y_c_687_n N_Y_c_704_n N_Y_c_757_p
+ N_Y_c_642_n N_Y_c_643_n N_Y_c_644_n N_Y_c_645_n N_Y_c_693_n N_Y_c_713_n
+ N_Y_c_646_n Y PM_SKY130_FD_SC_LP__NOR3B_4%Y
x_PM_SKY130_FD_SC_LP__NOR3B_4%VGND N_VGND_M1007_d N_VGND_M1016_s N_VGND_M1025_s
+ N_VGND_M1003_d N_VGND_M1022_d N_VGND_M1009_s N_VGND_M1019_s N_VGND_c_772_n
+ N_VGND_c_773_n N_VGND_c_774_n N_VGND_c_775_n N_VGND_c_776_n N_VGND_c_777_n
+ N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n
+ N_VGND_c_783_n N_VGND_c_784_n VGND N_VGND_c_785_n N_VGND_c_786_n
+ N_VGND_c_787_n N_VGND_c_788_n N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n
+ N_VGND_c_792_n N_VGND_c_793_n PM_SKY130_FD_SC_LP__NOR3B_4%VGND
cc_1 VNB N_C_N_M1013_g 0.00822276f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_2 VNB N_C_N_c_105_n 0.0206644f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.185
cc_3 VNB C_N 0.00446106f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C_N_c_107_n 0.0408719f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_5 VNB N_A_M1005_g 0.0212407f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_6 VNB N_A_M1016_g 0.0210533f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_7 VNB N_A_M1017_g 0.0214023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_M1025_g 0.0200596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_136_n 0.00132277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_c_137_n 0.0994482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_138_n 0.00342797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_c_139_n 0.00256805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A 0.00247834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_38_367#_M1002_g 0.0190482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_38_367#_M1003_g 0.0188632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_38_367#_M1015_g 0.0188632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_38_367#_M1022_g 0.0211677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_38_367#_c_226_n 0.0274314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_38_367#_c_227_n 0.031058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_38_367#_c_228_n 0.00119566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_38_367#_c_229_n 0.00133229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_38_367#_c_230_n 0.00131551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_38_367#_c_231_n 0.105293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_38_367#_c_232_n 0.0155939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_M1004_g 0.0213498f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_26 VNB N_B_M1000_g 0.00362641f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_27 VNB N_B_M1009_g 0.0191853f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.35
cc_28 VNB N_B_M1008_g 0.00350909f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.35
cc_29 VNB N_B_M1010_g 0.0193414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_M1012_g 0.00350659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_M1019_g 0.0224745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_M1024_g 0.00378138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_c_365_n 0.0858828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_366_n 0.00395591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_c_367_n 0.00122423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_443_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_640_n 0.00457497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_641_n 0.00321206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_642_n 0.0142399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_643_n 0.00200521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_644_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_645_n 0.00200198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_646_n 0.0024201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB Y 0.0259171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_772_n 0.00501153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_773_n 0.00436438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_774_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_775_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_776_n 3.20114e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_777_n 0.00429808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_778_n 3.20114e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_779_n 0.013077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_780_n 0.0253298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_781_n 0.0232161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_782_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_783_n 0.0167145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_784_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_785_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_786_n 0.015321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_787_n 0.015321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_788_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_789_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_790_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_791_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_792_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_793_n 0.33316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VPB N_C_N_M1013_g 0.0247245f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.465
cc_68 VPB N_A_c_141_n 0.0150696f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.515
cc_69 VPB N_A_c_142_n 0.0150524f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_70 VPB N_A_c_143_n 0.0150524f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.35
cc_71 VPB N_A_c_144_n 0.0186908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_c_137_n 0.0344234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_38_367#_c_233_n 0.0192473f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.35
cc_74 VPB N_A_38_367#_c_234_n 0.0152515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_38_367#_c_235_n 0.0152515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_38_367#_c_236_n 0.0153124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_38_367#_c_227_n 0.00230526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_38_367#_c_238_n 0.0494544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_38_367#_c_239_n 0.0129375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_38_367#_c_229_n 8.64304e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_38_367#_c_231_n 0.022123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_38_367#_c_242_n 0.0123255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_B_M1000_g 0.0185444f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.655
cc_84 VPB N_B_M1008_g 0.0184442f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.35
cc_85 VPB N_B_M1012_g 0.018426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_B_M1024_g 0.0235789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_444_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.35
cc_88 VPB N_VPWR_c_445_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_446_n 0.00737538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_447_n 0.017151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_448_n 0.012974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_449_n 0.012974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_450_n 0.0957238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_443_n 0.0495369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_452_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_453_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_454_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_211_367#_c_528_n 0.00947404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_576_367#_c_593_n 0.0083105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_576_367#_c_594_n 0.0326963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_Y_c_648_n 7.43414e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_Y_c_649_n 0.0210596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB Y 9.7145e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 N_C_N_c_105_n N_A_M1005_g 0.0155132f $X=0.71 $Y=1.185 $X2=0 $Y2=0
cc_105 C_N N_A_M1005_g 3.50142e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_106 N_C_N_M1013_g N_A_c_137_n 0.0287458f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_107 C_N N_A_c_137_n 0.00124111f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_108 N_C_N_c_107_n N_A_c_137_n 0.0114927f $X=0.55 $Y=1.35 $X2=0 $Y2=0
cc_109 C_N A 0.0236031f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_110 N_C_N_c_107_n A 6.24486e-19 $X=0.55 $Y=1.35 $X2=0 $Y2=0
cc_111 N_C_N_M1013_g N_A_38_367#_c_227_n 0.00465548f $X=0.55 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_C_N_c_105_n N_A_38_367#_c_227_n 0.00336606f $X=0.71 $Y=1.185 $X2=0
+ $Y2=0
cc_113 C_N N_A_38_367#_c_227_n 0.0251472f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_114 N_C_N_c_107_n N_A_38_367#_c_227_n 0.00836055f $X=0.55 $Y=1.35 $X2=0 $Y2=0
cc_115 N_C_N_M1013_g N_A_38_367#_c_239_n 0.0151374f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_116 C_N N_A_38_367#_c_239_n 0.0262423f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_117 N_C_N_c_107_n N_A_38_367#_c_239_n 0.0037534f $X=0.55 $Y=1.35 $X2=0 $Y2=0
cc_118 C_N N_A_38_367#_c_232_n 0.0110209f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_119 N_C_N_c_107_n N_A_38_367#_c_232_n 0.00708407f $X=0.55 $Y=1.35 $X2=0 $Y2=0
cc_120 N_C_N_c_107_n N_A_38_367#_c_242_n 0.00239209f $X=0.55 $Y=1.35 $X2=0 $Y2=0
cc_121 N_C_N_M1013_g N_VPWR_c_444_n 0.016366f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_122 N_C_N_M1013_g N_VPWR_c_447_n 0.00486043f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_123 N_C_N_M1013_g N_VPWR_c_443_n 0.00924348f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_124 N_C_N_c_105_n N_VGND_c_772_n 0.00399742f $X=0.71 $Y=1.185 $X2=0 $Y2=0
cc_125 N_C_N_c_105_n N_VGND_c_781_n 0.00585385f $X=0.71 $Y=1.185 $X2=0 $Y2=0
cc_126 N_C_N_c_105_n N_VGND_c_793_n 0.0118478f $X=0.71 $Y=1.185 $X2=0 $Y2=0
cc_127 N_A_M1025_g N_A_38_367#_M1002_g 0.0210713f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_128 N_A_c_141_n N_A_38_367#_c_239_n 0.0115424f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_129 N_A_c_142_n N_A_38_367#_c_239_n 0.0076791f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_130 N_A_c_143_n N_A_38_367#_c_239_n 0.0076791f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_131 N_A_c_144_n N_A_38_367#_c_239_n 0.0106725f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_132 N_A_c_137_n N_A_38_367#_c_239_n 0.0420295f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_133 N_A_c_138_n N_A_38_367#_c_239_n 0.0935688f $X=1.785 $Y=1.355 $X2=0 $Y2=0
cc_134 A N_A_38_367#_c_239_n 0.0194927f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A_c_136_n N_A_38_367#_c_228_n 0.012772f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_136 N_A_c_137_n N_A_38_367#_c_228_n 2.22064e-19 $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_137 N_A_c_136_n N_A_38_367#_c_229_n 0.00119237f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_138 N_A_c_137_n N_A_38_367#_c_229_n 0.00328997f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_139 N_A_M1025_g N_A_38_367#_c_231_n 0.0013464f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_140 N_A_c_136_n N_A_38_367#_c_231_n 2.9866e-19 $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_141 N_A_c_137_n N_A_38_367#_c_231_n 0.02491f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_142 N_A_c_141_n N_VPWR_c_444_n 0.0142032f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_143 N_A_c_142_n N_VPWR_c_444_n 6.95678e-19 $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_144 N_A_c_141_n N_VPWR_c_445_n 6.47302e-19 $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_145 N_A_c_142_n N_VPWR_c_445_n 0.0117424f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_146 N_A_c_143_n N_VPWR_c_445_n 0.0117345f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_147 N_A_c_144_n N_VPWR_c_445_n 6.19012e-19 $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_148 N_A_c_143_n N_VPWR_c_446_n 5.70917e-19 $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_149 N_A_c_144_n N_VPWR_c_446_n 0.0110361f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_150 N_A_c_141_n N_VPWR_c_448_n 0.00486043f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_151 N_A_c_142_n N_VPWR_c_448_n 0.00486043f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_152 N_A_c_143_n N_VPWR_c_449_n 0.00486043f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_153 N_A_c_144_n N_VPWR_c_449_n 0.00486043f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_154 N_A_c_141_n N_VPWR_c_443_n 0.00824727f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_155 N_A_c_142_n N_VPWR_c_443_n 0.00824727f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_156 N_A_c_143_n N_VPWR_c_443_n 0.00824727f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_157 N_A_c_144_n N_VPWR_c_443_n 0.004514f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_158 N_A_c_137_n N_A_211_367#_c_529_n 5.4695e-19 $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_159 N_A_c_142_n N_A_211_367#_c_530_n 0.0125125f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_160 N_A_c_143_n N_A_211_367#_c_530_n 0.0125125f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_161 N_A_c_137_n N_A_211_367#_c_530_n 4.8451e-19 $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_162 N_A_c_144_n N_A_211_367#_c_528_n 0.0123866f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_163 N_A_c_137_n N_A_211_367#_c_528_n 0.00134043f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_164 N_A_c_144_n N_A_211_367#_c_535_n 0.0137002f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A_c_137_n N_A_211_367#_c_535_n 5.4695e-19 $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_166 N_A_c_144_n N_A_576_367#_c_595_n 9.87213e-19 $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_167 N_A_M1016_g N_Y_c_651_n 0.0104467f $X=1.65 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A_M1017_g N_Y_c_651_n 0.0107139f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A_c_136_n N_Y_c_651_n 0.00978193f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_170 N_A_c_137_n N_Y_c_651_n 0.00177608f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_171 N_A_c_138_n N_Y_c_651_n 0.0267731f $X=1.785 $Y=1.355 $X2=0 $Y2=0
cc_172 N_A_c_137_n N_Y_c_656_n 6.23337e-19 $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_173 N_A_c_138_n N_Y_c_656_n 0.0185798f $X=1.785 $Y=1.355 $X2=0 $Y2=0
cc_174 N_A_M1025_g N_Y_c_640_n 0.0125778f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_175 N_A_c_136_n N_Y_c_640_n 0.0150012f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_176 N_A_c_137_n N_Y_c_640_n 5.06935e-19 $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_177 N_A_M1016_g N_Y_c_643_n 7.4342e-19 $X=1.65 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A_M1017_g N_Y_c_643_n 0.00521553f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A_c_136_n N_Y_c_643_n 0.0207928f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_180 N_A_c_137_n N_Y_c_643_n 0.00268352f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_181 N_A_M1005_g N_VGND_c_772_n 0.00257735f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_182 N_A_c_137_n N_VGND_c_772_n 0.00598147f $X=2.52 $Y=1.44 $X2=0 $Y2=0
cc_183 A N_VGND_c_772_n 0.00485564f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A_M1016_g N_VGND_c_773_n 0.00242526f $X=1.65 $Y=0.655 $X2=0 $Y2=0
cc_185 N_A_M1017_g N_VGND_c_773_n 0.00237608f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_186 N_A_M1017_g N_VGND_c_774_n 0.00585385f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_187 N_A_M1025_g N_VGND_c_774_n 0.00486043f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A_M1017_g N_VGND_c_775_n 6.24575e-19 $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A_M1025_g N_VGND_c_775_n 0.010031f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_190 N_A_M1005_g N_VGND_c_783_n 0.00585385f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A_M1016_g N_VGND_c_783_n 0.00585385f $X=1.65 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_M1005_g N_VGND_c_793_n 0.0107286f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A_M1016_g N_VGND_c_793_n 0.00644678f $X=1.65 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A_M1017_g N_VGND_c_793_n 0.00642981f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_M1025_g N_VGND_c_793_n 0.00824727f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A_38_367#_M1022_g N_B_M1004_g 0.029311f $X=4.31 $Y=0.655 $X2=0 $Y2=0
cc_197 N_A_38_367#_c_231_n N_B_M1000_g 0.0615891f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_198 N_A_38_367#_c_230_n N_B_c_365_n 7.5017e-19 $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_199 N_A_38_367#_c_231_n N_B_c_365_n 0.0241584f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_200 N_A_38_367#_M1022_g N_B_c_366_n 2.1494e-19 $X=4.31 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_38_367#_c_230_n N_B_c_366_n 0.0100744f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_202 N_A_38_367#_c_231_n N_B_c_366_n 6.58753e-19 $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_203 N_A_38_367#_c_239_n N_VPWR_M1013_d 0.00201607f $X=2.895 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_38_367#_c_239_n N_VPWR_M1014_s 0.00176891f $X=2.895 $Y=1.79 $X2=0
+ $Y2=0
cc_205 N_A_38_367#_c_239_n N_VPWR_M1021_s 0.00355171f $X=2.895 $Y=1.79 $X2=0
+ $Y2=0
cc_206 N_A_38_367#_c_239_n N_VPWR_c_444_n 0.0135931f $X=2.895 $Y=1.79 $X2=0
+ $Y2=0
cc_207 N_A_38_367#_c_233_n N_VPWR_c_446_n 0.00345279f $X=3.22 $Y=1.725 $X2=0
+ $Y2=0
cc_208 N_A_38_367#_c_238_n N_VPWR_c_447_n 0.0228053f $X=0.315 $Y=1.98 $X2=0
+ $Y2=0
cc_209 N_A_38_367#_c_233_n N_VPWR_c_450_n 0.00357877f $X=3.22 $Y=1.725 $X2=0
+ $Y2=0
cc_210 N_A_38_367#_c_234_n N_VPWR_c_450_n 0.00357877f $X=3.65 $Y=1.725 $X2=0
+ $Y2=0
cc_211 N_A_38_367#_c_235_n N_VPWR_c_450_n 0.00357877f $X=4.08 $Y=1.725 $X2=0
+ $Y2=0
cc_212 N_A_38_367#_c_236_n N_VPWR_c_450_n 0.00357877f $X=4.51 $Y=1.725 $X2=0
+ $Y2=0
cc_213 N_A_38_367#_M1013_s N_VPWR_c_443_n 0.00423245f $X=0.19 $Y=1.835 $X2=0
+ $Y2=0
cc_214 N_A_38_367#_c_233_n N_VPWR_c_443_n 0.0068216f $X=3.22 $Y=1.725 $X2=0
+ $Y2=0
cc_215 N_A_38_367#_c_234_n N_VPWR_c_443_n 0.00542194f $X=3.65 $Y=1.725 $X2=0
+ $Y2=0
cc_216 N_A_38_367#_c_235_n N_VPWR_c_443_n 0.00542194f $X=4.08 $Y=1.725 $X2=0
+ $Y2=0
cc_217 N_A_38_367#_c_236_n N_VPWR_c_443_n 0.00537654f $X=4.51 $Y=1.725 $X2=0
+ $Y2=0
cc_218 N_A_38_367#_c_238_n N_VPWR_c_443_n 0.0125522f $X=0.315 $Y=1.98 $X2=0
+ $Y2=0
cc_219 N_A_38_367#_c_239_n N_A_211_367#_M1001_d 0.00176461f $X=2.895 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_220 N_A_38_367#_c_239_n N_A_211_367#_M1020_d 0.00176461f $X=2.895 $Y=1.79
+ $X2=0 $Y2=0
cc_221 N_A_38_367#_c_239_n N_A_211_367#_c_529_n 0.0135055f $X=2.895 $Y=1.79
+ $X2=0 $Y2=0
cc_222 N_A_38_367#_c_239_n N_A_211_367#_c_530_n 0.0324646f $X=2.895 $Y=1.79
+ $X2=0 $Y2=0
cc_223 N_A_38_367#_c_233_n N_A_211_367#_c_528_n 0.0171083f $X=3.22 $Y=1.725
+ $X2=0 $Y2=0
cc_224 N_A_38_367#_c_234_n N_A_211_367#_c_528_n 0.0105479f $X=3.65 $Y=1.725
+ $X2=0 $Y2=0
cc_225 N_A_38_367#_c_235_n N_A_211_367#_c_528_n 0.0114768f $X=4.08 $Y=1.725
+ $X2=0 $Y2=0
cc_226 N_A_38_367#_c_236_n N_A_211_367#_c_528_n 0.0130923f $X=4.51 $Y=1.725
+ $X2=0 $Y2=0
cc_227 N_A_38_367#_c_239_n N_A_211_367#_c_528_n 0.0287157f $X=2.895 $Y=1.79
+ $X2=0 $Y2=0
cc_228 N_A_38_367#_c_231_n N_A_211_367#_c_528_n 8.86346e-19 $X=4.42 $Y=1.42
+ $X2=0 $Y2=0
cc_229 N_A_38_367#_c_239_n N_A_211_367#_c_535_n 0.0152326f $X=2.895 $Y=1.79
+ $X2=0 $Y2=0
cc_230 N_A_38_367#_c_236_n N_A_211_367#_c_548_n 0.00235178f $X=4.51 $Y=1.725
+ $X2=0 $Y2=0
cc_231 N_A_38_367#_c_239_n N_A_576_367#_M1006_s 0.00406843f $X=2.895 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_232 N_A_38_367#_c_233_n N_A_576_367#_c_595_n 0.0149547f $X=3.22 $Y=1.725
+ $X2=0 $Y2=0
cc_233 N_A_38_367#_c_234_n N_A_576_367#_c_595_n 0.0144853f $X=3.65 $Y=1.725
+ $X2=0 $Y2=0
cc_234 N_A_38_367#_c_235_n N_A_576_367#_c_599_n 0.00840109f $X=4.08 $Y=1.725
+ $X2=0 $Y2=0
cc_235 N_A_38_367#_c_236_n N_A_576_367#_c_599_n 0.00961806f $X=4.51 $Y=1.725
+ $X2=0 $Y2=0
cc_236 N_A_38_367#_c_235_n N_A_576_367#_c_601_n 0.00572851f $X=4.08 $Y=1.725
+ $X2=0 $Y2=0
cc_237 N_A_38_367#_c_236_n N_A_576_367#_c_601_n 0.00100996f $X=4.51 $Y=1.725
+ $X2=0 $Y2=0
cc_238 N_A_38_367#_M1002_g N_Y_c_640_n 0.0131471f $X=3.02 $Y=0.655 $X2=0 $Y2=0
cc_239 N_A_38_367#_c_239_n N_Y_c_640_n 0.00698972f $X=2.895 $Y=1.79 $X2=0 $Y2=0
cc_240 N_A_38_367#_c_228_n N_Y_c_640_n 0.012909f $X=2.98 $Y=1.505 $X2=0 $Y2=0
cc_241 N_A_38_367#_c_230_n N_Y_c_640_n 0.00520336f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_242 N_A_38_367#_c_231_n N_Y_c_640_n 0.00121703f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_243 N_A_38_367#_M1003_g N_Y_c_641_n 0.0131657f $X=3.45 $Y=0.655 $X2=0 $Y2=0
cc_244 N_A_38_367#_M1015_g N_Y_c_641_n 0.0126243f $X=3.88 $Y=0.655 $X2=0 $Y2=0
cc_245 N_A_38_367#_c_230_n N_Y_c_641_n 0.0469649f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_246 N_A_38_367#_c_231_n N_Y_c_641_n 0.00286055f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_247 N_A_38_367#_c_233_n N_Y_c_648_n 0.0011322f $X=3.22 $Y=1.725 $X2=0 $Y2=0
cc_248 N_A_38_367#_c_234_n N_Y_c_648_n 0.0140044f $X=3.65 $Y=1.725 $X2=0 $Y2=0
cc_249 N_A_38_367#_c_235_n N_Y_c_648_n 0.0142373f $X=4.08 $Y=1.725 $X2=0 $Y2=0
cc_250 N_A_38_367#_c_239_n N_Y_c_648_n 0.0100682f $X=2.895 $Y=1.79 $X2=0 $Y2=0
cc_251 N_A_38_367#_c_229_n N_Y_c_648_n 0.00163011f $X=2.98 $Y=1.705 $X2=0 $Y2=0
cc_252 N_A_38_367#_c_230_n N_Y_c_648_n 0.0915398f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_253 N_A_38_367#_c_231_n N_Y_c_648_n 0.0206792f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_254 N_A_38_367#_M1022_g N_Y_c_681_n 0.00908188f $X=4.31 $Y=0.655 $X2=0 $Y2=0
cc_255 N_A_38_367#_M1022_g N_Y_c_682_n 0.0132054f $X=4.31 $Y=0.655 $X2=0 $Y2=0
cc_256 N_A_38_367#_c_230_n N_Y_c_682_n 0.0137058f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_257 N_A_38_367#_c_231_n N_Y_c_682_n 0.0050641f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_258 N_A_38_367#_c_236_n N_Y_c_649_n 0.00816576f $X=4.51 $Y=1.725 $X2=0 $Y2=0
cc_259 N_A_38_367#_c_231_n N_Y_c_649_n 0.00395984f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_260 N_A_38_367#_M1022_g N_Y_c_687_n 6.18173e-19 $X=4.31 $Y=0.655 $X2=0 $Y2=0
cc_261 N_A_38_367#_c_230_n N_Y_c_644_n 0.0153881f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_262 N_A_38_367#_c_231_n N_Y_c_644_n 0.00296179f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_263 N_A_38_367#_M1022_g N_Y_c_645_n 0.00424531f $X=4.31 $Y=0.655 $X2=0 $Y2=0
cc_264 N_A_38_367#_c_230_n N_Y_c_645_n 0.0207877f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_265 N_A_38_367#_c_231_n N_Y_c_645_n 0.00296179f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_266 N_A_38_367#_c_231_n N_Y_c_693_n 0.00660333f $X=4.42 $Y=1.42 $X2=0 $Y2=0
cc_267 N_A_38_367#_M1002_g N_VGND_c_775_n 0.00993915f $X=3.02 $Y=0.655 $X2=0
+ $Y2=0
cc_268 N_A_38_367#_M1003_g N_VGND_c_775_n 6.0835e-19 $X=3.45 $Y=0.655 $X2=0
+ $Y2=0
cc_269 N_A_38_367#_M1002_g N_VGND_c_776_n 6.0835e-19 $X=3.02 $Y=0.655 $X2=0
+ $Y2=0
cc_270 N_A_38_367#_M1003_g N_VGND_c_776_n 0.0099749f $X=3.45 $Y=0.655 $X2=0
+ $Y2=0
cc_271 N_A_38_367#_M1015_g N_VGND_c_776_n 0.0101222f $X=3.88 $Y=0.655 $X2=0
+ $Y2=0
cc_272 N_A_38_367#_M1022_g N_VGND_c_776_n 6.88997e-19 $X=4.31 $Y=0.655 $X2=0
+ $Y2=0
cc_273 N_A_38_367#_M1022_g N_VGND_c_777_n 0.00451036f $X=4.31 $Y=0.655 $X2=0
+ $Y2=0
cc_274 N_A_38_367#_c_226_n N_VGND_c_781_n 0.0343027f $X=0.495 $Y=0.42 $X2=0
+ $Y2=0
cc_275 N_A_38_367#_M1002_g N_VGND_c_785_n 0.00486043f $X=3.02 $Y=0.655 $X2=0
+ $Y2=0
cc_276 N_A_38_367#_M1003_g N_VGND_c_785_n 0.00486043f $X=3.45 $Y=0.655 $X2=0
+ $Y2=0
cc_277 N_A_38_367#_M1015_g N_VGND_c_786_n 0.00486043f $X=3.88 $Y=0.655 $X2=0
+ $Y2=0
cc_278 N_A_38_367#_M1022_g N_VGND_c_786_n 0.0055654f $X=4.31 $Y=0.655 $X2=0
+ $Y2=0
cc_279 N_A_38_367#_M1007_s N_VGND_c_793_n 0.0040649f $X=0.37 $Y=0.235 $X2=0
+ $Y2=0
cc_280 N_A_38_367#_M1002_g N_VGND_c_793_n 0.00824727f $X=3.02 $Y=0.655 $X2=0
+ $Y2=0
cc_281 N_A_38_367#_M1003_g N_VGND_c_793_n 0.00824727f $X=3.45 $Y=0.655 $X2=0
+ $Y2=0
cc_282 N_A_38_367#_M1015_g N_VGND_c_793_n 0.00824727f $X=3.88 $Y=0.655 $X2=0
+ $Y2=0
cc_283 N_A_38_367#_M1022_g N_VGND_c_793_n 0.0103748f $X=4.31 $Y=0.655 $X2=0
+ $Y2=0
cc_284 N_A_38_367#_c_226_n N_VGND_c_793_n 0.0187726f $X=0.495 $Y=0.42 $X2=0
+ $Y2=0
cc_285 N_B_M1000_g N_VPWR_c_450_n 0.00357877f $X=4.94 $Y=2.465 $X2=0 $Y2=0
cc_286 N_B_M1008_g N_VPWR_c_450_n 0.00357877f $X=5.37 $Y=2.465 $X2=0 $Y2=0
cc_287 N_B_M1012_g N_VPWR_c_450_n 0.00357877f $X=5.8 $Y=2.465 $X2=0 $Y2=0
cc_288 N_B_M1024_g N_VPWR_c_450_n 0.00357877f $X=6.23 $Y=2.465 $X2=0 $Y2=0
cc_289 N_B_M1000_g N_VPWR_c_443_n 0.00536745f $X=4.94 $Y=2.465 $X2=0 $Y2=0
cc_290 N_B_M1008_g N_VPWR_c_443_n 0.0053512f $X=5.37 $Y=2.465 $X2=0 $Y2=0
cc_291 N_B_M1012_g N_VPWR_c_443_n 0.0053512f $X=5.8 $Y=2.465 $X2=0 $Y2=0
cc_292 N_B_M1024_g N_VPWR_c_443_n 0.00629771f $X=6.23 $Y=2.465 $X2=0 $Y2=0
cc_293 N_B_M1000_g N_A_211_367#_c_528_n 0.0105403f $X=4.94 $Y=2.465 $X2=0 $Y2=0
cc_294 N_B_M1008_g N_A_211_367#_c_550_n 0.0105896f $X=5.37 $Y=2.465 $X2=0 $Y2=0
cc_295 N_B_M1012_g N_A_211_367#_c_550_n 0.0114269f $X=5.8 $Y=2.465 $X2=0 $Y2=0
cc_296 N_B_M1000_g N_A_211_367#_c_548_n 0.0123455f $X=4.94 $Y=2.465 $X2=0 $Y2=0
cc_297 N_B_M1008_g N_A_211_367#_c_548_n 0.0093351f $X=5.37 $Y=2.465 $X2=0 $Y2=0
cc_298 N_B_M1012_g N_A_211_367#_c_548_n 6.15006e-19 $X=5.8 $Y=2.465 $X2=0 $Y2=0
cc_299 N_B_M1008_g N_A_211_367#_c_555_n 5.2821e-19 $X=5.37 $Y=2.465 $X2=0 $Y2=0
cc_300 N_B_M1012_g N_A_211_367#_c_555_n 0.00880696f $X=5.8 $Y=2.465 $X2=0 $Y2=0
cc_301 N_B_M1024_g N_A_211_367#_c_555_n 0.00935773f $X=6.23 $Y=2.465 $X2=0 $Y2=0
cc_302 N_B_M1000_g N_A_576_367#_c_599_n 0.00940986f $X=4.94 $Y=2.465 $X2=0 $Y2=0
cc_303 N_B_M1008_g N_A_576_367#_c_599_n 0.0103643f $X=5.37 $Y=2.465 $X2=0 $Y2=0
cc_304 N_B_M1012_g N_A_576_367#_c_605_n 0.0121057f $X=5.8 $Y=2.465 $X2=0 $Y2=0
cc_305 N_B_M1024_g N_A_576_367#_c_605_n 0.0121057f $X=6.23 $Y=2.465 $X2=0 $Y2=0
cc_306 N_B_M1004_g N_Y_c_681_n 6.18173e-19 $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_307 N_B_M1004_g N_Y_c_682_n 0.0129635f $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_308 N_B_c_366_n N_Y_c_682_n 0.00421253f $X=5.523 $Y=1.357 $X2=0 $Y2=0
cc_309 N_B_M1000_g N_Y_c_649_n 0.0121039f $X=4.94 $Y=2.465 $X2=0 $Y2=0
cc_310 N_B_M1008_g N_Y_c_649_n 0.0108682f $X=5.37 $Y=2.465 $X2=0 $Y2=0
cc_311 N_B_M1012_g N_Y_c_649_n 0.0108682f $X=5.8 $Y=2.465 $X2=0 $Y2=0
cc_312 N_B_M1024_g N_Y_c_649_n 0.0170787f $X=6.23 $Y=2.465 $X2=0 $Y2=0
cc_313 N_B_c_365_n N_Y_c_649_n 0.010715f $X=6.23 $Y=1.42 $X2=0 $Y2=0
cc_314 N_B_c_366_n N_Y_c_649_n 0.0974227f $X=5.523 $Y=1.357 $X2=0 $Y2=0
cc_315 N_B_M1004_g N_Y_c_687_n 0.00856802f $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_316 N_B_M1009_g N_Y_c_704_n 0.0122129f $X=5.3 $Y=0.655 $X2=0 $Y2=0
cc_317 N_B_M1010_g N_Y_c_704_n 0.0128965f $X=5.73 $Y=0.655 $X2=0 $Y2=0
cc_318 N_B_c_412_p N_Y_c_704_n 0.00660894f $X=6.05 $Y=1.42 $X2=0 $Y2=0
cc_319 N_B_c_365_n N_Y_c_704_n 6.36477e-19 $X=6.23 $Y=1.42 $X2=0 $Y2=0
cc_320 N_B_c_366_n N_Y_c_704_n 0.030935f $X=5.523 $Y=1.357 $X2=0 $Y2=0
cc_321 N_B_M1019_g N_Y_c_642_n 0.014442f $X=6.16 $Y=0.655 $X2=0 $Y2=0
cc_322 N_B_c_412_p N_Y_c_642_n 0.0115008f $X=6.05 $Y=1.42 $X2=0 $Y2=0
cc_323 N_B_c_365_n N_Y_c_642_n 0.00229216f $X=6.23 $Y=1.42 $X2=0 $Y2=0
cc_324 N_B_M1004_g N_Y_c_645_n 6.11592e-19 $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_325 N_B_M1004_g N_Y_c_713_n 5.79575e-19 $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_326 N_B_c_365_n N_Y_c_713_n 6.96874e-19 $X=6.23 $Y=1.42 $X2=0 $Y2=0
cc_327 N_B_c_366_n N_Y_c_713_n 0.0186516f $X=5.523 $Y=1.357 $X2=0 $Y2=0
cc_328 N_B_M1010_g N_Y_c_646_n 0.00199913f $X=5.73 $Y=0.655 $X2=0 $Y2=0
cc_329 N_B_c_412_p N_Y_c_646_n 0.0152561f $X=6.05 $Y=1.42 $X2=0 $Y2=0
cc_330 N_B_c_365_n N_Y_c_646_n 0.00285313f $X=6.23 $Y=1.42 $X2=0 $Y2=0
cc_331 N_B_M1019_g Y 0.00362658f $X=6.16 $Y=0.655 $X2=0 $Y2=0
cc_332 N_B_c_412_p Y 0.0138073f $X=6.05 $Y=1.42 $X2=0 $Y2=0
cc_333 N_B_c_365_n Y 0.016182f $X=6.23 $Y=1.42 $X2=0 $Y2=0
cc_334 N_B_M1004_g N_VGND_c_777_n 0.00451036f $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_335 N_B_M1004_g N_VGND_c_778_n 6.31488e-19 $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_336 N_B_M1009_g N_VGND_c_778_n 0.010537f $X=5.3 $Y=0.655 $X2=0 $Y2=0
cc_337 N_B_M1010_g N_VGND_c_778_n 0.0103898f $X=5.73 $Y=0.655 $X2=0 $Y2=0
cc_338 N_B_M1019_g N_VGND_c_778_n 5.75816e-19 $X=6.16 $Y=0.655 $X2=0 $Y2=0
cc_339 N_B_M1010_g N_VGND_c_780_n 6.0835e-19 $X=5.73 $Y=0.655 $X2=0 $Y2=0
cc_340 N_B_M1019_g N_VGND_c_780_n 0.0110384f $X=6.16 $Y=0.655 $X2=0 $Y2=0
cc_341 N_B_M1004_g N_VGND_c_787_n 0.0055654f $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_342 N_B_M1009_g N_VGND_c_787_n 0.00486043f $X=5.3 $Y=0.655 $X2=0 $Y2=0
cc_343 N_B_M1010_g N_VGND_c_788_n 0.00486043f $X=5.73 $Y=0.655 $X2=0 $Y2=0
cc_344 N_B_M1019_g N_VGND_c_788_n 0.00486043f $X=6.16 $Y=0.655 $X2=0 $Y2=0
cc_345 N_B_M1004_g N_VGND_c_793_n 0.0103748f $X=4.87 $Y=0.655 $X2=0 $Y2=0
cc_346 N_B_M1009_g N_VGND_c_793_n 0.00824727f $X=5.3 $Y=0.655 $X2=0 $Y2=0
cc_347 N_B_M1010_g N_VGND_c_793_n 0.00824727f $X=5.73 $Y=0.655 $X2=0 $Y2=0
cc_348 N_B_M1019_g N_VGND_c_793_n 0.00824727f $X=6.16 $Y=0.655 $X2=0 $Y2=0
cc_349 N_VPWR_c_443_n N_A_211_367#_M1001_d 0.00536823f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_350 N_VPWR_c_443_n N_A_211_367#_M1020_d 0.00408265f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_443_n N_A_211_367#_M1000_s 0.00225186f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_443_n N_A_211_367#_M1012_s 0.00225186f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_448_n N_A_211_367#_c_562_n 0.0117038f $X=1.46 $Y=3.33 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_443_n N_A_211_367#_c_562_n 0.00727431f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_355 N_VPWR_M1014_s N_A_211_367#_c_530_n 0.00336057f $X=1.485 $Y=1.835 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_445_n N_A_211_367#_c_530_n 0.0171443f $X=1.625 $Y=2.52 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_449_n N_A_211_367#_c_566_n 0.0117038f $X=2.32 $Y=3.33 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_443_n N_A_211_367#_c_566_n 0.00727431f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_359 N_VPWR_M1021_s N_A_211_367#_c_528_n 0.0060987f $X=2.345 $Y=1.835 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_446_n N_A_211_367#_c_528_n 0.0215105f $X=2.485 $Y=2.83 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_443_n N_A_211_367#_c_528_n 0.0166564f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_443_n N_A_211_367#_c_535_n 0.00237405f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_363 N_VPWR_c_443_n N_A_576_367#_M1006_s 0.00229095f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_364 N_VPWR_c_443_n N_A_576_367#_M1011_s 0.00225186f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_443_n N_A_576_367#_M1023_s 0.00223577f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_443_n N_A_576_367#_M1008_d 0.00223565f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_443_n N_A_576_367#_M1024_d 0.00215161f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_446_n N_A_576_367#_c_595_n 0.026781f $X=2.485 $Y=2.83 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_450_n N_A_576_367#_c_595_n 0.147462f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_370 N_VPWR_c_443_n N_A_576_367#_c_595_n 0.0940986f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_450_n N_A_576_367#_c_605_n 0.0363306f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_443_n N_A_576_367#_c_605_n 0.0237343f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_450_n N_A_576_367#_c_593_n 0.0179183f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_443_n N_A_576_367#_c_593_n 0.0101082f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_450_n N_A_576_367#_c_619_n 0.0125483f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_443_n N_A_576_367#_c_619_n 0.00739237f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_443_n N_Y_M1006_d 0.00225186f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_378 N_VPWR_c_443_n N_Y_M1018_d 0.00225186f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_379 N_A_211_367#_c_528_n N_A_576_367#_M1006_s 0.00719926f $X=4.99 $Y=2.41
+ $X2=-0.19 $Y2=1.655
cc_380 N_A_211_367#_c_528_n N_A_576_367#_M1011_s 0.00346119f $X=4.99 $Y=2.41
+ $X2=0 $Y2=0
cc_381 N_A_211_367#_c_528_n N_A_576_367#_M1023_s 0.00542592f $X=4.99 $Y=2.41
+ $X2=0 $Y2=0
cc_382 N_A_211_367#_c_550_n N_A_576_367#_M1008_d 0.00340214f $X=5.85 $Y=2.115
+ $X2=0 $Y2=0
cc_383 N_A_211_367#_c_528_n N_A_576_367#_c_595_n 0.0623731f $X=4.99 $Y=2.41
+ $X2=0 $Y2=0
cc_384 N_A_211_367#_M1000_s N_A_576_367#_c_599_n 0.00334014f $X=5.015 $Y=1.835
+ $X2=0 $Y2=0
cc_385 N_A_211_367#_c_528_n N_A_576_367#_c_599_n 0.0242378f $X=4.99 $Y=2.41
+ $X2=0 $Y2=0
cc_386 N_A_211_367#_c_550_n N_A_576_367#_c_599_n 0.0027272f $X=5.85 $Y=2.115
+ $X2=0 $Y2=0
cc_387 N_A_211_367#_c_548_n N_A_576_367#_c_599_n 0.0162722f $X=5.155 $Y=2.11
+ $X2=0 $Y2=0
cc_388 N_A_211_367#_c_550_n N_A_576_367#_c_630_n 0.0135898f $X=5.85 $Y=2.115
+ $X2=0 $Y2=0
cc_389 N_A_211_367#_M1012_s N_A_576_367#_c_605_n 0.00337788f $X=5.875 $Y=1.835
+ $X2=0 $Y2=0
cc_390 N_A_211_367#_c_555_n N_A_576_367#_c_605_n 0.0153963f $X=6.015 $Y=2.11
+ $X2=0 $Y2=0
cc_391 N_A_211_367#_c_528_n N_Y_M1006_d 0.00346119f $X=4.99 $Y=2.41 $X2=0 $Y2=0
cc_392 N_A_211_367#_c_528_n N_Y_M1018_d 0.00424197f $X=4.99 $Y=2.41 $X2=0 $Y2=0
cc_393 N_A_211_367#_c_528_n N_Y_c_648_n 0.0584969f $X=4.99 $Y=2.41 $X2=0 $Y2=0
cc_394 N_A_211_367#_M1000_s N_Y_c_649_n 0.00176773f $X=5.015 $Y=1.835 $X2=0
+ $Y2=0
cc_395 N_A_211_367#_M1012_s N_Y_c_649_n 0.00176773f $X=5.875 $Y=1.835 $X2=0
+ $Y2=0
cc_396 N_A_211_367#_c_528_n N_Y_c_649_n 0.0138935f $X=4.99 $Y=2.41 $X2=0 $Y2=0
cc_397 N_A_211_367#_c_550_n N_Y_c_649_n 0.0292216f $X=5.85 $Y=2.115 $X2=0 $Y2=0
cc_398 N_A_211_367#_c_548_n N_Y_c_649_n 0.0171443f $X=5.155 $Y=2.11 $X2=0 $Y2=0
cc_399 N_A_211_367#_c_555_n N_Y_c_649_n 0.0172972f $X=6.015 $Y=2.11 $X2=0 $Y2=0
cc_400 N_A_576_367#_c_595_n N_Y_M1006_d 0.00341909f $X=3.825 $Y=2.87 $X2=0 $Y2=0
cc_401 N_A_576_367#_c_599_n N_Y_M1018_d 0.00417318f $X=5.49 $Y=2.975 $X2=0 $Y2=0
cc_402 N_A_576_367#_M1011_s N_Y_c_648_n 0.00186947f $X=3.725 $Y=1.835 $X2=0
+ $Y2=0
cc_403 N_A_576_367#_M1023_s N_Y_c_649_n 0.00290659f $X=4.585 $Y=1.835 $X2=0
+ $Y2=0
cc_404 N_A_576_367#_M1008_d N_Y_c_649_n 0.00177204f $X=5.445 $Y=1.835 $X2=0
+ $Y2=0
cc_405 N_A_576_367#_M1024_d N_Y_c_649_n 0.00237563f $X=6.305 $Y=1.835 $X2=0
+ $Y2=0
cc_406 N_A_576_367#_c_594_n N_Y_c_649_n 0.0221758f $X=6.445 $Y=2.19 $X2=0 $Y2=0
cc_407 N_Y_c_651_n N_VGND_M1016_s 0.0050516f $X=2.21 $Y=0.93 $X2=0 $Y2=0
cc_408 N_Y_c_640_n N_VGND_M1025_s 0.00176461f $X=3.14 $Y=1.07 $X2=0 $Y2=0
cc_409 N_Y_c_641_n N_VGND_M1003_d 0.00176461f $X=4 $Y=1.07 $X2=0 $Y2=0
cc_410 N_Y_c_682_n N_VGND_M1022_d 0.00807729f $X=4.925 $Y=0.955 $X2=0 $Y2=0
cc_411 N_Y_c_704_n N_VGND_M1009_s 0.00331844f $X=5.84 $Y=0.955 $X2=0 $Y2=0
cc_412 N_Y_c_642_n N_VGND_M1019_s 0.00267403f $X=6.385 $Y=1.07 $X2=0 $Y2=0
cc_413 N_Y_c_651_n N_VGND_c_773_n 0.019584f $X=2.21 $Y=0.93 $X2=0 $Y2=0
cc_414 N_Y_c_747_p N_VGND_c_774_n 0.0138717f $X=2.375 $Y=0.42 $X2=0 $Y2=0
cc_415 N_Y_c_640_n N_VGND_c_775_n 0.0170777f $X=3.14 $Y=1.07 $X2=0 $Y2=0
cc_416 N_Y_c_641_n N_VGND_c_776_n 0.0170777f $X=4 $Y=1.07 $X2=0 $Y2=0
cc_417 N_Y_c_682_n N_VGND_c_777_n 0.0240821f $X=4.925 $Y=0.955 $X2=0 $Y2=0
cc_418 N_Y_c_704_n N_VGND_c_778_n 0.0170777f $X=5.84 $Y=0.955 $X2=0 $Y2=0
cc_419 N_Y_c_642_n N_VGND_c_780_n 0.0233388f $X=6.385 $Y=1.07 $X2=0 $Y2=0
cc_420 N_Y_c_753_p N_VGND_c_783_n 0.0151136f $X=1.435 $Y=0.42 $X2=0 $Y2=0
cc_421 N_Y_c_754_p N_VGND_c_785_n 0.0124525f $X=3.235 $Y=0.42 $X2=0 $Y2=0
cc_422 N_Y_c_681_n N_VGND_c_786_n 0.0153472f $X=4.095 $Y=0.42 $X2=0 $Y2=0
cc_423 N_Y_c_687_n N_VGND_c_787_n 0.0153472f $X=5.085 $Y=0.42 $X2=0 $Y2=0
cc_424 N_Y_c_757_p N_VGND_c_788_n 0.0124525f $X=5.945 $Y=0.42 $X2=0 $Y2=0
cc_425 N_Y_M1005_d N_VGND_c_793_n 0.00254326f $X=1.295 $Y=0.235 $X2=0 $Y2=0
cc_426 N_Y_M1017_d N_VGND_c_793_n 0.00376082f $X=2.235 $Y=0.235 $X2=0 $Y2=0
cc_427 N_Y_M1002_s N_VGND_c_793_n 0.00536646f $X=3.095 $Y=0.235 $X2=0 $Y2=0
cc_428 N_Y_M1015_s N_VGND_c_793_n 0.00380103f $X=3.955 $Y=0.235 $X2=0 $Y2=0
cc_429 N_Y_M1004_d N_VGND_c_793_n 0.00380103f $X=4.945 $Y=0.235 $X2=0 $Y2=0
cc_430 N_Y_M1010_d N_VGND_c_793_n 0.00536646f $X=5.805 $Y=0.235 $X2=0 $Y2=0
cc_431 N_Y_c_753_p N_VGND_c_793_n 0.0102248f $X=1.435 $Y=0.42 $X2=0 $Y2=0
cc_432 N_Y_c_651_n N_VGND_c_793_n 0.00965725f $X=2.21 $Y=0.93 $X2=0 $Y2=0
cc_433 N_Y_c_747_p N_VGND_c_793_n 0.00886411f $X=2.375 $Y=0.42 $X2=0 $Y2=0
cc_434 N_Y_c_754_p N_VGND_c_793_n 0.00730901f $X=3.235 $Y=0.42 $X2=0 $Y2=0
cc_435 N_Y_c_681_n N_VGND_c_793_n 0.00967594f $X=4.095 $Y=0.42 $X2=0 $Y2=0
cc_436 N_Y_c_687_n N_VGND_c_793_n 0.00967594f $X=5.085 $Y=0.42 $X2=0 $Y2=0
cc_437 N_Y_c_757_p N_VGND_c_793_n 0.00730901f $X=5.945 $Y=0.42 $X2=0 $Y2=0
cc_438 N_Y_c_643_n N_VGND_c_793_n 8.12449e-19 $X=2.375 $Y=0.93 $X2=0 $Y2=0
