* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfxbp_lp CLK D VGND VNB VPB VPWR Q Q_N
X0 a_1445_419# a_1507_321# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR a_1507_321# a_2062_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VGND a_1339_153# a_1742_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_2010_127# a_1507_321# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_455_85# a_615_93# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_1049_125# a_27_403# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_455_85# a_511_218# a_239_403# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 VPWR a_2062_367# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_1742_57# a_1339_153# a_1507_321# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_2168_127# a_1507_321# a_2062_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND D a_297_85# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_511_218# a_27_403# a_1049_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_2062_367# a_2436_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_349_323# a_615_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 a_349_323# a_27_403# a_455_85# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_2436_57# a_2062_367# Q_N VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1339_153# a_511_218# a_1445_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_1232_153# a_27_403# a_1339_153# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Q a_1507_321# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 a_27_403# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 VPWR a_1339_153# a_1507_321# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 Q a_1507_321# a_2010_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_763_119# a_455_85# a_615_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1339_153# a_511_218# a_615_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_125_85# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_27_403# CLK a_125_85# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_615_93# a_27_403# a_1339_153# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 VGND a_455_85# a_763_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_573_119# a_615_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VGND a_1507_321# a_2168_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VPWR D a_239_403# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X31 a_511_218# a_27_403# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 a_297_85# D a_239_403# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_239_403# a_27_403# a_455_85# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_455_85# a_511_218# a_573_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1232_153# a_1507_321# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
