* File: sky130_fd_sc_lp__or2_m.pxi.spice
* Created: Fri Aug 28 11:22:01 2020
* 
x_PM_SKY130_FD_SC_LP__OR2_M%B N_B_c_42_n N_B_c_43_n N_B_M1001_g N_B_c_49_n
+ N_B_M1004_g N_B_c_44_n N_B_c_45_n N_B_c_50_n B B N_B_c_47_n
+ PM_SKY130_FD_SC_LP__OR2_M%B
x_PM_SKY130_FD_SC_LP__OR2_M%A N_A_M1003_g N_A_M1002_g A N_A_c_84_n N_A_c_85_n
+ PM_SKY130_FD_SC_LP__OR2_M%A
x_PM_SKY130_FD_SC_LP__OR2_M%A_63_397# N_A_63_397#_M1001_d N_A_63_397#_M1004_s
+ N_A_63_397#_c_123_n N_A_63_397#_M1005_g N_A_63_397#_M1000_g
+ N_A_63_397#_c_125_n N_A_63_397#_c_119_n N_A_63_397#_c_120_n
+ N_A_63_397#_c_121_n N_A_63_397#_c_126_n N_A_63_397#_c_122_n
+ N_A_63_397#_c_128_n N_A_63_397#_c_129_n PM_SKY130_FD_SC_LP__OR2_M%A_63_397#
x_PM_SKY130_FD_SC_LP__OR2_M%VPWR N_VPWR_M1002_d N_VPWR_c_186_n VPWR
+ N_VPWR_c_187_n N_VPWR_c_188_n N_VPWR_c_185_n N_VPWR_c_190_n
+ PM_SKY130_FD_SC_LP__OR2_M%VPWR
x_PM_SKY130_FD_SC_LP__OR2_M%X N_X_M1005_d N_X_M1000_d X X X X X X X
+ PM_SKY130_FD_SC_LP__OR2_M%X
x_PM_SKY130_FD_SC_LP__OR2_M%VGND N_VGND_M1001_s N_VGND_M1003_d N_VGND_c_222_n
+ N_VGND_c_223_n N_VGND_c_224_n N_VGND_c_225_n VGND N_VGND_c_226_n
+ N_VGND_c_227_n N_VGND_c_228_n PM_SKY130_FD_SC_LP__OR2_M%VGND
cc_1 VNB N_B_c_42_n 0.0188576f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.725
cc_2 VNB N_B_c_43_n 0.0222812f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.765
cc_3 VNB N_B_c_44_n 0.0426915f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.84
cc_4 VNB N_B_c_45_n 0.0237561f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.435
cc_5 VNB B 0.00775901f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B_c_47_n 0.0369799f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.93
cc_7 VNB N_A_M1003_g 0.0378f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.765
cc_8 VNB N_A_M1002_g 0.0107867f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.195
cc_9 VNB N_A_c_84_n 0.0375039f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.84
cc_10 VNB N_A_c_85_n 0.00339651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_63_397#_M1005_g 0.0642298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_63_397#_c_119_n 0.00143385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_63_397#_c_120_n 0.00749167f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.93
cc_14 VNB N_A_63_397#_c_121_n 0.00345824f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.93
cc_15 VNB N_A_63_397#_c_122_n 0.00641091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_185_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.8
cc_17 VNB X 0.0490669f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.195
cc_18 VNB N_VGND_c_222_n 0.0142907f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.195
cc_19 VNB N_VGND_c_223_n 0.00441053f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.84
cc_20 VNB N_VGND_c_224_n 0.0181538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_225_n 0.00439692f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.435
cc_22 VNB N_VGND_c_226_n 0.0189732f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_VGND_c_227_n 0.131773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_228_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VPB N_B_c_42_n 0.00491218f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.725
cc_26 VPB N_B_c_49_n 0.0181974f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.875
cc_27 VPB N_B_c_50_n 0.0386439f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.8
cc_28 VPB N_A_M1002_g 0.0251169f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.195
cc_29 VPB N_A_63_397#_c_123_n 0.0422346f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.195
cc_30 VPB N_A_63_397#_M1005_g 0.0382546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_63_397#_c_125_n 0.0106479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_63_397#_c_126_n 0.00857164f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.93
cc_33 VPB N_A_63_397#_c_122_n 8.26908e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_63_397#_c_128_n 0.00615759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_63_397#_c_129_n 0.0517737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_186_n 0.018794f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.875
cc_37 VPB N_VPWR_c_187_n 0.0351191f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.915
cc_38 VPB N_VPWR_c_188_n 0.0194756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_185_n 0.0760514f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.8
cc_40 VPB N_VPWR_c_190_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_41 VPB X 0.0408935f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.195
cc_42 N_B_c_43_n N_A_M1003_g 0.0206232f $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_43 B N_A_M1003_g 0.00202482f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_44 N_B_c_47_n N_A_M1003_g 0.00396937f $X=0.27 $Y=0.93 $X2=0 $Y2=0
cc_45 N_B_c_42_n N_A_M1002_g 0.00443634f $X=0.36 $Y=1.725 $X2=0 $Y2=0
cc_46 N_B_c_50_n N_A_M1002_g 0.0522287f $X=0.655 $Y=1.8 $X2=0 $Y2=0
cc_47 N_B_c_50_n N_A_c_84_n 0.00196828f $X=0.655 $Y=1.8 $X2=0 $Y2=0
cc_48 B N_A_c_84_n 7.19452e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_49 N_B_c_47_n N_A_c_84_n 0.0169426f $X=0.27 $Y=0.93 $X2=0 $Y2=0
cc_50 N_B_c_44_n N_A_c_85_n 9.20069e-19 $X=0.585 $Y=0.84 $X2=0 $Y2=0
cc_51 N_B_c_50_n N_A_c_85_n 0.00156043f $X=0.655 $Y=1.8 $X2=0 $Y2=0
cc_52 B N_A_c_85_n 0.0103294f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_53 N_B_c_47_n N_A_c_85_n 0.00143887f $X=0.27 $Y=0.93 $X2=0 $Y2=0
cc_54 N_B_c_49_n N_A_63_397#_c_125_n 0.0162036f $X=0.655 $Y=1.875 $X2=0 $Y2=0
cc_55 N_B_c_43_n N_A_63_397#_c_119_n 0.0017418f $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_56 N_B_c_43_n N_A_63_397#_c_121_n 0.00300591f $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_57 B N_A_63_397#_c_121_n 0.00633017f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_B_c_49_n N_A_63_397#_c_128_n 0.0136228f $X=0.655 $Y=1.875 $X2=0 $Y2=0
cc_59 N_B_c_50_n N_A_63_397#_c_128_n 0.0307462f $X=0.655 $Y=1.8 $X2=0 $Y2=0
cc_60 B N_A_63_397#_c_128_n 9.70681e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_61 N_B_c_49_n N_A_63_397#_c_129_n 0.00636415f $X=0.655 $Y=1.875 $X2=0 $Y2=0
cc_62 N_B_c_49_n N_VPWR_c_185_n 9.23649e-19 $X=0.655 $Y=1.875 $X2=0 $Y2=0
cc_63 N_B_c_44_n N_VGND_c_222_n 0.00136711f $X=0.585 $Y=0.84 $X2=0 $Y2=0
cc_64 B N_VGND_c_222_n 0.0014801f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_65 N_B_c_43_n N_VGND_c_223_n 0.00328509f $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_66 N_B_c_44_n N_VGND_c_223_n 0.00534209f $X=0.585 $Y=0.84 $X2=0 $Y2=0
cc_67 B N_VGND_c_223_n 0.00589151f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_68 N_B_c_43_n N_VGND_c_224_n 0.00585385f $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_69 N_B_c_44_n N_VGND_c_224_n 5.38734e-19 $X=0.585 $Y=0.84 $X2=0 $Y2=0
cc_70 N_B_c_43_n N_VGND_c_227_n 0.0117471f $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_71 N_B_c_44_n N_VGND_c_227_n 0.0020757f $X=0.585 $Y=0.84 $X2=0 $Y2=0
cc_72 B N_VGND_c_227_n 0.00326316f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_A_63_397#_M1005_g 0.0738706f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_M1002_g N_A_63_397#_c_125_n 0.00432158f $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_A_63_397#_c_119_n 9.4709e-19 $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_A_63_397#_c_120_n 0.0142217f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_c_84_n N_A_63_397#_c_120_n 7.52443e-19 $X=0.86 $Y=1.32 $X2=0 $Y2=0
cc_78 N_A_c_85_n N_A_63_397#_c_120_n 0.00512801f $X=0.86 $Y=1.32 $X2=0 $Y2=0
cc_79 N_A_c_84_n N_A_63_397#_c_121_n 0.00474817f $X=0.86 $Y=1.32 $X2=0 $Y2=0
cc_80 N_A_c_85_n N_A_63_397#_c_121_n 0.0106208f $X=0.86 $Y=1.32 $X2=0 $Y2=0
cc_81 N_A_M1002_g N_A_63_397#_c_126_n 0.0148241f $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_82 N_A_M1003_g N_A_63_397#_c_122_n 0.0160141f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_c_85_n N_A_63_397#_c_122_n 0.0141363f $X=0.86 $Y=1.32 $X2=0 $Y2=0
cc_84 N_A_M1002_g N_A_63_397#_c_128_n 0.0100506f $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_85 N_A_c_84_n N_A_63_397#_c_128_n 0.00493599f $X=0.86 $Y=1.32 $X2=0 $Y2=0
cc_86 N_A_c_85_n N_A_63_397#_c_128_n 0.0176821f $X=0.86 $Y=1.32 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_A_63_397#_c_129_n 0.00965003f $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_88 N_A_M1002_g N_VPWR_c_186_n 9.84115e-19 $X=1.015 $Y=2.195 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VGND_c_224_n 0.00437852f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_M1003_g N_VGND_c_225_n 0.00156327f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_M1003_g N_VGND_c_227_n 0.00604796f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_63_397#_c_125_n A_146_397# 2.83863e-19 $X=0.78 $Y=2.94 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_63_397#_c_128_n A_146_397# 2.57373e-19 $X=0.945 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_63_397#_c_123_n N_VPWR_c_186_n 0.0182077f $X=1.37 $Y=2.85 $X2=0 $Y2=0
cc_95 N_A_63_397#_M1005_g N_VPWR_c_186_n 0.00666891f $X=1.445 $Y=0.445 $X2=0
+ $Y2=0
cc_96 N_A_63_397#_c_125_n N_VPWR_c_186_n 0.0496845f $X=0.78 $Y=2.94 $X2=0 $Y2=0
cc_97 N_A_63_397#_c_126_n N_VPWR_c_186_n 0.0157468f $X=1.205 $Y=1.83 $X2=0 $Y2=0
cc_98 N_A_63_397#_c_129_n N_VPWR_c_186_n 0.00508672f $X=0.78 $Y=2.85 $X2=0 $Y2=0
cc_99 N_A_63_397#_c_123_n N_VPWR_c_187_n 0.00445258f $X=1.37 $Y=2.85 $X2=0 $Y2=0
cc_100 N_A_63_397#_c_125_n N_VPWR_c_187_n 0.0167839f $X=0.78 $Y=2.94 $X2=0 $Y2=0
cc_101 N_A_63_397#_c_129_n N_VPWR_c_187_n 0.0059602f $X=0.78 $Y=2.85 $X2=0 $Y2=0
cc_102 N_A_63_397#_c_123_n N_VPWR_c_188_n 0.00550617f $X=1.37 $Y=2.85 $X2=0
+ $Y2=0
cc_103 N_A_63_397#_c_123_n N_VPWR_c_185_n 0.0106337f $X=1.37 $Y=2.85 $X2=0 $Y2=0
cc_104 N_A_63_397#_c_125_n N_VPWR_c_185_n 0.0108843f $X=0.78 $Y=2.94 $X2=0 $Y2=0
cc_105 N_A_63_397#_c_129_n N_VPWR_c_185_n 0.00806414f $X=0.78 $Y=2.85 $X2=0
+ $Y2=0
cc_106 N_A_63_397#_M1005_g X 0.0440414f $X=1.445 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_63_397#_c_119_n X 0.00204746f $X=0.8 $Y=0.51 $X2=0 $Y2=0
cc_108 N_A_63_397#_c_120_n X 0.0132066f $X=1.205 $Y=0.81 $X2=0 $Y2=0
cc_109 N_A_63_397#_c_126_n X 0.0132066f $X=1.205 $Y=1.83 $X2=0 $Y2=0
cc_110 N_A_63_397#_c_122_n X 0.0591676f $X=1.29 $Y=1.745 $X2=0 $Y2=0
cc_111 N_A_63_397#_c_128_n X 0.00366318f $X=0.945 $Y=2.02 $X2=0 $Y2=0
cc_112 N_A_63_397#_c_119_n N_VGND_c_224_n 0.008231f $X=0.8 $Y=0.51 $X2=0 $Y2=0
cc_113 N_A_63_397#_c_120_n N_VGND_c_224_n 0.00305343f $X=1.205 $Y=0.81 $X2=0
+ $Y2=0
cc_114 N_A_63_397#_M1005_g N_VGND_c_225_n 0.00288714f $X=1.445 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A_63_397#_c_120_n N_VGND_c_225_n 0.0149698f $X=1.205 $Y=0.81 $X2=0
+ $Y2=0
cc_116 N_A_63_397#_M1005_g N_VGND_c_226_n 0.00580462f $X=1.445 $Y=0.445 $X2=0
+ $Y2=0
cc_117 N_A_63_397#_c_120_n N_VGND_c_226_n 6.60115e-19 $X=1.205 $Y=0.81 $X2=0
+ $Y2=0
cc_118 N_A_63_397#_M1001_d N_VGND_c_227_n 0.00373063f $X=0.66 $Y=0.235 $X2=0
+ $Y2=0
cc_119 N_A_63_397#_M1005_g N_VGND_c_227_n 0.0115436f $X=1.445 $Y=0.445 $X2=0
+ $Y2=0
cc_120 N_A_63_397#_c_119_n N_VGND_c_227_n 0.00765087f $X=0.8 $Y=0.51 $X2=0 $Y2=0
cc_121 N_A_63_397#_c_120_n N_VGND_c_227_n 0.00702325f $X=1.205 $Y=0.81 $X2=0
+ $Y2=0
cc_122 N_VPWR_c_186_n X 0.0291033f $X=1.23 $Y=2.26 $X2=0 $Y2=0
cc_123 N_VPWR_c_188_n X 0.00623633f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_124 N_VPWR_c_185_n X 0.00710559f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_125 X N_VGND_c_226_n 0.00877924f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_126 N_X_M1005_d N_VGND_c_227_n 0.0042053f $X=1.52 $Y=0.235 $X2=0 $Y2=0
cc_127 X N_VGND_c_227_n 0.00770513f $X=1.595 $Y=0.47 $X2=0 $Y2=0
