* File: sky130_fd_sc_lp__xor2_2.pex.spice
* Created: Wed Sep  2 10:41:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR2_2%A 3 6 10 14 18 22 25 29 32 33 34 36 38 40 41
+ 42 45 52 53 55 59 60 62 63 68 74 75 78 83
c222 75 0 1.62796e-19 $X=2.35 $Y=1.51
c223 38 0 5.5472e-20 $X=3.83 $Y=1.355
c224 14 0 1.57015e-19 $X=2.35 $Y=0.745
r225 73 75 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.17 $Y=1.51
+ $X2=2.35 $Y2=1.51
r226 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.51 $X2=2.17 $Y2=1.51
r227 70 73 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.05 $Y=1.51
+ $X2=2.17 $Y2=1.51
r228 63 74 0.154333 $w=7.73e-07 $l=1e-08 $layer=LI1_cond $X=2.16 $Y=1.732
+ $X2=2.17 $Y2=1.732
r229 62 63 7.40797 $w=7.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.732
+ $X2=2.16 $Y2=1.732
r230 59 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.905 $Y=1.44
+ $X2=3.905 $Y2=1.605
r231 59 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.905 $Y=1.44
+ $X2=3.905 $Y2=1.275
r232 58 60 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.83 $Y=1.48
+ $X2=3.985 $Y2=1.48
r233 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.905
+ $Y=1.44 $X2=3.905 $Y2=1.44
r234 55 62 26.8611 $w=3.38e-07 $l=7.5e-07 $layer=LI1_cond $X=0.845 $Y=2.035
+ $X2=1.595 $Y2=2.035
r235 52 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.44
+ $X2=0.58 $Y2=1.605
r236 52 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.44
+ $X2=0.58 $Y2=1.275
r237 51 53 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.58 $Y=1.475
+ $X2=0.76 $Y2=1.475
r238 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.58
+ $Y=1.44 $X2=0.58 $Y2=1.44
r239 48 51 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.455 $Y=1.475
+ $X2=0.58 $Y2=1.475
r240 46 83 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.56 $Y=1.51
+ $X2=5.675 $Y2=1.51
r241 46 80 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.56 $Y=1.51 $X2=5.47
+ $Y2=1.51
r242 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.56
+ $Y=1.51 $X2=5.56 $Y2=1.51
r243 43 45 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.56 $Y=1.92
+ $X2=5.56 $Y2=1.51
r244 41 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.395 $Y=2.005
+ $X2=5.56 $Y2=1.92
r245 41 42 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=5.395 $Y=2.005
+ $X2=4.07 $Y2=2.005
r246 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.985 $Y=1.92
+ $X2=4.07 $Y2=2.005
r247 39 60 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.985 $Y=1.605
+ $X2=3.985 $Y2=1.48
r248 39 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.985 $Y=1.605
+ $X2=3.985 $Y2=1.92
r249 38 58 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.83 $Y=1.355
+ $X2=3.83 $Y2=1.48
r250 37 38 35.1212 $w=1.78e-07 $l=5.7e-07 $layer=LI1_cond $X=3.83 $Y=0.785
+ $X2=3.83 $Y2=1.355
r251 36 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=1.95
+ $X2=0.845 $Y2=2.035
r252 35 53 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.76 $Y=1.605
+ $X2=0.76 $Y2=1.475
r253 35 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.76 $Y=1.605
+ $X2=0.76 $Y2=1.95
r254 33 37 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.74 $Y=0.7
+ $X2=3.83 $Y2=0.785
r255 33 34 208.77 $w=1.68e-07 $l=3.2e-06 $layer=LI1_cond $X=3.74 $Y=0.7 $X2=0.54
+ $Y2=0.7
r256 32 48 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.455 $Y=1.345
+ $X2=0.455 $Y2=1.475
r257 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.455 $Y=0.785
+ $X2=0.54 $Y2=0.7
r258 31 32 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.455 $Y=0.785
+ $X2=0.455 $Y2=1.345
r259 27 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.675 $Y=1.345
+ $X2=5.675 $Y2=1.51
r260 27 29 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.675 $Y=1.345
+ $X2=5.675 $Y2=0.745
r261 23 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.675
+ $X2=5.47 $Y2=1.51
r262 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.47 $Y=1.675
+ $X2=5.47 $Y2=2.465
r263 22 78 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.995 $Y=0.745
+ $X2=3.995 $Y2=1.275
r264 18 79 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.86 $Y=2.465
+ $X2=3.86 $Y2=1.605
r265 12 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.345
+ $X2=2.35 $Y2=1.51
r266 12 14 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.35 $Y=1.345 $X2=2.35
+ $Y2=0.745
r267 8 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.675
+ $X2=2.05 $Y2=1.51
r268 8 10 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.05 $Y=1.675
+ $X2=2.05 $Y2=2.465
r269 6 69 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.67 $Y=2.465
+ $X2=0.67 $Y2=1.605
r270 3 68 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.67 $Y=0.745
+ $X2=0.67 $Y2=1.275
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%B 3 7 11 15 19 23 27 31 33 34 39 45 47 54 55
c143 55 0 5.5472e-20 $X=4.88 $Y=1.51
c144 45 0 1.62796e-19 $X=1.33 $Y=1.51
r145 54 63 2.76705 $w=6.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.62 $Y=1.51
+ $X2=4.62 $Y2=1.665
r146 53 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.79 $Y=1.51 $X2=4.88
+ $Y2=1.51
r147 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.79
+ $Y=1.51 $X2=4.79 $Y2=1.51
r148 51 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.45 $Y=1.51
+ $X2=4.79 $Y2=1.51
r149 49 51 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=4.425 $Y=1.51
+ $X2=4.45 $Y2=1.51
r150 46 47 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.53 $Y=1.51
+ $X2=1.69 $Y2=1.51
r151 44 46 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.33 $Y=1.51 $X2=1.53
+ $Y2=1.51
r152 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.33
+ $Y=1.51 $X2=1.33 $Y2=1.51
r153 41 44 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.1 $Y=1.51
+ $X2=1.33 $Y2=1.51
r154 39 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.665
r155 36 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r156 34 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r157 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=1.665
+ $X2=4.56 $Y2=1.665
r158 33 34 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=4.415 $Y=1.665
+ $X2=1.345 $Y2=1.665
r159 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.675
+ $X2=4.88 $Y2=1.51
r160 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.88 $Y=1.675
+ $X2=4.88 $Y2=2.465
r161 25 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.345
+ $X2=4.88 $Y2=1.51
r162 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.88 $Y=1.345 $X2=4.88
+ $Y2=0.745
r163 21 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.45 $Y=1.675
+ $X2=4.45 $Y2=1.51
r164 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.45 $Y=1.675
+ $X2=4.45 $Y2=2.465
r165 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.345
+ $X2=4.425 $Y2=1.51
r166 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.425 $Y=1.345
+ $X2=4.425 $Y2=0.745
r167 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.345
+ $X2=1.69 $Y2=1.51
r168 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.69 $Y=1.345 $X2=1.69
+ $Y2=0.745
r169 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.53 $Y=1.675
+ $X2=1.53 $Y2=1.51
r170 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.53 $Y=1.675
+ $X2=1.53 $Y2=2.465
r171 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.675
+ $X2=1.1 $Y2=1.51
r172 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.1 $Y=1.675 $X2=1.1
+ $Y2=2.465
r173 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.345
+ $X2=1.1 $Y2=1.51
r174 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.1 $Y=1.345 $X2=1.1
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%A_149_65# 1 2 3 10 12 15 17 19 22 24 30 33 35
+ 36 44 52
r115 51 52 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.405 $Y=1.44
+ $X2=3.43 $Y2=1.44
r116 50 51 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=3 $Y=1.44
+ $X2=3.405 $Y2=1.44
r117 49 50 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.975 $Y=1.44 $X2=3
+ $Y2=1.44
r118 45 49 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.865 $Y=1.44
+ $X2=2.975 $Y2=1.44
r119 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.44 $X2=2.865 $Y2=1.44
r120 36 39 4.32166 $w=2.38e-07 $l=9e-08 $layer=LI1_cond $X=1.31 $Y=2.375
+ $X2=1.31 $Y2=2.465
r121 34 35 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.615 $Y=1.605
+ $X2=2.615 $Y2=2.29
r122 33 44 10.4768 $w=2.73e-07 $l=2.5e-07 $layer=LI1_cond $X=2.615 $Y=1.467
+ $X2=2.865 $Y2=1.467
r123 33 34 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2.615 $Y=1.467
+ $X2=2.615 $Y2=1.605
r124 32 33 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.615 $Y=1.175
+ $X2=2.615 $Y2=1.33
r125 31 36 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.43 $Y=2.375
+ $X2=1.31 $Y2=2.375
r126 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.53 $Y=2.375
+ $X2=2.615 $Y2=2.29
r127 30 31 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.53 $Y=2.375
+ $X2=1.43 $Y2=2.375
r128 26 29 59.4556 $w=2.18e-07 $l=1.135e-06 $layer=LI1_cond $X=0.885 $Y=1.065
+ $X2=2.02 $Y2=1.065
r129 24 32 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.53 $Y=1.065
+ $X2=2.615 $Y2=1.175
r130 24 29 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=2.53 $Y=1.065
+ $X2=2.02 $Y2=1.065
r131 20 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.605
+ $X2=3.43 $Y2=1.44
r132 20 22 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.43 $Y=1.605
+ $X2=3.43 $Y2=2.465
r133 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.405 $Y=1.275
+ $X2=3.405 $Y2=1.44
r134 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.405 $Y=1.275
+ $X2=3.405 $Y2=0.745
r135 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3 $Y=1.605 $X2=3
+ $Y2=1.44
r136 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3 $Y=1.605 $X2=3
+ $Y2=2.465
r137 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.275
+ $X2=2.975 $Y2=1.44
r138 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.975 $Y=1.275
+ $X2=2.975 $Y2=0.745
r139 3 39 600 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.835 $X2=1.315 $Y2=2.465
r140 2 29 182 $w=1.7e-07 $l=8.32797e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.325 $X2=2.02 $Y2=1.04
r141 1 26 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=0.745
+ $Y=0.325 $X2=0.885 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%VPWR 1 2 3 4 15 18 21 23 26 28 30 35 45 46 52
+ 55 62
r85 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 62 65 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.175 $Y=3.025
+ $X2=5.175 $Y2=3.33
r87 59 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r88 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 55 58 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.155 $Y=3.025
+ $X2=4.155 $Y2=3.33
r90 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r91 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 46 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r93 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r94 43 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.34 $Y=3.33
+ $X2=5.175 $Y2=3.33
r95 43 45 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.34 $Y=3.33 $X2=6
+ $Y2=3.33
r96 42 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r98 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r100 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 36 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=3.33
+ $X2=2.265 $Y2=3.33
r102 36 38 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.43 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 35 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=4.155 $Y2=3.33
r104 35 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 34 53 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 34 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r107 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 31 49 4.79039 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.31 $Y2=3.33
r109 31 33 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.62 $Y=3.33 $X2=0.72
+ $Y2=3.33
r110 30 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=3.33
+ $X2=2.265 $Y2=3.33
r111 30 33 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.1 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 26 27 6.36223 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.437 $Y=2.455
+ $X2=0.437 $Y2=2.29
r115 24 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.155 $Y2=3.33
r116 23 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=5.175 $Y2=3.33
r117 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=4.32 $Y2=3.33
r118 19 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=3.245
+ $X2=2.265 $Y2=3.33
r119 19 21 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.265 $Y=3.245
+ $X2=2.265 $Y2=2.755
r120 18 49 3.27601 $w=3.65e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.437 $Y=3.245
+ $X2=0.31 $Y2=3.33
r121 17 26 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=0.437 $Y=2.472
+ $X2=0.437 $Y2=2.455
r122 17 18 24.4065 $w=3.63e-07 $l=7.73e-07 $layer=LI1_cond $X=0.437 $Y=2.472
+ $X2=0.437 $Y2=3.245
r123 15 27 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.38 $Y=1.985
+ $X2=0.38 $Y2=2.29
r124 4 62 600 $w=1.7e-07 $l=1.29534e-06 $layer=licon1_PDIFF $count=1 $X=4.955
+ $Y=1.835 $X2=5.175 $Y2=3.025
r125 3 55 600 $w=1.7e-07 $l=1.29534e-06 $layer=licon1_PDIFF $count=1 $X=3.935
+ $Y=1.835 $X2=4.155 $Y2=3.025
r126 2 21 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.835 $X2=2.265 $Y2=2.755
r127 1 26 300 $w=1.7e-07 $l=6.95414e-07 $layer=licon1_PDIFF $count=2 $X=0.295
+ $Y=1.835 $X2=0.455 $Y2=2.455
r128 1 15 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=0.295
+ $Y=1.835 $X2=0.42 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%A_149_367# 1 2 7 9 11 16
r23 16 18 6.3559 $w=3.28e-07 $l=1.82e-07 $layer=LI1_cond $X=1.765 $Y=2.755
+ $X2=1.765 $Y2=2.937
r24 12 14 3.14294 $w=2.75e-07 $l=1.15e-07 $layer=LI1_cond $X=1.02 $Y=2.937
+ $X2=0.905 $Y2=2.937
r25 11 18 1.82517 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=1.6 $Y=2.937
+ $X2=1.765 $Y2=2.937
r26 11 12 24.3061 $w=2.73e-07 $l=5.8e-07 $layer=LI1_cond $X=1.6 $Y=2.937
+ $X2=1.02 $Y2=2.937
r27 7 14 3.74419 $w=2.3e-07 $l=1.37e-07 $layer=LI1_cond $X=0.905 $Y=2.8
+ $X2=0.905 $Y2=2.937
r28 7 9 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.905 $Y=2.8
+ $X2=0.905 $Y2=2.455
r29 2 16 600 $w=1.7e-07 $l=9.96795e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.835 $X2=1.765 $Y2=2.755
r30 1 14 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.745
+ $Y=1.835 $X2=0.885 $Y2=2.91
r31 1 9 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=0.745
+ $Y=1.835 $X2=0.885 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%A_532_367# 1 2 3 4 13 14 19 25
r42 24 25 9.3668 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=2.837
+ $X2=3.81 $Y2=2.837
r43 17 19 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.665 $Y=2.685
+ $X2=5.685 $Y2=2.685
r44 17 25 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.665 $Y=2.685
+ $X2=3.81 $Y2=2.685
r45 14 22 10.7103 $w=4.75e-07 $l=4.17e-07 $layer=LI1_cond $X=3.202 $Y=2.837
+ $X2=2.785 $Y2=2.837
r46 13 24 1.813 $w=4.73e-07 $l=7.2e-08 $layer=LI1_cond $X=3.573 $Y=2.837
+ $X2=3.645 $Y2=2.837
r47 13 14 9.342 $w=4.73e-07 $l=3.71e-07 $layer=LI1_cond $X=3.573 $Y=2.837
+ $X2=3.202 $Y2=2.837
r48 4 19 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=5.545
+ $Y=1.835 $X2=5.685 $Y2=2.685
r49 3 17 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=1.835 $X2=4.665 $Y2=2.685
r50 2 24 600 $w=1.7e-07 $l=1.0176e-06 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.835 $X2=3.645 $Y2=2.785
r51 1 22 600 $w=1.7e-07 $l=1.02059e-06 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.835 $X2=2.785 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%X 1 2 3 11 13 16 17 18 23 25 27 29 30 31 38
+ 40
c94 23 0 1.57015e-19 $X=3.295 $Y=1.057
r95 38 40 2.21624 $w=2.58e-07 $l=5e-08 $layer=LI1_cond $X=6.025 $Y=1.245
+ $X2=6.025 $Y2=1.295
r96 30 31 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=6.025 $Y=1.665
+ $X2=6.025 $Y2=2.035
r97 29 38 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=1.16
+ $X2=6.025 $Y2=1.245
r98 29 30 15.6466 $w=2.58e-07 $l=3.53e-07 $layer=LI1_cond $X=6.025 $Y=1.312
+ $X2=6.025 $Y2=1.665
r99 29 40 0.75352 $w=2.58e-07 $l=1.7e-08 $layer=LI1_cond $X=6.025 $Y=1.312
+ $X2=6.025 $Y2=1.295
r100 27 51 5.27022 $w=5.44e-07 $l=2.35e-07 $layer=LI1_cond $X=4.8 $Y=0.925
+ $X2=4.8 $Y2=1.16
r101 27 47 5.49449 $w=5.44e-07 $l=2.45e-07 $layer=LI1_cond $X=4.8 $Y=0.925
+ $X2=4.8 $Y2=0.68
r102 26 31 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=6.025 $Y=2.26
+ $X2=6.025 $Y2=2.035
r103 21 23 5.68071 $w=2.03e-07 $l=1.05e-07 $layer=LI1_cond $X=3.19 $Y=1.057
+ $X2=3.295 $Y2=1.057
r104 19 51 7.68949 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=5.125 $Y=1.16
+ $X2=4.8 $Y2=1.16
r105 18 29 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.895 $Y=1.16
+ $X2=6.025 $Y2=1.16
r106 18 19 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.895 $Y=1.16
+ $X2=5.125 $Y2=1.16
r107 16 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.895 $Y=2.345
+ $X2=6.025 $Y2=2.26
r108 16 17 164.08 $w=1.68e-07 $l=2.515e-06 $layer=LI1_cond $X=5.895 $Y=2.345
+ $X2=3.38 $Y2=2.345
r109 14 23 1.83547 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=3.295 $Y=1.16
+ $X2=3.295 $Y2=1.057
r110 14 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.295 $Y=1.16
+ $X2=3.295 $Y2=1.84
r111 13 25 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=2.005
+ $X2=3.215 $Y2=1.84
r112 11 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.215 $Y=2.26
+ $X2=3.38 $Y2=2.345
r113 11 13 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.215 $Y=2.26
+ $X2=3.215 $Y2=2.005
r114 3 13 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=3.075
+ $Y=1.835 $X2=3.215 $Y2=2.005
r115 2 47 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=4.5
+ $Y=0.325 $X2=4.64 $Y2=0.68
r116 1 21 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=3.05
+ $Y=0.325 $X2=3.19 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%VGND 1 2 3 4 5 16 18 22 26 28 32 34 36 39 40
+ 41 47 51 63 66 70
r73 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r74 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r75 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r76 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r77 58 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r78 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r79 55 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r80 55 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r81 54 57 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r82 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r83 52 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=0 $X2=3.7
+ $Y2=0
r84 52 54 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.865 $Y=0 $X2=4.08
+ $Y2=0
r85 51 69 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=6.017
+ $Y2=0
r86 51 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.52
+ $Y2=0
r87 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r88 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r89 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.645
+ $Y2=0
r90 47 49 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.16
+ $Y2=0
r91 46 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r92 46 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r93 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r94 43 60 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.262
+ $Y2=0
r95 43 45 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=1.2
+ $Y2=0
r96 41 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r97 41 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r98 39 45 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.23 $Y=0 $X2=1.2
+ $Y2=0
r99 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=0 $X2=1.395
+ $Y2=0
r100 38 49 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=2.16
+ $Y2=0
r101 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.395
+ $Y2=0
r102 34 69 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=6.017 $Y2=0
r103 34 36 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=5.96 $Y2=0.47
r104 30 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085 $X2=3.7
+ $Y2=0
r105 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.36
r106 29 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.645
+ $Y2=0
r107 28 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.7
+ $Y2=0
r108 28 29 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.535 $Y=0
+ $X2=2.81 $Y2=0
r109 24 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0
r110 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0.36
r111 20 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0
r112 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0.36
r113 16 60 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.262 $Y2=0
r114 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.36 $Y2=0.36
r115 5 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.75
+ $Y=0.325 $X2=5.96 $Y2=0.47
r116 4 32 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=3.48
+ $Y=0.325 $X2=3.7 $Y2=0.36
r117 3 26 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.325 $X2=2.645 $Y2=0.36
r118 2 22 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.325 $X2=1.395 $Y2=0.36
r119 1 18 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.195 $X2=0.36 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_2%A_814_65# 1 2 9 11 12 13
r30 13 15 3.17341 $w=5.19e-07 $l=1.35e-07 $layer=LI1_cond $X=5.3 $Y=0.34 $X2=5.3
+ $Y2=0.475
r31 11 13 7.39147 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=5.3 $Y2=0.34
r32 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=4.305 $Y2=0.34
r33 7 12 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=4.197 $Y=0.425
+ $X2=4.305 $Y2=0.34
r34 7 9 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=4.197 $Y=0.425
+ $X2=4.197 $Y2=0.45
r35 2 15 60.6667 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_NDIFF $count=3 $X=4.955
+ $Y=0.325 $X2=5.46 $Y2=0.475
r36 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.07
+ $Y=0.325 $X2=4.21 $Y2=0.45
.ends

