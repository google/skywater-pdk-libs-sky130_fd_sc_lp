* File: sky130_fd_sc_lp__or2b_lp.pxi.spice
* Created: Fri Aug 28 11:22:42 2020
* 
x_PM_SKY130_FD_SC_LP__OR2B_LP%B_N N_B_N_M1006_g N_B_N_M1011_g N_B_N_M1002_g
+ N_B_N_c_71_n N_B_N_c_72_n B_N B_N N_B_N_c_74_n PM_SKY130_FD_SC_LP__OR2B_LP%B_N
x_PM_SKY130_FD_SC_LP__OR2B_LP%A_30_57# N_A_30_57#_M1006_s N_A_30_57#_M1011_s
+ N_A_30_57#_c_106_n N_A_30_57#_M1007_g N_A_30_57#_c_107_n N_A_30_57#_M1008_g
+ N_A_30_57#_M1005_g N_A_30_57#_c_109_n N_A_30_57#_c_110_n N_A_30_57#_c_111_n
+ N_A_30_57#_c_112_n N_A_30_57#_c_113_n N_A_30_57#_c_114_n
+ PM_SKY130_FD_SC_LP__OR2B_LP%A_30_57#
x_PM_SKY130_FD_SC_LP__OR2B_LP%A N_A_c_171_n N_A_M1001_g N_A_c_172_n N_A_c_173_n
+ N_A_M1010_g N_A_c_174_n N_A_M1009_g N_A_c_175_n N_A_c_176_n N_A_c_182_n
+ N_A_c_177_n A A A A N_A_c_178_n N_A_c_179_n PM_SKY130_FD_SC_LP__OR2B_LP%A
x_PM_SKY130_FD_SC_LP__OR2B_LP%A_290_409# N_A_290_409#_M1008_d
+ N_A_290_409#_M1005_s N_A_290_409#_M1003_g N_A_290_409#_M1000_g
+ N_A_290_409#_M1004_g N_A_290_409#_c_237_n N_A_290_409#_c_238_n
+ N_A_290_409#_c_247_n N_A_290_409#_c_239_n N_A_290_409#_c_240_n
+ N_A_290_409#_c_248_n N_A_290_409#_c_241_n N_A_290_409#_c_242_n
+ N_A_290_409#_c_243_n N_A_290_409#_c_244_n
+ PM_SKY130_FD_SC_LP__OR2B_LP%A_290_409#
x_PM_SKY130_FD_SC_LP__OR2B_LP%VPWR N_VPWR_M1011_d N_VPWR_M1010_d N_VPWR_c_322_n
+ N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n VPWR N_VPWR_c_326_n
+ N_VPWR_c_321_n N_VPWR_c_328_n PM_SKY130_FD_SC_LP__OR2B_LP%VPWR
x_PM_SKY130_FD_SC_LP__OR2B_LP%X N_X_M1004_d N_X_M1000_d X X X X X X X X
+ PM_SKY130_FD_SC_LP__OR2B_LP%X
x_PM_SKY130_FD_SC_LP__OR2B_LP%VGND N_VGND_M1002_d N_VGND_M1009_d N_VGND_c_377_n
+ N_VGND_c_378_n VGND N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n
+ N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n PM_SKY130_FD_SC_LP__OR2B_LP%VGND
cc_1 VNB N_B_N_M1006_g 0.0387204f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.495
cc_2 VNB N_B_N_M1002_g 0.0310648f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=0.495
cc_3 VNB N_B_N_c_71_n 0.0173685f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.325
cc_4 VNB N_B_N_c_72_n 0.00461971f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.845
cc_5 VNB B_N 2.87194e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_B_N_c_74_n 0.0308344f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.34
cc_7 VNB N_A_30_57#_c_106_n 0.0164502f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.545
cc_8 VNB N_A_30_57#_c_107_n 0.0160666f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=0.495
cc_9 VNB N_A_30_57#_M1005_g 0.0115644f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.325
cc_10 VNB N_A_30_57#_c_109_n 0.0240181f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_11 VNB N_A_30_57#_c_110_n 0.0335117f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.34
cc_12 VNB N_A_30_57#_c_111_n 0.0157643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_30_57#_c_112_n 0.00994965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_30_57#_c_113_n 0.0125723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_30_57#_c_114_n 0.0951568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_c_171_n 0.0137713f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.175
cc_17 VNB N_A_c_172_n 0.00751286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_c_173_n 0.00859552f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.845
cc_19 VNB N_A_c_174_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=0.495
cc_20 VNB N_A_c_175_n 0.0169794f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.618
cc_21 VNB N_A_c_176_n 0.0189696f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.845
cc_22 VNB N_A_c_177_n 0.00492764f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_23 VNB N_A_c_178_n 0.0143196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_179_n 0.00509927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_290_409#_M1003_g 0.0184847f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.175
cc_26 VNB N_A_290_409#_M1004_g 0.0229371f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.845
cc_27 VNB N_A_290_409#_c_237_n 0.0232427f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.34
cc_28 VNB N_A_290_409#_c_238_n 0.0318468f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.295
cc_29 VNB N_A_290_409#_c_239_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_290_409#_c_240_n 0.0147354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_290_409#_c_241_n 0.00875615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_290_409#_c_242_n 0.00424321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_290_409#_c_243_n 0.00425815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_290_409#_c_244_n 0.0276599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_321_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB X 0.0694043f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.545
cc_37 VNB N_VGND_c_377_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.175
cc_38 VNB N_VGND_c_378_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.325
cc_39 VNB N_VGND_c_379_n 0.0276759f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.845
cc_40 VNB N_VGND_c_380_n 0.0357921f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.34
cc_41 VNB N_VGND_c_381_n 0.0292623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_382_n 0.237872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_383_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_384_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_B_N_M1011_g 0.0391252f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_46 VPB N_B_N_c_72_n 0.0295448f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.845
cc_47 VPB B_N 0.00194915f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_48 VPB N_A_30_57#_M1005_g 0.0466264f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.325
cc_49 VPB N_A_30_57#_c_110_n 0.0601925f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.34
cc_50 VPB N_A_M1010_g 0.0263386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_c_176_n 0.00469138f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.845
cc_52 VPB N_A_c_182_n 0.0143495f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_53 VPB N_A_c_179_n 0.00451746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_290_409#_M1000_g 0.0483082f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.325
cc_55 VPB N_A_290_409#_c_238_n 3.76079e-19 $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.295
cc_56 VPB N_A_290_409#_c_247_n 0.0143204f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.665
cc_57 VPB N_A_290_409#_c_248_n 0.00702064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_290_409#_c_241_n 0.0126765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_322_n 0.0238024f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=0.495
cc_60 VPB N_VPWR_c_323_n 0.0108039f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.845
cc_61 VPB N_VPWR_c_324_n 0.0481455f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.34
cc_62 VPB N_VPWR_c_325_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.34
cc_63 VPB N_VPWR_c_326_n 0.0219546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_321_n 0.0864302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_328_n 0.0256278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB X 0.0217749f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_67 VPB X 0.0389141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB X 0.0123879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 N_B_N_M1002_g N_A_30_57#_c_106_n 0.0147173f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_70 N_B_N_M1006_g N_A_30_57#_c_109_n 0.01276f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_71 N_B_N_M1002_g N_A_30_57#_c_109_n 0.00193397f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_72 N_B_N_M1006_g N_A_30_57#_c_110_n 0.0347577f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_73 B_N N_A_30_57#_c_110_n 0.0496126f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B_N_M1006_g N_A_30_57#_c_111_n 0.0111106f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_75 N_B_N_M1002_g N_A_30_57#_c_111_n 0.0123667f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_76 N_B_N_c_71_n N_A_30_57#_c_111_n 2.06304e-19 $X=0.69 $Y=1.325 $X2=0 $Y2=0
cc_77 B_N N_A_30_57#_c_111_n 0.0246251f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_78 N_B_N_M1006_g N_A_30_57#_c_112_n 0.00513266f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_79 N_B_N_M1002_g N_A_30_57#_c_113_n 0.00177929f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_80 B_N N_A_30_57#_c_113_n 0.0154308f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_81 N_B_N_c_74_n N_A_30_57#_c_113_n 7.10774e-19 $X=0.725 $Y=1.34 $X2=0 $Y2=0
cc_82 N_B_N_M1002_g N_A_30_57#_c_114_n 0.0283808f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_83 B_N N_A_30_57#_c_114_n 0.0013408f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B_N_c_74_n N_A_30_57#_c_114_n 0.00739135f $X=0.725 $Y=1.34 $X2=0 $Y2=0
cc_85 N_B_N_M1011_g N_VPWR_c_322_n 0.0231779f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_86 N_B_N_c_71_n N_VPWR_c_322_n 0.00154385f $X=0.69 $Y=1.325 $X2=0 $Y2=0
cc_87 N_B_N_c_72_n N_VPWR_c_322_n 0.00158413f $X=0.662 $Y=1.845 $X2=0 $Y2=0
cc_88 B_N N_VPWR_c_322_n 0.0193328f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B_N_M1011_g N_VPWR_c_321_n 0.0149833f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_90 N_B_N_M1011_g N_VPWR_c_328_n 0.00802402f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_91 N_B_N_M1006_g N_VGND_c_377_n 0.00189426f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_92 N_B_N_M1002_g N_VGND_c_377_n 0.0106455f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_93 N_B_N_M1006_g N_VGND_c_379_n 0.00502664f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_94 N_B_N_M1002_g N_VGND_c_379_n 0.00445056f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_95 N_B_N_M1006_g N_VGND_c_382_n 0.00628724f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_96 N_B_N_M1002_g N_VGND_c_382_n 0.0041956f $X=0.87 $Y=0.495 $X2=0 $Y2=0
cc_97 N_A_30_57#_c_107_n N_A_c_171_n 0.00898345f $X=1.69 $Y=0.825 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_30_57#_c_114_n N_A_c_173_n 0.00898345f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_30_57#_c_114_n N_A_c_175_n 0.00351518f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_30_57#_M1005_g N_A_c_182_n 0.0479845f $X=1.86 $Y=2.545 $X2=0 $Y2=0
cc_101 N_A_30_57#_c_114_n N_A_c_178_n 0.0508993f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_30_57#_c_114_n N_A_c_179_n 0.0126671f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_30_57#_M1005_g N_A_290_409#_c_247_n 0.0192487f $X=1.86 $Y=2.545 $X2=0
+ $Y2=0
cc_104 N_A_30_57#_c_106_n N_A_290_409#_c_239_n 0.00212449f $X=1.3 $Y=0.825 $X2=0
+ $Y2=0
cc_105 N_A_30_57#_c_107_n N_A_290_409#_c_239_n 0.0134923f $X=1.69 $Y=0.825 $X2=0
+ $Y2=0
cc_106 N_A_30_57#_c_113_n N_A_290_409#_c_239_n 0.00304084f $X=1.35 $Y=0.99 $X2=0
+ $Y2=0
cc_107 N_A_30_57#_c_114_n N_A_290_409#_c_239_n 0.00128561f $X=1.69 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_30_57#_M1005_g N_A_290_409#_c_248_n 0.00472934f $X=1.86 $Y=2.545
+ $X2=0 $Y2=0
cc_109 N_A_30_57#_c_113_n N_A_290_409#_c_248_n 0.00313051f $X=1.35 $Y=0.99 $X2=0
+ $Y2=0
cc_110 N_A_30_57#_c_114_n N_A_290_409#_c_248_n 0.00655008f $X=1.69 $Y=1.16 $X2=0
+ $Y2=0
cc_111 N_A_30_57#_M1005_g N_A_290_409#_c_241_n 0.0184058f $X=1.86 $Y=2.545 $X2=0
+ $Y2=0
cc_112 N_A_30_57#_c_113_n N_A_290_409#_c_241_n 0.0313457f $X=1.35 $Y=0.99 $X2=0
+ $Y2=0
cc_113 N_A_30_57#_c_114_n N_A_290_409#_c_241_n 0.0189241f $X=1.69 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_A_30_57#_c_113_n N_A_290_409#_c_242_n 0.0135189f $X=1.35 $Y=0.99 $X2=0
+ $Y2=0
cc_115 N_A_30_57#_c_114_n N_A_290_409#_c_242_n 0.0115646f $X=1.69 $Y=1.16 $X2=0
+ $Y2=0
cc_116 N_A_30_57#_c_110_n N_VPWR_c_322_n 0.0272606f $X=0.295 $Y=2.19 $X2=0 $Y2=0
cc_117 N_A_30_57#_M1005_g N_VPWR_c_324_n 0.00714077f $X=1.86 $Y=2.545 $X2=0
+ $Y2=0
cc_118 N_A_30_57#_M1005_g N_VPWR_c_321_n 0.012733f $X=1.86 $Y=2.545 $X2=0 $Y2=0
cc_119 N_A_30_57#_c_110_n N_VPWR_c_321_n 0.0095959f $X=0.295 $Y=2.19 $X2=0 $Y2=0
cc_120 N_A_30_57#_c_110_n N_VPWR_c_328_n 0.0167213f $X=0.295 $Y=2.19 $X2=0 $Y2=0
cc_121 N_A_30_57#_c_106_n N_VGND_c_377_n 0.0106034f $X=1.3 $Y=0.825 $X2=0 $Y2=0
cc_122 N_A_30_57#_c_107_n N_VGND_c_377_n 0.00188152f $X=1.69 $Y=0.825 $X2=0
+ $Y2=0
cc_123 N_A_30_57#_c_109_n N_VGND_c_377_n 0.0127138f $X=0.295 $Y=0.495 $X2=0
+ $Y2=0
cc_124 N_A_30_57#_c_111_n N_VGND_c_377_n 0.0169449f $X=1.185 $Y=0.91 $X2=0 $Y2=0
cc_125 N_A_30_57#_c_113_n N_VGND_c_377_n 0.00335429f $X=1.35 $Y=0.99 $X2=0 $Y2=0
cc_126 N_A_30_57#_c_109_n N_VGND_c_379_n 0.0220321f $X=0.295 $Y=0.495 $X2=0
+ $Y2=0
cc_127 N_A_30_57#_c_106_n N_VGND_c_380_n 0.00445056f $X=1.3 $Y=0.825 $X2=0 $Y2=0
cc_128 N_A_30_57#_c_107_n N_VGND_c_380_n 0.00440121f $X=1.69 $Y=0.825 $X2=0
+ $Y2=0
cc_129 N_A_30_57#_c_106_n N_VGND_c_382_n 0.00425382f $X=1.3 $Y=0.825 $X2=0 $Y2=0
cc_130 N_A_30_57#_c_107_n N_VGND_c_382_n 0.00781382f $X=1.69 $Y=0.825 $X2=0
+ $Y2=0
cc_131 N_A_30_57#_c_109_n N_VGND_c_382_n 0.0125808f $X=0.295 $Y=0.495 $X2=0
+ $Y2=0
cc_132 N_A_30_57#_c_111_n N_VGND_c_382_n 0.0152008f $X=1.185 $Y=0.91 $X2=0 $Y2=0
cc_133 N_A_30_57#_c_113_n N_VGND_c_382_n 0.00931021f $X=1.35 $Y=0.99 $X2=0 $Y2=0
cc_134 N_A_30_57#_c_114_n N_VGND_c_382_n 2.55086e-19 $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_174_n N_A_290_409#_M1003_g 0.0115242f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_136 N_A_M1010_g N_A_290_409#_M1000_g 0.0123786f $X=2.35 $Y=2.545 $X2=0 $Y2=0
cc_137 N_A_c_182_n N_A_290_409#_M1000_g 0.00487136f $X=2.39 $Y=1.885 $X2=0 $Y2=0
cc_138 N_A_c_179_n N_A_290_409#_M1000_g 0.00424593f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_139 N_A_c_177_n N_A_290_409#_c_237_n 0.0115242f $X=2.48 $Y=0.855 $X2=0 $Y2=0
cc_140 N_A_c_176_n N_A_290_409#_c_238_n 0.00487136f $X=2.39 $Y=1.72 $X2=0 $Y2=0
cc_141 N_A_c_178_n N_A_290_409#_c_238_n 0.0115242f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_142 N_A_c_179_n N_A_290_409#_c_238_n 0.002012f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_143 N_A_M1010_g N_A_290_409#_c_247_n 9.16379e-19 $X=2.35 $Y=2.545 $X2=0 $Y2=0
cc_144 N_A_c_182_n N_A_290_409#_c_247_n 4.00383e-19 $X=2.39 $Y=1.885 $X2=0 $Y2=0
cc_145 N_A_c_171_n N_A_290_409#_c_239_n 0.00997923f $X=2.12 $Y=0.78 $X2=0 $Y2=0
cc_146 N_A_c_173_n N_A_290_409#_c_239_n 0.00501241f $X=2.195 $Y=0.855 $X2=0
+ $Y2=0
cc_147 N_A_c_174_n N_A_290_409#_c_239_n 0.00161255f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_148 N_A_c_172_n N_A_290_409#_c_240_n 0.011861f $X=2.405 $Y=0.855 $X2=0 $Y2=0
cc_149 N_A_c_173_n N_A_290_409#_c_240_n 0.00825744f $X=2.195 $Y=0.855 $X2=0
+ $Y2=0
cc_150 N_A_c_175_n N_A_290_409#_c_240_n 0.00680017f $X=2.39 $Y=1.215 $X2=0 $Y2=0
cc_151 N_A_c_177_n N_A_290_409#_c_240_n 0.00757543f $X=2.48 $Y=0.855 $X2=0 $Y2=0
cc_152 N_A_c_178_n N_A_290_409#_c_240_n 5.71378e-19 $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_153 N_A_c_179_n N_A_290_409#_c_240_n 0.037145f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_154 N_A_c_176_n N_A_290_409#_c_248_n 4.00383e-19 $X=2.39 $Y=1.72 $X2=0 $Y2=0
cc_155 N_A_c_175_n N_A_290_409#_c_241_n 0.0027441f $X=2.39 $Y=1.215 $X2=0 $Y2=0
cc_156 N_A_c_178_n N_A_290_409#_c_241_n 7.11508e-19 $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_157 N_A_c_179_n N_A_290_409#_c_241_n 0.12903f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_158 N_A_c_173_n N_A_290_409#_c_242_n 0.00131872f $X=2.195 $Y=0.855 $X2=0
+ $Y2=0
cc_159 N_A_c_179_n N_A_290_409#_c_242_n 0.00215865f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_160 N_A_c_175_n N_A_290_409#_c_243_n 0.0023621f $X=2.39 $Y=1.215 $X2=0 $Y2=0
cc_161 N_A_c_179_n N_A_290_409#_c_243_n 0.0166193f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_162 N_A_c_175_n N_A_290_409#_c_244_n 0.0115242f $X=2.39 $Y=1.215 $X2=0 $Y2=0
cc_163 N_A_c_179_n N_A_290_409#_c_244_n 0.0012554f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_164 N_A_c_179_n N_VPWR_M1010_d 0.00873031f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_165 N_A_M1010_g N_VPWR_c_323_n 0.00925841f $X=2.35 $Y=2.545 $X2=0 $Y2=0
cc_166 N_A_c_179_n N_VPWR_c_323_n 0.0687883f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_167 N_A_M1010_g N_VPWR_c_324_n 0.00595064f $X=2.35 $Y=2.545 $X2=0 $Y2=0
cc_168 N_A_c_179_n N_VPWR_c_324_n 0.0139974f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_169 N_A_M1010_g N_VPWR_c_321_n 0.00803281f $X=2.35 $Y=2.545 $X2=0 $Y2=0
cc_170 N_A_c_179_n N_VPWR_c_321_n 0.0164665f $X=2.39 $Y=1.38 $X2=0 $Y2=0
cc_171 N_A_c_179_n A_397_409# 0.00896584f $X=2.39 $Y=1.38 $X2=-0.19 $Y2=-0.245
cc_172 N_A_c_171_n N_VGND_c_378_n 0.00200313f $X=2.12 $Y=0.78 $X2=0 $Y2=0
cc_173 N_A_c_174_n N_VGND_c_378_n 0.0114587f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_174 N_A_c_171_n N_VGND_c_380_n 0.00502664f $X=2.12 $Y=0.78 $X2=0 $Y2=0
cc_175 N_A_c_172_n N_VGND_c_380_n 4.57848e-19 $X=2.405 $Y=0.855 $X2=0 $Y2=0
cc_176 N_A_c_174_n N_VGND_c_380_n 0.00445056f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_177 N_A_c_171_n N_VGND_c_382_n 0.00942073f $X=2.12 $Y=0.78 $X2=0 $Y2=0
cc_178 N_A_c_172_n N_VGND_c_382_n 6.33118e-19 $X=2.405 $Y=0.855 $X2=0 $Y2=0
cc_179 N_A_c_174_n N_VGND_c_382_n 0.00796275f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_180 N_A_290_409#_c_248_n N_VPWR_c_322_n 0.0458292f $X=1.595 $Y=2.19 $X2=0
+ $Y2=0
cc_181 N_A_290_409#_M1000_g N_VPWR_c_323_n 0.0245466f $X=3.165 $Y=2.545 $X2=0
+ $Y2=0
cc_182 N_A_290_409#_c_238_n N_VPWR_c_323_n 0.0013627f $X=3.012 $Y=1.358 $X2=0
+ $Y2=0
cc_183 N_A_290_409#_c_243_n N_VPWR_c_323_n 0.00903485f $X=3 $Y=1.03 $X2=0 $Y2=0
cc_184 N_A_290_409#_c_247_n N_VPWR_c_324_n 0.0287481f $X=1.595 $Y=2.9 $X2=0
+ $Y2=0
cc_185 N_A_290_409#_M1000_g N_VPWR_c_326_n 0.00769046f $X=3.165 $Y=2.545 $X2=0
+ $Y2=0
cc_186 N_A_290_409#_M1000_g N_VPWR_c_321_n 0.0141514f $X=3.165 $Y=2.545 $X2=0
+ $Y2=0
cc_187 N_A_290_409#_c_247_n N_VPWR_c_321_n 0.0161599f $X=1.595 $Y=2.9 $X2=0
+ $Y2=0
cc_188 N_A_290_409#_M1003_g X 0.00207391f $X=2.91 $Y=0.495 $X2=0 $Y2=0
cc_189 N_A_290_409#_M1004_g X 0.0146991f $X=3.3 $Y=0.495 $X2=0 $Y2=0
cc_190 N_A_290_409#_c_237_n X 0.00625895f $X=3.3 $Y=0.94 $X2=0 $Y2=0
cc_191 N_A_290_409#_c_238_n X 0.0218629f $X=3.012 $Y=1.358 $X2=0 $Y2=0
cc_192 N_A_290_409#_c_243_n X 0.0501798f $X=3 $Y=1.03 $X2=0 $Y2=0
cc_193 N_A_290_409#_c_244_n X 0.0122687f $X=3 $Y=1.03 $X2=0 $Y2=0
cc_194 N_A_290_409#_M1000_g X 0.0150217f $X=3.165 $Y=2.545 $X2=0 $Y2=0
cc_195 N_A_290_409#_M1000_g X 0.00557033f $X=3.165 $Y=2.545 $X2=0 $Y2=0
cc_196 N_A_290_409#_c_239_n N_VGND_c_377_n 0.013209f $X=1.905 $Y=0.495 $X2=0
+ $Y2=0
cc_197 N_A_290_409#_M1003_g N_VGND_c_378_n 0.0117579f $X=2.91 $Y=0.495 $X2=0
+ $Y2=0
cc_198 N_A_290_409#_M1004_g N_VGND_c_378_n 0.00201912f $X=3.3 $Y=0.495 $X2=0
+ $Y2=0
cc_199 N_A_290_409#_c_239_n N_VGND_c_378_n 0.0141909f $X=1.905 $Y=0.495 $X2=0
+ $Y2=0
cc_200 N_A_290_409#_c_240_n N_VGND_c_378_n 0.0190137f $X=2.835 $Y=0.95 $X2=0
+ $Y2=0
cc_201 N_A_290_409#_c_243_n N_VGND_c_378_n 0.00188705f $X=3 $Y=1.03 $X2=0 $Y2=0
cc_202 N_A_290_409#_c_239_n N_VGND_c_380_n 0.0248273f $X=1.905 $Y=0.495 $X2=0
+ $Y2=0
cc_203 N_A_290_409#_M1003_g N_VGND_c_381_n 0.00445056f $X=2.91 $Y=0.495 $X2=0
+ $Y2=0
cc_204 N_A_290_409#_M1004_g N_VGND_c_381_n 0.00502664f $X=3.3 $Y=0.495 $X2=0
+ $Y2=0
cc_205 N_A_290_409#_M1003_g N_VGND_c_382_n 0.00433746f $X=2.91 $Y=0.495 $X2=0
+ $Y2=0
cc_206 N_A_290_409#_M1004_g N_VGND_c_382_n 0.0101479f $X=3.3 $Y=0.495 $X2=0
+ $Y2=0
cc_207 N_A_290_409#_c_239_n N_VGND_c_382_n 0.0140042f $X=1.905 $Y=0.495 $X2=0
+ $Y2=0
cc_208 N_A_290_409#_c_243_n N_VGND_c_382_n 0.0102007f $X=3 $Y=1.03 $X2=0 $Y2=0
cc_209 N_VPWR_c_326_n X 0.030123f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_210 N_VPWR_c_321_n X 0.017224f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_323_n X 0.0701565f $X=2.9 $Y=2.19 $X2=0 $Y2=0
cc_212 X N_VGND_c_378_n 0.0134093f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_213 X N_VGND_c_381_n 0.024392f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_214 X N_VGND_c_382_n 0.0139351f $X=3.515 $Y=0.47 $X2=0 $Y2=0
