* File: sky130_fd_sc_lp__a41o_4.pex.spice
* Created: Wed Sep  2 09:29:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41O_4%A_100_23# 1 2 3 12 16 20 24 28 32 36 40 42 52
+ 55 56 60 64 68 76
r116 73 74 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.005 $Y=1.49
+ $X2=1.435 $Y2=1.49
r117 68 69 18.392 $w=1.99e-07 $l=3e-07 $layer=LI1_cond $X=2.487 $Y=1.49
+ $X2=2.487 $Y2=1.79
r118 62 64 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.03 $Y=1.875
+ $X2=3.03 $Y2=1.98
r119 58 67 0.067832 $w=3.3e-07 $l=1.13e-07 $layer=LI1_cond $X=2.605 $Y=0.85
+ $X2=2.492 $Y2=0.85
r120 58 60 44.8754 $w=3.28e-07 $l=1.285e-06 $layer=LI1_cond $X=2.605 $Y=0.85
+ $X2=3.89 $Y2=0.85
r121 57 69 1.66034 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=2.595 $Y=1.79
+ $X2=2.487 $Y2=1.79
r122 56 62 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.865 $Y=1.79
+ $X2=3.03 $Y2=1.875
r123 56 57 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.865 $Y=1.79
+ $X2=2.595 $Y2=1.79
r124 55 68 4.91046 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.487 $Y=1.405
+ $X2=2.487 $Y2=1.49
r125 54 67 7.13466 $w=2.2e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.487 $Y=1.015
+ $X2=2.492 $Y2=0.85
r126 54 55 20.9048 $w=2.13e-07 $l=3.9e-07 $layer=LI1_cond $X=2.487 $Y=1.015
+ $X2=2.487 $Y2=1.405
r127 50 67 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.492 $Y=0.685
+ $X2=2.492 $Y2=0.85
r128 50 52 13.5732 $w=2.23e-07 $l=2.65e-07 $layer=LI1_cond $X=2.492 $Y=0.685
+ $X2=2.492 $Y2=0.42
r129 49 76 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.775 $Y=1.49
+ $X2=1.865 $Y2=1.49
r130 49 74 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.775 $Y=1.49
+ $X2=1.435 $Y2=1.49
r131 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.775
+ $Y=1.49 $X2=1.775 $Y2=1.49
r132 45 73 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.755 $Y=1.49
+ $X2=1.005 $Y2=1.49
r133 45 70 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.755 $Y=1.49
+ $X2=0.575 $Y2=1.49
r134 44 48 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.755 $Y=1.49
+ $X2=1.775 $Y2=1.49
r135 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.755
+ $Y=1.49 $X2=0.755 $Y2=1.49
r136 42 68 1.66034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.38 $Y=1.49
+ $X2=2.487 $Y2=1.49
r137 42 48 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.38 $Y=1.49
+ $X2=1.775 $Y2=1.49
r138 38 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.655
+ $X2=1.865 $Y2=1.49
r139 38 40 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.865 $Y=1.655
+ $X2=1.865 $Y2=2.465
r140 34 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.325
+ $X2=1.865 $Y2=1.49
r141 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.865 $Y=1.325
+ $X2=1.865 $Y2=0.665
r142 30 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.655
+ $X2=1.435 $Y2=1.49
r143 30 32 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.435 $Y=1.655
+ $X2=1.435 $Y2=2.465
r144 26 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.325
+ $X2=1.435 $Y2=1.49
r145 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.435 $Y=1.325
+ $X2=1.435 $Y2=0.665
r146 22 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.655
+ $X2=1.005 $Y2=1.49
r147 22 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.005 $Y=1.655
+ $X2=1.005 $Y2=2.465
r148 18 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.325
+ $X2=1.005 $Y2=1.49
r149 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.005 $Y=1.325
+ $X2=1.005 $Y2=0.665
r150 14 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.655
+ $X2=0.575 $Y2=1.49
r151 14 16 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.575 $Y=1.655
+ $X2=0.575 $Y2=2.465
r152 10 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.325
+ $X2=0.575 $Y2=1.49
r153 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.575 $Y=1.325
+ $X2=0.575 $Y2=0.665
r154 3 64 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.89
+ $Y=1.835 $X2=3.03 $Y2=1.98
r155 2 60 182 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_NDIFF $count=1 $X=3.75
+ $Y=0.235 $X2=3.89 $Y2=0.85
r156 1 67 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=2.37
+ $Y=0.245 $X2=2.51 $Y2=0.96
r157 1 52 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.37
+ $Y=0.245 $X2=2.51 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%B1 1 3 4 6 9 13 15 16 23
c51 23 0 2.3832e-19 $X=2.86 $Y=1.36
c52 16 0 1.72668e-20 $X=3.6 $Y=1.295
r53 23 25 55.7267 $w=3.33e-07 $l=3.85e-07 $layer=POLY_cond $X=2.86 $Y=1.357
+ $X2=3.245 $Y2=1.357
r54 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.86
+ $Y=1.36 $X2=2.86 $Y2=1.36
r55 21 23 6.51351 $w=3.33e-07 $l=4.5e-08 $layer=POLY_cond $X=2.815 $Y=1.357
+ $X2=2.86 $Y2=1.357
r56 20 21 13.027 $w=3.33e-07 $l=9e-08 $layer=POLY_cond $X=2.725 $Y=1.357
+ $X2=2.815 $Y2=1.357
r57 15 16 16.2698 $w=3.38e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.6 $Y2=1.365
r58 15 24 8.8128 $w=3.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.86 $Y2=1.365
r59 11 25 21.4384 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=3.245 $Y=1.525
+ $X2=3.245 $Y2=1.357
r60 11 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.245 $Y=1.525 $X2=3.245
+ $Y2=2.465
r61 7 21 21.4384 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=2.815 $Y=1.525
+ $X2=2.815 $Y2=1.357
r62 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.815 $Y=1.525 $X2=2.815
+ $Y2=2.465
r63 4 20 21.4384 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=2.725 $Y=1.19
+ $X2=2.725 $Y2=1.357
r64 4 6 168.7 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.725 $Y=1.19 $X2=2.725
+ $Y2=0.665
r65 1 20 62.2402 $w=3.33e-07 $l=4.3e-07 $layer=POLY_cond $X=2.295 $Y=1.357
+ $X2=2.725 $Y2=1.357
r66 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.295 $Y=1.195
+ $X2=2.295 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A1 1 3 6 8 10 13 15 16 24
c50 16 0 2.55659e-19 $X=4.56 $Y=1.295
c51 13 0 1.72668e-20 $X=4.105 $Y=2.465
r52 22 24 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.055 $Y=1.35
+ $X2=4.105 $Y2=1.35
r53 19 22 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.675 $Y=1.35
+ $X2=4.055 $Y2=1.35
r54 15 16 15.5196 $w=3.73e-07 $l=5.05e-07 $layer=LI1_cond $X=4.055 $Y=1.397
+ $X2=4.56 $Y2=1.397
r55 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.055
+ $Y=1.35 $X2=4.055 $Y2=1.35
r56 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.515
+ $X2=4.105 $Y2=1.35
r57 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.105 $Y=1.515
+ $X2=4.105 $Y2=2.465
r58 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.185
+ $X2=4.105 $Y2=1.35
r59 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.105 $Y=1.185
+ $X2=4.105 $Y2=0.655
r60 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.675 $Y=1.515
+ $X2=3.675 $Y2=1.35
r61 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.675 $Y=1.515
+ $X2=3.675 $Y2=2.465
r62 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.675 $Y=1.185
+ $X2=3.675 $Y2=1.35
r63 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.675 $Y=1.185
+ $X2=3.675 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A2 1 3 6 8 10 13 15 23
r45 21 23 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.99 $Y=1.35 $X2=5.01
+ $Y2=1.35
r46 19 21 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=4.965 $Y=1.35
+ $X2=4.99 $Y2=1.35
r47 17 19 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.535 $Y=1.35
+ $X2=4.965 $Y2=1.35
r48 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.35 $X2=4.99 $Y2=1.35
r49 11 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.01 $Y=1.515
+ $X2=5.01 $Y2=1.35
r50 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.01 $Y=1.515
+ $X2=5.01 $Y2=2.465
r51 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=1.35
r52 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=0.655
r53 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.535 $Y=1.515
+ $X2=4.535 $Y2=1.35
r54 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.535 $Y=1.515
+ $X2=4.535 $Y2=2.465
r55 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.535 $Y=1.185
+ $X2=4.535 $Y2=1.35
r56 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.535 $Y=1.185
+ $X2=4.535 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A3 3 7 9 11 12 13 14 16 17 18
c53 18 0 1.81092e-19 $X=6 $Y=1.295
r54 25 26 6.84227 $w=3.17e-07 $l=4.5e-08 $layer=POLY_cond $X=5.87 $Y=1.35
+ $X2=5.915 $Y2=1.35
r55 23 25 32.6909 $w=3.17e-07 $l=2.15e-07 $layer=POLY_cond $X=5.655 $Y=1.35
+ $X2=5.87 $Y2=1.35
r56 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.655
+ $Y=1.35 $X2=5.655 $Y2=1.35
r57 21 23 32.6909 $w=3.17e-07 $l=2.15e-07 $layer=POLY_cond $X=5.44 $Y=1.35
+ $X2=5.655 $Y2=1.35
r58 18 24 12.8256 $w=3.08e-07 $l=3.45e-07 $layer=LI1_cond $X=6 $Y=1.365
+ $X2=5.655 $Y2=1.365
r59 17 24 5.0187 $w=3.08e-07 $l=1.35e-07 $layer=LI1_cond $X=5.52 $Y=1.365
+ $X2=5.655 $Y2=1.365
r60 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.345 $Y=1.185
+ $X2=6.345 $Y2=0.655
r61 13 26 24.856 $w=3.17e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.99 $Y=1.26
+ $X2=5.915 $Y2=1.35
r62 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.27 $Y=1.26
+ $X2=6.345 $Y2=1.185
r63 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.27 $Y=1.26
+ $X2=5.99 $Y2=1.26
r64 9 26 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.185
+ $X2=5.915 $Y2=1.35
r65 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.915 $Y=1.185
+ $X2=5.915 $Y2=0.655
r66 5 25 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.87 $Y=1.515
+ $X2=5.87 $Y2=1.35
r67 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.87 $Y=1.515 $X2=5.87
+ $Y2=2.465
r68 1 21 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.44 $Y=1.515
+ $X2=5.44 $Y2=1.35
r69 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.44 $Y=1.515 $X2=5.44
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A4 3 5 6 9 13 17 19 20 21 28
c46 13 0 6.9427e-20 $X=6.775 $Y=0.655
c47 5 0 4.5713e-21 $X=6.655 $Y=1.62
r48 28 30 12.2542 $w=3.54e-07 $l=9e-08 $layer=POLY_cond $X=7.115 $Y=1.51
+ $X2=7.205 $Y2=1.51
r49 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.115
+ $Y=1.49 $X2=7.115 $Y2=1.49
r50 26 28 46.2938 $w=3.54e-07 $l=3.4e-07 $layer=POLY_cond $X=6.775 $Y=1.51
+ $X2=7.115 $Y2=1.51
r51 25 26 6.12712 $w=3.54e-07 $l=4.5e-08 $layer=POLY_cond $X=6.73 $Y=1.51
+ $X2=6.775 $Y2=1.51
r52 21 29 10.2615 $w=3.63e-07 $l=3.25e-07 $layer=LI1_cond $X=7.44 $Y=1.392
+ $X2=7.115 $Y2=1.392
r53 20 29 4.89394 $w=3.63e-07 $l=1.55e-07 $layer=LI1_cond $X=6.96 $Y=1.392
+ $X2=7.115 $Y2=1.392
r54 19 20 15.1554 $w=3.63e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.392
+ $X2=6.96 $Y2=1.392
r55 15 30 22.9014 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=7.205 $Y=1.325
+ $X2=7.205 $Y2=1.51
r56 15 17 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.205 $Y=1.325
+ $X2=7.205 $Y2=0.655
r57 11 26 22.9014 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=6.775 $Y=1.325
+ $X2=6.775 $Y2=1.51
r58 11 13 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.775 $Y=1.325
+ $X2=6.775 $Y2=0.655
r59 7 25 22.9014 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=6.73 $Y=1.695
+ $X2=6.73 $Y2=1.51
r60 7 9 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.73 $Y=1.695 $X2=6.73
+ $Y2=2.465
r61 5 25 26.5778 $w=3.54e-07 $l=1.42653e-07 $layer=POLY_cond $X=6.655 $Y=1.62
+ $X2=6.73 $Y2=1.51
r62 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.655 $Y=1.62
+ $X2=6.375 $Y2=1.62
r63 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.3 $Y=1.695
+ $X2=6.375 $Y2=1.62
r64 1 3 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.3 $Y=1.695 $X2=6.3
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%VPWR 1 2 3 4 5 6 7 22 24 30 36 42 48 52 56 62
+ 67 68 69 70 71 73 78 90 97 98 104 107 110 113
c120 36 0 9.43259e-20 $X=2.08 $Y=1.98
r121 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r124 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r126 98 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r127 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r128 95 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.68 $Y=3.33
+ $X2=6.515 $Y2=3.33
r129 95 97 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.68 $Y=3.33
+ $X2=7.44 $Y2=3.33
r130 94 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r131 94 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r132 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r133 91 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=3.33
+ $X2=5.655 $Y2=3.33
r134 91 93 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.82 $Y=3.33 $X2=6
+ $Y2=3.33
r135 90 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.35 $Y=3.33
+ $X2=6.515 $Y2=3.33
r136 90 93 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.35 $Y=3.33 $X2=6
+ $Y2=3.33
r137 89 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r138 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r139 86 108 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.16 $Y2=3.33
r140 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r141 83 107 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.092 $Y2=3.33
r142 83 85 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 82 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r144 82 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r145 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r146 79 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.22 $Y2=3.33
r147 79 81 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.68 $Y2=3.33
r148 78 107 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.95 $Y=3.33
+ $X2=2.092 $Y2=3.33
r149 78 81 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.95 $Y=3.33
+ $X2=1.68 $Y2=3.33
r150 77 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r151 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r152 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r153 74 101 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.262 $Y2=3.33
r154 74 76 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.72 $Y2=3.33
r155 73 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.22 $Y2=3.33
r156 73 76 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r157 71 89 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 71 86 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r159 69 88 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r160 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.77 $Y2=3.33
r161 67 85 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=3.6 $Y2=3.33
r162 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=3.89 $Y2=3.33
r163 66 88 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.055 $Y=3.33
+ $X2=4.56 $Y2=3.33
r164 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=3.33
+ $X2=3.89 $Y2=3.33
r165 62 65 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.515 $Y=2.18
+ $X2=6.515 $Y2=2.95
r166 60 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.515 $Y=3.245
+ $X2=6.515 $Y2=3.33
r167 60 65 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.515 $Y=3.245
+ $X2=6.515 $Y2=2.95
r168 56 59 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=5.655 $Y=2.18
+ $X2=5.655 $Y2=2.95
r169 54 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=3.33
r170 54 59 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=2.95
r171 53 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=4.77 $Y2=3.33
r172 52 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.655 $Y2=3.33
r173 52 53 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=4.935 $Y2=3.33
r174 48 51 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.77 $Y=2.18
+ $X2=4.77 $Y2=2.95
r175 46 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=3.33
r176 46 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=2.95
r177 42 45 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.89 $Y=2.18
+ $X2=3.89 $Y2=2.95
r178 40 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=3.245
+ $X2=3.89 $Y2=3.33
r179 40 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.89 $Y=3.245
+ $X2=3.89 $Y2=2.95
r180 36 39 39.2235 $w=2.83e-07 $l=9.7e-07 $layer=LI1_cond $X=2.092 $Y=1.98
+ $X2=2.092 $Y2=2.95
r181 34 107 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.092 $Y=3.245
+ $X2=2.092 $Y2=3.33
r182 34 39 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=2.092 $Y=3.245
+ $X2=2.092 $Y2=2.95
r183 30 33 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.22 $Y=2.18
+ $X2=1.22 $Y2=2.95
r184 28 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r185 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.95
r186 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.36 $Y=2.18
+ $X2=0.36 $Y2=2.95
r187 22 101 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.262 $Y2=3.33
r188 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.36 $Y2=2.95
r189 7 65 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.375
+ $Y=1.835 $X2=6.515 $Y2=2.95
r190 7 62 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=6.375
+ $Y=1.835 $X2=6.515 $Y2=2.18
r191 6 59 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.515
+ $Y=1.835 $X2=5.655 $Y2=2.95
r192 6 56 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=5.515
+ $Y=1.835 $X2=5.655 $Y2=2.18
r193 5 51 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=4.61
+ $Y=1.835 $X2=4.77 $Y2=2.95
r194 5 48 400 $w=1.7e-07 $l=4.17403e-07 $layer=licon1_PDIFF $count=1 $X=4.61
+ $Y=1.835 $X2=4.77 $Y2=2.18
r195 4 45 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.75
+ $Y=1.835 $X2=3.89 $Y2=2.95
r196 4 42 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=3.75
+ $Y=1.835 $X2=3.89 $Y2=2.18
r197 3 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=2.95
r198 3 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=1.98
r199 2 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=2.95
r200 2 30 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=2.18
r201 1 27 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=2.95
r202 1 24 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%X 1 2 3 4 13 15 16 19 23 27 29 33 37 42 43 44
+ 45 49 51
r58 49 51 2.52097 $w=3.18e-07 $l=7e-08 $layer=LI1_cond $X=0.26 $Y=1.225 $X2=0.26
+ $Y2=1.295
r59 44 49 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.14 $X2=0.26
+ $Y2=1.225
r60 44 45 13.073 $w=3.18e-07 $l=3.63e-07 $layer=LI1_cond $X=0.26 $Y=1.302
+ $X2=0.26 $Y2=1.665
r61 44 51 0.252097 $w=3.18e-07 $l=7e-09 $layer=LI1_cond $X=0.26 $Y=1.302
+ $X2=0.26 $Y2=1.295
r62 41 45 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=0.26 $Y=1.755 $X2=0.26
+ $Y2=1.665
r63 37 39 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=1.667 $Y=1.98
+ $X2=1.667 $Y2=2.91
r64 35 37 2.81708 $w=2.23e-07 $l=5.5e-08 $layer=LI1_cond $X=1.667 $Y=1.925
+ $X2=1.667 $Y2=1.98
r65 31 33 32.5245 $w=2.23e-07 $l=6.35e-07 $layer=LI1_cond $X=1.667 $Y=1.055
+ $X2=1.667 $Y2=0.42
r66 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.885 $Y=1.84
+ $X2=0.79 $Y2=1.84
r67 29 35 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.555 $Y=1.84
+ $X2=1.667 $Y2=1.925
r68 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.555 $Y=1.84
+ $X2=0.885 $Y2=1.84
r69 28 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.885 $Y=1.14
+ $X2=0.79 $Y2=1.14
r70 27 31 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.555 $Y=1.14
+ $X2=1.667 $Y2=1.055
r71 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.555 $Y=1.14
+ $X2=0.885 $Y2=1.14
r72 23 25 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.79 $Y=1.98
+ $X2=0.79 $Y2=2.91
r73 21 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=1.925
+ $X2=0.79 $Y2=1.84
r74 21 23 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=0.79 $Y=1.925
+ $X2=0.79 $Y2=1.98
r75 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=1.055
+ $X2=0.79 $Y2=1.14
r76 17 19 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.79 $Y=1.055
+ $X2=0.79 $Y2=0.42
r77 16 41 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=0.42 $Y=1.84
+ $X2=0.26 $Y2=1.755
r78 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.695 $Y=1.84
+ $X2=0.79 $Y2=1.84
r79 15 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.695 $Y=1.84
+ $X2=0.42 $Y2=1.84
r80 14 44 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.42 $Y=1.14 $X2=0.26
+ $Y2=1.14
r81 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.695 $Y=1.14
+ $X2=0.79 $Y2=1.14
r82 13 14 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.695 $Y=1.14
+ $X2=0.42 $Y2=1.14
r83 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=2.91
r84 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=1.98
r85 3 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.835 $X2=0.79 $Y2=2.91
r86 3 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.835 $X2=0.79 $Y2=1.98
r87 2 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.245 $X2=1.65 $Y2=0.42
r88 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.65
+ $Y=0.245 $X2=0.79 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A_495_367# 1 2 3 4 5 6 19 21 23 26 29 30 33
+ 37 41 45 49 53 57 65 66 67
r78 57 59 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=6.98 $Y=1.98 $X2=6.98
+ $Y2=2.91
r79 55 57 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=6.98 $Y=1.925
+ $X2=6.98 $Y2=1.98
r80 54 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.18 $Y=1.84
+ $X2=6.085 $Y2=1.84
r81 53 55 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.85 $Y=1.84
+ $X2=6.98 $Y2=1.925
r82 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.85 $Y=1.84
+ $X2=6.18 $Y2=1.84
r83 49 51 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.085 $Y=1.98
+ $X2=6.085 $Y2=2.91
r84 47 67 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=1.925
+ $X2=6.085 $Y2=1.84
r85 47 49 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.085 $Y=1.925
+ $X2=6.085 $Y2=1.98
r86 46 66 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.32 $Y=1.84
+ $X2=5.215 $Y2=1.84
r87 45 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.99 $Y=1.84
+ $X2=6.085 $Y2=1.84
r88 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.99 $Y=1.84
+ $X2=5.32 $Y2=1.84
r89 41 43 49.1169 $w=2.08e-07 $l=9.3e-07 $layer=LI1_cond $X=5.215 $Y=1.98
+ $X2=5.215 $Y2=2.91
r90 39 66 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=1.925
+ $X2=5.215 $Y2=1.84
r91 39 41 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=5.215 $Y=1.925
+ $X2=5.215 $Y2=1.98
r92 38 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.415 $Y=1.84
+ $X2=4.32 $Y2=1.84
r93 37 66 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.11 $Y=1.84
+ $X2=5.215 $Y2=1.84
r94 37 38 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.11 $Y=1.84
+ $X2=4.415 $Y2=1.84
r95 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.32 $Y=1.98
+ $X2=4.32 $Y2=2.91
r96 31 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.32 $Y=1.925
+ $X2=4.32 $Y2=1.84
r97 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.32 $Y=1.925
+ $X2=4.32 $Y2=1.98
r98 29 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.225 $Y=1.84
+ $X2=4.32 $Y2=1.84
r99 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.225 $Y=1.84
+ $X2=3.555 $Y2=1.84
r100 26 64 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=2.905
+ $X2=3.46 $Y2=2.99
r101 26 28 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=3.46 $Y=2.905
+ $X2=3.46 $Y2=1.98
r102 25 30 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.46 $Y=1.925
+ $X2=3.555 $Y2=1.84
r103 25 28 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=3.46 $Y=1.925
+ $X2=3.46 $Y2=1.98
r104 24 62 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.695 $Y=2.99
+ $X2=2.565 $Y2=2.99
r105 23 64 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.365 $Y=2.99
+ $X2=3.46 $Y2=2.99
r106 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.365 $Y=2.99
+ $X2=2.695 $Y2=2.99
r107 19 62 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=2.905
+ $X2=2.565 $Y2=2.99
r108 19 21 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=2.565 $Y=2.905
+ $X2=2.565 $Y2=2.21
r109 6 59 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=1.835 $X2=6.945 $Y2=2.91
r110 6 57 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=1.835 $X2=6.945 $Y2=1.98
r111 5 51 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.945
+ $Y=1.835 $X2=6.085 $Y2=2.91
r112 5 49 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.945
+ $Y=1.835 $X2=6.085 $Y2=1.98
r113 4 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.085
+ $Y=1.835 $X2=5.225 $Y2=2.91
r114 4 41 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.085
+ $Y=1.835 $X2=5.225 $Y2=1.98
r115 3 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=2.91
r116 3 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=1.98
r117 2 64 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.835 $X2=3.46 $Y2=2.91
r118 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.835 $X2=3.46 $Y2=1.98
r119 1 62 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.835 $X2=2.6 $Y2=2.91
r120 1 21 400 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.835 $X2=2.6 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 42 44 56 65 66 72 75
r105 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r106 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r107 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r108 66 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r109 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r110 63 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=0 $X2=6.99
+ $Y2=0
r111 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.155 $Y=0
+ $X2=7.44 $Y2=0
r112 62 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r113 61 62 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r114 58 61 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=6.48
+ $Y2=0
r115 58 59 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r116 56 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.99
+ $Y2=0
r117 56 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.48
+ $Y2=0
r118 55 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r119 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r120 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r121 52 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r122 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r123 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r124 49 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r125 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r126 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r127 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r128 45 69 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.262 $Y2=0
r129 45 47 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.72 $Y2=0
r130 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r131 44 47 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r132 42 62 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=6.48
+ $Y2=0
r133 42 59 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r134 40 54 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0
+ $X2=2.64 $Y2=0
r135 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.94
+ $Y2=0
r136 39 58 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.12
+ $Y2=0
r137 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.94
+ $Y2=0
r138 37 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=1.68
+ $Y2=0
r139 37 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=2.08
+ $Y2=0
r140 36 54 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.64
+ $Y2=0
r141 36 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.08
+ $Y2=0
r142 32 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0
r143 32 34 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0.535
r144 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0
r145 28 30 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.41
r146 24 38 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r147 24 26 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.39
r148 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r149 20 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.37
r150 16 69 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.262 $Y2=0
r151 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.36 $Y2=0.39
r152 5 34 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=6.85
+ $Y=0.235 $X2=6.99 $Y2=0.535
r153 4 30 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.245 $X2=2.94 $Y2=0.41
r154 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.94
+ $Y=0.245 $X2=2.08 $Y2=0.39
r155 2 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.245 $X2=1.22 $Y2=0.37
r156 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.235
+ $Y=0.245 $X2=0.36 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A_667_47# 1 2 3 10 14 15 18
r29 16 23 3.54615 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=4.425 $Y=0.89
+ $X2=4.29 $Y2=0.89
r30 16 18 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=4.425 $Y=0.89
+ $X2=5.18 $Y2=0.89
r31 15 23 3.28347 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.29 $Y=0.765
+ $X2=4.29 $Y2=0.89
r32 14 21 3.28347 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.29 $Y=0.505
+ $X2=4.29 $Y2=0.38
r33 14 15 11.0976 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.29 $Y=0.505
+ $X2=4.29 $Y2=0.765
r34 10 21 3.54615 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=0.38
+ $X2=4.29 $Y2=0.38
r35 10 12 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.155 $Y=0.38
+ $X2=3.46 $Y2=0.38
r36 3 18 182 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.18 $Y2=0.88
r37 2 23 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.235 $X2=4.32 $Y2=0.875
r38 2 21 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.235 $X2=4.32 $Y2=0.42
r39 1 12 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.235 $X2=3.46 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A_922_47# 1 2 11
r16 8 11 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=4.75 $Y=0.43
+ $X2=6.13 $Y2=0.43
r17 2 11 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.235 $X2=6.13 $Y2=0.43
r18 1 8 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=4.61
+ $Y=0.235 $X2=4.75 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_4%A_1115_47# 1 2 3 10 16 18 22 24
c33 10 0 4.5713e-21 $X=6.405 $Y=0.902
r34 20 22 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=7.455 $Y=0.87
+ $X2=7.455 $Y2=0.42
r35 19 24 5.68576 $w=2.22e-07 $l=1.49164e-07 $layer=LI1_cond $X=6.655 $Y=0.955
+ $X2=6.53 $Y2=0.902
r36 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.325 $Y=0.955
+ $X2=7.455 $Y2=0.87
r37 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.325 $Y=0.955
+ $X2=6.655 $Y2=0.955
r38 14 24 0.926478 $w=2.5e-07 $l=1.37e-07 $layer=LI1_cond $X=6.53 $Y=0.765
+ $X2=6.53 $Y2=0.902
r39 14 16 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=6.53 $Y=0.765
+ $X2=6.53 $Y2=0.42
r40 10 24 5.68576 $w=2.22e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=0.902
+ $X2=6.53 $Y2=0.902
r41 10 12 29.5444 $w=2.73e-07 $l=7.05e-07 $layer=LI1_cond $X=6.405 $Y=0.902
+ $X2=5.7 $Y2=0.902
r42 3 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.28
+ $Y=0.235 $X2=7.42 $Y2=0.42
r43 2 16 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.42
+ $Y=0.235 $X2=6.56 $Y2=0.42
r44 1 12 182 $w=1.7e-07 $l=7.04734e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.7 $Y2=0.88
.ends

