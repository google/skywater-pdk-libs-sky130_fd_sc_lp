* File: sky130_fd_sc_lp__a2111oi_m.pex.spice
* Created: Wed Sep  2 09:17:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111OI_M%D1 3 7 11 12 13 14 15 16 17 24
r35 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.375 $X2=0.61 $Y2=1.375
r36 16 17 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=2.405
+ $X2=0.665 $Y2=2.775
r37 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.665 $Y2=2.405
r38 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=1.665
+ $X2=0.665 $Y2=2.035
r39 14 25 11.936 $w=2.78e-07 $l=2.9e-07 $layer=LI1_cond $X=0.665 $Y=1.665
+ $X2=0.665 $Y2=1.375
r40 13 25 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=0.665 $Y=1.295
+ $X2=0.665 $Y2=1.375
r41 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.61 $Y=1.715
+ $X2=0.61 $Y2=1.375
r42 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.715
+ $X2=0.61 $Y2=1.88
r43 10 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.21
+ $X2=0.61 $Y2=1.375
r44 7 12 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=0.7 $Y=2.875 $X2=0.7
+ $Y2=1.88
r45 3 10 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.7 $Y=0.445 $X2=0.7
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%C1 3 7 11 12 13 14 15 20 21
r40 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.06 $X2=1.15 $Y2=1.06
r41 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=2.035
r42 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.665
r43 13 21 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.06
r44 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.15 $Y=1.4 $X2=1.15
+ $Y2=1.06
r45 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.4
+ $X2=1.15 $Y2=1.565
r46 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=0.895
+ $X2=1.15 $Y2=1.06
r47 7 10 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.13 $Y=0.445
+ $X2=1.13 $Y2=0.895
r48 3 12 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=1.06 $Y=2.875
+ $X2=1.06 $Y2=1.565
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%B1 3 7 12 16 17 18 23
r46 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.45 $X2=1.69 $Y2=1.45
r47 17 18 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=2.035
r48 17 24 13.2475 $w=1.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.45
r49 16 24 9.5505 $w=1.78e-07 $l=1.55e-07 $layer=LI1_cond $X=1.685 $Y=1.295
+ $X2=1.685 $Y2=1.45
r50 15 23 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.285
+ $X2=1.69 $Y2=1.45
r51 12 23 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.69 $Y=1.805
+ $X2=1.69 $Y2=1.45
r52 9 12 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.42 $Y=1.88 $X2=1.69
+ $Y2=1.88
r53 7 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.71 $Y=0.445
+ $X2=1.71 $Y2=1.285
r54 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=1.955 $X2=1.42
+ $Y2=1.88
r55 1 3 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.42 $Y=1.955 $X2=1.42
+ $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%A1 1 3 7 11 14 15 16 21
r41 15 16 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=2.035
r42 15 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.69 $X2=2.23 $Y2=1.69
r43 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.295
+ $X2=2.195 $Y2=1.665
r44 13 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.525
+ $X2=2.23 $Y2=1.69
r45 11 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=2.03
+ $X2=2.23 $Y2=1.69
r46 7 13 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=2.14 $Y=0.445
+ $X2=2.14 $Y2=1.525
r47 1 11 94.4124 $w=1.94e-07 $l=4.5215e-07 $layer=POLY_cond $X=1.85 $Y=2.345
+ $X2=2.23 $Y2=2.187
r48 1 3 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.85 $Y=2.345 $X2=1.85
+ $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%A2 3 5 7 8 9 10 11 13 16 17 18 19 20 21 28
r38 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.085
+ $Y=1.12 $X2=3.085 $Y2=1.12
r39 20 21 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.102 $Y=1.665
+ $X2=3.102 $Y2=2.035
r40 19 20 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.102 $Y=1.295
+ $X2=3.102 $Y2=1.665
r41 19 29 9.46785 $w=2.03e-07 $l=1.75e-07 $layer=LI1_cond $X=3.102 $Y=1.295
+ $X2=3.102 $Y2=1.12
r42 18 29 10.5499 $w=2.03e-07 $l=1.95e-07 $layer=LI1_cond $X=3.102 $Y=0.925
+ $X2=3.102 $Y2=1.12
r43 17 18 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.102 $Y=0.555
+ $X2=3.102 $Y2=0.925
r44 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.085 $Y=1.46
+ $X2=3.085 $Y2=1.12
r45 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.46
+ $X2=3.085 $Y2=1.625
r46 14 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.085 $Y=1.105
+ $X2=3.085 $Y2=1.12
r47 13 16 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.995 $Y=2.405
+ $X2=2.995 $Y2=1.625
r48 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.92 $Y=2.48
+ $X2=2.995 $Y2=2.405
r49 10 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.92 $Y=2.48
+ $X2=2.575 $Y2=2.48
r50 8 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.92 $Y=1.03
+ $X2=3.085 $Y2=1.105
r51 8 9 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.92 $Y=1.03
+ $X2=2.575 $Y2=1.03
r52 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.5 $Y=2.555
+ $X2=2.575 $Y2=2.48
r53 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.5 $Y=2.555 $X2=2.5
+ $Y2=2.875
r54 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.5 $Y=0.955
+ $X2=2.575 $Y2=1.03
r55 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.5 $Y=0.955 $X2=2.5
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%Y 1 2 3 12 14 15 16 20 22 28
r48 22 28 5.48116 $w=3.45e-07 $l=1.55e-07 $layer=LI1_cond $X=0.827 $Y=0.555
+ $X2=0.827 $Y2=0.71
r49 22 25 1.5913 $w=3.45e-07 $l=4.5e-08 $layer=LI1_cond $X=0.827 $Y=0.555
+ $X2=0.827 $Y2=0.51
r50 18 20 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.925 $Y=0.625
+ $X2=1.925 $Y2=0.51
r51 17 28 4.88813 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.02 $Y=0.71
+ $X2=0.827 $Y2=0.71
r52 16 18 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.82 $Y=0.71
+ $X2=1.925 $Y2=0.625
r53 16 17 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.82 $Y=0.71 $X2=1.02
+ $Y2=0.71
r54 14 28 3.53623 $w=3.45e-07 $l=2.36778e-07 $layer=LI1_cond $X=0.635 $Y=0.81
+ $X2=0.827 $Y2=0.71
r55 14 15 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.635 $Y=0.81
+ $X2=0.345 $Y2=0.81
r56 10 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.25 $Y=0.895
+ $X2=0.345 $Y2=0.81
r57 10 12 111.785 $w=1.88e-07 $l=1.915e-06 $layer=LI1_cond $X=0.25 $Y=0.895
+ $X2=0.25 $Y2=2.81
r58 3 12 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.665 $X2=0.26 $Y2=2.81
r59 2 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.235 $X2=1.925 $Y2=0.51
r60 1 25 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.235 $X2=0.915 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%A_299_533# 1 2 9 11 12 13
c30 9 0 1.69038e-19 $X=1.635 $Y=2.81
r31 13 16 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.715 $Y=2.57
+ $X2=2.715 $Y2=2.81
r32 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=2.57
+ $X2=2.715 $Y2=2.57
r33 11 12 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.55 $Y=2.57
+ $X2=1.74 $Y2=2.57
r34 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.635 $Y=2.655
+ $X2=1.74 $Y2=2.57
r35 7 9 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.635 $Y=2.655
+ $X2=1.635 $Y2=2.81
r36 2 16 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.665 $X2=2.715 $Y2=2.81
r37 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.665 $X2=1.635 $Y2=2.81
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%VPWR 1 6 8 10 20 21 24
r39 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.085 $Y2=3.33
r43 18 20 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=2.085 $Y2=3.33
r47 10 16 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=3.245
+ $X2=2.085 $Y2=3.33
r52 4 6 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.085 $Y=3.245
+ $X2=2.085 $Y2=2.94
r53 1 6 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=2.665 $X2=2.085 $Y2=2.94
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_M%VGND 1 2 3 10 12 14 18 22 24 26 33 34 40
+ 43
r48 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r51 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 34 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r53 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 31 43 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=2.715
+ $Y2=0
r55 31 33 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=3.12
+ $Y2=0
r56 27 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.365
+ $Y2=0
r57 27 29 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.68
+ $Y2=0
r58 26 43 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.61 $Y=0 $X2=2.715
+ $Y2=0
r59 26 29 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.61 $Y=0 $X2=1.68
+ $Y2=0
r60 24 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r61 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r62 24 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r63 20 43 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0
r64 20 22 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0.38
r65 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0
r66 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0.36
r67 15 37 3.49867 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r68 14 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.365
+ $Y2=0
r69 14 15 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=0.455
+ $Y2=0
r70 10 37 3.34522 $w=1.9e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.227 $Y2=0
r71 10 12 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.36 $Y=0.085
+ $X2=0.36 $Y2=0.38
r72 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.235 $X2=2.715 $Y2=0.38
r73 2 18 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=1.205
+ $Y=0.235 $X2=1.365 $Y2=0.36
r74 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.38
.ends

