* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4_2 A B C D VGND VNB VPB VPWR X
X0 VPWR A a_72_49# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_72_49# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_72_49# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 X a_72_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_72_49# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_72_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_227_49# C a_335_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_335_49# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_72_49# A a_155_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR C a_72_49# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_72_49# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_155_49# B a_227_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
