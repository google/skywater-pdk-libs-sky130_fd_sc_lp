* File: sky130_fd_sc_lp__xor2_lp.pex.spice
* Created: Wed Sep  2 10:41:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR2_LP%A_84_93# 1 2 9 13 17 20 21 22 25 29 31 33 34
+ 36 39 41 44
c109 41 0 1.53328e-19 $X=0.82 $Y=1.73
c110 34 0 1.96367e-20 $X=2.925 $Y=0.915
r111 45 46 27.4756 $w=3.07e-07 $l=1.75e-07 $layer=POLY_cond $X=0.495 $Y=1.73
+ $X2=0.67 $Y2=1.73
r112 39 48 24.3355 $w=3.07e-07 $l=1.55e-07 $layer=POLY_cond $X=0.7 $Y=1.73
+ $X2=0.855 $Y2=1.73
r113 39 46 4.7101 $w=3.07e-07 $l=3e-08 $layer=POLY_cond $X=0.7 $Y=1.73 $X2=0.67
+ $Y2=1.73
r114 38 41 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.7 $Y=1.73 $X2=0.82
+ $Y2=1.73
r115 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.73 $X2=0.7 $Y2=1.73
r116 35 36 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.53 $Y=1 $X2=3.53
+ $Y2=2.04
r117 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=0.915
+ $X2=3.53 $Y2=1
r118 33 34 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.445 $Y=0.915
+ $X2=2.925 $Y2=0.915
r119 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=2.125
+ $X2=2.56 $Y2=2.125
r120 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=2.125
+ $X2=3.53 $Y2=2.04
r121 31 32 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.445 $Y=2.125
+ $X2=2.725 $Y2=2.125
r122 27 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.76 $Y=0.83
+ $X2=2.925 $Y2=0.915
r123 27 29 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.76 $Y=0.83
+ $X2=2.76 $Y2=0.55
r124 23 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=2.21
+ $X2=2.56 $Y2=2.125
r125 23 25 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.56 $Y=2.21
+ $X2=2.56 $Y2=2.9
r126 21 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=2.125
+ $X2=2.56 $Y2=2.125
r127 21 22 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=2.395 $Y=2.125
+ $X2=0.905 $Y2=2.125
r128 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.82 $Y=2.04
+ $X2=0.905 $Y2=2.125
r129 19 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=1.895
+ $X2=0.82 $Y2=1.73
r130 19 20 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.82 $Y=1.895
+ $X2=0.82 $Y2=2.04
r131 15 48 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.855 $Y=1.565
+ $X2=0.855 $Y2=1.73
r132 15 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.855 $Y=1.565
+ $X2=0.855 $Y2=0.805
r133 11 46 7.67377 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=1.895
+ $X2=0.67 $Y2=1.73
r134 11 13 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.67 $Y=1.895
+ $X2=0.67 $Y2=2.595
r135 7 45 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.565
+ $X2=0.495 $Y2=1.73
r136 7 9 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=1.565
+ $X2=0.495 $Y2=0.805
r137 2 44 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.06 $X2=2.56 $Y2=2.205
r138 2 25 400 $w=1.7e-07 $l=9.09615e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.06 $X2=2.56 $Y2=2.9
r139 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.34 $X2=2.76 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_LP%A 1 3 6 7 10 14 18 22 24 25 29 32 33 37 46
+ 54
c105 37 0 5.85314e-20 $X=1.735 $Y=1.46
c106 7 0 3.47863e-19 $X=1.325 $Y=1.55
r107 45 46 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.285 $Y=1.345
+ $X2=3.335 $Y2=1.345
r108 38 54 9.92865 $w=5.63e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.577
+ $X2=1.9 $Y2=1.577
r109 37 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.735 $Y=1.46
+ $X2=1.735 $Y2=1.55
r110 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.735 $Y=1.46
+ $X2=1.735 $Y2=1.295
r111 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.46 $X2=1.735 $Y2=1.46
r112 33 38 1.16432 $w=5.63e-07 $l=5.5e-08 $layer=LI1_cond $X=1.68 $Y=1.577
+ $X2=1.735 $Y2=1.577
r113 32 33 10.1614 $w=5.63e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.577
+ $X2=1.68 $Y2=1.577
r114 30 45 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.1 $Y=1.345
+ $X2=3.285 $Y2=1.345
r115 30 42 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.1 $Y=1.345
+ $X2=2.975 $Y2=1.345
r116 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.345 $X2=3.1 $Y2=1.345
r117 27 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.1 $Y=1.69
+ $X2=3.1 $Y2=1.345
r118 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.935 $Y=1.775
+ $X2=3.1 $Y2=1.69
r119 25 54 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.935 $Y=1.775
+ $X2=1.9 $Y2=1.775
r120 20 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=1.18
+ $X2=3.335 $Y2=1.345
r121 20 22 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.335 $Y=1.18
+ $X2=3.335 $Y2=0.55
r122 16 45 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.51
+ $X2=3.285 $Y2=1.345
r123 16 18 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=3.285 $Y=1.51
+ $X2=3.285 $Y2=2.56
r124 12 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.18
+ $X2=2.975 $Y2=1.345
r125 12 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.975 $Y=1.18
+ $X2=2.975 $Y2=0.55
r126 10 39 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.645 $Y=0.805
+ $X2=1.645 $Y2=1.295
r127 6 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.55
+ $X2=1.735 $Y2=1.55
r128 6 7 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.57 $Y=1.55
+ $X2=1.325 $Y2=1.55
r129 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.25 $Y=1.625
+ $X2=1.325 $Y2=1.55
r130 4 24 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.25 $Y=1.625
+ $X2=1.25 $Y2=1.955
r131 1 24 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.2 $Y=2.08 $X2=1.2
+ $Y2=1.955
r132 1 3 99.292 $w=2.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.2 $Y=2.08 $X2=1.2
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_LP%B 3 5 6 7 9 10 11 15 19 20 22 24 25 27 31 33
+ 34 37 39
c86 15 0 1.96367e-20 $X=2.155 $Y=0.55
r87 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=1.345
+ $X2=2.455 $Y2=1.51
r88 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.455
+ $Y=1.345 $X2=2.455 $Y2=1.345
r89 34 38 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=1.345
+ $X2=2.455 $Y2=1.345
r90 25 27 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.825 $Y=1.985
+ $X2=2.825 $Y2=2.56
r91 22 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.545 $Y=0.835
+ $X2=2.545 $Y2=0.91
r92 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.545 $Y=0.835
+ $X2=2.545 $Y2=0.55
r93 21 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.44 $Y=1.91
+ $X2=2.365 $Y2=1.91
r94 20 25 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=2.7 $Y=1.91
+ $X2=2.825 $Y2=1.985
r95 20 21 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.7 $Y=1.91 $X2=2.44
+ $Y2=1.91
r96 19 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.365 $Y=1.835
+ $X2=2.365 $Y2=1.91
r97 19 39 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.365 $Y=1.835
+ $X2=2.365 $Y2=1.51
r98 16 31 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.455 $Y=0.91
+ $X2=2.545 $Y2=0.91
r99 16 28 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.455 $Y=0.91 $X2=2.155
+ $Y2=0.91
r100 16 37 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.455 $Y=0.985
+ $X2=2.455 $Y2=1.345
r101 13 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.155 $Y=0.835
+ $X2=2.155 $Y2=0.91
r102 13 15 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.155 $Y=0.835
+ $X2=2.155 $Y2=0.55
r103 12 15 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.155 $Y=0.255
+ $X2=2.155 $Y2=0.55
r104 10 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.29 $Y=1.91
+ $X2=2.365 $Y2=1.91
r105 10 11 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.29 $Y=1.91
+ $X2=1.855 $Y2=1.91
r106 7 11 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=1.73 $Y=1.985
+ $X2=1.855 $Y2=1.91
r107 7 9 117.608 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.595
r108 5 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.08 $Y=0.18
+ $X2=2.155 $Y2=0.255
r109 5 6 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.08 $Y=0.18 $X2=1.36
+ $Y2=0.18
r110 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.285 $Y=0.255
+ $X2=1.36 $Y2=0.18
r111 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.285 $Y=0.255
+ $X2=1.285 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_LP%X 1 2 7 8 10 15 17 18 19 20 31
c44 15 0 1.94535e-19 $X=1.07 $Y=0.805
c45 7 0 5.85314e-20 $X=0.735 $Y=1.3
r46 32 41 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=0.34 $Y=2.29 $X2=0.34
+ $Y2=2.24
r47 31 39 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=0.24 $Y=2.035 $X2=0.24
+ $Y2=2.075
r48 19 20 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.34 $Y=2.405
+ $X2=0.34 $Y2=2.775
r49 19 32 3.08211 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.34 $Y=2.405
+ $X2=0.34 $Y2=2.29
r50 18 41 3.83254 $w=4.28e-07 $l=1.43e-07 $layer=LI1_cond $X=0.34 $Y=2.097
+ $X2=0.34 $Y2=2.24
r51 18 39 3.06767 $w=4.28e-07 $l=2.2e-08 $layer=LI1_cond $X=0.34 $Y=2.097
+ $X2=0.34 $Y2=2.075
r52 18 31 1.15244 $w=2.28e-07 $l=2.3e-08 $layer=LI1_cond $X=0.24 $Y=2.012
+ $X2=0.24 $Y2=2.035
r53 17 18 17.3869 $w=2.28e-07 $l=3.47e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.012
r54 12 15 6.50043 $w=4.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.82 $Y=0.805
+ $X2=1.07 $Y2=0.805
r55 11 17 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=1.385
+ $X2=0.24 $Y2=1.665
r56 9 12 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.82 $Y=1.035 $X2=0.82
+ $Y2=0.805
r57 9 10 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.82 $Y=1.035
+ $X2=0.82 $Y2=1.215
r58 8 11 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.3
+ $X2=0.24 $Y2=1.385
r59 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.735 $Y=1.3
+ $X2=0.82 $Y2=1.215
r60 7 8 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.735 $Y=1.3 $X2=0.355
+ $Y2=1.3
r61 2 41 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=2.095 $X2=0.39 $Y2=2.24
r62 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.595 $X2=1.07 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_LP%A_159_419# 1 2 9 14 16
r30 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=2.475
+ $X2=0.935 $Y2=2.475
r31 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=2.475
+ $X2=1.995 $Y2=2.475
r32 9 10 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.83 $Y=2.475 $X2=1.1
+ $Y2=2.475
r33 2 16 300 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_PDIFF $count=2 $X=1.855
+ $Y=2.095 $X2=1.995 $Y2=2.555
r34 1 14 300 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_PDIFF $count=2 $X=0.795
+ $Y=2.095 $X2=0.935 $Y2=2.555
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_LP%VPWR 1 2 9 11 13 16 17 18 27 36
r43 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 33 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 27 35 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.612 $Y2=3.33
r49 27 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 26 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 21 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 18 33 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 18 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 16 25 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.465 $Y2=3.33
r59 15 29 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.63 $Y=3.33 $X2=1.68
+ $Y2=3.33
r60 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=3.33
+ $X2=1.465 $Y2=3.33
r61 11 35 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.612 $Y2=3.33
r62 11 13 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.55 $Y2=2.555
r63 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=3.245
+ $X2=1.465 $Y2=3.33
r64 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.465 $Y=3.245
+ $X2=1.465 $Y2=2.925
r65 2 13 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=3.41
+ $Y=2.06 $X2=3.55 $Y2=2.555
r66 1 9 600 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=2.095 $X2=1.465 $Y2=2.925
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_LP%VGND 1 2 3 10 12 16 18 20 23 24 25 34 46
r48 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r49 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 40 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r51 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r53 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r54 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r55 34 45 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.612
+ $Y2=0
r56 34 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.12
+ $Y2=0
r57 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r59 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r60 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r61 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r62 27 42 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r63 27 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r64 25 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r65 25 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r66 23 32 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.68
+ $Y2=0
r67 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.94
+ $Y2=0
r68 22 36 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.16
+ $Y2=0
r69 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=1.94
+ $Y2=0
r70 18 45 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.612 $Y2=0
r71 18 20 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.55 $Y=0.085 $X2=3.55
+ $Y2=0.485
r72 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r73 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.55
r74 10 42 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r75 10 12 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.805
r76 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.34 $X2=3.55 $Y2=0.485
r77 2 16 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.595 $X2=1.94 $Y2=0.55
r78 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.595 $X2=0.28 $Y2=0.805
.ends

