* File: sky130_fd_sc_lp__dlxbp_lp2.pex.spice
* Created: Fri Aug 28 10:28:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%D 3 7 11 15 17 18 19 23
c37 18 0 7.01416e-20 $X=0.72 $Y=1.295
r38 18 19 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.67 $Y=1.275
+ $X2=0.67 $Y2=1.665
r39 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.275 $X2=0.67 $Y2=1.275
r40 16 23 29.5381 $w=4.8e-07 $l=2.65e-07 $layer=POLY_cond $X=0.69 $Y=1.54
+ $X2=0.69 $Y2=1.275
r41 16 17 38.9835 $w=4.8e-07 $l=2.4e-07 $layer=POLY_cond $X=0.69 $Y=1.54
+ $X2=0.69 $Y2=1.78
r42 15 23 1.67197 $w=4.8e-07 $l=1.5e-08 $layer=POLY_cond $X=0.69 $Y=1.26
+ $X2=0.69 $Y2=1.275
r43 7 17 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.575 $Y=2.545
+ $X2=0.575 $Y2=1.78
r44 1 15 24.2025 $w=4.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=1.11
+ $X2=0.675 $Y2=1.26
r45 1 11 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.855 $Y=1.11
+ $X2=0.855 $Y2=0.495
r46 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.495 $Y=1.11
+ $X2=0.495 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%GATE 3 7 11 13 14 22
c50 7 0 7.01416e-20 $X=1.315 $Y=0.495
r51 20 22 4.39203 $w=6.7e-07 $l=5.5e-08 $layer=POLY_cond $X=1.675 $Y=1.51
+ $X2=1.73 $Y2=1.51
r52 19 20 28.7479 $w=6.7e-07 $l=3.6e-07 $layer=POLY_cond $X=1.315 $Y=1.51
+ $X2=1.675 $Y2=1.51
r53 17 19 3.99276 $w=6.7e-07 $l=5e-08 $layer=POLY_cond $X=1.265 $Y=1.51
+ $X2=1.315 $Y2=1.51
r54 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.665
r55 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.34 $X2=1.73 $Y2=1.34
r56 9 20 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.675 $Y=1.175
+ $X2=1.675 $Y2=1.51
r57 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.675 $Y=1.175
+ $X2=1.675 $Y2=0.495
r58 5 19 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.315 $Y=1.175
+ $X2=1.315 $Y2=1.51
r59 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.315 $Y=1.175
+ $X2=1.315 $Y2=0.495
r60 1 17 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.265 $Y=1.845
+ $X2=1.265 $Y2=1.51
r61 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.265 $Y=1.845 $X2=1.265
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%A_278_409# 1 2 9 13 17 21 25 28 29 30 31
+ 35 37 38 41 42 48 57
r129 53 55 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.665 $Y=1.33
+ $X2=2.85 $Y2=1.33
r130 51 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.935 $Y=1.33
+ $X2=3.025 $Y2=1.33
r131 51 55 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=2.935 $Y=1.33
+ $X2=2.85 $Y2=1.33
r132 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.935
+ $Y=1.33 $X2=2.935 $Y2=1.33
r133 47 48 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=2.19
+ $X2=1.695 $Y2=2.19
r134 44 47 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.3 $Y=2.19
+ $X2=1.53 $Y2=2.19
r135 42 59 7.77419 $w=2.48e-07 $l=4e-08 $layer=POLY_cond $X=3.99 $Y=1.59
+ $X2=3.95 $Y2=1.59
r136 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.99
+ $Y=1.59 $X2=3.99 $Y2=1.59
r137 39 50 12.2471 $w=2.59e-07 $l=2.6e-07 $layer=LI1_cond $X=2.935 $Y=1.59
+ $X2=2.935 $Y2=1.33
r138 39 41 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=3.1 $Y=1.59 $X2=3.99
+ $Y2=1.59
r139 37 39 9.21269 $w=2.59e-07 $l=2.0106e-07 $layer=LI1_cond $X=3.015 $Y=1.755
+ $X2=2.935 $Y2=1.59
r140 37 38 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.015 $Y=1.755
+ $X2=3.015 $Y2=2.185
r141 33 35 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.89 $Y=0.825
+ $X2=1.89 $Y2=0.495
r142 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.93 $Y=2.27
+ $X2=3.015 $Y2=2.185
r143 31 48 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.93 $Y=2.27
+ $X2=1.695 $Y2=2.27
r144 29 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.89 $Y2=0.825
r145 29 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.385 $Y2=0.91
r146 28 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=2.025
+ $X2=1.3 $Y2=2.19
r147 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.3 $Y=0.995
+ $X2=1.385 $Y2=0.91
r148 27 28 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=1.3 $Y=0.995
+ $X2=1.3 $Y2=2.025
r149 23 42 70.9395 $w=2.48e-07 $l=4.39829e-07 $layer=POLY_cond $X=4.355 $Y=1.425
+ $X2=3.99 $Y2=1.59
r150 23 25 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.355 $Y=1.425
+ $X2=4.355 $Y2=0.485
r151 19 59 2.63694 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.755
+ $X2=3.95 $Y2=1.59
r152 19 21 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.95 $Y=1.755
+ $X2=3.95 $Y2=2.465
r153 15 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.025 $Y=1.165
+ $X2=3.025 $Y2=1.33
r154 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.025 $Y=1.165
+ $X2=3.025 $Y2=0.485
r155 11 55 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.495
+ $X2=2.85 $Y2=1.33
r156 11 13 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.85 $Y=1.495
+ $X2=2.85 $Y2=2.195
r157 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.165
+ $X2=2.665 $Y2=1.33
r158 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.665 $Y=1.165
+ $X2=2.665 $Y2=0.485
r159 2 47 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.39
+ $Y=2.045 $X2=1.53 $Y2=2.19
r160 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.285 $X2=1.89 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%A_27_57# 1 2 7 12 13 15 20 21 25 26 29 33
+ 34 35
c73 15 0 5.80817e-20 $X=3.455 $Y=0.485
r74 35 37 8.96345 $w=3.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.295 $Y=2.62
+ $X2=0.295 $Y2=2.9
r75 33 34 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.295 $Y=2.19
+ $X2=0.295 $Y2=2.025
r76 31 34 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=0.2 $Y=0.725 $X2=0.2
+ $Y2=2.025
r77 29 31 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.28 $Y=0.495
+ $X2=0.28 $Y2=0.725
r78 26 41 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=2.115 $Y=2.9
+ $X2=2.115 $Y2=3.14
r79 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=2.9 $X2=2.115 $Y2=2.9
r80 23 25 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.115 $Y=2.705
+ $X2=2.115 $Y2=2.9
r81 22 35 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.475 $Y=2.62
+ $X2=0.295 $Y2=2.62
r82 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.95 $Y=2.62
+ $X2=2.115 $Y2=2.705
r83 21 22 96.2299 $w=1.68e-07 $l=1.475e-06 $layer=LI1_cond $X=1.95 $Y=2.62
+ $X2=0.475 $Y2=2.62
r84 20 35 2.72105 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.295 $Y=2.535
+ $X2=0.295 $Y2=2.62
r85 19 33 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.295 $Y=2.205
+ $X2=0.295 $Y2=2.19
r86 19 20 10.5641 $w=3.58e-07 $l=3.3e-07 $layer=LI1_cond $X=0.295 $Y=2.205
+ $X2=0.295 $Y2=2.535
r87 13 15 679.415 $w=1.5e-07 $l=1.325e-06 $layer=POLY_cond $X=3.455 $Y=1.81
+ $X2=3.455 $Y2=0.485
r88 10 12 149.072 $w=2.5e-07 $l=6e-07 $layer=POLY_cond $X=3.46 $Y=3.065 $X2=3.46
+ $Y2=2.465
r89 9 13 29.876 $w=2.42e-07 $l=1.5248e-07 $layer=POLY_cond $X=3.46 $Y=1.96
+ $X2=3.455 $Y2=1.81
r90 9 12 125.469 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.46 $Y=1.96
+ $X2=3.46 $Y2=2.465
r91 8 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=3.14
+ $X2=2.115 $Y2=3.14
r92 7 10 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.335 $Y=3.14
+ $X2=3.46 $Y2=3.065
r93 7 8 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=3.335 $Y=3.14
+ $X2=2.28 $Y2=3.14
r94 2 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.045 $X2=0.31 $Y2=2.9
r95 2 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.045 $X2=0.31 $Y2=2.19
r96 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%A_461_55# 1 2 9 12 16 19 22 25 26 28 29 33
+ 35 36 39 41
c98 36 0 2.47412e-20 $X=4.42 $Y=1.64
c99 33 0 5.80817e-20 $X=2.585 $Y=1.84
r100 39 45 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.64
+ $X2=4.805 $Y2=1.805
r101 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.805
+ $Y=1.64 $X2=4.805 $Y2=1.64
r102 36 38 18.7131 $w=2.51e-07 $l=3.85e-07 $layer=LI1_cond $X=4.42 $Y=1.64
+ $X2=4.805 $Y2=1.64
r103 30 33 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.37 $Y=1.84
+ $X2=2.585 $Y2=1.84
r104 28 36 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=1.475
+ $X2=4.42 $Y2=1.64
r105 27 28 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.42 $Y=1.145
+ $X2=4.42 $Y2=1.475
r106 26 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.905 $Y=0.98
+ $X2=3.905 $Y2=0.815
r107 25 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=0.98
+ $X2=3.74 $Y2=0.98
r108 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.905
+ $Y=0.98 $X2=3.905 $Y2=0.98
r109 22 27 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.335 $Y=0.98
+ $X2=4.42 $Y2=1.145
r110 22 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.335 $Y=0.98
+ $X2=3.905 $Y2=0.98
r111 21 29 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0.9
+ $X2=2.45 $Y2=0.9
r112 21 35 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=2.615 $Y=0.9
+ $X2=3.74 $Y2=0.9
r113 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=1.675
+ $X2=2.37 $Y2=1.84
r114 18 29 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.37 $Y=0.985
+ $X2=2.45 $Y2=0.9
r115 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.37 $Y=0.985
+ $X2=2.37 $Y2=1.675
r116 14 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.815
+ $X2=2.45 $Y2=0.9
r117 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.45 $Y=0.815
+ $X2=2.45 $Y2=0.49
r118 12 45 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.765 $Y=2.465
+ $X2=4.765 $Y2=1.805
r119 9 41 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.845 $Y=0.485
+ $X2=3.845 $Y2=0.815
r120 2 33 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.695 $X2=2.585 $Y2=1.84
r121 1 16 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.275 $X2=2.45 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%A_934_29# 1 2 7 9 10 11 13 16 20 22 23 26
+ 30 34 38 42 52 54 56 58 60 62 69 70 72 73
c153 54 0 1.99266e-19 $X=6.275 $Y=1.72
c154 10 0 2.47412e-20 $X=5.21 $Y=0.845
r155 83 85 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=5.285 $Y=1.64
+ $X2=5.335 $Y2=1.64
r156 73 85 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=5.645 $Y=1.64
+ $X2=5.335 $Y2=1.64
r157 72 75 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=5.65 $Y=1.64 $X2=5.65
+ $Y2=1.72
r158 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.645
+ $Y=1.64 $X2=5.645 $Y2=1.64
r159 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.755
+ $Y=1.06 $X2=6.755 $Y2=1.06
r160 67 69 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.755 $Y=1.4
+ $X2=6.755 $Y2=1.06
r161 66 69 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.755 $Y=0.945
+ $X2=6.755 $Y2=1.06
r162 62 64 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.44 $Y=2.11
+ $X2=6.44 $Y2=2.82
r163 60 67 16.7087 $w=2.3e-07 $l=4.03943e-07 $layer=LI1_cond $X=6.44 $Y=1.805
+ $X2=6.755 $Y2=1.602
r164 60 62 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.44 $Y=1.805
+ $X2=6.44 $Y2=2.11
r165 56 66 37.4414 $w=1.45e-07 $l=4.45e-07 $layer=LI1_cond $X=6.31 $Y=0.86
+ $X2=6.755 $Y2=0.86
r166 56 58 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.31 $Y=0.775
+ $X2=6.31 $Y2=0.49
r167 55 75 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.81 $Y=1.72
+ $X2=5.65 $Y2=1.72
r168 54 60 9.60724 $w=2.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.275 $Y=1.72
+ $X2=6.44 $Y2=1.805
r169 54 55 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.275 $Y=1.72
+ $X2=5.81 $Y2=1.72
r170 45 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.755 $Y=1.045
+ $X2=6.755 $Y2=1.06
r171 45 47 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.755 $Y=0.97
+ $X2=7.085 $Y2=0.97
r172 40 52 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.235 $Y=0.895
+ $X2=8.235 $Y2=0.97
r173 40 42 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=8.235 $Y=0.895
+ $X2=8.235 $Y2=0.495
r174 36 52 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=8.185 $Y=0.97
+ $X2=8.235 $Y2=0.97
r175 36 50 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=8.185 $Y=0.97
+ $X2=7.875 $Y2=0.97
r176 36 38 320.505 $w=2.5e-07 $l=1.29e-06 $layer=POLY_cond $X=8.185 $Y=1.045
+ $X2=8.185 $Y2=2.335
r177 32 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.875 $Y=0.895
+ $X2=7.875 $Y2=0.97
r178 32 34 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.875 $Y=0.895
+ $X2=7.875 $Y2=0.495
r179 28 50 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=7.655 $Y=0.97
+ $X2=7.875 $Y2=0.97
r180 28 48 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.655 $Y=0.97
+ $X2=7.445 $Y2=0.97
r181 28 30 320.505 $w=2.5e-07 $l=1.29e-06 $layer=POLY_cond $X=7.655 $Y=1.045
+ $X2=7.655 $Y2=2.335
r182 24 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.445 $Y=0.895
+ $X2=7.445 $Y2=0.97
r183 24 26 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.445 $Y=0.895
+ $X2=7.445 $Y2=0.495
r184 23 47 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.16 $Y=0.97
+ $X2=7.085 $Y2=0.97
r185 22 48 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.37 $Y=0.97
+ $X2=7.445 $Y2=0.97
r186 22 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.37 $Y=0.97
+ $X2=7.16 $Y2=0.97
r187 18 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.085 $Y=0.895
+ $X2=7.085 $Y2=0.97
r188 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.085 $Y=0.895
+ $X2=7.085 $Y2=0.495
r189 14 85 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.335 $Y=1.805
+ $X2=5.335 $Y2=1.64
r190 14 16 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.335 $Y=1.805
+ $X2=5.335 $Y2=2.465
r191 13 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.475
+ $X2=5.285 $Y2=1.64
r192 12 13 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.285 $Y=0.92
+ $X2=5.285 $Y2=1.475
r193 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.21 $Y=0.845
+ $X2=5.285 $Y2=0.92
r194 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=5.21 $Y=0.845
+ $X2=4.82 $Y2=0.845
r195 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.745 $Y=0.77
+ $X2=4.82 $Y2=0.845
r196 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.745 $Y=0.77
+ $X2=4.745 $Y2=0.485
r197 2 64 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.965 $X2=6.44 $Y2=2.82
r198 2 62 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.965 $X2=6.44 $Y2=2.11
r199 1 58 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.17
+ $Y=0.275 $X2=6.31 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%A_784_55# 1 2 7 9 10 11 12 14 19 21 22 26
+ 28 30 33 34 35 37 38 42 43 47 50
c113 47 0 1.99266e-19 $X=6.185 $Y=1.29
r114 47 51 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.185 $Y=1.29
+ $X2=6.185 $Y2=1.455
r115 47 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.185 $Y=1.29
+ $X2=6.185 $Y2=1.125
r116 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.185
+ $Y=1.29 $X2=6.185 $Y2=1.29
r117 43 46 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.185 $Y=1.21
+ $X2=6.185 $Y2=1.29
r118 39 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=1.21
+ $X2=5.225 $Y2=1.21
r119 38 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.02 $Y=1.21
+ $X2=6.185 $Y2=1.21
r120 38 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.02 $Y=1.21
+ $X2=5.31 $Y2=1.21
r121 36 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=1.295
+ $X2=5.225 $Y2=1.21
r122 36 37 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=5.225 $Y=1.295
+ $X2=5.225 $Y2=2.815
r123 34 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=1.21
+ $X2=5.225 $Y2=1.21
r124 34 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.14 $Y=1.21
+ $X2=4.855 $Y2=1.21
r125 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.77 $Y=1.125
+ $X2=4.855 $Y2=1.21
r126 32 33 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.77 $Y=0.635
+ $X2=4.77 $Y2=1.125
r127 31 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=2.9
+ $X2=4.295 $Y2=2.9
r128 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=2.9
+ $X2=5.225 $Y2=2.815
r129 30 31 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.14 $Y=2.9
+ $X2=4.46 $Y2=2.9
r130 26 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=2.815
+ $X2=4.295 $Y2=2.9
r131 26 28 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=4.295 $Y=2.815
+ $X2=4.295 $Y2=2.11
r132 22 32 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.685 $Y=0.485
+ $X2=4.77 $Y2=0.635
r133 22 24 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=4.685 $Y=0.485
+ $X2=4.14 $Y2=0.485
r134 19 51 250.938 $w=2.5e-07 $l=1.01e-06 $layer=POLY_cond $X=6.175 $Y=2.465
+ $X2=6.175 $Y2=1.455
r135 15 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.095 $Y=0.92
+ $X2=6.095 $Y2=0.845
r136 15 50 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=6.095 $Y=0.92
+ $X2=6.095 $Y2=1.125
r137 12 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.095 $Y=0.77
+ $X2=6.095 $Y2=0.845
r138 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.095 $Y=0.77
+ $X2=6.095 $Y2=0.485
r139 10 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.02 $Y=0.845
+ $X2=6.095 $Y2=0.845
r140 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.02 $Y=0.845
+ $X2=5.81 $Y2=0.845
r141 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.735 $Y=0.77
+ $X2=5.81 $Y2=0.845
r142 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.735 $Y=0.77
+ $X2=5.735 $Y2=0.485
r143 2 41 400 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=4.075
+ $Y=1.965 $X2=4.295 $Y2=2.82
r144 2 28 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=4.075
+ $Y=1.965 $X2=4.295 $Y2=2.11
r145 1 24 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.275 $X2=4.14 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%A_1662_57# 1 2 9 13 17 21 25 29 33 36 39
r50 38 39 4.82966 $w=4.99e-07 $l=5e-08 $layer=POLY_cond $X=9.225 $Y=1.425
+ $X2=9.275 $Y2=1.425
r51 34 38 18.8357 $w=4.99e-07 $l=1.95e-07 $layer=POLY_cond $X=9.03 $Y=1.425
+ $X2=9.225 $Y2=1.425
r52 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.03
+ $Y=1.255 $X2=9.03 $Y2=1.255
r53 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.03 $Y=1.59
+ $X2=9.03 $Y2=1.255
r54 30 36 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=1.675
+ $X2=8.45 $Y2=1.675
r55 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.865 $Y=1.675
+ $X2=9.03 $Y2=1.59
r56 29 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.865 $Y=1.675
+ $X2=8.615 $Y2=1.675
r57 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.45 $Y=1.98 $X2=8.45
+ $Y2=2.69
r58 23 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=1.76 $X2=8.45
+ $Y2=1.675
r59 23 25 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=8.45 $Y=1.76
+ $X2=8.45 $Y2=1.98
r60 19 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=1.59 $X2=8.45
+ $Y2=1.675
r61 19 21 38.2402 $w=3.28e-07 $l=1.095e-06 $layer=LI1_cond $X=8.45 $Y=1.59
+ $X2=8.45 $Y2=0.495
r62 15 39 29.9439 $w=4.99e-07 $l=4.64839e-07 $layer=POLY_cond $X=9.585 $Y=1.09
+ $X2=9.275 $Y2=1.425
r63 15 17 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=9.585 $Y=1.09
+ $X2=9.585 $Y2=0.67
r64 11 39 18.9214 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.275 $Y=1.76
+ $X2=9.275 $Y2=1.425
r65 11 13 195.036 $w=2.5e-07 $l=7.85e-07 $layer=POLY_cond $X=9.275 $Y=1.76
+ $X2=9.275 $Y2=2.545
r66 7 38 31.3575 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.225 $Y=1.09
+ $X2=9.225 $Y2=1.425
r67 7 9 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=9.225 $Y=1.09
+ $X2=9.225 $Y2=0.67
r68 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.31
+ $Y=1.835 $X2=8.45 $Y2=2.69
r69 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.31
+ $Y=1.835 $X2=8.45 $Y2=1.98
r70 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.31
+ $Y=0.285 $X2=8.45 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%VPWR 1 2 3 4 5 18 22 26 30 34 38 43 44 45
+ 51 58 63 73 74 77 80 83 86
r90 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r91 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r92 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r93 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r94 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r95 74 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r96 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r97 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=3.33
+ $X2=9.01 $Y2=3.33
r98 71 73 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=9.175 $Y=3.33
+ $X2=9.84 $Y2=3.33
r99 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r100 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r101 67 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r102 67 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r103 66 69 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r104 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r105 64 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=3.33
+ $X2=5.655 $Y2=3.33
r106 64 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.82 $Y=3.33 $X2=6
+ $Y2=3.33
r107 63 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 63 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.44 $Y2=3.33
r109 62 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r111 59 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=3.33
+ $X2=3.195 $Y2=3.33
r112 59 61 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 58 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.655 $Y2=3.33
r114 58 61 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 57 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 54 57 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 53 56 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 51 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=3.33
+ $X2=3.195 $Y2=3.33
r121 51 56 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.03 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 49 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 45 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r125 45 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r126 43 48 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.92 $Y2=3.33
r128 42 53 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.92 $Y2=3.33
r130 38 41 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.01 $Y=2.19
+ $X2=9.01 $Y2=2.9
r131 36 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=3.245
+ $X2=9.01 $Y2=3.33
r132 36 41 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=9.01 $Y=3.245
+ $X2=9.01 $Y2=2.9
r133 35 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 34 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=9.01 $Y2=3.33
r135 34 35 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=8.085 $Y2=3.33
r136 30 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.92 $Y=1.98
+ $X2=7.92 $Y2=2.69
r137 28 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r138 28 33 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.69
r139 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=3.33
r140 24 26 38.2402 $w=3.28e-07 $l=1.095e-06 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=2.15
r141 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=3.245
+ $X2=3.195 $Y2=3.33
r142 20 22 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.195 $Y=3.245
+ $X2=3.195 $Y2=2.76
r143 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=3.33
r144 16 18 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=3.05
r145 5 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.865
+ $Y=2.045 $X2=9.01 $Y2=2.9
r146 5 38 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.865
+ $Y=2.045 $X2=9.01 $Y2=2.19
r147 4 33 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.835 $X2=7.92 $Y2=2.69
r148 4 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.835 $X2=7.92 $Y2=1.98
r149 3 26 300 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_PDIFF $count=2 $X=5.46
+ $Y=1.965 $X2=5.655 $Y2=2.15
r150 2 22 600 $w=1.7e-07 $l=1.16984e-06 $layer=licon1_PDIFF $count=1 $X=2.975
+ $Y=1.695 $X2=3.195 $Y2=2.76
r151 1 18 600 $w=1.7e-07 $l=1.10956e-06 $layer=licon1_PDIFF $count=1 $X=0.7
+ $Y=2.045 $X2=0.92 $Y2=3.05
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%Q 1 2 7 13 14 15 16 17 36
r39 16 17 7.49192 $w=4.53e-07 $l=2.85e-07 $layer=LI1_cond $X=7.327 $Y=2.405
+ $X2=7.327 $Y2=2.69
r40 15 16 11.1722 $w=4.53e-07 $l=4.25e-07 $layer=LI1_cond $X=7.327 $Y=1.98
+ $X2=7.327 $Y2=2.405
r41 14 15 8.28054 $w=4.53e-07 $l=3.15e-07 $layer=LI1_cond $X=7.327 $Y=1.665
+ $X2=7.327 $Y2=1.98
r42 14 23 6.78216 $w=4.53e-07 $l=2.58e-07 $layer=LI1_cond $X=7.327 $Y=1.665
+ $X2=7.327 $Y2=1.407
r43 13 23 2.94419 $w=4.53e-07 $l=1.12e-07 $layer=LI1_cond $X=7.327 $Y=1.295
+ $X2=7.327 $Y2=1.407
r44 13 36 7.93754 $w=4.53e-07 $l=1.15e-07 $layer=LI1_cond $X=7.327 $Y=1.295
+ $X2=7.327 $Y2=1.18
r45 11 36 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.185 $Y=0.595
+ $X2=7.185 $Y2=1.18
r46 7 11 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.1 $Y=0.43
+ $X2=7.185 $Y2=0.595
r47 7 9 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=7.1 $Y=0.43 $X2=6.87
+ $Y2=0.43
r48 2 17 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.835 $X2=7.39 $Y2=2.69
r49 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.835 $X2=7.39 $Y2=1.98
r50 1 9 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.725
+ $Y=0.285 $X2=6.87 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%Q_N 1 2 7 8 9 10 11 12 13 36
r15 22 36 2.1185 $w=5.46e-07 $l=1.34907e-07 $layer=LI1_cond $X=9.8 $Y=2.025
+ $X2=9.67 $Y2=2.035
r16 13 45 2.79304 $w=5.46e-07 $l=1.25e-07 $layer=LI1_cond $X=9.67 $Y=2.775
+ $X2=9.67 $Y2=2.9
r17 12 13 8.2674 $w=5.46e-07 $l=3.7e-07 $layer=LI1_cond $X=9.67 $Y=2.405
+ $X2=9.67 $Y2=2.775
r18 12 39 4.80403 $w=5.46e-07 $l=2.15e-07 $layer=LI1_cond $X=9.67 $Y=2.405
+ $X2=9.67 $Y2=2.19
r19 11 39 2.63663 $w=5.46e-07 $l=1.18e-07 $layer=LI1_cond $X=9.67 $Y=2.072
+ $X2=9.67 $Y2=2.19
r20 11 36 0.82674 $w=5.46e-07 $l=3.7e-08 $layer=LI1_cond $X=9.67 $Y=2.072
+ $X2=9.67 $Y2=2.035
r21 11 22 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=9.8 $Y=1.987 $X2=9.8
+ $Y2=2.025
r22 10 11 11.245 $w=3.28e-07 $l=3.22e-07 $layer=LI1_cond $X=9.8 $Y=1.665 $X2=9.8
+ $Y2=1.987
r23 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.8 $Y=1.295 $X2=9.8
+ $Y2=1.665
r24 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.8 $Y=0.925 $X2=9.8
+ $Y2=1.295
r25 8 27 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.8 $Y=0.925 $X2=9.8
+ $Y2=0.67
r26 7 27 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=9.8 $Y=0.555 $X2=9.8
+ $Y2=0.67
r27 2 45 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.4
+ $Y=2.045 $X2=9.54 $Y2=2.9
r28 2 39 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.4
+ $Y=2.045 $X2=9.54 $Y2=2.19
r29 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.46 $X2=9.8 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBP_LP2%VGND 1 2 3 4 5 18 20 24 28 32 36 39 40 41
+ 43 48 60 66 67 70 73 76 79
r113 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r114 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r115 71 74 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r116 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 67 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=8.88
+ $Y2=0
r118 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r119 64 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.01
+ $Y2=0
r120 64 66 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.84
+ $Y2=0
r121 63 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r122 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r123 60 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=0 $X2=9.01
+ $Y2=0
r124 60 62 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=8.845 $Y=0
+ $X2=7.92 $Y2=0
r125 59 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r126 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r127 56 59 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=7.44 $Y2=0
r128 55 58 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r129 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r130 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=0 $X2=5.2
+ $Y2=0
r131 53 55 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.365 $Y=0
+ $X2=5.52 $Y2=0
r132 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r133 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r134 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.24
+ $Y2=0
r135 49 51 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.6
+ $Y2=0
r136 48 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.2
+ $Y2=0
r137 48 51 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=5.035 $Y=0
+ $X2=3.6 $Y2=0
r138 46 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r139 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r140 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r141 43 45 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r142 41 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r143 41 52 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r144 41 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r145 39 58 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.495 $Y=0 $X2=7.44
+ $Y2=0
r146 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.495 $Y=0 $X2=7.66
+ $Y2=0
r147 38 62 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.825 $Y=0 $X2=7.92
+ $Y2=0
r148 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=0 $X2=7.66
+ $Y2=0
r149 34 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0
r150 34 36 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0.67
r151 30 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.66 $Y=0.085
+ $X2=7.66 $Y2=0
r152 30 32 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.66 $Y=0.085
+ $X2=7.66 $Y2=0.495
r153 26 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.2 $Y=0.085 $X2=5.2
+ $Y2=0
r154 26 28 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.2 $Y=0.085 $X2=5.2
+ $Y2=0.485
r155 22 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=0.085
+ $X2=3.24 $Y2=0
r156 22 24 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.24 $Y=0.085 $X2=3.24
+ $Y2=0.485
r157 21 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r158 20 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=0 $X2=3.24
+ $Y2=0
r159 20 21 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.075 $Y=0
+ $X2=1.235 $Y2=0
r160 16 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r161 16 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.455
r162 5 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.865
+ $Y=0.46 $X2=9.01 $Y2=0.67
r163 4 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.52
+ $Y=0.285 $X2=7.66 $Y2=0.495
r164 3 28 182 $w=1.7e-07 $l=4.73498e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.275 $X2=5.2 $Y2=0.485
r165 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.1
+ $Y=0.275 $X2=3.24 $Y2=0.485
r166 1 18 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.285 $X2=1.07 $Y2=0.455
.ends

