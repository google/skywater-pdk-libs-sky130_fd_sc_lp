* File: sky130_fd_sc_lp__a211oi_2.pex.spice
* Created: Wed Sep  2 09:18:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211OI_2%C1 1 3 6 8 10 13 15 16 24
r41 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.545 $Y=1.375
+ $X2=0.975 $Y2=1.375
r42 20 23 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.34 $Y=1.375
+ $X2=0.545 $Y2=1.375
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.375 $X2=0.34 $Y2=1.375
r44 16 21 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.375
r45 15 21 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.375
r46 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.54
+ $X2=0.975 $Y2=1.375
r47 11 13 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.975 $Y=1.54
+ $X2=0.975 $Y2=2.465
r48 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.21
+ $X2=0.975 $Y2=1.375
r49 8 10 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.975 $Y=1.21
+ $X2=0.975 $Y2=0.665
r50 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.54
+ $X2=0.545 $Y2=1.375
r51 4 6 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.545 $Y=1.54
+ $X2=0.545 $Y2=2.465
r52 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.21
+ $X2=0.545 $Y2=1.375
r53 1 3 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.545 $Y=1.21
+ $X2=0.545 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%B1 3 7 11 15 17 18 26
c50 18 0 1.60609e-19 $X=1.68 $Y=1.665
r51 24 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.62 $Y=1.51
+ $X2=1.835 $Y2=1.51
r52 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.51 $X2=1.62 $Y2=1.51
r53 21 24 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.405 $Y=1.51
+ $X2=1.62 $Y2=1.51
r54 18 25 2.12759 $w=3.23e-07 $l=6e-08 $layer=LI1_cond $X=1.68 $Y=1.587 $X2=1.62
+ $Y2=1.587
r55 17 25 14.8931 $w=3.23e-07 $l=4.2e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.62 $Y2=1.587
r56 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.675
+ $X2=1.835 $Y2=1.51
r57 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.835 $Y=1.675
+ $X2=1.835 $Y2=2.465
r58 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.345
+ $X2=1.835 $Y2=1.51
r59 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.835 $Y=1.345
+ $X2=1.835 $Y2=0.665
r60 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.675
+ $X2=1.405 $Y2=1.51
r61 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.405 $Y=1.675
+ $X2=1.405 $Y2=2.465
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.345
+ $X2=1.405 $Y2=1.51
r63 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.405 $Y=1.345
+ $X2=1.405 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%A2 3 7 11 15 22 25 26 27 28 35
c56 35 0 1.60609e-19 $X=3.375 $Y=1.51
c57 15 0 1.51646e-19 $X=3.375 $Y=2.465
r58 27 28 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.582
+ $X2=2.64 $Y2=1.582
r59 25 28 3.02731 $w=3.33e-07 $l=8.8e-08 $layer=LI1_cond $X=2.728 $Y=1.582
+ $X2=2.64 $Y2=1.582
r60 25 26 8.1966 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=2.728 $Y=1.582
+ $X2=2.895 $Y2=1.582
r61 23 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.285 $Y=1.51
+ $X2=3.375 $Y2=1.51
r62 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.285
+ $Y=1.51 $X2=3.285 $Y2=1.51
r63 20 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.945 $Y=1.51
+ $X2=3.285 $Y2=1.51
r64 20 31 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.945 $Y=1.51
+ $X2=2.785 $Y2=1.51
r65 19 22 20.9495 $w=1.78e-07 $l=3.4e-07 $layer=LI1_cond $X=2.945 $Y=1.505
+ $X2=3.285 $Y2=1.505
r66 19 26 3.08081 $w=1.78e-07 $l=5e-08 $layer=LI1_cond $X=2.945 $Y=1.505
+ $X2=2.895 $Y2=1.505
r67 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.945
+ $Y=1.51 $X2=2.945 $Y2=1.51
r68 13 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.675
+ $X2=3.375 $Y2=1.51
r69 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.375 $Y=1.675
+ $X2=3.375 $Y2=2.465
r70 9 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.345
+ $X2=3.375 $Y2=1.51
r71 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.375 $Y=1.345 $X2=3.375
+ $Y2=0.745
r72 5 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=1.675
+ $X2=2.945 $Y2=1.51
r73 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.945 $Y=1.675
+ $X2=2.945 $Y2=2.465
r74 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.345
+ $X2=2.785 $Y2=1.51
r75 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.785 $Y=1.345 $X2=2.785
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%A1 1 3 6 10 12 14 15 20 21 27
r48 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.44 $X2=4.53 $Y2=1.44
r49 27 29 27.8575 $w=3.72e-07 $l=2.15e-07 $layer=POLY_cond $X=4.315 $Y=1.475
+ $X2=4.53 $Y2=1.475
r50 26 27 10.3656 $w=3.72e-07 $l=8e-08 $layer=POLY_cond $X=4.235 $Y=1.475
+ $X2=4.315 $Y2=1.475
r51 21 30 9.60369 $w=2.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.58 $Y=1.665
+ $X2=4.58 $Y2=1.44
r52 20 30 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.58 $Y=1.295
+ $X2=4.58 $Y2=1.44
r53 18 26 44.0538 $w=3.72e-07 $l=3.4e-07 $layer=POLY_cond $X=3.895 $Y=1.475
+ $X2=4.235 $Y2=1.475
r54 18 24 11.6613 $w=3.72e-07 $l=9e-08 $layer=POLY_cond $X=3.895 $Y=1.475
+ $X2=3.805 $Y2=1.475
r55 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.895
+ $Y=1.51 $X2=3.895 $Y2=1.51
r56 15 30 3.11056 $w=1.8e-07 $l=1.64317e-07 $layer=LI1_cond $X=4.445 $Y=1.505
+ $X2=4.58 $Y2=1.44
r57 15 17 33.8889 $w=1.78e-07 $l=5.5e-07 $layer=LI1_cond $X=4.445 $Y=1.505
+ $X2=3.895 $Y2=1.505
r58 12 27 24.0971 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=4.315 $Y=1.275
+ $X2=4.315 $Y2=1.475
r59 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.315 $Y=1.275
+ $X2=4.315 $Y2=0.745
r60 8 26 24.0971 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=4.235 $Y=1.675
+ $X2=4.235 $Y2=1.475
r61 8 10 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.235 $Y=1.675
+ $X2=4.235 $Y2=2.465
r62 4 24 24.0971 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.805 $Y=1.675
+ $X2=3.805 $Y2=1.475
r63 4 6 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.805 $Y=1.675
+ $X2=3.805 $Y2=2.465
r64 1 24 24.0971 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.805 $Y=1.275
+ $X2=3.805 $Y2=1.475
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.805 $Y=1.275
+ $X2=3.805 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%A_41_367# 1 2 3 10 12 14 18 20 24 29
r32 22 24 21.2759 $w=2.58e-07 $l=4.8e-07 $layer=LI1_cond $X=2.085 $Y=2.905
+ $X2=2.085 $Y2=2.425
r33 21 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.285 $Y=2.99
+ $X2=1.19 $Y2=2.99
r34 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=2.085 $Y2=2.905
r35 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=1.285 $Y2=2.99
r36 16 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=2.905
+ $X2=1.19 $Y2=2.99
r37 16 18 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=1.19 $Y=2.905
+ $X2=1.19 $Y2=2.085
r38 15 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.425 $Y=2.99
+ $X2=0.295 $Y2=2.99
r39 14 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=1.19 $Y2=2.99
r40 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=0.425 $Y2=2.99
r41 10 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.295 $Y=2.905
+ $X2=0.295 $Y2=2.99
r42 10 12 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.295 $Y=2.905
+ $X2=0.295 $Y2=2.085
r43 3 24 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.425
r44 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.91
r45 2 18 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.085
r46 1 27 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.91
r47 1 12 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%Y 1 2 3 4 15 19 23 25 29 31 33 34 35 39
r60 34 35 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=0.555
+ $X2=1.645 $Y2=0.925
r61 34 39 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.645 $Y=0.555
+ $X2=1.645 $Y2=0.42
r62 32 35 7.20277 $w=2.38e-07 $l=1.5e-07 $layer=LI1_cond $X=1.645 $Y=1.075
+ $X2=1.645 $Y2=0.925
r63 32 33 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.075
+ $X2=1.645 $Y2=1.16
r64 27 29 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.1 $Y=1.075
+ $X2=4.1 $Y2=0.68
r65 26 33 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.765 $Y=1.16
+ $X2=1.645 $Y2=1.16
r66 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.935 $Y=1.16
+ $X2=4.1 $Y2=1.075
r67 25 26 141.572 $w=1.68e-07 $l=2.17e-06 $layer=LI1_cond $X=3.935 $Y=1.16
+ $X2=1.765 $Y2=1.16
r68 24 31 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=1.16
+ $X2=0.76 $Y2=1.16
r69 23 33 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.525 $Y=1.16
+ $X2=1.645 $Y2=1.16
r70 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.525 $Y=1.16
+ $X2=0.925 $Y2=1.16
r71 19 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.76 $Y=1.97
+ $X2=0.76 $Y2=2.65
r72 17 31 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=1.245
+ $X2=0.76 $Y2=1.16
r73 17 19 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=0.76 $Y=1.245
+ $X2=0.76 $Y2=1.97
r74 13 31 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.725 $Y=1.075
+ $X2=0.76 $Y2=1.16
r75 13 15 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=0.725 $Y=1.075
+ $X2=0.725 $Y2=0.42
r76 4 21 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.65
r77 4 19 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=1.97
r78 3 29 91 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.325 $X2=4.1 $Y2=0.68
r79 2 39 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.48
+ $Y=0.245 $X2=1.62 $Y2=0.42
r80 1 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.62
+ $Y=0.245 $X2=0.76 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%A_296_367# 1 2 3 12 14 15 18 20 24 28
c41 28 0 1.51646e-19 $X=3.16 $Y=1.85
r42 31 32 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=3.16 $Y=1.98
+ $X2=3.16 $Y2=2.005
r43 28 31 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=3.16 $Y=1.85
+ $X2=3.16 $Y2=1.98
r44 24 26 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.02 $Y=1.98
+ $X2=4.02 $Y2=2.91
r45 22 24 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=4.02 $Y=1.935
+ $X2=4.02 $Y2=1.98
r46 21 28 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.255 $Y=1.85 $X2=3.16
+ $Y2=1.85
r47 20 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.925 $Y=1.85
+ $X2=4.02 $Y2=1.935
r48 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.925 $Y=1.85
+ $X2=3.255 $Y2=1.85
r49 16 32 4.96172 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=2.09
+ $X2=3.16 $Y2=2.005
r50 16 18 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=3.16 $Y=2.09
+ $X2=3.16 $Y2=2.455
r51 14 32 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.065 $Y=2.005 $X2=3.16
+ $Y2=2.005
r52 14 15 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=3.065 $Y=2.005
+ $X2=1.785 $Y2=2.005
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=2.09
+ $X2=1.785 $Y2=2.005
r54 10 12 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.62 $Y=2.09 $X2=1.62
+ $Y2=2.095
r55 3 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.835 $X2=4.02 $Y2=2.91
r56 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.835 $X2=4.02 $Y2=1.98
r57 2 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.835 $X2=3.16 $Y2=1.98
r58 2 18 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=3.02
+ $Y=1.835 $X2=3.16 $Y2=2.455
r59 1 12 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%VPWR 1 2 3 12 16 20 22 26 28 33 38 44 47 51
r64 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r65 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r66 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 42 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r68 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r70 39 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.59 $Y2=3.33
r71 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=4.08 $Y2=3.33
r72 38 50 4.59886 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.542 $Y2=3.33
r73 38 41 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.08 $Y2=3.33
r74 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r75 37 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r77 34 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.73 $Y2=3.33
r78 34 36 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 33 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.59 $Y2=3.33
r80 33 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.12 $Y2=3.33
r81 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r82 28 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.73 $Y2=3.33
r83 28 30 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 26 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r85 26 31 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 22 25 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=4.45 $Y=2.005
+ $X2=4.45 $Y2=2.95
r87 20 50 3.16731 $w=3.3e-07 $l=1.27609e-07 $layer=LI1_cond $X=4.45 $Y=3.245
+ $X2=4.542 $Y2=3.33
r88 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.45 $Y=3.245
+ $X2=4.45 $Y2=2.95
r89 16 19 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=3.59 $Y=2.19
+ $X2=3.59 $Y2=2.95
r90 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=3.33
r91 14 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=2.95
r92 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=3.33
r93 10 12 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=2.38
r94 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.835 $X2=4.45 $Y2=2.95
r95 3 22 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.835 $X2=4.45 $Y2=2.005
r96 2 19 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.835 $X2=3.59 $Y2=2.95
r97 2 16 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.835 $X2=3.59 $Y2=2.19
r98 1 12 300 $w=1.7e-07 $l=6.04276e-07 $layer=licon1_PDIFF $count=2 $X=2.605
+ $Y=1.835 $X2=2.73 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%VGND 1 2 3 4 13 15 19 23 27 30 31 32 34 43
+ 52 53 59 62
r66 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r67 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r69 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r70 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r71 50 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r72 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r73 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r74 47 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.08
+ $Y2=0
r75 47 49 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.6
+ $Y2=0
r76 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r77 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r78 43 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.08
+ $Y2=0
r79 43 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r80 42 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r81 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r82 39 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.19
+ $Y2=0
r83 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.68
+ $Y2=0
r84 38 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r85 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r86 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 35 56 4.03203 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r88 35 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r89 34 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.19
+ $Y2=0
r90 34 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.72
+ $Y2=0
r91 32 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r92 32 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r93 30 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.68
+ $Y2=0
r94 30 31 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.075
+ $Y2=0
r95 29 45 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.64
+ $Y2=0
r96 29 31 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.075
+ $Y2=0
r97 25 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r98 25 27 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.45
r99 21 31 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0
r100 21 23 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0.39
r101 17 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=0.085
+ $X2=1.19 $Y2=0
r102 17 19 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.19 $Y=0.085
+ $X2=1.19 $Y2=0.39
r103 13 56 3.18019 $w=2.6e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.212 $Y2=0
r104 13 15 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.39
r105 4 27 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.325 $X2=3.08 $Y2=0.45
r106 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.91
+ $Y=0.245 $X2=2.05 $Y2=0.39
r107 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.05
+ $Y=0.245 $X2=1.19 $Y2=0.39
r108 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.205
+ $Y=0.245 $X2=0.33 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_2%A_489_65# 1 2 3 12 14 15 19 20 21 24
r43 22 24 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=4.565 $Y=0.425
+ $X2=4.565 $Y2=0.47
r44 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.435 $Y=0.34
+ $X2=4.565 $Y2=0.425
r45 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.435 $Y=0.34
+ $X2=3.755 $Y2=0.34
r46 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.59 $Y=0.735
+ $X2=3.59 $Y2=0.45
r47 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.59 $Y=0.425
+ $X2=3.755 $Y2=0.34
r48 16 19 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.59 $Y=0.425
+ $X2=3.59 $Y2=0.45
r49 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.425 $Y=0.82
+ $X2=3.59 $Y2=0.735
r50 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.425 $Y=0.82
+ $X2=2.735 $Y2=0.82
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.57 $Y=0.735
+ $X2=2.735 $Y2=0.82
r52 10 12 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.57 $Y=0.735
+ $X2=2.57 $Y2=0.47
r53 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.39
+ $Y=0.325 $X2=4.53 $Y2=0.47
r54 2 19 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.45
+ $Y=0.325 $X2=3.59 $Y2=0.45
r55 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.325 $X2=2.57 $Y2=0.47
.ends

