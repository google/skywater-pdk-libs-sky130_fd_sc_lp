* File: sky130_fd_sc_lp__nand2b_1.spice
* Created: Fri Aug 28 10:47:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2b_1.pex.spice"
.subckt sky130_fd_sc_lp__nand2b_1  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_N_M1000_g N_A_40_367#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0854 AS=0.1113 PD=0.8 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1003 A_269_47# N_B_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.1708 PD=1.05 PS=1.6 NRD=7.14 NRS=11.424 M=1 R=5.6 SA=75000.4 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_A_40_367#_M1001_g A_269_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2856 AS=0.0882 PD=2.36 PS=1.05 NRD=4.992 NRS=7.14 M=1 R=5.6 SA=75000.8
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A_N_M1004_g N_A_40_367#_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=46.886 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.285075 PD=1.54 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_40_367#_M1005_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__nand2b_1.pxi.spice"
*
.ends
*
*
