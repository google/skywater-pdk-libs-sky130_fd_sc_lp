* File: sky130_fd_sc_lp__and4b_m.pex.spice
* Created: Fri Aug 28 10:08:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4B_M%A_N 3 5 6 7 9 12 13 16 17
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.14 $X2=0.385 $Y2=1.14
r40 13 17 3.40061 $w=5.08e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.31
+ $X2=0.385 $Y2=1.31
r41 12 16 100.545 $w=3.3e-07 $l=5.75e-07 $layer=POLY_cond $X=0.385 $Y=1.715
+ $X2=0.385 $Y2=1.14
r42 11 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=0.975
+ $X2=0.385 $Y2=1.14
r43 7 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1 $Y=1.865 $X2=1
+ $Y2=2.195
r44 6 12 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.55 $Y=1.79
+ $X2=0.385 $Y2=1.715
r45 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=1.79
+ $X2=1 $Y2=1.865
r46 5 6 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.925 $Y=1.79
+ $X2=0.55 $Y2=1.79
r47 3 11 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.475 $Y=0.485
+ $X2=0.475 $Y2=0.975
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%A_27_55# 1 2 9 10 11 12 14 15 17 18 20 22 23
+ 26 30 32 33 36 41 42 45
c79 22 0 1.27692e-19 $X=0.925 $Y=0.805
r80 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=0.97 $X2=0.925 $Y2=0.97
r81 39 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=1.745
+ $X2=0.925 $Y2=1.83
r82 39 41 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.925 $Y=1.745
+ $X2=0.925 $Y2=0.97
r83 38 41 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.925 $Y=0.875
+ $X2=0.925 $Y2=0.97
r84 34 45 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.785 $Y=1.83
+ $X2=0.925 $Y2=1.83
r85 34 36 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=0.785 $Y=1.915
+ $X2=0.785 $Y2=2.13
r86 32 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.84 $Y=0.79
+ $X2=0.925 $Y2=0.875
r87 32 33 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.84 $Y=0.79
+ $X2=0.345 $Y2=0.79
r88 28 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.25 $Y=0.705
+ $X2=0.345 $Y2=0.79
r89 28 30 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=0.25 $Y=0.705
+ $X2=0.25 $Y2=0.55
r90 24 26 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.36 $Y=1.8 $X2=1.46
+ $Y2=1.8
r91 23 42 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.925 $Y=1.325
+ $X2=0.925 $Y2=0.97
r92 22 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=0.805
+ $X2=0.925 $Y2=0.97
r93 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.54 $Y=0.255
+ $X2=1.54 $Y2=0.575
r94 15 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.46 $Y=1.875
+ $X2=1.46 $Y2=1.8
r95 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.46 $Y=1.875
+ $X2=1.46 $Y2=2.195
r96 14 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.36 $Y=1.725
+ $X2=1.36 $Y2=1.8
r97 13 14 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.36 $Y=1.475
+ $X2=1.36 $Y2=1.725
r98 12 23 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.09 $Y=1.4
+ $X2=0.925 $Y2=1.325
r99 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.285 $Y=1.4
+ $X2=1.36 $Y2=1.475
r100 11 12 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.285 $Y=1.4
+ $X2=1.09 $Y2=1.4
r101 9 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.465 $Y=0.18
+ $X2=1.54 $Y2=0.255
r102 9 10 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.465 $Y=0.18
+ $X2=1.09 $Y2=0.18
r103 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.015 $Y=0.255
+ $X2=1.09 $Y2=0.18
r104 7 22 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.015 $Y=0.255
+ $X2=1.015 $Y2=0.805
r105 2 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.985 $X2=0.785 $Y2=2.13
r106 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.275 $X2=0.26 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%B 3 7 9 10 11 16
c34 9 0 1.27692e-19 $X=1.68 $Y=0.555
r35 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.32
+ $X2=1.81 $Y2=1.485
r36 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.32
+ $X2=1.81 $Y2=1.155
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.32 $X2=1.81 $Y2=1.32
r38 11 17 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=1.745 $Y=1.295
+ $X2=1.745 $Y2=1.32
r39 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.745 $Y=0.925
+ $X2=1.745 $Y2=1.295
r40 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.745 $Y=0.555
+ $X2=1.745 $Y2=0.925
r41 7 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.9 $Y=2.195 $X2=1.9
+ $Y2=1.485
r42 3 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.9 $Y=0.575 $X2=1.9
+ $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%C 3 6 9 10 11 12 13 14 19
c38 9 0 5.41121e-20 $X=2.35 $Y=0.895
r39 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.35
+ $Y=1.06 $X2=2.35 $Y2=1.06
r40 14 20 7.52289 $w=3.58e-07 $l=2.35e-07 $layer=LI1_cond $X=2.255 $Y=1.295
+ $X2=2.255 $Y2=1.06
r41 13 20 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=2.255 $Y=0.925
+ $X2=2.255 $Y2=1.06
r42 12 13 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.255 $Y=0.555
+ $X2=2.255 $Y2=0.925
r43 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.35 $Y=1.4 $X2=2.35
+ $Y2=1.06
r44 10 11 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.4
+ $X2=2.35 $Y2=1.565
r45 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=0.895
+ $X2=2.35 $Y2=1.06
r46 6 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.345 $Y=2.195
+ $X2=2.345 $Y2=1.565
r47 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.26 $Y=0.575 $X2=2.26
+ $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%D 3 6 9 10 11 12 13 17
c34 12 0 5.41121e-20 $X=3.12 $Y=0.925
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.89
+ $Y=1.06 $X2=2.89 $Y2=1.06
r36 13 18 6.7706 $w=3.98e-07 $l=2.35e-07 $layer=LI1_cond $X=3.005 $Y=1.295
+ $X2=3.005 $Y2=1.06
r37 12 18 3.8895 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=3.005 $Y=0.925
+ $X2=3.005 $Y2=1.06
r38 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.89 $Y=1.4 $X2=2.89
+ $Y2=1.06
r39 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=1.4
+ $X2=2.89 $Y2=1.565
r40 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=0.895
+ $X2=2.89 $Y2=1.06
r41 6 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.8 $Y=2.195 $X2=2.8
+ $Y2=1.565
r42 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.8 $Y=0.575 $X2=2.8
+ $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%A_240_73# 1 2 3 10 14 17 20 24 26 27 29 31
+ 40
r71 38 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.645 $Y=2.94
+ $X2=2.645 $Y2=2.85
r72 29 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=2.94 $X2=2.645 $Y2=2.94
r73 29 31 38.29 $w=2.08e-07 $l=7.25e-07 $layer=LI1_cond $X=2.585 $Y=2.855
+ $X2=2.585 $Y2=2.13
r74 28 31 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.585 $Y=1.915
+ $X2=2.585 $Y2=2.13
r75 26 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.48 $Y=1.83
+ $X2=2.585 $Y2=1.915
r76 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.48 $Y=1.83 $X2=1.78
+ $Y2=1.83
r77 22 27 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.675 $Y=1.83
+ $X2=1.78 $Y2=1.83
r78 22 32 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.675 $Y=1.83
+ $X2=1.315 $Y2=1.83
r79 22 24 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.675 $Y=1.915
+ $X2=1.675 $Y2=2.13
r80 18 32 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=1.745
+ $X2=1.315 $Y2=1.83
r81 18 20 64.5024 $w=1.88e-07 $l=1.105e-06 $layer=LI1_cond $X=1.315 $Y=1.745
+ $X2=1.315 $Y2=0.64
r82 14 17 830.681 $w=1.5e-07 $l=1.62e-06 $layer=POLY_cond $X=3.34 $Y=0.575
+ $X2=3.34 $Y2=2.195
r83 12 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.34 $Y=2.775
+ $X2=3.34 $Y2=2.195
r84 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=2.85
+ $X2=2.645 $Y2=2.85
r85 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.265 $Y=2.85
+ $X2=3.34 $Y2=2.775
r86 10 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.265 $Y=2.85
+ $X2=2.81 $Y2=2.85
r87 3 31 600 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.985 $X2=2.585 $Y2=2.13
r88 2 24 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.985 $X2=1.675 $Y2=2.13
r89 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.365 $X2=1.325 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%VPWR 1 2 3 12 16 20 23 24 25 27 32 42 43 46
+ 49
r46 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r50 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.125 $Y2=3.33
r53 37 39 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 33 46 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.215 $Y2=3.33
r57 33 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.96 $Y=3.33
+ $X2=2.125 $Y2=3.33
r59 32 35 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 30 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 27 46 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.11 $Y=3.33
+ $X2=1.215 $Y2=3.33
r63 27 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.11 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 25 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 25 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 23 39 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=3.095 $Y2=3.33
r68 22 42 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r69 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.2 $Y=3.33
+ $X2=3.095 $Y2=3.33
r70 18 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.095 $Y2=3.33
r71 18 20 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.095 $Y2=2.26
r72 14 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=3.33
r73 14 16 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=2.26
r74 10 46 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=3.245
+ $X2=1.215 $Y2=3.33
r75 10 12 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=1.215 $Y=3.245
+ $X2=1.215 $Y2=2.26
r76 3 20 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.985 $X2=3.095 $Y2=2.26
r77 2 16 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.985 $X2=2.125 $Y2=2.26
r78 1 12 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.985 $X2=1.215 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%X 1 2 7 8 9 10 11 12 13
r9 12 13 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.567 $Y=2.405
+ $X2=3.567 $Y2=2.775
r10 12 34 13.486 $w=2.33e-07 $l=2.75e-07 $layer=LI1_cond $X=3.567 $Y=2.405
+ $X2=3.567 $Y2=2.13
r11 11 34 4.65881 $w=2.33e-07 $l=9.5e-08 $layer=LI1_cond $X=3.567 $Y=2.035
+ $X2=3.567 $Y2=2.13
r12 10 11 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.567 $Y=1.665
+ $X2=3.567 $Y2=2.035
r13 9 10 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.567 $Y=1.295
+ $X2=3.567 $Y2=1.665
r14 8 9 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.567 $Y=0.925
+ $X2=3.567 $Y2=1.295
r15 7 8 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.567 $Y=0.555
+ $X2=3.567 $Y2=0.925
r16 2 34 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.985 $X2=3.555 $Y2=2.13
r17 1 7 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.365 $X2=3.555 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_M%VGND 1 2 9 13 16 17 18 20 33 34 37
r46 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r48 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r49 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r52 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r54 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r55 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r58 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r59 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r61 16 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.64
+ $Y2=0
r62 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=3.015
+ $Y2=0
r63 15 33 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.6
+ $Y2=0
r64 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.015
+ $Y2=0
r65 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0
r66 11 13 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0.51
r67 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r68 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0.42
r69 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.365 $X2=3.015 $Y2=0.51
r70 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.275 $X2=0.69 $Y2=0.42
.ends

