* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_80_21# A3 a_356_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.631e+11p pd=6.41e+06u as=3.843e+11p ps=3.13e+06u
M1001 VGND A2 a_267_47# VNB nshort w=840000u l=150000u
+  ad=8.988e+11p pd=5.5e+06u as=6.174e+11p ps=4.83e+06u
M1002 VPWR a_80_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=9.828e+11p pd=6.6e+06u as=3.339e+11p ps=3.05e+06u
M1003 VGND a_80_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1004 VPWR B1 a_80_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_267_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_267_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.717e+11p pd=3.11e+06u as=0p ps=0u
M1007 a_591_47# B1 a_267_47# VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1008 a_80_21# C1 a_591_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1009 a_80_21# C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_356_367# A2 a_267_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_267_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
