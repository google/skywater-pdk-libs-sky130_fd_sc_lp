* NGSPICE file created from sky130_fd_sc_lp__sdfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 VPWR RESET_B a_229_491# VPB phighvt w=640000u l=150000u
+  ad=2.7924e+12p pd=2.209e+07u as=5.389e+11p ps=5.28e+06u
M1001 a_1406_399# a_1278_529# VGND VNB nshort w=640000u l=150000u
+  ad=3.2785e+11p pd=2.31e+06u as=1.64372e+12p ps=1.392e+07u
M1002 a_2226_127# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 a_1278_529# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1004 VPWR a_1870_127# a_2370_351# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1005 a_1278_529# a_857_367# a_229_491# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1870_127# a_1080_47# a_1406_399# VPB phighvt w=840000u l=150000u
+  ad=2.688e+11p pd=2.43e+06u as=2.352e+11p ps=2.24e+06u
M1007 a_1509_127# a_1406_399# a_1437_127# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1008 a_1437_127# a_857_367# a_1278_529# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1009 VGND RESET_B a_1509_127# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_565_59# D a_229_491# VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.708e+11p ps=3.99e+06u
M1011 VGND a_1870_127# a_2370_351# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 VPWR a_2064_101# a_2022_533# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 VPWR a_1870_127# a_2064_101# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1014 a_562_491# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1015 a_278_59# a_113_63# a_565_59# VNB nshort w=420000u l=150000u
+  ad=2.751e+11p pd=2.99e+06u as=0p ps=0u
M1016 a_1870_127# a_857_367# a_1406_399# VNB nshort w=640000u l=150000u
+  ad=3.662e+11p pd=2.5e+06u as=0p ps=0u
M1017 a_2022_127# a_1080_47# a_1870_127# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1018 a_229_491# D a_562_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1080_47# a_857_367# VGND VNB nshort w=840000u l=150000u
+  ad=3.679e+11p pd=2.7e+06u as=0p ps=0u
M1020 a_1278_529# a_1080_47# a_229_491# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_113_63# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1022 a_1080_47# a_857_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1023 a_857_367# CLK_N VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1024 a_2022_533# a_857_367# a_1870_127# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_2370_351# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1026 a_361_59# SCD a_278_59# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1027 a_1364_529# a_1080_47# a_1278_529# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1028 a_229_491# SCE a_361_59# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_2064_101# a_2022_127# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_2064_101# a_1870_127# a_2226_127# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1031 Q a_2370_351# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1032 a_312_491# a_113_63# a_229_491# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1033 a_2064_101# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND RESET_B a_278_59# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_857_367# CLK_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1036 VPWR a_1406_399# a_1364_529# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR SCD a_312_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1406_399# a_1278_529# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_113_63# SCE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

