* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 VPWR a_1252_451# a_1836_47# VPB phighvt w=640000u l=150000u
+  ad=2.1846e+12p pd=1.806e+07u as=1.696e+11p ps=1.81e+06u
M1001 VPWR RESET_B a_318_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1002 a_318_535# D a_483_78# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.799e+11p ps=1.97e+06u
M1003 VPWR CLK a_27_101# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1004 a_573_535# a_27_101# a_318_535# VNB nshort w=420000u l=150000u
+  ad=2.31e+11p pd=1.94e+06u as=0p ps=0u
M1005 VPWR a_1399_473# a_1357_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_667_535# a_27_101# a_573_535# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.457e+11p ps=2.85e+06u
M1007 a_709_411# a_573_535# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 VPWR a_709_411# a_667_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND CLK a_27_101# VNB nshort w=420000u l=150000u
+  ad=1.3485e+12p pd=1.194e+07u as=1.113e+11p ps=1.37e+06u
M1010 a_573_535# a_196_464# a_318_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_573_535# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1399_125# a_27_101# a_1252_451# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=2.991e+11p ps=2.4e+06u
M1013 VGND a_1252_451# a_1836_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1014 a_883_119# a_709_411# a_811_119# VNB nshort w=420000u l=150000u
+  ad=1.704e+11p pd=1.74e+06u as=8.82e+10p ps=1.26e+06u
M1015 a_1357_535# a_196_464# a_1252_451# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.43e+06u
M1016 VPWR a_1252_451# a_1399_473# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1017 a_709_411# a_573_535# VGND VNB nshort w=640000u l=150000u
+  ad=2.912e+11p pd=2.19e+06u as=0p ps=0u
M1018 a_1399_473# a_1252_451# a_1593_125# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1019 a_196_464# a_27_101# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1020 a_1252_451# a_196_464# a_709_411# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_196_464# a_27_101# VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1022 Q a_1836_47# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1023 a_811_119# a_196_464# a_573_535# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_1399_473# a_1399_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_1836_47# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_318_535# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND RESET_B a_883_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1593_125# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q a_1836_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1030 a_1252_451# a_27_101# a_709_411# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1399_473# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_483_78# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1836_47# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
