* File: sky130_fd_sc_lp__invlp_8.spice
* Created: Fri Aug 28 10:40:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__invlp_8.pex.spice"
.subckt sky130_fd_sc_lp__invlp_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_A_114_53#_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75006.9 A=0.126 P=1.98 MULT=1
MM1004 N_A_114_53#_M1001_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75006.4 A=0.126 P=1.98 MULT=1
MM1011 N_A_114_53#_M1011_d N_A_M1011_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75006
+ A=0.126 P=1.98 MULT=1
MM1013 N_A_114_53#_M1011_d N_A_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75005.6 A=0.126 P=1.98 MULT=1
MM1015 N_A_114_53#_M1015_d N_A_M1015_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75005.1 A=0.126 P=1.98 MULT=1
MM1016 N_A_114_53#_M1015_d N_A_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75004.7 A=0.126 P=1.98 MULT=1
MM1022 N_A_114_53#_M1022_d N_A_M1022_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_A_114_53#_M1022_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1000_d N_A_M1002_g N_A_114_53#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_A_114_53#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1 SB=75003
+ A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1007_d N_A_M1009_g N_A_114_53#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.5
+ SB=75002.6 A=0.126 P=1.98 MULT=1
MM1014 N_Y_M1014_d N_A_M1014_g N_A_114_53#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.9
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1025 N_Y_M1014_d N_A_M1025_g N_A_114_53#_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75005.4
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1026 N_Y_M1026_d N_A_M1026_g N_A_114_53#_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75005.9
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1027 N_Y_M1026_d N_A_M1027_g N_A_114_53#_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75006.4
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1023 N_A_114_53#_M1027_s N_A_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.2394 PD=1.19 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75006.9 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_114_367#_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75006.9 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_114_367#_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.4 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1006_d N_A_M1010_g N_A_114_367#_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1 SB=75006
+ A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g N_A_114_367#_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1020 N_VPWR_M1017_d N_A_M1020_g N_A_114_367#_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_A_114_367#_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.1764 PD=1.68 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1028 N_VPWR_M1021_d N_A_M1028_g N_A_114_367#_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.1764 PD=1.68 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_A_114_367#_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1005_d N_A_M1008_g N_A_114_367#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_A_114_367#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1018 N_Y_M1012_d N_A_M1018_g N_A_114_367#_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.6
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1019_d N_A_M1019_g N_A_114_367#_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1024 N_Y_M1019_d N_A_M1024_g N_A_114_367#_M1024_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.5
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1030 N_Y_M1030_d N_A_M1030_g N_A_114_367#_M1024_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.1764 PD=1.61 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75005.9
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1031 N_Y_M1030_d N_A_M1031_g N_A_114_367#_M1031_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.1764 PD=1.61 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g N_A_114_367#_M1031_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.0319 P=19.85
*
.include "sky130_fd_sc_lp__invlp_8.pxi.spice"
*
.ends
*
*
