* File: sky130_fd_sc_lp__fa_m.pex.spice
* Created: Wed Sep  2 09:53:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FA_M%A_80_241# 1 2 9 13 17 21 23 27 31 35 36 39 40
+ 43
c95 35 0 1.99168e-19 $X=5.45 $Y=1.45
c96 27 0 1.28278e-19 $X=1.635 $Y=0.92
c97 9 0 3.38977e-20 $X=0.475 $Y=2.045
r98 40 46 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.37
+ $X2=0.587 $Y2=1.535
r99 40 45 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.37
+ $X2=0.587 $Y2=1.205
r100 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.37 $X2=0.61 $Y2=1.37
r101 36 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.45 $Y=1.45
+ $X2=5.45 $Y2=1.615
r102 36 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.45 $Y=1.45
+ $X2=5.45 $Y2=1.285
r103 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.45
+ $Y=1.45 $X2=5.45 $Y2=1.45
r104 33 43 4.56482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=1.45
+ $X2=1.635 $Y2=1.45
r105 33 35 238.128 $w=1.68e-07 $l=3.65e-06 $layer=LI1_cond $X=1.8 $Y=1.45
+ $X2=5.45 $Y2=1.45
r106 29 43 1.76929 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=1.535
+ $X2=1.635 $Y2=1.45
r107 29 31 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=1.635 $Y=1.535
+ $X2=1.635 $Y2=1.98
r108 25 43 1.76929 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=1.365
+ $X2=1.635 $Y2=1.45
r109 25 27 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.635 $Y=1.365
+ $X2=1.635 $Y2=0.92
r110 24 39 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.695 $Y=1.45
+ $X2=0.61 $Y2=1.37
r111 23 43 4.56482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=1.45
+ $X2=1.635 $Y2=1.45
r112 23 24 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.47 $Y=1.45
+ $X2=0.695 $Y2=1.45
r113 21 49 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.43 $Y=2.165
+ $X2=5.43 $Y2=1.615
r114 17 48 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.43 $Y=0.805
+ $X2=5.43 $Y2=1.285
r115 13 45 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.63 $Y=0.835
+ $X2=0.63 $Y2=1.205
r116 9 46 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.475 $Y=2.045
+ $X2=0.475 $Y2=1.535
r117 2 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.835 $X2=1.635 $Y2=1.98
r118 1 27 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.625 $X2=1.635 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%B 3 6 9 11 13 14 18 22 26 30 33 34 35 36 39 42
+ 43 46 47 49 54 55 56 62 65 67 72 79
c142 43 0 3.38977e-20 $X=1.415 $Y=2.425
c143 42 0 7.74325e-20 $X=2.135 $Y=2.425
c144 39 0 1.25016e-19 $X=1.25 $Y=2.79
c145 11 0 1.73635e-19 $X=2.945 $Y=1.665
r146 65 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=2.7
+ $X2=3.525 $Y2=2.535
r147 56 79 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=2.805
+ $X2=3.69 $Y2=2.805
r148 56 72 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.525 $Y=2.805
+ $X2=3.5 $Y2=2.805
r149 56 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.525
+ $Y=2.7 $X2=3.525 $Y2=2.7
r150 55 72 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.12 $Y=2.805
+ $X2=3.5 $Y2=2.805
r151 54 55 14.5572 $w=3.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=2.805
+ $X2=3.12 $Y2=2.805
r152 52 54 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=2.805
+ $X2=2.64 $Y2=2.805
r153 49 52 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.22 $Y=2.425
+ $X2=2.22 $Y2=2.805
r154 47 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.35 $Y=2.91
+ $X2=6.35 $Y2=2.745
r155 46 79 173.54 $w=1.68e-07 $l=2.66e-06 $layer=LI1_cond $X=6.35 $Y=2.91
+ $X2=3.69 $Y2=2.91
r156 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.35
+ $Y=2.91 $X2=6.35 $Y2=2.91
r157 42 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=2.425
+ $X2=2.22 $Y2=2.425
r158 42 43 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.135 $Y=2.425
+ $X2=1.415 $Y2=2.425
r159 40 62 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.25 $Y=2.79
+ $X2=1.42 $Y2=2.79
r160 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=2.79 $X2=1.25 $Y2=2.79
r161 37 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=2.51
+ $X2=1.415 $Y2=2.425
r162 37 39 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.25 $Y=2.51
+ $X2=1.25 $Y2=2.79
r163 33 70 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.26 $Y=2.165
+ $X2=6.26 $Y2=2.745
r164 30 33 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=6.26 $Y=0.805
+ $X2=6.26 $Y2=2.165
r165 24 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.14 $Y=1.665
+ $X2=4.14 $Y2=1.59
r166 24 26 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=4.14 $Y=1.665
+ $X2=4.14 $Y2=2.165
r167 20 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.14 $Y=1.515
+ $X2=4.14 $Y2=1.59
r168 20 22 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.14 $Y=1.515
+ $X2=4.14 $Y2=0.805
r169 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=1.59
+ $X2=3.435 $Y2=1.59
r170 18 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.065 $Y=1.59
+ $X2=4.14 $Y2=1.59
r171 18 19 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.065 $Y=1.59
+ $X2=3.51 $Y2=1.59
r172 16 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.435 $Y=1.665
+ $X2=3.435 $Y2=1.59
r173 16 67 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.435 $Y=1.665
+ $X2=3.435 $Y2=2.535
r174 15 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.02 $Y=1.59
+ $X2=2.945 $Y2=1.59
r175 14 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.36 $Y=1.59
+ $X2=3.435 $Y2=1.59
r176 14 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.36 $Y=1.59
+ $X2=3.02 $Y2=1.59
r177 11 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=1.665
+ $X2=2.945 $Y2=1.59
r178 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.945 $Y=1.665
+ $X2=2.945 $Y2=1.985
r179 7 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=1.515
+ $X2=2.945 $Y2=1.59
r180 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.945 $Y=1.515
+ $X2=2.945 $Y2=0.835
r181 3 6 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=1.42 $Y=0.835
+ $X2=1.42 $Y2=2.045
r182 1 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=2.625
+ $X2=1.42 $Y2=2.79
r183 1 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.42 $Y=2.625
+ $X2=1.42 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%CIN 3 6 7 8 11 14 15 19 22 25 26 27 30 31
c75 30 0 1.25016e-19 $X=1.87 $Y=2.9
c76 19 0 1.99168e-19 $X=5.9 $Y=0.805
r77 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.87
+ $Y=2.9 $X2=1.87 $Y2=2.9
r78 27 31 5.83904 $w=3.73e-07 $l=1.9e-07 $layer=LI1_cond $X=1.68 $Y=2.877
+ $X2=1.87 $Y2=2.877
r79 25 30 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.87 $Y=3.075
+ $X2=1.87 $Y2=2.9
r80 24 30 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=2.735
+ $X2=1.87 $Y2=2.9
r81 19 22 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=5.9 $Y=0.805
+ $X2=5.9 $Y2=2.165
r82 17 22 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=5.9 $Y=3.075 $X2=5.9
+ $Y2=2.165
r83 16 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.645 $Y=3.15
+ $X2=4.57 $Y2=3.15
r84 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.825 $Y=3.15
+ $X2=5.9 $Y2=3.075
r85 15 16 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=5.825 $Y=3.15
+ $X2=4.645 $Y2=3.15
r86 11 14 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=4.57 $Y=0.805
+ $X2=4.57 $Y2=2.165
r87 9 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.57 $Y=3.075
+ $X2=4.57 $Y2=3.15
r88 9 14 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.57 $Y=3.075
+ $X2=4.57 $Y2=2.165
r89 8 25 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.035 $Y=3.15
+ $X2=1.87 $Y2=3.075
r90 7 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.495 $Y=3.15
+ $X2=4.57 $Y2=3.15
r91 7 8 1261.4 $w=1.5e-07 $l=2.46e-06 $layer=POLY_cond $X=4.495 $Y=3.15
+ $X2=2.035 $Y2=3.15
r92 6 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.85 $Y=2.045
+ $X2=1.85 $Y2=2.735
r93 3 6 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=1.85 $Y=0.835
+ $X2=1.85 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%A 3 5 7 8 11 16 17 21 23 25 29 31 35 37 38 39
+ 40 44 50
c118 29 0 2.00703e-19 $X=6.62 $Y=0.805
c119 16 0 1.28278e-19 $X=2.36 $Y=0.835
c120 11 0 7.74325e-20 $X=2.28 $Y=2.045
r121 47 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=0.35
+ $X2=2.33 $Y2=0.515
r122 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=0.35 $X2=2.33 $Y2=0.35
r123 44 47 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.33 $Y=0.18
+ $X2=2.33 $Y2=0.35
r124 40 48 7.56934 $w=2.74e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=0.452
+ $X2=2.33 $Y2=0.452
r125 40 50 4.22604 $w=3.75e-07 $l=1.02e-07 $layer=LI1_cond $X=2.16 $Y=0.452
+ $X2=2.058 $Y2=0.452
r126 39 50 11.6166 $w=3.73e-07 $l=3.78e-07 $layer=LI1_cond $X=1.68 $Y=0.452
+ $X2=2.058 $Y2=0.452
r127 38 39 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.452
+ $X2=1.68 $Y2=0.452
r128 33 35 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=2.28 $Y=1.23 $X2=2.36
+ $Y2=1.23
r129 29 31 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=6.62 $Y=0.805
+ $X2=6.62 $Y2=2.165
r130 27 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.62 $Y=0.255
+ $X2=6.62 $Y2=0.805
r131 26 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.075 $Y=0.18 $X2=5
+ $Y2=0.18
r132 25 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.545 $Y=0.18
+ $X2=6.62 $Y2=0.255
r133 25 26 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=6.545 $Y=0.18
+ $X2=5.075 $Y2=0.18
r134 21 23 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=5 $Y=0.805 $X2=5
+ $Y2=2.165
r135 19 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5 $Y=0.255 $X2=5
+ $Y2=0.18
r136 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5 $Y=0.255 $X2=5
+ $Y2=0.805
r137 18 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=0.18
+ $X2=2.33 $Y2=0.18
r138 17 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.925 $Y=0.18 $X2=5
+ $Y2=0.18
r139 17 18 1246.02 $w=1.5e-07 $l=2.43e-06 $layer=POLY_cond $X=4.925 $Y=0.18
+ $X2=2.495 $Y2=0.18
r140 16 49 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.36 $Y=0.835
+ $X2=2.36 $Y2=0.515
r141 14 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.155
+ $X2=2.36 $Y2=1.23
r142 14 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.36 $Y=1.155
+ $X2=2.36 $Y2=0.835
r143 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=1.305
+ $X2=2.28 $Y2=1.23
r144 9 11 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.28 $Y=1.305
+ $X2=2.28 $Y2=2.045
r145 7 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=0.18
+ $X2=2.33 $Y2=0.18
r146 7 8 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=2.165 $Y=0.18
+ $X2=1.135 $Y2=0.18
r147 3 5 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=1.06 $Y=0.835
+ $X2=1.06 $Y2=2.045
r148 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.06 $Y=0.255
+ $X2=1.135 $Y2=0.18
r149 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.06 $Y=0.255
+ $X2=1.06 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%A_1101_119# 1 2 8 11 14 16 17 18 19 29 32 33 35
r58 33 35 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.092 $Y=1.29
+ $X2=7.092 $Y2=1.125
r59 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.07
+ $Y=1.29 $X2=7.07 $Y2=1.29
r60 27 29 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.685 $Y=2.08
+ $X2=5.88 $Y2=2.08
r61 20 24 14.3034 $w=2.9e-07 $l=4.25699e-07 $layer=LI1_cond $X=5.965 $Y=1.21
+ $X2=5.772 $Y2=0.87
r62 19 32 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=1.21
+ $X2=7.07 $Y2=1.21
r63 19 20 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.985 $Y=1.21
+ $X2=5.965 $Y2=1.21
r64 18 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.88 $Y=1.915
+ $X2=5.88 $Y2=2.08
r65 17 20 5.64745 $w=2.9e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.88 $Y=1.295
+ $X2=5.965 $Y2=1.21
r66 17 18 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.88 $Y=1.295
+ $X2=5.88 $Y2=1.915
r67 14 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.205 $Y=2.165
+ $X2=7.205 $Y2=1.795
r68 11 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.05 $Y=0.805
+ $X2=7.05 $Y2=1.125
r69 8 16 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=7.092 $Y=1.608
+ $X2=7.092 $Y2=1.795
r70 7 33 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=7.092 $Y=1.312
+ $X2=7.092 $Y2=1.29
r71 7 8 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=7.092 $Y=1.312
+ $X2=7.092 $Y2=1.608
r72 2 27 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.955 $X2=5.685 $Y2=2.08
r73 1 24 182 $w=1.7e-07 $l=3.5373e-07 $layer=licon1_NDIFF $count=1 $X=5.505
+ $Y=0.595 $X2=5.685 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%COUT 1 2 11 13 14 15 16 17
r12 16 17 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.405
+ $X2=0.25 $Y2=2.775
r13 15 16 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=0.25 $Y=1.98
+ $X2=0.25 $Y2=2.405
r14 14 15 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=1.98
r15 13 14 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r16 8 13 15.7608 $w=1.88e-07 $l=2.7e-07 $layer=LI1_cond $X=0.25 $Y=1.025
+ $X2=0.25 $Y2=1.295
r17 7 11 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.25 $Y=0.86
+ $X2=0.415 $Y2=0.86
r18 7 8 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.25 $Y=0.86 $X2=0.25
+ $Y2=1.025
r19 2 15 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r20 1 11 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.29
+ $Y=0.625 $X2=0.415 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%VPWR 1 2 3 4 5 18 20 22 26 28 31 33 39 41 43 48
+ 49 50 52 65 66 69
c101 66 0 2.58091e-20 $X=7.44 $Y=3.33
r102 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r105 62 63 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 60 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 59 62 344.471 $w=1.68e-07 $l=5.28e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 59 60 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 57 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r110 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 55 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 52 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r114 52 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r115 50 63 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=6.48 $Y2=3.33
r116 50 60 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 48 62 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.83 $Y=3.33
+ $X2=6.48 $Y2=3.33
r118 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=3.33
+ $X2=6.915 $Y2=3.33
r119 47 65 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7 $Y=3.33 $X2=7.44
+ $Y2=3.33
r120 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=3.33 $X2=6.915
+ $Y2=3.33
r121 45 46 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.835 $Y=2.51
+ $X2=6.835 $Y2=2.595
r122 43 45 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.835 $Y=2.23
+ $X2=6.835 $Y2=2.51
r123 39 40 9.56863 $w=2.04e-07 $l=1.6e-07 $layer=LI1_cond $X=3.93 $Y=2.35
+ $X2=3.93 $Y2=2.51
r124 38 39 7.17647 $w=2.04e-07 $l=1.2e-07 $layer=LI1_cond $X=3.93 $Y=2.23
+ $X2=3.93 $Y2=2.35
r125 33 35 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.65 $Y=2.15 $X2=2.65
+ $Y2=2.35
r126 31 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=3.245
+ $X2=6.915 $Y2=3.33
r127 31 46 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.915 $Y=3.245
+ $X2=6.915 $Y2=2.595
r128 29 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.89 $Y=2.51
+ $X2=4.785 $Y2=2.51
r129 28 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=2.51
+ $X2=6.835 $Y2=2.51
r130 28 29 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=6.67 $Y=2.51
+ $X2=4.89 $Y2=2.51
r131 24 41 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.425
+ $X2=4.785 $Y2=2.51
r132 24 26 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=4.785 $Y=2.425
+ $X2=4.785 $Y2=2.23
r133 23 40 1.80669 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.04 $Y=2.51
+ $X2=3.93 $Y2=2.51
r134 22 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.68 $Y=2.51
+ $X2=4.785 $Y2=2.51
r135 22 23 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.68 $Y=2.51
+ $X2=4.04 $Y2=2.51
r136 21 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.35
+ $X2=2.65 $Y2=2.35
r137 20 39 1.80669 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.82 $Y=2.35
+ $X2=3.93 $Y2=2.35
r138 20 21 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=3.82 $Y=2.35
+ $X2=2.815 $Y2=2.35
r139 16 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r140 16 18 39.6371 $w=3.28e-07 $l=1.135e-06 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.11
r141 5 43 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=6.695
+ $Y=1.955 $X2=6.835 $Y2=2.23
r142 4 26 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.955 $X2=4.785 $Y2=2.23
r143 3 38 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=3.8
+ $Y=1.955 $X2=3.925 $Y2=2.23
r144 2 33 600 $w=1.7e-07 $l=4.38349e-07 $layer=licon1_PDIFF $count=1 $X=2.355
+ $Y=1.835 $X2=2.65 $Y2=2.15
r145 1 18 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%A_385_367# 1 2 7 9 14
c21 14 0 1.73635e-19 $X=3.16 $Y=1.8
r22 14 17 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=3.16 $Y=1.8 $X2=3.16
+ $Y2=1.92
r23 9 12 9.50649 $w=2.08e-07 $l=1.8e-07 $layer=LI1_cond $X=2.065 $Y=1.8
+ $X2=2.065 $Y2=1.98
r24 8 9 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.17 $Y=1.8 $X2=2.065
+ $Y2=1.8
r25 7 14 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.055 $Y=1.8 $X2=3.16
+ $Y2=1.8
r26 7 8 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.055 $Y=1.8 $X2=2.17
+ $Y2=1.8
r27 2 17 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.775 $X2=3.16 $Y2=1.92
r28 1 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=1.835 $X2=2.065 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%A_843_391# 1 2 9 11 12 15
r23 13 15 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=5.215 $Y=1.885
+ $X2=5.215 $Y2=2.08
r24 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.11 $Y=1.8
+ $X2=5.215 $Y2=1.885
r25 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.11 $Y=1.8 $X2=4.46
+ $Y2=1.8
r26 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.355 $Y=1.885
+ $X2=4.46 $Y2=1.8
r27 7 9 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=4.355 $Y=1.885
+ $X2=4.355 $Y2=2.08
r28 2 15 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=5.075
+ $Y=1.955 $X2=5.215 $Y2=2.08
r29 1 9 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.215
+ $Y=1.955 $X2=4.355 $Y2=2.08
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%SUM 1 2 10 13 14 15 16 17
c14 10 0 1.74894e-19 $X=7.43 $Y=0.84
r15 16 17 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.43 $Y=2.405
+ $X2=7.43 $Y2=2.775
r16 15 16 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.43 $Y=2.035
+ $X2=7.43 $Y2=2.405
r17 14 15 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.43 $Y=1.665
+ $X2=7.43 $Y2=2.035
r18 13 14 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.43 $Y=1.295
+ $X2=7.43 $Y2=1.665
r19 11 13 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=7.43 $Y=0.945
+ $X2=7.43 $Y2=1.295
r20 10 11 1.31963 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=7.43 $Y=0.84
+ $X2=7.43 $Y2=0.945
r21 8 10 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=0.84
+ $X2=7.43 $Y2=0.84
r22 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.955 $X2=7.42 $Y2=2.1
r23 1 8 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.595 $X2=7.265 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%VGND 1 2 3 4 5 18 21 24 28 32 35 36 40 43 44 46
+ 47 49 50 52 53 54 79 80
r84 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r85 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r86 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r87 74 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r88 73 76 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r89 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r90 71 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r91 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r92 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r93 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r94 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r95 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r96 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r97 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r98 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r99 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r100 54 71 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r101 54 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r102 52 76 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.73 $Y=0 $X2=6.48
+ $Y2=0
r103 52 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.73 $Y=0 $X2=6.825
+ $Y2=0
r104 51 79 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.92 $Y=0 $X2=7.44
+ $Y2=0
r105 51 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.92 $Y=0 $X2=6.825
+ $Y2=0
r106 49 70 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.62 $Y=0 $X2=4.56
+ $Y2=0
r107 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=0 $X2=4.785
+ $Y2=0
r108 48 73 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.95 $Y=0 $X2=5.04
+ $Y2=0
r109 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.95 $Y=0 $X2=4.785
+ $Y2=0
r110 46 67 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.6
+ $Y2=0
r111 46 47 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.925
+ $Y2=0
r112 45 70 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.03 $Y=0 $X2=4.56
+ $Y2=0
r113 45 47 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.03 $Y=0 $X2=3.925
+ $Y2=0
r114 43 64 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.64
+ $Y2=0
r115 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.76
+ $Y2=0
r116 42 67 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=3.6
+ $Y2=0
r117 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.76
+ $Y2=0
r118 38 40 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=2.68 $Y=0.74 $X2=2.76
+ $Y2=0.74
r119 35 57 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.72
+ $Y2=0
r120 35 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.835
+ $Y2=0
r121 34 61 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.2
+ $Y2=0
r122 34 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.835
+ $Y2=0
r123 30 53 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.825 $Y=0.085
+ $X2=6.825 $Y2=0
r124 30 32 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=6.825 $Y=0.085
+ $X2=6.825 $Y2=0.74
r125 26 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=0.085
+ $X2=4.785 $Y2=0
r126 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.785 $Y=0.085
+ $X2=4.785 $Y2=0.72
r127 22 47 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r128 22 24 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.74
r129 21 40 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.76 $Y=0.645 $X2=2.76
+ $Y2=0.74
r130 20 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0
r131 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0.645
r132 16 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.085
+ $X2=0.835 $Y2=0
r133 16 18 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=0.835 $Y=0.085
+ $X2=0.835 $Y2=0.77
r134 5 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.595 $X2=6.835 $Y2=0.74
r135 4 28 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.645
+ $Y=0.595 $X2=4.785 $Y2=0.72
r136 3 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.8
+ $Y=0.595 $X2=3.925 $Y2=0.74
r137 2 38 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.625 $X2=2.68 $Y2=0.75
r138 1 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.705
+ $Y=0.625 $X2=0.845 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%A_385_125# 1 2 7 11 14
r26 14 16 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.145 $Y=0.92
+ $X2=2.145 $Y2=1.1
r27 9 11 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=3.16 $Y=1.015
+ $X2=3.16 $Y2=0.9
r28 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=1.1 $X2=2.145
+ $Y2=1.1
r29 7 9 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.055 $Y=1.1
+ $X2=3.16 $Y2=1.015
r30 7 8 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.055 $Y=1.1 $X2=2.31
+ $Y2=1.1
r31 2 11 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.625 $X2=3.16 $Y2=0.9
r32 1 14 182 $w=1.7e-07 $l=3.89776e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.625 $X2=2.145 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__FA_M%A_843_119# 1 2 9 11 12 15
r18 13 15 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=5.225 $Y=1.005
+ $X2=5.225 $Y2=0.87
r19 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.13 $Y=1.09
+ $X2=5.225 $Y2=1.005
r20 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.13 $Y=1.09 $X2=4.44
+ $Y2=1.09
r21 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.345 $Y=1.005
+ $X2=4.44 $Y2=1.09
r22 7 9 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=4.345 $Y=1.005
+ $X2=4.345 $Y2=0.87
r23 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.075
+ $Y=0.595 $X2=5.215 $Y2=0.87
r24 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.595 $X2=4.355 $Y2=0.87
.ends

