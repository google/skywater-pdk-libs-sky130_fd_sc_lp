* File: sky130_fd_sc_lp__dlxbp_lp2.spice
* Created: Wed Sep  2 09:48:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxbp_lp2.pex.spice"
.subckt sky130_fd_sc_lp__dlxbp_lp2  VNB VPB D GATE VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1011 A_114_57# N_D_M1011_g N_A_27_57#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g A_114_57# VNB NSHORT L=0.15 W=0.42 AD=0.0651
+ AS=0.0441 PD=0.73 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1021 A_278_57# N_GATE_M1021_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0651 PD=0.63 PS=0.73 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_278_409#_M1012_d N_GATE_M1012_g A_278_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_548_55# N_A_278_409#_M1003_g N_A_461_55#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_278_409#_M1020_g A_548_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1006 A_706_55# N_A_27_57#_M1006_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_784_55#_M1007_d N_A_461_55#_M1007_g A_706_55# VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1013 A_886_55# N_A_278_409#_M1013_g N_A_784_55#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_934_29#_M1014_g A_886_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.1764 AS=0.0504 PD=1.26 PS=0.66 NRD=68.568 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1022 A_1162_55# N_A_784_55#_M1022_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1764 PD=0.63 PS=1.26 NRD=14.28 NRS=91.428 M=1 R=2.8 SA=75003.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_934_29#_M1024_d N_A_784_55#_M1024_g A_1162_55# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_1432_57# N_A_934_29#_M1002_g N_Q_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_934_29#_M1025_g A_1432_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_1590_57# N_A_934_29#_M1004_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_1662_57#_M1008_d N_A_934_29#_M1008_g A_1590_57# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_1860_92# N_A_1662_57#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_Q_N_M1017_d N_A_1662_57#_M1017_g A_1860_92# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_D_M1018_g N_A_27_57#_M1018_s VPB PHIGHVT L=0.25 W=1
+ AD=0.24175 AS=0.285 PD=1.59 PS=2.57 NRD=16.7253 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1005 N_A_278_409#_M1005_d N_GATE_M1005_g N_VPWR_M1018_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.24175 PD=2.57 PS=1.59 NRD=0 NRS=16.7253 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1019 N_VPWR_M1019_d N_A_278_409#_M1019_g N_A_461_55#_M1019_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.203625 AS=0.285 PD=1.63 PS=2.57 NRD=29.2742 NRS=0 M=1 R=4
+ SA=125000 SB=125003 A=0.25 P=2.5 MULT=1
MM1027 A_717_393# N_A_27_57#_M1027_g N_VPWR_M1019_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.203625 PD=1.24 PS=1.63 NRD=12.7853 NRS=0 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1009 N_A_784_55#_M1009_d N_A_278_409#_M1009_g A_717_393# VPB PHIGHVT L=0.25
+ W=1 AD=0.2825 AS=0.12 PD=1.565 PS=1.24 NRD=15.7403 NRS=12.7853 M=1 R=4
+ SA=125001 SB=125002 A=0.25 P=2.5 MULT=1
MM1016 A_978_393# N_A_461_55#_M1016_g N_A_784_55#_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.2825 PD=1.32 PS=1.565 NRD=20.6653 NRS=40.3653 M=1 R=4 SA=125002
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_934_29#_M1001_g A_978_393# VPB PHIGHVT L=0.25 W=1
+ AD=0.295 AS=0.16 PD=1.59 PS=1.32 NRD=10.8153 NRS=20.6653 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1023 N_A_934_29#_M1023_d N_A_784_55#_M1023_g N_VPWR_M1001_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.295 PD=2.57 PS=1.59 NRD=0 NRS=50.2153 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1010 N_VPWR_M1010_d N_A_934_29#_M1010_g N_Q_M1010_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1026 N_A_1662_57#_M1026_d N_A_934_29#_M1026_g N_VPWR_M1010_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1028 N_Q_N_M1028_d N_A_1662_57#_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX29_noxref VNB VPB NWDIODE A=20.1386 P=24.93
*
.include "sky130_fd_sc_lp__dlxbp_lp2.pxi.spice"
*
.ends
*
*
