* File: sky130_fd_sc_lp__o211ai_lp.spice
* Created: Fri Aug 28 11:03:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o211ai_lp  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_38_57#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1197 PD=0.86 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_38_57#_M1005_d N_A2_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 A_329_57# N_B1_M1001_g N_A_38_57#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_C1_M1002_g A_329_57# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 A_137_409# N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1003 N_Y_M1003_d N_A2_M1003_g A_137_409# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.12 PD=1.32 PS=1.24 NRD=7.8603 NRS=12.7853 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_Y_M1003_d VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.16 PD=1.32 PS=1.32 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1000 N_Y_M1000_d N_C1_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=7.8603 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__o211ai_lp.pxi.spice"
*
.ends
*
*
