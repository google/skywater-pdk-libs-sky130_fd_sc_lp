* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or3b_2 A B C_N VGND VNB VPB VPWR X
X0 VPWR a_195_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_33_131# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_33_131# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 X a_195_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_195_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_195_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_448_385# B a_520_385# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_520_385# a_33_131# a_195_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_33_131# a_195_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND A a_195_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_195_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR A a_448_385# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
